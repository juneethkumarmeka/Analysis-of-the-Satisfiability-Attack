module basic_3000_30000_3500_15_levels_10xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
and U0 (N_0,In_2796,In_88);
nand U1 (N_1,In_1798,In_1074);
and U2 (N_2,In_2405,In_860);
xor U3 (N_3,In_2137,In_1511);
or U4 (N_4,In_1280,In_277);
nand U5 (N_5,In_763,In_1766);
xnor U6 (N_6,In_1556,In_703);
nand U7 (N_7,In_2719,In_202);
nand U8 (N_8,In_2615,In_2426);
xnor U9 (N_9,In_1481,In_1000);
or U10 (N_10,In_1252,In_2202);
xor U11 (N_11,In_1056,In_2253);
nor U12 (N_12,In_1985,In_1097);
nor U13 (N_13,In_2403,In_1599);
xnor U14 (N_14,In_2538,In_2156);
or U15 (N_15,In_1760,In_2204);
nand U16 (N_16,In_2490,In_1306);
or U17 (N_17,In_2820,In_262);
nor U18 (N_18,In_305,In_2610);
and U19 (N_19,In_2114,In_832);
xnor U20 (N_20,In_1976,In_2513);
and U21 (N_21,In_760,In_2386);
nand U22 (N_22,In_304,In_2505);
xor U23 (N_23,In_2563,In_359);
or U24 (N_24,In_1064,In_2678);
xnor U25 (N_25,In_996,In_292);
xor U26 (N_26,In_2762,In_1674);
nand U27 (N_27,In_1992,In_961);
nand U28 (N_28,In_1523,In_389);
nand U29 (N_29,In_81,In_510);
or U30 (N_30,In_1112,In_932);
and U31 (N_31,In_1486,In_1989);
and U32 (N_32,In_607,In_853);
nor U33 (N_33,In_1968,In_2173);
and U34 (N_34,In_999,In_1089);
nand U35 (N_35,In_2718,In_2457);
xnor U36 (N_36,In_784,In_1507);
xor U37 (N_37,In_1452,In_361);
and U38 (N_38,In_1218,In_1355);
or U39 (N_39,In_501,In_185);
nor U40 (N_40,In_1585,In_1349);
xnor U41 (N_41,In_2412,In_2266);
nand U42 (N_42,In_274,In_275);
nand U43 (N_43,In_683,In_1963);
or U44 (N_44,In_1971,In_2811);
nor U45 (N_45,In_2010,In_32);
xor U46 (N_46,In_1126,In_851);
nand U47 (N_47,In_1838,In_2948);
xnor U48 (N_48,In_933,In_689);
xnor U49 (N_49,In_576,In_1625);
or U50 (N_50,In_1623,In_2933);
nor U51 (N_51,In_2081,In_2486);
nand U52 (N_52,In_2641,In_1878);
or U53 (N_53,In_72,In_645);
or U54 (N_54,In_1849,In_2371);
and U55 (N_55,In_236,In_1258);
nand U56 (N_56,In_1909,In_138);
or U57 (N_57,In_2712,In_634);
nand U58 (N_58,In_556,In_1151);
or U59 (N_59,In_2668,In_1794);
nor U60 (N_60,In_690,In_1464);
and U61 (N_61,In_2778,In_1865);
xnor U62 (N_62,In_1844,In_2982);
nor U63 (N_63,In_1808,In_1758);
and U64 (N_64,In_858,In_400);
or U65 (N_65,In_1288,In_1113);
nand U66 (N_66,In_2182,In_987);
or U67 (N_67,In_499,In_707);
nor U68 (N_68,In_2663,In_1608);
and U69 (N_69,In_699,In_1604);
or U70 (N_70,In_2991,In_883);
nand U71 (N_71,In_2210,In_931);
or U72 (N_72,In_1465,In_2223);
xnor U73 (N_73,In_412,In_1555);
xnor U74 (N_74,In_313,In_2746);
xnor U75 (N_75,In_11,In_2675);
xnor U76 (N_76,In_2591,In_272);
nand U77 (N_77,In_2042,In_840);
or U78 (N_78,In_696,In_2877);
and U79 (N_79,In_2738,In_1006);
nor U80 (N_80,In_158,In_1517);
nor U81 (N_81,In_2344,In_2469);
nand U82 (N_82,In_887,In_2485);
nand U83 (N_83,In_2111,In_1477);
nor U84 (N_84,In_1207,In_943);
xnor U85 (N_85,In_727,In_1630);
and U86 (N_86,In_925,In_793);
xnor U87 (N_87,In_546,In_1803);
and U88 (N_88,In_2879,In_2364);
nor U89 (N_89,In_823,In_1330);
xnor U90 (N_90,In_1539,In_2704);
or U91 (N_91,In_1160,In_415);
or U92 (N_92,In_1718,In_44);
or U93 (N_93,In_929,In_2925);
nor U94 (N_94,In_1594,In_190);
nor U95 (N_95,In_2914,In_1079);
or U96 (N_96,In_2556,In_698);
and U97 (N_97,In_2453,In_2191);
and U98 (N_98,In_263,In_2074);
nand U99 (N_99,In_801,In_1809);
or U100 (N_100,In_1129,In_2450);
nor U101 (N_101,In_2614,In_1924);
nor U102 (N_102,In_1364,In_568);
and U103 (N_103,In_1712,In_579);
and U104 (N_104,In_2440,In_1372);
or U105 (N_105,In_284,In_43);
nand U106 (N_106,In_1225,In_2909);
xor U107 (N_107,In_2126,In_1051);
nand U108 (N_108,In_1281,In_1236);
and U109 (N_109,In_124,In_162);
and U110 (N_110,In_24,In_533);
and U111 (N_111,In_1916,In_1810);
xnor U112 (N_112,In_928,In_2783);
nand U113 (N_113,In_19,In_2262);
xnor U114 (N_114,In_592,In_2656);
nand U115 (N_115,In_759,In_1036);
or U116 (N_116,In_895,In_635);
or U117 (N_117,In_1859,In_1341);
nor U118 (N_118,In_718,In_746);
or U119 (N_119,In_2826,In_2727);
and U120 (N_120,In_2441,In_939);
xor U121 (N_121,In_2587,In_2922);
nor U122 (N_122,In_2154,In_2978);
xnor U123 (N_123,In_256,In_1133);
xor U124 (N_124,In_136,In_2955);
nand U125 (N_125,In_2717,In_1125);
nand U126 (N_126,In_289,In_2072);
nor U127 (N_127,In_1842,In_2789);
and U128 (N_128,In_658,In_1884);
or U129 (N_129,In_49,In_1209);
nor U130 (N_130,In_729,In_1607);
nor U131 (N_131,In_2268,In_1614);
nor U132 (N_132,In_1731,In_2546);
and U133 (N_133,In_564,In_2157);
or U134 (N_134,In_994,In_2047);
nand U135 (N_135,In_2056,In_1186);
nand U136 (N_136,In_2821,In_156);
xnor U137 (N_137,In_2708,In_2819);
xor U138 (N_138,In_80,In_435);
nand U139 (N_139,In_2448,In_2121);
xnor U140 (N_140,In_1374,In_1531);
nor U141 (N_141,In_1118,In_1804);
or U142 (N_142,In_524,In_672);
xnor U143 (N_143,In_1384,In_1152);
nor U144 (N_144,In_2572,In_2217);
and U145 (N_145,In_2996,In_721);
nand U146 (N_146,In_2912,In_845);
nor U147 (N_147,In_2264,In_2805);
nor U148 (N_148,In_573,In_100);
or U149 (N_149,In_2644,In_2999);
xor U150 (N_150,In_505,In_173);
and U151 (N_151,In_306,In_2807);
nor U152 (N_152,In_294,In_1580);
and U153 (N_153,In_2054,In_2270);
xnor U154 (N_154,In_2671,In_62);
or U155 (N_155,In_633,In_740);
xor U156 (N_156,In_2929,In_2517);
nor U157 (N_157,In_332,In_1038);
nor U158 (N_158,In_945,In_1296);
nand U159 (N_159,In_1759,In_2152);
nand U160 (N_160,In_90,In_2153);
nor U161 (N_161,In_2176,In_1860);
and U162 (N_162,In_1168,In_103);
nand U163 (N_163,In_1039,In_2093);
nor U164 (N_164,In_2582,In_664);
xnor U165 (N_165,In_150,In_196);
xnor U166 (N_166,In_204,In_1843);
and U167 (N_167,In_2545,In_2129);
nand U168 (N_168,In_2932,In_991);
and U169 (N_169,In_1080,In_1853);
nor U170 (N_170,In_927,In_627);
xnor U171 (N_171,In_1790,In_1744);
nor U172 (N_172,In_2281,In_930);
xor U173 (N_173,In_2541,In_2810);
nor U174 (N_174,In_1220,In_2395);
xnor U175 (N_175,In_270,In_2686);
or U176 (N_176,In_1774,In_2477);
xnor U177 (N_177,In_938,In_2684);
xor U178 (N_178,In_2363,In_2389);
nor U179 (N_179,In_1443,In_349);
and U180 (N_180,In_2761,In_717);
nand U181 (N_181,In_1498,In_1195);
xnor U182 (N_182,In_2941,In_1012);
xnor U183 (N_183,In_1346,In_787);
and U184 (N_184,In_439,In_1504);
nand U185 (N_185,In_2798,In_2903);
and U186 (N_186,In_406,In_1215);
and U187 (N_187,In_2406,In_2532);
nand U188 (N_188,In_364,In_2001);
and U189 (N_189,In_1096,In_2331);
or U190 (N_190,In_1619,In_1387);
and U191 (N_191,In_2215,In_449);
or U192 (N_192,In_382,In_2677);
and U193 (N_193,In_286,In_2327);
nand U194 (N_194,In_2442,In_2588);
nand U195 (N_195,In_668,In_399);
and U196 (N_196,In_1969,In_2526);
and U197 (N_197,In_526,In_1197);
nand U198 (N_198,In_820,In_241);
and U199 (N_199,In_2082,In_497);
nand U200 (N_200,In_2414,In_557);
xnor U201 (N_201,In_86,In_2004);
nand U202 (N_202,In_2425,In_953);
or U203 (N_203,In_2062,In_1738);
nor U204 (N_204,In_813,In_45);
and U205 (N_205,In_575,In_1870);
nor U206 (N_206,In_542,In_583);
xnor U207 (N_207,In_611,In_553);
nand U208 (N_208,In_985,In_488);
or U209 (N_209,In_1568,In_1627);
nor U210 (N_210,In_992,In_747);
xnor U211 (N_211,In_653,In_2889);
nand U212 (N_212,In_1381,In_2236);
xor U213 (N_213,In_2958,In_360);
or U214 (N_214,In_1169,In_50);
nand U215 (N_215,In_2068,In_955);
or U216 (N_216,In_2317,In_500);
and U217 (N_217,In_1073,In_495);
and U218 (N_218,In_530,In_563);
or U219 (N_219,In_2483,In_323);
nor U220 (N_220,In_1240,In_458);
and U221 (N_221,In_1470,In_309);
nand U222 (N_222,In_2979,In_2891);
nor U223 (N_223,In_1796,In_393);
and U224 (N_224,In_2231,In_383);
or U225 (N_225,In_1034,In_2252);
nand U226 (N_226,In_2755,In_551);
and U227 (N_227,In_2136,In_2989);
nand U228 (N_228,In_1973,In_477);
and U229 (N_229,In_1093,In_2737);
xnor U230 (N_230,In_1622,In_520);
or U231 (N_231,In_2051,In_2658);
and U232 (N_232,In_792,In_2860);
nand U233 (N_233,In_937,In_1388);
and U234 (N_234,In_1401,In_1727);
or U235 (N_235,In_1418,In_2906);
nand U236 (N_236,In_1121,In_897);
and U237 (N_237,In_1515,In_252);
nand U238 (N_238,In_1673,In_1065);
xnor U239 (N_239,In_416,In_2435);
xnor U240 (N_240,In_947,In_2333);
and U241 (N_241,In_1597,In_1213);
or U242 (N_242,In_1882,In_321);
nor U243 (N_243,In_2185,In_1565);
or U244 (N_244,In_1845,In_203);
or U245 (N_245,In_129,In_1243);
or U246 (N_246,In_1132,In_2692);
xor U247 (N_247,In_1763,In_1193);
xor U248 (N_248,In_450,In_585);
or U249 (N_249,In_1370,In_914);
or U250 (N_250,In_1104,In_659);
or U251 (N_251,In_334,In_1410);
nand U252 (N_252,In_1869,In_2581);
nand U253 (N_253,In_1660,In_69);
or U254 (N_254,In_1995,In_2823);
nand U255 (N_255,In_2520,In_2649);
or U256 (N_256,In_2276,In_1950);
nand U257 (N_257,In_594,In_1905);
nand U258 (N_258,In_1473,In_215);
and U259 (N_259,In_1017,In_2949);
and U260 (N_260,In_1540,In_2183);
nor U261 (N_261,In_1538,In_1378);
and U262 (N_262,In_2574,In_1183);
xnor U263 (N_263,In_1543,In_2674);
and U264 (N_264,In_258,In_1035);
or U265 (N_265,In_2626,In_1307);
xnor U266 (N_266,In_1230,In_2940);
xor U267 (N_267,In_414,In_2800);
nand U268 (N_268,In_1553,In_1728);
and U269 (N_269,In_351,In_1805);
nand U270 (N_270,In_529,In_598);
and U271 (N_271,In_1695,In_1016);
nor U272 (N_272,In_2928,In_260);
nor U273 (N_273,In_1488,In_2624);
and U274 (N_274,In_259,In_7);
nand U275 (N_275,In_2873,In_1704);
xor U276 (N_276,In_584,In_1491);
and U277 (N_277,In_2035,In_1600);
or U278 (N_278,In_200,In_1211);
xnor U279 (N_279,In_723,In_2709);
nor U280 (N_280,In_2244,In_538);
xnor U281 (N_281,In_1161,In_2196);
nand U282 (N_282,In_1595,In_1566);
nor U283 (N_283,In_1545,In_205);
xor U284 (N_284,In_2080,In_2087);
nand U285 (N_285,In_113,In_2335);
nand U286 (N_286,In_2046,In_2300);
or U287 (N_287,In_2107,In_1899);
or U288 (N_288,In_268,In_1512);
xor U289 (N_289,In_2831,In_622);
nand U290 (N_290,In_1764,In_2464);
nand U291 (N_291,In_1244,In_1835);
and U292 (N_292,In_1455,In_1888);
and U293 (N_293,In_2007,In_2437);
nand U294 (N_294,In_2701,In_1693);
and U295 (N_295,In_806,In_2473);
or U296 (N_296,In_963,In_1255);
nor U297 (N_297,In_2354,In_2599);
xnor U298 (N_298,In_2492,In_2049);
nand U299 (N_299,In_197,In_1544);
nand U300 (N_300,In_394,In_989);
and U301 (N_301,In_2027,In_2870);
xor U302 (N_302,In_2551,In_1533);
and U303 (N_303,In_1049,In_1821);
xnor U304 (N_304,In_1967,In_2697);
and U305 (N_305,In_797,In_261);
or U306 (N_306,In_2954,In_2);
nand U307 (N_307,In_1886,In_713);
nor U308 (N_308,In_1771,In_1925);
nand U309 (N_309,In_971,In_1671);
or U310 (N_310,In_1437,In_397);
and U311 (N_311,In_1044,In_599);
nand U312 (N_312,In_881,In_1047);
or U313 (N_313,In_2659,In_448);
nand U314 (N_314,In_348,In_421);
nor U315 (N_315,In_443,In_1548);
nand U316 (N_316,In_1644,In_1441);
nor U317 (N_317,In_1351,In_1226);
nor U318 (N_318,In_1938,In_974);
or U319 (N_319,In_2288,In_386);
nor U320 (N_320,In_755,In_1714);
xnor U321 (N_321,In_493,In_251);
or U322 (N_322,In_983,In_1628);
xor U323 (N_323,In_2645,In_965);
nand U324 (N_324,In_2060,In_1416);
and U325 (N_325,In_2646,In_2994);
nand U326 (N_326,In_1856,In_1653);
or U327 (N_327,In_2222,In_771);
and U328 (N_328,In_1857,In_2601);
xnor U329 (N_329,In_340,In_1881);
or U330 (N_330,In_2953,In_850);
or U331 (N_331,In_403,In_1454);
xnor U332 (N_332,In_2924,In_151);
nor U333 (N_333,In_977,In_593);
nand U334 (N_334,In_582,In_1075);
and U335 (N_335,In_1270,In_1266);
nand U336 (N_336,In_2085,In_193);
xnor U337 (N_337,In_273,In_1601);
or U338 (N_338,In_2140,In_1534);
nor U339 (N_339,In_405,In_1);
xor U340 (N_340,In_1302,In_436);
and U341 (N_341,In_408,In_1677);
and U342 (N_342,In_1191,In_2420);
nand U343 (N_343,In_2854,In_1633);
xor U344 (N_344,In_997,In_1641);
or U345 (N_345,In_1469,In_1147);
xor U346 (N_346,In_1110,In_1179);
nand U347 (N_347,In_2211,In_46);
nor U348 (N_348,In_2346,In_61);
nand U349 (N_349,In_475,In_1818);
xnor U350 (N_350,In_169,In_2401);
and U351 (N_351,In_917,In_2104);
xor U352 (N_352,In_2297,In_1363);
xnor U353 (N_353,In_1357,In_28);
nor U354 (N_354,In_1689,In_998);
nand U355 (N_355,In_817,In_369);
and U356 (N_356,In_871,In_339);
or U357 (N_357,In_1793,In_2433);
xnor U358 (N_358,In_1423,In_271);
nand U359 (N_359,In_1785,In_2391);
xnor U360 (N_360,In_1020,In_2634);
nand U361 (N_361,In_2181,In_1740);
and U362 (N_362,In_2689,In_2938);
xnor U363 (N_363,In_1516,In_2744);
or U364 (N_364,In_904,In_2206);
xor U365 (N_365,In_1530,In_879);
nor U366 (N_366,In_1509,In_2757);
or U367 (N_367,In_1127,In_726);
and U368 (N_368,In_1022,In_1837);
or U369 (N_369,In_1159,In_1814);
xnor U370 (N_370,In_2964,In_1334);
xnor U371 (N_371,In_1576,In_401);
or U372 (N_372,In_1383,In_206);
and U373 (N_373,In_508,In_2977);
nor U374 (N_374,In_2199,In_1164);
xor U375 (N_375,In_988,In_1956);
nand U376 (N_376,In_765,In_368);
and U377 (N_377,In_1972,In_1977);
xnor U378 (N_378,In_367,In_1405);
xnor U379 (N_379,In_2419,In_1339);
nand U380 (N_380,In_671,In_2372);
nor U381 (N_381,In_410,In_1439);
nor U382 (N_382,In_2228,In_1780);
or U383 (N_383,In_1299,In_2053);
and U384 (N_384,In_374,In_2670);
nor U385 (N_385,In_2775,In_2586);
xnor U386 (N_386,In_2163,In_2250);
and U387 (N_387,In_1048,In_1668);
nor U388 (N_388,In_597,In_1659);
nand U389 (N_389,In_76,In_99);
and U390 (N_390,In_1134,In_852);
and U391 (N_391,In_2748,In_307);
xor U392 (N_392,In_2621,In_1932);
nor U393 (N_393,In_2937,In_528);
nor U394 (N_394,In_1392,In_935);
and U395 (N_395,In_1298,In_1008);
xnor U396 (N_396,In_2462,In_1267);
nor U397 (N_397,In_1715,In_749);
or U398 (N_398,In_473,In_680);
xnor U399 (N_399,In_126,In_2872);
and U400 (N_400,In_745,In_2523);
or U401 (N_401,In_1910,In_2133);
nor U402 (N_402,In_1007,In_2155);
nor U403 (N_403,In_1292,In_637);
nor U404 (N_404,In_1479,In_33);
nand U405 (N_405,In_2455,In_224);
nand U406 (N_406,In_1942,In_1224);
xnor U407 (N_407,In_1250,In_1639);
xor U408 (N_408,In_451,In_1834);
nand U409 (N_409,In_209,In_485);
or U410 (N_410,In_2079,In_1400);
nor U411 (N_411,In_722,In_504);
or U412 (N_412,In_2201,In_1333);
or U413 (N_413,In_2740,In_379);
and U414 (N_414,In_2503,In_291);
nor U415 (N_415,In_467,In_968);
nor U416 (N_416,In_2917,In_1431);
or U417 (N_417,In_1547,In_1058);
nor U418 (N_418,In_2552,In_859);
nand U419 (N_419,In_131,In_882);
or U420 (N_420,In_1792,In_249);
nor U421 (N_421,In_1584,In_2071);
and U422 (N_422,In_666,In_2986);
or U423 (N_423,In_221,In_1993);
nor U424 (N_424,In_1018,In_753);
xnor U425 (N_425,In_1496,In_1260);
nor U426 (N_426,In_381,In_1911);
xor U427 (N_427,In_580,In_384);
nor U428 (N_428,In_1935,In_1107);
and U429 (N_429,In_934,In_1305);
nor U430 (N_430,In_327,In_2562);
nand U431 (N_431,In_1755,In_1440);
and U432 (N_432,In_1786,In_2274);
nand U433 (N_433,In_2257,In_245);
and U434 (N_434,In_2186,In_1912);
nor U435 (N_435,In_949,In_1930);
nor U436 (N_436,In_506,In_461);
xor U437 (N_437,In_1811,In_77);
nand U438 (N_438,In_2690,In_2431);
and U439 (N_439,In_78,In_1246);
nor U440 (N_440,In_350,In_1707);
nor U441 (N_441,In_1365,In_1490);
nand U442 (N_442,In_2801,In_1045);
xor U443 (N_443,In_2939,In_828);
xnor U444 (N_444,In_2065,In_130);
or U445 (N_445,In_2905,In_2487);
nor U446 (N_446,In_2606,In_232);
xnor U447 (N_447,In_1245,In_160);
or U448 (N_448,In_697,In_2827);
nor U449 (N_449,In_1920,In_1124);
xnor U450 (N_450,In_958,In_549);
or U451 (N_451,In_1923,In_1573);
nand U452 (N_452,In_388,In_398);
nand U453 (N_453,In_237,In_2816);
xor U454 (N_454,In_590,In_2897);
xor U455 (N_455,In_2102,In_2305);
xnor U456 (N_456,In_775,In_907);
and U457 (N_457,In_2747,In_1948);
xor U458 (N_458,In_2238,In_1887);
nand U459 (N_459,In_812,In_2983);
nand U460 (N_460,In_2410,In_1228);
nand U461 (N_461,In_842,In_515);
and U462 (N_462,In_378,In_2495);
nor U463 (N_463,In_1889,In_1554);
or U464 (N_464,In_2303,In_1140);
and U465 (N_465,In_2703,In_2184);
and U466 (N_466,In_2549,In_2751);
or U467 (N_467,In_1730,In_180);
or U468 (N_468,In_2661,In_2326);
and U469 (N_469,In_1960,In_2825);
or U470 (N_470,In_2693,In_2162);
nand U471 (N_471,In_975,In_1558);
xnor U472 (N_472,In_2369,In_2749);
or U473 (N_473,In_572,In_27);
xnor U474 (N_474,In_2600,In_1602);
or U475 (N_475,In_700,In_2648);
or U476 (N_476,In_704,In_1749);
and U477 (N_477,In_1596,In_2622);
nand U478 (N_478,In_2030,In_2310);
xnor U479 (N_479,In_391,In_1269);
xnor U480 (N_480,In_1475,In_1907);
nor U481 (N_481,In_854,In_1918);
nand U482 (N_482,In_2390,In_1583);
nor U483 (N_483,In_2997,In_2029);
or U484 (N_484,In_1407,In_1901);
xnor U485 (N_485,In_1389,In_1783);
nor U486 (N_486,In_217,In_2654);
or U487 (N_487,In_6,In_1666);
nor U488 (N_488,In_525,In_1577);
xnor U489 (N_489,In_1522,In_14);
nor U490 (N_490,In_157,In_222);
nand U491 (N_491,In_2566,In_51);
or U492 (N_492,In_380,In_2205);
nor U493 (N_493,In_2839,In_868);
and U494 (N_494,In_287,In_872);
xnor U495 (N_495,In_1332,In_1949);
nand U496 (N_496,In_239,In_2830);
or U497 (N_497,In_324,In_2759);
nand U498 (N_498,In_1753,In_163);
xor U499 (N_499,In_2017,In_818);
and U500 (N_500,In_712,In_293);
or U501 (N_501,In_2164,In_2255);
or U502 (N_502,In_1004,In_780);
nor U503 (N_503,In_40,In_2141);
xnor U504 (N_504,In_2968,In_1954);
or U505 (N_505,In_2285,In_1412);
nand U506 (N_506,In_1521,In_2899);
xnor U507 (N_507,In_899,In_1696);
xor U508 (N_508,In_2491,In_1189);
and U509 (N_509,In_1343,In_1768);
nor U510 (N_510,In_36,In_2314);
nor U511 (N_511,In_396,In_2976);
or U512 (N_512,In_73,In_2845);
or U513 (N_513,In_344,In_1591);
nor U514 (N_514,In_2076,In_1885);
xnor U515 (N_515,In_10,In_869);
nor U516 (N_516,In_2290,In_2033);
or U517 (N_517,In_2479,In_2512);
nand U518 (N_518,In_2221,In_419);
nand U519 (N_519,In_1494,In_2560);
nand U520 (N_520,In_1432,In_1767);
or U521 (N_521,In_2669,In_2868);
or U522 (N_522,In_824,In_654);
or U523 (N_523,In_2832,In_1733);
or U524 (N_524,In_2760,In_164);
and U525 (N_525,In_320,In_2411);
nor U526 (N_526,In_2247,In_2786);
nand U527 (N_527,In_365,In_1836);
or U528 (N_528,In_702,In_2148);
xor U529 (N_529,In_1570,In_1997);
and U530 (N_530,In_95,In_954);
nand U531 (N_531,In_2892,In_1769);
nor U532 (N_532,In_1831,In_827);
and U533 (N_533,In_110,In_923);
nand U534 (N_534,In_1959,In_1552);
or U535 (N_535,In_2880,In_2808);
or U536 (N_536,In_1986,In_1451);
and U537 (N_537,In_1482,In_2275);
xor U538 (N_538,In_1222,In_2734);
and U539 (N_539,In_1114,In_581);
nand U540 (N_540,In_896,In_2874);
or U541 (N_541,In_1829,In_2110);
nor U542 (N_542,In_660,In_1647);
or U543 (N_543,In_2643,In_2000);
xor U544 (N_544,In_1770,In_2066);
and U545 (N_545,In_2251,In_1291);
nand U546 (N_546,In_681,In_950);
xor U547 (N_547,In_808,In_1024);
nor U548 (N_548,In_316,In_1615);
nor U549 (N_549,In_2396,In_2192);
nand U550 (N_550,In_1902,In_541);
nor U551 (N_551,In_2197,In_2788);
nand U552 (N_552,In_59,In_464);
and U553 (N_553,In_1679,In_2028);
xor U554 (N_554,In_519,In_1166);
nand U555 (N_555,In_695,In_1979);
or U556 (N_556,In_1264,In_1640);
nand U557 (N_557,In_1561,In_632);
nor U558 (N_558,In_770,In_839);
nor U559 (N_559,In_425,In_905);
or U560 (N_560,In_1171,In_679);
nand U561 (N_561,In_547,In_1756);
nor U562 (N_562,In_2097,In_2966);
nand U563 (N_563,In_822,In_2888);
xor U564 (N_564,In_2394,In_87);
nor U565 (N_565,In_1157,In_385);
or U566 (N_566,In_1311,In_1812);
nor U567 (N_567,In_2213,In_144);
nand U568 (N_568,In_2857,In_2302);
nand U569 (N_569,In_1485,In_2263);
nor U570 (N_570,In_107,In_2226);
or U571 (N_571,In_2752,In_764);
and U572 (N_572,In_518,In_798);
nor U573 (N_573,In_816,In_2119);
and U574 (N_574,In_1342,In_1867);
and U575 (N_575,In_2910,In_1459);
nor U576 (N_576,In_1026,In_1719);
nor U577 (N_577,In_1943,In_2018);
xor U578 (N_578,In_329,In_642);
nor U579 (N_579,In_1221,In_1210);
nor U580 (N_580,In_1646,In_498);
and U581 (N_581,In_1550,In_1415);
nor U582 (N_582,In_650,In_1077);
and U583 (N_583,In_2267,In_213);
and U584 (N_584,In_1356,In_1088);
nand U585 (N_585,In_2856,In_2584);
nor U586 (N_586,In_2842,In_1314);
nor U587 (N_587,In_1433,In_2355);
xor U588 (N_588,In_874,In_1068);
or U589 (N_589,In_1419,In_417);
xnor U590 (N_590,In_4,In_2973);
or U591 (N_591,In_34,In_2175);
nand U592 (N_592,In_2299,In_2324);
nand U593 (N_593,In_2320,In_2935);
or U594 (N_594,In_1537,In_856);
nand U595 (N_595,In_1994,In_2402);
xnor U596 (N_596,In_1503,In_1564);
nand U597 (N_597,In_1456,In_1046);
nor U598 (N_598,In_1717,In_2232);
or U599 (N_599,In_1434,In_1385);
nor U600 (N_600,In_1176,In_2043);
and U601 (N_601,In_2992,In_670);
or U602 (N_602,In_31,In_1656);
nor U603 (N_603,In_1892,In_1621);
or U604 (N_604,In_377,In_978);
nand U605 (N_605,In_2040,In_571);
nor U606 (N_606,In_2515,In_684);
nand U607 (N_607,In_2777,In_2635);
xnor U608 (N_608,In_12,In_1527);
nor U609 (N_609,In_1069,In_2044);
or U610 (N_610,In_1137,In_1941);
xor U611 (N_611,In_2048,In_1864);
and U612 (N_612,In_1706,In_2679);
or U613 (N_613,In_2459,In_2397);
xor U614 (N_614,In_2174,In_1202);
xor U615 (N_615,In_266,In_687);
nor U616 (N_616,In_1216,In_815);
and U617 (N_617,In_1231,In_2430);
nand U618 (N_618,In_1541,In_2618);
nor U619 (N_619,In_208,In_2967);
and U620 (N_620,In_2502,In_302);
nand U621 (N_621,In_1052,In_912);
or U622 (N_622,In_1880,In_1130);
nor U623 (N_623,In_281,In_2585);
xor U624 (N_624,In_2045,In_976);
xor U625 (N_625,In_1263,In_1593);
nor U626 (N_626,In_548,In_478);
or U627 (N_627,In_1120,In_1487);
and U628 (N_628,In_2234,In_2898);
or U629 (N_629,In_2100,In_1807);
and U630 (N_630,In_2179,In_1223);
xnor U631 (N_631,In_783,In_951);
and U632 (N_632,In_1688,In_919);
xor U633 (N_633,In_2779,In_494);
and U634 (N_634,In_876,In_1289);
and U635 (N_635,In_1513,In_231);
and U636 (N_636,In_491,In_2116);
nand U637 (N_637,In_2439,In_2501);
nand U638 (N_638,In_766,In_1376);
nand U639 (N_639,In_1071,In_1832);
or U640 (N_640,In_2714,In_424);
and U641 (N_641,In_2339,In_1198);
and U642 (N_642,In_1395,In_736);
nand U643 (N_643,In_1725,In_1736);
nor U644 (N_644,In_1906,In_1340);
and U645 (N_645,In_288,In_2144);
nor U646 (N_646,In_2529,In_2038);
nor U647 (N_647,In_115,In_2347);
nor U648 (N_648,In_1055,In_1855);
xnor U649 (N_649,In_2200,In_2682);
nor U650 (N_650,In_2286,In_739);
nor U651 (N_651,In_226,In_908);
and U652 (N_652,In_1722,In_2280);
xor U653 (N_653,In_2537,In_94);
nor U654 (N_654,In_186,In_2248);
nand U655 (N_655,In_716,In_849);
xor U656 (N_656,In_890,In_1921);
or U657 (N_657,In_1061,In_29);
nor U658 (N_658,In_1066,In_2094);
nor U659 (N_659,In_1362,In_2423);
nor U660 (N_660,In_1279,In_982);
or U661 (N_661,In_0,In_1397);
or U662 (N_662,In_2052,In_2328);
or U663 (N_663,In_2518,In_145);
xor U664 (N_664,In_471,In_315);
or U665 (N_665,In_2672,In_2258);
nor U666 (N_666,In_2417,In_1895);
xnor U667 (N_667,In_1915,In_511);
nor U668 (N_668,In_355,In_629);
xnor U669 (N_669,In_2169,In_407);
nand U670 (N_670,In_47,In_647);
nand U671 (N_671,In_1560,In_1275);
xor U672 (N_672,In_1322,In_1190);
nand U673 (N_673,In_805,In_1840);
or U674 (N_674,In_2313,In_2957);
nand U675 (N_675,In_2595,In_651);
nand U676 (N_676,In_1420,In_814);
or U677 (N_677,In_655,In_2309);
or U678 (N_678,In_1675,In_2160);
and U679 (N_679,In_1303,In_1146);
and U680 (N_680,In_1192,In_2273);
xor U681 (N_681,In_1447,In_2947);
nor U682 (N_682,In_1345,In_490);
xnor U683 (N_683,In_1732,In_432);
or U684 (N_684,In_693,In_9);
or U685 (N_685,In_2316,In_2665);
nor U686 (N_686,In_1360,In_922);
and U687 (N_687,In_120,In_1103);
or U688 (N_688,In_1021,In_2057);
nor U689 (N_689,In_2525,In_174);
nand U690 (N_690,In_1457,In_586);
nor U691 (N_691,In_880,In_1635);
or U692 (N_692,In_2378,In_2329);
xnor U693 (N_693,In_404,In_1824);
and U694 (N_694,In_264,In_1739);
nor U695 (N_695,In_1773,In_1109);
nand U696 (N_696,In_371,In_1449);
nand U697 (N_697,In_2629,In_885);
nand U698 (N_698,In_96,In_314);
nor U699 (N_699,In_146,In_544);
nor U700 (N_700,In_2063,In_2083);
and U701 (N_701,In_480,In_2246);
or U702 (N_702,In_2304,In_2936);
xnor U703 (N_703,In_514,In_2383);
or U704 (N_704,In_1287,In_2229);
and U705 (N_705,In_1002,In_543);
nand U706 (N_706,In_1508,In_2836);
xnor U707 (N_707,In_1238,In_819);
nor U708 (N_708,In_2539,In_2544);
xnor U709 (N_709,In_1700,In_1282);
nor U710 (N_710,In_618,In_2233);
xnor U711 (N_711,In_71,In_522);
and U712 (N_712,In_2887,In_1295);
nor U713 (N_713,In_1027,In_2338);
nor U714 (N_714,In_1970,In_2804);
xnor U715 (N_715,In_1462,In_165);
and U716 (N_716,In_630,In_387);
and U717 (N_717,In_1196,In_921);
xor U718 (N_718,In_1347,In_1315);
and U719 (N_719,In_1891,In_1734);
nor U720 (N_720,In_1526,In_2829);
xor U721 (N_721,In_427,In_2271);
nor U722 (N_722,In_2334,In_1931);
nor U723 (N_723,In_2950,In_2471);
and U724 (N_724,In_1578,In_1106);
and U725 (N_725,In_2489,In_198);
xnor U726 (N_726,In_16,In_2128);
nor U727 (N_727,In_708,In_317);
nor U728 (N_728,In_1698,In_1185);
nand U729 (N_729,In_2866,In_1634);
nand U730 (N_730,In_453,In_1436);
nor U731 (N_731,In_1908,In_149);
xor U732 (N_732,In_1524,In_118);
nand U733 (N_733,In_2059,In_83);
or U734 (N_734,In_2368,In_2969);
or U735 (N_735,In_48,In_1751);
and U736 (N_736,In_1319,In_1682);
or U737 (N_737,In_2195,In_1435);
or U738 (N_738,In_2500,In_2447);
xnor U739 (N_739,In_176,In_466);
and U740 (N_740,In_1546,In_1100);
and U741 (N_741,In_886,In_75);
xor U742 (N_742,In_1964,In_2765);
xor U743 (N_743,In_2177,In_1368);
and U744 (N_744,In_2108,In_2876);
xnor U745 (N_745,In_342,In_1101);
nand U746 (N_746,In_1478,In_1086);
nand U747 (N_747,In_1787,In_429);
nand U748 (N_748,In_250,In_188);
and U749 (N_749,In_1019,In_2294);
and U750 (N_750,In_1138,In_952);
and U751 (N_751,In_2135,In_30);
nor U752 (N_752,In_212,In_1424);
nor U753 (N_753,In_1359,In_1784);
and U754 (N_754,In_2931,In_2833);
nor U755 (N_755,In_2985,In_437);
xor U756 (N_756,In_1371,In_1799);
and U757 (N_757,In_2376,In_159);
and U758 (N_758,In_2847,In_2676);
and U759 (N_759,In_502,In_2178);
nand U760 (N_760,In_1237,In_1861);
and U761 (N_761,In_2564,In_2451);
or U762 (N_762,In_1788,In_2337);
nor U763 (N_763,In_959,In_390);
nand U764 (N_764,In_2429,In_2416);
and U765 (N_765,In_1825,In_2878);
nor U766 (N_766,In_602,In_2428);
nand U767 (N_767,In_444,In_308);
nand U768 (N_768,In_1928,In_2726);
nor U769 (N_769,In_1254,In_1468);
nand U770 (N_770,In_1316,In_2521);
or U771 (N_771,In_1934,In_2741);
or U772 (N_772,In_2636,In_2667);
xor U773 (N_773,In_2806,In_2569);
or U774 (N_774,In_758,In_1324);
nor U775 (N_775,In_1283,In_152);
xnor U776 (N_776,In_535,In_2357);
nand U777 (N_777,In_774,In_238);
nand U778 (N_778,In_1676,In_1830);
nor U779 (N_779,In_2167,In_1241);
nor U780 (N_780,In_248,In_1632);
xnor U781 (N_781,In_1813,In_1119);
nor U782 (N_782,In_2791,In_111);
nand U783 (N_783,In_85,In_2975);
nor U784 (N_784,In_836,In_1284);
or U785 (N_785,In_2466,In_137);
and U786 (N_786,In_625,In_751);
and U787 (N_787,In_1265,In_2332);
xnor U788 (N_788,In_1900,In_2387);
nor U789 (N_789,In_768,In_1257);
nor U790 (N_790,In_1500,In_311);
or U791 (N_791,In_661,In_2103);
or U792 (N_792,In_23,In_1354);
nor U793 (N_793,In_1702,In_2632);
nor U794 (N_794,In_1642,In_2598);
xor U795 (N_795,In_345,In_1380);
and U796 (N_796,In_980,In_1067);
xor U797 (N_797,In_1670,In_2041);
nor U798 (N_798,In_2956,In_619);
nor U799 (N_799,In_559,In_1273);
and U800 (N_800,In_2037,In_2227);
and U801 (N_801,In_2120,In_1858);
nand U802 (N_802,In_1613,In_540);
and U803 (N_803,In_588,In_2336);
nor U804 (N_804,In_2318,In_1806);
or U805 (N_805,In_1369,In_257);
and U806 (N_806,In_2350,In_566);
xnor U807 (N_807,In_1446,In_2550);
and U808 (N_808,In_1678,In_1217);
nand U809 (N_809,In_2578,In_2409);
or U810 (N_810,In_940,In_1054);
xor U811 (N_811,In_2988,In_2476);
xnor U812 (N_812,In_667,In_1610);
nand U813 (N_813,In_846,In_2627);
xnor U814 (N_814,In_143,In_2715);
nor U815 (N_815,In_1060,In_13);
xnor U816 (N_816,In_2261,In_2113);
nand U817 (N_817,In_2013,In_516);
nand U818 (N_818,In_967,In_463);
nor U819 (N_819,In_2240,In_641);
xnor U820 (N_820,In_1586,In_2882);
nand U821 (N_821,In_1782,In_1532);
nor U822 (N_822,In_2852,In_799);
or U823 (N_823,In_26,In_2702);
nor U824 (N_824,In_1876,In_2617);
and U825 (N_825,In_2691,In_2014);
nand U826 (N_826,In_1629,In_829);
and U827 (N_827,In_2034,In_2871);
xor U828 (N_828,In_322,In_2944);
nor U829 (N_829,In_395,In_1329);
nand U830 (N_830,In_714,In_1145);
nor U831 (N_831,In_2086,In_1212);
xor U832 (N_832,In_1833,In_2209);
nor U833 (N_833,In_1111,In_1765);
and U834 (N_834,In_2509,In_2352);
and U835 (N_835,In_1234,In_1274);
nand U836 (N_836,In_1519,In_440);
and U837 (N_837,In_685,In_1181);
xnor U838 (N_838,In_1414,In_2012);
nor U839 (N_839,In_2050,In_861);
nor U840 (N_840,In_2496,In_2132);
nor U841 (N_841,In_2998,In_2282);
nand U842 (N_842,In_2558,In_2952);
or U843 (N_843,In_155,In_70);
nand U844 (N_844,In_1579,In_608);
xnor U845 (N_845,In_2022,In_1875);
nor U846 (N_846,In_2639,In_1598);
and U847 (N_847,In_748,In_866);
or U848 (N_848,In_1499,In_2838);
and U849 (N_849,In_1952,In_375);
nor U850 (N_850,In_2239,In_1795);
xor U851 (N_851,In_358,In_276);
xor U852 (N_852,In_2696,In_646);
xnor U853 (N_853,In_2130,In_1862);
or U854 (N_854,In_1172,In_993);
and U855 (N_855,In_686,In_133);
xnor U856 (N_856,In_2722,In_2292);
nor U857 (N_857,In_2965,In_2099);
and U858 (N_858,In_1493,In_1272);
nor U859 (N_859,In_1214,In_2296);
nor U860 (N_860,In_2117,In_2769);
nor U861 (N_861,In_2602,In_2720);
nor U862 (N_862,In_2444,In_1822);
nor U863 (N_863,In_789,In_1582);
and U864 (N_864,In_648,In_1390);
nor U865 (N_865,In_843,In_1091);
or U866 (N_866,In_878,In_1847);
or U867 (N_867,In_2750,In_1939);
nand U868 (N_868,In_1259,In_915);
nor U869 (N_869,In_181,In_1951);
xnor U870 (N_870,In_2498,In_454);
nand U871 (N_871,In_1729,In_2680);
or U872 (N_872,In_253,In_2571);
and U873 (N_873,In_1413,In_1394);
or U874 (N_874,In_1571,In_235);
xnor U875 (N_875,In_803,In_2031);
nand U876 (N_876,In_626,In_1894);
nor U877 (N_877,In_1476,In_772);
or U878 (N_878,In_225,In_2926);
and U879 (N_879,In_2092,In_2724);
nor U880 (N_880,In_1898,In_172);
nand U881 (N_881,In_2384,In_2923);
nand U882 (N_882,In_2790,In_2377);
or U883 (N_883,In_1846,In_1996);
nand U884 (N_884,In_2449,In_972);
nor U885 (N_885,In_1382,In_1497);
and U886 (N_886,In_1082,In_2025);
nand U887 (N_887,In_2101,In_2647);
and U888 (N_888,In_229,In_191);
nand U889 (N_889,In_777,In_1286);
nand U890 (N_890,In_1762,In_2064);
and U891 (N_891,In_2519,In_1772);
and U892 (N_892,In_1318,In_1603);
xor U893 (N_893,In_117,In_1426);
xor U894 (N_894,In_1699,In_906);
xor U895 (N_895,In_733,In_1775);
nand U896 (N_896,In_1178,In_1663);
xnor U897 (N_897,In_656,In_1940);
or U898 (N_898,In_2468,In_1271);
nor U899 (N_899,In_2036,In_1863);
xor U900 (N_900,In_2124,In_643);
nand U901 (N_901,In_1325,In_657);
xnor U902 (N_902,In_2235,In_1297);
or U903 (N_903,In_2745,In_1205);
nor U904 (N_904,In_1425,In_1852);
and U905 (N_905,In_1685,In_1098);
or U906 (N_906,In_2818,In_639);
and U907 (N_907,In_964,In_300);
nor U908 (N_908,In_1463,In_68);
nand U909 (N_909,In_610,In_2835);
or U910 (N_910,In_2577,In_1823);
nor U911 (N_911,In_844,In_1944);
nor U912 (N_912,In_1966,In_2834);
and U913 (N_913,In_210,In_1495);
nand U914 (N_914,In_2890,In_1742);
or U915 (N_915,In_1800,In_2930);
nor U916 (N_916,In_735,In_2728);
nand U917 (N_917,In_848,In_1386);
nand U918 (N_918,In_1946,In_2754);
and U919 (N_919,In_1877,In_166);
xor U920 (N_920,In_2105,In_2883);
and U921 (N_921,In_920,In_470);
nor U922 (N_922,In_561,In_2407);
and U923 (N_923,In_1711,In_1686);
nand U924 (N_924,In_1510,In_280);
or U925 (N_925,In_677,In_1072);
nand U926 (N_926,In_605,In_1293);
nand U927 (N_927,In_2342,In_2188);
nand U928 (N_928,In_278,In_1200);
nor U929 (N_929,In_179,In_2723);
nand U930 (N_930,In_2172,In_41);
nand U931 (N_931,In_2711,In_1331);
or U932 (N_932,In_2149,In_409);
and U933 (N_933,In_1344,In_1797);
xor U934 (N_934,In_1638,In_1957);
nor U935 (N_935,In_569,In_489);
xor U936 (N_936,In_194,In_1981);
and U937 (N_937,In_153,In_1094);
nor U938 (N_938,In_1664,In_2458);
and U939 (N_939,In_2803,In_2815);
or U940 (N_940,In_558,In_1059);
or U941 (N_941,In_333,In_2542);
and U942 (N_942,In_93,In_725);
and U943 (N_943,In_343,In_192);
or U944 (N_944,In_220,In_2039);
xnor U945 (N_945,In_1321,In_1518);
xnor U946 (N_946,In_2962,In_674);
and U947 (N_947,In_1309,In_1201);
xor U948 (N_948,In_532,In_761);
nor U949 (N_949,In_1023,In_64);
xor U950 (N_950,In_995,In_1165);
nand U951 (N_951,In_513,In_441);
nand U952 (N_952,In_2974,In_1542);
xnor U953 (N_953,In_2139,In_127);
and U954 (N_954,In_123,In_1883);
nand U955 (N_955,In_1396,In_2488);
or U956 (N_956,In_2730,In_2006);
and U957 (N_957,In_2349,In_1162);
and U958 (N_958,In_1980,In_1958);
nand U959 (N_959,In_1697,In_1816);
and U960 (N_960,In_1285,In_195);
or U961 (N_961,In_1148,In_1743);
or U962 (N_962,In_2776,In_2289);
nand U963 (N_963,In_1328,In_1175);
nand U964 (N_964,In_826,In_2472);
or U965 (N_965,In_1745,In_552);
nand U966 (N_966,In_2366,In_1050);
xnor U967 (N_967,In_1590,In_161);
or U968 (N_968,In_2608,In_171);
nor U969 (N_969,In_1820,In_2536);
and U970 (N_970,In_125,In_1815);
and U971 (N_971,In_1789,In_570);
xor U972 (N_972,In_1983,In_199);
xnor U973 (N_973,In_2700,In_1249);
xnor U974 (N_974,In_1326,In_18);
xnor U975 (N_975,In_2091,In_2687);
or U976 (N_976,In_692,In_1277);
nand U977 (N_977,In_187,In_301);
nor U978 (N_978,In_487,In_2002);
xor U979 (N_979,In_2125,In_603);
or U980 (N_980,In_214,In_531);
xnor U981 (N_981,In_1897,In_2088);
nor U982 (N_982,In_830,In_875);
and U983 (N_983,In_2628,In_1551);
or U984 (N_984,In_354,In_644);
or U985 (N_985,In_2158,In_247);
or U986 (N_986,In_108,In_785);
or U987 (N_987,In_2652,In_242);
xor U988 (N_988,In_2568,In_2597);
and U989 (N_989,In_710,In_2095);
and U990 (N_990,In_2146,In_2681);
and U991 (N_991,In_601,In_2846);
nor U992 (N_992,In_1444,In_8);
or U993 (N_993,In_2993,In_2633);
nand U994 (N_994,In_1438,In_1262);
or U995 (N_995,In_1654,In_1350);
and U996 (N_996,In_2408,In_894);
xnor U997 (N_997,In_1428,In_52);
xnor U998 (N_998,In_1204,In_433);
nand U999 (N_999,In_833,In_738);
nor U1000 (N_1000,In_455,In_1645);
nor U1001 (N_1001,In_2707,In_457);
xnor U1002 (N_1002,In_296,In_1651);
nor U1003 (N_1003,In_2920,In_2090);
nor U1004 (N_1004,In_2374,In_1042);
xor U1005 (N_1005,In_2579,In_2138);
nor U1006 (N_1006,In_1631,In_428);
and U1007 (N_1007,In_420,In_2353);
xor U1008 (N_1008,In_565,In_767);
nor U1009 (N_1009,In_2078,In_1575);
and U1010 (N_1010,In_589,In_2494);
and U1011 (N_1011,In_865,In_228);
and U1012 (N_1012,In_1011,In_1251);
nor U1013 (N_1013,In_1399,In_2548);
xor U1014 (N_1014,In_2424,In_2524);
nand U1015 (N_1015,In_2147,In_521);
or U1016 (N_1016,In_2824,In_1502);
nor U1017 (N_1017,In_2853,In_1926);
or U1018 (N_1018,In_1149,In_776);
or U1019 (N_1019,In_2865,In_613);
nor U1020 (N_1020,In_1721,In_1705);
nor U1021 (N_1021,In_2214,In_2864);
nand U1022 (N_1022,In_616,In_2380);
and U1023 (N_1023,In_916,In_299);
nor U1024 (N_1024,In_678,In_1135);
nand U1025 (N_1025,In_577,In_2919);
nor U1026 (N_1026,In_2055,In_2308);
nand U1027 (N_1027,In_550,In_732);
or U1028 (N_1028,In_402,In_2822);
or U1029 (N_1029,In_1665,In_2260);
and U1030 (N_1030,In_1057,In_2341);
or U1031 (N_1031,In_2604,In_1528);
and U1032 (N_1032,In_2540,In_2287);
nand U1033 (N_1033,In_1652,In_2881);
nor U1034 (N_1034,In_731,In_2279);
nor U1035 (N_1035,In_1999,In_474);
nand U1036 (N_1036,In_1988,In_1637);
nor U1037 (N_1037,In_1987,In_1975);
nand U1038 (N_1038,In_154,In_2980);
xnor U1039 (N_1039,In_2650,In_1826);
nand U1040 (N_1040,In_1974,In_2522);
xnor U1041 (N_1041,In_290,In_1649);
or U1042 (N_1042,In_2620,In_1616);
and U1043 (N_1043,In_669,In_1874);
nor U1044 (N_1044,In_2554,In_2736);
or U1045 (N_1045,In_1117,In_1710);
nor U1046 (N_1046,In_2609,In_1317);
nor U1047 (N_1047,In_2203,In_456);
nor U1048 (N_1048,In_2573,In_1187);
or U1049 (N_1049,In_1242,In_2109);
xor U1050 (N_1050,In_2143,In_2886);
nand U1051 (N_1051,In_479,In_170);
nand U1052 (N_1052,In_2946,In_1953);
or U1053 (N_1053,In_2504,In_821);
or U1054 (N_1054,In_2683,In_1460);
xnor U1055 (N_1055,In_121,In_2224);
or U1056 (N_1056,In_2642,In_537);
xor U1057 (N_1057,In_503,In_1965);
and U1058 (N_1058,In_1208,In_1115);
and U1059 (N_1059,In_1802,In_756);
or U1060 (N_1060,In_55,In_754);
xnor U1061 (N_1061,In_2851,In_1030);
and U1062 (N_1062,In_2972,In_484);
nand U1063 (N_1063,In_1105,In_104);
nand U1064 (N_1064,In_1562,In_1662);
nor U1065 (N_1065,In_2166,In_1791);
or U1066 (N_1066,In_884,In_2900);
xnor U1067 (N_1067,In_1612,In_1471);
nor U1068 (N_1068,In_512,In_2699);
nand U1069 (N_1069,In_37,In_2764);
nor U1070 (N_1070,In_790,In_901);
or U1071 (N_1071,In_183,In_54);
xnor U1072 (N_1072,In_867,In_265);
or U1073 (N_1073,In_1690,In_2772);
xor U1074 (N_1074,In_1559,In_705);
nand U1075 (N_1075,In_1962,In_142);
xnor U1076 (N_1076,In_2771,In_2660);
or U1077 (N_1077,In_2907,In_2927);
and U1078 (N_1078,In_2841,In_2553);
or U1079 (N_1079,In_2535,In_335);
nor U1080 (N_1080,In_373,In_132);
or U1081 (N_1081,In_139,In_1501);
or U1082 (N_1082,In_337,In_1839);
nand U1083 (N_1083,In_63,In_2813);
and U1084 (N_1084,In_1092,In_2547);
or U1085 (N_1085,In_1041,In_662);
or U1086 (N_1086,In_1741,In_2123);
xor U1087 (N_1087,In_682,In_2913);
nor U1088 (N_1088,In_545,In_957);
or U1089 (N_1089,In_2561,In_2916);
xor U1090 (N_1090,In_1170,In_423);
or U1091 (N_1091,In_1053,In_2630);
nor U1092 (N_1092,In_469,In_218);
xnor U1093 (N_1093,In_800,In_2514);
or U1094 (N_1094,In_1708,In_2773);
or U1095 (N_1095,In_701,In_2508);
or U1096 (N_1096,In_353,In_2893);
and U1097 (N_1097,In_1040,In_1312);
or U1098 (N_1098,In_312,In_2218);
xnor U1099 (N_1099,In_2970,In_728);
and U1100 (N_1100,In_1361,In_778);
nand U1101 (N_1101,In_2452,In_1484);
xor U1102 (N_1102,In_2445,In_2921);
xnor U1103 (N_1103,In_2662,In_2758);
xor U1104 (N_1104,In_325,In_1828);
nor U1105 (N_1105,In_66,In_2194);
xor U1106 (N_1106,In_3,In_2706);
nand U1107 (N_1107,In_1448,In_2767);
xnor U1108 (N_1108,In_1142,In_1991);
or U1109 (N_1109,In_2655,In_175);
nand U1110 (N_1110,In_1445,In_606);
xor U1111 (N_1111,In_2020,In_2901);
nand U1112 (N_1112,In_2673,In_60);
nand U1113 (N_1113,In_1589,In_2793);
xor U1114 (N_1114,In_1182,In_422);
nand U1115 (N_1115,In_20,In_962);
nor U1116 (N_1116,In_1536,In_857);
or U1117 (N_1117,In_460,In_2307);
nand U1118 (N_1118,In_2145,In_2528);
nand U1119 (N_1119,In_911,In_2283);
and U1120 (N_1120,In_442,In_216);
xnor U1121 (N_1121,In_2067,In_1720);
xor U1122 (N_1122,In_1872,In_1890);
nor U1123 (N_1123,In_57,In_1587);
nor U1124 (N_1124,In_948,In_1403);
xnor U1125 (N_1125,In_2766,In_2474);
nand U1126 (N_1126,In_782,In_53);
xor U1127 (N_1127,In_2705,In_1001);
nand U1128 (N_1128,In_447,In_2446);
nor U1129 (N_1129,In_979,In_2971);
xnor U1130 (N_1130,In_2293,In_2603);
nor U1131 (N_1131,In_459,In_1232);
and U1132 (N_1132,In_2768,In_2325);
and U1133 (N_1133,In_1037,In_2077);
nor U1134 (N_1134,In_2565,In_2651);
xor U1135 (N_1135,In_2859,In_2295);
nand U1136 (N_1136,In_141,In_1871);
or U1137 (N_1137,In_1750,In_1154);
nand U1138 (N_1138,In_1937,In_2306);
and U1139 (N_1139,In_182,In_1854);
xor U1140 (N_1140,In_1879,In_2189);
nor U1141 (N_1141,In_2084,In_2259);
and U1142 (N_1142,In_1005,In_946);
xor U1143 (N_1143,In_1003,In_2422);
xnor U1144 (N_1144,In_2589,In_2475);
xor U1145 (N_1145,In_140,In_89);
nand U1146 (N_1146,In_1492,In_2575);
xnor U1147 (N_1147,In_1373,In_1624);
or U1148 (N_1148,In_1144,In_1483);
nand U1149 (N_1149,In_788,In_285);
nand U1150 (N_1150,In_303,In_168);
and U1151 (N_1151,In_2918,In_1417);
nand U1152 (N_1152,In_2731,In_370);
nand U1153 (N_1153,In_2315,In_363);
nand U1154 (N_1154,In_615,In_1131);
and U1155 (N_1155,In_298,In_574);
nor U1156 (N_1156,In_638,In_1658);
nand U1157 (N_1157,In_2482,In_2089);
or U1158 (N_1158,In_2534,In_189);
nand U1159 (N_1159,In_2207,In_2003);
nand U1160 (N_1160,In_1779,In_1617);
xnor U1161 (N_1161,In_1116,In_411);
nor U1162 (N_1162,In_1514,In_1929);
nor U1163 (N_1163,In_1474,In_114);
xnor U1164 (N_1164,In_1984,In_472);
and U1165 (N_1165,In_2653,In_1726);
xnor U1166 (N_1166,In_2527,In_1636);
nand U1167 (N_1167,In_2781,In_2902);
and U1168 (N_1168,In_1998,In_612);
nor U1169 (N_1169,In_2567,In_888);
or U1170 (N_1170,In_2592,In_2159);
nor U1171 (N_1171,In_1087,In_328);
nor U1172 (N_1172,In_119,In_1694);
or U1173 (N_1173,In_663,In_2345);
xnor U1174 (N_1174,In_1393,In_101);
nor U1175 (N_1175,In_1158,In_1893);
xor U1176 (N_1176,In_709,In_1851);
xnor U1177 (N_1177,In_623,In_219);
or U1178 (N_1178,In_1123,In_1320);
xnor U1179 (N_1179,In_2625,In_873);
and U1180 (N_1180,In_847,In_1927);
xnor U1181 (N_1181,In_903,In_2638);
or U1182 (N_1182,In_2298,In_1480);
or U1183 (N_1183,In_2795,In_554);
and U1184 (N_1184,In_2848,In_2869);
or U1185 (N_1185,In_2379,In_913);
xnor U1186 (N_1186,In_1961,In_2454);
nand U1187 (N_1187,In_1406,In_2005);
nor U1188 (N_1188,In_240,In_614);
nor U1189 (N_1189,In_2242,In_438);
nand U1190 (N_1190,In_2436,In_1421);
and U1191 (N_1191,In_2118,In_2319);
and U1192 (N_1192,In_539,In_1398);
or U1193 (N_1193,In_91,In_1155);
and U1194 (N_1194,In_109,In_631);
or U1195 (N_1195,In_1184,In_1866);
or U1196 (N_1196,In_2301,In_79);
and U1197 (N_1197,In_2510,In_2312);
nor U1198 (N_1198,In_492,In_604);
xnor U1199 (N_1199,In_1626,In_1535);
and U1200 (N_1200,In_595,In_825);
nand U1201 (N_1201,In_1922,In_326);
and U1202 (N_1202,In_2904,In_2356);
or U1203 (N_1203,In_1301,In_773);
xnor U1204 (N_1204,In_483,In_2122);
nor U1205 (N_1205,In_246,In_1310);
nand U1206 (N_1206,In_426,In_838);
xnor U1207 (N_1207,In_1095,In_1801);
nor U1208 (N_1208,In_1352,In_1083);
or U1209 (N_1209,In_1817,In_1163);
nand U1210 (N_1210,In_730,In_990);
and U1211 (N_1211,In_1010,In_864);
xnor U1212 (N_1212,In_67,In_970);
nand U1213 (N_1213,In_1737,In_2142);
nor U1214 (N_1214,In_762,In_2607);
or U1215 (N_1215,In_1102,In_2106);
nor U1216 (N_1216,In_2461,In_2583);
or U1217 (N_1217,In_831,In_567);
nand U1218 (N_1218,In_1409,In_1156);
and U1219 (N_1219,In_621,In_1348);
nor U1220 (N_1220,In_742,In_2792);
xor U1221 (N_1221,In_809,In_2787);
nand U1222 (N_1222,In_640,In_523);
xor U1223 (N_1223,In_2373,In_1025);
and U1224 (N_1224,In_628,In_1990);
nand U1225 (N_1225,In_2688,In_2212);
xnor U1226 (N_1226,In_2943,In_2134);
or U1227 (N_1227,In_1466,In_1043);
xnor U1228 (N_1228,In_1408,In_1335);
or U1229 (N_1229,In_2951,In_2348);
and U1230 (N_1230,In_58,In_2580);
xnor U1231 (N_1231,In_1982,In_184);
nand U1232 (N_1232,In_1701,In_2570);
xnor U1233 (N_1233,In_2637,In_135);
xnor U1234 (N_1234,In_2254,In_1290);
or U1235 (N_1235,In_893,In_2096);
xor U1236 (N_1236,In_2180,In_1684);
nand U1237 (N_1237,In_392,In_2365);
nor U1238 (N_1238,In_1429,In_1122);
nor U1239 (N_1239,In_1850,In_796);
or U1240 (N_1240,In_1261,In_1375);
xor U1241 (N_1241,In_2024,In_2460);
and U1242 (N_1242,In_2151,In_2507);
and U1243 (N_1243,In_112,In_207);
and U1244 (N_1244,In_2995,In_2237);
nor U1245 (N_1245,In_694,In_1581);
nand U1246 (N_1246,In_1919,In_2291);
nand U1247 (N_1247,In_468,In_1761);
nand U1248 (N_1248,In_2388,In_1945);
or U1249 (N_1249,In_2171,In_1143);
nand U1250 (N_1250,In_376,In_1323);
and U1251 (N_1251,In_84,In_2895);
nor U1252 (N_1252,In_960,In_2216);
nor U1253 (N_1253,In_941,In_2467);
xnor U1254 (N_1254,In_609,In_1472);
or U1255 (N_1255,In_944,In_2733);
nand U1256 (N_1256,In_2594,In_918);
xnor U1257 (N_1257,In_1606,In_2543);
and U1258 (N_1258,In_1525,In_233);
and U1259 (N_1259,In_1461,In_2862);
nor U1260 (N_1260,In_2375,In_2415);
nor U1261 (N_1261,In_1028,In_2193);
and U1262 (N_1262,In_1467,In_1203);
nor U1263 (N_1263,In_234,In_2942);
or U1264 (N_1264,In_2061,In_1239);
nand U1265 (N_1265,In_1868,In_1955);
or U1266 (N_1266,In_1248,In_106);
nand U1267 (N_1267,In_1691,In_2098);
or U1268 (N_1268,In_555,In_1735);
and U1269 (N_1269,In_2404,In_1569);
nor U1270 (N_1270,In_1757,In_22);
nor U1271 (N_1271,In_2593,In_673);
and U1272 (N_1272,In_741,In_600);
xor U1273 (N_1273,In_331,In_1778);
nor U1274 (N_1274,In_1070,In_1136);
nand U1275 (N_1275,In_1338,In_1620);
and U1276 (N_1276,In_2321,In_750);
nand U1277 (N_1277,In_2716,In_791);
nand U1278 (N_1278,In_2150,In_909);
nor U1279 (N_1279,In_255,In_318);
nand U1280 (N_1280,In_1650,In_25);
xnor U1281 (N_1281,In_1247,In_1709);
and U1282 (N_1282,In_1752,In_1206);
nor U1283 (N_1283,In_42,In_676);
nor U1284 (N_1284,In_2343,In_2915);
nor U1285 (N_1285,In_2009,In_1703);
and U1286 (N_1286,In_724,In_1167);
or U1287 (N_1287,In_1141,In_2360);
or U1288 (N_1288,In_2695,In_2058);
and U1289 (N_1289,In_2230,In_719);
nor U1290 (N_1290,In_134,In_1657);
or U1291 (N_1291,In_2959,In_2666);
or U1292 (N_1292,In_910,In_2438);
or U1293 (N_1293,In_2616,In_1062);
xor U1294 (N_1294,In_1180,In_2480);
or U1295 (N_1295,In_462,In_1776);
or U1296 (N_1296,In_496,In_1489);
nand U1297 (N_1297,In_2559,In_97);
nand U1298 (N_1298,In_1723,In_2867);
nand U1299 (N_1299,In_1680,In_2187);
nand U1300 (N_1300,In_2362,In_65);
and U1301 (N_1301,In_1873,In_578);
nor U1302 (N_1302,In_1848,In_1746);
nor U1303 (N_1303,In_98,In_1681);
nand U1304 (N_1304,In_711,In_2443);
nand U1305 (N_1305,In_744,In_15);
nand U1306 (N_1306,In_1672,In_56);
nand U1307 (N_1307,In_779,In_1574);
xor U1308 (N_1308,In_2075,In_1358);
nor U1309 (N_1309,In_1411,In_1084);
nor U1310 (N_1310,In_1377,In_1150);
nand U1311 (N_1311,In_2493,In_2269);
or U1312 (N_1312,In_1300,In_1327);
nor U1313 (N_1313,In_900,In_1450);
nor U1314 (N_1314,In_445,In_346);
xor U1315 (N_1315,In_587,In_1278);
xnor U1316 (N_1316,In_691,In_898);
xnor U1317 (N_1317,In_21,In_283);
nand U1318 (N_1318,In_2497,In_39);
xor U1319 (N_1319,In_1014,In_244);
or U1320 (N_1320,In_1529,In_2008);
nor U1321 (N_1321,In_1713,In_752);
or U1322 (N_1322,In_675,In_341);
nor U1323 (N_1323,In_942,In_2023);
and U1324 (N_1324,In_2277,In_319);
nor U1325 (N_1325,In_1430,In_2799);
xor U1326 (N_1326,In_1031,In_2351);
nor U1327 (N_1327,In_2015,In_1336);
nor U1328 (N_1328,In_1353,In_1692);
or U1329 (N_1329,In_1013,In_2190);
nor U1330 (N_1330,In_1913,In_148);
and U1331 (N_1331,In_431,In_2908);
nor U1332 (N_1332,In_617,In_1304);
or U1333 (N_1333,In_38,In_517);
nand U1334 (N_1334,In_1557,In_889);
or U1335 (N_1335,In_243,In_1563);
or U1336 (N_1336,In_841,In_891);
or U1337 (N_1337,In_1549,In_737);
nor U1338 (N_1338,In_1724,In_1936);
xor U1339 (N_1339,In_1669,In_122);
nor U1340 (N_1340,In_507,In_2710);
nor U1341 (N_1341,In_2784,In_902);
nor U1342 (N_1342,In_2619,In_82);
or U1343 (N_1343,In_1667,In_1914);
xor U1344 (N_1344,In_2516,In_2470);
or U1345 (N_1345,In_476,In_167);
and U1346 (N_1346,In_1177,In_2170);
or U1347 (N_1347,In_1904,In_536);
nor U1348 (N_1348,In_2278,In_2698);
nand U1349 (N_1349,In_560,In_2990);
and U1350 (N_1350,In_2812,In_102);
or U1351 (N_1351,In_794,In_562);
and U1352 (N_1352,In_810,In_2713);
nor U1353 (N_1353,In_1505,In_413);
xor U1354 (N_1354,In_1404,In_1747);
nor U1355 (N_1355,In_2725,In_279);
xnor U1356 (N_1356,In_2127,In_2817);
xnor U1357 (N_1357,In_1716,In_1947);
or U1358 (N_1358,In_2945,In_2265);
or U1359 (N_1359,In_807,In_786);
or U1360 (N_1360,In_591,In_2850);
nor U1361 (N_1361,In_2358,In_2605);
and U1362 (N_1362,In_1085,In_2463);
or U1363 (N_1363,In_336,In_2894);
and U1364 (N_1364,In_2241,In_2249);
nor U1365 (N_1365,In_1572,In_743);
and U1366 (N_1366,In_1661,In_1367);
or U1367 (N_1367,In_1032,In_2685);
nor U1368 (N_1368,In_2168,In_2398);
nor U1369 (N_1369,In_1427,In_1520);
and U1370 (N_1370,In_811,In_2657);
and U1371 (N_1371,In_1253,In_2112);
or U1372 (N_1372,In_1567,In_2370);
or U1373 (N_1373,In_649,In_2418);
xnor U1374 (N_1374,In_2785,In_2245);
nand U1375 (N_1375,In_2855,In_509);
xnor U1376 (N_1376,In_2456,In_330);
xnor U1377 (N_1377,In_2732,In_1219);
nand U1378 (N_1378,In_2911,In_1337);
and U1379 (N_1379,In_834,In_2385);
and U1380 (N_1380,In_2011,In_2770);
nand U1381 (N_1381,In_105,In_2330);
xnor U1382 (N_1382,In_2809,In_2763);
nand U1383 (N_1383,In_227,In_362);
nand U1384 (N_1384,In_2961,In_1781);
nor U1385 (N_1385,In_795,In_2478);
and U1386 (N_1386,In_2802,In_2721);
xnor U1387 (N_1387,In_973,In_2272);
or U1388 (N_1388,In_267,In_1827);
nor U1389 (N_1389,In_1308,In_863);
and U1390 (N_1390,In_1933,In_223);
or U1391 (N_1391,In_2465,In_534);
nor U1392 (N_1392,In_2612,In_2576);
nor U1393 (N_1393,In_2381,In_1108);
xor U1394 (N_1394,In_254,In_310);
and U1395 (N_1395,In_92,In_17);
or U1396 (N_1396,In_1506,In_1402);
nor U1397 (N_1397,In_870,In_1090);
nand U1398 (N_1398,In_715,In_486);
xnor U1399 (N_1399,In_1128,In_2797);
xor U1400 (N_1400,In_1029,In_2393);
and U1401 (N_1401,In_1063,In_201);
and U1402 (N_1402,In_147,In_1588);
xnor U1403 (N_1403,In_282,In_1978);
xor U1404 (N_1404,In_2533,In_1754);
nor U1405 (N_1405,In_527,In_2963);
nor U1406 (N_1406,In_734,In_1235);
nor U1407 (N_1407,In_430,In_2219);
or U1408 (N_1408,In_2400,In_2884);
nand U1409 (N_1409,In_2220,In_1081);
nor U1410 (N_1410,In_2782,In_2399);
xnor U1411 (N_1411,In_802,In_418);
or U1412 (N_1412,In_2987,In_2960);
nor U1413 (N_1413,In_2837,In_297);
xnor U1414 (N_1414,In_706,In_2694);
nor U1415 (N_1415,In_2311,In_2323);
and U1416 (N_1416,In_956,In_2596);
nand U1417 (N_1417,In_1643,In_1174);
and U1418 (N_1418,In_1076,In_1687);
xnor U1419 (N_1419,In_652,In_1611);
nor U1420 (N_1420,In_924,In_2753);
xor U1421 (N_1421,In_2026,In_269);
nor U1422 (N_1422,In_2208,In_757);
and U1423 (N_1423,In_178,In_636);
xnor U1424 (N_1424,In_1227,In_2631);
or U1425 (N_1425,In_128,In_347);
xor U1426 (N_1426,In_2555,In_2413);
xor U1427 (N_1427,In_295,In_984);
and U1428 (N_1428,In_837,In_804);
nor U1429 (N_1429,In_1458,In_2640);
and U1430 (N_1430,In_2611,In_2284);
nand U1431 (N_1431,In_1153,In_2743);
and U1432 (N_1432,In_482,In_1903);
nand U1433 (N_1433,In_338,In_1078);
nand U1434 (N_1434,In_1188,In_2530);
and U1435 (N_1435,In_5,In_2774);
nand U1436 (N_1436,In_1276,In_2115);
and U1437 (N_1437,In_2499,In_2828);
nor U1438 (N_1438,In_1592,In_2382);
nand U1439 (N_1439,In_1366,In_2421);
xor U1440 (N_1440,In_1294,In_1379);
nor U1441 (N_1441,In_1896,In_966);
xnor U1442 (N_1442,In_2069,In_877);
or U1443 (N_1443,In_1233,In_1139);
nor U1444 (N_1444,In_1256,In_665);
nor U1445 (N_1445,In_2623,In_2896);
or U1446 (N_1446,In_356,In_1648);
nor U1447 (N_1447,In_688,In_2613);
nand U1448 (N_1448,In_2735,In_781);
nor U1449 (N_1449,In_1015,In_2756);
and U1450 (N_1450,In_1841,In_892);
or U1451 (N_1451,In_769,In_1748);
or U1452 (N_1452,In_2359,In_352);
nand U1453 (N_1453,In_2256,In_2019);
or U1454 (N_1454,In_969,In_986);
and U1455 (N_1455,In_2225,In_624);
xor U1456 (N_1456,In_481,In_2165);
xor U1457 (N_1457,In_2814,In_2511);
nand U1458 (N_1458,In_2739,In_1819);
or U1459 (N_1459,In_2070,In_2794);
and U1460 (N_1460,In_2340,In_1268);
or U1461 (N_1461,In_2885,In_2198);
nand U1462 (N_1462,In_2729,In_230);
nand U1463 (N_1463,In_1229,In_1194);
xnor U1464 (N_1464,In_452,In_116);
and U1465 (N_1465,In_177,In_1391);
nand U1466 (N_1466,In_2863,In_2506);
and U1467 (N_1467,In_2016,In_2590);
nor U1468 (N_1468,In_2432,In_2322);
and U1469 (N_1469,In_372,In_465);
and U1470 (N_1470,In_2849,In_2531);
and U1471 (N_1471,In_1609,In_835);
nor U1472 (N_1472,In_2843,In_35);
or U1473 (N_1473,In_620,In_2161);
xor U1474 (N_1474,In_2032,In_1033);
nor U1475 (N_1475,In_1099,In_2664);
nand U1476 (N_1476,In_936,In_2481);
nand U1477 (N_1477,In_1683,In_2875);
and U1478 (N_1478,In_2427,In_2984);
nor U1479 (N_1479,In_434,In_446);
and U1480 (N_1480,In_1605,In_1009);
xor U1481 (N_1481,In_366,In_2131);
and U1482 (N_1482,In_2484,In_1173);
nand U1483 (N_1483,In_1453,In_2434);
nand U1484 (N_1484,In_2243,In_74);
and U1485 (N_1485,In_2021,In_2934);
xnor U1486 (N_1486,In_1199,In_2742);
nand U1487 (N_1487,In_2367,In_2981);
or U1488 (N_1488,In_2858,In_211);
and U1489 (N_1489,In_2780,In_2557);
nor U1490 (N_1490,In_1655,In_1917);
or U1491 (N_1491,In_2392,In_1777);
nand U1492 (N_1492,In_2840,In_1313);
nand U1493 (N_1493,In_1618,In_720);
nor U1494 (N_1494,In_2361,In_926);
xnor U1495 (N_1495,In_855,In_2861);
nor U1496 (N_1496,In_1442,In_981);
and U1497 (N_1497,In_2844,In_862);
and U1498 (N_1498,In_2073,In_596);
and U1499 (N_1499,In_1422,In_357);
nand U1500 (N_1500,In_689,In_1063);
nor U1501 (N_1501,In_130,In_458);
nor U1502 (N_1502,In_2323,In_1262);
and U1503 (N_1503,In_2187,In_2453);
and U1504 (N_1504,In_137,In_255);
nand U1505 (N_1505,In_2124,In_928);
and U1506 (N_1506,In_1116,In_1278);
nand U1507 (N_1507,In_1859,In_2511);
or U1508 (N_1508,In_2408,In_2406);
or U1509 (N_1509,In_498,In_2300);
or U1510 (N_1510,In_2104,In_1476);
nand U1511 (N_1511,In_974,In_985);
and U1512 (N_1512,In_1287,In_270);
nor U1513 (N_1513,In_2165,In_1771);
and U1514 (N_1514,In_2793,In_493);
nor U1515 (N_1515,In_286,In_2839);
nor U1516 (N_1516,In_2231,In_565);
xor U1517 (N_1517,In_1579,In_143);
or U1518 (N_1518,In_584,In_942);
nand U1519 (N_1519,In_279,In_2794);
xor U1520 (N_1520,In_516,In_1662);
or U1521 (N_1521,In_1671,In_914);
nand U1522 (N_1522,In_1202,In_804);
or U1523 (N_1523,In_548,In_2812);
and U1524 (N_1524,In_2195,In_134);
nand U1525 (N_1525,In_2372,In_2244);
xor U1526 (N_1526,In_497,In_1039);
nand U1527 (N_1527,In_2718,In_212);
or U1528 (N_1528,In_1031,In_2509);
or U1529 (N_1529,In_949,In_953);
xor U1530 (N_1530,In_286,In_676);
and U1531 (N_1531,In_1486,In_1411);
and U1532 (N_1532,In_2262,In_2268);
nand U1533 (N_1533,In_2842,In_1745);
nor U1534 (N_1534,In_1466,In_1770);
or U1535 (N_1535,In_2117,In_2294);
and U1536 (N_1536,In_422,In_1850);
or U1537 (N_1537,In_278,In_1704);
and U1538 (N_1538,In_1601,In_618);
xor U1539 (N_1539,In_2174,In_691);
or U1540 (N_1540,In_1293,In_783);
nand U1541 (N_1541,In_753,In_954);
xor U1542 (N_1542,In_2035,In_1967);
xnor U1543 (N_1543,In_1280,In_2658);
xnor U1544 (N_1544,In_2072,In_2942);
or U1545 (N_1545,In_2061,In_1219);
or U1546 (N_1546,In_1439,In_2100);
or U1547 (N_1547,In_1065,In_859);
and U1548 (N_1548,In_1357,In_1991);
xnor U1549 (N_1549,In_672,In_678);
nor U1550 (N_1550,In_846,In_395);
xnor U1551 (N_1551,In_1799,In_1550);
nand U1552 (N_1552,In_1887,In_2140);
xor U1553 (N_1553,In_395,In_871);
or U1554 (N_1554,In_2045,In_2314);
and U1555 (N_1555,In_1118,In_1465);
xor U1556 (N_1556,In_1939,In_559);
or U1557 (N_1557,In_2328,In_1142);
and U1558 (N_1558,In_1779,In_2243);
and U1559 (N_1559,In_2272,In_2723);
or U1560 (N_1560,In_319,In_2665);
xnor U1561 (N_1561,In_2606,In_959);
and U1562 (N_1562,In_1067,In_801);
nor U1563 (N_1563,In_577,In_1437);
nor U1564 (N_1564,In_2478,In_2087);
xnor U1565 (N_1565,In_2914,In_111);
and U1566 (N_1566,In_2556,In_1930);
and U1567 (N_1567,In_403,In_2588);
xor U1568 (N_1568,In_1449,In_2110);
nor U1569 (N_1569,In_2123,In_1476);
xor U1570 (N_1570,In_2873,In_2234);
and U1571 (N_1571,In_1197,In_955);
and U1572 (N_1572,In_70,In_445);
xor U1573 (N_1573,In_899,In_76);
xor U1574 (N_1574,In_2257,In_68);
nand U1575 (N_1575,In_1518,In_145);
nand U1576 (N_1576,In_2865,In_1538);
and U1577 (N_1577,In_2254,In_2828);
nand U1578 (N_1578,In_1220,In_153);
nand U1579 (N_1579,In_2737,In_896);
or U1580 (N_1580,In_101,In_2710);
nand U1581 (N_1581,In_1887,In_1038);
xnor U1582 (N_1582,In_1190,In_2297);
or U1583 (N_1583,In_2412,In_856);
or U1584 (N_1584,In_317,In_1152);
xor U1585 (N_1585,In_1373,In_256);
nor U1586 (N_1586,In_1269,In_2044);
or U1587 (N_1587,In_1303,In_2390);
nor U1588 (N_1588,In_220,In_2583);
nand U1589 (N_1589,In_2949,In_2883);
and U1590 (N_1590,In_2598,In_1275);
and U1591 (N_1591,In_2487,In_1262);
nor U1592 (N_1592,In_1392,In_940);
xor U1593 (N_1593,In_1740,In_822);
nand U1594 (N_1594,In_1689,In_2190);
and U1595 (N_1595,In_1698,In_682);
xor U1596 (N_1596,In_2557,In_1320);
or U1597 (N_1597,In_2267,In_1808);
xnor U1598 (N_1598,In_762,In_2567);
nand U1599 (N_1599,In_576,In_2798);
xnor U1600 (N_1600,In_2241,In_1425);
nor U1601 (N_1601,In_2649,In_1460);
or U1602 (N_1602,In_906,In_8);
or U1603 (N_1603,In_2597,In_1249);
nand U1604 (N_1604,In_1981,In_1364);
or U1605 (N_1605,In_2104,In_2086);
nor U1606 (N_1606,In_974,In_2663);
nand U1607 (N_1607,In_1819,In_1513);
and U1608 (N_1608,In_163,In_2849);
xor U1609 (N_1609,In_1312,In_1714);
or U1610 (N_1610,In_2528,In_1525);
or U1611 (N_1611,In_38,In_1862);
nand U1612 (N_1612,In_824,In_2010);
nor U1613 (N_1613,In_1604,In_990);
xor U1614 (N_1614,In_444,In_338);
nand U1615 (N_1615,In_2534,In_754);
nand U1616 (N_1616,In_1269,In_2999);
and U1617 (N_1617,In_1209,In_1028);
nand U1618 (N_1618,In_1216,In_1844);
and U1619 (N_1619,In_2759,In_285);
nand U1620 (N_1620,In_974,In_1491);
nand U1621 (N_1621,In_2683,In_574);
xor U1622 (N_1622,In_1425,In_1095);
nor U1623 (N_1623,In_527,In_1915);
or U1624 (N_1624,In_1518,In_1572);
xnor U1625 (N_1625,In_2610,In_2812);
or U1626 (N_1626,In_736,In_413);
xnor U1627 (N_1627,In_1643,In_561);
xor U1628 (N_1628,In_890,In_1086);
nand U1629 (N_1629,In_2737,In_1244);
and U1630 (N_1630,In_129,In_2968);
nand U1631 (N_1631,In_976,In_376);
xor U1632 (N_1632,In_635,In_891);
xnor U1633 (N_1633,In_2752,In_1584);
nor U1634 (N_1634,In_1069,In_1107);
nand U1635 (N_1635,In_27,In_2762);
nor U1636 (N_1636,In_1135,In_1185);
or U1637 (N_1637,In_1193,In_1932);
nand U1638 (N_1638,In_717,In_1029);
and U1639 (N_1639,In_2386,In_1574);
xor U1640 (N_1640,In_193,In_1335);
nand U1641 (N_1641,In_2411,In_2734);
nor U1642 (N_1642,In_2897,In_1491);
or U1643 (N_1643,In_2366,In_1803);
and U1644 (N_1644,In_81,In_1037);
nor U1645 (N_1645,In_1038,In_2943);
or U1646 (N_1646,In_953,In_1801);
and U1647 (N_1647,In_1374,In_1431);
xor U1648 (N_1648,In_2349,In_494);
and U1649 (N_1649,In_2402,In_317);
or U1650 (N_1650,In_906,In_2392);
and U1651 (N_1651,In_2376,In_1670);
nor U1652 (N_1652,In_207,In_2217);
or U1653 (N_1653,In_1722,In_2108);
nor U1654 (N_1654,In_1415,In_1546);
nor U1655 (N_1655,In_1187,In_85);
xor U1656 (N_1656,In_2602,In_2811);
nor U1657 (N_1657,In_54,In_2796);
nor U1658 (N_1658,In_1524,In_2054);
and U1659 (N_1659,In_178,In_508);
nand U1660 (N_1660,In_2522,In_2830);
xnor U1661 (N_1661,In_1010,In_461);
xor U1662 (N_1662,In_2637,In_916);
nand U1663 (N_1663,In_353,In_2972);
and U1664 (N_1664,In_2083,In_1070);
xor U1665 (N_1665,In_1266,In_2296);
xnor U1666 (N_1666,In_2050,In_907);
nor U1667 (N_1667,In_2507,In_1223);
nand U1668 (N_1668,In_155,In_1307);
xor U1669 (N_1669,In_1582,In_2312);
or U1670 (N_1670,In_940,In_1085);
nand U1671 (N_1671,In_1280,In_2953);
nor U1672 (N_1672,In_382,In_2179);
nand U1673 (N_1673,In_616,In_841);
and U1674 (N_1674,In_959,In_1317);
nand U1675 (N_1675,In_1806,In_752);
and U1676 (N_1676,In_411,In_871);
xnor U1677 (N_1677,In_1139,In_1897);
xnor U1678 (N_1678,In_2020,In_731);
and U1679 (N_1679,In_1064,In_1201);
or U1680 (N_1680,In_1937,In_2825);
nor U1681 (N_1681,In_1525,In_2028);
nand U1682 (N_1682,In_2590,In_1681);
nor U1683 (N_1683,In_2141,In_1432);
nor U1684 (N_1684,In_1551,In_1895);
nor U1685 (N_1685,In_1521,In_2661);
and U1686 (N_1686,In_1183,In_1967);
xor U1687 (N_1687,In_2866,In_198);
xor U1688 (N_1688,In_1242,In_1978);
nand U1689 (N_1689,In_2819,In_101);
or U1690 (N_1690,In_1147,In_2178);
nor U1691 (N_1691,In_2166,In_2048);
or U1692 (N_1692,In_239,In_720);
nand U1693 (N_1693,In_847,In_2531);
nand U1694 (N_1694,In_765,In_2178);
xor U1695 (N_1695,In_2245,In_2306);
nand U1696 (N_1696,In_975,In_583);
nand U1697 (N_1697,In_630,In_139);
or U1698 (N_1698,In_2250,In_71);
or U1699 (N_1699,In_2587,In_631);
and U1700 (N_1700,In_2968,In_1803);
xnor U1701 (N_1701,In_2075,In_518);
nand U1702 (N_1702,In_1358,In_2340);
nand U1703 (N_1703,In_1693,In_2248);
nor U1704 (N_1704,In_672,In_2589);
nor U1705 (N_1705,In_1908,In_987);
xor U1706 (N_1706,In_687,In_1398);
and U1707 (N_1707,In_868,In_958);
or U1708 (N_1708,In_2975,In_182);
nand U1709 (N_1709,In_2746,In_1893);
nor U1710 (N_1710,In_74,In_2068);
nor U1711 (N_1711,In_1417,In_1823);
and U1712 (N_1712,In_1964,In_566);
nand U1713 (N_1713,In_1678,In_1494);
or U1714 (N_1714,In_2782,In_2161);
and U1715 (N_1715,In_913,In_1328);
or U1716 (N_1716,In_2555,In_1949);
nand U1717 (N_1717,In_24,In_1359);
nand U1718 (N_1718,In_1847,In_1144);
or U1719 (N_1719,In_1725,In_647);
and U1720 (N_1720,In_1347,In_630);
and U1721 (N_1721,In_1519,In_1439);
nor U1722 (N_1722,In_1257,In_233);
nand U1723 (N_1723,In_799,In_1840);
nand U1724 (N_1724,In_707,In_2345);
nand U1725 (N_1725,In_2259,In_168);
nand U1726 (N_1726,In_2593,In_846);
xnor U1727 (N_1727,In_1118,In_362);
nor U1728 (N_1728,In_304,In_242);
and U1729 (N_1729,In_1456,In_137);
xor U1730 (N_1730,In_2739,In_231);
or U1731 (N_1731,In_2695,In_1808);
nor U1732 (N_1732,In_2794,In_1445);
nor U1733 (N_1733,In_2982,In_2487);
or U1734 (N_1734,In_1665,In_1688);
xnor U1735 (N_1735,In_2741,In_2801);
or U1736 (N_1736,In_2481,In_1592);
nor U1737 (N_1737,In_970,In_839);
xor U1738 (N_1738,In_485,In_2785);
or U1739 (N_1739,In_1921,In_552);
nor U1740 (N_1740,In_1203,In_2132);
xor U1741 (N_1741,In_1185,In_606);
xor U1742 (N_1742,In_1923,In_975);
nor U1743 (N_1743,In_890,In_2000);
nor U1744 (N_1744,In_2510,In_2528);
nand U1745 (N_1745,In_1154,In_1502);
nand U1746 (N_1746,In_2283,In_2733);
xor U1747 (N_1747,In_764,In_1667);
xnor U1748 (N_1748,In_2329,In_2501);
and U1749 (N_1749,In_411,In_757);
or U1750 (N_1750,In_733,In_2204);
nand U1751 (N_1751,In_2721,In_2716);
xnor U1752 (N_1752,In_2144,In_1594);
nand U1753 (N_1753,In_843,In_544);
nand U1754 (N_1754,In_179,In_408);
xnor U1755 (N_1755,In_2905,In_2663);
or U1756 (N_1756,In_2479,In_2761);
or U1757 (N_1757,In_2536,In_2862);
nand U1758 (N_1758,In_990,In_1637);
and U1759 (N_1759,In_1450,In_2810);
nor U1760 (N_1760,In_1707,In_1998);
xor U1761 (N_1761,In_2392,In_1291);
nand U1762 (N_1762,In_2636,In_593);
nor U1763 (N_1763,In_2673,In_963);
nand U1764 (N_1764,In_963,In_292);
xor U1765 (N_1765,In_793,In_2390);
and U1766 (N_1766,In_739,In_2780);
nor U1767 (N_1767,In_2838,In_558);
and U1768 (N_1768,In_1945,In_1808);
and U1769 (N_1769,In_2771,In_2696);
xnor U1770 (N_1770,In_388,In_1915);
or U1771 (N_1771,In_695,In_2514);
nand U1772 (N_1772,In_618,In_2381);
and U1773 (N_1773,In_450,In_1015);
nor U1774 (N_1774,In_1447,In_1894);
xnor U1775 (N_1775,In_2527,In_2982);
or U1776 (N_1776,In_1423,In_2338);
or U1777 (N_1777,In_679,In_554);
nand U1778 (N_1778,In_2158,In_2593);
xnor U1779 (N_1779,In_1547,In_1793);
and U1780 (N_1780,In_1605,In_2906);
and U1781 (N_1781,In_1499,In_1888);
nor U1782 (N_1782,In_2422,In_464);
nand U1783 (N_1783,In_1780,In_738);
or U1784 (N_1784,In_1106,In_1839);
nor U1785 (N_1785,In_2129,In_2794);
and U1786 (N_1786,In_389,In_1479);
and U1787 (N_1787,In_2806,In_1421);
and U1788 (N_1788,In_2786,In_154);
xor U1789 (N_1789,In_620,In_726);
xnor U1790 (N_1790,In_653,In_1278);
or U1791 (N_1791,In_2038,In_1529);
nand U1792 (N_1792,In_1837,In_1428);
or U1793 (N_1793,In_2396,In_1792);
xnor U1794 (N_1794,In_2010,In_1976);
xor U1795 (N_1795,In_668,In_307);
and U1796 (N_1796,In_1763,In_1353);
or U1797 (N_1797,In_1550,In_2518);
or U1798 (N_1798,In_2454,In_273);
nor U1799 (N_1799,In_326,In_2147);
xor U1800 (N_1800,In_1836,In_1346);
nor U1801 (N_1801,In_2142,In_2539);
xnor U1802 (N_1802,In_1309,In_529);
and U1803 (N_1803,In_2312,In_31);
nand U1804 (N_1804,In_391,In_1359);
nand U1805 (N_1805,In_2830,In_144);
and U1806 (N_1806,In_521,In_374);
xnor U1807 (N_1807,In_2341,In_2112);
nand U1808 (N_1808,In_51,In_2959);
xnor U1809 (N_1809,In_2506,In_1402);
nor U1810 (N_1810,In_2185,In_2415);
or U1811 (N_1811,In_657,In_1705);
nand U1812 (N_1812,In_2129,In_2319);
nor U1813 (N_1813,In_2882,In_139);
and U1814 (N_1814,In_814,In_458);
xnor U1815 (N_1815,In_640,In_893);
nand U1816 (N_1816,In_1230,In_1869);
or U1817 (N_1817,In_195,In_160);
xor U1818 (N_1818,In_2832,In_1276);
and U1819 (N_1819,In_1641,In_297);
and U1820 (N_1820,In_1513,In_1066);
nand U1821 (N_1821,In_481,In_2946);
and U1822 (N_1822,In_954,In_2445);
xor U1823 (N_1823,In_1313,In_2203);
or U1824 (N_1824,In_2785,In_2102);
or U1825 (N_1825,In_2549,In_1414);
nor U1826 (N_1826,In_1990,In_1266);
and U1827 (N_1827,In_1402,In_648);
and U1828 (N_1828,In_1908,In_2197);
and U1829 (N_1829,In_2945,In_1781);
nor U1830 (N_1830,In_20,In_459);
or U1831 (N_1831,In_2326,In_1292);
or U1832 (N_1832,In_837,In_2839);
nor U1833 (N_1833,In_2028,In_1038);
nand U1834 (N_1834,In_1636,In_1001);
or U1835 (N_1835,In_1781,In_766);
and U1836 (N_1836,In_2729,In_2073);
and U1837 (N_1837,In_1530,In_518);
and U1838 (N_1838,In_657,In_2632);
nor U1839 (N_1839,In_2556,In_1367);
xnor U1840 (N_1840,In_1938,In_2652);
nand U1841 (N_1841,In_1433,In_735);
nor U1842 (N_1842,In_2541,In_941);
or U1843 (N_1843,In_705,In_1686);
nor U1844 (N_1844,In_379,In_1447);
or U1845 (N_1845,In_225,In_1633);
or U1846 (N_1846,In_321,In_1223);
or U1847 (N_1847,In_1891,In_1782);
or U1848 (N_1848,In_2573,In_2497);
and U1849 (N_1849,In_350,In_599);
xnor U1850 (N_1850,In_1546,In_297);
nand U1851 (N_1851,In_670,In_2038);
or U1852 (N_1852,In_2036,In_2200);
nor U1853 (N_1853,In_1548,In_242);
nor U1854 (N_1854,In_2734,In_1168);
or U1855 (N_1855,In_741,In_1512);
nand U1856 (N_1856,In_1160,In_2905);
and U1857 (N_1857,In_1486,In_728);
or U1858 (N_1858,In_462,In_2288);
nor U1859 (N_1859,In_118,In_2246);
nor U1860 (N_1860,In_1828,In_1936);
xnor U1861 (N_1861,In_2401,In_669);
nor U1862 (N_1862,In_1347,In_1038);
nor U1863 (N_1863,In_794,In_1304);
and U1864 (N_1864,In_653,In_475);
nor U1865 (N_1865,In_931,In_1546);
xor U1866 (N_1866,In_1677,In_107);
nor U1867 (N_1867,In_1214,In_1029);
and U1868 (N_1868,In_1224,In_1517);
xnor U1869 (N_1869,In_2417,In_2798);
nor U1870 (N_1870,In_404,In_1466);
or U1871 (N_1871,In_200,In_1950);
or U1872 (N_1872,In_2299,In_851);
nand U1873 (N_1873,In_2105,In_2514);
xor U1874 (N_1874,In_1262,In_1759);
nand U1875 (N_1875,In_2405,In_243);
nand U1876 (N_1876,In_911,In_2186);
or U1877 (N_1877,In_2060,In_1587);
and U1878 (N_1878,In_1902,In_1201);
nor U1879 (N_1879,In_2313,In_825);
xnor U1880 (N_1880,In_2936,In_106);
and U1881 (N_1881,In_509,In_447);
and U1882 (N_1882,In_1201,In_1759);
or U1883 (N_1883,In_2750,In_812);
nor U1884 (N_1884,In_2167,In_1744);
xnor U1885 (N_1885,In_756,In_137);
xor U1886 (N_1886,In_513,In_2064);
nand U1887 (N_1887,In_442,In_1826);
and U1888 (N_1888,In_1200,In_2223);
xnor U1889 (N_1889,In_2576,In_2981);
nor U1890 (N_1890,In_1472,In_1157);
xor U1891 (N_1891,In_1756,In_2952);
xnor U1892 (N_1892,In_823,In_2880);
xnor U1893 (N_1893,In_2405,In_2864);
xnor U1894 (N_1894,In_2847,In_54);
xnor U1895 (N_1895,In_2483,In_1790);
and U1896 (N_1896,In_2123,In_2511);
nor U1897 (N_1897,In_1777,In_906);
nor U1898 (N_1898,In_375,In_1624);
xor U1899 (N_1899,In_1365,In_1773);
nand U1900 (N_1900,In_2334,In_2161);
or U1901 (N_1901,In_1969,In_582);
or U1902 (N_1902,In_548,In_1565);
and U1903 (N_1903,In_1962,In_967);
nand U1904 (N_1904,In_51,In_1938);
and U1905 (N_1905,In_63,In_2042);
or U1906 (N_1906,In_1581,In_2505);
nor U1907 (N_1907,In_2133,In_306);
nor U1908 (N_1908,In_2019,In_1114);
xnor U1909 (N_1909,In_1543,In_2673);
xor U1910 (N_1910,In_2760,In_2061);
nand U1911 (N_1911,In_2713,In_1862);
nor U1912 (N_1912,In_924,In_1946);
and U1913 (N_1913,In_2358,In_76);
nand U1914 (N_1914,In_487,In_2722);
nand U1915 (N_1915,In_151,In_69);
nand U1916 (N_1916,In_328,In_2889);
or U1917 (N_1917,In_968,In_646);
or U1918 (N_1918,In_1015,In_2306);
or U1919 (N_1919,In_1749,In_2504);
and U1920 (N_1920,In_1187,In_2446);
or U1921 (N_1921,In_656,In_2268);
nor U1922 (N_1922,In_2708,In_2193);
or U1923 (N_1923,In_2833,In_1228);
xnor U1924 (N_1924,In_323,In_813);
nand U1925 (N_1925,In_439,In_1159);
and U1926 (N_1926,In_2218,In_1540);
or U1927 (N_1927,In_1012,In_1459);
nand U1928 (N_1928,In_2300,In_645);
or U1929 (N_1929,In_1938,In_2707);
and U1930 (N_1930,In_530,In_528);
nor U1931 (N_1931,In_1407,In_1210);
nand U1932 (N_1932,In_1566,In_825);
nand U1933 (N_1933,In_926,In_891);
nand U1934 (N_1934,In_873,In_1406);
or U1935 (N_1935,In_580,In_187);
nand U1936 (N_1936,In_2966,In_2636);
xnor U1937 (N_1937,In_1030,In_1874);
or U1938 (N_1938,In_2776,In_475);
and U1939 (N_1939,In_1860,In_2897);
nor U1940 (N_1940,In_762,In_1580);
nand U1941 (N_1941,In_2888,In_1991);
xor U1942 (N_1942,In_918,In_150);
and U1943 (N_1943,In_1426,In_607);
xor U1944 (N_1944,In_126,In_2240);
and U1945 (N_1945,In_812,In_575);
or U1946 (N_1946,In_1007,In_2193);
xnor U1947 (N_1947,In_1552,In_583);
xor U1948 (N_1948,In_2046,In_332);
xor U1949 (N_1949,In_2715,In_725);
or U1950 (N_1950,In_2665,In_2093);
xor U1951 (N_1951,In_2266,In_867);
or U1952 (N_1952,In_862,In_1082);
or U1953 (N_1953,In_1197,In_722);
nor U1954 (N_1954,In_2871,In_793);
nand U1955 (N_1955,In_2879,In_2449);
xnor U1956 (N_1956,In_806,In_612);
and U1957 (N_1957,In_1184,In_2745);
xnor U1958 (N_1958,In_578,In_2847);
nand U1959 (N_1959,In_695,In_1641);
and U1960 (N_1960,In_1369,In_2182);
or U1961 (N_1961,In_2962,In_458);
xor U1962 (N_1962,In_1807,In_263);
and U1963 (N_1963,In_193,In_312);
nor U1964 (N_1964,In_2224,In_2062);
or U1965 (N_1965,In_872,In_2957);
nand U1966 (N_1966,In_1189,In_1707);
or U1967 (N_1967,In_2524,In_1288);
nor U1968 (N_1968,In_1836,In_6);
nor U1969 (N_1969,In_948,In_2321);
nor U1970 (N_1970,In_236,In_2777);
nand U1971 (N_1971,In_1035,In_2966);
and U1972 (N_1972,In_1735,In_1720);
or U1973 (N_1973,In_1412,In_2521);
and U1974 (N_1974,In_1186,In_507);
xnor U1975 (N_1975,In_2304,In_1068);
nor U1976 (N_1976,In_979,In_1497);
and U1977 (N_1977,In_1007,In_2029);
and U1978 (N_1978,In_2410,In_2552);
nor U1979 (N_1979,In_103,In_1712);
and U1980 (N_1980,In_2290,In_2843);
and U1981 (N_1981,In_648,In_644);
nand U1982 (N_1982,In_2736,In_473);
nor U1983 (N_1983,In_775,In_1484);
nand U1984 (N_1984,In_601,In_2077);
and U1985 (N_1985,In_1519,In_837);
or U1986 (N_1986,In_1967,In_244);
or U1987 (N_1987,In_1371,In_2457);
and U1988 (N_1988,In_772,In_1110);
nor U1989 (N_1989,In_136,In_429);
nand U1990 (N_1990,In_745,In_2339);
xnor U1991 (N_1991,In_2547,In_2332);
xor U1992 (N_1992,In_2017,In_1158);
and U1993 (N_1993,In_1535,In_865);
nand U1994 (N_1994,In_119,In_2315);
or U1995 (N_1995,In_229,In_1075);
xor U1996 (N_1996,In_153,In_114);
nor U1997 (N_1997,In_1216,In_475);
and U1998 (N_1998,In_2664,In_1635);
nor U1999 (N_1999,In_981,In_95);
nand U2000 (N_2000,N_1037,N_975);
and U2001 (N_2001,N_1359,N_117);
or U2002 (N_2002,N_1374,N_881);
nor U2003 (N_2003,N_1155,N_1235);
xor U2004 (N_2004,N_1441,N_1454);
or U2005 (N_2005,N_524,N_883);
nor U2006 (N_2006,N_1408,N_567);
nand U2007 (N_2007,N_26,N_226);
xnor U2008 (N_2008,N_185,N_686);
xnor U2009 (N_2009,N_731,N_356);
and U2010 (N_2010,N_175,N_403);
or U2011 (N_2011,N_45,N_357);
or U2012 (N_2012,N_537,N_987);
and U2013 (N_2013,N_1822,N_304);
xnor U2014 (N_2014,N_1332,N_1941);
or U2015 (N_2015,N_257,N_194);
xor U2016 (N_2016,N_781,N_688);
xor U2017 (N_2017,N_1327,N_1532);
or U2018 (N_2018,N_153,N_1225);
nor U2019 (N_2019,N_934,N_780);
and U2020 (N_2020,N_846,N_825);
and U2021 (N_2021,N_25,N_1743);
nand U2022 (N_2022,N_189,N_1852);
nand U2023 (N_2023,N_1602,N_187);
nor U2024 (N_2024,N_1466,N_806);
or U2025 (N_2025,N_1178,N_1856);
xnor U2026 (N_2026,N_698,N_1913);
nand U2027 (N_2027,N_103,N_1336);
and U2028 (N_2028,N_751,N_1476);
nor U2029 (N_2029,N_1994,N_1043);
and U2030 (N_2030,N_321,N_1540);
or U2031 (N_2031,N_1618,N_1817);
nand U2032 (N_2032,N_1613,N_1224);
and U2033 (N_2033,N_124,N_1715);
or U2034 (N_2034,N_1529,N_1293);
nor U2035 (N_2035,N_108,N_917);
or U2036 (N_2036,N_213,N_1003);
or U2037 (N_2037,N_1075,N_1048);
and U2038 (N_2038,N_711,N_1619);
xnor U2039 (N_2039,N_1786,N_1232);
xnor U2040 (N_2040,N_363,N_1766);
xor U2041 (N_2041,N_1106,N_1152);
and U2042 (N_2042,N_1751,N_1967);
nand U2043 (N_2043,N_1319,N_12);
or U2044 (N_2044,N_1858,N_1203);
or U2045 (N_2045,N_967,N_1682);
nand U2046 (N_2046,N_683,N_211);
nor U2047 (N_2047,N_699,N_1603);
nor U2048 (N_2048,N_912,N_1552);
nand U2049 (N_2049,N_1735,N_663);
or U2050 (N_2050,N_1512,N_1304);
and U2051 (N_2051,N_1382,N_1830);
and U2052 (N_2052,N_690,N_1537);
nand U2053 (N_2053,N_1773,N_1827);
or U2054 (N_2054,N_1947,N_513);
xor U2055 (N_2055,N_366,N_417);
xnor U2056 (N_2056,N_736,N_1939);
or U2057 (N_2057,N_1579,N_40);
xnor U2058 (N_2058,N_1616,N_629);
xor U2059 (N_2059,N_1975,N_633);
nand U2060 (N_2060,N_1121,N_51);
and U2061 (N_2061,N_756,N_1796);
or U2062 (N_2062,N_374,N_1849);
and U2063 (N_2063,N_1657,N_890);
nand U2064 (N_2064,N_1689,N_34);
or U2065 (N_2065,N_260,N_876);
and U2066 (N_2066,N_469,N_1549);
and U2067 (N_2067,N_148,N_1711);
xor U2068 (N_2068,N_292,N_1397);
or U2069 (N_2069,N_1996,N_1626);
nor U2070 (N_2070,N_140,N_1760);
nor U2071 (N_2071,N_702,N_966);
and U2072 (N_2072,N_868,N_556);
xor U2073 (N_2073,N_441,N_1311);
or U2074 (N_2074,N_330,N_241);
nand U2075 (N_2075,N_1890,N_380);
nor U2076 (N_2076,N_986,N_499);
xnor U2077 (N_2077,N_1742,N_1451);
or U2078 (N_2078,N_922,N_1874);
or U2079 (N_2079,N_677,N_1713);
nor U2080 (N_2080,N_765,N_453);
xnor U2081 (N_2081,N_1038,N_997);
nor U2082 (N_2082,N_1222,N_1191);
and U2083 (N_2083,N_794,N_464);
nand U2084 (N_2084,N_381,N_337);
nor U2085 (N_2085,N_1999,N_1060);
nand U2086 (N_2086,N_1197,N_1325);
and U2087 (N_2087,N_1957,N_168);
and U2088 (N_2088,N_64,N_877);
or U2089 (N_2089,N_1204,N_1964);
nand U2090 (N_2090,N_771,N_583);
nand U2091 (N_2091,N_826,N_860);
or U2092 (N_2092,N_691,N_268);
nor U2093 (N_2093,N_1686,N_1472);
xor U2094 (N_2094,N_763,N_801);
nor U2095 (N_2095,N_1872,N_623);
nand U2096 (N_2096,N_1675,N_1103);
nand U2097 (N_2097,N_335,N_1439);
xnor U2098 (N_2098,N_1192,N_1058);
and U2099 (N_2099,N_1193,N_1493);
nand U2100 (N_2100,N_1024,N_1406);
nor U2101 (N_2101,N_1463,N_1386);
and U2102 (N_2102,N_67,N_1503);
or U2103 (N_2103,N_1158,N_1691);
or U2104 (N_2104,N_730,N_306);
xnor U2105 (N_2105,N_1312,N_869);
nand U2106 (N_2106,N_599,N_1568);
xnor U2107 (N_2107,N_899,N_750);
nor U2108 (N_2108,N_1244,N_160);
nor U2109 (N_2109,N_1400,N_1380);
and U2110 (N_2110,N_143,N_578);
xnor U2111 (N_2111,N_1650,N_1068);
nor U2112 (N_2112,N_1535,N_1292);
xor U2113 (N_2113,N_224,N_1880);
and U2114 (N_2114,N_421,N_1298);
nand U2115 (N_2115,N_1693,N_1143);
xor U2116 (N_2116,N_113,N_1169);
nand U2117 (N_2117,N_276,N_1917);
xnor U2118 (N_2118,N_1694,N_414);
xor U2119 (N_2119,N_830,N_1708);
xnor U2120 (N_2120,N_416,N_1378);
and U2121 (N_2121,N_1119,N_1623);
nand U2122 (N_2122,N_1356,N_1099);
and U2123 (N_2123,N_775,N_289);
xor U2124 (N_2124,N_760,N_1139);
nor U2125 (N_2125,N_139,N_1801);
nor U2126 (N_2126,N_666,N_53);
xor U2127 (N_2127,N_1342,N_615);
xnor U2128 (N_2128,N_1847,N_48);
nand U2129 (N_2129,N_59,N_101);
and U2130 (N_2130,N_1710,N_1718);
nand U2131 (N_2131,N_486,N_15);
nand U2132 (N_2132,N_1054,N_866);
and U2133 (N_2133,N_924,N_120);
nand U2134 (N_2134,N_1351,N_1974);
or U2135 (N_2135,N_1923,N_1810);
xor U2136 (N_2136,N_1110,N_1851);
nand U2137 (N_2137,N_938,N_1839);
nor U2138 (N_2138,N_483,N_1213);
nand U2139 (N_2139,N_905,N_563);
and U2140 (N_2140,N_1296,N_11);
xor U2141 (N_2141,N_72,N_1745);
xnor U2142 (N_2142,N_1318,N_1663);
nor U2143 (N_2143,N_1948,N_1412);
nand U2144 (N_2144,N_1971,N_1545);
xnor U2145 (N_2145,N_398,N_271);
and U2146 (N_2146,N_1164,N_575);
and U2147 (N_2147,N_1114,N_624);
xor U2148 (N_2148,N_295,N_115);
nor U2149 (N_2149,N_785,N_1940);
xnor U2150 (N_2150,N_580,N_454);
nor U2151 (N_2151,N_1173,N_1525);
nand U2152 (N_2152,N_1528,N_258);
xor U2153 (N_2153,N_1744,N_776);
nor U2154 (N_2154,N_521,N_498);
xnor U2155 (N_2155,N_1826,N_1092);
or U2156 (N_2156,N_114,N_1286);
and U2157 (N_2157,N_465,N_1183);
xnor U2158 (N_2158,N_1415,N_1358);
or U2159 (N_2159,N_1343,N_548);
nor U2160 (N_2160,N_859,N_201);
xnor U2161 (N_2161,N_66,N_586);
and U2162 (N_2162,N_1490,N_1883);
or U2163 (N_2163,N_1376,N_1362);
xor U2164 (N_2164,N_753,N_635);
nor U2165 (N_2165,N_36,N_1081);
xnor U2166 (N_2166,N_1598,N_1145);
xor U2167 (N_2167,N_1233,N_1085);
and U2168 (N_2168,N_1278,N_1302);
nand U2169 (N_2169,N_1624,N_1930);
nor U2170 (N_2170,N_1901,N_584);
nand U2171 (N_2171,N_689,N_1803);
xnor U2172 (N_2172,N_95,N_525);
xnor U2173 (N_2173,N_823,N_1987);
or U2174 (N_2174,N_1864,N_1128);
and U2175 (N_2175,N_61,N_961);
and U2176 (N_2176,N_485,N_1069);
nor U2177 (N_2177,N_1738,N_661);
and U2178 (N_2178,N_310,N_1953);
nand U2179 (N_2179,N_549,N_1515);
or U2180 (N_2180,N_252,N_1214);
nor U2181 (N_2181,N_1248,N_1868);
xor U2182 (N_2182,N_1017,N_810);
and U2183 (N_2183,N_1869,N_1129);
and U2184 (N_2184,N_1458,N_1909);
nand U2185 (N_2185,N_618,N_1083);
xnor U2186 (N_2186,N_553,N_1254);
or U2187 (N_2187,N_837,N_69);
nand U2188 (N_2188,N_104,N_1435);
nand U2189 (N_2189,N_121,N_747);
and U2190 (N_2190,N_1599,N_1414);
nor U2191 (N_2191,N_1877,N_1889);
and U2192 (N_2192,N_871,N_1554);
nor U2193 (N_2193,N_407,N_972);
nor U2194 (N_2194,N_950,N_565);
or U2195 (N_2195,N_331,N_77);
xnor U2196 (N_2196,N_190,N_1335);
and U2197 (N_2197,N_1679,N_212);
nor U2198 (N_2198,N_1992,N_713);
or U2199 (N_2199,N_861,N_1641);
nand U2200 (N_2200,N_216,N_679);
and U2201 (N_2201,N_1459,N_766);
and U2202 (N_2202,N_350,N_1669);
nand U2203 (N_2203,N_1289,N_438);
nand U2204 (N_2204,N_960,N_1445);
nand U2205 (N_2205,N_1934,N_594);
nand U2206 (N_2206,N_1565,N_1820);
or U2207 (N_2207,N_1671,N_470);
nand U2208 (N_2208,N_1600,N_1984);
nand U2209 (N_2209,N_1063,N_78);
nor U2210 (N_2210,N_770,N_333);
nor U2211 (N_2211,N_184,N_1775);
and U2212 (N_2212,N_1688,N_475);
nand U2213 (N_2213,N_297,N_621);
and U2214 (N_2214,N_1942,N_803);
or U2215 (N_2215,N_610,N_718);
nor U2216 (N_2216,N_1305,N_913);
or U2217 (N_2217,N_259,N_562);
nand U2218 (N_2218,N_491,N_1239);
or U2219 (N_2219,N_569,N_1645);
nor U2220 (N_2220,N_543,N_982);
xnor U2221 (N_2221,N_432,N_1431);
nand U2222 (N_2222,N_723,N_1991);
xor U2223 (N_2223,N_237,N_1405);
or U2224 (N_2224,N_272,N_654);
nand U2225 (N_2225,N_1309,N_1091);
xnor U2226 (N_2226,N_1511,N_92);
or U2227 (N_2227,N_1230,N_1746);
nand U2228 (N_2228,N_551,N_1523);
nand U2229 (N_2229,N_1496,N_1195);
nor U2230 (N_2230,N_444,N_1465);
nor U2231 (N_2231,N_1592,N_449);
and U2232 (N_2232,N_301,N_1281);
nand U2233 (N_2233,N_1547,N_1731);
nand U2234 (N_2234,N_405,N_1842);
or U2235 (N_2235,N_1837,N_238);
nor U2236 (N_2236,N_606,N_1073);
nand U2237 (N_2237,N_340,N_1840);
nand U2238 (N_2238,N_1094,N_1577);
and U2239 (N_2239,N_1135,N_571);
or U2240 (N_2240,N_1906,N_1383);
and U2241 (N_2241,N_1871,N_595);
or U2242 (N_2242,N_1098,N_1768);
or U2243 (N_2243,N_1491,N_996);
nor U2244 (N_2244,N_1208,N_10);
or U2245 (N_2245,N_250,N_75);
nand U2246 (N_2246,N_375,N_1097);
or U2247 (N_2247,N_93,N_1159);
or U2248 (N_2248,N_1120,N_307);
nand U2249 (N_2249,N_164,N_620);
or U2250 (N_2250,N_1390,N_197);
and U2251 (N_2251,N_1709,N_327);
and U2252 (N_2252,N_941,N_445);
and U2253 (N_2253,N_334,N_456);
xnor U2254 (N_2254,N_1597,N_458);
nor U2255 (N_2255,N_755,N_1285);
nand U2256 (N_2256,N_1628,N_1015);
nand U2257 (N_2257,N_362,N_1521);
and U2258 (N_2258,N_1495,N_625);
and U2259 (N_2259,N_1702,N_318);
nand U2260 (N_2260,N_99,N_696);
or U2261 (N_2261,N_1935,N_734);
xor U2262 (N_2262,N_210,N_428);
and U2263 (N_2263,N_1273,N_1564);
nor U2264 (N_2264,N_1680,N_448);
and U2265 (N_2265,N_70,N_1566);
nand U2266 (N_2266,N_943,N_1988);
nor U2267 (N_2267,N_1714,N_1190);
or U2268 (N_2268,N_903,N_530);
nor U2269 (N_2269,N_809,N_1265);
or U2270 (N_2270,N_354,N_740);
nand U2271 (N_2271,N_488,N_743);
nor U2272 (N_2272,N_1583,N_1497);
nor U2273 (N_2273,N_1522,N_1620);
or U2274 (N_2274,N_429,N_1369);
xnor U2275 (N_2275,N_32,N_1313);
or U2276 (N_2276,N_1064,N_1902);
nand U2277 (N_2277,N_523,N_648);
and U2278 (N_2278,N_952,N_1524);
nand U2279 (N_2279,N_332,N_1998);
nand U2280 (N_2280,N_631,N_887);
nand U2281 (N_2281,N_361,N_16);
nand U2282 (N_2282,N_1697,N_1426);
and U2283 (N_2283,N_1571,N_102);
nand U2284 (N_2284,N_1785,N_792);
or U2285 (N_2285,N_1347,N_1968);
xor U2286 (N_2286,N_918,N_954);
nand U2287 (N_2287,N_744,N_1417);
xnor U2288 (N_2288,N_928,N_1654);
nor U2289 (N_2289,N_1268,N_910);
and U2290 (N_2290,N_389,N_1250);
nand U2291 (N_2291,N_681,N_1102);
nor U2292 (N_2292,N_865,N_1381);
or U2293 (N_2293,N_450,N_1464);
xnor U2294 (N_2294,N_1402,N_544);
or U2295 (N_2295,N_1956,N_286);
nor U2296 (N_2296,N_1487,N_1379);
nor U2297 (N_2297,N_157,N_864);
xnor U2298 (N_2298,N_596,N_774);
and U2299 (N_2299,N_795,N_1841);
xor U2300 (N_2300,N_853,N_653);
nand U2301 (N_2301,N_487,N_1020);
xnor U2302 (N_2302,N_24,N_616);
nor U2303 (N_2303,N_822,N_1946);
xnor U2304 (N_2304,N_1301,N_1093);
nor U2305 (N_2305,N_1019,N_128);
or U2306 (N_2306,N_91,N_29);
xor U2307 (N_2307,N_1557,N_1588);
nor U2308 (N_2308,N_1256,N_1717);
nand U2309 (N_2309,N_515,N_1053);
xor U2310 (N_2310,N_1366,N_1115);
and U2311 (N_2311,N_685,N_1506);
or U2312 (N_2312,N_1737,N_1750);
and U2313 (N_2313,N_1432,N_850);
or U2314 (N_2314,N_1084,N_1574);
or U2315 (N_2315,N_670,N_1300);
nor U2316 (N_2316,N_1531,N_540);
xor U2317 (N_2317,N_7,N_1976);
and U2318 (N_2318,N_684,N_1704);
nor U2319 (N_2319,N_715,N_325);
nand U2320 (N_2320,N_1829,N_1368);
nor U2321 (N_2321,N_1189,N_531);
nor U2322 (N_2322,N_273,N_999);
or U2323 (N_2323,N_1185,N_1610);
nor U2324 (N_2324,N_1320,N_1026);
xnor U2325 (N_2325,N_1678,N_855);
nand U2326 (N_2326,N_1891,N_159);
and U2327 (N_2327,N_283,N_1299);
or U2328 (N_2328,N_558,N_974);
xnor U2329 (N_2329,N_669,N_1134);
xor U2330 (N_2330,N_1790,N_1217);
or U2331 (N_2331,N_908,N_430);
nor U2332 (N_2332,N_798,N_607);
xnor U2333 (N_2333,N_886,N_285);
or U2334 (N_2334,N_1642,N_1919);
or U2335 (N_2335,N_1252,N_1527);
nor U2336 (N_2336,N_674,N_1050);
and U2337 (N_2337,N_1629,N_1672);
or U2338 (N_2338,N_1206,N_1072);
nand U2339 (N_2339,N_516,N_1959);
or U2340 (N_2340,N_1945,N_1848);
nor U2341 (N_2341,N_105,N_435);
or U2342 (N_2342,N_1517,N_927);
xor U2343 (N_2343,N_1137,N_1653);
nor U2344 (N_2344,N_1478,N_1033);
and U2345 (N_2345,N_979,N_94);
or U2346 (N_2346,N_1259,N_1799);
or U2347 (N_2347,N_137,N_1067);
and U2348 (N_2348,N_915,N_1898);
nor U2349 (N_2349,N_290,N_642);
or U2350 (N_2350,N_1881,N_1283);
xor U2351 (N_2351,N_1448,N_161);
and U2352 (N_2352,N_1154,N_1587);
xnor U2353 (N_2353,N_341,N_1622);
xnor U2354 (N_2354,N_1365,N_1133);
xor U2355 (N_2355,N_338,N_948);
xor U2356 (N_2356,N_1692,N_254);
xor U2357 (N_2357,N_207,N_667);
xnor U2358 (N_2358,N_1253,N_265);
and U2359 (N_2359,N_719,N_694);
or U2360 (N_2360,N_1260,N_1831);
xnor U2361 (N_2361,N_1684,N_839);
xnor U2362 (N_2362,N_1853,N_1646);
nor U2363 (N_2363,N_1394,N_1627);
or U2364 (N_2364,N_650,N_559);
or U2365 (N_2365,N_1958,N_1882);
or U2366 (N_2366,N_1410,N_1486);
nor U2367 (N_2367,N_505,N_446);
xnor U2368 (N_2368,N_1569,N_873);
or U2369 (N_2369,N_460,N_937);
xnor U2370 (N_2370,N_579,N_1255);
nand U2371 (N_2371,N_1352,N_1427);
nand U2372 (N_2372,N_358,N_821);
nand U2373 (N_2373,N_443,N_958);
nand U2374 (N_2374,N_710,N_1467);
and U2375 (N_2375,N_1409,N_901);
and U2376 (N_2376,N_856,N_1986);
or U2377 (N_2377,N_1823,N_302);
or U2378 (N_2378,N_401,N_697);
nor U2379 (N_2379,N_222,N_141);
nor U2380 (N_2380,N_848,N_712);
and U2381 (N_2381,N_930,N_1360);
or U2382 (N_2382,N_1551,N_879);
nand U2383 (N_2383,N_1809,N_925);
nor U2384 (N_2384,N_646,N_342);
nand U2385 (N_2385,N_1648,N_1924);
nor U2386 (N_2386,N_181,N_1601);
and U2387 (N_2387,N_1635,N_1411);
or U2388 (N_2388,N_1407,N_518);
and U2389 (N_2389,N_1716,N_529);
nand U2390 (N_2390,N_1797,N_1228);
or U2391 (N_2391,N_973,N_976);
xnor U2392 (N_2392,N_716,N_1113);
and U2393 (N_2393,N_779,N_935);
xor U2394 (N_2394,N_500,N_202);
xor U2395 (N_2395,N_1644,N_672);
nand U2396 (N_2396,N_1944,N_1074);
or U2397 (N_2397,N_145,N_135);
and U2398 (N_2398,N_1447,N_1167);
xnor U2399 (N_2399,N_1000,N_1995);
nor U2400 (N_2400,N_1161,N_379);
xnor U2401 (N_2401,N_796,N_983);
or U2402 (N_2402,N_969,N_1863);
or U2403 (N_2403,N_208,N_234);
nor U2404 (N_2404,N_326,N_264);
or U2405 (N_2405,N_39,N_1350);
and U2406 (N_2406,N_1388,N_1078);
nor U2407 (N_2407,N_402,N_1550);
and U2408 (N_2408,N_1754,N_787);
xor U2409 (N_2409,N_344,N_1510);
xor U2410 (N_2410,N_1031,N_1899);
nand U2411 (N_2411,N_1168,N_142);
nor U2412 (N_2412,N_1210,N_1245);
xnor U2413 (N_2413,N_1052,N_1850);
xor U2414 (N_2414,N_628,N_527);
xnor U2415 (N_2415,N_1655,N_1961);
xnor U2416 (N_2416,N_1677,N_1886);
nor U2417 (N_2417,N_277,N_284);
and U2418 (N_2418,N_1662,N_1422);
nor U2419 (N_2419,N_673,N_311);
nand U2420 (N_2420,N_1334,N_965);
xor U2421 (N_2421,N_1720,N_981);
and U2422 (N_2422,N_1770,N_1904);
nand U2423 (N_2423,N_1209,N_1044);
or U2424 (N_2424,N_1361,N_1605);
nand U2425 (N_2425,N_130,N_1982);
xnor U2426 (N_2426,N_1741,N_294);
xor U2427 (N_2427,N_1498,N_151);
and U2428 (N_2428,N_109,N_1440);
nand U2429 (N_2429,N_1326,N_1187);
or U2430 (N_2430,N_1543,N_1219);
or U2431 (N_2431,N_923,N_668);
and U2432 (N_2432,N_1148,N_1008);
nand U2433 (N_2433,N_1212,N_30);
or U2434 (N_2434,N_54,N_1387);
xnor U2435 (N_2435,N_1815,N_299);
nand U2436 (N_2436,N_1955,N_627);
xor U2437 (N_2437,N_1895,N_1546);
or U2438 (N_2438,N_591,N_461);
xnor U2439 (N_2439,N_778,N_1734);
or U2440 (N_2440,N_1739,N_1040);
xnor U2441 (N_2441,N_637,N_501);
xnor U2442 (N_2442,N_962,N_526);
or U2443 (N_2443,N_1127,N_1520);
nand U2444 (N_2444,N_1355,N_1725);
nor U2445 (N_2445,N_1771,N_1166);
nor U2446 (N_2446,N_1845,N_1375);
nor U2447 (N_2447,N_1802,N_1727);
or U2448 (N_2448,N_1444,N_1032);
nand U2449 (N_2449,N_305,N_1896);
nor U2450 (N_2450,N_231,N_1581);
nor U2451 (N_2451,N_1908,N_410);
nand U2452 (N_2452,N_1251,N_1969);
nor U2453 (N_2453,N_1395,N_1246);
or U2454 (N_2454,N_777,N_611);
nand U2455 (N_2455,N_746,N_1866);
or U2456 (N_2456,N_56,N_626);
or U2457 (N_2457,N_415,N_727);
nor U2458 (N_2458,N_968,N_1276);
nor U2459 (N_2459,N_134,N_851);
nand U2460 (N_2460,N_1218,N_1485);
xor U2461 (N_2461,N_154,N_817);
nand U2462 (N_2462,N_71,N_949);
or U2463 (N_2463,N_1978,N_814);
nor U2464 (N_2464,N_22,N_847);
or U2465 (N_2465,N_1501,N_1556);
or U2466 (N_2466,N_198,N_1249);
xnor U2467 (N_2467,N_163,N_811);
or U2468 (N_2468,N_1142,N_119);
and U2469 (N_2469,N_1983,N_1261);
and U2470 (N_2470,N_1471,N_1514);
nor U2471 (N_2471,N_1474,N_20);
xnor U2472 (N_2472,N_1196,N_1595);
nand U2473 (N_2473,N_1772,N_1297);
and U2474 (N_2474,N_1834,N_634);
xor U2475 (N_2475,N_799,N_582);
nand U2476 (N_2476,N_1756,N_1962);
xor U2477 (N_2477,N_1860,N_1157);
nand U2478 (N_2478,N_1783,N_123);
nand U2479 (N_2479,N_1668,N_1401);
nand U2480 (N_2480,N_1198,N_1372);
nand U2481 (N_2481,N_589,N_14);
xnor U2482 (N_2482,N_1077,N_282);
and U2483 (N_2483,N_385,N_1789);
and U2484 (N_2484,N_1095,N_1065);
xor U2485 (N_2485,N_640,N_1617);
or U2486 (N_2486,N_1502,N_1416);
nor U2487 (N_2487,N_1291,N_1314);
and U2488 (N_2488,N_19,N_79);
xor U2489 (N_2489,N_1341,N_1787);
or U2490 (N_2490,N_1649,N_1780);
and U2491 (N_2491,N_555,N_1036);
nand U2492 (N_2492,N_35,N_1582);
xor U2493 (N_2493,N_1791,N_246);
and U2494 (N_2494,N_1205,N_757);
nand U2495 (N_2495,N_225,N_18);
and U2496 (N_2496,N_831,N_312);
nor U2497 (N_2497,N_1703,N_482);
nand U2498 (N_2498,N_959,N_395);
or U2499 (N_2499,N_619,N_936);
nand U2500 (N_2500,N_1371,N_452);
nand U2501 (N_2501,N_1434,N_343);
or U2502 (N_2502,N_1794,N_0);
and U2503 (N_2503,N_1696,N_560);
and U2504 (N_2504,N_1670,N_1461);
and U2505 (N_2505,N_1354,N_98);
xnor U2506 (N_2506,N_782,N_1966);
nor U2507 (N_2507,N_474,N_1492);
xnor U2508 (N_2508,N_827,N_1509);
xor U2509 (N_2509,N_1377,N_1450);
or U2510 (N_2510,N_269,N_291);
and U2511 (N_2511,N_1483,N_717);
and U2512 (N_2512,N_1774,N_1279);
nand U2513 (N_2513,N_977,N_1534);
or U2514 (N_2514,N_1269,N_1176);
or U2515 (N_2515,N_1980,N_682);
and U2516 (N_2516,N_1712,N_1345);
or U2517 (N_2517,N_44,N_1533);
or U2518 (N_2518,N_220,N_1221);
or U2519 (N_2519,N_155,N_322);
and U2520 (N_2520,N_1585,N_991);
xor U2521 (N_2521,N_1997,N_1322);
xor U2522 (N_2522,N_319,N_50);
and U2523 (N_2523,N_1240,N_1938);
nor U2524 (N_2524,N_550,N_630);
and U2525 (N_2525,N_52,N_253);
and U2526 (N_2526,N_639,N_931);
nor U2527 (N_2527,N_479,N_564);
and U2528 (N_2528,N_156,N_281);
nand U2529 (N_2529,N_5,N_1057);
xor U2530 (N_2530,N_1736,N_152);
nand U2531 (N_2531,N_1606,N_904);
and U2532 (N_2532,N_651,N_761);
xnor U2533 (N_2533,N_1442,N_182);
or U2534 (N_2534,N_1242,N_1667);
nor U2535 (N_2535,N_1538,N_1526);
xnor U2536 (N_2536,N_97,N_1636);
or U2537 (N_2537,N_1460,N_144);
nor U2538 (N_2538,N_369,N_835);
or U2539 (N_2539,N_503,N_1324);
or U2540 (N_2540,N_1398,N_1494);
nand U2541 (N_2541,N_721,N_1055);
and U2542 (N_2542,N_784,N_1022);
and U2543 (N_2543,N_23,N_106);
or U2544 (N_2544,N_1757,N_680);
nor U2545 (N_2545,N_243,N_590);
nor U2546 (N_2546,N_174,N_665);
nor U2547 (N_2547,N_1005,N_1002);
nor U2548 (N_2548,N_1719,N_221);
xnor U2549 (N_2549,N_1647,N_179);
nor U2550 (N_2550,N_1722,N_926);
nor U2551 (N_2551,N_722,N_1721);
or U2552 (N_2552,N_31,N_833);
and U2553 (N_2553,N_1887,N_348);
nand U2554 (N_2554,N_1685,N_956);
and U2555 (N_2555,N_228,N_995);
nor U2556 (N_2556,N_309,N_1201);
nand U2557 (N_2557,N_328,N_1634);
xor U2558 (N_2558,N_110,N_517);
nor U2559 (N_2559,N_90,N_612);
and U2560 (N_2560,N_245,N_209);
and U2561 (N_2561,N_63,N_162);
nor U2562 (N_2562,N_539,N_1596);
xnor U2563 (N_2563,N_707,N_1973);
nand U2564 (N_2564,N_1862,N_1014);
xnor U2565 (N_2565,N_1661,N_1813);
nand U2566 (N_2566,N_3,N_1);
or U2567 (N_2567,N_724,N_1784);
nand U2568 (N_2568,N_199,N_1700);
and U2569 (N_2569,N_1855,N_166);
nor U2570 (N_2570,N_535,N_1748);
xor U2571 (N_2571,N_1630,N_1082);
and U2572 (N_2572,N_392,N_1726);
or U2573 (N_2573,N_1473,N_1160);
nor U2574 (N_2574,N_1006,N_1184);
and U2575 (N_2575,N_714,N_1846);
or U2576 (N_2576,N_532,N_368);
nor U2577 (N_2577,N_434,N_376);
or U2578 (N_2578,N_725,N_1270);
xor U2579 (N_2579,N_1066,N_953);
nor U2580 (N_2580,N_720,N_1788);
nand U2581 (N_2581,N_1900,N_1274);
nand U2582 (N_2582,N_73,N_1331);
nor U2583 (N_2583,N_506,N_442);
nor U2584 (N_2584,N_1165,N_481);
xor U2585 (N_2585,N_1468,N_1070);
nor U2586 (N_2586,N_1989,N_1151);
or U2587 (N_2587,N_118,N_978);
nor U2588 (N_2588,N_660,N_236);
xnor U2589 (N_2589,N_1202,N_783);
or U2590 (N_2590,N_574,N_472);
and U2591 (N_2591,N_1364,N_1104);
nor U2592 (N_2592,N_581,N_43);
nor U2593 (N_2593,N_1612,N_1284);
nor U2594 (N_2594,N_597,N_1805);
or U2595 (N_2595,N_1812,N_17);
or U2596 (N_2596,N_1211,N_1660);
or U2597 (N_2597,N_909,N_867);
xor U2598 (N_2598,N_1972,N_1280);
nand U2599 (N_2599,N_424,N_214);
or U2600 (N_2600,N_1330,N_695);
and U2601 (N_2601,N_400,N_463);
and U2602 (N_2602,N_6,N_984);
nor U2603 (N_2603,N_1666,N_459);
or U2604 (N_2604,N_129,N_622);
and U2605 (N_2605,N_832,N_932);
and U2606 (N_2606,N_1117,N_836);
nor U2607 (N_2607,N_1138,N_57);
nand U2608 (N_2608,N_336,N_1767);
or U2609 (N_2609,N_372,N_447);
or U2610 (N_2610,N_480,N_1927);
or U2611 (N_2611,N_1544,N_100);
or U2612 (N_2612,N_738,N_418);
nor U2613 (N_2613,N_1272,N_955);
nor U2614 (N_2614,N_1828,N_298);
xnor U2615 (N_2615,N_764,N_1707);
xnor U2616 (N_2616,N_1340,N_1089);
or U2617 (N_2617,N_1080,N_1306);
nor U2618 (N_2618,N_1965,N_1590);
or U2619 (N_2619,N_745,N_1267);
nor U2620 (N_2620,N_902,N_1243);
and U2621 (N_2621,N_1271,N_1793);
nor U2622 (N_2622,N_180,N_546);
nand U2623 (N_2623,N_992,N_436);
nand U2624 (N_2624,N_1724,N_1056);
xor U2625 (N_2625,N_566,N_1611);
and U2626 (N_2626,N_739,N_1079);
xor U2627 (N_2627,N_520,N_195);
nand U2628 (N_2628,N_1963,N_1023);
nand U2629 (N_2629,N_437,N_1979);
or U2630 (N_2630,N_1854,N_433);
xnor U2631 (N_2631,N_1643,N_788);
and U2632 (N_2632,N_87,N_364);
or U2633 (N_2633,N_200,N_467);
nor U2634 (N_2634,N_1937,N_408);
nand U2635 (N_2635,N_1981,N_455);
xnor U2636 (N_2636,N_1404,N_1317);
nand U2637 (N_2637,N_645,N_1111);
nand U2638 (N_2638,N_1141,N_1194);
nor U2639 (N_2639,N_1162,N_1449);
and U2640 (N_2640,N_288,N_1125);
nor U2641 (N_2641,N_68,N_1951);
or U2642 (N_2642,N_495,N_240);
nand U2643 (N_2643,N_1455,N_62);
and U2644 (N_2644,N_808,N_844);
or U2645 (N_2645,N_1548,N_1519);
xor U2646 (N_2646,N_1761,N_229);
nand U2647 (N_2647,N_1123,N_1396);
and U2648 (N_2648,N_872,N_1393);
nand U2649 (N_2649,N_1118,N_193);
nand U2650 (N_2650,N_116,N_1100);
nor U2651 (N_2651,N_1664,N_1029);
xor U2652 (N_2652,N_1607,N_317);
xnor U2653 (N_2653,N_1753,N_186);
and U2654 (N_2654,N_793,N_863);
nor U2655 (N_2655,N_1687,N_1076);
nand U2656 (N_2656,N_37,N_382);
nor U2657 (N_2657,N_1508,N_898);
and U2658 (N_2658,N_1584,N_215);
or U2659 (N_2659,N_1763,N_1876);
and U2660 (N_2660,N_907,N_843);
and U2661 (N_2661,N_897,N_409);
xnor U2662 (N_2662,N_1107,N_383);
xor U2663 (N_2663,N_21,N_1475);
nand U2664 (N_2664,N_492,N_440);
nor U2665 (N_2665,N_88,N_287);
nor U2666 (N_2666,N_1798,N_896);
nand U2667 (N_2667,N_536,N_1216);
and U2668 (N_2668,N_1257,N_701);
nor U2669 (N_2669,N_1457,N_478);
nand U2670 (N_2670,N_638,N_643);
and U2671 (N_2671,N_1391,N_790);
nor U2672 (N_2672,N_852,N_700);
nor U2673 (N_2673,N_497,N_1188);
or U2674 (N_2674,N_880,N_916);
and U2675 (N_2675,N_373,N_920);
or U2676 (N_2676,N_1749,N_617);
nor U2677 (N_2677,N_1572,N_1857);
and U2678 (N_2678,N_1013,N_1329);
or U2679 (N_2679,N_248,N_749);
xor U2680 (N_2680,N_1418,N_1004);
xor U2681 (N_2681,N_1928,N_1061);
xnor U2682 (N_2682,N_192,N_613);
xor U2683 (N_2683,N_1456,N_404);
nor U2684 (N_2684,N_1413,N_963);
nand U2685 (N_2685,N_58,N_947);
and U2686 (N_2686,N_875,N_1621);
nor U2687 (N_2687,N_576,N_352);
nor U2688 (N_2688,N_1096,N_1516);
nand U2689 (N_2689,N_1781,N_1960);
xnor U2690 (N_2690,N_391,N_1237);
nor U2691 (N_2691,N_732,N_280);
and U2692 (N_2692,N_76,N_33);
nor U2693 (N_2693,N_1423,N_693);
nand U2694 (N_2694,N_845,N_1370);
nand U2695 (N_2695,N_985,N_223);
and U2696 (N_2696,N_413,N_1765);
nor U2697 (N_2697,N_568,N_994);
nor U2698 (N_2698,N_547,N_218);
or U2699 (N_2699,N_111,N_1594);
nand U2700 (N_2700,N_1752,N_1912);
nand U2701 (N_2701,N_1907,N_1925);
xor U2702 (N_2702,N_1262,N_1348);
and U2703 (N_2703,N_1832,N_545);
and U2704 (N_2704,N_133,N_1488);
nand U2705 (N_2705,N_494,N_541);
and U2706 (N_2706,N_1021,N_598);
and U2707 (N_2707,N_1042,N_46);
nand U2708 (N_2708,N_807,N_227);
nor U2709 (N_2709,N_313,N_1640);
xnor U2710 (N_2710,N_1016,N_1949);
xnor U2711 (N_2711,N_1373,N_854);
nor U2712 (N_2712,N_1425,N_878);
nand U2713 (N_2713,N_577,N_768);
nand U2714 (N_2714,N_1045,N_2);
nand U2715 (N_2715,N_55,N_561);
or U2716 (N_2716,N_1652,N_692);
nand U2717 (N_2717,N_1747,N_1806);
nand U2718 (N_2718,N_1504,N_819);
nand U2719 (N_2719,N_1295,N_862);
or U2720 (N_2720,N_1795,N_1170);
nor U2721 (N_2721,N_1541,N_1695);
and U2722 (N_2722,N_1580,N_204);
xnor U2723 (N_2723,N_528,N_1163);
nand U2724 (N_2724,N_664,N_1929);
and U2725 (N_2725,N_1762,N_1130);
and U2726 (N_2726,N_178,N_1266);
and U2727 (N_2727,N_1604,N_1489);
or U2728 (N_2728,N_1690,N_998);
nand U2729 (N_2729,N_980,N_1699);
and U2730 (N_2730,N_1282,N_993);
xor U2731 (N_2731,N_773,N_1446);
nor U2732 (N_2732,N_1698,N_614);
nor U2733 (N_2733,N_1769,N_316);
or U2734 (N_2734,N_1918,N_1367);
or U2735 (N_2735,N_279,N_1764);
or U2736 (N_2736,N_451,N_1659);
or U2737 (N_2737,N_1140,N_1438);
nor U2738 (N_2738,N_324,N_1778);
xnor U2739 (N_2739,N_27,N_1041);
and U2740 (N_2740,N_1333,N_150);
or U2741 (N_2741,N_1888,N_945);
or U2742 (N_2742,N_1625,N_601);
nand U2743 (N_2743,N_708,N_802);
and U2744 (N_2744,N_351,N_127);
and U2745 (N_2745,N_125,N_1885);
nor U2746 (N_2746,N_360,N_1172);
xor U2747 (N_2747,N_183,N_1589);
nand U2748 (N_2748,N_605,N_813);
nor U2749 (N_2749,N_347,N_1171);
nand U2750 (N_2750,N_849,N_65);
or U2751 (N_2751,N_1560,N_320);
nor U2752 (N_2752,N_641,N_1051);
nand U2753 (N_2753,N_158,N_592);
or U2754 (N_2754,N_1484,N_1915);
nor U2755 (N_2755,N_89,N_588);
or U2756 (N_2756,N_1559,N_426);
or U2757 (N_2757,N_1816,N_509);
xor U2758 (N_2758,N_767,N_255);
nor U2759 (N_2759,N_1873,N_1665);
or U2760 (N_2760,N_1001,N_1452);
nor U2761 (N_2761,N_1843,N_726);
xor U2762 (N_2762,N_1288,N_647);
and U2763 (N_2763,N_1639,N_1182);
xnor U2764 (N_2764,N_267,N_1507);
and U2765 (N_2765,N_1153,N_800);
nor U2766 (N_2766,N_1807,N_838);
xnor U2767 (N_2767,N_1859,N_1561);
xnor U2768 (N_2768,N_371,N_86);
nor U2769 (N_2769,N_1223,N_112);
and U2770 (N_2770,N_906,N_1215);
nor U2771 (N_2771,N_346,N_786);
xor U2772 (N_2772,N_275,N_1615);
xor U2773 (N_2773,N_1836,N_1954);
nor U2774 (N_2774,N_754,N_1263);
nor U2775 (N_2775,N_656,N_169);
nand U2776 (N_2776,N_1943,N_1800);
and U2777 (N_2777,N_60,N_1567);
xor U2778 (N_2778,N_812,N_911);
and U2779 (N_2779,N_422,N_1730);
and U2780 (N_2780,N_1570,N_552);
nand U2781 (N_2781,N_772,N_293);
xor U2782 (N_2782,N_370,N_655);
and U2783 (N_2783,N_493,N_1328);
or U2784 (N_2784,N_1818,N_964);
xor U2785 (N_2785,N_315,N_1419);
xnor U2786 (N_2786,N_419,N_74);
and U2787 (N_2787,N_81,N_946);
nand U2788 (N_2788,N_235,N_13);
and U2789 (N_2789,N_874,N_1825);
xnor U2790 (N_2790,N_476,N_818);
xor U2791 (N_2791,N_1985,N_83);
nor U2792 (N_2792,N_1903,N_9);
and U2793 (N_2793,N_900,N_1555);
nor U2794 (N_2794,N_1062,N_1144);
nor U2795 (N_2795,N_1136,N_1838);
xor U2796 (N_2796,N_323,N_1658);
or U2797 (N_2797,N_274,N_1200);
xnor U2798 (N_2798,N_261,N_1027);
nand U2799 (N_2799,N_1156,N_511);
nor U2800 (N_2800,N_1303,N_1363);
or U2801 (N_2801,N_1732,N_841);
and U2802 (N_2802,N_314,N_733);
and U2803 (N_2803,N_957,N_329);
and U2804 (N_2804,N_232,N_534);
xnor U2805 (N_2805,N_251,N_1729);
nor U2806 (N_2806,N_386,N_1952);
nor U2807 (N_2807,N_171,N_570);
or U2808 (N_2808,N_1275,N_468);
nand U2809 (N_2809,N_1573,N_1453);
or U2810 (N_2810,N_573,N_1861);
and U2811 (N_2811,N_951,N_1733);
xor U2812 (N_2812,N_49,N_1116);
nand U2813 (N_2813,N_1310,N_394);
nor U2814 (N_2814,N_1776,N_173);
xor U2815 (N_2815,N_1344,N_1884);
nor U2816 (N_2816,N_1443,N_687);
and U2817 (N_2817,N_1150,N_1047);
nor U2818 (N_2818,N_38,N_196);
xnor U2819 (N_2819,N_41,N_1892);
and U2820 (N_2820,N_652,N_1911);
and U2821 (N_2821,N_510,N_939);
or U2822 (N_2822,N_1681,N_728);
nor U2823 (N_2823,N_882,N_1146);
and U2824 (N_2824,N_149,N_1878);
and U2825 (N_2825,N_1477,N_632);
xnor U2826 (N_2826,N_4,N_1804);
or U2827 (N_2827,N_729,N_296);
xnor U2828 (N_2828,N_484,N_1220);
xor U2829 (N_2829,N_1936,N_1294);
xor U2830 (N_2830,N_1910,N_703);
and U2831 (N_2831,N_399,N_1403);
nor U2832 (N_2832,N_1542,N_929);
or U2833 (N_2833,N_678,N_791);
or U2834 (N_2834,N_136,N_933);
xor U2835 (N_2835,N_1049,N_1088);
nor U2836 (N_2836,N_752,N_249);
nor U2837 (N_2837,N_572,N_858);
or U2838 (N_2838,N_519,N_270);
or U2839 (N_2839,N_557,N_471);
nor U2840 (N_2840,N_406,N_1631);
nand U2841 (N_2841,N_1247,N_593);
xor U2842 (N_2842,N_1920,N_365);
nand U2843 (N_2843,N_411,N_1231);
and U2844 (N_2844,N_1177,N_349);
xor U2845 (N_2845,N_893,N_1337);
and U2846 (N_2846,N_1059,N_191);
or U2847 (N_2847,N_762,N_244);
nand U2848 (N_2848,N_427,N_1614);
and U2849 (N_2849,N_585,N_1108);
or U2850 (N_2850,N_1905,N_1226);
or U2851 (N_2851,N_359,N_1500);
xnor U2852 (N_2852,N_247,N_1701);
nor U2853 (N_2853,N_1513,N_1632);
and U2854 (N_2854,N_1132,N_1034);
and U2855 (N_2855,N_1931,N_1993);
nor U2856 (N_2856,N_671,N_1035);
and U2857 (N_2857,N_1833,N_895);
nand U2858 (N_2858,N_233,N_676);
and U2859 (N_2859,N_504,N_1357);
or U2860 (N_2860,N_1287,N_266);
or U2861 (N_2861,N_759,N_1147);
xnor U2862 (N_2862,N_824,N_1437);
and U2863 (N_2863,N_1740,N_1424);
xor U2864 (N_2864,N_1518,N_1633);
and U2865 (N_2865,N_1656,N_944);
xnor U2866 (N_2866,N_891,N_1346);
or U2867 (N_2867,N_587,N_820);
xor U2868 (N_2868,N_431,N_1428);
xnor U2869 (N_2869,N_42,N_602);
xor U2870 (N_2870,N_1576,N_658);
or U2871 (N_2871,N_1637,N_1811);
xor U2872 (N_2872,N_816,N_704);
or U2873 (N_2873,N_439,N_705);
or U2874 (N_2874,N_741,N_1349);
nor U2875 (N_2875,N_278,N_1420);
nand U2876 (N_2876,N_1009,N_1124);
and U2877 (N_2877,N_804,N_1539);
and U2878 (N_2878,N_1315,N_1338);
xor U2879 (N_2879,N_80,N_609);
xnor U2880 (N_2880,N_709,N_1018);
or U2881 (N_2881,N_748,N_206);
xnor U2882 (N_2882,N_1462,N_1175);
nor U2883 (N_2883,N_1608,N_554);
or U2884 (N_2884,N_353,N_1339);
and U2885 (N_2885,N_466,N_1385);
xnor U2886 (N_2886,N_649,N_1821);
or U2887 (N_2887,N_8,N_1011);
nor U2888 (N_2888,N_205,N_1926);
nand U2889 (N_2889,N_1536,N_769);
xnor U2890 (N_2890,N_970,N_892);
xnor U2891 (N_2891,N_262,N_1012);
or U2892 (N_2892,N_1086,N_203);
nand U2893 (N_2893,N_1932,N_1593);
xnor U2894 (N_2894,N_1553,N_263);
xor U2895 (N_2895,N_489,N_1779);
nor U2896 (N_2896,N_1323,N_1728);
xor U2897 (N_2897,N_940,N_420);
nand U2898 (N_2898,N_308,N_1867);
nand U2899 (N_2899,N_805,N_1429);
nor U2900 (N_2900,N_1112,N_1824);
nand U2901 (N_2901,N_82,N_706);
or U2902 (N_2902,N_396,N_1025);
or U2903 (N_2903,N_1990,N_1392);
xor U2904 (N_2904,N_507,N_1782);
xnor U2905 (N_2905,N_1353,N_1705);
nand U2906 (N_2906,N_1258,N_1897);
and U2907 (N_2907,N_122,N_1236);
xor U2908 (N_2908,N_1007,N_397);
nand U2909 (N_2909,N_742,N_1480);
xor U2910 (N_2910,N_1563,N_1087);
nor U2911 (N_2911,N_496,N_789);
nor U2912 (N_2912,N_303,N_1835);
or U2913 (N_2913,N_172,N_1470);
and U2914 (N_2914,N_1922,N_888);
xor U2915 (N_2915,N_219,N_1179);
nand U2916 (N_2916,N_1039,N_870);
or U2917 (N_2917,N_1030,N_815);
and U2918 (N_2918,N_659,N_457);
xor U2919 (N_2919,N_96,N_604);
nor U2920 (N_2920,N_1308,N_1105);
nor U2921 (N_2921,N_1844,N_1609);
and U2922 (N_2922,N_1307,N_502);
and U2923 (N_2923,N_1436,N_170);
and U2924 (N_2924,N_146,N_1101);
and U2925 (N_2925,N_1290,N_885);
nand U2926 (N_2926,N_737,N_1950);
nand U2927 (N_2927,N_1122,N_1758);
and U2928 (N_2928,N_126,N_1241);
nor U2929 (N_2929,N_473,N_1469);
nor U2930 (N_2930,N_107,N_1384);
and U2931 (N_2931,N_914,N_542);
or U2932 (N_2932,N_828,N_921);
nor U2933 (N_2933,N_533,N_1562);
nand U2934 (N_2934,N_603,N_1389);
nor U2935 (N_2935,N_988,N_1481);
xnor U2936 (N_2936,N_355,N_388);
xor U2937 (N_2937,N_797,N_1819);
xor U2938 (N_2938,N_1199,N_242);
nand U2939 (N_2939,N_1264,N_608);
and U2940 (N_2940,N_85,N_522);
and U2941 (N_2941,N_1421,N_1186);
or U2942 (N_2942,N_1651,N_1321);
and U2943 (N_2943,N_1792,N_378);
and U2944 (N_2944,N_1586,N_829);
and U2945 (N_2945,N_1109,N_644);
or U2946 (N_2946,N_857,N_1673);
nor U2947 (N_2947,N_1126,N_1977);
and U2948 (N_2948,N_490,N_840);
or U2949 (N_2949,N_1071,N_1174);
and U2950 (N_2950,N_1399,N_1638);
xor U2951 (N_2951,N_842,N_28);
nor U2952 (N_2952,N_675,N_147);
and U2953 (N_2953,N_894,N_1879);
or U2954 (N_2954,N_1482,N_1914);
or U2955 (N_2955,N_1814,N_1808);
xnor U2956 (N_2956,N_538,N_377);
nor U2957 (N_2957,N_165,N_84);
nor U2958 (N_2958,N_1870,N_1575);
or U2959 (N_2959,N_1530,N_367);
nor U2960 (N_2960,N_230,N_942);
nor U2961 (N_2961,N_1131,N_1916);
nor U2962 (N_2962,N_1046,N_971);
xor U2963 (N_2963,N_1028,N_990);
and U2964 (N_2964,N_477,N_339);
xor U2965 (N_2965,N_1894,N_1090);
or U2966 (N_2966,N_132,N_662);
xnor U2967 (N_2967,N_1674,N_131);
xnor U2968 (N_2968,N_1238,N_384);
nor U2969 (N_2969,N_1970,N_256);
and U2970 (N_2970,N_462,N_412);
or U2971 (N_2971,N_188,N_884);
or U2972 (N_2972,N_1499,N_345);
and U2973 (N_2973,N_514,N_1430);
and U2974 (N_2974,N_889,N_1181);
and U2975 (N_2975,N_423,N_834);
nor U2976 (N_2976,N_989,N_735);
xnor U2977 (N_2977,N_390,N_1755);
or U2978 (N_2978,N_1207,N_636);
nor U2979 (N_2979,N_1180,N_1316);
nor U2980 (N_2980,N_300,N_138);
nor U2981 (N_2981,N_1676,N_1433);
or U2982 (N_2982,N_512,N_758);
or U2983 (N_2983,N_600,N_239);
xor U2984 (N_2984,N_1578,N_1227);
and U2985 (N_2985,N_508,N_1591);
nand U2986 (N_2986,N_177,N_1865);
and U2987 (N_2987,N_393,N_1759);
and U2988 (N_2988,N_1893,N_1723);
and U2989 (N_2989,N_176,N_167);
xnor U2990 (N_2990,N_1234,N_657);
nand U2991 (N_2991,N_1921,N_1875);
and U2992 (N_2992,N_1277,N_47);
xor U2993 (N_2993,N_1479,N_1933);
and U2994 (N_2994,N_1706,N_1149);
nor U2995 (N_2995,N_1777,N_919);
or U2996 (N_2996,N_387,N_1505);
xor U2997 (N_2997,N_1010,N_1229);
xor U2998 (N_2998,N_1558,N_1683);
and U2999 (N_2999,N_425,N_217);
xor U3000 (N_3000,N_1827,N_1145);
and U3001 (N_3001,N_258,N_1712);
nor U3002 (N_3002,N_89,N_1853);
or U3003 (N_3003,N_1362,N_1473);
and U3004 (N_3004,N_203,N_1592);
and U3005 (N_3005,N_453,N_504);
nor U3006 (N_3006,N_1157,N_369);
or U3007 (N_3007,N_1853,N_1059);
xnor U3008 (N_3008,N_1000,N_907);
xor U3009 (N_3009,N_126,N_1729);
or U3010 (N_3010,N_1254,N_822);
xor U3011 (N_3011,N_1674,N_839);
nand U3012 (N_3012,N_804,N_1925);
xnor U3013 (N_3013,N_1891,N_1940);
and U3014 (N_3014,N_503,N_182);
xor U3015 (N_3015,N_713,N_944);
or U3016 (N_3016,N_1937,N_1950);
and U3017 (N_3017,N_945,N_1433);
nor U3018 (N_3018,N_1955,N_632);
and U3019 (N_3019,N_1634,N_975);
or U3020 (N_3020,N_92,N_18);
nand U3021 (N_3021,N_574,N_1603);
nor U3022 (N_3022,N_1496,N_709);
or U3023 (N_3023,N_635,N_407);
nand U3024 (N_3024,N_322,N_711);
or U3025 (N_3025,N_978,N_1274);
and U3026 (N_3026,N_1088,N_15);
nor U3027 (N_3027,N_1300,N_1330);
and U3028 (N_3028,N_1494,N_165);
or U3029 (N_3029,N_947,N_1380);
nand U3030 (N_3030,N_1059,N_196);
or U3031 (N_3031,N_17,N_929);
nand U3032 (N_3032,N_1255,N_1417);
and U3033 (N_3033,N_1567,N_1841);
nor U3034 (N_3034,N_969,N_1490);
and U3035 (N_3035,N_37,N_1888);
nand U3036 (N_3036,N_1551,N_290);
nor U3037 (N_3037,N_318,N_1922);
or U3038 (N_3038,N_985,N_1566);
nor U3039 (N_3039,N_1296,N_504);
nor U3040 (N_3040,N_1378,N_1392);
or U3041 (N_3041,N_373,N_1148);
and U3042 (N_3042,N_786,N_1136);
and U3043 (N_3043,N_659,N_1183);
and U3044 (N_3044,N_326,N_863);
xnor U3045 (N_3045,N_1030,N_1004);
nor U3046 (N_3046,N_1614,N_1165);
nor U3047 (N_3047,N_954,N_1728);
nand U3048 (N_3048,N_673,N_329);
xnor U3049 (N_3049,N_789,N_267);
nand U3050 (N_3050,N_430,N_1739);
or U3051 (N_3051,N_1769,N_541);
and U3052 (N_3052,N_946,N_394);
or U3053 (N_3053,N_538,N_1515);
or U3054 (N_3054,N_1290,N_93);
nor U3055 (N_3055,N_1482,N_181);
or U3056 (N_3056,N_1060,N_886);
or U3057 (N_3057,N_1674,N_1930);
xor U3058 (N_3058,N_1629,N_1321);
and U3059 (N_3059,N_249,N_1387);
and U3060 (N_3060,N_1663,N_891);
or U3061 (N_3061,N_724,N_226);
nor U3062 (N_3062,N_301,N_1215);
or U3063 (N_3063,N_65,N_219);
xnor U3064 (N_3064,N_139,N_209);
and U3065 (N_3065,N_97,N_984);
nand U3066 (N_3066,N_913,N_1116);
and U3067 (N_3067,N_1077,N_395);
nand U3068 (N_3068,N_374,N_1632);
xnor U3069 (N_3069,N_691,N_623);
and U3070 (N_3070,N_32,N_1598);
nand U3071 (N_3071,N_1380,N_193);
nand U3072 (N_3072,N_450,N_216);
and U3073 (N_3073,N_415,N_849);
nor U3074 (N_3074,N_287,N_465);
xor U3075 (N_3075,N_1295,N_1108);
xnor U3076 (N_3076,N_1053,N_804);
nand U3077 (N_3077,N_1437,N_1218);
nand U3078 (N_3078,N_1614,N_748);
nor U3079 (N_3079,N_846,N_815);
nor U3080 (N_3080,N_1395,N_113);
xnor U3081 (N_3081,N_107,N_145);
xnor U3082 (N_3082,N_683,N_797);
or U3083 (N_3083,N_967,N_1221);
and U3084 (N_3084,N_1694,N_1745);
or U3085 (N_3085,N_242,N_1969);
nand U3086 (N_3086,N_544,N_1595);
xnor U3087 (N_3087,N_183,N_552);
nor U3088 (N_3088,N_1929,N_1535);
xnor U3089 (N_3089,N_1877,N_8);
or U3090 (N_3090,N_1164,N_100);
nor U3091 (N_3091,N_700,N_912);
or U3092 (N_3092,N_1299,N_1868);
nand U3093 (N_3093,N_819,N_736);
nand U3094 (N_3094,N_1937,N_276);
nand U3095 (N_3095,N_82,N_1295);
nand U3096 (N_3096,N_1595,N_729);
xor U3097 (N_3097,N_875,N_132);
nor U3098 (N_3098,N_1504,N_659);
nand U3099 (N_3099,N_703,N_1411);
nand U3100 (N_3100,N_6,N_150);
and U3101 (N_3101,N_692,N_1823);
or U3102 (N_3102,N_1610,N_1063);
nand U3103 (N_3103,N_979,N_895);
xor U3104 (N_3104,N_265,N_1914);
nor U3105 (N_3105,N_589,N_1180);
nor U3106 (N_3106,N_1199,N_297);
nand U3107 (N_3107,N_369,N_492);
and U3108 (N_3108,N_310,N_1835);
and U3109 (N_3109,N_836,N_1365);
xnor U3110 (N_3110,N_100,N_1047);
nand U3111 (N_3111,N_1969,N_969);
or U3112 (N_3112,N_1353,N_422);
and U3113 (N_3113,N_659,N_641);
xor U3114 (N_3114,N_309,N_317);
xnor U3115 (N_3115,N_1419,N_1745);
and U3116 (N_3116,N_1291,N_1387);
or U3117 (N_3117,N_1183,N_32);
and U3118 (N_3118,N_452,N_543);
xor U3119 (N_3119,N_452,N_1310);
xor U3120 (N_3120,N_1580,N_1504);
and U3121 (N_3121,N_1209,N_229);
or U3122 (N_3122,N_627,N_644);
and U3123 (N_3123,N_1145,N_604);
nor U3124 (N_3124,N_48,N_758);
and U3125 (N_3125,N_1033,N_1511);
nand U3126 (N_3126,N_1930,N_1059);
or U3127 (N_3127,N_1286,N_1974);
nor U3128 (N_3128,N_485,N_1160);
and U3129 (N_3129,N_198,N_1914);
nand U3130 (N_3130,N_1716,N_1000);
xor U3131 (N_3131,N_353,N_808);
and U3132 (N_3132,N_389,N_80);
xor U3133 (N_3133,N_128,N_417);
or U3134 (N_3134,N_1018,N_1378);
xnor U3135 (N_3135,N_765,N_726);
nand U3136 (N_3136,N_1448,N_349);
and U3137 (N_3137,N_752,N_342);
xor U3138 (N_3138,N_1745,N_959);
xnor U3139 (N_3139,N_49,N_59);
nor U3140 (N_3140,N_1512,N_1511);
xnor U3141 (N_3141,N_391,N_1347);
nor U3142 (N_3142,N_922,N_753);
or U3143 (N_3143,N_639,N_146);
nor U3144 (N_3144,N_1907,N_266);
xnor U3145 (N_3145,N_624,N_1248);
xnor U3146 (N_3146,N_1553,N_170);
nor U3147 (N_3147,N_453,N_1294);
nor U3148 (N_3148,N_937,N_1458);
nor U3149 (N_3149,N_440,N_899);
or U3150 (N_3150,N_295,N_965);
and U3151 (N_3151,N_867,N_1720);
nand U3152 (N_3152,N_979,N_1891);
xor U3153 (N_3153,N_1326,N_378);
xnor U3154 (N_3154,N_1739,N_825);
and U3155 (N_3155,N_799,N_508);
xnor U3156 (N_3156,N_20,N_756);
and U3157 (N_3157,N_248,N_1339);
nand U3158 (N_3158,N_1423,N_831);
xor U3159 (N_3159,N_639,N_482);
nor U3160 (N_3160,N_1972,N_1952);
xnor U3161 (N_3161,N_297,N_458);
nor U3162 (N_3162,N_1861,N_306);
and U3163 (N_3163,N_1027,N_472);
nand U3164 (N_3164,N_139,N_1725);
and U3165 (N_3165,N_647,N_829);
and U3166 (N_3166,N_630,N_1169);
or U3167 (N_3167,N_148,N_1240);
nor U3168 (N_3168,N_1941,N_885);
nor U3169 (N_3169,N_379,N_784);
and U3170 (N_3170,N_1108,N_90);
nand U3171 (N_3171,N_1558,N_470);
or U3172 (N_3172,N_765,N_292);
nand U3173 (N_3173,N_387,N_541);
and U3174 (N_3174,N_1447,N_1887);
xnor U3175 (N_3175,N_1153,N_1008);
nand U3176 (N_3176,N_1155,N_644);
xor U3177 (N_3177,N_1294,N_163);
nand U3178 (N_3178,N_1146,N_213);
nand U3179 (N_3179,N_1100,N_1626);
and U3180 (N_3180,N_656,N_6);
nor U3181 (N_3181,N_163,N_1910);
nor U3182 (N_3182,N_228,N_768);
nor U3183 (N_3183,N_570,N_153);
or U3184 (N_3184,N_354,N_794);
xor U3185 (N_3185,N_519,N_909);
nand U3186 (N_3186,N_1759,N_1462);
xor U3187 (N_3187,N_184,N_1332);
and U3188 (N_3188,N_953,N_1536);
xnor U3189 (N_3189,N_1169,N_941);
and U3190 (N_3190,N_1361,N_1250);
and U3191 (N_3191,N_503,N_593);
nor U3192 (N_3192,N_1059,N_628);
xnor U3193 (N_3193,N_1742,N_900);
nand U3194 (N_3194,N_602,N_1871);
xnor U3195 (N_3195,N_969,N_1362);
xnor U3196 (N_3196,N_1474,N_574);
or U3197 (N_3197,N_130,N_242);
nor U3198 (N_3198,N_949,N_122);
nand U3199 (N_3199,N_526,N_727);
and U3200 (N_3200,N_1774,N_994);
nand U3201 (N_3201,N_23,N_1993);
nand U3202 (N_3202,N_731,N_953);
and U3203 (N_3203,N_1809,N_240);
nor U3204 (N_3204,N_1873,N_1515);
nor U3205 (N_3205,N_617,N_202);
xnor U3206 (N_3206,N_1876,N_1039);
and U3207 (N_3207,N_363,N_1122);
or U3208 (N_3208,N_873,N_1975);
or U3209 (N_3209,N_1136,N_1336);
and U3210 (N_3210,N_494,N_1215);
nor U3211 (N_3211,N_1465,N_656);
xnor U3212 (N_3212,N_1276,N_1963);
and U3213 (N_3213,N_789,N_958);
xor U3214 (N_3214,N_1135,N_1045);
nand U3215 (N_3215,N_1510,N_1983);
or U3216 (N_3216,N_1878,N_1354);
nor U3217 (N_3217,N_973,N_1693);
and U3218 (N_3218,N_1126,N_1324);
or U3219 (N_3219,N_1062,N_1856);
or U3220 (N_3220,N_1191,N_479);
and U3221 (N_3221,N_1145,N_13);
and U3222 (N_3222,N_657,N_781);
nor U3223 (N_3223,N_829,N_212);
and U3224 (N_3224,N_1243,N_1090);
nand U3225 (N_3225,N_877,N_363);
nor U3226 (N_3226,N_1704,N_330);
and U3227 (N_3227,N_43,N_266);
or U3228 (N_3228,N_1128,N_564);
nor U3229 (N_3229,N_1805,N_55);
and U3230 (N_3230,N_959,N_1301);
nor U3231 (N_3231,N_1947,N_678);
and U3232 (N_3232,N_135,N_319);
xnor U3233 (N_3233,N_964,N_936);
xor U3234 (N_3234,N_1390,N_470);
or U3235 (N_3235,N_794,N_1052);
or U3236 (N_3236,N_1735,N_1241);
and U3237 (N_3237,N_343,N_317);
xor U3238 (N_3238,N_375,N_169);
or U3239 (N_3239,N_255,N_326);
or U3240 (N_3240,N_391,N_1777);
and U3241 (N_3241,N_1702,N_876);
and U3242 (N_3242,N_864,N_1115);
nor U3243 (N_3243,N_1491,N_676);
and U3244 (N_3244,N_488,N_106);
nor U3245 (N_3245,N_644,N_812);
nor U3246 (N_3246,N_1643,N_1472);
or U3247 (N_3247,N_924,N_1055);
nor U3248 (N_3248,N_730,N_1345);
nor U3249 (N_3249,N_689,N_1326);
or U3250 (N_3250,N_1574,N_1334);
and U3251 (N_3251,N_4,N_1525);
or U3252 (N_3252,N_1253,N_521);
nand U3253 (N_3253,N_1943,N_221);
and U3254 (N_3254,N_7,N_1330);
nor U3255 (N_3255,N_639,N_1038);
or U3256 (N_3256,N_798,N_1985);
or U3257 (N_3257,N_998,N_878);
and U3258 (N_3258,N_1530,N_1714);
and U3259 (N_3259,N_811,N_997);
xor U3260 (N_3260,N_1459,N_1904);
nand U3261 (N_3261,N_1371,N_345);
xor U3262 (N_3262,N_754,N_1261);
or U3263 (N_3263,N_162,N_1436);
nor U3264 (N_3264,N_1277,N_325);
nor U3265 (N_3265,N_1811,N_366);
and U3266 (N_3266,N_1458,N_802);
or U3267 (N_3267,N_1960,N_1824);
and U3268 (N_3268,N_848,N_200);
nand U3269 (N_3269,N_20,N_793);
nand U3270 (N_3270,N_14,N_882);
nor U3271 (N_3271,N_1049,N_153);
xnor U3272 (N_3272,N_1676,N_155);
nand U3273 (N_3273,N_1773,N_226);
or U3274 (N_3274,N_1909,N_1986);
nor U3275 (N_3275,N_68,N_1833);
and U3276 (N_3276,N_120,N_1993);
nand U3277 (N_3277,N_1492,N_1986);
and U3278 (N_3278,N_926,N_1571);
and U3279 (N_3279,N_1324,N_789);
and U3280 (N_3280,N_279,N_420);
xnor U3281 (N_3281,N_606,N_1904);
xor U3282 (N_3282,N_1395,N_381);
and U3283 (N_3283,N_1472,N_1551);
or U3284 (N_3284,N_173,N_474);
or U3285 (N_3285,N_403,N_1507);
or U3286 (N_3286,N_1321,N_1457);
and U3287 (N_3287,N_1242,N_1640);
nand U3288 (N_3288,N_839,N_464);
xnor U3289 (N_3289,N_1414,N_609);
nor U3290 (N_3290,N_1387,N_404);
xnor U3291 (N_3291,N_1767,N_140);
or U3292 (N_3292,N_394,N_722);
xor U3293 (N_3293,N_1782,N_1262);
xnor U3294 (N_3294,N_234,N_1158);
xor U3295 (N_3295,N_1369,N_1801);
or U3296 (N_3296,N_93,N_330);
nor U3297 (N_3297,N_428,N_1662);
and U3298 (N_3298,N_656,N_71);
xor U3299 (N_3299,N_1796,N_1819);
nor U3300 (N_3300,N_1964,N_1344);
nand U3301 (N_3301,N_947,N_1145);
and U3302 (N_3302,N_1058,N_1123);
nand U3303 (N_3303,N_247,N_447);
or U3304 (N_3304,N_993,N_1886);
or U3305 (N_3305,N_840,N_1322);
or U3306 (N_3306,N_1567,N_257);
nand U3307 (N_3307,N_1315,N_981);
xor U3308 (N_3308,N_1188,N_1927);
nor U3309 (N_3309,N_882,N_1280);
and U3310 (N_3310,N_63,N_797);
nor U3311 (N_3311,N_553,N_953);
and U3312 (N_3312,N_1271,N_1852);
nand U3313 (N_3313,N_96,N_768);
or U3314 (N_3314,N_1860,N_1609);
xor U3315 (N_3315,N_276,N_695);
nor U3316 (N_3316,N_1541,N_819);
or U3317 (N_3317,N_1788,N_1908);
nand U3318 (N_3318,N_1543,N_1150);
and U3319 (N_3319,N_162,N_198);
nor U3320 (N_3320,N_841,N_987);
nand U3321 (N_3321,N_308,N_1385);
or U3322 (N_3322,N_1391,N_949);
nand U3323 (N_3323,N_1417,N_1907);
nand U3324 (N_3324,N_1371,N_314);
xor U3325 (N_3325,N_233,N_1917);
nand U3326 (N_3326,N_383,N_1428);
nand U3327 (N_3327,N_3,N_1150);
or U3328 (N_3328,N_462,N_1081);
xor U3329 (N_3329,N_276,N_1800);
nand U3330 (N_3330,N_1987,N_1631);
or U3331 (N_3331,N_1866,N_590);
nand U3332 (N_3332,N_393,N_1489);
xnor U3333 (N_3333,N_397,N_470);
and U3334 (N_3334,N_1149,N_63);
or U3335 (N_3335,N_1395,N_1796);
nor U3336 (N_3336,N_1975,N_335);
nor U3337 (N_3337,N_171,N_1416);
or U3338 (N_3338,N_843,N_206);
xor U3339 (N_3339,N_1644,N_932);
or U3340 (N_3340,N_256,N_1764);
nor U3341 (N_3341,N_1299,N_227);
nor U3342 (N_3342,N_1776,N_618);
nor U3343 (N_3343,N_1383,N_933);
or U3344 (N_3344,N_729,N_80);
xnor U3345 (N_3345,N_497,N_943);
nand U3346 (N_3346,N_850,N_1314);
nor U3347 (N_3347,N_1648,N_1824);
xor U3348 (N_3348,N_1092,N_813);
xnor U3349 (N_3349,N_1451,N_1911);
nand U3350 (N_3350,N_138,N_1948);
and U3351 (N_3351,N_878,N_1497);
and U3352 (N_3352,N_486,N_295);
or U3353 (N_3353,N_1754,N_1860);
xnor U3354 (N_3354,N_1743,N_597);
and U3355 (N_3355,N_1771,N_1364);
or U3356 (N_3356,N_486,N_1533);
or U3357 (N_3357,N_1872,N_561);
nor U3358 (N_3358,N_14,N_522);
or U3359 (N_3359,N_23,N_268);
nand U3360 (N_3360,N_102,N_137);
nand U3361 (N_3361,N_27,N_1086);
nor U3362 (N_3362,N_1534,N_802);
nor U3363 (N_3363,N_1555,N_206);
or U3364 (N_3364,N_524,N_996);
nor U3365 (N_3365,N_1975,N_550);
and U3366 (N_3366,N_1998,N_287);
nor U3367 (N_3367,N_628,N_548);
nor U3368 (N_3368,N_320,N_303);
and U3369 (N_3369,N_1767,N_1522);
nand U3370 (N_3370,N_220,N_1720);
nand U3371 (N_3371,N_1398,N_1199);
and U3372 (N_3372,N_1247,N_1779);
or U3373 (N_3373,N_1199,N_1030);
and U3374 (N_3374,N_1765,N_896);
or U3375 (N_3375,N_906,N_706);
and U3376 (N_3376,N_1054,N_1872);
nor U3377 (N_3377,N_810,N_210);
nand U3378 (N_3378,N_264,N_1811);
nor U3379 (N_3379,N_151,N_850);
nand U3380 (N_3380,N_19,N_685);
nand U3381 (N_3381,N_971,N_345);
nor U3382 (N_3382,N_823,N_1914);
nand U3383 (N_3383,N_1172,N_1012);
nor U3384 (N_3384,N_733,N_323);
nor U3385 (N_3385,N_1335,N_1382);
nand U3386 (N_3386,N_1744,N_14);
and U3387 (N_3387,N_1930,N_1663);
or U3388 (N_3388,N_810,N_350);
and U3389 (N_3389,N_1468,N_1156);
and U3390 (N_3390,N_894,N_322);
xnor U3391 (N_3391,N_794,N_928);
nand U3392 (N_3392,N_35,N_717);
or U3393 (N_3393,N_577,N_1669);
and U3394 (N_3394,N_1752,N_312);
nand U3395 (N_3395,N_392,N_146);
and U3396 (N_3396,N_780,N_104);
or U3397 (N_3397,N_708,N_1970);
or U3398 (N_3398,N_1992,N_332);
nor U3399 (N_3399,N_722,N_974);
nor U3400 (N_3400,N_1823,N_1373);
nor U3401 (N_3401,N_1804,N_189);
nand U3402 (N_3402,N_1749,N_318);
nor U3403 (N_3403,N_1623,N_1758);
or U3404 (N_3404,N_150,N_1886);
and U3405 (N_3405,N_648,N_1436);
nand U3406 (N_3406,N_747,N_1860);
nor U3407 (N_3407,N_776,N_38);
nand U3408 (N_3408,N_1657,N_244);
and U3409 (N_3409,N_1879,N_1244);
nor U3410 (N_3410,N_1809,N_978);
and U3411 (N_3411,N_1762,N_1220);
xor U3412 (N_3412,N_1443,N_49);
or U3413 (N_3413,N_1497,N_906);
nor U3414 (N_3414,N_1131,N_1163);
xnor U3415 (N_3415,N_755,N_896);
nand U3416 (N_3416,N_1880,N_1902);
or U3417 (N_3417,N_1378,N_358);
or U3418 (N_3418,N_4,N_1680);
xor U3419 (N_3419,N_1074,N_1649);
nand U3420 (N_3420,N_1112,N_1022);
and U3421 (N_3421,N_1876,N_1611);
nand U3422 (N_3422,N_1697,N_791);
or U3423 (N_3423,N_714,N_174);
nor U3424 (N_3424,N_1662,N_1119);
xnor U3425 (N_3425,N_1767,N_48);
nand U3426 (N_3426,N_356,N_233);
nand U3427 (N_3427,N_65,N_948);
xnor U3428 (N_3428,N_1057,N_1417);
nand U3429 (N_3429,N_424,N_848);
xnor U3430 (N_3430,N_206,N_683);
xnor U3431 (N_3431,N_989,N_543);
nor U3432 (N_3432,N_649,N_839);
and U3433 (N_3433,N_375,N_30);
nor U3434 (N_3434,N_937,N_295);
nand U3435 (N_3435,N_458,N_783);
nand U3436 (N_3436,N_995,N_624);
nor U3437 (N_3437,N_875,N_492);
nand U3438 (N_3438,N_1929,N_1892);
and U3439 (N_3439,N_638,N_1182);
nor U3440 (N_3440,N_181,N_977);
and U3441 (N_3441,N_1019,N_1263);
and U3442 (N_3442,N_469,N_261);
or U3443 (N_3443,N_547,N_1053);
nor U3444 (N_3444,N_647,N_1504);
nand U3445 (N_3445,N_331,N_129);
and U3446 (N_3446,N_1453,N_717);
or U3447 (N_3447,N_1324,N_1699);
nor U3448 (N_3448,N_1168,N_1051);
xor U3449 (N_3449,N_63,N_568);
xor U3450 (N_3450,N_939,N_126);
or U3451 (N_3451,N_1683,N_101);
nand U3452 (N_3452,N_604,N_1120);
xnor U3453 (N_3453,N_190,N_508);
and U3454 (N_3454,N_1676,N_522);
xnor U3455 (N_3455,N_755,N_1798);
nand U3456 (N_3456,N_355,N_1432);
and U3457 (N_3457,N_531,N_1748);
or U3458 (N_3458,N_1333,N_1717);
xnor U3459 (N_3459,N_409,N_861);
or U3460 (N_3460,N_1799,N_1383);
and U3461 (N_3461,N_851,N_1532);
nand U3462 (N_3462,N_1083,N_771);
nand U3463 (N_3463,N_268,N_1020);
or U3464 (N_3464,N_946,N_1653);
and U3465 (N_3465,N_154,N_405);
and U3466 (N_3466,N_258,N_721);
or U3467 (N_3467,N_1011,N_1391);
xnor U3468 (N_3468,N_342,N_702);
nand U3469 (N_3469,N_1108,N_6);
or U3470 (N_3470,N_1341,N_547);
and U3471 (N_3471,N_1468,N_415);
nor U3472 (N_3472,N_1765,N_1716);
xnor U3473 (N_3473,N_1777,N_41);
or U3474 (N_3474,N_699,N_10);
or U3475 (N_3475,N_612,N_1707);
nand U3476 (N_3476,N_1369,N_706);
or U3477 (N_3477,N_12,N_258);
xor U3478 (N_3478,N_129,N_376);
and U3479 (N_3479,N_1232,N_1743);
nor U3480 (N_3480,N_568,N_433);
nor U3481 (N_3481,N_1587,N_1788);
or U3482 (N_3482,N_606,N_411);
and U3483 (N_3483,N_1773,N_316);
xor U3484 (N_3484,N_1636,N_309);
xnor U3485 (N_3485,N_1040,N_281);
nor U3486 (N_3486,N_1298,N_596);
and U3487 (N_3487,N_333,N_1920);
or U3488 (N_3488,N_1087,N_1247);
nand U3489 (N_3489,N_136,N_1298);
nor U3490 (N_3490,N_1831,N_182);
nand U3491 (N_3491,N_528,N_944);
nand U3492 (N_3492,N_1232,N_605);
xor U3493 (N_3493,N_121,N_1912);
nor U3494 (N_3494,N_1733,N_1857);
or U3495 (N_3495,N_235,N_1586);
xor U3496 (N_3496,N_532,N_779);
nand U3497 (N_3497,N_1807,N_648);
and U3498 (N_3498,N_791,N_802);
nand U3499 (N_3499,N_1184,N_1303);
or U3500 (N_3500,N_877,N_1461);
or U3501 (N_3501,N_1601,N_1038);
nor U3502 (N_3502,N_1042,N_465);
nand U3503 (N_3503,N_1410,N_94);
nor U3504 (N_3504,N_1758,N_553);
nor U3505 (N_3505,N_1288,N_1169);
xor U3506 (N_3506,N_1606,N_1892);
nor U3507 (N_3507,N_76,N_1501);
xnor U3508 (N_3508,N_481,N_274);
or U3509 (N_3509,N_701,N_1074);
and U3510 (N_3510,N_1297,N_623);
nor U3511 (N_3511,N_1317,N_276);
nor U3512 (N_3512,N_116,N_341);
or U3513 (N_3513,N_1903,N_137);
or U3514 (N_3514,N_1502,N_810);
and U3515 (N_3515,N_1804,N_70);
nand U3516 (N_3516,N_1547,N_1739);
nand U3517 (N_3517,N_737,N_1438);
and U3518 (N_3518,N_387,N_1450);
xor U3519 (N_3519,N_412,N_1751);
or U3520 (N_3520,N_687,N_1285);
xor U3521 (N_3521,N_450,N_829);
nand U3522 (N_3522,N_1957,N_824);
nand U3523 (N_3523,N_945,N_1933);
nor U3524 (N_3524,N_1502,N_1821);
nand U3525 (N_3525,N_635,N_1861);
or U3526 (N_3526,N_428,N_1996);
nand U3527 (N_3527,N_344,N_1862);
nand U3528 (N_3528,N_1642,N_788);
and U3529 (N_3529,N_889,N_1638);
and U3530 (N_3530,N_1038,N_1957);
or U3531 (N_3531,N_296,N_115);
and U3532 (N_3532,N_477,N_402);
nor U3533 (N_3533,N_219,N_1418);
or U3534 (N_3534,N_1589,N_1634);
nor U3535 (N_3535,N_1139,N_351);
nand U3536 (N_3536,N_660,N_238);
or U3537 (N_3537,N_1170,N_650);
xnor U3538 (N_3538,N_875,N_1638);
and U3539 (N_3539,N_1212,N_391);
nand U3540 (N_3540,N_1341,N_1844);
nand U3541 (N_3541,N_1626,N_1937);
nor U3542 (N_3542,N_1943,N_530);
and U3543 (N_3543,N_558,N_74);
and U3544 (N_3544,N_12,N_172);
xor U3545 (N_3545,N_509,N_442);
and U3546 (N_3546,N_1911,N_1616);
and U3547 (N_3547,N_844,N_380);
nand U3548 (N_3548,N_153,N_1742);
nand U3549 (N_3549,N_297,N_1249);
nand U3550 (N_3550,N_1302,N_368);
nand U3551 (N_3551,N_393,N_1024);
nor U3552 (N_3552,N_786,N_90);
and U3553 (N_3553,N_999,N_1184);
nor U3554 (N_3554,N_1347,N_81);
and U3555 (N_3555,N_737,N_855);
or U3556 (N_3556,N_335,N_317);
nand U3557 (N_3557,N_1782,N_984);
nor U3558 (N_3558,N_1437,N_890);
and U3559 (N_3559,N_841,N_210);
or U3560 (N_3560,N_170,N_518);
or U3561 (N_3561,N_59,N_1888);
and U3562 (N_3562,N_1176,N_363);
xor U3563 (N_3563,N_1912,N_1071);
or U3564 (N_3564,N_647,N_1726);
nor U3565 (N_3565,N_1838,N_433);
xnor U3566 (N_3566,N_1488,N_1575);
and U3567 (N_3567,N_1697,N_1972);
and U3568 (N_3568,N_371,N_1505);
nand U3569 (N_3569,N_422,N_1324);
or U3570 (N_3570,N_172,N_1910);
nand U3571 (N_3571,N_1306,N_665);
or U3572 (N_3572,N_1293,N_272);
nand U3573 (N_3573,N_1801,N_1491);
xor U3574 (N_3574,N_1006,N_693);
or U3575 (N_3575,N_918,N_1851);
xnor U3576 (N_3576,N_1000,N_813);
and U3577 (N_3577,N_484,N_1007);
xnor U3578 (N_3578,N_1827,N_1420);
or U3579 (N_3579,N_319,N_1627);
nor U3580 (N_3580,N_561,N_1916);
xnor U3581 (N_3581,N_448,N_1297);
and U3582 (N_3582,N_1629,N_781);
and U3583 (N_3583,N_340,N_1290);
nand U3584 (N_3584,N_1209,N_792);
nor U3585 (N_3585,N_1894,N_242);
nand U3586 (N_3586,N_1753,N_665);
xor U3587 (N_3587,N_1579,N_43);
or U3588 (N_3588,N_298,N_529);
nor U3589 (N_3589,N_458,N_514);
nand U3590 (N_3590,N_289,N_1416);
or U3591 (N_3591,N_1500,N_142);
and U3592 (N_3592,N_1846,N_486);
nand U3593 (N_3593,N_1236,N_1753);
xor U3594 (N_3594,N_810,N_1953);
and U3595 (N_3595,N_273,N_1909);
nand U3596 (N_3596,N_938,N_1888);
or U3597 (N_3597,N_67,N_717);
nand U3598 (N_3598,N_706,N_885);
nor U3599 (N_3599,N_1435,N_1365);
or U3600 (N_3600,N_1077,N_636);
xnor U3601 (N_3601,N_1055,N_119);
and U3602 (N_3602,N_434,N_394);
nor U3603 (N_3603,N_961,N_264);
xor U3604 (N_3604,N_1739,N_1452);
or U3605 (N_3605,N_1535,N_1581);
xnor U3606 (N_3606,N_1875,N_1974);
or U3607 (N_3607,N_962,N_1477);
xnor U3608 (N_3608,N_547,N_1367);
and U3609 (N_3609,N_1583,N_1975);
nand U3610 (N_3610,N_760,N_1887);
nor U3611 (N_3611,N_1709,N_1164);
xnor U3612 (N_3612,N_1806,N_473);
nand U3613 (N_3613,N_1484,N_8);
nand U3614 (N_3614,N_1010,N_341);
and U3615 (N_3615,N_176,N_1380);
or U3616 (N_3616,N_1401,N_238);
and U3617 (N_3617,N_1763,N_1453);
nand U3618 (N_3618,N_573,N_1030);
nand U3619 (N_3619,N_385,N_1896);
nand U3620 (N_3620,N_1294,N_205);
and U3621 (N_3621,N_381,N_606);
xnor U3622 (N_3622,N_1508,N_1240);
and U3623 (N_3623,N_984,N_1819);
nor U3624 (N_3624,N_101,N_1541);
xor U3625 (N_3625,N_545,N_1554);
xnor U3626 (N_3626,N_394,N_1049);
or U3627 (N_3627,N_411,N_810);
nor U3628 (N_3628,N_220,N_710);
and U3629 (N_3629,N_596,N_820);
and U3630 (N_3630,N_1033,N_819);
xnor U3631 (N_3631,N_567,N_20);
or U3632 (N_3632,N_974,N_767);
or U3633 (N_3633,N_262,N_720);
and U3634 (N_3634,N_691,N_1306);
or U3635 (N_3635,N_317,N_1057);
and U3636 (N_3636,N_1267,N_941);
nor U3637 (N_3637,N_530,N_218);
and U3638 (N_3638,N_865,N_1819);
nor U3639 (N_3639,N_294,N_1720);
nor U3640 (N_3640,N_48,N_1453);
or U3641 (N_3641,N_20,N_1114);
nor U3642 (N_3642,N_257,N_396);
nor U3643 (N_3643,N_1496,N_915);
nand U3644 (N_3644,N_1094,N_1148);
or U3645 (N_3645,N_1574,N_1065);
and U3646 (N_3646,N_210,N_447);
and U3647 (N_3647,N_974,N_102);
nor U3648 (N_3648,N_117,N_667);
and U3649 (N_3649,N_1232,N_334);
and U3650 (N_3650,N_1579,N_1671);
and U3651 (N_3651,N_1881,N_859);
nor U3652 (N_3652,N_112,N_343);
nand U3653 (N_3653,N_176,N_1483);
nand U3654 (N_3654,N_1236,N_561);
nor U3655 (N_3655,N_1088,N_590);
xnor U3656 (N_3656,N_1190,N_722);
and U3657 (N_3657,N_1981,N_1220);
and U3658 (N_3658,N_1498,N_588);
nor U3659 (N_3659,N_1103,N_29);
xnor U3660 (N_3660,N_67,N_200);
or U3661 (N_3661,N_342,N_1448);
nand U3662 (N_3662,N_1901,N_266);
nor U3663 (N_3663,N_96,N_521);
nand U3664 (N_3664,N_1673,N_848);
nor U3665 (N_3665,N_1515,N_1963);
or U3666 (N_3666,N_1670,N_990);
xor U3667 (N_3667,N_1575,N_1342);
nor U3668 (N_3668,N_901,N_1278);
xnor U3669 (N_3669,N_904,N_720);
nor U3670 (N_3670,N_1742,N_1818);
xor U3671 (N_3671,N_791,N_877);
nand U3672 (N_3672,N_256,N_1048);
xor U3673 (N_3673,N_271,N_803);
or U3674 (N_3674,N_585,N_624);
nand U3675 (N_3675,N_1793,N_1407);
and U3676 (N_3676,N_1332,N_1252);
or U3677 (N_3677,N_387,N_548);
nor U3678 (N_3678,N_995,N_1626);
nand U3679 (N_3679,N_783,N_0);
nand U3680 (N_3680,N_1836,N_1424);
nor U3681 (N_3681,N_254,N_1669);
nand U3682 (N_3682,N_1342,N_835);
and U3683 (N_3683,N_563,N_774);
or U3684 (N_3684,N_716,N_1739);
or U3685 (N_3685,N_115,N_613);
xnor U3686 (N_3686,N_889,N_725);
and U3687 (N_3687,N_941,N_993);
or U3688 (N_3688,N_1239,N_1445);
and U3689 (N_3689,N_791,N_408);
or U3690 (N_3690,N_446,N_1678);
nand U3691 (N_3691,N_1890,N_156);
or U3692 (N_3692,N_1244,N_862);
or U3693 (N_3693,N_1966,N_1863);
nor U3694 (N_3694,N_339,N_369);
and U3695 (N_3695,N_43,N_1778);
nand U3696 (N_3696,N_1967,N_946);
nor U3697 (N_3697,N_968,N_1622);
nand U3698 (N_3698,N_134,N_1032);
or U3699 (N_3699,N_324,N_1196);
nor U3700 (N_3700,N_697,N_18);
or U3701 (N_3701,N_505,N_479);
nor U3702 (N_3702,N_205,N_9);
nor U3703 (N_3703,N_1929,N_336);
xor U3704 (N_3704,N_1406,N_1951);
xor U3705 (N_3705,N_1414,N_1147);
nor U3706 (N_3706,N_1403,N_1607);
and U3707 (N_3707,N_1821,N_682);
nand U3708 (N_3708,N_1995,N_670);
and U3709 (N_3709,N_1216,N_567);
nand U3710 (N_3710,N_1750,N_1113);
and U3711 (N_3711,N_229,N_1543);
and U3712 (N_3712,N_283,N_642);
nand U3713 (N_3713,N_425,N_409);
xor U3714 (N_3714,N_263,N_916);
xnor U3715 (N_3715,N_346,N_1456);
and U3716 (N_3716,N_1032,N_838);
and U3717 (N_3717,N_1327,N_334);
nand U3718 (N_3718,N_1887,N_1241);
or U3719 (N_3719,N_1161,N_837);
nor U3720 (N_3720,N_1932,N_334);
nand U3721 (N_3721,N_1225,N_1901);
nor U3722 (N_3722,N_1957,N_1936);
and U3723 (N_3723,N_575,N_1162);
xnor U3724 (N_3724,N_1228,N_1001);
or U3725 (N_3725,N_1917,N_1717);
or U3726 (N_3726,N_528,N_1030);
xnor U3727 (N_3727,N_631,N_263);
and U3728 (N_3728,N_1857,N_1600);
nor U3729 (N_3729,N_1235,N_298);
xor U3730 (N_3730,N_443,N_702);
xnor U3731 (N_3731,N_1930,N_1807);
and U3732 (N_3732,N_638,N_967);
and U3733 (N_3733,N_960,N_1762);
and U3734 (N_3734,N_1080,N_452);
and U3735 (N_3735,N_224,N_539);
nand U3736 (N_3736,N_267,N_1691);
and U3737 (N_3737,N_1396,N_174);
xor U3738 (N_3738,N_578,N_434);
xor U3739 (N_3739,N_685,N_425);
or U3740 (N_3740,N_1886,N_755);
and U3741 (N_3741,N_885,N_585);
or U3742 (N_3742,N_160,N_1032);
or U3743 (N_3743,N_1490,N_435);
and U3744 (N_3744,N_902,N_736);
and U3745 (N_3745,N_1999,N_706);
nor U3746 (N_3746,N_1852,N_786);
nor U3747 (N_3747,N_1386,N_1580);
or U3748 (N_3748,N_1302,N_1705);
xnor U3749 (N_3749,N_258,N_195);
and U3750 (N_3750,N_45,N_1773);
and U3751 (N_3751,N_1202,N_1369);
xor U3752 (N_3752,N_566,N_183);
or U3753 (N_3753,N_1305,N_1533);
nor U3754 (N_3754,N_17,N_864);
nor U3755 (N_3755,N_794,N_1005);
xnor U3756 (N_3756,N_1229,N_603);
xnor U3757 (N_3757,N_900,N_1119);
and U3758 (N_3758,N_211,N_1989);
or U3759 (N_3759,N_408,N_1617);
and U3760 (N_3760,N_302,N_1857);
and U3761 (N_3761,N_592,N_952);
xor U3762 (N_3762,N_720,N_1310);
xor U3763 (N_3763,N_318,N_1589);
nor U3764 (N_3764,N_752,N_516);
nand U3765 (N_3765,N_1906,N_1367);
and U3766 (N_3766,N_1908,N_1697);
or U3767 (N_3767,N_354,N_1648);
nor U3768 (N_3768,N_1787,N_331);
nand U3769 (N_3769,N_1890,N_1429);
nand U3770 (N_3770,N_792,N_1793);
xor U3771 (N_3771,N_1210,N_1154);
and U3772 (N_3772,N_1698,N_1537);
or U3773 (N_3773,N_1491,N_563);
and U3774 (N_3774,N_173,N_789);
and U3775 (N_3775,N_1639,N_1964);
nand U3776 (N_3776,N_1582,N_1189);
nand U3777 (N_3777,N_805,N_1664);
nand U3778 (N_3778,N_1514,N_316);
and U3779 (N_3779,N_309,N_502);
xnor U3780 (N_3780,N_1280,N_1902);
or U3781 (N_3781,N_1288,N_1782);
or U3782 (N_3782,N_1030,N_918);
or U3783 (N_3783,N_1919,N_809);
and U3784 (N_3784,N_534,N_1259);
nor U3785 (N_3785,N_1089,N_793);
nor U3786 (N_3786,N_773,N_1662);
nand U3787 (N_3787,N_662,N_1916);
and U3788 (N_3788,N_1977,N_872);
xnor U3789 (N_3789,N_616,N_625);
nand U3790 (N_3790,N_1510,N_1214);
nand U3791 (N_3791,N_65,N_1576);
nand U3792 (N_3792,N_592,N_1585);
or U3793 (N_3793,N_1585,N_68);
and U3794 (N_3794,N_1085,N_1622);
nor U3795 (N_3795,N_936,N_1872);
xnor U3796 (N_3796,N_1187,N_1402);
and U3797 (N_3797,N_1441,N_1492);
or U3798 (N_3798,N_1958,N_825);
and U3799 (N_3799,N_622,N_492);
nand U3800 (N_3800,N_232,N_147);
or U3801 (N_3801,N_257,N_1459);
nor U3802 (N_3802,N_71,N_1893);
nand U3803 (N_3803,N_1367,N_704);
nand U3804 (N_3804,N_1184,N_740);
nand U3805 (N_3805,N_748,N_1054);
and U3806 (N_3806,N_901,N_1450);
and U3807 (N_3807,N_255,N_646);
nor U3808 (N_3808,N_1130,N_1036);
xor U3809 (N_3809,N_158,N_1675);
and U3810 (N_3810,N_1501,N_1677);
and U3811 (N_3811,N_724,N_162);
xnor U3812 (N_3812,N_1042,N_1977);
xor U3813 (N_3813,N_1935,N_1821);
and U3814 (N_3814,N_1788,N_1581);
xor U3815 (N_3815,N_246,N_723);
or U3816 (N_3816,N_782,N_1401);
nand U3817 (N_3817,N_510,N_1790);
nand U3818 (N_3818,N_1779,N_1175);
nor U3819 (N_3819,N_1829,N_764);
or U3820 (N_3820,N_1808,N_210);
nor U3821 (N_3821,N_75,N_1332);
nand U3822 (N_3822,N_689,N_1603);
and U3823 (N_3823,N_650,N_421);
or U3824 (N_3824,N_599,N_810);
nand U3825 (N_3825,N_1868,N_1450);
nor U3826 (N_3826,N_1804,N_34);
or U3827 (N_3827,N_376,N_974);
nor U3828 (N_3828,N_1788,N_511);
and U3829 (N_3829,N_675,N_1765);
and U3830 (N_3830,N_647,N_688);
or U3831 (N_3831,N_330,N_1377);
nand U3832 (N_3832,N_1486,N_508);
xnor U3833 (N_3833,N_605,N_921);
nor U3834 (N_3834,N_1792,N_881);
nand U3835 (N_3835,N_1974,N_241);
and U3836 (N_3836,N_1144,N_934);
nand U3837 (N_3837,N_1396,N_87);
nor U3838 (N_3838,N_162,N_1249);
or U3839 (N_3839,N_250,N_29);
or U3840 (N_3840,N_238,N_1476);
or U3841 (N_3841,N_1545,N_713);
nor U3842 (N_3842,N_504,N_1404);
nand U3843 (N_3843,N_1677,N_1390);
xor U3844 (N_3844,N_1407,N_1833);
or U3845 (N_3845,N_1702,N_1080);
nor U3846 (N_3846,N_935,N_302);
nand U3847 (N_3847,N_120,N_1187);
or U3848 (N_3848,N_700,N_730);
nor U3849 (N_3849,N_1009,N_1807);
and U3850 (N_3850,N_109,N_353);
nand U3851 (N_3851,N_368,N_1890);
or U3852 (N_3852,N_1823,N_82);
or U3853 (N_3853,N_366,N_922);
nand U3854 (N_3854,N_1271,N_878);
xnor U3855 (N_3855,N_41,N_1739);
nand U3856 (N_3856,N_1364,N_53);
nand U3857 (N_3857,N_908,N_366);
and U3858 (N_3858,N_778,N_424);
nor U3859 (N_3859,N_1883,N_783);
and U3860 (N_3860,N_946,N_1234);
nor U3861 (N_3861,N_306,N_815);
nand U3862 (N_3862,N_436,N_1634);
xor U3863 (N_3863,N_1288,N_584);
and U3864 (N_3864,N_1137,N_1172);
or U3865 (N_3865,N_1628,N_1061);
or U3866 (N_3866,N_1502,N_1399);
or U3867 (N_3867,N_1733,N_234);
or U3868 (N_3868,N_1824,N_243);
or U3869 (N_3869,N_894,N_1454);
nand U3870 (N_3870,N_805,N_41);
nor U3871 (N_3871,N_837,N_1334);
nand U3872 (N_3872,N_1082,N_71);
nand U3873 (N_3873,N_1016,N_210);
and U3874 (N_3874,N_1670,N_404);
nor U3875 (N_3875,N_1457,N_1732);
nor U3876 (N_3876,N_758,N_1511);
and U3877 (N_3877,N_569,N_1178);
nor U3878 (N_3878,N_34,N_862);
nor U3879 (N_3879,N_1483,N_1641);
nor U3880 (N_3880,N_1137,N_319);
nand U3881 (N_3881,N_224,N_310);
nor U3882 (N_3882,N_924,N_1282);
and U3883 (N_3883,N_1046,N_930);
nand U3884 (N_3884,N_1046,N_1736);
nand U3885 (N_3885,N_1308,N_474);
and U3886 (N_3886,N_1481,N_453);
and U3887 (N_3887,N_361,N_224);
or U3888 (N_3888,N_88,N_1863);
xor U3889 (N_3889,N_640,N_511);
or U3890 (N_3890,N_720,N_715);
or U3891 (N_3891,N_1530,N_1564);
or U3892 (N_3892,N_1721,N_432);
and U3893 (N_3893,N_1830,N_1966);
nand U3894 (N_3894,N_1162,N_1922);
nand U3895 (N_3895,N_1109,N_33);
nand U3896 (N_3896,N_466,N_1084);
xor U3897 (N_3897,N_154,N_1867);
and U3898 (N_3898,N_902,N_1947);
or U3899 (N_3899,N_1649,N_262);
nor U3900 (N_3900,N_1309,N_1841);
and U3901 (N_3901,N_1192,N_1758);
or U3902 (N_3902,N_956,N_489);
nor U3903 (N_3903,N_1499,N_1059);
or U3904 (N_3904,N_888,N_1355);
nor U3905 (N_3905,N_1378,N_958);
nand U3906 (N_3906,N_1298,N_427);
and U3907 (N_3907,N_1715,N_1294);
xnor U3908 (N_3908,N_1120,N_1149);
xor U3909 (N_3909,N_764,N_294);
nand U3910 (N_3910,N_678,N_735);
xor U3911 (N_3911,N_890,N_122);
or U3912 (N_3912,N_1513,N_247);
nand U3913 (N_3913,N_1427,N_1623);
nand U3914 (N_3914,N_364,N_1468);
nand U3915 (N_3915,N_1583,N_1829);
and U3916 (N_3916,N_796,N_736);
or U3917 (N_3917,N_626,N_1908);
nor U3918 (N_3918,N_937,N_1441);
nand U3919 (N_3919,N_1788,N_901);
or U3920 (N_3920,N_922,N_1015);
nand U3921 (N_3921,N_1011,N_486);
xor U3922 (N_3922,N_142,N_1884);
xor U3923 (N_3923,N_336,N_1940);
nor U3924 (N_3924,N_375,N_1599);
xnor U3925 (N_3925,N_456,N_1084);
xor U3926 (N_3926,N_1892,N_1894);
nand U3927 (N_3927,N_1847,N_483);
xnor U3928 (N_3928,N_637,N_1790);
xnor U3929 (N_3929,N_431,N_557);
and U3930 (N_3930,N_186,N_1401);
xnor U3931 (N_3931,N_1007,N_1170);
nor U3932 (N_3932,N_1965,N_457);
or U3933 (N_3933,N_944,N_364);
xnor U3934 (N_3934,N_1844,N_1240);
and U3935 (N_3935,N_60,N_1015);
or U3936 (N_3936,N_533,N_151);
and U3937 (N_3937,N_330,N_327);
xor U3938 (N_3938,N_399,N_663);
nand U3939 (N_3939,N_802,N_941);
or U3940 (N_3940,N_1191,N_1115);
xor U3941 (N_3941,N_1797,N_1176);
or U3942 (N_3942,N_277,N_1375);
nor U3943 (N_3943,N_1100,N_867);
nand U3944 (N_3944,N_1434,N_987);
nand U3945 (N_3945,N_1945,N_101);
and U3946 (N_3946,N_1925,N_1636);
xor U3947 (N_3947,N_75,N_545);
nand U3948 (N_3948,N_1049,N_1309);
or U3949 (N_3949,N_1330,N_69);
nand U3950 (N_3950,N_785,N_378);
or U3951 (N_3951,N_1154,N_190);
xor U3952 (N_3952,N_1835,N_1034);
or U3953 (N_3953,N_1865,N_981);
and U3954 (N_3954,N_1752,N_1270);
or U3955 (N_3955,N_726,N_21);
and U3956 (N_3956,N_488,N_917);
nor U3957 (N_3957,N_1555,N_1734);
nor U3958 (N_3958,N_824,N_1413);
and U3959 (N_3959,N_423,N_1866);
nand U3960 (N_3960,N_337,N_163);
nor U3961 (N_3961,N_1559,N_1143);
and U3962 (N_3962,N_1875,N_626);
xnor U3963 (N_3963,N_798,N_945);
nand U3964 (N_3964,N_1395,N_1123);
and U3965 (N_3965,N_1522,N_408);
and U3966 (N_3966,N_954,N_135);
xnor U3967 (N_3967,N_1518,N_1548);
or U3968 (N_3968,N_843,N_900);
or U3969 (N_3969,N_503,N_688);
xnor U3970 (N_3970,N_69,N_1251);
nor U3971 (N_3971,N_367,N_1225);
nor U3972 (N_3972,N_1745,N_1638);
or U3973 (N_3973,N_949,N_1473);
nand U3974 (N_3974,N_1066,N_920);
or U3975 (N_3975,N_1682,N_1042);
or U3976 (N_3976,N_75,N_122);
and U3977 (N_3977,N_1064,N_531);
xnor U3978 (N_3978,N_861,N_1298);
nand U3979 (N_3979,N_463,N_129);
nor U3980 (N_3980,N_898,N_717);
nor U3981 (N_3981,N_1232,N_133);
or U3982 (N_3982,N_1678,N_1846);
or U3983 (N_3983,N_30,N_1447);
nor U3984 (N_3984,N_723,N_761);
nor U3985 (N_3985,N_1032,N_1304);
nor U3986 (N_3986,N_1500,N_1995);
nand U3987 (N_3987,N_633,N_1073);
nand U3988 (N_3988,N_968,N_1190);
or U3989 (N_3989,N_1084,N_832);
nor U3990 (N_3990,N_480,N_356);
or U3991 (N_3991,N_1329,N_657);
or U3992 (N_3992,N_1283,N_1912);
xor U3993 (N_3993,N_1127,N_376);
or U3994 (N_3994,N_1225,N_1030);
and U3995 (N_3995,N_160,N_1683);
nor U3996 (N_3996,N_1444,N_752);
or U3997 (N_3997,N_1049,N_1832);
and U3998 (N_3998,N_1618,N_316);
and U3999 (N_3999,N_225,N_143);
or U4000 (N_4000,N_3597,N_3836);
nand U4001 (N_4001,N_3057,N_2584);
and U4002 (N_4002,N_3481,N_2239);
xor U4003 (N_4003,N_2296,N_3530);
nand U4004 (N_4004,N_3652,N_3326);
nand U4005 (N_4005,N_3152,N_3332);
nor U4006 (N_4006,N_3479,N_3825);
or U4007 (N_4007,N_3934,N_3684);
nand U4008 (N_4008,N_3919,N_3991);
nand U4009 (N_4009,N_2339,N_3519);
xnor U4010 (N_4010,N_2400,N_3942);
nor U4011 (N_4011,N_2777,N_2042);
xnor U4012 (N_4012,N_3715,N_2513);
xnor U4013 (N_4013,N_3722,N_3370);
and U4014 (N_4014,N_3429,N_3513);
xnor U4015 (N_4015,N_2890,N_2717);
nor U4016 (N_4016,N_2333,N_2297);
nor U4017 (N_4017,N_2149,N_3309);
nor U4018 (N_4018,N_3443,N_3685);
or U4019 (N_4019,N_2520,N_2194);
xor U4020 (N_4020,N_3725,N_3394);
nor U4021 (N_4021,N_2989,N_3639);
nor U4022 (N_4022,N_3829,N_2528);
xnor U4023 (N_4023,N_3213,N_2082);
nor U4024 (N_4024,N_3780,N_2656);
and U4025 (N_4025,N_2269,N_3924);
nand U4026 (N_4026,N_2228,N_3763);
or U4027 (N_4027,N_3195,N_3745);
xor U4028 (N_4028,N_3683,N_2608);
and U4029 (N_4029,N_2443,N_2594);
xnor U4030 (N_4030,N_3839,N_2801);
and U4031 (N_4031,N_3871,N_2576);
nor U4032 (N_4032,N_3704,N_2694);
or U4033 (N_4033,N_2848,N_3436);
or U4034 (N_4034,N_2366,N_2639);
nand U4035 (N_4035,N_2325,N_2776);
nor U4036 (N_4036,N_3746,N_2447);
nor U4037 (N_4037,N_3385,N_3830);
nand U4038 (N_4038,N_3622,N_3552);
nand U4039 (N_4039,N_3322,N_2987);
or U4040 (N_4040,N_3150,N_3849);
nand U4041 (N_4041,N_3800,N_2713);
nand U4042 (N_4042,N_2671,N_3637);
and U4043 (N_4043,N_3783,N_2986);
xnor U4044 (N_4044,N_2460,N_2940);
nand U4045 (N_4045,N_2346,N_2953);
and U4046 (N_4046,N_3252,N_2845);
or U4047 (N_4047,N_2309,N_2392);
and U4048 (N_4048,N_2418,N_3705);
nand U4049 (N_4049,N_3787,N_3416);
nand U4050 (N_4050,N_2234,N_2591);
nand U4051 (N_4051,N_3936,N_2062);
xnor U4052 (N_4052,N_3040,N_2032);
xnor U4053 (N_4053,N_2053,N_3419);
xor U4054 (N_4054,N_2078,N_3165);
xnor U4055 (N_4055,N_2287,N_3231);
or U4056 (N_4056,N_3188,N_2756);
or U4057 (N_4057,N_3382,N_3145);
xor U4058 (N_4058,N_3903,N_2859);
and U4059 (N_4059,N_2273,N_3857);
nand U4060 (N_4060,N_2831,N_2626);
xor U4061 (N_4061,N_2722,N_2715);
or U4062 (N_4062,N_3992,N_3233);
nand U4063 (N_4063,N_2841,N_2498);
or U4064 (N_4064,N_2470,N_3721);
and U4065 (N_4065,N_2539,N_2634);
nor U4066 (N_4066,N_2616,N_2484);
xor U4067 (N_4067,N_3888,N_3592);
nand U4068 (N_4068,N_3403,N_2463);
nand U4069 (N_4069,N_3617,N_2988);
nand U4070 (N_4070,N_3525,N_2266);
or U4071 (N_4071,N_3372,N_3182);
nand U4072 (N_4072,N_3041,N_2678);
or U4073 (N_4073,N_3455,N_2261);
or U4074 (N_4074,N_2969,N_3067);
nand U4075 (N_4075,N_2727,N_3889);
xor U4076 (N_4076,N_2453,N_2882);
nand U4077 (N_4077,N_2633,N_3036);
nor U4078 (N_4078,N_3980,N_3906);
nor U4079 (N_4079,N_3744,N_3535);
or U4080 (N_4080,N_3444,N_3719);
and U4081 (N_4081,N_2057,N_3316);
or U4082 (N_4082,N_3155,N_3069);
nor U4083 (N_4083,N_3944,N_2832);
xor U4084 (N_4084,N_3472,N_3303);
xnor U4085 (N_4085,N_2945,N_2721);
nor U4086 (N_4086,N_3365,N_3350);
xor U4087 (N_4087,N_3131,N_3738);
nor U4088 (N_4088,N_2157,N_3566);
or U4089 (N_4089,N_3373,N_2290);
nand U4090 (N_4090,N_2322,N_2701);
xnor U4091 (N_4091,N_3549,N_2730);
nand U4092 (N_4092,N_3494,N_3771);
nand U4093 (N_4093,N_3272,N_3070);
or U4094 (N_4094,N_2427,N_2462);
or U4095 (N_4095,N_3124,N_2654);
xor U4096 (N_4096,N_2536,N_2564);
nor U4097 (N_4097,N_3461,N_2158);
nand U4098 (N_4098,N_3968,N_3263);
nor U4099 (N_4099,N_2302,N_3022);
and U4100 (N_4100,N_3136,N_2016);
nand U4101 (N_4101,N_3805,N_2080);
nand U4102 (N_4102,N_2898,N_3969);
or U4103 (N_4103,N_2792,N_3709);
or U4104 (N_4104,N_2294,N_2972);
xor U4105 (N_4105,N_3895,N_3603);
xnor U4106 (N_4106,N_2330,N_2155);
nor U4107 (N_4107,N_2272,N_3890);
and U4108 (N_4108,N_2546,N_3079);
and U4109 (N_4109,N_2123,N_3467);
nand U4110 (N_4110,N_2602,N_2203);
and U4111 (N_4111,N_3009,N_2214);
or U4112 (N_4112,N_3623,N_3295);
nand U4113 (N_4113,N_2120,N_3961);
and U4114 (N_4114,N_3585,N_3445);
nand U4115 (N_4115,N_3669,N_3062);
or U4116 (N_4116,N_3514,N_2128);
or U4117 (N_4117,N_2110,N_2686);
xnor U4118 (N_4118,N_3790,N_3016);
or U4119 (N_4119,N_3014,N_3453);
and U4120 (N_4120,N_2387,N_3024);
xnor U4121 (N_4121,N_3293,N_3851);
nand U4122 (N_4122,N_3077,N_3149);
and U4123 (N_4123,N_2581,N_2775);
nand U4124 (N_4124,N_3522,N_2599);
or U4125 (N_4125,N_2574,N_3580);
nand U4126 (N_4126,N_3651,N_2950);
or U4127 (N_4127,N_2213,N_3562);
nand U4128 (N_4128,N_2965,N_3607);
nand U4129 (N_4129,N_2535,N_3733);
nor U4130 (N_4130,N_2049,N_2517);
or U4131 (N_4131,N_2191,N_3879);
or U4132 (N_4132,N_2852,N_2063);
xor U4133 (N_4133,N_3806,N_3846);
xor U4134 (N_4134,N_2352,N_2838);
nand U4135 (N_4135,N_2856,N_3135);
or U4136 (N_4136,N_2824,N_2136);
xor U4137 (N_4137,N_2122,N_3858);
nand U4138 (N_4138,N_2625,N_2834);
nor U4139 (N_4139,N_2970,N_2225);
or U4140 (N_4140,N_2642,N_3031);
and U4141 (N_4141,N_2005,N_2797);
and U4142 (N_4142,N_2281,N_2098);
nand U4143 (N_4143,N_2631,N_2148);
nand U4144 (N_4144,N_3731,N_3670);
and U4145 (N_4145,N_2091,N_2764);
nand U4146 (N_4146,N_2014,N_3624);
and U4147 (N_4147,N_2087,N_2647);
or U4148 (N_4148,N_2251,N_2344);
and U4149 (N_4149,N_2610,N_2755);
nor U4150 (N_4150,N_3943,N_3119);
nand U4151 (N_4151,N_2304,N_3171);
xnor U4152 (N_4152,N_2026,N_3544);
xnor U4153 (N_4153,N_3812,N_2499);
and U4154 (N_4154,N_3557,N_2981);
and U4155 (N_4155,N_3250,N_2025);
or U4156 (N_4156,N_3986,N_2113);
and U4157 (N_4157,N_3325,N_2449);
nor U4158 (N_4158,N_3071,N_3672);
xor U4159 (N_4159,N_3276,N_2544);
and U4160 (N_4160,N_3772,N_3491);
nand U4161 (N_4161,N_3148,N_2402);
nand U4162 (N_4162,N_2936,N_3172);
xnor U4163 (N_4163,N_3635,N_3834);
and U4164 (N_4164,N_3499,N_2033);
or U4165 (N_4165,N_3510,N_2072);
or U4166 (N_4166,N_2518,N_3007);
and U4167 (N_4167,N_3105,N_2648);
xnor U4168 (N_4168,N_3291,N_2794);
xor U4169 (N_4169,N_2259,N_3344);
and U4170 (N_4170,N_3246,N_2863);
xnor U4171 (N_4171,N_2055,N_2205);
and U4172 (N_4172,N_3743,N_3343);
nor U4173 (N_4173,N_2267,N_2808);
and U4174 (N_4174,N_2186,N_3046);
nand U4175 (N_4175,N_3859,N_2919);
and U4176 (N_4176,N_2420,N_2215);
nor U4177 (N_4177,N_2163,N_2334);
nand U4178 (N_4178,N_2623,N_3492);
and U4179 (N_4179,N_2660,N_3139);
and U4180 (N_4180,N_3407,N_3701);
or U4181 (N_4181,N_2614,N_2206);
nand U4182 (N_4182,N_2481,N_3634);
nor U4183 (N_4183,N_3984,N_2524);
or U4184 (N_4184,N_2922,N_2673);
and U4185 (N_4185,N_3560,N_2636);
and U4186 (N_4186,N_2508,N_2938);
xor U4187 (N_4187,N_3532,N_2900);
xnor U4188 (N_4188,N_3636,N_2935);
or U4189 (N_4189,N_2820,N_2628);
nor U4190 (N_4190,N_2587,N_2506);
and U4191 (N_4191,N_2682,N_3297);
and U4192 (N_4192,N_3959,N_3088);
or U4193 (N_4193,N_2397,N_2108);
and U4194 (N_4194,N_3261,N_2412);
nor U4195 (N_4195,N_3693,N_3275);
xor U4196 (N_4196,N_3848,N_3880);
and U4197 (N_4197,N_3034,N_3949);
nand U4198 (N_4198,N_2915,N_2468);
or U4199 (N_4199,N_2473,N_3748);
xnor U4200 (N_4200,N_3577,N_2358);
and U4201 (N_4201,N_2702,N_2283);
nor U4202 (N_4202,N_3129,N_2044);
or U4203 (N_4203,N_3822,N_3038);
nand U4204 (N_4204,N_2441,N_3586);
or U4205 (N_4205,N_2746,N_3084);
and U4206 (N_4206,N_2867,N_3534);
xor U4207 (N_4207,N_2632,N_2118);
xor U4208 (N_4208,N_3483,N_2012);
nand U4209 (N_4209,N_3905,N_3273);
and U4210 (N_4210,N_2644,N_2464);
or U4211 (N_4211,N_3758,N_2485);
xnor U4212 (N_4212,N_2391,N_3418);
xor U4213 (N_4213,N_3374,N_3832);
xnor U4214 (N_4214,N_2337,N_3337);
and U4215 (N_4215,N_2386,N_2169);
or U4216 (N_4216,N_2226,N_3321);
and U4217 (N_4217,N_3290,N_3223);
xor U4218 (N_4218,N_3940,N_3387);
xor U4219 (N_4219,N_2568,N_2328);
nand U4220 (N_4220,N_2074,N_2372);
and U4221 (N_4221,N_2939,N_2523);
nand U4222 (N_4222,N_2045,N_3244);
nor U4223 (N_4223,N_2753,N_2515);
nand U4224 (N_4224,N_3167,N_3778);
and U4225 (N_4225,N_2189,N_3573);
and U4226 (N_4226,N_3765,N_3567);
xor U4227 (N_4227,N_2723,N_3779);
or U4228 (N_4228,N_2132,N_3180);
or U4229 (N_4229,N_3947,N_2652);
and U4230 (N_4230,N_2849,N_3060);
xnor U4231 (N_4231,N_3909,N_2992);
nand U4232 (N_4232,N_2277,N_2600);
and U4233 (N_4233,N_3893,N_2604);
or U4234 (N_4234,N_3762,N_3564);
nand U4235 (N_4235,N_3141,N_2551);
and U4236 (N_4236,N_2990,N_3995);
or U4237 (N_4237,N_2300,N_2291);
nand U4238 (N_4238,N_2264,N_2347);
and U4239 (N_4239,N_3921,N_2478);
and U4240 (N_4240,N_3868,N_2252);
nor U4241 (N_4241,N_3799,N_2285);
nor U4242 (N_4242,N_2817,N_3807);
nand U4243 (N_4243,N_3663,N_2278);
xnor U4244 (N_4244,N_3808,N_3718);
or U4245 (N_4245,N_3698,N_3205);
or U4246 (N_4246,N_3185,N_2492);
nor U4247 (N_4247,N_2445,N_2127);
and U4248 (N_4248,N_2949,N_2635);
and U4249 (N_4249,N_2575,N_3368);
or U4250 (N_4250,N_3138,N_3682);
and U4251 (N_4251,N_3477,N_3692);
xor U4252 (N_4252,N_2216,N_2601);
xor U4253 (N_4253,N_2006,N_3656);
and U4254 (N_4254,N_2349,N_3608);
and U4255 (N_4255,N_3154,N_2116);
and U4256 (N_4256,N_2089,N_3442);
xor U4257 (N_4257,N_2177,N_3796);
and U4258 (N_4258,N_2173,N_3414);
nand U4259 (N_4259,N_2041,N_2703);
xnor U4260 (N_4260,N_2677,N_2643);
xor U4261 (N_4261,N_2708,N_2844);
or U4262 (N_4262,N_3015,N_2256);
xor U4263 (N_4263,N_2435,N_2477);
nor U4264 (N_4264,N_2140,N_2995);
or U4265 (N_4265,N_2582,N_2174);
and U4266 (N_4266,N_2367,N_2212);
and U4267 (N_4267,N_2279,N_2310);
xor U4268 (N_4268,N_2380,N_2338);
and U4269 (N_4269,N_3437,N_2415);
or U4270 (N_4270,N_3411,N_2408);
xnor U4271 (N_4271,N_2562,N_3827);
and U4272 (N_4272,N_3003,N_3896);
xor U4273 (N_4273,N_3177,N_2043);
or U4274 (N_4274,N_2847,N_2350);
or U4275 (N_4275,N_3578,N_3842);
or U4276 (N_4276,N_2172,N_2411);
or U4277 (N_4277,N_3476,N_3454);
nor U4278 (N_4278,N_2697,N_2018);
nand U4279 (N_4279,N_3509,N_3996);
nor U4280 (N_4280,N_3254,N_3466);
xnor U4281 (N_4281,N_2810,N_2036);
or U4282 (N_4282,N_3899,N_3723);
nor U4283 (N_4283,N_3019,N_3795);
nor U4284 (N_4284,N_3487,N_3262);
and U4285 (N_4285,N_2668,N_3190);
or U4286 (N_4286,N_3065,N_3686);
nor U4287 (N_4287,N_3985,N_2565);
or U4288 (N_4288,N_2001,N_3033);
or U4289 (N_4289,N_3794,N_2522);
nor U4290 (N_4290,N_2268,N_2241);
or U4291 (N_4291,N_2292,N_3420);
and U4292 (N_4292,N_3916,N_3626);
and U4293 (N_4293,N_2705,N_2961);
nor U4294 (N_4294,N_3887,N_2145);
xnor U4295 (N_4295,N_3742,N_2092);
xnor U4296 (N_4296,N_3313,N_3963);
nand U4297 (N_4297,N_2305,N_3517);
nor U4298 (N_4298,N_3753,N_2222);
xor U4299 (N_4299,N_2903,N_2857);
nor U4300 (N_4300,N_3080,N_2377);
nand U4301 (N_4301,N_2813,N_3100);
xor U4302 (N_4302,N_3111,N_3638);
nand U4303 (N_4303,N_3128,N_3941);
or U4304 (N_4304,N_3551,N_3432);
nand U4305 (N_4305,N_3075,N_3645);
or U4306 (N_4306,N_2021,N_2774);
nand U4307 (N_4307,N_3159,N_3927);
xor U4308 (N_4308,N_2250,N_2204);
xnor U4309 (N_4309,N_3937,N_3237);
nand U4310 (N_4310,N_2282,N_2627);
xnor U4311 (N_4311,N_3540,N_2918);
nand U4312 (N_4312,N_2262,N_2090);
and U4313 (N_4313,N_2426,N_2249);
xor U4314 (N_4314,N_3604,N_2665);
xor U4315 (N_4315,N_2833,N_2002);
and U4316 (N_4316,N_3773,N_2942);
nor U4317 (N_4317,N_3417,N_2571);
or U4318 (N_4318,N_2710,N_3099);
xor U4319 (N_4319,N_2670,N_2861);
and U4320 (N_4320,N_3631,N_2288);
and U4321 (N_4321,N_3486,N_3703);
nor U4322 (N_4322,N_2086,N_3595);
and U4323 (N_4323,N_3439,N_2183);
or U4324 (N_4324,N_3484,N_3094);
nand U4325 (N_4325,N_2910,N_2850);
nor U4326 (N_4326,N_2371,N_2580);
xor U4327 (N_4327,N_2343,N_2168);
nor U4328 (N_4328,N_2780,N_2680);
nand U4329 (N_4329,N_3083,N_3654);
and U4330 (N_4330,N_2303,N_3469);
nor U4331 (N_4331,N_3358,N_3831);
or U4332 (N_4332,N_3964,N_3542);
and U4333 (N_4333,N_3786,N_2690);
nand U4334 (N_4334,N_3086,N_2311);
and U4335 (N_4335,N_3955,N_2052);
nor U4336 (N_4336,N_3973,N_2583);
nand U4337 (N_4337,N_2886,N_2359);
nand U4338 (N_4338,N_2130,N_2280);
nand U4339 (N_4339,N_2176,N_3464);
nor U4340 (N_4340,N_2869,N_2319);
and U4341 (N_4341,N_2706,N_3271);
or U4342 (N_4342,N_3118,N_3098);
nor U4343 (N_4343,N_2760,N_3301);
xnor U4344 (N_4344,N_2618,N_3266);
nor U4345 (N_4345,N_2020,N_2803);
nand U4346 (N_4346,N_3948,N_2783);
and U4347 (N_4347,N_2892,N_2865);
xnor U4348 (N_4348,N_2048,N_3521);
nand U4349 (N_4349,N_2879,N_2691);
and U4350 (N_4350,N_2547,N_3629);
nand U4351 (N_4351,N_2795,N_3911);
xor U4352 (N_4352,N_3388,N_3383);
xnor U4353 (N_4353,N_2889,N_3881);
nor U4354 (N_4354,N_3448,N_3699);
and U4355 (N_4355,N_3130,N_2778);
nand U4356 (N_4356,N_3336,N_3625);
and U4357 (N_4357,N_3198,N_3093);
xnor U4358 (N_4358,N_3897,N_3010);
or U4359 (N_4359,N_3357,N_3950);
nor U4360 (N_4360,N_3930,N_2789);
or U4361 (N_4361,N_3389,N_3012);
xnor U4362 (N_4362,N_3081,N_3274);
nand U4363 (N_4363,N_3352,N_3122);
or U4364 (N_4364,N_3170,N_3866);
nand U4365 (N_4365,N_3667,N_3761);
xnor U4366 (N_4366,N_3528,N_3946);
xnor U4367 (N_4367,N_2738,N_2142);
nand U4368 (N_4368,N_3175,N_2487);
xnor U4369 (N_4369,N_2081,N_3306);
xor U4370 (N_4370,N_3408,N_2925);
and U4371 (N_4371,N_3101,N_3907);
and U4372 (N_4372,N_2271,N_3048);
nor U4373 (N_4373,N_3673,N_3052);
or U4374 (N_4374,N_3826,N_3039);
nand U4375 (N_4375,N_3446,N_2452);
nand U4376 (N_4376,N_3249,N_3757);
nand U4377 (N_4377,N_2067,N_2170);
xor U4378 (N_4378,N_3133,N_3657);
nor U4379 (N_4379,N_2236,N_2374);
nand U4380 (N_4380,N_2699,N_2812);
nor U4381 (N_4381,N_3431,N_2567);
nor U4382 (N_4382,N_3855,N_2870);
xnor U4383 (N_4383,N_2597,N_3163);
nand U4384 (N_4384,N_2926,N_3269);
nor U4385 (N_4385,N_2977,N_3501);
and U4386 (N_4386,N_3676,N_3650);
xnor U4387 (N_4387,N_3740,N_3558);
or U4388 (N_4388,N_3495,N_2413);
nor U4389 (N_4389,N_2491,N_3640);
nand U4390 (N_4390,N_3876,N_2743);
xor U4391 (N_4391,N_2003,N_3302);
nor U4392 (N_4392,N_3706,N_2154);
and U4393 (N_4393,N_3861,N_2274);
nor U4394 (N_4394,N_2554,N_2436);
and U4395 (N_4395,N_3828,N_3990);
and U4396 (N_4396,N_3875,N_2927);
nand U4397 (N_4397,N_3230,N_2355);
and U4398 (N_4398,N_2872,N_2029);
xnor U4399 (N_4399,N_3166,N_3283);
nor U4400 (N_4400,N_2566,N_2550);
nor U4401 (N_4401,N_2862,N_3219);
or U4402 (N_4402,N_3314,N_2537);
and U4403 (N_4403,N_2704,N_3914);
nor U4404 (N_4404,N_2975,N_3471);
nor U4405 (N_4405,N_3434,N_2933);
nand U4406 (N_4406,N_2807,N_3421);
and U4407 (N_4407,N_3376,N_2257);
or U4408 (N_4408,N_2902,N_3363);
and U4409 (N_4409,N_2968,N_3598);
nand U4410 (N_4410,N_2299,N_3983);
nand U4411 (N_4411,N_2751,N_2894);
nor U4412 (N_4412,N_2885,N_2707);
and U4413 (N_4413,N_3788,N_3406);
and U4414 (N_4414,N_2401,N_2585);
nand U4415 (N_4415,N_3256,N_3473);
nand U4416 (N_4416,N_3049,N_3835);
nand U4417 (N_4417,N_2548,N_2141);
nand U4418 (N_4418,N_3892,N_3220);
nor U4419 (N_4419,N_2017,N_2231);
and U4420 (N_4420,N_2980,N_3689);
nand U4421 (N_4421,N_3999,N_3369);
or U4422 (N_4422,N_2765,N_3194);
and U4423 (N_4423,N_3202,N_3860);
or U4424 (N_4424,N_2687,N_2416);
xnor U4425 (N_4425,N_3457,N_3559);
xnor U4426 (N_4426,N_3366,N_2672);
and U4427 (N_4427,N_2223,N_3707);
and U4428 (N_4428,N_2224,N_2907);
nor U4429 (N_4429,N_3335,N_2275);
nor U4430 (N_4430,N_2156,N_2024);
and U4431 (N_4431,N_2138,N_2790);
nand U4432 (N_4432,N_3952,N_2720);
xor U4433 (N_4433,N_2899,N_3465);
nand U4434 (N_4434,N_2318,N_3489);
and U4435 (N_4435,N_3653,N_3055);
or U4436 (N_4436,N_2896,N_2983);
xor U4437 (N_4437,N_3258,N_3214);
nand U4438 (N_4438,N_3137,N_3115);
nor U4439 (N_4439,N_3865,N_2716);
or U4440 (N_4440,N_2769,N_2512);
xnor U4441 (N_4441,N_3063,N_2860);
nor U4442 (N_4442,N_2891,N_2748);
and U4443 (N_4443,N_2908,N_3282);
or U4444 (N_4444,N_3798,N_2510);
xnor U4445 (N_4445,N_2577,N_3066);
nand U4446 (N_4446,N_3801,N_2645);
xor U4447 (N_4447,N_2260,N_2724);
nor U4448 (N_4448,N_2749,N_2152);
or U4449 (N_4449,N_2428,N_3209);
nor U4450 (N_4450,N_2754,N_2479);
nand U4451 (N_4451,N_3975,N_2240);
xor U4452 (N_4452,N_3324,N_2210);
or U4453 (N_4453,N_3588,N_3613);
and U4454 (N_4454,N_2624,N_3463);
or U4455 (N_4455,N_2093,N_2050);
nand U4456 (N_4456,N_2117,N_3384);
and U4457 (N_4457,N_3206,N_3179);
nand U4458 (N_4458,N_2454,N_2077);
nand U4459 (N_4459,N_2731,N_3158);
nand U4460 (N_4460,N_3345,N_2663);
nor U4461 (N_4461,N_3380,N_3193);
nand U4462 (N_4462,N_2920,N_2028);
nor U4463 (N_4463,N_2931,N_3413);
nand U4464 (N_4464,N_3221,N_2315);
nand U4465 (N_4465,N_3210,N_3878);
nand U4466 (N_4466,N_3460,N_3609);
or U4467 (N_4467,N_2784,N_3441);
nand U4468 (N_4468,N_3775,N_2175);
nor U4469 (N_4469,N_3161,N_3327);
nor U4470 (N_4470,N_3928,N_2973);
nor U4471 (N_4471,N_3023,N_2549);
or U4472 (N_4472,N_3545,N_2096);
nand U4473 (N_4473,N_3268,N_3570);
or U4474 (N_4474,N_2657,N_3089);
nand U4475 (N_4475,N_3134,N_2946);
or U4476 (N_4476,N_3561,N_2819);
and U4477 (N_4477,N_2301,N_2666);
xor U4478 (N_4478,N_2417,N_3767);
and U4479 (N_4479,N_2185,N_3393);
or U4480 (N_4480,N_2895,N_2955);
nand U4481 (N_4481,N_2010,N_3427);
nor U4482 (N_4482,N_2365,N_3251);
or U4483 (N_4483,N_3072,N_2497);
or U4484 (N_4484,N_2556,N_2773);
and U4485 (N_4485,N_3201,N_2320);
or U4486 (N_4486,N_2461,N_3506);
nand U4487 (N_4487,N_2519,N_3110);
nor U4488 (N_4488,N_2119,N_2388);
and U4489 (N_4489,N_2928,N_3279);
and U4490 (N_4490,N_2978,N_2237);
and U4491 (N_4491,N_2061,N_3183);
nand U4492 (N_4492,N_2974,N_3869);
xnor U4493 (N_4493,N_2770,N_3354);
nor U4494 (N_4494,N_2828,N_3462);
nand U4495 (N_4495,N_2617,N_3236);
xor U4496 (N_4496,N_3864,N_2736);
nor U4497 (N_4497,N_2569,N_2725);
nand U4498 (N_4498,N_3392,N_3811);
nand U4499 (N_4499,N_2084,N_2923);
xnor U4500 (N_4500,N_2102,N_2664);
or U4501 (N_4501,N_2818,N_3708);
or U4502 (N_4502,N_3212,N_3529);
or U4503 (N_4503,N_2410,N_3030);
nand U4504 (N_4504,N_2433,N_2192);
or U4505 (N_4505,N_2444,N_2558);
or U4506 (N_4506,N_2768,N_2188);
or U4507 (N_4507,N_2385,N_3348);
or U4508 (N_4508,N_2429,N_3096);
xnor U4509 (N_4509,N_2711,N_2313);
nand U4510 (N_4510,N_3833,N_3005);
xnor U4511 (N_4511,N_3993,N_2112);
or U4512 (N_4512,N_3847,N_3837);
nor U4513 (N_4513,N_2348,N_2153);
xor U4514 (N_4514,N_3668,N_3342);
xor U4515 (N_4515,N_3160,N_2166);
xor U4516 (N_4516,N_3064,N_3809);
or U4517 (N_4517,N_3541,N_3058);
nor U4518 (N_4518,N_3951,N_2115);
and U4519 (N_4519,N_3872,N_2502);
nor U4520 (N_4520,N_3176,N_3511);
and U4521 (N_4521,N_2662,N_3156);
xnor U4522 (N_4522,N_2917,N_2781);
xor U4523 (N_4523,N_3543,N_3768);
or U4524 (N_4524,N_2952,N_3601);
or U4525 (N_4525,N_2679,N_2255);
and U4526 (N_4526,N_3697,N_3132);
xor U4527 (N_4527,N_2467,N_2196);
nand U4528 (N_4528,N_3323,N_3341);
xor U4529 (N_4529,N_2134,N_3224);
nand U4530 (N_4530,N_3945,N_2182);
or U4531 (N_4531,N_3364,N_2009);
nor U4532 (N_4532,N_2384,N_3904);
nand U4533 (N_4533,N_2996,N_2866);
xor U4534 (N_4534,N_2151,N_3405);
or U4535 (N_4535,N_2085,N_3565);
or U4536 (N_4536,N_3423,N_3671);
and U4537 (N_4537,N_2382,N_2039);
xor U4538 (N_4538,N_2150,N_2037);
or U4539 (N_4539,N_3710,N_3310);
or U4540 (N_4540,N_2135,N_3000);
xor U4541 (N_4541,N_2094,N_3186);
nand U4542 (N_4542,N_3610,N_3076);
and U4543 (N_4543,N_3804,N_2286);
and U4544 (N_4544,N_2409,N_3315);
or U4545 (N_4545,N_3997,N_2396);
xor U4546 (N_4546,N_3583,N_2611);
xnor U4547 (N_4547,N_3264,N_2659);
or U4548 (N_4548,N_2465,N_3329);
xor U4549 (N_4549,N_2976,N_2971);
nor U4550 (N_4550,N_2219,N_2105);
and U4551 (N_4551,N_2489,N_3018);
xnor U4552 (N_4552,N_2864,N_2739);
or U4553 (N_4553,N_2312,N_2825);
or U4554 (N_4554,N_3346,N_3789);
or U4555 (N_4555,N_3108,N_2998);
nand U4556 (N_4556,N_2031,N_3884);
nand U4557 (N_4557,N_2414,N_2871);
nand U4558 (N_4558,N_3173,N_2437);
and U4559 (N_4559,N_2772,N_3422);
xnor U4560 (N_4560,N_3724,N_2160);
or U4561 (N_4561,N_2242,N_2308);
or U4562 (N_4562,N_3774,N_3841);
nor U4563 (N_4563,N_2941,N_2476);
and U4564 (N_4564,N_2004,N_3073);
and U4565 (N_4565,N_2107,N_2104);
nor U4566 (N_4566,N_3147,N_2543);
and U4567 (N_4567,N_2555,N_3929);
and U4568 (N_4568,N_3378,N_2674);
xor U4569 (N_4569,N_3355,N_2984);
nor U4570 (N_4570,N_2579,N_3785);
nor U4571 (N_4571,N_3028,N_2793);
nand U4572 (N_4572,N_3593,N_3215);
xor U4573 (N_4573,N_2620,N_2621);
and U4574 (N_4574,N_3255,N_3450);
xnor U4575 (N_4575,N_3011,N_2394);
and U4576 (N_4576,N_2425,N_3621);
nor U4577 (N_4577,N_2207,N_3569);
xnor U4578 (N_4578,N_3923,N_2321);
or U4579 (N_4579,N_3591,N_2370);
xor U4580 (N_4580,N_2752,N_3218);
and U4581 (N_4581,N_2712,N_2187);
nor U4582 (N_4582,N_2809,N_3933);
or U4583 (N_4583,N_2669,N_3480);
xor U4584 (N_4584,N_2162,N_2909);
or U4585 (N_4585,N_2405,N_2527);
nand U4586 (N_4586,N_3777,N_2329);
nand U4587 (N_4587,N_3690,N_2235);
nand U4588 (N_4588,N_2905,N_2501);
nor U4589 (N_4589,N_2612,N_2822);
or U4590 (N_4590,N_2901,N_3228);
nand U4591 (N_4591,N_3216,N_2336);
nand U4592 (N_4592,N_2779,N_2880);
and U4593 (N_4593,N_3524,N_3356);
or U4594 (N_4594,N_2184,N_2693);
nor U4595 (N_4595,N_3047,N_3447);
and U4596 (N_4596,N_2619,N_3957);
or U4597 (N_4597,N_3770,N_2211);
xor U4598 (N_4598,N_2378,N_2421);
or U4599 (N_4599,N_3582,N_2221);
or U4600 (N_4600,N_2873,N_2685);
or U4601 (N_4601,N_2466,N_2379);
or U4602 (N_4602,N_2361,N_3208);
and U4603 (N_4603,N_3920,N_3222);
nor U4604 (N_4604,N_2937,N_3278);
nor U4605 (N_4605,N_2040,N_2741);
or U4606 (N_4606,N_3987,N_3688);
xnor U4607 (N_4607,N_2419,N_2525);
and U4608 (N_4608,N_3106,N_3362);
nand U4609 (N_4609,N_2529,N_3883);
nand U4610 (N_4610,N_2858,N_2758);
xor U4611 (N_4611,N_2500,N_2851);
xor U4612 (N_4612,N_3425,N_2837);
nor U4613 (N_4613,N_2985,N_2830);
or U4614 (N_4614,N_2383,N_2689);
nand U4615 (N_4615,N_2199,N_3087);
xor U4616 (N_4616,N_3550,N_3459);
nand U4617 (N_4617,N_3270,N_2930);
xor U4618 (N_4618,N_2395,N_3120);
nand U4619 (N_4619,N_2904,N_2179);
and U4620 (N_4620,N_2013,N_3396);
nand U4621 (N_4621,N_2788,N_3340);
nand U4622 (N_4622,N_3318,N_3059);
xor U4623 (N_4623,N_3286,N_3284);
nand U4624 (N_4624,N_3885,N_3157);
or U4625 (N_4625,N_2836,N_3433);
or U4626 (N_4626,N_3289,N_3037);
nand U4627 (N_4627,N_3013,N_2622);
xnor U4628 (N_4628,N_2254,N_3584);
xor U4629 (N_4629,N_3611,N_3428);
or U4630 (N_4630,N_2314,N_3844);
xor U4631 (N_4631,N_3526,N_3803);
xor U4632 (N_4632,N_3781,N_2771);
or U4633 (N_4633,N_2109,N_3412);
or U4634 (N_4634,N_3938,N_2997);
xor U4635 (N_4635,N_3296,N_3971);
nand U4636 (N_4636,N_2364,N_2046);
nand U4637 (N_4637,N_3674,N_3197);
or U4638 (N_4638,N_3409,N_2609);
nand U4639 (N_4639,N_2403,N_3600);
or U4640 (N_4640,N_2967,N_2446);
xor U4641 (N_4641,N_3647,N_3485);
nand U4642 (N_4642,N_2165,N_2530);
and U4643 (N_4643,N_2734,N_3061);
nor U4644 (N_4644,N_2431,N_2197);
or U4645 (N_4645,N_3260,N_2369);
and U4646 (N_4646,N_3615,N_2563);
or U4647 (N_4647,N_2958,N_2233);
nor U4648 (N_4648,N_2650,N_2641);
nand U4649 (N_4649,N_2531,N_3211);
and U4650 (N_4650,N_2125,N_2966);
and U4651 (N_4651,N_3664,N_2561);
and U4652 (N_4652,N_2700,N_2557);
xor U4653 (N_4653,N_3204,N_2533);
xnor U4654 (N_4654,N_2071,N_2198);
nand U4655 (N_4655,N_2167,N_3109);
or U4656 (N_4656,N_3776,N_2605);
or U4657 (N_4657,N_3862,N_2786);
and U4658 (N_4658,N_3679,N_2593);
nor U4659 (N_4659,N_3838,N_3716);
or U4660 (N_4660,N_3845,N_2217);
nor U4661 (N_4661,N_2307,N_3694);
and U4662 (N_4662,N_2353,N_2883);
xnor U4663 (N_4663,N_3068,N_2114);
nor U4664 (N_4664,N_3229,N_3587);
nor U4665 (N_4665,N_2243,N_3680);
or U4666 (N_4666,N_2027,N_3438);
nor U4667 (N_4667,N_2757,N_3497);
or U4668 (N_4668,N_3979,N_2509);
xor U4669 (N_4669,N_3257,N_3292);
or U4670 (N_4670,N_3051,N_3143);
nor U4671 (N_4671,N_2814,N_2058);
xor U4672 (N_4672,N_3720,N_2064);
and U4673 (N_4673,N_3994,N_3643);
nand U4674 (N_4674,N_2295,N_2326);
xor U4675 (N_4675,N_2000,N_2696);
nand U4676 (N_4676,N_2331,N_3006);
xor U4677 (N_4677,N_2573,N_2066);
xnor U4678 (N_4678,N_3764,N_3649);
and U4679 (N_4679,N_3238,N_2332);
nand U4680 (N_4680,N_3754,N_2270);
and U4681 (N_4681,N_3044,N_3735);
and U4682 (N_4682,N_2034,N_3953);
xor U4683 (N_4683,N_3630,N_3908);
or U4684 (N_4684,N_3882,N_3901);
nor U4685 (N_4685,N_3982,N_3311);
nand U4686 (N_4686,N_2874,N_2737);
or U4687 (N_4687,N_3749,N_2253);
xnor U4688 (N_4688,N_3918,N_2422);
xor U4689 (N_4689,N_2881,N_3053);
xnor U4690 (N_4690,N_2914,N_2069);
or U4691 (N_4691,N_2060,N_3700);
nand U4692 (N_4692,N_2471,N_3241);
xor U4693 (N_4693,N_2876,N_3576);
nor U4694 (N_4694,N_3456,N_2335);
and U4695 (N_4695,N_2532,N_3988);
and U4696 (N_4696,N_3902,N_2227);
nand U4697 (N_4697,N_3853,N_2595);
and U4698 (N_4698,N_3713,N_2802);
nor U4699 (N_4699,N_3498,N_2448);
nand U4700 (N_4700,N_3142,N_3523);
or U4701 (N_4701,N_2960,N_3575);
and U4702 (N_4702,N_2826,N_3572);
or U4703 (N_4703,N_3816,N_2606);
nand U4704 (N_4704,N_3633,N_3140);
and U4705 (N_4705,N_2766,N_2887);
xnor U4706 (N_4706,N_2916,N_2785);
or U4707 (N_4707,N_2079,N_3415);
and U4708 (N_4708,N_3747,N_2787);
or U4709 (N_4709,N_3351,N_3300);
xor U4710 (N_4710,N_3225,N_3001);
and U4711 (N_4711,N_3042,N_3568);
and U4712 (N_4712,N_2103,N_2956);
nand U4713 (N_4713,N_3589,N_2655);
nor U4714 (N_4714,N_2022,N_3886);
xnor U4715 (N_4715,N_3863,N_3915);
or U4716 (N_4716,N_3755,N_2854);
nand U4717 (N_4717,N_2298,N_3579);
xnor U4718 (N_4718,N_2811,N_2316);
or U4719 (N_4719,N_3605,N_2596);
nor U4720 (N_4720,N_3870,N_2991);
nand U4721 (N_4721,N_3054,N_2398);
xnor U4722 (N_4722,N_2782,N_2456);
nor U4723 (N_4723,N_2846,N_2947);
nor U4724 (N_4724,N_2526,N_2276);
nand U4725 (N_4725,N_3935,N_3085);
nand U4726 (N_4726,N_3242,N_3029);
nor U4727 (N_4727,N_3184,N_3616);
nor U4728 (N_4728,N_3596,N_2180);
or U4729 (N_4729,N_3475,N_2796);
nand U4730 (N_4730,N_3107,N_2193);
nand U4731 (N_4731,N_3424,N_3304);
nand U4732 (N_4732,N_2229,N_3515);
nand U4733 (N_4733,N_2954,N_2008);
or U4734 (N_4734,N_2341,N_2244);
xor U4735 (N_4735,N_2356,N_3151);
nand U4736 (N_4736,N_2763,N_3103);
or U4737 (N_4737,N_2791,N_3873);
and U4738 (N_4738,N_3627,N_3153);
nand U4739 (N_4739,N_3732,N_3240);
xor U4740 (N_4740,N_2159,N_2327);
or U4741 (N_4741,N_2201,N_3817);
or U4742 (N_4742,N_2306,N_3127);
nand U4743 (N_4743,N_3972,N_3954);
nor U4744 (N_4744,N_3646,N_2121);
and U4745 (N_4745,N_3470,N_3168);
nor U4746 (N_4746,N_3691,N_3962);
nor U4747 (N_4747,N_3285,N_3594);
or U4748 (N_4748,N_2023,N_3533);
nand U4749 (N_4749,N_3500,N_2934);
nand U4750 (N_4750,N_2982,N_2559);
or U4751 (N_4751,N_2137,N_3430);
nand U4752 (N_4752,N_2126,N_3537);
nand U4753 (N_4753,N_2921,N_3741);
xor U4754 (N_4754,N_3925,N_2111);
and U4755 (N_4755,N_2957,N_2038);
nand U4756 (N_4756,N_3677,N_3662);
nor U4757 (N_4757,N_3675,N_3243);
nor U4758 (N_4758,N_2496,N_3199);
and U4759 (N_4759,N_3518,N_2944);
and U4760 (N_4760,N_3823,N_3717);
nand U4761 (N_4761,N_2613,N_3856);
nand U4762 (N_4762,N_2661,N_3203);
nor U4763 (N_4763,N_2442,N_2342);
nand U4764 (N_4764,N_2075,N_3730);
nor U4765 (N_4765,N_3555,N_3821);
nand U4766 (N_4766,N_3097,N_2994);
or U4767 (N_4767,N_3267,N_3217);
nand U4768 (N_4768,N_3478,N_3095);
and U4769 (N_4769,N_3850,N_3045);
or U4770 (N_4770,N_2829,N_3125);
nor U4771 (N_4771,N_3239,N_3312);
xor U4772 (N_4772,N_3922,N_2853);
and U4773 (N_4773,N_2545,N_3375);
xor U4774 (N_4774,N_2570,N_3410);
nand U4775 (N_4775,N_3377,N_3619);
nor U4776 (N_4776,N_2979,N_2258);
xnor U4777 (N_4777,N_2407,N_3553);
nor U4778 (N_4778,N_2051,N_3114);
nor U4779 (N_4779,N_3395,N_2144);
or U4780 (N_4780,N_3234,N_3966);
xnor U4781 (N_4781,N_2729,N_2450);
or U4782 (N_4782,N_2709,N_3091);
nand U4783 (N_4783,N_3714,N_3531);
xnor U4784 (N_4784,N_3820,N_2030);
nor U4785 (N_4785,N_3520,N_2929);
nor U4786 (N_4786,N_3331,N_2855);
or U4787 (N_4787,N_3612,N_3563);
and U4788 (N_4788,N_3894,N_2578);
nor U4789 (N_4789,N_3232,N_3998);
xor U4790 (N_4790,N_3035,N_3678);
nand U4791 (N_4791,N_3642,N_3112);
nand U4792 (N_4792,N_3751,N_3334);
and U4793 (N_4793,N_2875,N_2840);
xnor U4794 (N_4794,N_2139,N_2572);
and U4795 (N_4795,N_3404,N_2483);
and U4796 (N_4796,N_3328,N_3032);
nand U4797 (N_4797,N_3958,N_3655);
xor U4798 (N_4798,N_3641,N_2649);
nand U4799 (N_4799,N_2011,N_2054);
xor U4800 (N_4800,N_3288,N_3020);
and U4801 (N_4801,N_3333,N_2728);
or U4802 (N_4802,N_3632,N_3092);
xnor U4803 (N_4803,N_2598,N_2494);
or U4804 (N_4804,N_3736,N_2835);
xnor U4805 (N_4805,N_3981,N_3874);
or U4806 (N_4806,N_3898,N_2097);
nand U4807 (N_4807,N_3169,N_3867);
xor U4808 (N_4808,N_3792,N_2434);
xor U4809 (N_4809,N_2745,N_3400);
nor U4810 (N_4810,N_3294,N_3852);
nor U4811 (N_4811,N_3056,N_3280);
xor U4812 (N_4812,N_2317,N_2375);
and U4813 (N_4813,N_3602,N_3146);
nand U4814 (N_4814,N_2912,N_3644);
nand U4815 (N_4815,N_3960,N_2143);
and U4816 (N_4816,N_3931,N_3507);
xnor U4817 (N_4817,N_3305,N_3750);
xnor U4818 (N_4818,N_3164,N_2482);
xor U4819 (N_4819,N_3547,N_3727);
xnor U4820 (N_4820,N_3021,N_2218);
nor U4821 (N_4821,N_3265,N_3123);
or U4822 (N_4822,N_3025,N_3207);
nor U4823 (N_4823,N_3967,N_2323);
nand U4824 (N_4824,N_2220,N_3359);
nor U4825 (N_4825,N_3317,N_2095);
nor U4826 (N_4826,N_3760,N_2015);
nor U4827 (N_4827,N_2658,N_2459);
and U4828 (N_4828,N_2246,N_3665);
and U4829 (N_4829,N_2124,N_3116);
xnor U4830 (N_4830,N_3628,N_2430);
nor U4831 (N_4831,N_2451,N_2376);
and U4832 (N_4832,N_2815,N_3571);
and U4833 (N_4833,N_2068,N_3017);
nand U4834 (N_4834,N_3756,N_2683);
and U4835 (N_4835,N_3458,N_2698);
nand U4836 (N_4836,N_2590,N_3004);
or U4837 (N_4837,N_3815,N_3512);
and U4838 (N_4838,N_2560,N_3339);
or U4839 (N_4839,N_2475,N_3538);
nand U4840 (N_4840,N_2540,N_3398);
nand U4841 (N_4841,N_2248,N_2423);
or U4842 (N_4842,N_2056,N_2208);
nor U4843 (N_4843,N_2897,N_3505);
nand U4844 (N_4844,N_3939,N_3226);
nand U4845 (N_4845,N_2340,N_3162);
nor U4846 (N_4846,N_2588,N_3074);
and U4847 (N_4847,N_3956,N_3739);
xnor U4848 (N_4848,N_3298,N_2798);
xor U4849 (N_4849,N_3451,N_2284);
nand U4850 (N_4850,N_3308,N_3468);
nor U4851 (N_4851,N_3397,N_2354);
nand U4852 (N_4852,N_3658,N_2490);
nand U4853 (N_4853,N_2629,N_2245);
xor U4854 (N_4854,N_3493,N_3516);
and U4855 (N_4855,N_2877,N_2750);
xnor U4856 (N_4856,N_3253,N_3452);
or U4857 (N_4857,N_2474,N_2458);
or U4858 (N_4858,N_2542,N_2959);
xor U4859 (N_4859,N_3503,N_3917);
nor U4860 (N_4860,N_2230,N_2131);
or U4861 (N_4861,N_2681,N_3281);
nor U4862 (N_4862,N_3695,N_2603);
or U4863 (N_4863,N_3390,N_2842);
and U4864 (N_4864,N_3196,N_3361);
nor U4865 (N_4865,N_3508,N_3307);
and U4866 (N_4866,N_2432,N_2868);
nand U4867 (N_4867,N_3299,N_2202);
nor U4868 (N_4868,N_2740,N_3769);
xnor U4869 (N_4869,N_3711,N_3606);
xnor U4870 (N_4870,N_2638,N_3913);
or U4871 (N_4871,N_2171,N_2129);
and U4872 (N_4872,N_2806,N_3353);
nand U4873 (N_4873,N_3247,N_2913);
xor U4874 (N_4874,N_2507,N_2362);
and U4875 (N_4875,N_2265,N_3117);
and U4876 (N_4876,N_2238,N_2893);
nor U4877 (N_4877,N_3910,N_2035);
nand U4878 (N_4878,N_2161,N_2804);
xor U4879 (N_4879,N_3539,N_2839);
nand U4880 (N_4880,N_3527,N_3371);
nor U4881 (N_4881,N_3449,N_2747);
or U4882 (N_4882,N_2480,N_2503);
or U4883 (N_4883,N_2070,N_3912);
and U4884 (N_4884,N_3082,N_2100);
nand U4885 (N_4885,N_3401,N_3810);
nand U4886 (N_4886,N_2932,N_3581);
xor U4887 (N_4887,N_2726,N_2695);
nand U4888 (N_4888,N_3259,N_3737);
nor U4889 (N_4889,N_2521,N_3319);
or U4890 (N_4890,N_2488,N_2906);
nor U4891 (N_4891,N_2232,N_3729);
xor U4892 (N_4892,N_2363,N_2247);
nand U4893 (N_4893,N_3144,N_2106);
nand U4894 (N_4894,N_2744,N_2800);
xor U4895 (N_4895,N_3659,N_2164);
nor U4896 (N_4896,N_3504,N_2514);
and U4897 (N_4897,N_2504,N_3496);
and U4898 (N_4898,N_2293,N_2999);
nand U4899 (N_4899,N_2289,N_3752);
and U4900 (N_4900,N_2667,N_2538);
and U4901 (N_4901,N_3189,N_2963);
or U4902 (N_4902,N_3965,N_3090);
and U4903 (N_4903,N_2399,N_3126);
and U4904 (N_4904,N_3488,N_2742);
xor U4905 (N_4905,N_2653,N_2630);
or U4906 (N_4906,N_3702,N_2457);
xnor U4907 (N_4907,N_2181,N_3978);
nor U4908 (N_4908,N_3381,N_2146);
or U4909 (N_4909,N_3661,N_2732);
nand U4910 (N_4910,N_2586,N_2195);
and U4911 (N_4911,N_3078,N_2592);
or U4912 (N_4912,N_2200,N_3554);
or U4913 (N_4913,N_2823,N_2615);
nand U4914 (N_4914,N_3782,N_3840);
or U4915 (N_4915,N_3843,N_3712);
xor U4916 (N_4916,N_2962,N_3178);
or U4917 (N_4917,N_2147,N_3360);
nor U4918 (N_4918,N_2390,N_3970);
nand U4919 (N_4919,N_3113,N_3399);
nor U4920 (N_4920,N_2692,N_2511);
and U4921 (N_4921,N_2816,N_2007);
and U4922 (N_4922,N_2438,N_3696);
and U4923 (N_4923,N_2911,N_2493);
and U4924 (N_4924,N_3599,N_2404);
xnor U4925 (N_4925,N_3338,N_3548);
or U4926 (N_4926,N_2495,N_2684);
or U4927 (N_4927,N_2640,N_2714);
or U4928 (N_4928,N_3502,N_3614);
and U4929 (N_4929,N_3824,N_2733);
nor U4930 (N_4930,N_3681,N_3759);
nor U4931 (N_4931,N_3490,N_2964);
nor U4932 (N_4932,N_3349,N_3187);
nor U4933 (N_4933,N_2805,N_3802);
nand U4934 (N_4934,N_3192,N_2389);
xnor U4935 (N_4935,N_3191,N_3435);
and U4936 (N_4936,N_3043,N_3426);
nand U4937 (N_4937,N_3347,N_2099);
nor U4938 (N_4938,N_3027,N_3989);
nor U4939 (N_4939,N_2360,N_2505);
nand U4940 (N_4940,N_2178,N_2553);
nand U4941 (N_4941,N_3728,N_2209);
xnor U4942 (N_4942,N_2047,N_3402);
or U4943 (N_4943,N_2759,N_3819);
xor U4944 (N_4944,N_3556,N_2083);
nand U4945 (N_4945,N_2472,N_2637);
or U4946 (N_4946,N_3536,N_3121);
and U4947 (N_4947,N_3391,N_2133);
or U4948 (N_4948,N_3104,N_3002);
nand U4949 (N_4949,N_2821,N_3330);
and U4950 (N_4950,N_2345,N_3926);
and U4951 (N_4951,N_2534,N_2888);
or U4952 (N_4952,N_2190,N_2827);
and U4953 (N_4953,N_2676,N_2440);
nand U4954 (N_4954,N_2541,N_2059);
and U4955 (N_4955,N_3277,N_3379);
or U4956 (N_4956,N_3474,N_2406);
xnor U4957 (N_4957,N_2675,N_3793);
nor U4958 (N_4958,N_2439,N_2088);
or U4959 (N_4959,N_2076,N_2552);
and U4960 (N_4960,N_3620,N_3546);
and U4961 (N_4961,N_3248,N_3726);
xor U4962 (N_4962,N_2884,N_3784);
and U4963 (N_4963,N_2393,N_3174);
nor U4964 (N_4964,N_2455,N_2351);
nand U4965 (N_4965,N_2424,N_3227);
nor U4966 (N_4966,N_2607,N_3287);
and U4967 (N_4967,N_3026,N_3687);
and U4968 (N_4968,N_3974,N_3618);
and U4969 (N_4969,N_3854,N_3050);
nand U4970 (N_4970,N_2357,N_3245);
and U4971 (N_4971,N_2486,N_2718);
nand U4972 (N_4972,N_3235,N_2843);
and U4973 (N_4973,N_3102,N_2073);
xor U4974 (N_4974,N_2761,N_3891);
nand U4975 (N_4975,N_2101,N_2735);
xnor U4976 (N_4976,N_2381,N_3900);
or U4977 (N_4977,N_2924,N_2943);
or U4978 (N_4978,N_2373,N_3977);
nand U4979 (N_4979,N_2589,N_3797);
xor U4980 (N_4980,N_3367,N_2469);
or U4981 (N_4981,N_3976,N_3666);
nand U4982 (N_4982,N_3818,N_3181);
xnor U4983 (N_4983,N_3791,N_3320);
xor U4984 (N_4984,N_2688,N_2065);
or U4985 (N_4985,N_3574,N_3590);
xnor U4986 (N_4986,N_2368,N_3648);
or U4987 (N_4987,N_2646,N_3877);
or U4988 (N_4988,N_3813,N_2019);
or U4989 (N_4989,N_3386,N_2651);
and U4990 (N_4990,N_2762,N_3440);
xnor U4991 (N_4991,N_3932,N_2799);
xor U4992 (N_4992,N_2767,N_2878);
xnor U4993 (N_4993,N_2951,N_2324);
nand U4994 (N_4994,N_3008,N_3660);
nor U4995 (N_4995,N_3482,N_3734);
or U4996 (N_4996,N_3766,N_2948);
nor U4997 (N_4997,N_2263,N_2993);
nand U4998 (N_4998,N_3814,N_2719);
or U4999 (N_4999,N_2516,N_3200);
nor U5000 (N_5000,N_3758,N_2606);
or U5001 (N_5001,N_3466,N_2391);
and U5002 (N_5002,N_2021,N_2457);
nor U5003 (N_5003,N_3557,N_2228);
nand U5004 (N_5004,N_3668,N_3631);
or U5005 (N_5005,N_3775,N_3853);
or U5006 (N_5006,N_3777,N_2622);
nand U5007 (N_5007,N_2051,N_3591);
and U5008 (N_5008,N_2973,N_3279);
and U5009 (N_5009,N_3893,N_2901);
xor U5010 (N_5010,N_2953,N_2816);
nor U5011 (N_5011,N_2827,N_2063);
and U5012 (N_5012,N_3073,N_2289);
nand U5013 (N_5013,N_3814,N_3934);
nor U5014 (N_5014,N_3933,N_3665);
nor U5015 (N_5015,N_3909,N_2066);
or U5016 (N_5016,N_2164,N_2035);
or U5017 (N_5017,N_3678,N_2491);
nor U5018 (N_5018,N_3129,N_3885);
xnor U5019 (N_5019,N_3618,N_3186);
nand U5020 (N_5020,N_2754,N_3020);
nor U5021 (N_5021,N_2353,N_2229);
or U5022 (N_5022,N_2463,N_3855);
nand U5023 (N_5023,N_3235,N_2081);
or U5024 (N_5024,N_3229,N_3647);
nand U5025 (N_5025,N_3953,N_2485);
or U5026 (N_5026,N_2896,N_2066);
or U5027 (N_5027,N_3344,N_2350);
xnor U5028 (N_5028,N_3560,N_3716);
xor U5029 (N_5029,N_3084,N_2348);
nor U5030 (N_5030,N_2321,N_3857);
and U5031 (N_5031,N_3316,N_2373);
nor U5032 (N_5032,N_3203,N_3845);
or U5033 (N_5033,N_3907,N_2050);
or U5034 (N_5034,N_3628,N_3734);
nor U5035 (N_5035,N_3712,N_2777);
nand U5036 (N_5036,N_3668,N_3321);
xnor U5037 (N_5037,N_3262,N_2991);
and U5038 (N_5038,N_3981,N_3559);
or U5039 (N_5039,N_2010,N_2533);
nand U5040 (N_5040,N_2609,N_3795);
and U5041 (N_5041,N_3989,N_2534);
nand U5042 (N_5042,N_2510,N_2552);
or U5043 (N_5043,N_3185,N_2599);
xnor U5044 (N_5044,N_3933,N_2478);
nor U5045 (N_5045,N_3499,N_2583);
or U5046 (N_5046,N_3598,N_3949);
nand U5047 (N_5047,N_2223,N_3668);
nand U5048 (N_5048,N_3630,N_3091);
and U5049 (N_5049,N_2142,N_3484);
nor U5050 (N_5050,N_2873,N_3289);
nor U5051 (N_5051,N_3231,N_3040);
xor U5052 (N_5052,N_2216,N_2015);
or U5053 (N_5053,N_2582,N_3080);
nor U5054 (N_5054,N_3840,N_3272);
and U5055 (N_5055,N_2047,N_2162);
nor U5056 (N_5056,N_3407,N_3747);
xnor U5057 (N_5057,N_2021,N_3516);
nand U5058 (N_5058,N_3961,N_3414);
nor U5059 (N_5059,N_2225,N_3837);
and U5060 (N_5060,N_3716,N_3601);
and U5061 (N_5061,N_2761,N_3543);
xnor U5062 (N_5062,N_3317,N_2854);
nand U5063 (N_5063,N_3288,N_3080);
xor U5064 (N_5064,N_2052,N_2905);
and U5065 (N_5065,N_3936,N_2729);
or U5066 (N_5066,N_2688,N_3625);
and U5067 (N_5067,N_2801,N_2828);
nor U5068 (N_5068,N_2873,N_3741);
or U5069 (N_5069,N_2859,N_3636);
nand U5070 (N_5070,N_2946,N_2445);
and U5071 (N_5071,N_2141,N_3144);
nor U5072 (N_5072,N_2009,N_3760);
or U5073 (N_5073,N_3617,N_3136);
and U5074 (N_5074,N_3747,N_2918);
and U5075 (N_5075,N_2756,N_3101);
xor U5076 (N_5076,N_2564,N_2490);
or U5077 (N_5077,N_3782,N_2828);
and U5078 (N_5078,N_3439,N_3438);
nand U5079 (N_5079,N_2578,N_2254);
nand U5080 (N_5080,N_2371,N_2058);
and U5081 (N_5081,N_3083,N_2419);
or U5082 (N_5082,N_3731,N_3104);
nor U5083 (N_5083,N_3476,N_3059);
nor U5084 (N_5084,N_2705,N_3480);
xor U5085 (N_5085,N_3157,N_2163);
and U5086 (N_5086,N_2903,N_2017);
nand U5087 (N_5087,N_2712,N_3160);
nand U5088 (N_5088,N_2512,N_3707);
nand U5089 (N_5089,N_2500,N_2717);
and U5090 (N_5090,N_2392,N_2966);
xnor U5091 (N_5091,N_3360,N_3959);
nor U5092 (N_5092,N_2633,N_2677);
nor U5093 (N_5093,N_3006,N_3853);
and U5094 (N_5094,N_2242,N_3752);
and U5095 (N_5095,N_2556,N_2299);
and U5096 (N_5096,N_2453,N_2786);
xor U5097 (N_5097,N_2423,N_2059);
or U5098 (N_5098,N_2651,N_3625);
xnor U5099 (N_5099,N_2308,N_3900);
or U5100 (N_5100,N_3923,N_2811);
or U5101 (N_5101,N_2125,N_2732);
and U5102 (N_5102,N_2355,N_3527);
and U5103 (N_5103,N_2266,N_2997);
nand U5104 (N_5104,N_2202,N_3564);
nor U5105 (N_5105,N_2891,N_3042);
xor U5106 (N_5106,N_3632,N_3257);
nor U5107 (N_5107,N_2948,N_2230);
and U5108 (N_5108,N_3738,N_2028);
nor U5109 (N_5109,N_2256,N_3191);
or U5110 (N_5110,N_2894,N_2957);
and U5111 (N_5111,N_3005,N_3726);
and U5112 (N_5112,N_2124,N_3013);
nand U5113 (N_5113,N_3017,N_3603);
nand U5114 (N_5114,N_2789,N_3150);
nand U5115 (N_5115,N_2489,N_2517);
xnor U5116 (N_5116,N_3520,N_2343);
and U5117 (N_5117,N_2887,N_3424);
nor U5118 (N_5118,N_2132,N_2017);
nor U5119 (N_5119,N_3470,N_2340);
nor U5120 (N_5120,N_2306,N_2717);
nor U5121 (N_5121,N_2352,N_2776);
or U5122 (N_5122,N_3059,N_3248);
or U5123 (N_5123,N_3152,N_2093);
or U5124 (N_5124,N_3403,N_3896);
xnor U5125 (N_5125,N_2202,N_3938);
and U5126 (N_5126,N_3687,N_3067);
or U5127 (N_5127,N_2960,N_3316);
nand U5128 (N_5128,N_2413,N_3667);
nand U5129 (N_5129,N_3952,N_3155);
and U5130 (N_5130,N_2676,N_2818);
xnor U5131 (N_5131,N_2369,N_3231);
or U5132 (N_5132,N_3194,N_2381);
nand U5133 (N_5133,N_2210,N_3175);
or U5134 (N_5134,N_2582,N_2074);
xnor U5135 (N_5135,N_3414,N_3178);
nor U5136 (N_5136,N_3950,N_2581);
and U5137 (N_5137,N_2047,N_3242);
or U5138 (N_5138,N_3361,N_2242);
xnor U5139 (N_5139,N_3336,N_2161);
nand U5140 (N_5140,N_3393,N_2797);
and U5141 (N_5141,N_2134,N_2743);
xnor U5142 (N_5142,N_2317,N_3978);
nor U5143 (N_5143,N_3504,N_2920);
or U5144 (N_5144,N_2871,N_3766);
or U5145 (N_5145,N_3086,N_2133);
nand U5146 (N_5146,N_3125,N_2275);
nor U5147 (N_5147,N_3613,N_3069);
and U5148 (N_5148,N_3048,N_3929);
and U5149 (N_5149,N_3391,N_2006);
nand U5150 (N_5150,N_3824,N_3753);
xnor U5151 (N_5151,N_3470,N_2135);
nand U5152 (N_5152,N_2546,N_3272);
xor U5153 (N_5153,N_2165,N_3890);
or U5154 (N_5154,N_2713,N_2811);
or U5155 (N_5155,N_3572,N_2599);
and U5156 (N_5156,N_2058,N_2307);
nand U5157 (N_5157,N_2076,N_2116);
and U5158 (N_5158,N_2053,N_2909);
or U5159 (N_5159,N_2490,N_3369);
or U5160 (N_5160,N_2588,N_2010);
nand U5161 (N_5161,N_3555,N_2727);
and U5162 (N_5162,N_2953,N_3705);
nor U5163 (N_5163,N_3815,N_3043);
nor U5164 (N_5164,N_3607,N_3040);
or U5165 (N_5165,N_2855,N_2591);
or U5166 (N_5166,N_3142,N_2289);
or U5167 (N_5167,N_2236,N_3054);
nor U5168 (N_5168,N_2787,N_3943);
or U5169 (N_5169,N_2487,N_2512);
nor U5170 (N_5170,N_3592,N_2848);
nor U5171 (N_5171,N_2473,N_2893);
nor U5172 (N_5172,N_3930,N_3863);
nand U5173 (N_5173,N_3953,N_2191);
and U5174 (N_5174,N_2791,N_2361);
or U5175 (N_5175,N_2543,N_2526);
nand U5176 (N_5176,N_3600,N_3816);
nand U5177 (N_5177,N_3036,N_3436);
xnor U5178 (N_5178,N_2874,N_2879);
nand U5179 (N_5179,N_2032,N_2240);
or U5180 (N_5180,N_3213,N_2059);
nor U5181 (N_5181,N_3353,N_2085);
nor U5182 (N_5182,N_2109,N_2178);
nand U5183 (N_5183,N_2980,N_3045);
xor U5184 (N_5184,N_2096,N_3814);
or U5185 (N_5185,N_2071,N_2736);
or U5186 (N_5186,N_3970,N_2730);
or U5187 (N_5187,N_2388,N_2904);
or U5188 (N_5188,N_3864,N_3930);
or U5189 (N_5189,N_2679,N_3928);
nand U5190 (N_5190,N_2416,N_2974);
and U5191 (N_5191,N_2201,N_2920);
nor U5192 (N_5192,N_3203,N_3570);
nor U5193 (N_5193,N_3354,N_2341);
and U5194 (N_5194,N_3652,N_2867);
xnor U5195 (N_5195,N_3622,N_2004);
and U5196 (N_5196,N_2783,N_2329);
nor U5197 (N_5197,N_2042,N_2525);
nor U5198 (N_5198,N_2767,N_2631);
nor U5199 (N_5199,N_2973,N_2370);
nand U5200 (N_5200,N_2374,N_2508);
or U5201 (N_5201,N_3671,N_3870);
or U5202 (N_5202,N_3234,N_3433);
nand U5203 (N_5203,N_3199,N_3347);
or U5204 (N_5204,N_3332,N_3327);
nand U5205 (N_5205,N_3189,N_2084);
nand U5206 (N_5206,N_2978,N_3645);
xor U5207 (N_5207,N_3053,N_3247);
or U5208 (N_5208,N_2227,N_3681);
or U5209 (N_5209,N_3975,N_3473);
or U5210 (N_5210,N_3877,N_2869);
and U5211 (N_5211,N_2257,N_3786);
or U5212 (N_5212,N_2226,N_3186);
nand U5213 (N_5213,N_3517,N_2418);
xor U5214 (N_5214,N_2465,N_2040);
xnor U5215 (N_5215,N_2621,N_3851);
nand U5216 (N_5216,N_2753,N_2045);
and U5217 (N_5217,N_2658,N_3276);
nand U5218 (N_5218,N_3906,N_2646);
nor U5219 (N_5219,N_2335,N_2873);
and U5220 (N_5220,N_3373,N_2875);
xnor U5221 (N_5221,N_3189,N_3880);
nor U5222 (N_5222,N_3519,N_2517);
nand U5223 (N_5223,N_3131,N_2788);
and U5224 (N_5224,N_3152,N_3457);
and U5225 (N_5225,N_2947,N_2115);
nor U5226 (N_5226,N_2466,N_3429);
xor U5227 (N_5227,N_2100,N_2075);
nand U5228 (N_5228,N_2445,N_3473);
xor U5229 (N_5229,N_3266,N_3147);
nor U5230 (N_5230,N_2647,N_2747);
xnor U5231 (N_5231,N_2131,N_2368);
xor U5232 (N_5232,N_2718,N_2038);
nand U5233 (N_5233,N_2121,N_3523);
and U5234 (N_5234,N_2263,N_3319);
nor U5235 (N_5235,N_3527,N_3587);
nor U5236 (N_5236,N_3657,N_3084);
and U5237 (N_5237,N_3248,N_3135);
xnor U5238 (N_5238,N_2242,N_2831);
xnor U5239 (N_5239,N_2397,N_2083);
xnor U5240 (N_5240,N_3035,N_2997);
or U5241 (N_5241,N_2023,N_3153);
or U5242 (N_5242,N_3985,N_2522);
or U5243 (N_5243,N_2030,N_2305);
nor U5244 (N_5244,N_2172,N_2206);
or U5245 (N_5245,N_2101,N_2456);
nand U5246 (N_5246,N_3112,N_2360);
nor U5247 (N_5247,N_2572,N_3435);
nor U5248 (N_5248,N_2997,N_2779);
or U5249 (N_5249,N_2186,N_3688);
nand U5250 (N_5250,N_2825,N_3195);
nor U5251 (N_5251,N_2495,N_2750);
nor U5252 (N_5252,N_3196,N_2992);
xor U5253 (N_5253,N_2678,N_2830);
and U5254 (N_5254,N_3262,N_3805);
xor U5255 (N_5255,N_2358,N_3664);
and U5256 (N_5256,N_3784,N_2379);
or U5257 (N_5257,N_3564,N_2655);
and U5258 (N_5258,N_3579,N_2462);
xor U5259 (N_5259,N_2819,N_2271);
or U5260 (N_5260,N_2060,N_2732);
nand U5261 (N_5261,N_2112,N_3571);
nor U5262 (N_5262,N_2529,N_2535);
nand U5263 (N_5263,N_2576,N_2470);
xnor U5264 (N_5264,N_3520,N_3920);
nand U5265 (N_5265,N_3103,N_3845);
and U5266 (N_5266,N_2935,N_3872);
and U5267 (N_5267,N_2142,N_3525);
and U5268 (N_5268,N_2256,N_2692);
nor U5269 (N_5269,N_3561,N_3057);
and U5270 (N_5270,N_2875,N_3422);
nor U5271 (N_5271,N_2178,N_3628);
nand U5272 (N_5272,N_2580,N_2017);
nor U5273 (N_5273,N_3757,N_2120);
nand U5274 (N_5274,N_3638,N_2952);
nand U5275 (N_5275,N_2235,N_2221);
and U5276 (N_5276,N_3581,N_2432);
nor U5277 (N_5277,N_2824,N_3621);
and U5278 (N_5278,N_2058,N_3511);
and U5279 (N_5279,N_2499,N_2033);
xnor U5280 (N_5280,N_2627,N_2358);
nor U5281 (N_5281,N_2061,N_2383);
nor U5282 (N_5282,N_3671,N_3797);
and U5283 (N_5283,N_2262,N_3029);
nor U5284 (N_5284,N_3953,N_3141);
xnor U5285 (N_5285,N_3159,N_2989);
and U5286 (N_5286,N_3843,N_2442);
nand U5287 (N_5287,N_3411,N_3917);
nor U5288 (N_5288,N_3253,N_3498);
and U5289 (N_5289,N_3157,N_2891);
and U5290 (N_5290,N_2806,N_2909);
nor U5291 (N_5291,N_3448,N_3350);
and U5292 (N_5292,N_3415,N_3759);
or U5293 (N_5293,N_3570,N_2881);
and U5294 (N_5294,N_2628,N_3981);
or U5295 (N_5295,N_2081,N_3858);
nor U5296 (N_5296,N_3585,N_2729);
or U5297 (N_5297,N_2032,N_2918);
xor U5298 (N_5298,N_3231,N_3611);
or U5299 (N_5299,N_3342,N_3350);
and U5300 (N_5300,N_3680,N_2252);
nand U5301 (N_5301,N_2123,N_2245);
xnor U5302 (N_5302,N_2108,N_3100);
and U5303 (N_5303,N_2564,N_3818);
nor U5304 (N_5304,N_3418,N_3144);
nand U5305 (N_5305,N_3355,N_3857);
and U5306 (N_5306,N_2727,N_3816);
xnor U5307 (N_5307,N_3230,N_3597);
nand U5308 (N_5308,N_2826,N_3282);
nor U5309 (N_5309,N_3570,N_3787);
nor U5310 (N_5310,N_3674,N_2672);
xnor U5311 (N_5311,N_3892,N_2612);
xnor U5312 (N_5312,N_2719,N_2089);
nand U5313 (N_5313,N_2059,N_3197);
nor U5314 (N_5314,N_3377,N_3341);
or U5315 (N_5315,N_3405,N_2723);
nand U5316 (N_5316,N_3254,N_3016);
nor U5317 (N_5317,N_3004,N_2072);
and U5318 (N_5318,N_3258,N_2367);
xor U5319 (N_5319,N_2539,N_2686);
and U5320 (N_5320,N_2486,N_2152);
nor U5321 (N_5321,N_2958,N_3320);
nand U5322 (N_5322,N_3040,N_3610);
and U5323 (N_5323,N_2568,N_3257);
nor U5324 (N_5324,N_2069,N_2815);
nor U5325 (N_5325,N_2416,N_2318);
and U5326 (N_5326,N_2335,N_2543);
xnor U5327 (N_5327,N_3477,N_3761);
and U5328 (N_5328,N_3774,N_3344);
xnor U5329 (N_5329,N_2185,N_3154);
and U5330 (N_5330,N_2326,N_2892);
or U5331 (N_5331,N_3261,N_3247);
and U5332 (N_5332,N_3976,N_3864);
nor U5333 (N_5333,N_2183,N_3368);
nor U5334 (N_5334,N_2179,N_2363);
xnor U5335 (N_5335,N_2534,N_2381);
nand U5336 (N_5336,N_3537,N_2627);
nand U5337 (N_5337,N_2447,N_3900);
or U5338 (N_5338,N_3978,N_3605);
xor U5339 (N_5339,N_2202,N_2221);
nor U5340 (N_5340,N_2854,N_3497);
nor U5341 (N_5341,N_2509,N_3164);
nand U5342 (N_5342,N_3614,N_2926);
nand U5343 (N_5343,N_2082,N_2220);
nor U5344 (N_5344,N_2052,N_3242);
and U5345 (N_5345,N_2180,N_3610);
nor U5346 (N_5346,N_2907,N_2427);
xnor U5347 (N_5347,N_3983,N_3318);
xor U5348 (N_5348,N_3663,N_3159);
nor U5349 (N_5349,N_2302,N_3673);
or U5350 (N_5350,N_2134,N_3174);
nor U5351 (N_5351,N_3466,N_3728);
xor U5352 (N_5352,N_3677,N_2789);
nor U5353 (N_5353,N_3439,N_2725);
nand U5354 (N_5354,N_3787,N_3577);
nor U5355 (N_5355,N_3802,N_2562);
xor U5356 (N_5356,N_3192,N_3410);
xor U5357 (N_5357,N_2761,N_3817);
nand U5358 (N_5358,N_2930,N_3819);
or U5359 (N_5359,N_2480,N_3123);
and U5360 (N_5360,N_2007,N_2801);
or U5361 (N_5361,N_2808,N_3392);
xor U5362 (N_5362,N_2133,N_3676);
nor U5363 (N_5363,N_3616,N_3179);
xnor U5364 (N_5364,N_3576,N_2319);
and U5365 (N_5365,N_3473,N_2510);
or U5366 (N_5366,N_3889,N_3755);
and U5367 (N_5367,N_2547,N_3444);
nand U5368 (N_5368,N_3789,N_3368);
and U5369 (N_5369,N_2901,N_2568);
nor U5370 (N_5370,N_3786,N_3578);
nand U5371 (N_5371,N_3527,N_2209);
nand U5372 (N_5372,N_3076,N_2092);
nor U5373 (N_5373,N_2248,N_2246);
nor U5374 (N_5374,N_3460,N_3166);
or U5375 (N_5375,N_3907,N_2387);
nand U5376 (N_5376,N_3814,N_2743);
nor U5377 (N_5377,N_3475,N_3362);
and U5378 (N_5378,N_2370,N_3861);
nand U5379 (N_5379,N_2428,N_2391);
and U5380 (N_5380,N_3568,N_3046);
nor U5381 (N_5381,N_3590,N_2867);
nand U5382 (N_5382,N_3255,N_3161);
xor U5383 (N_5383,N_2366,N_2122);
xnor U5384 (N_5384,N_2344,N_2843);
and U5385 (N_5385,N_2080,N_2124);
nor U5386 (N_5386,N_2370,N_2679);
nand U5387 (N_5387,N_2517,N_2993);
and U5388 (N_5388,N_3694,N_3309);
xnor U5389 (N_5389,N_2018,N_2184);
nand U5390 (N_5390,N_3404,N_2316);
nor U5391 (N_5391,N_3167,N_3281);
nor U5392 (N_5392,N_3154,N_3899);
and U5393 (N_5393,N_2415,N_3889);
xor U5394 (N_5394,N_3080,N_3051);
and U5395 (N_5395,N_2804,N_2904);
nand U5396 (N_5396,N_2352,N_2227);
nand U5397 (N_5397,N_3388,N_3979);
and U5398 (N_5398,N_2122,N_2423);
nand U5399 (N_5399,N_2845,N_3043);
nand U5400 (N_5400,N_3529,N_2057);
and U5401 (N_5401,N_2252,N_3960);
xor U5402 (N_5402,N_3433,N_3079);
nand U5403 (N_5403,N_2330,N_2277);
nor U5404 (N_5404,N_3282,N_3072);
and U5405 (N_5405,N_2306,N_2479);
nor U5406 (N_5406,N_3321,N_3915);
or U5407 (N_5407,N_3786,N_2054);
nand U5408 (N_5408,N_3795,N_2099);
nor U5409 (N_5409,N_3503,N_2634);
and U5410 (N_5410,N_3764,N_3972);
xnor U5411 (N_5411,N_2563,N_2333);
nor U5412 (N_5412,N_3519,N_2595);
nor U5413 (N_5413,N_3817,N_2420);
xnor U5414 (N_5414,N_2760,N_3133);
nor U5415 (N_5415,N_2357,N_2787);
nor U5416 (N_5416,N_3555,N_3503);
nand U5417 (N_5417,N_3081,N_2002);
nand U5418 (N_5418,N_2610,N_2506);
nor U5419 (N_5419,N_3719,N_2784);
and U5420 (N_5420,N_2831,N_2598);
nand U5421 (N_5421,N_2959,N_2606);
or U5422 (N_5422,N_3432,N_2282);
nand U5423 (N_5423,N_3224,N_2893);
nor U5424 (N_5424,N_3396,N_2061);
xor U5425 (N_5425,N_3185,N_2901);
nor U5426 (N_5426,N_3807,N_2228);
or U5427 (N_5427,N_2296,N_2914);
nand U5428 (N_5428,N_2629,N_3917);
and U5429 (N_5429,N_3194,N_3681);
or U5430 (N_5430,N_3587,N_3040);
nor U5431 (N_5431,N_3142,N_3765);
nor U5432 (N_5432,N_3040,N_2166);
and U5433 (N_5433,N_2389,N_3511);
nand U5434 (N_5434,N_2739,N_2238);
or U5435 (N_5435,N_3792,N_3655);
nand U5436 (N_5436,N_2792,N_3315);
or U5437 (N_5437,N_2104,N_3479);
nand U5438 (N_5438,N_2699,N_2980);
and U5439 (N_5439,N_2958,N_3399);
nand U5440 (N_5440,N_2501,N_2751);
and U5441 (N_5441,N_2225,N_3715);
xnor U5442 (N_5442,N_2030,N_3686);
nand U5443 (N_5443,N_3996,N_2611);
nand U5444 (N_5444,N_3831,N_2067);
and U5445 (N_5445,N_2269,N_3492);
nor U5446 (N_5446,N_2026,N_2005);
and U5447 (N_5447,N_3294,N_3244);
nor U5448 (N_5448,N_2065,N_2299);
and U5449 (N_5449,N_2252,N_2181);
xnor U5450 (N_5450,N_3449,N_3286);
and U5451 (N_5451,N_3999,N_3746);
and U5452 (N_5452,N_3173,N_3993);
and U5453 (N_5453,N_3208,N_3859);
or U5454 (N_5454,N_3378,N_2704);
or U5455 (N_5455,N_2759,N_2087);
xor U5456 (N_5456,N_2263,N_3828);
nor U5457 (N_5457,N_2576,N_2812);
nand U5458 (N_5458,N_2769,N_2381);
and U5459 (N_5459,N_3607,N_3075);
xor U5460 (N_5460,N_3633,N_2865);
xor U5461 (N_5461,N_2115,N_2843);
and U5462 (N_5462,N_2019,N_2462);
and U5463 (N_5463,N_3011,N_2718);
xnor U5464 (N_5464,N_2754,N_3327);
and U5465 (N_5465,N_3375,N_2653);
and U5466 (N_5466,N_3049,N_3037);
or U5467 (N_5467,N_2331,N_2907);
xnor U5468 (N_5468,N_3902,N_2998);
nor U5469 (N_5469,N_2354,N_2088);
and U5470 (N_5470,N_3073,N_3322);
or U5471 (N_5471,N_3567,N_2536);
xor U5472 (N_5472,N_3909,N_2651);
or U5473 (N_5473,N_3849,N_3066);
or U5474 (N_5474,N_3805,N_3011);
nand U5475 (N_5475,N_3492,N_2948);
nor U5476 (N_5476,N_2760,N_3392);
nor U5477 (N_5477,N_3500,N_2720);
nand U5478 (N_5478,N_3114,N_2455);
nor U5479 (N_5479,N_2122,N_2348);
and U5480 (N_5480,N_2065,N_2087);
and U5481 (N_5481,N_3960,N_2832);
and U5482 (N_5482,N_3042,N_3155);
nor U5483 (N_5483,N_2120,N_2177);
nor U5484 (N_5484,N_3515,N_3854);
and U5485 (N_5485,N_2683,N_2687);
xor U5486 (N_5486,N_3371,N_3394);
and U5487 (N_5487,N_2553,N_3637);
and U5488 (N_5488,N_2352,N_2030);
nor U5489 (N_5489,N_3420,N_3102);
nor U5490 (N_5490,N_3832,N_3578);
or U5491 (N_5491,N_2212,N_3878);
or U5492 (N_5492,N_3227,N_2879);
xor U5493 (N_5493,N_3941,N_2357);
nand U5494 (N_5494,N_2329,N_2752);
and U5495 (N_5495,N_3082,N_3950);
and U5496 (N_5496,N_3711,N_3858);
nor U5497 (N_5497,N_2418,N_2953);
xnor U5498 (N_5498,N_2818,N_2447);
xor U5499 (N_5499,N_3499,N_2377);
nor U5500 (N_5500,N_2171,N_2521);
and U5501 (N_5501,N_2326,N_2714);
nand U5502 (N_5502,N_2489,N_2435);
or U5503 (N_5503,N_2192,N_2191);
nor U5504 (N_5504,N_3730,N_2745);
nor U5505 (N_5505,N_2261,N_3055);
nand U5506 (N_5506,N_3962,N_3652);
xor U5507 (N_5507,N_2857,N_2431);
or U5508 (N_5508,N_2200,N_3351);
nor U5509 (N_5509,N_2476,N_3867);
xnor U5510 (N_5510,N_3116,N_2135);
nor U5511 (N_5511,N_3082,N_2590);
xor U5512 (N_5512,N_3132,N_3062);
or U5513 (N_5513,N_3081,N_3080);
nor U5514 (N_5514,N_2315,N_2794);
xor U5515 (N_5515,N_3157,N_3977);
and U5516 (N_5516,N_2931,N_2938);
nor U5517 (N_5517,N_3289,N_3612);
nand U5518 (N_5518,N_3699,N_2593);
xnor U5519 (N_5519,N_2895,N_2172);
nor U5520 (N_5520,N_3711,N_2330);
or U5521 (N_5521,N_2998,N_3794);
nor U5522 (N_5522,N_2199,N_2180);
nand U5523 (N_5523,N_3498,N_3835);
nand U5524 (N_5524,N_2905,N_3375);
xor U5525 (N_5525,N_2918,N_3710);
xnor U5526 (N_5526,N_2669,N_3174);
xor U5527 (N_5527,N_3034,N_3232);
nand U5528 (N_5528,N_3907,N_2907);
nand U5529 (N_5529,N_2210,N_3264);
and U5530 (N_5530,N_3299,N_2447);
xnor U5531 (N_5531,N_3250,N_2584);
xor U5532 (N_5532,N_2216,N_3655);
xor U5533 (N_5533,N_2792,N_2698);
xor U5534 (N_5534,N_3184,N_3114);
nand U5535 (N_5535,N_3130,N_2955);
nand U5536 (N_5536,N_2171,N_3022);
or U5537 (N_5537,N_3257,N_2161);
or U5538 (N_5538,N_3922,N_3526);
xnor U5539 (N_5539,N_2911,N_3768);
xor U5540 (N_5540,N_2021,N_2250);
or U5541 (N_5541,N_3667,N_2081);
nor U5542 (N_5542,N_3715,N_3174);
and U5543 (N_5543,N_3964,N_3691);
or U5544 (N_5544,N_3564,N_3026);
nor U5545 (N_5545,N_3811,N_2138);
nand U5546 (N_5546,N_2826,N_3876);
and U5547 (N_5547,N_2018,N_2610);
xnor U5548 (N_5548,N_2296,N_2268);
xor U5549 (N_5549,N_2208,N_2356);
and U5550 (N_5550,N_3356,N_3914);
and U5551 (N_5551,N_2001,N_3996);
xor U5552 (N_5552,N_2904,N_2294);
and U5553 (N_5553,N_2026,N_2596);
and U5554 (N_5554,N_2665,N_2028);
xnor U5555 (N_5555,N_2199,N_3100);
xor U5556 (N_5556,N_2058,N_2728);
nand U5557 (N_5557,N_3816,N_3566);
and U5558 (N_5558,N_2701,N_2748);
nor U5559 (N_5559,N_3076,N_3646);
nor U5560 (N_5560,N_3947,N_3562);
or U5561 (N_5561,N_2721,N_3517);
nand U5562 (N_5562,N_3060,N_2182);
and U5563 (N_5563,N_3309,N_2337);
and U5564 (N_5564,N_2012,N_3705);
or U5565 (N_5565,N_3509,N_2110);
and U5566 (N_5566,N_2989,N_3274);
or U5567 (N_5567,N_2453,N_2292);
nand U5568 (N_5568,N_2858,N_2826);
xor U5569 (N_5569,N_2052,N_2721);
or U5570 (N_5570,N_3506,N_2136);
and U5571 (N_5571,N_3380,N_2038);
and U5572 (N_5572,N_3500,N_3023);
and U5573 (N_5573,N_2724,N_2380);
nor U5574 (N_5574,N_3404,N_2676);
or U5575 (N_5575,N_2478,N_2681);
nor U5576 (N_5576,N_3654,N_2404);
nand U5577 (N_5577,N_2831,N_2538);
nand U5578 (N_5578,N_3189,N_2849);
nor U5579 (N_5579,N_3606,N_3519);
nand U5580 (N_5580,N_3881,N_3211);
nor U5581 (N_5581,N_2902,N_3531);
or U5582 (N_5582,N_3669,N_3061);
or U5583 (N_5583,N_2622,N_2427);
or U5584 (N_5584,N_3636,N_3632);
nand U5585 (N_5585,N_2060,N_2642);
and U5586 (N_5586,N_3684,N_3685);
nor U5587 (N_5587,N_3905,N_2059);
or U5588 (N_5588,N_2412,N_2278);
nor U5589 (N_5589,N_3550,N_3058);
nand U5590 (N_5590,N_2893,N_2113);
and U5591 (N_5591,N_2983,N_3528);
and U5592 (N_5592,N_3890,N_3442);
nor U5593 (N_5593,N_3278,N_3570);
nand U5594 (N_5594,N_3748,N_2889);
or U5595 (N_5595,N_3628,N_3198);
and U5596 (N_5596,N_3520,N_2651);
and U5597 (N_5597,N_2629,N_3850);
nor U5598 (N_5598,N_2045,N_3327);
or U5599 (N_5599,N_2939,N_2503);
xor U5600 (N_5600,N_3355,N_3668);
and U5601 (N_5601,N_3265,N_3721);
nor U5602 (N_5602,N_3055,N_2643);
nand U5603 (N_5603,N_2797,N_2934);
and U5604 (N_5604,N_2246,N_3435);
and U5605 (N_5605,N_2701,N_3392);
nand U5606 (N_5606,N_3625,N_2761);
nand U5607 (N_5607,N_2887,N_2741);
or U5608 (N_5608,N_3452,N_3875);
or U5609 (N_5609,N_3317,N_2559);
or U5610 (N_5610,N_3162,N_3274);
xor U5611 (N_5611,N_3046,N_3368);
or U5612 (N_5612,N_2131,N_3850);
or U5613 (N_5613,N_3859,N_2231);
xor U5614 (N_5614,N_2452,N_2425);
nor U5615 (N_5615,N_2302,N_3167);
and U5616 (N_5616,N_3102,N_3941);
or U5617 (N_5617,N_3844,N_2919);
or U5618 (N_5618,N_2927,N_3116);
and U5619 (N_5619,N_3733,N_2777);
nand U5620 (N_5620,N_2100,N_3914);
or U5621 (N_5621,N_3295,N_2389);
nor U5622 (N_5622,N_3416,N_3880);
nor U5623 (N_5623,N_3539,N_2491);
nor U5624 (N_5624,N_3469,N_3064);
and U5625 (N_5625,N_2179,N_3281);
xnor U5626 (N_5626,N_3110,N_2882);
and U5627 (N_5627,N_3402,N_3455);
nand U5628 (N_5628,N_3290,N_3900);
nand U5629 (N_5629,N_3356,N_2388);
or U5630 (N_5630,N_3132,N_2785);
nand U5631 (N_5631,N_2958,N_2176);
xnor U5632 (N_5632,N_2186,N_2678);
xnor U5633 (N_5633,N_3327,N_3181);
and U5634 (N_5634,N_3245,N_2589);
and U5635 (N_5635,N_2220,N_3796);
and U5636 (N_5636,N_3942,N_2423);
nor U5637 (N_5637,N_2902,N_2628);
or U5638 (N_5638,N_3669,N_3937);
nor U5639 (N_5639,N_2211,N_3058);
nand U5640 (N_5640,N_2162,N_3473);
nor U5641 (N_5641,N_2703,N_2102);
or U5642 (N_5642,N_3053,N_2938);
and U5643 (N_5643,N_3747,N_2339);
xor U5644 (N_5644,N_3659,N_2309);
or U5645 (N_5645,N_3176,N_2692);
and U5646 (N_5646,N_2875,N_2690);
xor U5647 (N_5647,N_2721,N_2505);
nand U5648 (N_5648,N_2525,N_2527);
nor U5649 (N_5649,N_3299,N_3568);
or U5650 (N_5650,N_3002,N_2069);
xor U5651 (N_5651,N_3366,N_2275);
xor U5652 (N_5652,N_2648,N_3071);
or U5653 (N_5653,N_2892,N_2121);
or U5654 (N_5654,N_3030,N_2369);
or U5655 (N_5655,N_2327,N_3940);
nand U5656 (N_5656,N_3435,N_2909);
or U5657 (N_5657,N_2766,N_3186);
nor U5658 (N_5658,N_2121,N_3505);
nand U5659 (N_5659,N_2552,N_3969);
and U5660 (N_5660,N_3847,N_3234);
xnor U5661 (N_5661,N_2324,N_3323);
nand U5662 (N_5662,N_2740,N_2074);
or U5663 (N_5663,N_2552,N_3829);
and U5664 (N_5664,N_2486,N_2281);
nor U5665 (N_5665,N_3239,N_2920);
nand U5666 (N_5666,N_2653,N_3251);
xor U5667 (N_5667,N_3339,N_2592);
and U5668 (N_5668,N_3679,N_3775);
and U5669 (N_5669,N_3964,N_3180);
xor U5670 (N_5670,N_2542,N_2512);
nand U5671 (N_5671,N_2820,N_3852);
and U5672 (N_5672,N_2419,N_3258);
or U5673 (N_5673,N_2166,N_3411);
or U5674 (N_5674,N_2716,N_3763);
and U5675 (N_5675,N_3774,N_3057);
or U5676 (N_5676,N_2980,N_3290);
nor U5677 (N_5677,N_2552,N_2186);
and U5678 (N_5678,N_2955,N_2663);
or U5679 (N_5679,N_2677,N_2064);
nand U5680 (N_5680,N_2358,N_2943);
or U5681 (N_5681,N_3848,N_2638);
nand U5682 (N_5682,N_3492,N_2993);
nand U5683 (N_5683,N_2275,N_2962);
or U5684 (N_5684,N_3576,N_3121);
nand U5685 (N_5685,N_2372,N_2689);
nand U5686 (N_5686,N_2471,N_3581);
xnor U5687 (N_5687,N_3819,N_2322);
and U5688 (N_5688,N_3841,N_3914);
or U5689 (N_5689,N_2447,N_3858);
or U5690 (N_5690,N_3485,N_2084);
and U5691 (N_5691,N_3752,N_2304);
nor U5692 (N_5692,N_2851,N_2214);
nor U5693 (N_5693,N_2319,N_2763);
nand U5694 (N_5694,N_3768,N_2021);
xor U5695 (N_5695,N_2072,N_3710);
or U5696 (N_5696,N_3009,N_2726);
xnor U5697 (N_5697,N_3163,N_2870);
nor U5698 (N_5698,N_2767,N_3255);
nand U5699 (N_5699,N_3349,N_2515);
xnor U5700 (N_5700,N_3844,N_2669);
xor U5701 (N_5701,N_2122,N_2911);
and U5702 (N_5702,N_2768,N_3050);
nand U5703 (N_5703,N_3793,N_2849);
or U5704 (N_5704,N_2227,N_3846);
xnor U5705 (N_5705,N_3978,N_2934);
xor U5706 (N_5706,N_2703,N_2234);
nand U5707 (N_5707,N_2482,N_2455);
nand U5708 (N_5708,N_2617,N_2498);
or U5709 (N_5709,N_3036,N_3574);
xor U5710 (N_5710,N_2618,N_3316);
nor U5711 (N_5711,N_3041,N_2685);
nand U5712 (N_5712,N_2463,N_3924);
or U5713 (N_5713,N_2746,N_2213);
nand U5714 (N_5714,N_2508,N_3993);
nor U5715 (N_5715,N_2847,N_2719);
or U5716 (N_5716,N_2800,N_2132);
nand U5717 (N_5717,N_3668,N_2582);
or U5718 (N_5718,N_2557,N_3022);
nand U5719 (N_5719,N_2414,N_3631);
xnor U5720 (N_5720,N_3464,N_2161);
nor U5721 (N_5721,N_3538,N_3756);
and U5722 (N_5722,N_3125,N_2139);
nor U5723 (N_5723,N_2323,N_3029);
and U5724 (N_5724,N_2260,N_2086);
nor U5725 (N_5725,N_3841,N_2280);
xor U5726 (N_5726,N_2868,N_2422);
xor U5727 (N_5727,N_2668,N_3122);
nor U5728 (N_5728,N_2786,N_3030);
nor U5729 (N_5729,N_3652,N_2247);
and U5730 (N_5730,N_3757,N_2302);
xnor U5731 (N_5731,N_3582,N_2170);
and U5732 (N_5732,N_3593,N_2332);
and U5733 (N_5733,N_2814,N_2683);
or U5734 (N_5734,N_3843,N_2898);
nor U5735 (N_5735,N_3208,N_2934);
or U5736 (N_5736,N_3883,N_2712);
nor U5737 (N_5737,N_3944,N_3599);
nor U5738 (N_5738,N_2969,N_2362);
xor U5739 (N_5739,N_3830,N_2064);
nand U5740 (N_5740,N_3169,N_2088);
xnor U5741 (N_5741,N_3511,N_2223);
or U5742 (N_5742,N_2075,N_2330);
nand U5743 (N_5743,N_3247,N_2210);
nor U5744 (N_5744,N_3123,N_3080);
and U5745 (N_5745,N_3431,N_3729);
nand U5746 (N_5746,N_2802,N_2640);
nor U5747 (N_5747,N_2882,N_3571);
xnor U5748 (N_5748,N_2057,N_2777);
nor U5749 (N_5749,N_3740,N_2281);
nor U5750 (N_5750,N_2021,N_3281);
and U5751 (N_5751,N_2900,N_3163);
xnor U5752 (N_5752,N_2610,N_3340);
nand U5753 (N_5753,N_3601,N_3845);
xor U5754 (N_5754,N_2635,N_2017);
and U5755 (N_5755,N_3831,N_3611);
or U5756 (N_5756,N_2411,N_2352);
or U5757 (N_5757,N_2185,N_2426);
xnor U5758 (N_5758,N_2293,N_3764);
nand U5759 (N_5759,N_3598,N_2281);
xor U5760 (N_5760,N_3316,N_2006);
nor U5761 (N_5761,N_3533,N_2005);
xnor U5762 (N_5762,N_2014,N_2638);
nand U5763 (N_5763,N_2185,N_3061);
nor U5764 (N_5764,N_2287,N_3583);
and U5765 (N_5765,N_3513,N_3915);
xor U5766 (N_5766,N_2334,N_3977);
xor U5767 (N_5767,N_3095,N_2330);
and U5768 (N_5768,N_2564,N_2578);
xnor U5769 (N_5769,N_2326,N_3336);
and U5770 (N_5770,N_2205,N_3312);
or U5771 (N_5771,N_2530,N_2184);
or U5772 (N_5772,N_2123,N_3819);
and U5773 (N_5773,N_2477,N_2464);
nor U5774 (N_5774,N_3978,N_3195);
or U5775 (N_5775,N_2700,N_2369);
nor U5776 (N_5776,N_2937,N_3574);
xor U5777 (N_5777,N_3687,N_3864);
and U5778 (N_5778,N_2576,N_2238);
xor U5779 (N_5779,N_3202,N_3290);
xor U5780 (N_5780,N_2269,N_2326);
nor U5781 (N_5781,N_2276,N_2172);
and U5782 (N_5782,N_2740,N_2574);
nor U5783 (N_5783,N_3479,N_2180);
nand U5784 (N_5784,N_2724,N_3833);
and U5785 (N_5785,N_2207,N_3167);
xnor U5786 (N_5786,N_2274,N_2490);
nor U5787 (N_5787,N_3517,N_3873);
or U5788 (N_5788,N_2234,N_2539);
xor U5789 (N_5789,N_3424,N_2456);
nor U5790 (N_5790,N_2060,N_2108);
and U5791 (N_5791,N_2832,N_2393);
nand U5792 (N_5792,N_2995,N_2135);
nor U5793 (N_5793,N_2755,N_3994);
nand U5794 (N_5794,N_2453,N_3630);
and U5795 (N_5795,N_3840,N_3126);
or U5796 (N_5796,N_2329,N_2775);
nand U5797 (N_5797,N_3879,N_2543);
xnor U5798 (N_5798,N_3423,N_3526);
or U5799 (N_5799,N_2618,N_3166);
or U5800 (N_5800,N_2238,N_3455);
and U5801 (N_5801,N_2476,N_3195);
nor U5802 (N_5802,N_3682,N_2116);
xor U5803 (N_5803,N_2009,N_2280);
nor U5804 (N_5804,N_3042,N_3812);
nor U5805 (N_5805,N_2753,N_2593);
and U5806 (N_5806,N_3071,N_3866);
and U5807 (N_5807,N_3108,N_3313);
nor U5808 (N_5808,N_3415,N_2490);
nor U5809 (N_5809,N_2436,N_3139);
nand U5810 (N_5810,N_2268,N_2977);
xnor U5811 (N_5811,N_2785,N_3029);
xor U5812 (N_5812,N_3941,N_2654);
or U5813 (N_5813,N_2069,N_2252);
nand U5814 (N_5814,N_3788,N_3736);
nand U5815 (N_5815,N_2534,N_2257);
nand U5816 (N_5816,N_2952,N_2093);
or U5817 (N_5817,N_3109,N_2469);
nand U5818 (N_5818,N_2447,N_2241);
or U5819 (N_5819,N_3037,N_2885);
nand U5820 (N_5820,N_2257,N_2846);
nand U5821 (N_5821,N_3302,N_3202);
or U5822 (N_5822,N_3378,N_3482);
nor U5823 (N_5823,N_3662,N_2550);
and U5824 (N_5824,N_3523,N_3655);
nand U5825 (N_5825,N_3894,N_2826);
xor U5826 (N_5826,N_3859,N_2717);
nor U5827 (N_5827,N_2006,N_2918);
or U5828 (N_5828,N_2639,N_3723);
nor U5829 (N_5829,N_3612,N_3687);
and U5830 (N_5830,N_2730,N_3405);
xor U5831 (N_5831,N_2563,N_3188);
or U5832 (N_5832,N_3345,N_2506);
or U5833 (N_5833,N_2273,N_3929);
or U5834 (N_5834,N_2732,N_2213);
nand U5835 (N_5835,N_3437,N_3936);
or U5836 (N_5836,N_3445,N_2808);
and U5837 (N_5837,N_3008,N_2169);
and U5838 (N_5838,N_3787,N_2299);
nor U5839 (N_5839,N_3382,N_2412);
nand U5840 (N_5840,N_2545,N_3188);
and U5841 (N_5841,N_2181,N_3509);
nor U5842 (N_5842,N_3268,N_3309);
xnor U5843 (N_5843,N_3133,N_3485);
nor U5844 (N_5844,N_2248,N_3065);
and U5845 (N_5845,N_3312,N_2179);
nand U5846 (N_5846,N_2152,N_3894);
nor U5847 (N_5847,N_3934,N_2409);
xnor U5848 (N_5848,N_3982,N_3827);
and U5849 (N_5849,N_3560,N_3547);
nand U5850 (N_5850,N_3319,N_2297);
and U5851 (N_5851,N_2170,N_3777);
and U5852 (N_5852,N_2218,N_3541);
xnor U5853 (N_5853,N_2030,N_3771);
and U5854 (N_5854,N_2000,N_3316);
nor U5855 (N_5855,N_3542,N_3527);
or U5856 (N_5856,N_2913,N_3318);
xnor U5857 (N_5857,N_3979,N_2615);
nand U5858 (N_5858,N_2069,N_3917);
nand U5859 (N_5859,N_2600,N_3768);
and U5860 (N_5860,N_3197,N_3971);
or U5861 (N_5861,N_2672,N_3275);
nand U5862 (N_5862,N_2576,N_3538);
xor U5863 (N_5863,N_3234,N_3031);
xor U5864 (N_5864,N_2636,N_2781);
nand U5865 (N_5865,N_2260,N_3360);
nand U5866 (N_5866,N_3107,N_2321);
nor U5867 (N_5867,N_2871,N_3604);
xor U5868 (N_5868,N_3240,N_3054);
and U5869 (N_5869,N_2859,N_2306);
and U5870 (N_5870,N_3596,N_2594);
or U5871 (N_5871,N_3863,N_2413);
and U5872 (N_5872,N_3498,N_2732);
nand U5873 (N_5873,N_2327,N_2333);
nand U5874 (N_5874,N_3752,N_3148);
or U5875 (N_5875,N_3832,N_2942);
nor U5876 (N_5876,N_2879,N_2643);
or U5877 (N_5877,N_3718,N_3651);
nor U5878 (N_5878,N_3091,N_2566);
or U5879 (N_5879,N_3227,N_3919);
and U5880 (N_5880,N_2537,N_2259);
and U5881 (N_5881,N_2683,N_2507);
nor U5882 (N_5882,N_2686,N_2872);
xor U5883 (N_5883,N_3522,N_3381);
nand U5884 (N_5884,N_2062,N_3928);
or U5885 (N_5885,N_3940,N_3338);
nand U5886 (N_5886,N_3458,N_3926);
and U5887 (N_5887,N_3724,N_2931);
xor U5888 (N_5888,N_3019,N_2527);
and U5889 (N_5889,N_2220,N_2180);
xnor U5890 (N_5890,N_3288,N_2276);
xor U5891 (N_5891,N_2168,N_2786);
nand U5892 (N_5892,N_2461,N_3983);
nand U5893 (N_5893,N_2702,N_3129);
nor U5894 (N_5894,N_3683,N_2966);
nand U5895 (N_5895,N_2308,N_3967);
xor U5896 (N_5896,N_2522,N_3449);
or U5897 (N_5897,N_3751,N_2939);
nand U5898 (N_5898,N_3256,N_3651);
and U5899 (N_5899,N_3728,N_3571);
nor U5900 (N_5900,N_3037,N_3890);
nand U5901 (N_5901,N_3017,N_2960);
nor U5902 (N_5902,N_2007,N_3433);
or U5903 (N_5903,N_3823,N_3855);
or U5904 (N_5904,N_3572,N_2859);
nand U5905 (N_5905,N_3795,N_2259);
nand U5906 (N_5906,N_3110,N_2560);
nand U5907 (N_5907,N_3132,N_3933);
xnor U5908 (N_5908,N_3779,N_3325);
nor U5909 (N_5909,N_3096,N_3144);
and U5910 (N_5910,N_2285,N_2110);
nor U5911 (N_5911,N_2744,N_3875);
nor U5912 (N_5912,N_3171,N_3287);
nor U5913 (N_5913,N_2169,N_2221);
nand U5914 (N_5914,N_3907,N_3812);
nor U5915 (N_5915,N_3674,N_2740);
xnor U5916 (N_5916,N_3772,N_3100);
or U5917 (N_5917,N_2767,N_2384);
xnor U5918 (N_5918,N_2808,N_3095);
xnor U5919 (N_5919,N_2015,N_2474);
nor U5920 (N_5920,N_2120,N_2271);
nand U5921 (N_5921,N_2572,N_2419);
or U5922 (N_5922,N_2923,N_3089);
or U5923 (N_5923,N_3906,N_3345);
and U5924 (N_5924,N_3362,N_3945);
xnor U5925 (N_5925,N_3826,N_3374);
xor U5926 (N_5926,N_2482,N_3873);
nand U5927 (N_5927,N_2697,N_3784);
nand U5928 (N_5928,N_2459,N_2306);
or U5929 (N_5929,N_2427,N_3358);
xor U5930 (N_5930,N_2422,N_2589);
and U5931 (N_5931,N_2810,N_3595);
and U5932 (N_5932,N_3190,N_2402);
nor U5933 (N_5933,N_2718,N_3129);
nand U5934 (N_5934,N_3211,N_2168);
or U5935 (N_5935,N_3629,N_2168);
xor U5936 (N_5936,N_3140,N_3300);
nand U5937 (N_5937,N_2113,N_3357);
and U5938 (N_5938,N_3871,N_3044);
or U5939 (N_5939,N_2460,N_3974);
nand U5940 (N_5940,N_2319,N_3808);
or U5941 (N_5941,N_2227,N_3664);
nor U5942 (N_5942,N_3971,N_2207);
or U5943 (N_5943,N_3161,N_2284);
xnor U5944 (N_5944,N_2828,N_2856);
or U5945 (N_5945,N_2583,N_2064);
nor U5946 (N_5946,N_2229,N_3129);
nand U5947 (N_5947,N_2313,N_2769);
and U5948 (N_5948,N_3911,N_2352);
nand U5949 (N_5949,N_2334,N_2485);
nand U5950 (N_5950,N_3933,N_3857);
or U5951 (N_5951,N_2937,N_2887);
xor U5952 (N_5952,N_3335,N_2226);
and U5953 (N_5953,N_2796,N_2922);
xnor U5954 (N_5954,N_3372,N_3455);
nand U5955 (N_5955,N_3535,N_2741);
and U5956 (N_5956,N_3504,N_2811);
and U5957 (N_5957,N_2888,N_3936);
xor U5958 (N_5958,N_2008,N_2222);
or U5959 (N_5959,N_3429,N_2896);
nand U5960 (N_5960,N_2160,N_3552);
nor U5961 (N_5961,N_3199,N_2870);
nand U5962 (N_5962,N_3095,N_3829);
xnor U5963 (N_5963,N_3296,N_2681);
and U5964 (N_5964,N_3995,N_2719);
or U5965 (N_5965,N_3994,N_3321);
and U5966 (N_5966,N_3137,N_3640);
and U5967 (N_5967,N_2597,N_2395);
xnor U5968 (N_5968,N_3812,N_3423);
nand U5969 (N_5969,N_3020,N_3142);
nand U5970 (N_5970,N_2818,N_2372);
and U5971 (N_5971,N_2010,N_2942);
and U5972 (N_5972,N_3253,N_3533);
xnor U5973 (N_5973,N_3240,N_3034);
xnor U5974 (N_5974,N_2639,N_2677);
and U5975 (N_5975,N_3775,N_3110);
xor U5976 (N_5976,N_2873,N_3274);
xnor U5977 (N_5977,N_2637,N_2448);
xor U5978 (N_5978,N_2496,N_2573);
xor U5979 (N_5979,N_2857,N_2398);
nor U5980 (N_5980,N_3888,N_3069);
or U5981 (N_5981,N_3472,N_2207);
and U5982 (N_5982,N_2153,N_3442);
nand U5983 (N_5983,N_3134,N_3385);
nand U5984 (N_5984,N_3250,N_3097);
xnor U5985 (N_5985,N_3678,N_2743);
nand U5986 (N_5986,N_3699,N_3751);
nor U5987 (N_5987,N_2192,N_3755);
and U5988 (N_5988,N_2369,N_3877);
and U5989 (N_5989,N_2803,N_3641);
xor U5990 (N_5990,N_2053,N_3356);
nand U5991 (N_5991,N_2742,N_3692);
xnor U5992 (N_5992,N_3360,N_3988);
and U5993 (N_5993,N_2372,N_3540);
and U5994 (N_5994,N_2755,N_3194);
and U5995 (N_5995,N_2302,N_3042);
or U5996 (N_5996,N_3615,N_3172);
xor U5997 (N_5997,N_3758,N_2148);
nand U5998 (N_5998,N_2159,N_2280);
and U5999 (N_5999,N_3134,N_2064);
or U6000 (N_6000,N_5282,N_5102);
and U6001 (N_6001,N_5040,N_4802);
and U6002 (N_6002,N_5112,N_4959);
or U6003 (N_6003,N_4638,N_5538);
xnor U6004 (N_6004,N_5274,N_4907);
or U6005 (N_6005,N_5150,N_5350);
nor U6006 (N_6006,N_5823,N_4604);
and U6007 (N_6007,N_5595,N_5807);
or U6008 (N_6008,N_4986,N_4195);
and U6009 (N_6009,N_4215,N_4019);
nand U6010 (N_6010,N_4782,N_4749);
and U6011 (N_6011,N_5370,N_5141);
xor U6012 (N_6012,N_5652,N_4819);
or U6013 (N_6013,N_5613,N_4866);
nand U6014 (N_6014,N_4261,N_5531);
and U6015 (N_6015,N_5480,N_4091);
nor U6016 (N_6016,N_5001,N_4614);
or U6017 (N_6017,N_5589,N_5748);
or U6018 (N_6018,N_5263,N_4369);
and U6019 (N_6019,N_4750,N_4473);
xnor U6020 (N_6020,N_4378,N_5320);
or U6021 (N_6021,N_4271,N_4376);
or U6022 (N_6022,N_5573,N_4021);
xnor U6023 (N_6023,N_5325,N_5798);
nor U6024 (N_6024,N_4260,N_4106);
nand U6025 (N_6025,N_5215,N_4384);
or U6026 (N_6026,N_4694,N_5338);
nor U6027 (N_6027,N_4512,N_5007);
nand U6028 (N_6028,N_5657,N_5433);
xor U6029 (N_6029,N_5624,N_5683);
nand U6030 (N_6030,N_5923,N_4067);
or U6031 (N_6031,N_5138,N_4223);
and U6032 (N_6032,N_4693,N_4045);
nand U6033 (N_6033,N_5241,N_5444);
or U6034 (N_6034,N_4014,N_4930);
and U6035 (N_6035,N_4781,N_4504);
and U6036 (N_6036,N_4375,N_5261);
xor U6037 (N_6037,N_5213,N_5121);
xnor U6038 (N_6038,N_5938,N_5580);
xnor U6039 (N_6039,N_5786,N_5578);
or U6040 (N_6040,N_5388,N_4560);
nand U6041 (N_6041,N_4400,N_4851);
or U6042 (N_6042,N_5742,N_5303);
nor U6043 (N_6043,N_5954,N_4258);
and U6044 (N_6044,N_5010,N_4649);
nor U6045 (N_6045,N_4336,N_4612);
and U6046 (N_6046,N_4017,N_4575);
nand U6047 (N_6047,N_5249,N_4152);
xnor U6048 (N_6048,N_4104,N_5094);
and U6049 (N_6049,N_5314,N_5077);
or U6050 (N_6050,N_4948,N_5212);
or U6051 (N_6051,N_4797,N_5206);
nand U6052 (N_6052,N_5650,N_5794);
xnor U6053 (N_6053,N_4358,N_4762);
and U6054 (N_6054,N_4643,N_5781);
or U6055 (N_6055,N_5585,N_4134);
nor U6056 (N_6056,N_5855,N_5542);
xor U6057 (N_6057,N_5925,N_5708);
and U6058 (N_6058,N_4310,N_4367);
and U6059 (N_6059,N_5336,N_5686);
xor U6060 (N_6060,N_5266,N_5041);
or U6061 (N_6061,N_4875,N_5571);
nand U6062 (N_6062,N_4572,N_4302);
nor U6063 (N_6063,N_5851,N_4294);
nor U6064 (N_6064,N_5301,N_5161);
xor U6065 (N_6065,N_4999,N_5119);
and U6066 (N_6066,N_5701,N_4777);
nand U6067 (N_6067,N_5557,N_5561);
nand U6068 (N_6068,N_5020,N_5479);
xor U6069 (N_6069,N_4304,N_5791);
nor U6070 (N_6070,N_4549,N_5948);
or U6071 (N_6071,N_4314,N_4641);
or U6072 (N_6072,N_4080,N_5892);
or U6073 (N_6073,N_5057,N_5525);
nand U6074 (N_6074,N_5026,N_5231);
xnor U6075 (N_6075,N_4583,N_4668);
nor U6076 (N_6076,N_5262,N_4318);
and U6077 (N_6077,N_5332,N_5620);
and U6078 (N_6078,N_4900,N_4506);
or U6079 (N_6079,N_5247,N_5098);
nand U6080 (N_6080,N_4899,N_5551);
nor U6081 (N_6081,N_5123,N_4684);
nor U6082 (N_6082,N_5827,N_4611);
or U6083 (N_6083,N_5003,N_5867);
and U6084 (N_6084,N_4074,N_4984);
and U6085 (N_6085,N_5897,N_4626);
xnor U6086 (N_6086,N_5767,N_4130);
or U6087 (N_6087,N_4234,N_4420);
xor U6088 (N_6088,N_5836,N_4574);
nor U6089 (N_6089,N_5167,N_4500);
or U6090 (N_6090,N_5013,N_4128);
xnor U6091 (N_6091,N_4941,N_5185);
nor U6092 (N_6092,N_5083,N_4298);
and U6093 (N_6093,N_4177,N_5464);
nand U6094 (N_6094,N_4517,N_5497);
or U6095 (N_6095,N_5875,N_5016);
nand U6096 (N_6096,N_4450,N_5131);
xor U6097 (N_6097,N_5104,N_5108);
or U6098 (N_6098,N_5698,N_4897);
xor U6099 (N_6099,N_5272,N_5011);
nand U6100 (N_6100,N_4639,N_4100);
nand U6101 (N_6101,N_4590,N_4193);
nor U6102 (N_6102,N_5608,N_4278);
xnor U6103 (N_6103,N_5873,N_5841);
xor U6104 (N_6104,N_4006,N_4410);
and U6105 (N_6105,N_4936,N_5508);
or U6106 (N_6106,N_4228,N_4865);
and U6107 (N_6107,N_5680,N_5177);
nand U6108 (N_6108,N_4446,N_4608);
nand U6109 (N_6109,N_4053,N_5635);
nand U6110 (N_6110,N_5152,N_5244);
and U6111 (N_6111,N_4265,N_4121);
nor U6112 (N_6112,N_5940,N_4279);
and U6113 (N_6113,N_4287,N_4334);
xor U6114 (N_6114,N_4327,N_4343);
nand U6115 (N_6115,N_5059,N_4390);
and U6116 (N_6116,N_4700,N_5801);
xnor U6117 (N_6117,N_5712,N_5991);
nand U6118 (N_6118,N_4386,N_4370);
nor U6119 (N_6119,N_4032,N_5127);
or U6120 (N_6120,N_5824,N_5736);
xor U6121 (N_6121,N_4337,N_4853);
nor U6122 (N_6122,N_4438,N_4084);
and U6123 (N_6123,N_4631,N_4826);
and U6124 (N_6124,N_5988,N_4775);
xnor U6125 (N_6125,N_4116,N_4415);
and U6126 (N_6126,N_5248,N_4515);
nand U6127 (N_6127,N_5245,N_4648);
xor U6128 (N_6128,N_4124,N_5339);
nor U6129 (N_6129,N_5431,N_4994);
or U6130 (N_6130,N_5250,N_4497);
and U6131 (N_6131,N_4451,N_5820);
or U6132 (N_6132,N_4509,N_5176);
nor U6133 (N_6133,N_5151,N_4027);
nand U6134 (N_6134,N_4704,N_4435);
nor U6135 (N_6135,N_4259,N_4389);
nor U6136 (N_6136,N_5258,N_5158);
nor U6137 (N_6137,N_4245,N_5465);
xnor U6138 (N_6138,N_4792,N_5967);
nand U6139 (N_6139,N_5236,N_4022);
nand U6140 (N_6140,N_5481,N_4811);
nor U6141 (N_6141,N_4677,N_5866);
and U6142 (N_6142,N_5027,N_4945);
or U6143 (N_6143,N_5772,N_4498);
or U6144 (N_6144,N_4548,N_4181);
and U6145 (N_6145,N_4711,N_5776);
nand U6146 (N_6146,N_5745,N_5290);
xor U6147 (N_6147,N_4320,N_5037);
nand U6148 (N_6148,N_4013,N_4728);
nand U6149 (N_6149,N_4556,N_5612);
or U6150 (N_6150,N_4541,N_4946);
nor U6151 (N_6151,N_5474,N_4809);
or U6152 (N_6152,N_5628,N_5296);
nand U6153 (N_6153,N_4879,N_4636);
nand U6154 (N_6154,N_4189,N_4492);
xnor U6155 (N_6155,N_4886,N_5472);
or U6156 (N_6156,N_5567,N_4272);
or U6157 (N_6157,N_4605,N_4731);
nor U6158 (N_6158,N_4399,N_4843);
or U6159 (N_6159,N_4666,N_5496);
and U6160 (N_6160,N_4697,N_4081);
nor U6161 (N_6161,N_4413,N_4003);
nand U6162 (N_6162,N_5276,N_4239);
nor U6163 (N_6163,N_5126,N_4606);
nand U6164 (N_6164,N_4250,N_4267);
nor U6165 (N_6165,N_4974,N_5023);
nand U6166 (N_6166,N_5974,N_4913);
xor U6167 (N_6167,N_4800,N_5068);
nand U6168 (N_6168,N_4931,N_5305);
nand U6169 (N_6169,N_5694,N_5868);
or U6170 (N_6170,N_4447,N_5033);
nor U6171 (N_6171,N_4528,N_5936);
nor U6172 (N_6172,N_4197,N_5756);
nor U6173 (N_6173,N_5019,N_4043);
and U6174 (N_6174,N_5584,N_5269);
nand U6175 (N_6175,N_4321,N_4301);
or U6176 (N_6176,N_5294,N_4571);
xor U6177 (N_6177,N_5645,N_4673);
xnor U6178 (N_6178,N_4785,N_5977);
or U6179 (N_6179,N_5616,N_4589);
or U6180 (N_6180,N_5385,N_4524);
nand U6181 (N_6181,N_4566,N_4996);
xnor U6182 (N_6182,N_4980,N_5396);
and U6183 (N_6183,N_4712,N_4915);
nand U6184 (N_6184,N_5216,N_4530);
or U6185 (N_6185,N_4408,N_5467);
or U6186 (N_6186,N_4698,N_4965);
and U6187 (N_6187,N_5529,N_4150);
and U6188 (N_6188,N_4368,N_5420);
and U6189 (N_6189,N_5688,N_5941);
nand U6190 (N_6190,N_4962,N_5513);
or U6191 (N_6191,N_5091,N_4458);
nand U6192 (N_6192,N_4145,N_4854);
or U6193 (N_6193,N_4676,N_4182);
and U6194 (N_6194,N_4881,N_5728);
nand U6195 (N_6195,N_5409,N_5278);
or U6196 (N_6196,N_5195,N_4493);
xnor U6197 (N_6197,N_5775,N_5356);
xnor U6198 (N_6198,N_5644,N_5283);
nand U6199 (N_6199,N_4646,N_5184);
xnor U6200 (N_6200,N_4065,N_4998);
nand U6201 (N_6201,N_4820,N_5872);
or U6202 (N_6202,N_5235,N_5349);
nor U6203 (N_6203,N_4538,N_5082);
nor U6204 (N_6204,N_5207,N_5171);
nand U6205 (N_6205,N_4490,N_5522);
and U6206 (N_6206,N_4448,N_5252);
and U6207 (N_6207,N_5452,N_5975);
xnor U6208 (N_6208,N_5710,N_5267);
or U6209 (N_6209,N_5870,N_5861);
nand U6210 (N_6210,N_4804,N_4041);
and U6211 (N_6211,N_4071,N_5362);
nand U6212 (N_6212,N_4578,N_5572);
nor U6213 (N_6213,N_4817,N_5035);
and U6214 (N_6214,N_5625,N_4277);
nand U6215 (N_6215,N_4703,N_5379);
and U6216 (N_6216,N_5143,N_5166);
nor U6217 (N_6217,N_5074,N_5360);
or U6218 (N_6218,N_4659,N_4387);
nand U6219 (N_6219,N_5711,N_4967);
xor U6220 (N_6220,N_5746,N_4862);
nor U6221 (N_6221,N_5859,N_4202);
and U6222 (N_6222,N_4093,N_4937);
xnor U6223 (N_6223,N_4520,N_5913);
and U6224 (N_6224,N_4786,N_5878);
nor U6225 (N_6225,N_4194,N_4144);
and U6226 (N_6226,N_4374,N_4034);
nand U6227 (N_6227,N_4107,N_5306);
and U6228 (N_6228,N_4254,N_5056);
nor U6229 (N_6229,N_4755,N_4850);
nand U6230 (N_6230,N_4455,N_4233);
and U6231 (N_6231,N_5880,N_4772);
xor U6232 (N_6232,N_4868,N_4395);
and U6233 (N_6233,N_4339,N_4291);
xnor U6234 (N_6234,N_4266,N_5980);
xnor U6235 (N_6235,N_4089,N_4799);
and U6236 (N_6236,N_5257,N_4559);
or U6237 (N_6237,N_5295,N_5512);
and U6238 (N_6238,N_5355,N_4653);
and U6239 (N_6239,N_5502,N_5730);
nand U6240 (N_6240,N_4727,N_5424);
nor U6241 (N_6241,N_4264,N_5456);
nor U6242 (N_6242,N_4838,N_5381);
xnor U6243 (N_6243,N_5631,N_4158);
nor U6244 (N_6244,N_5477,N_4769);
xor U6245 (N_6245,N_4280,N_5051);
and U6246 (N_6246,N_4131,N_4839);
and U6247 (N_6247,N_5753,N_4825);
and U6248 (N_6248,N_5342,N_4122);
or U6249 (N_6249,N_5802,N_5443);
nor U6250 (N_6250,N_5270,N_5142);
or U6251 (N_6251,N_4429,N_4629);
or U6252 (N_6252,N_5982,N_4870);
nand U6253 (N_6253,N_5197,N_5958);
nor U6254 (N_6254,N_5739,N_4437);
or U6255 (N_6255,N_5888,N_5675);
nand U6256 (N_6256,N_5406,N_4169);
or U6257 (N_6257,N_4991,N_4940);
or U6258 (N_6258,N_4184,N_4833);
and U6259 (N_6259,N_5107,N_5667);
nand U6260 (N_6260,N_5829,N_5894);
xnor U6261 (N_6261,N_4592,N_5637);
nor U6262 (N_6262,N_4213,N_4981);
and U6263 (N_6263,N_4315,N_4747);
nand U6264 (N_6264,N_5603,N_5425);
nor U6265 (N_6265,N_4508,N_4029);
or U6266 (N_6266,N_5187,N_4475);
nand U6267 (N_6267,N_5440,N_4411);
xor U6268 (N_6268,N_5163,N_5434);
nor U6269 (N_6269,N_5706,N_5159);
nor U6270 (N_6270,N_5337,N_5676);
and U6271 (N_6271,N_4523,N_5660);
nand U6272 (N_6272,N_4580,N_4964);
and U6273 (N_6273,N_4024,N_4544);
xor U6274 (N_6274,N_5656,N_5760);
and U6275 (N_6275,N_4191,N_4105);
nor U6276 (N_6276,N_4129,N_5576);
or U6277 (N_6277,N_4503,N_4004);
nor U6278 (N_6278,N_5081,N_5854);
nor U6279 (N_6279,N_4163,N_4766);
nand U6280 (N_6280,N_5653,N_4424);
and U6281 (N_6281,N_4114,N_4126);
and U6282 (N_6282,N_4737,N_5032);
xor U6283 (N_6283,N_5633,N_4622);
nor U6284 (N_6284,N_4028,N_5703);
or U6285 (N_6285,N_5254,N_5071);
nor U6286 (N_6286,N_4401,N_5681);
or U6287 (N_6287,N_5953,N_4244);
nand U6288 (N_6288,N_5816,N_4050);
and U6289 (N_6289,N_4642,N_5401);
and U6290 (N_6290,N_4689,N_5462);
and U6291 (N_6291,N_4049,N_4360);
nand U6292 (N_6292,N_5393,N_4655);
or U6293 (N_6293,N_4633,N_5340);
or U6294 (N_6294,N_5981,N_5963);
xnor U6295 (N_6295,N_5933,N_5664);
or U6296 (N_6296,N_5049,N_5815);
or U6297 (N_6297,N_5946,N_4869);
or U6298 (N_6298,N_4779,N_5671);
and U6299 (N_6299,N_4678,N_4922);
nor U6300 (N_6300,N_5907,N_4829);
or U6301 (N_6301,N_5630,N_4474);
nand U6302 (N_6302,N_5034,N_5932);
and U6303 (N_6303,N_5601,N_4674);
xnor U6304 (N_6304,N_4793,N_5788);
nor U6305 (N_6305,N_5234,N_4467);
xor U6306 (N_6306,N_5658,N_5915);
nor U6307 (N_6307,N_4885,N_4031);
nor U6308 (N_6308,N_5436,N_4364);
nand U6309 (N_6309,N_5693,N_5366);
or U6310 (N_6310,N_4351,N_5117);
xnor U6311 (N_6311,N_5281,N_4142);
nor U6312 (N_6312,N_4432,N_5417);
and U6313 (N_6313,N_4292,N_4748);
nand U6314 (N_6314,N_5028,N_4742);
or U6315 (N_6315,N_5521,N_5541);
or U6316 (N_6316,N_4722,N_4361);
xor U6317 (N_6317,N_5917,N_4569);
or U6318 (N_6318,N_5426,N_5376);
and U6319 (N_6319,N_4925,N_4060);
and U6320 (N_6320,N_5455,N_5715);
nand U6321 (N_6321,N_4086,N_4909);
nor U6322 (N_6322,N_4919,N_4317);
nor U6323 (N_6323,N_5780,N_4224);
nand U6324 (N_6324,N_4303,N_5103);
nor U6325 (N_6325,N_5983,N_5367);
and U6326 (N_6326,N_4859,N_4350);
xnor U6327 (N_6327,N_4932,N_4393);
or U6328 (N_6328,N_4662,N_5952);
or U6329 (N_6329,N_4978,N_4903);
nand U6330 (N_6330,N_5375,N_5476);
or U6331 (N_6331,N_4103,N_5640);
or U6332 (N_6332,N_4468,N_5598);
or U6333 (N_6333,N_4595,N_4836);
and U6334 (N_6334,N_4300,N_4718);
nand U6335 (N_6335,N_5805,N_4893);
and U6336 (N_6336,N_5709,N_4346);
nand U6337 (N_6337,N_4090,N_4667);
nand U6338 (N_6338,N_5491,N_4097);
nand U6339 (N_6339,N_5564,N_4273);
and U6340 (N_6340,N_5116,N_4864);
nand U6341 (N_6341,N_4877,N_4835);
nand U6342 (N_6342,N_5469,N_5864);
and U6343 (N_6343,N_4308,N_5144);
nor U6344 (N_6344,N_5662,N_4229);
nand U6345 (N_6345,N_5731,N_5587);
xor U6346 (N_6346,N_5804,N_5389);
or U6347 (N_6347,N_5473,N_4412);
xor U6348 (N_6348,N_5810,N_4852);
or U6349 (N_6349,N_4917,N_5789);
nand U6350 (N_6350,N_5607,N_4539);
and U6351 (N_6351,N_4968,N_5714);
or U6352 (N_6352,N_5965,N_5725);
or U6353 (N_6353,N_4961,N_4230);
or U6354 (N_6354,N_5383,N_5009);
nor U6355 (N_6355,N_4882,N_4204);
nand U6356 (N_6356,N_4225,N_5666);
nor U6357 (N_6357,N_5606,N_4546);
and U6358 (N_6358,N_4009,N_5507);
nor U6359 (N_6359,N_5209,N_5485);
nor U6360 (N_6360,N_5412,N_5225);
or U6361 (N_6361,N_4658,N_4510);
and U6362 (N_6362,N_5149,N_5682);
and U6363 (N_6363,N_4935,N_4815);
or U6364 (N_6364,N_4331,N_5445);
nor U6365 (N_6365,N_5992,N_4989);
xnor U6366 (N_6366,N_5583,N_5345);
and U6367 (N_6367,N_4719,N_4421);
nand U6368 (N_6368,N_4562,N_4617);
nand U6369 (N_6369,N_4491,N_4288);
nor U6370 (N_6370,N_4950,N_4414);
and U6371 (N_6371,N_4275,N_5313);
or U6372 (N_6372,N_5287,N_5504);
and U6373 (N_6373,N_4660,N_5911);
and U6374 (N_6374,N_4768,N_4927);
and U6375 (N_6375,N_4721,N_5649);
nand U6376 (N_6376,N_5895,N_5304);
nor U6377 (N_6377,N_5596,N_5945);
and U6378 (N_6378,N_4068,N_4840);
or U6379 (N_6379,N_4247,N_5487);
nor U6380 (N_6380,N_4231,N_4058);
nand U6381 (N_6381,N_4138,N_4814);
or U6382 (N_6382,N_5415,N_4582);
xor U6383 (N_6383,N_4844,N_4613);
nor U6384 (N_6384,N_4969,N_4284);
nand U6385 (N_6385,N_4746,N_4044);
xor U6386 (N_6386,N_4831,N_4016);
nand U6387 (N_6387,N_5839,N_5944);
and U6388 (N_6388,N_4469,N_5732);
or U6389 (N_6389,N_4724,N_4198);
nor U6390 (N_6390,N_5297,N_4471);
nand U6391 (N_6391,N_5699,N_5826);
xnor U6392 (N_6392,N_5903,N_4756);
xnor U6393 (N_6393,N_5240,N_5066);
and U6394 (N_6394,N_5792,N_5845);
nor U6395 (N_6395,N_5070,N_5993);
or U6396 (N_6396,N_5602,N_5468);
or U6397 (N_6397,N_5852,N_4416);
xor U6398 (N_6398,N_5246,N_4286);
and U6399 (N_6399,N_5222,N_5080);
xnor U6400 (N_6400,N_5271,N_5749);
and U6401 (N_6401,N_4619,N_4880);
nor U6402 (N_6402,N_5806,N_5463);
or U6403 (N_6403,N_4990,N_4398);
nor U6404 (N_6404,N_5744,N_5405);
nand U6405 (N_6405,N_5901,N_5545);
and U6406 (N_6406,N_5654,N_5299);
and U6407 (N_6407,N_5368,N_5428);
or U6408 (N_6408,N_4236,N_4216);
nand U6409 (N_6409,N_4669,N_4738);
or U6410 (N_6410,N_4063,N_4736);
and U6411 (N_6411,N_5951,N_4701);
nand U6412 (N_6412,N_5787,N_5833);
nand U6413 (N_6413,N_4976,N_5621);
nand U6414 (N_6414,N_5761,N_5201);
or U6415 (N_6415,N_5790,N_4168);
xor U6416 (N_6416,N_4010,N_5626);
nand U6417 (N_6417,N_5553,N_5369);
nor U6418 (N_6418,N_5713,N_5819);
and U6419 (N_6419,N_4521,N_5526);
xnor U6420 (N_6420,N_4127,N_4640);
nor U6421 (N_6421,N_4997,N_4363);
xnor U6422 (N_6422,N_5704,N_4135);
and U6423 (N_6423,N_4661,N_5186);
nor U6424 (N_6424,N_4912,N_5461);
nor U6425 (N_6425,N_5782,N_5947);
nor U6426 (N_6426,N_5054,N_5489);
xnor U6427 (N_6427,N_4108,N_5677);
xnor U6428 (N_6428,N_5237,N_4645);
or U6429 (N_6429,N_4430,N_5435);
or U6430 (N_6430,N_5135,N_5453);
or U6431 (N_6431,N_4837,N_4076);
xor U6432 (N_6432,N_5733,N_5500);
xnor U6433 (N_6433,N_5550,N_4120);
nor U6434 (N_6434,N_4872,N_5492);
and U6435 (N_6435,N_4238,N_4342);
or U6436 (N_6436,N_4042,N_5972);
nor U6437 (N_6437,N_5770,N_4519);
or U6438 (N_6438,N_5348,N_4249);
or U6439 (N_6439,N_5264,N_5985);
nor U6440 (N_6440,N_5814,N_4344);
xor U6441 (N_6441,N_4349,N_5005);
nor U6442 (N_6442,N_5960,N_5466);
and U6443 (N_6443,N_5311,N_5734);
nand U6444 (N_6444,N_4488,N_4957);
xnor U6445 (N_6445,N_5063,N_5618);
nand U6446 (N_6446,N_4269,N_5976);
and U6447 (N_6447,N_4699,N_4581);
nand U6448 (N_6448,N_5086,N_4443);
and U6449 (N_6449,N_5322,N_5097);
nor U6450 (N_6450,N_4561,N_4325);
xor U6451 (N_6451,N_4312,N_5397);
nand U6452 (N_6452,N_4944,N_5853);
or U6453 (N_6453,N_4289,N_4253);
nor U6454 (N_6454,N_5527,N_4118);
nor U6455 (N_6455,N_4211,N_5717);
nor U6456 (N_6456,N_5343,N_5413);
xnor U6457 (N_6457,N_4079,N_4563);
and U6458 (N_6458,N_5002,N_5588);
xnor U6459 (N_6459,N_4175,N_5488);
xnor U6460 (N_6460,N_4396,N_5210);
nor U6461 (N_6461,N_5145,N_5471);
and U6462 (N_6462,N_5078,N_4462);
nor U6463 (N_6463,N_4557,N_5022);
nor U6464 (N_6464,N_5909,N_4757);
or U6465 (N_6465,N_5575,N_5031);
and U6466 (N_6466,N_5403,N_4427);
nor U6467 (N_6467,N_4082,N_4494);
nor U6468 (N_6468,N_4218,N_4888);
nand U6469 (N_6469,N_4955,N_5335);
and U6470 (N_6470,N_5846,N_4453);
nor U6471 (N_6471,N_4920,N_4898);
xor U6472 (N_6472,N_4516,N_4001);
nand U6473 (N_6473,N_4603,N_4205);
or U6474 (N_6474,N_4297,N_5619);
and U6475 (N_6475,N_5562,N_5268);
or U6476 (N_6476,N_4309,N_4140);
xor U6477 (N_6477,N_5090,N_4828);
or U6478 (N_6478,N_4863,N_5196);
xor U6479 (N_6479,N_4148,N_5534);
nor U6480 (N_6480,N_4217,N_5926);
nor U6481 (N_6481,N_4373,N_5844);
xnor U6482 (N_6482,N_4484,N_4070);
and U6483 (N_6483,N_4487,N_4005);
nand U6484 (N_6484,N_4600,N_5537);
and U6485 (N_6485,N_4979,N_4949);
nand U6486 (N_6486,N_4183,N_4345);
xor U6487 (N_6487,N_4858,N_5987);
or U6488 (N_6488,N_5524,N_4176);
nand U6489 (N_6489,N_5723,N_5498);
and U6490 (N_6490,N_4137,N_4274);
nand U6491 (N_6491,N_5130,N_5604);
nor U6492 (N_6492,N_4155,N_5935);
xor U6493 (N_6493,N_4507,N_5300);
xor U6494 (N_6494,N_5228,N_5884);
or U6495 (N_6495,N_4867,N_4276);
and U6496 (N_6496,N_4774,N_4759);
nor U6497 (N_6497,N_4348,N_4064);
nor U6498 (N_6498,N_5890,N_4607);
nand U6499 (N_6499,N_5840,N_5232);
nor U6500 (N_6500,N_5611,N_5673);
xnor U6501 (N_6501,N_5865,N_4534);
nand U6502 (N_6502,N_5726,N_4422);
nand U6503 (N_6503,N_5523,N_5419);
nand U6504 (N_6504,N_5110,N_4476);
nand U6505 (N_6505,N_5690,N_5994);
nor U6506 (N_6506,N_4834,N_5877);
xor U6507 (N_6507,N_4499,N_5778);
and U6508 (N_6508,N_4977,N_4861);
nor U6509 (N_6509,N_5483,N_5400);
xnor U6510 (N_6510,N_5641,N_4085);
nor U6511 (N_6511,N_4002,N_4048);
xor U6512 (N_6512,N_4784,N_5326);
and U6513 (N_6513,N_5691,N_4716);
xnor U6514 (N_6514,N_5341,N_4243);
or U6515 (N_6515,N_4733,N_4123);
or U6516 (N_6516,N_5908,N_4760);
nor U6517 (N_6517,N_4418,N_5949);
nor U6518 (N_6518,N_4672,N_4609);
and U6519 (N_6519,N_4382,N_4132);
nor U6520 (N_6520,N_4167,N_4052);
nand U6521 (N_6521,N_4096,N_5797);
nor U6522 (N_6522,N_4440,N_4615);
xor U6523 (N_6523,N_4405,N_5887);
nand U6524 (N_6524,N_4904,N_4650);
nor U6525 (N_6525,N_4178,N_4026);
nand U6526 (N_6526,N_5449,N_5594);
and U6527 (N_6527,N_4255,N_4299);
nand U6528 (N_6528,N_5114,N_5881);
and U6529 (N_6529,N_5610,N_5904);
nand U6530 (N_6530,N_4725,N_4452);
xnor U6531 (N_6531,N_4039,N_4388);
nand U6532 (N_6532,N_4921,N_4537);
and U6533 (N_6533,N_5065,N_5838);
and U6534 (N_6534,N_5220,N_4982);
or U6535 (N_6535,N_4165,N_5238);
nand U6536 (N_6536,N_4773,N_5517);
xor U6537 (N_6537,N_4663,N_5192);
xor U6538 (N_6538,N_4906,N_4729);
nor U6539 (N_6539,N_4735,N_4685);
xnor U6540 (N_6540,N_4441,N_5219);
nor U6541 (N_6541,N_5421,N_5800);
nand U6542 (N_6542,N_4813,N_5718);
xor U6543 (N_6543,N_4270,N_4188);
xnor U6544 (N_6544,N_4803,N_5458);
xnor U6545 (N_6545,N_5555,N_4072);
or U6546 (N_6546,N_4371,N_5202);
nand U6547 (N_6547,N_4381,N_5702);
xnor U6548 (N_6548,N_4092,N_5871);
and U6549 (N_6549,N_5076,N_5593);
xnor U6550 (N_6550,N_5679,N_4732);
nand U6551 (N_6551,N_4975,N_4226);
and U6552 (N_6552,N_4993,N_5885);
xnor U6553 (N_6553,N_5998,N_4873);
nand U6554 (N_6554,N_5950,N_4496);
nor U6555 (N_6555,N_5494,N_5685);
nor U6556 (N_6556,N_5170,N_5347);
and U6557 (N_6557,N_5392,N_5955);
nor U6558 (N_6558,N_4485,N_4161);
nor U6559 (N_6559,N_5316,N_5979);
xnor U6560 (N_6560,N_4856,N_4956);
nor U6561 (N_6561,N_4486,N_4652);
and U6562 (N_6562,N_5180,N_5591);
xor U6563 (N_6563,N_4240,N_5779);
nor U6564 (N_6564,N_4187,N_4745);
xor U6565 (N_6565,N_4268,N_5391);
nand U6566 (N_6566,N_5291,N_5148);
nor U6567 (N_6567,N_5099,N_5361);
or U6568 (N_6568,N_4531,N_5700);
or U6569 (N_6569,N_4306,N_5784);
or U6570 (N_6570,N_5156,N_5191);
or U6571 (N_6571,N_5817,N_5763);
and U6572 (N_6572,N_5139,N_5747);
xnor U6573 (N_6573,N_4180,N_4190);
and U6574 (N_6574,N_5659,N_4824);
and U6575 (N_6575,N_5309,N_5200);
nand U6576 (N_6576,N_5705,N_4354);
xnor U6577 (N_6577,N_4634,N_5162);
nand U6578 (N_6578,N_4692,N_4754);
or U6579 (N_6579,N_5879,N_4456);
and U6580 (N_6580,N_4513,N_5357);
or U6581 (N_6581,N_5224,N_5046);
xnor U6582 (N_6582,N_5378,N_5622);
xor U6583 (N_6583,N_4845,N_5284);
nor U6584 (N_6584,N_4338,N_5317);
xor U6585 (N_6585,N_4201,N_5891);
or U6586 (N_6586,N_5758,N_5095);
xnor U6587 (N_6587,N_4657,N_5582);
xor U6588 (N_6588,N_5793,N_4632);
nor U6589 (N_6589,N_5364,N_4439);
nor U6590 (N_6590,N_4758,N_5547);
nand U6591 (N_6591,N_4366,N_5432);
nor U6592 (N_6592,N_5762,N_5125);
and U6593 (N_6593,N_5910,N_4200);
nand U6594 (N_6594,N_5429,N_5451);
xor U6595 (N_6595,N_5646,N_4584);
nand U6596 (N_6596,N_5179,N_4057);
xnor U6597 (N_6597,N_4133,N_5918);
nor U6598 (N_6598,N_4015,N_4514);
xnor U6599 (N_6599,N_5073,N_4807);
nor U6600 (N_6600,N_4847,N_5106);
nor U6601 (N_6601,N_5533,N_5964);
or U6602 (N_6602,N_5905,N_5765);
or U6603 (N_6603,N_4166,N_5253);
nand U6604 (N_6604,N_5124,N_4094);
xnor U6605 (N_6605,N_4088,N_4536);
and U6606 (N_6606,N_5048,N_5989);
nor U6607 (N_6607,N_5182,N_5638);
or U6608 (N_6608,N_4307,N_4564);
nand U6609 (N_6609,N_5021,N_5566);
xor U6610 (N_6610,N_5330,N_5505);
nor U6611 (N_6611,N_5856,N_4252);
nor U6612 (N_6612,N_4206,N_4527);
or U6613 (N_6613,N_5757,N_5025);
or U6614 (N_6614,N_4551,N_5414);
xor U6615 (N_6615,N_5223,N_5832);
nand U6616 (N_6616,N_4543,N_4651);
nor U6617 (N_6617,N_5101,N_4355);
nand U6618 (N_6618,N_5600,N_4489);
and U6619 (N_6619,N_5661,N_5017);
nand U6620 (N_6620,N_4789,N_5906);
xnor U6621 (N_6621,N_4734,N_5321);
nor U6622 (N_6622,N_4220,N_5052);
nor U6623 (N_6623,N_4710,N_5629);
and U6624 (N_6624,N_5198,N_5874);
xor U6625 (N_6625,N_5999,N_5648);
xor U6626 (N_6626,N_5934,N_5259);
nand U6627 (N_6627,N_4923,N_5539);
and U6628 (N_6628,N_4313,N_5217);
nor U6629 (N_6629,N_4235,N_4472);
nand U6630 (N_6630,N_5922,N_5689);
nor U6631 (N_6631,N_4533,N_4333);
nand U6632 (N_6632,N_4832,N_4040);
or U6633 (N_6633,N_5153,N_5100);
and U6634 (N_6634,N_4780,N_4630);
xnor U6635 (N_6635,N_4848,N_4753);
nand U6636 (N_6636,N_4056,N_5410);
and U6637 (N_6637,N_4383,N_4884);
xnor U6638 (N_6638,N_5737,N_5129);
nand U6639 (N_6639,N_4542,N_4796);
and U6640 (N_6640,N_4585,N_4708);
and U6641 (N_6641,N_4599,N_4916);
nor U6642 (N_6642,N_4540,N_4461);
xor U6643 (N_6643,N_5168,N_4573);
and U6644 (N_6644,N_5136,N_5175);
nand U6645 (N_6645,N_5047,N_4928);
and U6646 (N_6646,N_4908,N_5298);
nor U6647 (N_6647,N_5697,N_5796);
and U6648 (N_6648,N_5862,N_5692);
xor U6649 (N_6649,N_4380,N_5863);
or U6650 (N_6650,N_5014,N_4077);
and U6651 (N_6651,N_4199,N_5279);
nand U6652 (N_6652,N_5377,N_5442);
and U6653 (N_6653,N_4172,N_5111);
and U6654 (N_6654,N_4740,N_5275);
or U6655 (N_6655,N_5373,N_5809);
and U6656 (N_6656,N_5189,N_5984);
and U6657 (N_6657,N_4285,N_4918);
xnor U6658 (N_6658,N_5821,N_4394);
and U6659 (N_6659,N_4890,N_5351);
xor U6660 (N_6660,N_5754,N_5857);
and U6661 (N_6661,N_5799,N_4723);
or U6662 (N_6662,N_5506,N_5921);
nor U6663 (N_6663,N_5569,N_5695);
or U6664 (N_6664,N_4816,N_4203);
or U6665 (N_6665,N_5837,N_5024);
nor U6666 (N_6666,N_4237,N_4971);
nand U6667 (N_6667,N_5535,N_4707);
and U6668 (N_6668,N_5454,N_5755);
and U6669 (N_6669,N_5785,N_4970);
xnor U6670 (N_6670,N_5012,N_5546);
or U6671 (N_6671,N_5006,N_5831);
nor U6672 (N_6672,N_4511,N_4332);
and U6673 (N_6673,N_4464,N_4889);
xor U6674 (N_6674,N_4359,N_4340);
nor U6675 (N_6675,N_5475,N_5053);
or U6676 (N_6676,N_5882,N_4117);
and U6677 (N_6677,N_5331,N_4688);
or U6678 (N_6678,N_4709,N_4905);
or U6679 (N_6679,N_4392,N_5060);
or U6680 (N_6680,N_5720,N_5140);
nand U6681 (N_6681,N_5614,N_4593);
xor U6682 (N_6682,N_5642,N_4214);
nand U6683 (N_6683,N_4047,N_5727);
or U6684 (N_6684,N_4576,N_4665);
xor U6685 (N_6685,N_4874,N_4690);
or U6686 (N_6686,N_4185,N_4157);
and U6687 (N_6687,N_4987,N_4162);
nand U6688 (N_6688,N_4257,N_5674);
xnor U6689 (N_6689,N_5193,N_5590);
or U6690 (N_6690,N_5423,N_4554);
nand U6691 (N_6691,N_4319,N_4480);
xnor U6692 (N_6692,N_4579,N_5307);
and U6693 (N_6693,N_5501,N_4159);
nand U6694 (N_6694,N_5165,N_5286);
nor U6695 (N_6695,N_5015,N_4914);
nand U6696 (N_6696,N_5924,N_5242);
nand U6697 (N_6697,N_4377,N_5643);
or U6698 (N_6698,N_5427,N_5828);
nor U6699 (N_6699,N_5243,N_4445);
or U6700 (N_6700,N_4212,N_5665);
and U6701 (N_6701,N_5178,N_4391);
nor U6702 (N_6702,N_4404,N_4143);
and U6703 (N_6703,N_4683,N_5324);
xor U6704 (N_6704,N_4153,N_5312);
and U6705 (N_6705,N_5447,N_4419);
xor U6706 (N_6706,N_4952,N_4098);
nand U6707 (N_6707,N_4171,N_4227);
and U6708 (N_6708,N_5858,N_5115);
or U6709 (N_6709,N_5605,N_5134);
nor U6710 (N_6710,N_4101,N_5511);
nor U6711 (N_6711,N_4656,N_5055);
or U6712 (N_6712,N_5825,N_5769);
or U6713 (N_6713,N_5764,N_4055);
and U6714 (N_6714,N_5996,N_5061);
nor U6715 (N_6715,N_5226,N_5227);
nor U6716 (N_6716,N_5639,N_5615);
nor U6717 (N_6717,N_5743,N_5230);
or U6718 (N_6718,N_4938,N_4365);
nand U6719 (N_6719,N_4173,N_4352);
or U6720 (N_6720,N_5668,N_5556);
nor U6721 (N_6721,N_5777,N_5315);
and U6722 (N_6722,N_4726,N_4156);
nor U6723 (N_6723,N_4362,N_5499);
nor U6724 (N_6724,N_5532,N_5365);
xor U6725 (N_6725,N_4330,N_4610);
nor U6726 (N_6726,N_5072,N_4036);
nand U6727 (N_6727,N_5457,N_4895);
nor U6728 (N_6728,N_5916,N_5029);
xor U6729 (N_6729,N_4702,N_5233);
nor U6730 (N_6730,N_5822,N_5554);
or U6731 (N_6731,N_4281,N_4311);
xnor U6732 (N_6732,N_4625,N_4624);
and U6733 (N_6733,N_5374,N_4147);
xnor U6734 (N_6734,N_4596,N_4470);
xnor U6735 (N_6735,N_4810,N_4767);
nor U6736 (N_6736,N_5724,N_5599);
or U6737 (N_6737,N_5430,N_5155);
or U6738 (N_6738,N_4403,N_4620);
xor U6739 (N_6739,N_4588,N_5289);
or U6740 (N_6740,N_5199,N_5670);
xnor U6741 (N_6741,N_4011,N_5835);
nand U6742 (N_6742,N_5058,N_4808);
nand U6743 (N_6743,N_5045,N_4141);
and U6744 (N_6744,N_5842,N_5751);
nor U6745 (N_6745,N_4532,N_5721);
nor U6746 (N_6746,N_5735,N_4675);
xor U6747 (N_6747,N_4518,N_5188);
nand U6748 (N_6748,N_4846,N_4290);
nand U6749 (N_6749,N_5956,N_5902);
nand U6750 (N_6750,N_4020,N_4686);
nor U6751 (N_6751,N_4597,N_5969);
and U6752 (N_6752,N_5265,N_4963);
nand U6753 (N_6753,N_5157,N_4425);
or U6754 (N_6754,N_5169,N_5133);
and U6755 (N_6755,N_4457,N_4483);
or U6756 (N_6756,N_5172,N_5722);
xnor U6757 (N_6757,N_5203,N_5795);
xnor U6758 (N_6758,N_5719,N_4705);
nor U6759 (N_6759,N_4397,N_5869);
nand U6760 (N_6760,N_5930,N_5586);
nand U6761 (N_6761,N_4951,N_4628);
and U6762 (N_6762,N_4958,N_5574);
xor U6763 (N_6763,N_4887,N_4062);
nand U6764 (N_6764,N_5404,N_4878);
and U6765 (N_6765,N_5408,N_5318);
nor U6766 (N_6766,N_4444,N_5543);
nor U6767 (N_6767,N_5929,N_4798);
nor U6768 (N_6768,N_4787,N_4988);
or U6769 (N_6769,N_5132,N_4822);
and U6770 (N_6770,N_5218,N_5229);
and U6771 (N_6771,N_5422,N_5548);
or U6772 (N_6772,N_4842,N_5516);
nand U6773 (N_6773,N_5482,N_5678);
or U6774 (N_6774,N_5085,N_4046);
and U6775 (N_6775,N_5803,N_5372);
or U6776 (N_6776,N_4763,N_5536);
and U6777 (N_6777,N_5808,N_4111);
nor U6778 (N_6778,N_5087,N_4008);
nor U6779 (N_6779,N_4567,N_5493);
nand U6780 (N_6780,N_5096,N_5850);
nor U6781 (N_6781,N_5062,N_4752);
and U6782 (N_6782,N_4442,N_5514);
nand U6783 (N_6783,N_4460,N_5883);
or U6784 (N_6784,N_4764,N_5914);
and U6785 (N_6785,N_5937,N_5812);
or U6786 (N_6786,N_4434,N_4776);
or U6787 (N_6787,N_5597,N_5122);
nor U6788 (N_6788,N_5570,N_5919);
or U6789 (N_6789,N_5036,N_5239);
or U6790 (N_6790,N_5893,N_4841);
nand U6791 (N_6791,N_5696,N_4857);
nor U6792 (N_6792,N_4125,N_5448);
nand U6793 (N_6793,N_4305,N_4018);
and U6794 (N_6794,N_4102,N_5004);
and U6795 (N_6795,N_5147,N_5581);
or U6796 (N_6796,N_5768,N_5627);
nor U6797 (N_6797,N_4431,N_4565);
nand U6798 (N_6798,N_4293,N_5280);
xnor U6799 (N_6799,N_5707,N_4644);
or U6800 (N_6800,N_5260,N_4783);
and U6801 (N_6801,N_4637,N_5860);
xor U6802 (N_6802,N_5293,N_4478);
nor U6803 (N_6803,N_5920,N_4482);
or U6804 (N_6804,N_5371,N_5592);
or U6805 (N_6805,N_5813,N_5818);
nor U6806 (N_6806,N_5050,N_5251);
xor U6807 (N_6807,N_5285,N_4849);
nand U6808 (N_6808,N_5503,N_5559);
nor U6809 (N_6809,N_5687,N_4196);
and U6810 (N_6810,N_4322,N_5038);
xor U6811 (N_6811,N_5438,N_4910);
nor U6812 (N_6812,N_4682,N_5847);
or U6813 (N_6813,N_4248,N_4407);
xnor U6814 (N_6814,N_5310,N_4449);
nand U6815 (N_6815,N_4942,N_4730);
nand U6816 (N_6816,N_5510,N_5579);
nor U6817 (N_6817,N_5319,N_5039);
nor U6818 (N_6818,N_5323,N_4695);
nor U6819 (N_6819,N_4883,N_4896);
or U6820 (N_6820,N_5849,N_4207);
nand U6821 (N_6821,N_5113,N_4221);
nor U6822 (N_6822,N_4552,N_5774);
or U6823 (N_6823,N_5636,N_4025);
xnor U6824 (N_6824,N_4051,N_4558);
nand U6825 (N_6825,N_4061,N_4222);
xnor U6826 (N_6826,N_5896,N_4929);
nand U6827 (N_6827,N_5327,N_5990);
or U6828 (N_6828,N_5484,N_5402);
xor U6829 (N_6829,N_4409,N_4119);
nand U6830 (N_6830,N_4947,N_5470);
xor U6831 (N_6831,N_5939,N_4671);
nor U6832 (N_6832,N_5146,N_5450);
nor U6833 (N_6833,N_4139,N_5387);
and U6834 (N_6834,N_4465,N_4525);
nor U6835 (N_6835,N_4892,N_5384);
and U6836 (N_6836,N_4679,N_4256);
and U6837 (N_6837,N_5128,N_5834);
nand U6838 (N_6838,N_4739,N_5997);
nor U6839 (N_6839,N_4555,N_4219);
xnor U6840 (N_6840,N_5609,N_4966);
nor U6841 (N_6841,N_5759,N_4295);
or U6842 (N_6842,N_4691,N_4066);
and U6843 (N_6843,N_4924,N_4995);
nor U6844 (N_6844,N_5043,N_4179);
nand U6845 (N_6845,N_4477,N_5394);
nor U6846 (N_6846,N_5970,N_4000);
and U6847 (N_6847,N_4526,N_5577);
xnor U6848 (N_6848,N_4324,N_5486);
xnor U6849 (N_6849,N_5549,N_4209);
nand U6850 (N_6850,N_5478,N_4616);
or U6851 (N_6851,N_5292,N_5655);
nor U6852 (N_6852,N_5978,N_4232);
or U6853 (N_6853,N_5651,N_5352);
nand U6854 (N_6854,N_5518,N_4417);
xnor U6855 (N_6855,N_4242,N_4501);
and U6856 (N_6856,N_4263,N_5623);
or U6857 (N_6857,N_5540,N_4765);
nand U6858 (N_6858,N_5973,N_4326);
and U6859 (N_6859,N_4505,N_5520);
nand U6860 (N_6860,N_4587,N_4670);
or U6861 (N_6861,N_5344,N_4481);
xnor U6862 (N_6862,N_5441,N_4522);
nand U6863 (N_6863,N_4830,N_5354);
or U6864 (N_6864,N_4113,N_5986);
xor U6865 (N_6865,N_5211,N_5565);
and U6866 (N_6866,N_5672,N_4078);
or U6867 (N_6867,N_5030,N_5962);
nor U6868 (N_6868,N_4876,N_4192);
or U6869 (N_6869,N_4033,N_4805);
nor U6870 (N_6870,N_4023,N_4164);
and U6871 (N_6871,N_4149,N_5811);
xor U6872 (N_6872,N_5183,N_5181);
nand U6873 (N_6873,N_4794,N_4030);
xor U6874 (N_6874,N_4827,N_5912);
nor U6875 (N_6875,N_4109,N_5411);
nand U6876 (N_6876,N_4761,N_5137);
xnor U6877 (N_6877,N_5900,N_5558);
and U6878 (N_6878,N_5966,N_5084);
nor U6879 (N_6879,N_5899,N_5959);
or U6880 (N_6880,N_4618,N_5563);
nand U6881 (N_6881,N_5437,N_4871);
or U6882 (N_6882,N_5044,N_4806);
nor U6883 (N_6883,N_5328,N_4911);
and U6884 (N_6884,N_4939,N_4770);
and U6885 (N_6885,N_4983,N_5961);
xor U6886 (N_6886,N_4426,N_5407);
nor U6887 (N_6887,N_5519,N_4680);
and U6888 (N_6888,N_4054,N_5750);
xnor U6889 (N_6889,N_5079,N_5018);
or U6890 (N_6890,N_4788,N_5255);
or U6891 (N_6891,N_4075,N_4347);
and U6892 (N_6892,N_4795,N_5208);
or U6893 (N_6893,N_4771,N_5771);
xor U6894 (N_6894,N_5221,N_4357);
or U6895 (N_6895,N_5164,N_5359);
nand U6896 (N_6896,N_4087,N_5386);
and U6897 (N_6897,N_4007,N_4791);
nand U6898 (N_6898,N_5353,N_5490);
or U6899 (N_6899,N_5174,N_4647);
or U6900 (N_6900,N_4664,N_5684);
or U6901 (N_6901,N_4035,N_4329);
xnor U6902 (N_6902,N_4099,N_4943);
nand U6903 (N_6903,N_5783,N_4433);
or U6904 (N_6904,N_4623,N_5075);
nand U6905 (N_6905,N_5560,N_4570);
nand U6906 (N_6906,N_4594,N_4073);
or U6907 (N_6907,N_4627,N_4186);
nand U6908 (N_6908,N_4241,N_5390);
xor U6909 (N_6909,N_5830,N_4423);
or U6910 (N_6910,N_5898,N_4495);
nor U6911 (N_6911,N_4894,N_5634);
nor U6912 (N_6912,N_4635,N_4316);
and U6913 (N_6913,N_4463,N_4741);
or U6914 (N_6914,N_5346,N_5876);
or U6915 (N_6915,N_4602,N_5927);
nand U6916 (N_6916,N_4706,N_5398);
and U6917 (N_6917,N_4115,N_5495);
nor U6918 (N_6918,N_4547,N_4479);
xor U6919 (N_6919,N_4174,N_4012);
xnor U6920 (N_6920,N_5741,N_5118);
nand U6921 (N_6921,N_4428,N_4778);
xor U6922 (N_6922,N_4170,N_5843);
nand U6923 (N_6923,N_5439,N_4601);
xor U6924 (N_6924,N_5214,N_5105);
xnor U6925 (N_6925,N_4720,N_5460);
or U6926 (N_6926,N_5382,N_4146);
nand U6927 (N_6927,N_5889,N_5302);
nand U6928 (N_6928,N_4568,N_5109);
and U6929 (N_6929,N_4545,N_5716);
xor U6930 (N_6930,N_4353,N_5399);
nand U6931 (N_6931,N_4717,N_5204);
nand U6932 (N_6932,N_4654,N_4283);
xnor U6933 (N_6933,N_5848,N_4083);
nand U6934 (N_6934,N_5738,N_5092);
and U6935 (N_6935,N_5277,N_4372);
nor U6936 (N_6936,N_4954,N_4902);
and U6937 (N_6937,N_5971,N_4550);
and U6938 (N_6938,N_5173,N_5766);
and U6939 (N_6939,N_4713,N_5190);
nor U6940 (N_6940,N_5669,N_4926);
nor U6941 (N_6941,N_5288,N_4459);
xor U6942 (N_6942,N_4901,N_4696);
and U6943 (N_6943,N_5617,N_5509);
xor U6944 (N_6944,N_4714,N_4743);
xor U6945 (N_6945,N_5154,N_4821);
and U6946 (N_6946,N_5334,N_5000);
and U6947 (N_6947,N_4262,N_4436);
or U6948 (N_6948,N_5088,N_5333);
xnor U6949 (N_6949,N_4112,N_4402);
nand U6950 (N_6950,N_4038,N_4687);
xnor U6951 (N_6951,N_4454,N_5093);
and U6952 (N_6952,N_4818,N_5886);
xnor U6953 (N_6953,N_4591,N_5544);
nand U6954 (N_6954,N_5528,N_4356);
and U6955 (N_6955,N_4335,N_4341);
or U6956 (N_6956,N_4210,N_5968);
and U6957 (N_6957,N_4323,N_4095);
nand U6958 (N_6958,N_5308,N_4379);
xor U6959 (N_6959,N_4681,N_4282);
xor U6960 (N_6960,N_5663,N_4801);
nor U6961 (N_6961,N_5089,N_5380);
or U6962 (N_6962,N_4985,N_4110);
xnor U6963 (N_6963,N_4972,N_5928);
nor U6964 (N_6964,N_5160,N_5647);
or U6965 (N_6965,N_4160,N_4860);
nor U6966 (N_6966,N_5064,N_4934);
nor U6967 (N_6967,N_5740,N_4992);
or U6968 (N_6968,N_5120,N_4208);
nor U6969 (N_6969,N_4855,N_4960);
or U6970 (N_6970,N_5363,N_4535);
or U6971 (N_6971,N_4385,N_5273);
xor U6972 (N_6972,N_4715,N_4037);
and U6973 (N_6973,N_5957,N_5395);
xnor U6974 (N_6974,N_4466,N_5995);
or U6975 (N_6975,N_5530,N_4406);
or U6976 (N_6976,N_4933,N_5552);
and U6977 (N_6977,N_5358,N_5632);
or U6978 (N_6978,N_5446,N_5069);
and U6979 (N_6979,N_5067,N_5459);
nand U6980 (N_6980,N_4529,N_4069);
nor U6981 (N_6981,N_4328,N_5042);
xnor U6982 (N_6982,N_4891,N_4502);
or U6983 (N_6983,N_5008,N_5515);
and U6984 (N_6984,N_5942,N_4812);
or U6985 (N_6985,N_4251,N_4823);
and U6986 (N_6986,N_4151,N_5256);
or U6987 (N_6987,N_5752,N_4059);
nor U6988 (N_6988,N_4586,N_5418);
and U6989 (N_6989,N_5329,N_5205);
or U6990 (N_6990,N_4953,N_4246);
nor U6991 (N_6991,N_5568,N_4973);
nand U6992 (N_6992,N_5729,N_4598);
nand U6993 (N_6993,N_5416,N_4136);
xnor U6994 (N_6994,N_5773,N_4296);
and U6995 (N_6995,N_4790,N_5931);
nand U6996 (N_6996,N_5943,N_4751);
nor U6997 (N_6997,N_4744,N_4553);
or U6998 (N_6998,N_4621,N_4154);
and U6999 (N_6999,N_4577,N_5194);
nor U7000 (N_7000,N_5849,N_4702);
nand U7001 (N_7001,N_4635,N_5335);
xor U7002 (N_7002,N_4773,N_4839);
and U7003 (N_7003,N_4612,N_4090);
xor U7004 (N_7004,N_4331,N_4066);
xnor U7005 (N_7005,N_5523,N_5454);
or U7006 (N_7006,N_5744,N_4930);
nor U7007 (N_7007,N_5265,N_4263);
nand U7008 (N_7008,N_4633,N_4699);
xor U7009 (N_7009,N_4453,N_4393);
xnor U7010 (N_7010,N_4461,N_5308);
nand U7011 (N_7011,N_4635,N_5234);
or U7012 (N_7012,N_5499,N_4732);
and U7013 (N_7013,N_5454,N_5033);
and U7014 (N_7014,N_5192,N_5574);
or U7015 (N_7015,N_4588,N_5010);
or U7016 (N_7016,N_5623,N_4656);
xor U7017 (N_7017,N_5202,N_5217);
xnor U7018 (N_7018,N_4647,N_5939);
and U7019 (N_7019,N_5406,N_5282);
nand U7020 (N_7020,N_5674,N_4611);
nand U7021 (N_7021,N_4359,N_4354);
xnor U7022 (N_7022,N_5389,N_5019);
and U7023 (N_7023,N_4062,N_4727);
and U7024 (N_7024,N_5090,N_5443);
nor U7025 (N_7025,N_5746,N_4284);
nand U7026 (N_7026,N_5250,N_5779);
xnor U7027 (N_7027,N_4054,N_5290);
and U7028 (N_7028,N_5167,N_5467);
nand U7029 (N_7029,N_4093,N_4242);
nor U7030 (N_7030,N_5656,N_4426);
or U7031 (N_7031,N_4326,N_4421);
nor U7032 (N_7032,N_4142,N_4323);
nor U7033 (N_7033,N_5961,N_4357);
nand U7034 (N_7034,N_4808,N_4290);
nor U7035 (N_7035,N_4014,N_5133);
xnor U7036 (N_7036,N_5789,N_4154);
nor U7037 (N_7037,N_4545,N_5067);
and U7038 (N_7038,N_5465,N_4451);
or U7039 (N_7039,N_4471,N_5745);
and U7040 (N_7040,N_4280,N_4818);
xor U7041 (N_7041,N_4130,N_5699);
nor U7042 (N_7042,N_5424,N_5675);
nand U7043 (N_7043,N_4549,N_4419);
and U7044 (N_7044,N_4590,N_4426);
nor U7045 (N_7045,N_5409,N_5791);
nor U7046 (N_7046,N_5290,N_5509);
xor U7047 (N_7047,N_5849,N_5489);
and U7048 (N_7048,N_5718,N_4417);
nor U7049 (N_7049,N_4987,N_5650);
nand U7050 (N_7050,N_5658,N_5776);
xor U7051 (N_7051,N_4065,N_4684);
nand U7052 (N_7052,N_4638,N_4662);
and U7053 (N_7053,N_4363,N_5994);
nand U7054 (N_7054,N_4561,N_5291);
and U7055 (N_7055,N_4417,N_5845);
nand U7056 (N_7056,N_5344,N_4958);
or U7057 (N_7057,N_5556,N_5831);
or U7058 (N_7058,N_5666,N_4203);
nor U7059 (N_7059,N_5068,N_5143);
or U7060 (N_7060,N_4566,N_5225);
or U7061 (N_7061,N_5897,N_4485);
nand U7062 (N_7062,N_5537,N_5175);
xnor U7063 (N_7063,N_5593,N_5416);
xnor U7064 (N_7064,N_4793,N_5581);
and U7065 (N_7065,N_4934,N_5451);
nand U7066 (N_7066,N_4987,N_5883);
and U7067 (N_7067,N_5435,N_5342);
nand U7068 (N_7068,N_4422,N_4721);
and U7069 (N_7069,N_4604,N_4524);
nand U7070 (N_7070,N_4173,N_5383);
xnor U7071 (N_7071,N_4712,N_4540);
and U7072 (N_7072,N_4567,N_5046);
nand U7073 (N_7073,N_4706,N_4806);
xor U7074 (N_7074,N_4078,N_4981);
xnor U7075 (N_7075,N_5153,N_5469);
and U7076 (N_7076,N_5816,N_5087);
nor U7077 (N_7077,N_5275,N_4362);
or U7078 (N_7078,N_5390,N_4586);
nor U7079 (N_7079,N_4852,N_4444);
xor U7080 (N_7080,N_5869,N_5520);
xor U7081 (N_7081,N_4327,N_4757);
xor U7082 (N_7082,N_5153,N_4813);
or U7083 (N_7083,N_4034,N_4825);
and U7084 (N_7084,N_4035,N_4217);
nor U7085 (N_7085,N_4823,N_4640);
and U7086 (N_7086,N_4364,N_5517);
or U7087 (N_7087,N_5122,N_5747);
and U7088 (N_7088,N_4202,N_4660);
and U7089 (N_7089,N_4095,N_4437);
nand U7090 (N_7090,N_5747,N_5724);
or U7091 (N_7091,N_4879,N_5672);
nor U7092 (N_7092,N_5723,N_4859);
nand U7093 (N_7093,N_5391,N_5088);
nand U7094 (N_7094,N_4357,N_5908);
nor U7095 (N_7095,N_4224,N_5371);
and U7096 (N_7096,N_5467,N_5042);
or U7097 (N_7097,N_4719,N_5309);
or U7098 (N_7098,N_5814,N_5502);
nor U7099 (N_7099,N_4012,N_5567);
nor U7100 (N_7100,N_4201,N_5895);
or U7101 (N_7101,N_4357,N_5991);
nand U7102 (N_7102,N_4587,N_5593);
xnor U7103 (N_7103,N_4598,N_4939);
xnor U7104 (N_7104,N_5089,N_5360);
nand U7105 (N_7105,N_4081,N_4629);
xnor U7106 (N_7106,N_5971,N_5809);
nand U7107 (N_7107,N_4506,N_5355);
or U7108 (N_7108,N_4274,N_5010);
xor U7109 (N_7109,N_5503,N_4068);
xor U7110 (N_7110,N_4193,N_5451);
xnor U7111 (N_7111,N_5544,N_5475);
and U7112 (N_7112,N_5050,N_5029);
xor U7113 (N_7113,N_5575,N_4931);
xnor U7114 (N_7114,N_4099,N_5499);
and U7115 (N_7115,N_4518,N_5763);
or U7116 (N_7116,N_4015,N_4201);
nor U7117 (N_7117,N_4887,N_5242);
xor U7118 (N_7118,N_5632,N_4256);
and U7119 (N_7119,N_4821,N_5008);
nand U7120 (N_7120,N_4686,N_5879);
nor U7121 (N_7121,N_5940,N_4149);
and U7122 (N_7122,N_5647,N_4408);
nand U7123 (N_7123,N_4160,N_4482);
or U7124 (N_7124,N_5550,N_4734);
nand U7125 (N_7125,N_5120,N_4944);
nor U7126 (N_7126,N_5984,N_5623);
xnor U7127 (N_7127,N_5251,N_5456);
nand U7128 (N_7128,N_4729,N_5025);
and U7129 (N_7129,N_5681,N_5017);
and U7130 (N_7130,N_4986,N_4426);
xnor U7131 (N_7131,N_4441,N_5603);
and U7132 (N_7132,N_4225,N_4676);
nor U7133 (N_7133,N_5461,N_4590);
xor U7134 (N_7134,N_5273,N_5026);
nor U7135 (N_7135,N_5549,N_5290);
nand U7136 (N_7136,N_4470,N_4864);
nand U7137 (N_7137,N_4864,N_4878);
and U7138 (N_7138,N_5666,N_5728);
nand U7139 (N_7139,N_5216,N_5915);
and U7140 (N_7140,N_4376,N_4804);
or U7141 (N_7141,N_5873,N_5815);
nor U7142 (N_7142,N_5618,N_5513);
or U7143 (N_7143,N_5871,N_5091);
nand U7144 (N_7144,N_5100,N_5283);
nor U7145 (N_7145,N_5722,N_5016);
xnor U7146 (N_7146,N_5964,N_4776);
nor U7147 (N_7147,N_4819,N_5220);
or U7148 (N_7148,N_4473,N_4417);
xnor U7149 (N_7149,N_4604,N_5043);
or U7150 (N_7150,N_5278,N_4252);
nand U7151 (N_7151,N_4938,N_4450);
xnor U7152 (N_7152,N_5612,N_5554);
nor U7153 (N_7153,N_4314,N_4098);
xor U7154 (N_7154,N_5551,N_5016);
or U7155 (N_7155,N_5493,N_4032);
and U7156 (N_7156,N_5010,N_5705);
xnor U7157 (N_7157,N_4577,N_5829);
nand U7158 (N_7158,N_4096,N_4458);
nand U7159 (N_7159,N_5096,N_4085);
nor U7160 (N_7160,N_4948,N_4251);
xnor U7161 (N_7161,N_4793,N_5466);
nand U7162 (N_7162,N_5817,N_4006);
or U7163 (N_7163,N_5772,N_5187);
or U7164 (N_7164,N_5258,N_4721);
xor U7165 (N_7165,N_5636,N_4964);
nand U7166 (N_7166,N_4585,N_5581);
or U7167 (N_7167,N_5610,N_5037);
nand U7168 (N_7168,N_5756,N_5599);
or U7169 (N_7169,N_5662,N_5159);
or U7170 (N_7170,N_4624,N_4059);
xnor U7171 (N_7171,N_4663,N_4893);
nor U7172 (N_7172,N_5504,N_5330);
and U7173 (N_7173,N_5069,N_5077);
or U7174 (N_7174,N_5893,N_4247);
nor U7175 (N_7175,N_4317,N_4493);
nand U7176 (N_7176,N_4220,N_4785);
nor U7177 (N_7177,N_5407,N_5658);
xor U7178 (N_7178,N_4109,N_5834);
nor U7179 (N_7179,N_5244,N_5050);
or U7180 (N_7180,N_4358,N_5178);
xor U7181 (N_7181,N_4431,N_4911);
and U7182 (N_7182,N_4864,N_5420);
or U7183 (N_7183,N_4744,N_4268);
xor U7184 (N_7184,N_4604,N_4155);
xor U7185 (N_7185,N_4917,N_4363);
or U7186 (N_7186,N_5759,N_5974);
nand U7187 (N_7187,N_4621,N_4547);
xor U7188 (N_7188,N_4627,N_4368);
or U7189 (N_7189,N_4593,N_4577);
and U7190 (N_7190,N_5954,N_4674);
nor U7191 (N_7191,N_5807,N_4437);
xor U7192 (N_7192,N_5840,N_4246);
xnor U7193 (N_7193,N_5751,N_4225);
xnor U7194 (N_7194,N_4682,N_4502);
nand U7195 (N_7195,N_4973,N_4358);
nor U7196 (N_7196,N_4709,N_4093);
xnor U7197 (N_7197,N_4221,N_4585);
or U7198 (N_7198,N_5011,N_4427);
nor U7199 (N_7199,N_5644,N_5127);
nand U7200 (N_7200,N_5490,N_5470);
xor U7201 (N_7201,N_4268,N_4544);
or U7202 (N_7202,N_5569,N_5308);
nand U7203 (N_7203,N_4095,N_4500);
nor U7204 (N_7204,N_4044,N_4083);
xor U7205 (N_7205,N_5439,N_4325);
or U7206 (N_7206,N_4183,N_4870);
xnor U7207 (N_7207,N_5338,N_5319);
and U7208 (N_7208,N_4990,N_4537);
nor U7209 (N_7209,N_5046,N_5643);
xnor U7210 (N_7210,N_5754,N_5482);
nor U7211 (N_7211,N_5878,N_5084);
xor U7212 (N_7212,N_4208,N_4109);
xnor U7213 (N_7213,N_4428,N_4849);
or U7214 (N_7214,N_5670,N_5802);
and U7215 (N_7215,N_5286,N_5785);
xnor U7216 (N_7216,N_4336,N_4361);
nor U7217 (N_7217,N_4522,N_5426);
or U7218 (N_7218,N_5716,N_5294);
nand U7219 (N_7219,N_4453,N_4396);
and U7220 (N_7220,N_5180,N_4261);
and U7221 (N_7221,N_5275,N_5220);
xor U7222 (N_7222,N_5344,N_4653);
nor U7223 (N_7223,N_5695,N_5010);
nand U7224 (N_7224,N_5243,N_5877);
nor U7225 (N_7225,N_4190,N_4118);
nand U7226 (N_7226,N_4368,N_5830);
nor U7227 (N_7227,N_4906,N_5620);
or U7228 (N_7228,N_4824,N_5203);
nor U7229 (N_7229,N_4040,N_5315);
and U7230 (N_7230,N_5271,N_4565);
and U7231 (N_7231,N_5974,N_4483);
and U7232 (N_7232,N_4241,N_4643);
or U7233 (N_7233,N_5120,N_4782);
and U7234 (N_7234,N_4745,N_5835);
nor U7235 (N_7235,N_4979,N_5346);
nand U7236 (N_7236,N_4753,N_4059);
nand U7237 (N_7237,N_4207,N_5482);
nor U7238 (N_7238,N_5452,N_5547);
nor U7239 (N_7239,N_5040,N_5970);
or U7240 (N_7240,N_4230,N_5038);
nor U7241 (N_7241,N_5460,N_4074);
and U7242 (N_7242,N_4369,N_5051);
and U7243 (N_7243,N_5685,N_5317);
nand U7244 (N_7244,N_5005,N_4212);
xnor U7245 (N_7245,N_5908,N_5442);
nand U7246 (N_7246,N_5226,N_4415);
nand U7247 (N_7247,N_4814,N_5803);
xor U7248 (N_7248,N_5417,N_5410);
and U7249 (N_7249,N_4787,N_4840);
xnor U7250 (N_7250,N_4699,N_5980);
nand U7251 (N_7251,N_4258,N_4327);
nand U7252 (N_7252,N_4205,N_5552);
nor U7253 (N_7253,N_4173,N_5726);
nor U7254 (N_7254,N_4980,N_5055);
or U7255 (N_7255,N_4875,N_4655);
nor U7256 (N_7256,N_4859,N_4566);
nand U7257 (N_7257,N_4379,N_5572);
xnor U7258 (N_7258,N_5549,N_4532);
or U7259 (N_7259,N_5984,N_5678);
nand U7260 (N_7260,N_4254,N_5983);
nor U7261 (N_7261,N_5103,N_5687);
nor U7262 (N_7262,N_4675,N_4710);
and U7263 (N_7263,N_5642,N_4816);
nor U7264 (N_7264,N_5184,N_5849);
and U7265 (N_7265,N_4641,N_4363);
and U7266 (N_7266,N_5577,N_4076);
xnor U7267 (N_7267,N_5876,N_4327);
nand U7268 (N_7268,N_5964,N_5824);
nand U7269 (N_7269,N_5012,N_5014);
and U7270 (N_7270,N_5677,N_4164);
nand U7271 (N_7271,N_4381,N_4815);
or U7272 (N_7272,N_4032,N_5194);
nor U7273 (N_7273,N_5947,N_4134);
and U7274 (N_7274,N_5406,N_5896);
xnor U7275 (N_7275,N_5291,N_5069);
or U7276 (N_7276,N_5750,N_5980);
xor U7277 (N_7277,N_4581,N_5546);
xor U7278 (N_7278,N_5260,N_5052);
nor U7279 (N_7279,N_4171,N_4451);
or U7280 (N_7280,N_4520,N_5867);
and U7281 (N_7281,N_5998,N_4833);
nor U7282 (N_7282,N_5765,N_5928);
and U7283 (N_7283,N_5455,N_4340);
nand U7284 (N_7284,N_5341,N_5292);
xnor U7285 (N_7285,N_4203,N_4322);
xor U7286 (N_7286,N_5918,N_4661);
or U7287 (N_7287,N_5085,N_5000);
or U7288 (N_7288,N_5878,N_4875);
or U7289 (N_7289,N_4285,N_4785);
or U7290 (N_7290,N_5663,N_4996);
nor U7291 (N_7291,N_5716,N_5307);
nor U7292 (N_7292,N_4578,N_4120);
xor U7293 (N_7293,N_4057,N_5143);
nand U7294 (N_7294,N_4906,N_4501);
xor U7295 (N_7295,N_5007,N_5652);
or U7296 (N_7296,N_5339,N_4168);
and U7297 (N_7297,N_5233,N_4976);
nor U7298 (N_7298,N_4795,N_4574);
nor U7299 (N_7299,N_5705,N_4154);
or U7300 (N_7300,N_4175,N_5527);
and U7301 (N_7301,N_4132,N_4209);
nand U7302 (N_7302,N_4037,N_5729);
nand U7303 (N_7303,N_5611,N_4764);
and U7304 (N_7304,N_5915,N_5726);
xnor U7305 (N_7305,N_5648,N_5171);
nor U7306 (N_7306,N_4218,N_5562);
nand U7307 (N_7307,N_4449,N_5372);
nand U7308 (N_7308,N_4153,N_4019);
xnor U7309 (N_7309,N_5725,N_4955);
nor U7310 (N_7310,N_5064,N_4467);
xor U7311 (N_7311,N_5363,N_4323);
nor U7312 (N_7312,N_5001,N_5947);
or U7313 (N_7313,N_4137,N_5772);
or U7314 (N_7314,N_4682,N_5004);
nor U7315 (N_7315,N_4436,N_4715);
and U7316 (N_7316,N_4457,N_4950);
nor U7317 (N_7317,N_5025,N_4946);
or U7318 (N_7318,N_5634,N_4579);
nand U7319 (N_7319,N_5378,N_5726);
nand U7320 (N_7320,N_5455,N_5326);
or U7321 (N_7321,N_5650,N_5208);
or U7322 (N_7322,N_4860,N_5094);
xor U7323 (N_7323,N_4841,N_4531);
nor U7324 (N_7324,N_5358,N_5995);
nor U7325 (N_7325,N_4474,N_5379);
xor U7326 (N_7326,N_5214,N_4854);
and U7327 (N_7327,N_4475,N_5986);
nand U7328 (N_7328,N_5526,N_5483);
nand U7329 (N_7329,N_4619,N_4031);
and U7330 (N_7330,N_5089,N_4015);
nor U7331 (N_7331,N_4796,N_5514);
or U7332 (N_7332,N_5397,N_5982);
nand U7333 (N_7333,N_5262,N_5828);
xnor U7334 (N_7334,N_4541,N_5513);
nor U7335 (N_7335,N_5464,N_5660);
or U7336 (N_7336,N_4755,N_5930);
xnor U7337 (N_7337,N_5441,N_5931);
nand U7338 (N_7338,N_4022,N_5880);
nand U7339 (N_7339,N_5886,N_4608);
nand U7340 (N_7340,N_4842,N_4383);
and U7341 (N_7341,N_4573,N_4665);
xor U7342 (N_7342,N_4027,N_5814);
nor U7343 (N_7343,N_5871,N_5938);
or U7344 (N_7344,N_4267,N_5504);
xnor U7345 (N_7345,N_4384,N_5989);
and U7346 (N_7346,N_4005,N_5220);
xnor U7347 (N_7347,N_5085,N_5468);
nor U7348 (N_7348,N_5886,N_5739);
nand U7349 (N_7349,N_5541,N_5292);
and U7350 (N_7350,N_5752,N_4301);
nor U7351 (N_7351,N_4677,N_4705);
nor U7352 (N_7352,N_4969,N_4793);
nand U7353 (N_7353,N_4684,N_4340);
and U7354 (N_7354,N_4295,N_5255);
nand U7355 (N_7355,N_5534,N_4070);
or U7356 (N_7356,N_4203,N_4255);
and U7357 (N_7357,N_4892,N_4007);
and U7358 (N_7358,N_4692,N_5402);
nor U7359 (N_7359,N_5455,N_4791);
nor U7360 (N_7360,N_4852,N_5051);
and U7361 (N_7361,N_4171,N_4922);
and U7362 (N_7362,N_5140,N_5192);
xnor U7363 (N_7363,N_5571,N_4286);
or U7364 (N_7364,N_5322,N_5493);
nor U7365 (N_7365,N_4896,N_4356);
and U7366 (N_7366,N_5719,N_5167);
and U7367 (N_7367,N_5264,N_4293);
nor U7368 (N_7368,N_5487,N_5084);
and U7369 (N_7369,N_4171,N_5242);
xor U7370 (N_7370,N_5829,N_4589);
or U7371 (N_7371,N_5971,N_5235);
nand U7372 (N_7372,N_5977,N_5309);
nor U7373 (N_7373,N_4982,N_5598);
xnor U7374 (N_7374,N_5426,N_5452);
nand U7375 (N_7375,N_5158,N_4993);
xnor U7376 (N_7376,N_5064,N_5015);
nand U7377 (N_7377,N_4308,N_4280);
and U7378 (N_7378,N_5728,N_5671);
xnor U7379 (N_7379,N_4168,N_5087);
or U7380 (N_7380,N_5810,N_4821);
and U7381 (N_7381,N_5331,N_5235);
xor U7382 (N_7382,N_5653,N_5751);
and U7383 (N_7383,N_5361,N_5653);
nor U7384 (N_7384,N_5496,N_4938);
nor U7385 (N_7385,N_5567,N_5898);
nand U7386 (N_7386,N_5927,N_4707);
and U7387 (N_7387,N_4464,N_4058);
nand U7388 (N_7388,N_5793,N_4855);
nor U7389 (N_7389,N_5145,N_4250);
and U7390 (N_7390,N_4454,N_4817);
nor U7391 (N_7391,N_4931,N_5012);
nor U7392 (N_7392,N_4633,N_5741);
xnor U7393 (N_7393,N_5720,N_4274);
and U7394 (N_7394,N_5067,N_5336);
xnor U7395 (N_7395,N_4318,N_5797);
nand U7396 (N_7396,N_5665,N_4946);
xnor U7397 (N_7397,N_4081,N_4480);
xor U7398 (N_7398,N_4655,N_5497);
nor U7399 (N_7399,N_4809,N_5800);
nor U7400 (N_7400,N_5069,N_4623);
nand U7401 (N_7401,N_5392,N_4125);
or U7402 (N_7402,N_5172,N_4118);
nor U7403 (N_7403,N_5499,N_5438);
xnor U7404 (N_7404,N_5249,N_4628);
and U7405 (N_7405,N_5256,N_4509);
nand U7406 (N_7406,N_5454,N_5424);
xor U7407 (N_7407,N_4398,N_5663);
nor U7408 (N_7408,N_4601,N_5930);
or U7409 (N_7409,N_5154,N_4568);
xor U7410 (N_7410,N_4921,N_4914);
xnor U7411 (N_7411,N_5765,N_4173);
or U7412 (N_7412,N_4507,N_5046);
and U7413 (N_7413,N_5202,N_5805);
xor U7414 (N_7414,N_5891,N_4464);
nor U7415 (N_7415,N_5046,N_4786);
or U7416 (N_7416,N_4347,N_5396);
or U7417 (N_7417,N_5044,N_4020);
and U7418 (N_7418,N_5194,N_5147);
xnor U7419 (N_7419,N_5281,N_4748);
nand U7420 (N_7420,N_5194,N_4146);
nor U7421 (N_7421,N_4513,N_4209);
nand U7422 (N_7422,N_4952,N_5286);
and U7423 (N_7423,N_4635,N_4938);
and U7424 (N_7424,N_5232,N_5615);
nor U7425 (N_7425,N_4035,N_4940);
xnor U7426 (N_7426,N_4089,N_5937);
nor U7427 (N_7427,N_5217,N_5422);
nor U7428 (N_7428,N_4425,N_4864);
nand U7429 (N_7429,N_5301,N_4923);
or U7430 (N_7430,N_5493,N_5047);
xor U7431 (N_7431,N_4767,N_4071);
xnor U7432 (N_7432,N_4219,N_5542);
nand U7433 (N_7433,N_4320,N_5937);
nand U7434 (N_7434,N_4639,N_4699);
xnor U7435 (N_7435,N_5472,N_5698);
nor U7436 (N_7436,N_4356,N_4587);
and U7437 (N_7437,N_4558,N_5983);
and U7438 (N_7438,N_5758,N_4284);
nand U7439 (N_7439,N_4068,N_5973);
nand U7440 (N_7440,N_5246,N_5354);
or U7441 (N_7441,N_4450,N_4223);
and U7442 (N_7442,N_5753,N_5492);
or U7443 (N_7443,N_5830,N_5545);
xor U7444 (N_7444,N_4403,N_5410);
nor U7445 (N_7445,N_4738,N_5816);
nor U7446 (N_7446,N_5798,N_5410);
or U7447 (N_7447,N_4104,N_5624);
xor U7448 (N_7448,N_4575,N_4130);
and U7449 (N_7449,N_4869,N_5777);
or U7450 (N_7450,N_4093,N_4719);
nor U7451 (N_7451,N_4056,N_4048);
nand U7452 (N_7452,N_4591,N_5023);
xnor U7453 (N_7453,N_4981,N_4246);
xor U7454 (N_7454,N_5755,N_4864);
xnor U7455 (N_7455,N_4180,N_5113);
nand U7456 (N_7456,N_5824,N_5244);
nand U7457 (N_7457,N_5140,N_5307);
nand U7458 (N_7458,N_5401,N_4356);
nor U7459 (N_7459,N_4596,N_4051);
xnor U7460 (N_7460,N_5357,N_5564);
or U7461 (N_7461,N_5867,N_4365);
nand U7462 (N_7462,N_5608,N_5921);
nor U7463 (N_7463,N_5700,N_4044);
nand U7464 (N_7464,N_5935,N_5898);
or U7465 (N_7465,N_4144,N_4328);
xor U7466 (N_7466,N_5179,N_5656);
xor U7467 (N_7467,N_5159,N_5789);
xor U7468 (N_7468,N_4339,N_5151);
and U7469 (N_7469,N_4745,N_5111);
xnor U7470 (N_7470,N_5173,N_5230);
nand U7471 (N_7471,N_4794,N_4607);
or U7472 (N_7472,N_5467,N_4980);
or U7473 (N_7473,N_5027,N_5832);
xor U7474 (N_7474,N_4420,N_5452);
nand U7475 (N_7475,N_5009,N_5102);
nor U7476 (N_7476,N_5911,N_5888);
xnor U7477 (N_7477,N_4336,N_4959);
nand U7478 (N_7478,N_5575,N_5354);
nand U7479 (N_7479,N_4083,N_4812);
and U7480 (N_7480,N_5357,N_5158);
xnor U7481 (N_7481,N_5369,N_5507);
and U7482 (N_7482,N_4351,N_5657);
or U7483 (N_7483,N_5674,N_5074);
and U7484 (N_7484,N_4267,N_5255);
xnor U7485 (N_7485,N_4640,N_4019);
and U7486 (N_7486,N_5852,N_4567);
or U7487 (N_7487,N_5139,N_4420);
nor U7488 (N_7488,N_5863,N_5652);
nand U7489 (N_7489,N_4052,N_4535);
nor U7490 (N_7490,N_4096,N_5692);
nand U7491 (N_7491,N_5329,N_4253);
xnor U7492 (N_7492,N_4673,N_5958);
xnor U7493 (N_7493,N_4313,N_5148);
xor U7494 (N_7494,N_5936,N_5871);
nor U7495 (N_7495,N_5986,N_5246);
or U7496 (N_7496,N_5836,N_4154);
or U7497 (N_7497,N_5908,N_4453);
nor U7498 (N_7498,N_4759,N_5199);
nor U7499 (N_7499,N_5221,N_5460);
or U7500 (N_7500,N_4015,N_4059);
xor U7501 (N_7501,N_5033,N_4613);
and U7502 (N_7502,N_5108,N_4268);
and U7503 (N_7503,N_4215,N_5577);
and U7504 (N_7504,N_4820,N_5017);
nor U7505 (N_7505,N_4559,N_4684);
nor U7506 (N_7506,N_4946,N_5847);
nor U7507 (N_7507,N_5447,N_5350);
or U7508 (N_7508,N_5628,N_4250);
xor U7509 (N_7509,N_5937,N_4158);
and U7510 (N_7510,N_4448,N_4173);
and U7511 (N_7511,N_4513,N_4191);
nand U7512 (N_7512,N_4351,N_4611);
nand U7513 (N_7513,N_4511,N_5428);
nand U7514 (N_7514,N_4841,N_5373);
or U7515 (N_7515,N_4046,N_4421);
nor U7516 (N_7516,N_4654,N_5146);
nand U7517 (N_7517,N_5875,N_4618);
nor U7518 (N_7518,N_5632,N_5001);
nor U7519 (N_7519,N_4758,N_5277);
and U7520 (N_7520,N_5868,N_5433);
nand U7521 (N_7521,N_4808,N_5413);
xor U7522 (N_7522,N_5577,N_4868);
and U7523 (N_7523,N_5088,N_4341);
and U7524 (N_7524,N_5147,N_5084);
nor U7525 (N_7525,N_4471,N_5525);
or U7526 (N_7526,N_4982,N_5358);
nand U7527 (N_7527,N_5698,N_4212);
nand U7528 (N_7528,N_5997,N_4706);
nand U7529 (N_7529,N_5369,N_4728);
xnor U7530 (N_7530,N_5529,N_5953);
nand U7531 (N_7531,N_5420,N_5404);
nand U7532 (N_7532,N_5760,N_4477);
or U7533 (N_7533,N_4831,N_5947);
nor U7534 (N_7534,N_5545,N_4884);
and U7535 (N_7535,N_5645,N_4388);
nor U7536 (N_7536,N_4061,N_5151);
nor U7537 (N_7537,N_4519,N_5809);
nand U7538 (N_7538,N_4578,N_5918);
nand U7539 (N_7539,N_5964,N_4803);
xor U7540 (N_7540,N_5236,N_5250);
nand U7541 (N_7541,N_4310,N_5137);
nand U7542 (N_7542,N_4806,N_4338);
nor U7543 (N_7543,N_5891,N_4287);
or U7544 (N_7544,N_4313,N_5657);
nor U7545 (N_7545,N_4643,N_4780);
xnor U7546 (N_7546,N_5288,N_5537);
or U7547 (N_7547,N_4350,N_4562);
and U7548 (N_7548,N_5213,N_5144);
nand U7549 (N_7549,N_4461,N_4965);
nor U7550 (N_7550,N_5249,N_4088);
xor U7551 (N_7551,N_4653,N_4085);
and U7552 (N_7552,N_5733,N_5373);
nor U7553 (N_7553,N_5056,N_5141);
or U7554 (N_7554,N_5425,N_5223);
or U7555 (N_7555,N_5113,N_5603);
nor U7556 (N_7556,N_5327,N_5387);
and U7557 (N_7557,N_5085,N_4176);
nand U7558 (N_7558,N_5730,N_5189);
nand U7559 (N_7559,N_4576,N_4088);
or U7560 (N_7560,N_4205,N_5654);
and U7561 (N_7561,N_4379,N_5228);
nor U7562 (N_7562,N_5052,N_4779);
nor U7563 (N_7563,N_4689,N_5495);
xnor U7564 (N_7564,N_5043,N_5691);
nand U7565 (N_7565,N_4866,N_4716);
nor U7566 (N_7566,N_5225,N_5816);
xnor U7567 (N_7567,N_4845,N_5820);
nand U7568 (N_7568,N_4308,N_5784);
nor U7569 (N_7569,N_5558,N_5389);
xor U7570 (N_7570,N_5597,N_4034);
nor U7571 (N_7571,N_4561,N_4743);
nand U7572 (N_7572,N_5400,N_4612);
and U7573 (N_7573,N_5471,N_4967);
or U7574 (N_7574,N_4431,N_5825);
xor U7575 (N_7575,N_5743,N_5198);
nor U7576 (N_7576,N_4411,N_5640);
nor U7577 (N_7577,N_4702,N_4562);
xnor U7578 (N_7578,N_5717,N_5519);
nand U7579 (N_7579,N_4637,N_5865);
or U7580 (N_7580,N_5369,N_5564);
nor U7581 (N_7581,N_4306,N_5207);
nand U7582 (N_7582,N_5868,N_4680);
xor U7583 (N_7583,N_5366,N_4607);
or U7584 (N_7584,N_5123,N_4410);
or U7585 (N_7585,N_5347,N_5390);
nor U7586 (N_7586,N_4675,N_4891);
or U7587 (N_7587,N_4629,N_4909);
nor U7588 (N_7588,N_4159,N_4846);
and U7589 (N_7589,N_5566,N_5315);
or U7590 (N_7590,N_5073,N_5898);
nand U7591 (N_7591,N_4584,N_4751);
and U7592 (N_7592,N_5101,N_4959);
nor U7593 (N_7593,N_5360,N_5596);
xnor U7594 (N_7594,N_5331,N_4313);
nor U7595 (N_7595,N_5575,N_4036);
xnor U7596 (N_7596,N_4353,N_5008);
or U7597 (N_7597,N_5718,N_4108);
nor U7598 (N_7598,N_4954,N_5425);
and U7599 (N_7599,N_5981,N_5772);
nor U7600 (N_7600,N_4050,N_5866);
or U7601 (N_7601,N_5155,N_4240);
xor U7602 (N_7602,N_5614,N_5713);
nor U7603 (N_7603,N_5283,N_5634);
nor U7604 (N_7604,N_4596,N_5013);
nor U7605 (N_7605,N_4942,N_4107);
nand U7606 (N_7606,N_5770,N_4657);
xor U7607 (N_7607,N_5948,N_5455);
and U7608 (N_7608,N_5410,N_5902);
and U7609 (N_7609,N_5759,N_4479);
or U7610 (N_7610,N_4532,N_5020);
and U7611 (N_7611,N_5347,N_4494);
xnor U7612 (N_7612,N_4944,N_4581);
and U7613 (N_7613,N_5913,N_5311);
nand U7614 (N_7614,N_5910,N_5422);
nand U7615 (N_7615,N_4843,N_4343);
nand U7616 (N_7616,N_5488,N_5269);
nand U7617 (N_7617,N_5059,N_5042);
or U7618 (N_7618,N_4604,N_4273);
xnor U7619 (N_7619,N_4788,N_4477);
and U7620 (N_7620,N_5730,N_5107);
or U7621 (N_7621,N_4868,N_5236);
xor U7622 (N_7622,N_5357,N_4122);
or U7623 (N_7623,N_5716,N_5536);
xor U7624 (N_7624,N_4205,N_4662);
xnor U7625 (N_7625,N_5611,N_5154);
nor U7626 (N_7626,N_5296,N_5957);
nand U7627 (N_7627,N_4481,N_5890);
xnor U7628 (N_7628,N_4092,N_5413);
or U7629 (N_7629,N_4307,N_4894);
nor U7630 (N_7630,N_5695,N_4978);
and U7631 (N_7631,N_5393,N_4531);
and U7632 (N_7632,N_4983,N_4132);
or U7633 (N_7633,N_5778,N_5228);
nor U7634 (N_7634,N_4223,N_5442);
or U7635 (N_7635,N_4958,N_4224);
and U7636 (N_7636,N_4175,N_4688);
or U7637 (N_7637,N_5631,N_5484);
nand U7638 (N_7638,N_4420,N_5383);
or U7639 (N_7639,N_5947,N_4105);
nor U7640 (N_7640,N_4899,N_5577);
nand U7641 (N_7641,N_4336,N_5754);
or U7642 (N_7642,N_5122,N_5799);
nor U7643 (N_7643,N_5371,N_4008);
xnor U7644 (N_7644,N_4038,N_5080);
or U7645 (N_7645,N_5557,N_4209);
nor U7646 (N_7646,N_4532,N_4858);
and U7647 (N_7647,N_4543,N_5231);
nor U7648 (N_7648,N_5002,N_4164);
nand U7649 (N_7649,N_5729,N_4422);
and U7650 (N_7650,N_4369,N_4982);
nand U7651 (N_7651,N_5894,N_5705);
or U7652 (N_7652,N_4043,N_4535);
nand U7653 (N_7653,N_4750,N_4007);
xor U7654 (N_7654,N_4089,N_4148);
nand U7655 (N_7655,N_4487,N_4641);
and U7656 (N_7656,N_5730,N_4753);
xnor U7657 (N_7657,N_5068,N_5862);
or U7658 (N_7658,N_5923,N_5646);
and U7659 (N_7659,N_4426,N_5276);
and U7660 (N_7660,N_5141,N_5994);
xor U7661 (N_7661,N_5932,N_4661);
xor U7662 (N_7662,N_5409,N_5482);
nor U7663 (N_7663,N_5257,N_5330);
or U7664 (N_7664,N_4077,N_5457);
xor U7665 (N_7665,N_4395,N_4250);
or U7666 (N_7666,N_4801,N_5576);
and U7667 (N_7667,N_4724,N_5583);
nand U7668 (N_7668,N_4150,N_5462);
or U7669 (N_7669,N_4486,N_5454);
nand U7670 (N_7670,N_5734,N_4047);
and U7671 (N_7671,N_4792,N_4272);
nand U7672 (N_7672,N_5715,N_4541);
and U7673 (N_7673,N_5112,N_4918);
nor U7674 (N_7674,N_4437,N_5014);
xnor U7675 (N_7675,N_5181,N_5460);
or U7676 (N_7676,N_4787,N_4171);
and U7677 (N_7677,N_4877,N_5701);
or U7678 (N_7678,N_4989,N_5397);
nor U7679 (N_7679,N_5616,N_5765);
nand U7680 (N_7680,N_5358,N_5391);
and U7681 (N_7681,N_5745,N_4003);
or U7682 (N_7682,N_4498,N_5758);
nor U7683 (N_7683,N_5859,N_5595);
and U7684 (N_7684,N_5390,N_5625);
and U7685 (N_7685,N_5566,N_4229);
and U7686 (N_7686,N_5162,N_4897);
nand U7687 (N_7687,N_4426,N_4420);
nor U7688 (N_7688,N_5310,N_5793);
and U7689 (N_7689,N_4715,N_4172);
or U7690 (N_7690,N_5925,N_4233);
and U7691 (N_7691,N_4090,N_4372);
nand U7692 (N_7692,N_4975,N_5962);
nor U7693 (N_7693,N_5591,N_5282);
or U7694 (N_7694,N_4167,N_5369);
xnor U7695 (N_7695,N_4223,N_5441);
xor U7696 (N_7696,N_4248,N_4715);
nor U7697 (N_7697,N_5308,N_5537);
and U7698 (N_7698,N_5794,N_4179);
and U7699 (N_7699,N_5377,N_4873);
xnor U7700 (N_7700,N_5473,N_4032);
xor U7701 (N_7701,N_5667,N_4037);
nor U7702 (N_7702,N_4392,N_5323);
xnor U7703 (N_7703,N_4389,N_5841);
xor U7704 (N_7704,N_5206,N_4603);
nand U7705 (N_7705,N_5872,N_5326);
or U7706 (N_7706,N_4488,N_4511);
nor U7707 (N_7707,N_5810,N_5692);
and U7708 (N_7708,N_5188,N_4738);
xor U7709 (N_7709,N_5091,N_4269);
or U7710 (N_7710,N_4766,N_5448);
and U7711 (N_7711,N_4096,N_4516);
and U7712 (N_7712,N_5559,N_5270);
or U7713 (N_7713,N_5929,N_5777);
and U7714 (N_7714,N_5344,N_4702);
nor U7715 (N_7715,N_4488,N_4999);
nor U7716 (N_7716,N_5072,N_4718);
and U7717 (N_7717,N_5221,N_5558);
or U7718 (N_7718,N_5952,N_4609);
or U7719 (N_7719,N_5942,N_4571);
and U7720 (N_7720,N_4743,N_5738);
nand U7721 (N_7721,N_5530,N_4000);
xor U7722 (N_7722,N_4031,N_4290);
or U7723 (N_7723,N_5094,N_5000);
nor U7724 (N_7724,N_4684,N_4919);
nand U7725 (N_7725,N_5167,N_4603);
xor U7726 (N_7726,N_4179,N_4824);
or U7727 (N_7727,N_5380,N_5656);
xor U7728 (N_7728,N_4644,N_4689);
nand U7729 (N_7729,N_4589,N_4953);
nor U7730 (N_7730,N_5974,N_5379);
or U7731 (N_7731,N_4689,N_4322);
and U7732 (N_7732,N_4739,N_4281);
nor U7733 (N_7733,N_5688,N_5091);
or U7734 (N_7734,N_5157,N_4427);
nand U7735 (N_7735,N_5414,N_5817);
xor U7736 (N_7736,N_4934,N_5617);
xor U7737 (N_7737,N_5748,N_4170);
xor U7738 (N_7738,N_5604,N_4874);
and U7739 (N_7739,N_5818,N_5675);
nand U7740 (N_7740,N_5360,N_4884);
nor U7741 (N_7741,N_4054,N_4528);
nor U7742 (N_7742,N_5422,N_5944);
xnor U7743 (N_7743,N_5838,N_4961);
xnor U7744 (N_7744,N_5789,N_5869);
or U7745 (N_7745,N_4839,N_5958);
nor U7746 (N_7746,N_4106,N_5373);
nand U7747 (N_7747,N_4482,N_4331);
nor U7748 (N_7748,N_5290,N_5613);
nand U7749 (N_7749,N_4853,N_4981);
xor U7750 (N_7750,N_4065,N_4912);
and U7751 (N_7751,N_5729,N_4147);
nor U7752 (N_7752,N_5755,N_4642);
and U7753 (N_7753,N_5450,N_4886);
nor U7754 (N_7754,N_5274,N_4095);
nor U7755 (N_7755,N_4257,N_4603);
nand U7756 (N_7756,N_5100,N_4669);
and U7757 (N_7757,N_4824,N_5185);
xnor U7758 (N_7758,N_5010,N_4914);
and U7759 (N_7759,N_4964,N_5976);
nor U7760 (N_7760,N_5026,N_5882);
nor U7761 (N_7761,N_5036,N_5122);
or U7762 (N_7762,N_4736,N_4663);
nor U7763 (N_7763,N_4250,N_5349);
and U7764 (N_7764,N_5120,N_4533);
xnor U7765 (N_7765,N_4664,N_4065);
xor U7766 (N_7766,N_4700,N_5375);
xnor U7767 (N_7767,N_4284,N_5726);
nor U7768 (N_7768,N_4018,N_5390);
and U7769 (N_7769,N_5171,N_5304);
nor U7770 (N_7770,N_5020,N_5840);
xor U7771 (N_7771,N_5589,N_5012);
or U7772 (N_7772,N_4855,N_4415);
nor U7773 (N_7773,N_4660,N_4093);
nand U7774 (N_7774,N_4973,N_5336);
or U7775 (N_7775,N_5603,N_5347);
or U7776 (N_7776,N_4400,N_4578);
or U7777 (N_7777,N_5014,N_5779);
and U7778 (N_7778,N_4719,N_5457);
nor U7779 (N_7779,N_5564,N_4159);
or U7780 (N_7780,N_4677,N_4164);
or U7781 (N_7781,N_4594,N_4190);
nand U7782 (N_7782,N_4120,N_5827);
or U7783 (N_7783,N_4444,N_5226);
and U7784 (N_7784,N_5724,N_4967);
nor U7785 (N_7785,N_4372,N_5168);
nand U7786 (N_7786,N_4553,N_4579);
and U7787 (N_7787,N_4882,N_4753);
xor U7788 (N_7788,N_5293,N_5078);
nor U7789 (N_7789,N_5544,N_4213);
nor U7790 (N_7790,N_4131,N_5963);
nand U7791 (N_7791,N_5578,N_4101);
xnor U7792 (N_7792,N_4649,N_5949);
or U7793 (N_7793,N_5699,N_4367);
nor U7794 (N_7794,N_4413,N_4250);
xnor U7795 (N_7795,N_5319,N_4733);
nand U7796 (N_7796,N_5123,N_4071);
or U7797 (N_7797,N_4545,N_5065);
and U7798 (N_7798,N_5827,N_4192);
nand U7799 (N_7799,N_4375,N_4640);
and U7800 (N_7800,N_5338,N_5425);
and U7801 (N_7801,N_5238,N_4431);
nor U7802 (N_7802,N_4970,N_4278);
or U7803 (N_7803,N_4137,N_4930);
nor U7804 (N_7804,N_5610,N_4195);
or U7805 (N_7805,N_4125,N_5304);
and U7806 (N_7806,N_5002,N_4130);
xor U7807 (N_7807,N_5101,N_5552);
or U7808 (N_7808,N_5983,N_5905);
nor U7809 (N_7809,N_4303,N_5471);
nand U7810 (N_7810,N_4700,N_4385);
xor U7811 (N_7811,N_5764,N_4047);
nor U7812 (N_7812,N_4273,N_5123);
and U7813 (N_7813,N_5425,N_4656);
xnor U7814 (N_7814,N_5709,N_5014);
nand U7815 (N_7815,N_4294,N_4917);
nand U7816 (N_7816,N_5279,N_5108);
or U7817 (N_7817,N_5549,N_5170);
nand U7818 (N_7818,N_4917,N_5150);
or U7819 (N_7819,N_5366,N_5649);
or U7820 (N_7820,N_5878,N_5705);
xor U7821 (N_7821,N_4858,N_4691);
nand U7822 (N_7822,N_5814,N_5177);
nor U7823 (N_7823,N_4361,N_4320);
nand U7824 (N_7824,N_4716,N_5019);
xnor U7825 (N_7825,N_4595,N_5794);
or U7826 (N_7826,N_4537,N_4126);
and U7827 (N_7827,N_4481,N_5741);
nor U7828 (N_7828,N_5981,N_4477);
nor U7829 (N_7829,N_5069,N_5146);
and U7830 (N_7830,N_4722,N_5354);
nor U7831 (N_7831,N_5072,N_4578);
nor U7832 (N_7832,N_5289,N_4674);
nor U7833 (N_7833,N_4088,N_4163);
and U7834 (N_7834,N_4086,N_5614);
and U7835 (N_7835,N_4160,N_5108);
and U7836 (N_7836,N_5082,N_4596);
nor U7837 (N_7837,N_4507,N_5917);
and U7838 (N_7838,N_4863,N_4589);
or U7839 (N_7839,N_4210,N_5340);
and U7840 (N_7840,N_5768,N_4767);
nor U7841 (N_7841,N_5797,N_4217);
nand U7842 (N_7842,N_5223,N_4903);
xnor U7843 (N_7843,N_4469,N_4190);
or U7844 (N_7844,N_5229,N_4206);
nor U7845 (N_7845,N_4724,N_5722);
nor U7846 (N_7846,N_4337,N_4748);
nor U7847 (N_7847,N_5886,N_4046);
or U7848 (N_7848,N_4521,N_4457);
or U7849 (N_7849,N_4813,N_4878);
nor U7850 (N_7850,N_5079,N_5895);
nand U7851 (N_7851,N_5412,N_5854);
nor U7852 (N_7852,N_4679,N_5381);
nand U7853 (N_7853,N_4989,N_5757);
and U7854 (N_7854,N_5799,N_5097);
xor U7855 (N_7855,N_4030,N_4881);
nand U7856 (N_7856,N_5449,N_5694);
nor U7857 (N_7857,N_4609,N_5446);
and U7858 (N_7858,N_5319,N_4087);
nand U7859 (N_7859,N_4013,N_4154);
nor U7860 (N_7860,N_5663,N_4567);
nand U7861 (N_7861,N_4993,N_5662);
nor U7862 (N_7862,N_4739,N_5302);
nor U7863 (N_7863,N_4545,N_4092);
nand U7864 (N_7864,N_4113,N_5577);
and U7865 (N_7865,N_5508,N_5879);
nand U7866 (N_7866,N_5780,N_4524);
nor U7867 (N_7867,N_5139,N_4194);
xor U7868 (N_7868,N_5439,N_5007);
xor U7869 (N_7869,N_5310,N_5006);
and U7870 (N_7870,N_5109,N_5596);
nor U7871 (N_7871,N_4252,N_5116);
nor U7872 (N_7872,N_4406,N_4358);
nor U7873 (N_7873,N_5911,N_5628);
or U7874 (N_7874,N_4176,N_5841);
or U7875 (N_7875,N_4840,N_4387);
and U7876 (N_7876,N_5653,N_4416);
nor U7877 (N_7877,N_5448,N_4886);
nor U7878 (N_7878,N_5343,N_5723);
or U7879 (N_7879,N_5667,N_4531);
or U7880 (N_7880,N_4407,N_5312);
nand U7881 (N_7881,N_4944,N_4741);
xor U7882 (N_7882,N_4855,N_4220);
nand U7883 (N_7883,N_4245,N_4472);
and U7884 (N_7884,N_5037,N_5410);
or U7885 (N_7885,N_5758,N_4343);
xnor U7886 (N_7886,N_4467,N_4267);
and U7887 (N_7887,N_4132,N_5303);
or U7888 (N_7888,N_4765,N_5710);
xor U7889 (N_7889,N_4039,N_4759);
and U7890 (N_7890,N_4154,N_4295);
and U7891 (N_7891,N_5490,N_4990);
xnor U7892 (N_7892,N_5440,N_5198);
or U7893 (N_7893,N_4770,N_4331);
or U7894 (N_7894,N_5683,N_5042);
or U7895 (N_7895,N_4750,N_5612);
or U7896 (N_7896,N_5379,N_5966);
nand U7897 (N_7897,N_4481,N_4685);
nand U7898 (N_7898,N_4128,N_5470);
and U7899 (N_7899,N_5596,N_4800);
or U7900 (N_7900,N_4108,N_4298);
nand U7901 (N_7901,N_4390,N_4674);
and U7902 (N_7902,N_5463,N_4667);
or U7903 (N_7903,N_5654,N_4691);
nand U7904 (N_7904,N_4313,N_5293);
or U7905 (N_7905,N_5292,N_5231);
xnor U7906 (N_7906,N_5369,N_5931);
or U7907 (N_7907,N_5432,N_4096);
and U7908 (N_7908,N_5728,N_5083);
nand U7909 (N_7909,N_5182,N_5185);
nor U7910 (N_7910,N_5885,N_5089);
and U7911 (N_7911,N_4222,N_4783);
nand U7912 (N_7912,N_5811,N_4615);
and U7913 (N_7913,N_4284,N_4551);
or U7914 (N_7914,N_4800,N_5756);
nand U7915 (N_7915,N_4040,N_5293);
nor U7916 (N_7916,N_5472,N_4833);
or U7917 (N_7917,N_4414,N_4724);
xor U7918 (N_7918,N_5115,N_5530);
or U7919 (N_7919,N_4533,N_5543);
nand U7920 (N_7920,N_4427,N_4860);
or U7921 (N_7921,N_5828,N_4617);
or U7922 (N_7922,N_4513,N_4640);
nor U7923 (N_7923,N_4383,N_5168);
or U7924 (N_7924,N_5760,N_5752);
and U7925 (N_7925,N_4084,N_5715);
xnor U7926 (N_7926,N_5994,N_5655);
xnor U7927 (N_7927,N_5904,N_4050);
or U7928 (N_7928,N_5212,N_4954);
nand U7929 (N_7929,N_4613,N_4957);
nor U7930 (N_7930,N_5112,N_5602);
nand U7931 (N_7931,N_5224,N_4339);
nand U7932 (N_7932,N_5932,N_5336);
xor U7933 (N_7933,N_4639,N_5281);
nor U7934 (N_7934,N_5368,N_5418);
nand U7935 (N_7935,N_5635,N_5754);
or U7936 (N_7936,N_5878,N_4535);
and U7937 (N_7937,N_4788,N_5196);
and U7938 (N_7938,N_4190,N_4189);
xnor U7939 (N_7939,N_5157,N_5288);
xnor U7940 (N_7940,N_4061,N_4666);
nor U7941 (N_7941,N_4159,N_5571);
or U7942 (N_7942,N_4220,N_4659);
nand U7943 (N_7943,N_5199,N_5540);
or U7944 (N_7944,N_4673,N_4208);
and U7945 (N_7945,N_5955,N_4809);
and U7946 (N_7946,N_4598,N_4399);
nor U7947 (N_7947,N_5670,N_4405);
xnor U7948 (N_7948,N_5946,N_5889);
and U7949 (N_7949,N_5659,N_4206);
xor U7950 (N_7950,N_4281,N_4990);
or U7951 (N_7951,N_4439,N_4010);
nand U7952 (N_7952,N_4616,N_4127);
and U7953 (N_7953,N_4784,N_5879);
or U7954 (N_7954,N_4047,N_4294);
or U7955 (N_7955,N_4670,N_4762);
nor U7956 (N_7956,N_5374,N_5998);
nor U7957 (N_7957,N_4954,N_4727);
xor U7958 (N_7958,N_5253,N_4002);
or U7959 (N_7959,N_5005,N_5381);
and U7960 (N_7960,N_4692,N_4840);
xnor U7961 (N_7961,N_5134,N_4802);
nor U7962 (N_7962,N_4257,N_4347);
nor U7963 (N_7963,N_5979,N_5772);
xor U7964 (N_7964,N_4939,N_5429);
or U7965 (N_7965,N_4742,N_5425);
or U7966 (N_7966,N_4134,N_5747);
nor U7967 (N_7967,N_4627,N_4548);
or U7968 (N_7968,N_4295,N_4089);
nand U7969 (N_7969,N_5136,N_5448);
or U7970 (N_7970,N_4069,N_4277);
or U7971 (N_7971,N_4662,N_5986);
or U7972 (N_7972,N_5820,N_4084);
or U7973 (N_7973,N_4825,N_4548);
nand U7974 (N_7974,N_5543,N_5313);
xor U7975 (N_7975,N_5921,N_5744);
xor U7976 (N_7976,N_4226,N_5659);
xor U7977 (N_7977,N_4542,N_5118);
nand U7978 (N_7978,N_4131,N_5395);
or U7979 (N_7979,N_5458,N_5999);
and U7980 (N_7980,N_4466,N_4244);
xnor U7981 (N_7981,N_5750,N_5432);
and U7982 (N_7982,N_5489,N_5720);
xnor U7983 (N_7983,N_5494,N_5366);
xnor U7984 (N_7984,N_4050,N_5942);
nand U7985 (N_7985,N_4165,N_4311);
xnor U7986 (N_7986,N_4665,N_5009);
xor U7987 (N_7987,N_5260,N_5344);
xnor U7988 (N_7988,N_5635,N_4575);
and U7989 (N_7989,N_5518,N_5668);
or U7990 (N_7990,N_4081,N_5674);
or U7991 (N_7991,N_5896,N_4543);
nand U7992 (N_7992,N_4585,N_4587);
and U7993 (N_7993,N_5923,N_4426);
and U7994 (N_7994,N_4697,N_5022);
and U7995 (N_7995,N_5160,N_5010);
nand U7996 (N_7996,N_4780,N_4558);
and U7997 (N_7997,N_5115,N_5330);
xor U7998 (N_7998,N_5782,N_5028);
or U7999 (N_7999,N_4949,N_4708);
or U8000 (N_8000,N_6861,N_7505);
or U8001 (N_8001,N_6512,N_7145);
xor U8002 (N_8002,N_7993,N_6938);
xnor U8003 (N_8003,N_7517,N_6980);
xor U8004 (N_8004,N_6846,N_7875);
or U8005 (N_8005,N_6684,N_6180);
and U8006 (N_8006,N_6478,N_7708);
or U8007 (N_8007,N_7473,N_6013);
nand U8008 (N_8008,N_6933,N_7114);
nand U8009 (N_8009,N_6887,N_6853);
nor U8010 (N_8010,N_6648,N_7658);
nor U8011 (N_8011,N_6185,N_6146);
nor U8012 (N_8012,N_7839,N_7846);
or U8013 (N_8013,N_6667,N_6396);
xor U8014 (N_8014,N_7812,N_6934);
nor U8015 (N_8015,N_6497,N_7397);
and U8016 (N_8016,N_7332,N_6636);
or U8017 (N_8017,N_6754,N_6564);
nor U8018 (N_8018,N_7841,N_7766);
and U8019 (N_8019,N_7444,N_7238);
and U8020 (N_8020,N_7956,N_7244);
and U8021 (N_8021,N_6895,N_6401);
xnor U8022 (N_8022,N_6014,N_6447);
and U8023 (N_8023,N_6457,N_6311);
and U8024 (N_8024,N_6438,N_7992);
nor U8025 (N_8025,N_6350,N_7831);
nand U8026 (N_8026,N_6331,N_6434);
and U8027 (N_8027,N_7110,N_7698);
nor U8028 (N_8028,N_6238,N_7175);
or U8029 (N_8029,N_7489,N_7929);
nand U8030 (N_8030,N_7325,N_6620);
nor U8031 (N_8031,N_6202,N_6380);
nand U8032 (N_8032,N_6763,N_7240);
nand U8033 (N_8033,N_6612,N_6417);
nand U8034 (N_8034,N_7746,N_7322);
nor U8035 (N_8035,N_7163,N_7520);
and U8036 (N_8036,N_7524,N_7609);
nand U8037 (N_8037,N_7748,N_6702);
nand U8038 (N_8038,N_7646,N_6394);
nor U8039 (N_8039,N_6699,N_6000);
nand U8040 (N_8040,N_7883,N_7387);
and U8041 (N_8041,N_7030,N_7945);
nand U8042 (N_8042,N_7633,N_7734);
nor U8043 (N_8043,N_6217,N_6493);
xnor U8044 (N_8044,N_7765,N_6627);
nand U8045 (N_8045,N_6161,N_7369);
xnor U8046 (N_8046,N_7394,N_7869);
nor U8047 (N_8047,N_7068,N_6662);
nor U8048 (N_8048,N_7578,N_7177);
or U8049 (N_8049,N_6413,N_7006);
and U8050 (N_8050,N_7303,N_6642);
nand U8051 (N_8051,N_7196,N_6558);
or U8052 (N_8052,N_6506,N_7521);
and U8053 (N_8053,N_7009,N_6496);
nor U8054 (N_8054,N_7176,N_6208);
nor U8055 (N_8055,N_7800,N_6097);
nor U8056 (N_8056,N_6461,N_7095);
nor U8057 (N_8057,N_6539,N_6927);
or U8058 (N_8058,N_7446,N_6542);
and U8059 (N_8059,N_6357,N_7057);
nand U8060 (N_8060,N_6130,N_7773);
nand U8061 (N_8061,N_6163,N_7208);
and U8062 (N_8062,N_6544,N_6373);
nand U8063 (N_8063,N_7591,N_7179);
or U8064 (N_8064,N_6525,N_7378);
nor U8065 (N_8065,N_6147,N_7349);
nand U8066 (N_8066,N_6116,N_7648);
xnor U8067 (N_8067,N_6982,N_6724);
nand U8068 (N_8068,N_6638,N_6068);
or U8069 (N_8069,N_7552,N_7126);
and U8070 (N_8070,N_6640,N_6035);
nor U8071 (N_8071,N_6969,N_6428);
nor U8072 (N_8072,N_7543,N_7485);
nand U8073 (N_8073,N_6986,N_6759);
or U8074 (N_8074,N_6309,N_6235);
and U8075 (N_8075,N_6641,N_7226);
and U8076 (N_8076,N_6826,N_6864);
or U8077 (N_8077,N_6440,N_6067);
xnor U8078 (N_8078,N_6753,N_6231);
xnor U8079 (N_8079,N_7863,N_7361);
nor U8080 (N_8080,N_6837,N_6211);
nand U8081 (N_8081,N_6418,N_7930);
and U8082 (N_8082,N_7630,N_7724);
or U8083 (N_8083,N_7085,N_6098);
nand U8084 (N_8084,N_6928,N_6463);
xnor U8085 (N_8085,N_6446,N_7854);
nor U8086 (N_8086,N_7239,N_7689);
nor U8087 (N_8087,N_6752,N_7575);
xor U8088 (N_8088,N_7504,N_7039);
xnor U8089 (N_8089,N_6550,N_7702);
and U8090 (N_8090,N_7070,N_6888);
nand U8091 (N_8091,N_7144,N_6198);
or U8092 (N_8092,N_6788,N_7016);
or U8093 (N_8093,N_7036,N_6994);
or U8094 (N_8094,N_6689,N_7440);
xor U8095 (N_8095,N_6297,N_6171);
or U8096 (N_8096,N_7173,N_6923);
nand U8097 (N_8097,N_6218,N_7008);
nand U8098 (N_8098,N_6675,N_7732);
xnor U8099 (N_8099,N_6141,N_7873);
nand U8100 (N_8100,N_7069,N_6624);
and U8101 (N_8101,N_6424,N_7222);
xor U8102 (N_8102,N_6820,N_6960);
xor U8103 (N_8103,N_7204,N_6604);
or U8104 (N_8104,N_7355,N_7117);
or U8105 (N_8105,N_7097,N_6420);
nand U8106 (N_8106,N_6771,N_6028);
nor U8107 (N_8107,N_6165,N_7275);
nand U8108 (N_8108,N_6017,N_6793);
nand U8109 (N_8109,N_6959,N_7838);
nand U8110 (N_8110,N_7100,N_7935);
nor U8111 (N_8111,N_7075,N_7522);
nor U8112 (N_8112,N_6731,N_6288);
and U8113 (N_8113,N_7687,N_6502);
xnor U8114 (N_8114,N_7823,N_6491);
or U8115 (N_8115,N_7205,N_7770);
and U8116 (N_8116,N_6678,N_6568);
or U8117 (N_8117,N_6561,N_7174);
nand U8118 (N_8118,N_6166,N_7178);
nand U8119 (N_8119,N_7342,N_7640);
nor U8120 (N_8120,N_7487,N_7852);
nor U8121 (N_8121,N_6695,N_7666);
nor U8122 (N_8122,N_6132,N_7395);
and U8123 (N_8123,N_6975,N_7872);
nor U8124 (N_8124,N_6956,N_6630);
nand U8125 (N_8125,N_7169,N_6749);
nor U8126 (N_8126,N_6546,N_7903);
nand U8127 (N_8127,N_6918,N_7082);
xnor U8128 (N_8128,N_7649,N_7664);
or U8129 (N_8129,N_7399,N_6510);
nand U8130 (N_8130,N_7978,N_7788);
nand U8131 (N_8131,N_7931,N_7101);
or U8132 (N_8132,N_6138,N_7871);
nor U8133 (N_8133,N_6486,N_7847);
and U8134 (N_8134,N_6230,N_7199);
nand U8135 (N_8135,N_7248,N_7570);
and U8136 (N_8136,N_7492,N_7155);
and U8137 (N_8137,N_6666,N_7374);
nand U8138 (N_8138,N_7683,N_6325);
nand U8139 (N_8139,N_7262,N_7775);
xnor U8140 (N_8140,N_7932,N_6079);
xor U8141 (N_8141,N_6043,N_6857);
xnor U8142 (N_8142,N_6511,N_7076);
nor U8143 (N_8143,N_7802,N_6643);
nor U8144 (N_8144,N_7086,N_6178);
nor U8145 (N_8145,N_6626,N_7413);
and U8146 (N_8146,N_7321,N_6992);
nand U8147 (N_8147,N_7460,N_7403);
and U8148 (N_8148,N_6006,N_6681);
nor U8149 (N_8149,N_6455,N_6445);
nor U8150 (N_8150,N_6450,N_6131);
xnor U8151 (N_8151,N_7231,N_6814);
or U8152 (N_8152,N_7712,N_6884);
or U8153 (N_8153,N_6037,N_6280);
nor U8154 (N_8154,N_6056,N_7880);
or U8155 (N_8155,N_7421,N_6914);
nor U8156 (N_8156,N_6600,N_6266);
or U8157 (N_8157,N_6562,N_7379);
nor U8158 (N_8158,N_7813,N_6860);
and U8159 (N_8159,N_6393,N_6725);
and U8160 (N_8160,N_6522,N_7739);
xor U8161 (N_8161,N_6634,N_7891);
or U8162 (N_8162,N_7799,N_7499);
nor U8163 (N_8163,N_7456,N_7895);
nand U8164 (N_8164,N_7621,N_6809);
nor U8165 (N_8165,N_6811,N_6338);
or U8166 (N_8166,N_7143,N_7138);
or U8167 (N_8167,N_7285,N_7628);
nor U8168 (N_8168,N_7373,N_7357);
and U8169 (N_8169,N_6189,N_6984);
and U8170 (N_8170,N_6777,N_7362);
nor U8171 (N_8171,N_7922,N_7962);
or U8172 (N_8172,N_7152,N_6863);
or U8173 (N_8173,N_6275,N_7639);
and U8174 (N_8174,N_6877,N_7434);
nor U8175 (N_8175,N_6194,N_6475);
xnor U8176 (N_8176,N_6874,N_6748);
xor U8177 (N_8177,N_7498,N_6770);
xor U8178 (N_8178,N_7140,N_7777);
nand U8179 (N_8179,N_6528,N_7827);
nor U8180 (N_8180,N_7583,N_7571);
nand U8181 (N_8181,N_6354,N_6532);
xor U8182 (N_8182,N_7386,N_6804);
nor U8183 (N_8183,N_6136,N_7881);
xor U8184 (N_8184,N_6517,N_7488);
nor U8185 (N_8185,N_7477,N_6925);
nor U8186 (N_8186,N_6520,N_7051);
xor U8187 (N_8187,N_7263,N_7319);
nand U8188 (N_8188,N_7072,N_6588);
or U8189 (N_8189,N_7741,N_6036);
nor U8190 (N_8190,N_6796,N_6388);
xnor U8191 (N_8191,N_7162,N_7425);
nand U8192 (N_8192,N_6876,N_6154);
and U8193 (N_8193,N_6560,N_6785);
and U8194 (N_8194,N_7506,N_7503);
or U8195 (N_8195,N_6983,N_6993);
and U8196 (N_8196,N_7315,N_7428);
xor U8197 (N_8197,N_6535,N_6063);
nand U8198 (N_8198,N_6945,N_7717);
xnor U8199 (N_8199,N_7610,N_6492);
and U8200 (N_8200,N_7682,N_7849);
and U8201 (N_8201,N_7330,N_7066);
and U8202 (N_8202,N_6436,N_7195);
nor U8203 (N_8203,N_6946,N_7731);
or U8204 (N_8204,N_6714,N_7921);
nand U8205 (N_8205,N_7298,N_7896);
nand U8206 (N_8206,N_7122,N_6677);
xor U8207 (N_8207,N_6303,N_7718);
xor U8208 (N_8208,N_7229,N_6987);
xor U8209 (N_8209,N_6069,N_7705);
or U8210 (N_8210,N_6299,N_7261);
nor U8211 (N_8211,N_7518,N_6172);
or U8212 (N_8212,N_7294,N_6214);
and U8213 (N_8213,N_6893,N_6016);
nand U8214 (N_8214,N_7366,N_7572);
and U8215 (N_8215,N_6090,N_6848);
xnor U8216 (N_8216,N_7946,N_6422);
and U8217 (N_8217,N_6781,N_7055);
and U8218 (N_8218,N_6690,N_7866);
or U8219 (N_8219,N_7040,N_7000);
and U8220 (N_8220,N_7964,N_7455);
nor U8221 (N_8221,N_6283,N_7359);
xnor U8222 (N_8222,N_6365,N_7098);
and U8223 (N_8223,N_6849,N_6301);
or U8224 (N_8224,N_7784,N_7848);
and U8225 (N_8225,N_7912,N_7508);
and U8226 (N_8226,N_7118,N_6411);
or U8227 (N_8227,N_6023,N_6187);
nand U8228 (N_8228,N_7808,N_7651);
nor U8229 (N_8229,N_6792,N_7018);
or U8230 (N_8230,N_7474,N_7451);
nor U8231 (N_8231,N_7423,N_6381);
xnor U8232 (N_8232,N_7265,N_7180);
or U8233 (N_8233,N_7585,N_7783);
nor U8234 (N_8234,N_6730,N_6227);
nand U8235 (N_8235,N_6829,N_7119);
nor U8236 (N_8236,N_6322,N_6766);
or U8237 (N_8237,N_7202,N_7120);
nor U8238 (N_8238,N_7620,N_7678);
nor U8239 (N_8239,N_6272,N_7184);
and U8240 (N_8240,N_7182,N_7314);
xor U8241 (N_8241,N_6663,N_7096);
or U8242 (N_8242,N_7532,N_7886);
nand U8243 (N_8243,N_7638,N_7674);
or U8244 (N_8244,N_6158,N_7480);
nand U8245 (N_8245,N_6025,N_7998);
nand U8246 (N_8246,N_7052,N_7125);
and U8247 (N_8247,N_6534,N_7304);
nand U8248 (N_8248,N_6609,N_7590);
or U8249 (N_8249,N_6419,N_7778);
xnor U8250 (N_8250,N_6372,N_6371);
xor U8251 (N_8251,N_6533,N_7551);
and U8252 (N_8252,N_7554,N_7519);
xor U8253 (N_8253,N_7859,N_6654);
or U8254 (N_8254,N_6318,N_6489);
and U8255 (N_8255,N_6500,N_7692);
nor U8256 (N_8256,N_7020,N_7690);
or U8257 (N_8257,N_7360,N_6433);
nand U8258 (N_8258,N_7433,N_7569);
or U8259 (N_8259,N_6088,N_6536);
nand U8260 (N_8260,N_7415,N_7172);
nor U8261 (N_8261,N_7562,N_6278);
nor U8262 (N_8262,N_7787,N_7448);
and U8263 (N_8263,N_6935,N_6990);
or U8264 (N_8264,N_6182,N_6981);
nor U8265 (N_8265,N_6064,N_6578);
or U8266 (N_8266,N_7496,N_6976);
or U8267 (N_8267,N_6479,N_7221);
xor U8268 (N_8268,N_6767,N_7789);
xnor U8269 (N_8269,N_7277,N_6637);
and U8270 (N_8270,N_7232,N_7889);
xor U8271 (N_8271,N_7546,N_6773);
xor U8272 (N_8272,N_7441,N_6742);
and U8273 (N_8273,N_7206,N_6289);
nand U8274 (N_8274,N_7959,N_6692);
xnor U8275 (N_8275,N_6051,N_7376);
nor U8276 (N_8276,N_6355,N_6647);
nor U8277 (N_8277,N_6042,N_7555);
nand U8278 (N_8278,N_7971,N_6889);
nor U8279 (N_8279,N_6207,N_6705);
xor U8280 (N_8280,N_6469,N_6285);
nand U8281 (N_8281,N_6239,N_6740);
or U8282 (N_8282,N_7862,N_6940);
or U8283 (N_8283,N_7760,N_7406);
or U8284 (N_8284,N_7242,N_7807);
xor U8285 (N_8285,N_6921,N_7171);
and U8286 (N_8286,N_6062,N_6349);
or U8287 (N_8287,N_7865,N_7112);
xnor U8288 (N_8288,N_6269,N_6591);
xor U8289 (N_8289,N_6170,N_7707);
nand U8290 (N_8290,N_6800,N_6515);
xor U8291 (N_8291,N_6751,N_6686);
and U8292 (N_8292,N_7478,N_7588);
nor U8293 (N_8293,N_7986,N_7233);
xor U8294 (N_8294,N_7824,N_7464);
and U8295 (N_8295,N_6629,N_7745);
or U8296 (N_8296,N_6252,N_6423);
and U8297 (N_8297,N_6720,N_7656);
and U8298 (N_8298,N_6314,N_7219);
xor U8299 (N_8299,N_6802,N_7410);
and U8300 (N_8300,N_6570,N_6452);
xor U8301 (N_8301,N_7160,N_6222);
nor U8302 (N_8302,N_7795,N_6747);
nor U8303 (N_8303,N_7257,N_6490);
nor U8304 (N_8304,N_7836,N_6177);
nor U8305 (N_8305,N_7771,N_7673);
or U8306 (N_8306,N_7123,N_6205);
xnor U8307 (N_8307,N_6842,N_6795);
xor U8308 (N_8308,N_6547,N_6957);
nor U8309 (N_8309,N_6339,N_7200);
and U8310 (N_8310,N_7894,N_6144);
and U8311 (N_8311,N_7671,N_7370);
nor U8312 (N_8312,N_7918,N_7539);
nor U8313 (N_8313,N_7280,N_6094);
nor U8314 (N_8314,N_6460,N_6870);
or U8315 (N_8315,N_7427,N_6726);
and U8316 (N_8316,N_7906,N_6429);
and U8317 (N_8317,N_6237,N_6585);
or U8318 (N_8318,N_6631,N_7985);
or U8319 (N_8319,N_6086,N_7350);
and U8320 (N_8320,N_7127,N_6002);
and U8321 (N_8321,N_6320,N_6430);
or U8322 (N_8322,N_7194,N_6593);
nand U8323 (N_8323,N_6845,N_6179);
xnor U8324 (N_8324,N_7353,N_6223);
nand U8325 (N_8325,N_6468,N_6917);
nor U8326 (N_8326,N_7589,N_6364);
and U8327 (N_8327,N_6385,N_7038);
nand U8328 (N_8328,N_6657,N_7302);
xnor U8329 (N_8329,N_6149,N_6482);
xnor U8330 (N_8330,N_7928,N_7393);
and U8331 (N_8331,N_7438,N_6294);
nor U8332 (N_8332,N_6526,N_7104);
xnor U8333 (N_8333,N_7346,N_7801);
xor U8334 (N_8334,N_6680,N_6351);
nand U8335 (N_8335,N_7367,N_7471);
nand U8336 (N_8336,N_6234,N_7853);
and U8337 (N_8337,N_6890,N_6831);
nand U8338 (N_8338,N_6833,N_7034);
and U8339 (N_8339,N_6264,N_7927);
nand U8340 (N_8340,N_7274,N_7635);
nand U8341 (N_8341,N_7267,N_7568);
nor U8342 (N_8342,N_7384,N_7241);
nor U8343 (N_8343,N_7763,N_7452);
xnor U8344 (N_8344,N_7121,N_6108);
nand U8345 (N_8345,N_7391,N_6875);
and U8346 (N_8346,N_7974,N_6603);
xnor U8347 (N_8347,N_7181,N_7259);
nor U8348 (N_8348,N_6672,N_7412);
nand U8349 (N_8349,N_7031,N_7048);
or U8350 (N_8350,N_7574,N_6519);
xnor U8351 (N_8351,N_6193,N_7027);
xnor U8352 (N_8352,N_6022,N_7706);
or U8353 (N_8353,N_6153,N_6703);
nand U8354 (N_8354,N_6465,N_7967);
xor U8355 (N_8355,N_7402,N_7965);
or U8356 (N_8356,N_6736,N_6480);
nand U8357 (N_8357,N_7025,N_7901);
or U8358 (N_8358,N_7501,N_7805);
nor U8359 (N_8359,N_6257,N_6370);
xor U8360 (N_8360,N_6772,N_6378);
nor U8361 (N_8361,N_7913,N_6324);
nor U8362 (N_8362,N_6145,N_7026);
nand U8363 (N_8363,N_6527,N_6076);
xor U8364 (N_8364,N_6229,N_7252);
nor U8365 (N_8365,N_7614,N_6661);
and U8366 (N_8366,N_7669,N_7876);
nand U8367 (N_8367,N_7354,N_6554);
or U8368 (N_8368,N_6389,N_6464);
and U8369 (N_8369,N_7939,N_6942);
or U8370 (N_8370,N_6538,N_6871);
and U8371 (N_8371,N_6655,N_7972);
nor U8372 (N_8372,N_6854,N_7223);
or U8373 (N_8373,N_6973,N_6685);
and U8374 (N_8374,N_7916,N_7790);
nand U8375 (N_8375,N_6369,N_6516);
nand U8376 (N_8376,N_7253,N_7329);
or U8377 (N_8377,N_7786,N_7481);
nor U8378 (N_8378,N_7491,N_6007);
nand U8379 (N_8379,N_7538,N_7017);
and U8380 (N_8380,N_7715,N_6970);
nor U8381 (N_8381,N_6467,N_6844);
nand U8382 (N_8382,N_6020,N_6139);
or U8383 (N_8383,N_7653,N_6008);
nand U8384 (N_8384,N_7652,N_7850);
nor U8385 (N_8385,N_7467,N_6403);
nand U8386 (N_8386,N_7401,N_6432);
or U8387 (N_8387,N_6856,N_6117);
nor U8388 (N_8388,N_7542,N_6409);
and U8389 (N_8389,N_7168,N_7215);
and U8390 (N_8390,N_6101,N_7953);
and U8391 (N_8391,N_6531,N_6867);
nor U8392 (N_8392,N_6045,N_7544);
or U8393 (N_8393,N_6922,N_6965);
nor U8394 (N_8394,N_7502,N_6580);
nand U8395 (N_8395,N_6236,N_6072);
xnor U8396 (N_8396,N_7797,N_7989);
nor U8397 (N_8397,N_7714,N_6209);
nor U8398 (N_8398,N_7388,N_7576);
nor U8399 (N_8399,N_6225,N_6807);
nand U8400 (N_8400,N_6739,N_7214);
xnor U8401 (N_8401,N_6839,N_7166);
and U8402 (N_8402,N_7284,N_6952);
nand U8403 (N_8403,N_7540,N_6099);
xnor U8404 (N_8404,N_6951,N_6184);
and U8405 (N_8405,N_7597,N_7268);
or U8406 (N_8406,N_6316,N_7400);
xor U8407 (N_8407,N_7958,N_7820);
nor U8408 (N_8408,N_7564,N_6581);
xnor U8409 (N_8409,N_6616,N_7917);
or U8410 (N_8410,N_7197,N_6671);
xor U8411 (N_8411,N_6551,N_6114);
and U8412 (N_8412,N_6410,N_7536);
nand U8413 (N_8413,N_6553,N_6633);
nor U8414 (N_8414,N_7286,N_7382);
nor U8415 (N_8415,N_7759,N_6204);
nor U8416 (N_8416,N_6213,N_7622);
or U8417 (N_8417,N_6883,N_6451);
or U8418 (N_8418,N_6083,N_6212);
or U8419 (N_8419,N_6015,N_6815);
or U8420 (N_8420,N_7728,N_6881);
nor U8421 (N_8421,N_7884,N_7087);
and U8422 (N_8422,N_6226,N_7843);
xor U8423 (N_8423,N_6737,N_7952);
nor U8424 (N_8424,N_6050,N_6483);
xnor U8425 (N_8425,N_6812,N_6346);
nor U8426 (N_8426,N_7513,N_6886);
or U8427 (N_8427,N_7147,N_6174);
nand U8428 (N_8428,N_7577,N_7563);
or U8429 (N_8429,N_6374,N_6004);
nand U8430 (N_8430,N_6670,N_7465);
or U8431 (N_8431,N_7469,N_7511);
xnor U8432 (N_8432,N_6852,N_6038);
and U8433 (N_8433,N_7645,N_7015);
or U8434 (N_8434,N_6586,N_7115);
nand U8435 (N_8435,N_6789,N_6721);
nor U8436 (N_8436,N_7529,N_6347);
xor U8437 (N_8437,N_7819,N_7851);
and U8438 (N_8438,N_6206,N_7490);
nor U8439 (N_8439,N_7341,N_7149);
or U8440 (N_8440,N_6783,N_7968);
or U8441 (N_8441,N_7670,N_6717);
or U8442 (N_8442,N_6985,N_7212);
or U8443 (N_8443,N_7798,N_7861);
and U8444 (N_8444,N_7022,N_7293);
and U8445 (N_8445,N_7882,N_7925);
or U8446 (N_8446,N_6425,N_6133);
and U8447 (N_8447,N_6614,N_7270);
xor U8448 (N_8448,N_6120,N_7398);
nand U8449 (N_8449,N_6071,N_7631);
nand U8450 (N_8450,N_6691,N_7510);
nand U8451 (N_8451,N_7201,N_7981);
and U8452 (N_8452,N_6905,N_7459);
nor U8453 (N_8453,N_7207,N_7750);
nand U8454 (N_8454,N_6995,N_7721);
nand U8455 (N_8455,N_7716,N_6248);
and U8456 (N_8456,N_6127,N_7390);
or U8457 (N_8457,N_7407,N_6618);
nand U8458 (N_8458,N_7601,N_6825);
nand U8459 (N_8459,N_7581,N_7874);
and U8460 (N_8460,N_6011,N_7336);
xor U8461 (N_8461,N_6948,N_7537);
xor U8462 (N_8462,N_6317,N_7436);
nor U8463 (N_8463,N_7364,N_6251);
nand U8464 (N_8464,N_7713,N_7579);
and U8465 (N_8465,N_7973,N_7059);
xnor U8466 (N_8466,N_7318,N_6334);
and U8467 (N_8467,N_6112,N_7926);
nor U8468 (N_8468,N_6077,N_7081);
or U8469 (N_8469,N_7755,N_7988);
xnor U8470 (N_8470,N_6906,N_7324);
and U8471 (N_8471,N_6727,N_6010);
or U8472 (N_8472,N_6404,N_7753);
and U8473 (N_8473,N_6150,N_6862);
nand U8474 (N_8474,N_7693,N_7791);
and U8475 (N_8475,N_6950,N_6769);
or U8476 (N_8476,N_7632,N_6961);
xnor U8477 (N_8477,N_6477,N_7316);
nand U8478 (N_8478,N_6298,N_6216);
nand U8479 (N_8479,N_7634,N_6091);
and U8480 (N_8480,N_6416,N_6868);
and U8481 (N_8481,N_7032,N_7439);
nor U8482 (N_8482,N_7740,N_6494);
and U8483 (N_8483,N_7347,N_6448);
xor U8484 (N_8484,N_6653,N_7044);
xnor U8485 (N_8485,N_7722,N_7541);
and U8486 (N_8486,N_6649,N_7078);
and U8487 (N_8487,N_6024,N_7470);
or U8488 (N_8488,N_7558,N_7107);
or U8489 (N_8489,N_6897,N_6646);
nand U8490 (N_8490,N_7192,N_6111);
nor U8491 (N_8491,N_6221,N_7957);
nor U8492 (N_8492,N_6996,N_6601);
nor U8493 (N_8493,N_6032,N_7761);
or U8494 (N_8494,N_6613,N_7334);
or U8495 (N_8495,N_6947,N_6287);
nor U8496 (N_8496,N_6929,N_7785);
and U8497 (N_8497,N_6244,N_7949);
or U8498 (N_8498,N_6215,N_6955);
or U8499 (N_8499,N_6265,N_6332);
nor U8500 (N_8500,N_7338,N_6105);
or U8501 (N_8501,N_6449,N_6258);
nand U8502 (N_8502,N_6348,N_6164);
and U8503 (N_8503,N_6160,N_7028);
nand U8504 (N_8504,N_7816,N_6344);
xor U8505 (N_8505,N_6018,N_6328);
xnor U8506 (N_8506,N_7879,N_6220);
and U8507 (N_8507,N_6472,N_7942);
xnor U8508 (N_8508,N_7063,N_7997);
xor U8509 (N_8509,N_7047,N_7567);
nand U8510 (N_8510,N_7516,N_7157);
or U8511 (N_8511,N_6694,N_7767);
or U8512 (N_8512,N_7963,N_7902);
xor U8513 (N_8513,N_6060,N_6557);
nand U8514 (N_8514,N_7091,N_6119);
nor U8515 (N_8515,N_7613,N_6384);
xor U8516 (N_8516,N_6192,N_7327);
nor U8517 (N_8517,N_7530,N_7067);
nor U8518 (N_8518,N_7764,N_7604);
xor U8519 (N_8519,N_7190,N_6444);
nand U8520 (N_8520,N_7099,N_7050);
xor U8521 (N_8521,N_7396,N_6254);
and U8522 (N_8522,N_7146,N_6142);
and U8523 (N_8523,N_6697,N_6391);
or U8524 (N_8524,N_7897,N_6784);
nand U8525 (N_8525,N_7593,N_7218);
or U8526 (N_8526,N_6974,N_6949);
xnor U8527 (N_8527,N_6594,N_7776);
and U8528 (N_8528,N_6650,N_7695);
nand U8529 (N_8529,N_7420,N_6488);
nand U8530 (N_8530,N_6556,N_7266);
xnor U8531 (N_8531,N_6054,N_6247);
and U8532 (N_8532,N_6819,N_7435);
nand U8533 (N_8533,N_6201,N_7535);
nor U8534 (N_8534,N_6352,N_6967);
nand U8535 (N_8535,N_7005,N_6723);
nor U8536 (N_8536,N_6891,N_7549);
nand U8537 (N_8537,N_7408,N_6659);
nand U8538 (N_8538,N_6823,N_6092);
nor U8539 (N_8539,N_7447,N_6989);
xor U8540 (N_8540,N_6597,N_7271);
or U8541 (N_8541,N_6572,N_7203);
or U8542 (N_8542,N_7595,N_7213);
and U8543 (N_8543,N_7250,N_6402);
or U8544 (N_8544,N_6733,N_6732);
nor U8545 (N_8545,N_6760,N_6920);
and U8546 (N_8546,N_7662,N_6832);
or U8547 (N_8547,N_6173,N_6508);
nand U8548 (N_8548,N_6865,N_7062);
and U8549 (N_8549,N_7363,N_7461);
xor U8550 (N_8550,N_7994,N_7089);
or U8551 (N_8551,N_6128,N_7723);
xnor U8552 (N_8552,N_6828,N_6310);
xor U8553 (N_8553,N_6963,N_6728);
nor U8554 (N_8554,N_7148,N_6379);
nand U8555 (N_8555,N_7561,N_7860);
nand U8556 (N_8556,N_7003,N_6397);
xor U8557 (N_8557,N_6047,N_7385);
or U8558 (N_8558,N_7943,N_6798);
nor U8559 (N_8559,N_7806,N_6583);
or U8560 (N_8560,N_7686,N_6499);
nand U8561 (N_8561,N_6523,N_7264);
nor U8562 (N_8562,N_6836,N_7547);
and U8563 (N_8563,N_7887,N_7855);
or U8564 (N_8564,N_6679,N_7291);
xnor U8565 (N_8565,N_6904,N_7580);
nand U8566 (N_8566,N_6459,N_6135);
and U8567 (N_8567,N_6827,N_6255);
xor U8568 (N_8568,N_6687,N_7372);
xor U8569 (N_8569,N_6608,N_7642);
xnor U8570 (N_8570,N_6281,N_7779);
and U8571 (N_8571,N_6134,N_7983);
nand U8572 (N_8572,N_7220,N_7948);
nor U8573 (N_8573,N_6505,N_7079);
or U8574 (N_8574,N_6701,N_6276);
or U8575 (N_8575,N_6924,N_7830);
or U8576 (N_8576,N_7680,N_6121);
and U8577 (N_8577,N_6151,N_7996);
or U8578 (N_8578,N_6027,N_7371);
or U8579 (N_8579,N_6053,N_6065);
or U8580 (N_8580,N_7054,N_7703);
and U8581 (N_8581,N_6375,N_6652);
and U8582 (N_8582,N_6242,N_7616);
nand U8583 (N_8583,N_6911,N_6872);
nor U8584 (N_8584,N_6639,N_6414);
or U8585 (N_8585,N_7966,N_7211);
and U8586 (N_8586,N_6610,N_7660);
xnor U8587 (N_8587,N_6152,N_7225);
xor U8588 (N_8588,N_6907,N_6080);
or U8589 (N_8589,N_7150,N_6049);
nand U8590 (N_8590,N_6543,N_7033);
nor U8591 (N_8591,N_6110,N_6755);
nor U8592 (N_8592,N_6319,N_7061);
nor U8593 (N_8593,N_7296,N_7450);
nor U8594 (N_8594,N_7345,N_6390);
and U8595 (N_8595,N_7064,N_7483);
nor U8596 (N_8596,N_6958,N_6595);
and U8597 (N_8597,N_6758,N_7463);
or U8598 (N_8598,N_7377,N_7493);
nor U8599 (N_8599,N_7624,N_6293);
and U8600 (N_8600,N_7476,N_6787);
or U8601 (N_8601,N_6162,N_6034);
or U8602 (N_8602,N_6282,N_6715);
or U8603 (N_8603,N_7629,N_7911);
and U8604 (N_8604,N_7920,N_6873);
and U8605 (N_8605,N_6061,N_6003);
nor U8606 (N_8606,N_7186,N_6830);
or U8607 (N_8607,N_7113,N_7258);
and U8608 (N_8608,N_6582,N_7858);
nor U8609 (N_8609,N_6356,N_7701);
and U8610 (N_8610,N_6979,N_6622);
nor U8611 (N_8611,N_7584,N_7907);
or U8612 (N_8612,N_6143,N_7210);
or U8613 (N_8613,N_6458,N_7527);
xnor U8614 (N_8614,N_6599,N_7010);
and U8615 (N_8615,N_7352,N_7193);
and U8616 (N_8616,N_7982,N_6308);
nand U8617 (N_8617,N_7037,N_7725);
nand U8618 (N_8618,N_6126,N_6782);
or U8619 (N_8619,N_7600,N_6368);
or U8620 (N_8620,N_6471,N_7961);
nor U8621 (N_8621,N_7941,N_7818);
or U8622 (N_8622,N_7405,N_7295);
and U8623 (N_8623,N_6041,N_7137);
nor U8624 (N_8624,N_7606,N_7924);
and U8625 (N_8625,N_6866,N_7923);
nor U8626 (N_8626,N_6249,N_7077);
xnor U8627 (N_8627,N_6669,N_6360);
nand U8628 (N_8628,N_7608,N_6470);
nand U8629 (N_8629,N_7738,N_6291);
or U8630 (N_8630,N_7979,N_7699);
and U8631 (N_8631,N_7742,N_6190);
nand U8632 (N_8632,N_7710,N_7368);
nor U8633 (N_8633,N_6939,N_6668);
and U8634 (N_8634,N_6503,N_6466);
xor U8635 (N_8635,N_6474,N_7313);
xor U8636 (N_8636,N_6210,N_6001);
xor U8637 (N_8637,N_6926,N_7641);
or U8638 (N_8638,N_6834,N_7249);
nor U8639 (N_8639,N_7165,N_7605);
nor U8640 (N_8640,N_7424,N_6421);
xnor U8641 (N_8641,N_6046,N_7810);
xnor U8642 (N_8642,N_7747,N_6387);
and U8643 (N_8643,N_6033,N_7685);
and U8644 (N_8644,N_6456,N_7209);
nor U8645 (N_8645,N_6183,N_6159);
and U8646 (N_8646,N_7358,N_7890);
nand U8647 (N_8647,N_7073,N_7661);
xnor U8648 (N_8648,N_7247,N_7736);
xor U8649 (N_8649,N_7774,N_7418);
or U8650 (N_8650,N_7216,N_7936);
and U8651 (N_8651,N_6988,N_6245);
or U8652 (N_8652,N_7158,N_7696);
nand U8653 (N_8653,N_6169,N_6892);
xnor U8654 (N_8654,N_7893,N_6607);
or U8655 (N_8655,N_6824,N_6693);
nand U8656 (N_8656,N_7757,N_7243);
nor U8657 (N_8657,N_7512,N_6228);
xnor U8658 (N_8658,N_6665,N_7023);
and U8659 (N_8659,N_7691,N_7665);
nand U8660 (N_8660,N_6954,N_7803);
nor U8661 (N_8661,N_6337,N_6882);
xnor U8662 (N_8662,N_7161,N_6953);
xor U8663 (N_8663,N_6333,N_7733);
xor U8664 (N_8664,N_7888,N_6919);
and U8665 (N_8665,N_6292,N_6507);
xor U8666 (N_8666,N_7596,N_6084);
xnor U8667 (N_8667,N_7442,N_7289);
and U8668 (N_8668,N_7479,N_6611);
and U8669 (N_8669,N_7383,N_7758);
nor U8670 (N_8670,N_6623,N_7307);
nor U8671 (N_8671,N_6361,N_7281);
or U8672 (N_8672,N_6262,N_7904);
or U8673 (N_8673,N_7351,N_7781);
xnor U8674 (N_8674,N_7677,N_7139);
and U8675 (N_8675,N_7627,N_6899);
and U8676 (N_8676,N_6880,N_7709);
xnor U8677 (N_8677,N_6093,N_6540);
or U8678 (N_8678,N_7058,N_6790);
xnor U8679 (N_8679,N_7556,N_6321);
nor U8680 (N_8680,N_6514,N_7305);
xnor U8681 (N_8681,N_6878,N_6859);
or U8682 (N_8682,N_6074,N_7272);
or U8683 (N_8683,N_7944,N_7422);
nor U8684 (N_8684,N_6577,N_7043);
and U8685 (N_8685,N_6707,N_6200);
nor U8686 (N_8686,N_6521,N_7344);
xnor U8687 (N_8687,N_6850,N_6305);
nor U8688 (N_8688,N_7153,N_6628);
and U8689 (N_8689,N_6453,N_7323);
nor U8690 (N_8690,N_7106,N_7654);
nor U8691 (N_8691,N_7500,N_7938);
or U8692 (N_8692,N_6625,N_7011);
xor U8693 (N_8693,N_7782,N_6029);
and U8694 (N_8694,N_7533,N_6123);
and U8695 (N_8695,N_7102,N_7915);
and U8696 (N_8696,N_7484,N_7142);
nor U8697 (N_8697,N_6541,N_6735);
nand U8698 (N_8698,N_6358,N_7328);
and U8699 (N_8699,N_7131,N_7817);
and U8700 (N_8700,N_6596,N_6805);
and U8701 (N_8701,N_6605,N_7655);
or U8702 (N_8702,N_7458,N_6999);
nand U8703 (N_8703,N_7029,N_7833);
and U8704 (N_8704,N_6199,N_6304);
nand U8705 (N_8705,N_6012,N_6263);
or U8706 (N_8706,N_7255,N_6797);
or U8707 (N_8707,N_7688,N_7004);
xnor U8708 (N_8708,N_6683,N_7375);
xnor U8709 (N_8709,N_6106,N_6399);
and U8710 (N_8710,N_6619,N_6155);
nand U8711 (N_8711,N_6273,N_7780);
xor U8712 (N_8712,N_7276,N_7246);
nand U8713 (N_8713,N_7910,N_7720);
or U8714 (N_8714,N_7431,N_6224);
nand U8715 (N_8715,N_7309,N_7804);
nand U8716 (N_8716,N_7237,N_7809);
or U8717 (N_8717,N_6026,N_6779);
xor U8718 (N_8718,N_7188,N_7898);
and U8719 (N_8719,N_6780,N_6589);
xor U8720 (N_8720,N_6256,N_7980);
or U8721 (N_8721,N_7885,N_6296);
and U8722 (N_8722,N_6765,N_6821);
nor U8723 (N_8723,N_7870,N_7151);
xor U8724 (N_8724,N_6901,N_6395);
nand U8725 (N_8725,N_7657,N_7111);
xnor U8726 (N_8726,N_7103,N_7007);
xor U8727 (N_8727,N_6327,N_7337);
nand U8728 (N_8728,N_6575,N_6259);
xnor U8729 (N_8729,N_6109,N_7092);
or U8730 (N_8730,N_7411,N_6658);
nor U8731 (N_8731,N_6089,N_7905);
and U8732 (N_8732,N_6571,N_6484);
or U8733 (N_8733,N_7637,N_6070);
or U8734 (N_8734,N_6057,N_6722);
and U8735 (N_8735,N_7339,N_7462);
xnor U8736 (N_8736,N_7001,N_7553);
nor U8737 (N_8737,N_7729,N_6267);
or U8738 (N_8738,N_6813,N_7534);
and U8739 (N_8739,N_6757,N_7586);
and U8740 (N_8740,N_6427,N_7840);
xor U8741 (N_8741,N_6803,N_7129);
xnor U8742 (N_8742,N_6768,N_6738);
xor U8743 (N_8743,N_6362,N_7735);
nand U8744 (N_8744,N_7432,N_6977);
nor U8745 (N_8745,N_6635,N_6756);
and U8746 (N_8746,N_7409,N_7864);
xor U8747 (N_8747,N_6592,N_7024);
xor U8748 (N_8748,N_6481,N_6052);
and U8749 (N_8749,N_6443,N_7550);
nor U8750 (N_8750,N_6087,N_6944);
nand U8751 (N_8751,N_7602,N_6698);
nand U8752 (N_8752,N_7084,N_6392);
or U8753 (N_8753,N_6073,N_6383);
or U8754 (N_8754,N_7308,N_7466);
or U8755 (N_8755,N_6261,N_6778);
nor U8756 (N_8756,N_7227,N_7650);
xor U8757 (N_8757,N_6991,N_7468);
nor U8758 (N_8758,N_6188,N_7719);
xnor U8759 (N_8759,N_6095,N_7623);
and U8760 (N_8760,N_7083,N_6566);
nand U8761 (N_8761,N_6363,N_7299);
and U8762 (N_8762,N_6125,N_7443);
and U8763 (N_8763,N_6406,N_6806);
or U8764 (N_8764,N_7752,N_7603);
nor U8765 (N_8765,N_7672,N_7834);
or U8766 (N_8766,N_7937,N_6019);
nand U8767 (N_8767,N_6219,N_7130);
or U8768 (N_8768,N_6343,N_7947);
or U8769 (N_8769,N_7290,N_6966);
and U8770 (N_8770,N_7940,N_6962);
nand U8771 (N_8771,N_7977,N_6590);
nor U8772 (N_8772,N_6869,N_7183);
and U8773 (N_8773,N_6233,N_6367);
nor U8774 (N_8774,N_7743,N_7002);
xnor U8775 (N_8775,N_7392,N_7235);
nand U8776 (N_8776,N_6518,N_7909);
xnor U8777 (N_8777,N_7230,N_6816);
nor U8778 (N_8778,N_6196,N_6435);
or U8779 (N_8779,N_6118,N_7486);
nand U8780 (N_8780,N_6791,N_7256);
nand U8781 (N_8781,N_6931,N_7611);
and U8782 (N_8782,N_7515,N_6102);
nand U8783 (N_8783,N_7279,N_6910);
nor U8784 (N_8784,N_6059,N_6157);
nor U8785 (N_8785,N_7626,N_7071);
nor U8786 (N_8786,N_6407,N_7198);
and U8787 (N_8787,N_7663,N_6576);
xor U8788 (N_8788,N_7260,N_7381);
nand U8789 (N_8789,N_7557,N_6858);
nor U8790 (N_8790,N_6277,N_6943);
nand U8791 (N_8791,N_6801,N_6279);
or U8792 (N_8792,N_7046,N_7525);
and U8793 (N_8793,N_6377,N_6567);
nor U8794 (N_8794,N_7531,N_7124);
nor U8795 (N_8795,N_7514,N_6548);
or U8796 (N_8796,N_6300,N_6932);
nor U8797 (N_8797,N_7042,N_7236);
nand U8798 (N_8798,N_7311,N_6181);
or U8799 (N_8799,N_6615,N_6840);
nand U8800 (N_8800,N_6021,N_6167);
and U8801 (N_8801,N_7035,N_6085);
and U8802 (N_8802,N_6799,N_7141);
or U8803 (N_8803,N_7768,N_6997);
or U8804 (N_8804,N_7116,N_7074);
nand U8805 (N_8805,N_7133,N_7105);
xnor U8806 (N_8806,N_7643,N_7300);
xor U8807 (N_8807,N_6232,N_6412);
nor U8808 (N_8808,N_7414,N_7494);
and U8809 (N_8809,N_7644,N_6137);
nand U8810 (N_8810,N_6908,N_6066);
or U8811 (N_8811,N_6606,N_7065);
xnor U8812 (N_8812,N_6555,N_7587);
xnor U8813 (N_8813,N_7528,N_7019);
nor U8814 (N_8814,N_6454,N_6529);
and U8815 (N_8815,N_7793,N_7615);
nor U8816 (N_8816,N_7592,N_6718);
nor U8817 (N_8817,N_7815,N_6175);
or U8818 (N_8818,N_6473,N_7594);
xor U8819 (N_8819,N_7991,N_6326);
nand U8820 (N_8820,N_7449,N_7333);
and U8821 (N_8821,N_6838,N_6081);
and U8822 (N_8822,N_6745,N_6268);
xnor U8823 (N_8823,N_6674,N_7751);
or U8824 (N_8824,N_6243,N_7697);
nand U8825 (N_8825,N_6441,N_7273);
xnor U8826 (N_8826,N_7744,N_6711);
nand U8827 (N_8827,N_7288,N_6078);
nand U8828 (N_8828,N_6260,N_6122);
nand U8829 (N_8829,N_6719,N_6336);
nor U8830 (N_8830,N_6851,N_6913);
nor U8831 (N_8831,N_6808,N_7796);
or U8832 (N_8832,N_6253,N_7618);
or U8833 (N_8833,N_7228,N_7109);
and U8834 (N_8834,N_6900,N_6103);
and U8835 (N_8835,N_6100,N_7348);
or U8836 (N_8836,N_6916,N_7429);
xnor U8837 (N_8837,N_6729,N_6545);
or U8838 (N_8838,N_7080,N_6898);
nand U8839 (N_8839,N_6656,N_6250);
nand U8840 (N_8840,N_7730,N_6971);
and U8841 (N_8841,N_6552,N_6313);
or U8842 (N_8842,N_6794,N_6513);
or U8843 (N_8843,N_7829,N_6382);
xor U8844 (N_8844,N_7737,N_6978);
xnor U8845 (N_8845,N_7832,N_6909);
xor U8846 (N_8846,N_6284,N_6565);
and U8847 (N_8847,N_6431,N_6487);
nand U8848 (N_8848,N_6621,N_7343);
or U8849 (N_8849,N_7934,N_7599);
nor U8850 (N_8850,N_7821,N_7619);
nand U8851 (N_8851,N_7625,N_7108);
and U8852 (N_8852,N_7283,N_6295);
and U8853 (N_8853,N_6442,N_7509);
and U8854 (N_8854,N_7573,N_6644);
nor U8855 (N_8855,N_6706,N_6485);
nor U8856 (N_8856,N_6746,N_7794);
nor U8857 (N_8857,N_6645,N_6176);
nor U8858 (N_8858,N_6439,N_6195);
nor U8859 (N_8859,N_7132,N_7426);
nand U8860 (N_8860,N_6696,N_6498);
nand U8861 (N_8861,N_7762,N_7856);
xnor U8862 (N_8862,N_6039,N_6835);
or U8863 (N_8863,N_7868,N_7012);
and U8864 (N_8864,N_7548,N_7021);
and U8865 (N_8865,N_7607,N_7857);
nor U8866 (N_8866,N_6573,N_6329);
or U8867 (N_8867,N_6290,N_6903);
xnor U8868 (N_8868,N_7088,N_6040);
nand U8869 (N_8869,N_7134,N_7559);
and U8870 (N_8870,N_6107,N_6673);
or U8871 (N_8871,N_6191,N_7598);
nand U8872 (N_8872,N_7090,N_6342);
or U8873 (N_8873,N_7845,N_7482);
nand U8874 (N_8874,N_6750,N_7659);
xor U8875 (N_8875,N_6340,N_6688);
and U8876 (N_8876,N_7726,N_6902);
or U8877 (N_8877,N_7170,N_7049);
nand U8878 (N_8878,N_6764,N_7475);
nand U8879 (N_8879,N_6660,N_7507);
and U8880 (N_8880,N_6129,N_6082);
nand U8881 (N_8881,N_7404,N_7454);
and U8882 (N_8882,N_7955,N_7380);
nand U8883 (N_8883,N_6524,N_7310);
nand U8884 (N_8884,N_7749,N_7975);
xnor U8885 (N_8885,N_6307,N_6156);
or U8886 (N_8886,N_6312,N_6274);
nand U8887 (N_8887,N_7269,N_6408);
nor U8888 (N_8888,N_7837,N_7224);
nand U8889 (N_8889,N_7356,N_7056);
or U8890 (N_8890,N_7497,N_6335);
and U8891 (N_8891,N_7769,N_7668);
and U8892 (N_8892,N_6822,N_6569);
or U8893 (N_8893,N_7093,N_6712);
nor U8894 (N_8894,N_7189,N_6855);
nand U8895 (N_8895,N_7340,N_6704);
xor U8896 (N_8896,N_7312,N_6786);
or U8897 (N_8897,N_7164,N_6894);
and U8898 (N_8898,N_7754,N_7053);
or U8899 (N_8899,N_7976,N_7191);
and U8900 (N_8900,N_6847,N_6912);
nor U8901 (N_8901,N_6437,N_7041);
or U8902 (N_8902,N_7317,N_7320);
nor U8903 (N_8903,N_6400,N_7234);
xor U8904 (N_8904,N_6044,N_7582);
and U8905 (N_8905,N_7990,N_7060);
nor U8906 (N_8906,N_7136,N_7292);
or U8907 (N_8907,N_6587,N_7416);
xnor U8908 (N_8908,N_6936,N_7684);
and U8909 (N_8909,N_7301,N_7185);
or U8910 (N_8910,N_7306,N_6140);
and U8911 (N_8911,N_6632,N_7811);
xor U8912 (N_8912,N_7844,N_7419);
xor U8913 (N_8913,N_7681,N_7704);
nand U8914 (N_8914,N_6598,N_6241);
and U8915 (N_8915,N_6972,N_6197);
or U8916 (N_8916,N_6761,N_7331);
xnor U8917 (N_8917,N_6549,N_6941);
and U8918 (N_8918,N_7245,N_6405);
nor U8919 (N_8919,N_7933,N_6462);
xor U8920 (N_8920,N_7984,N_7675);
nand U8921 (N_8921,N_6345,N_7814);
and U8922 (N_8922,N_7156,N_7526);
and U8923 (N_8923,N_7999,N_7878);
or U8924 (N_8924,N_7014,N_6398);
xnor U8925 (N_8925,N_7919,N_6376);
xor U8926 (N_8926,N_7899,N_6817);
xor U8927 (N_8927,N_6186,N_6602);
nor U8928 (N_8928,N_7914,N_7326);
xor U8929 (N_8929,N_7842,N_6058);
or U8930 (N_8930,N_6708,N_6168);
nand U8931 (N_8931,N_6741,N_7251);
or U8932 (N_8932,N_6359,N_6713);
xor U8933 (N_8933,N_6286,N_7217);
or U8934 (N_8934,N_7612,N_6810);
nor U8935 (N_8935,N_6270,N_6386);
nand U8936 (N_8936,N_6501,N_6341);
nor U8937 (N_8937,N_6495,N_6302);
nor U8938 (N_8938,N_6009,N_6676);
xor U8939 (N_8939,N_6776,N_7792);
nand U8940 (N_8940,N_7877,N_6762);
or U8941 (N_8941,N_6885,N_6075);
or U8942 (N_8942,N_7960,N_6271);
and U8943 (N_8943,N_7094,N_7835);
nor U8944 (N_8944,N_6651,N_7254);
or U8945 (N_8945,N_6896,N_6366);
nand U8946 (N_8946,N_7969,N_6306);
and U8947 (N_8947,N_6203,N_7472);
xor U8948 (N_8948,N_7900,N_7951);
xnor U8949 (N_8949,N_7187,N_7159);
xnor U8950 (N_8950,N_7826,N_6682);
xnor U8951 (N_8951,N_6330,N_7297);
nor U8952 (N_8952,N_7647,N_6716);
xor U8953 (N_8953,N_6700,N_7995);
xnor U8954 (N_8954,N_7453,N_6055);
or U8955 (N_8955,N_6579,N_6509);
or U8956 (N_8956,N_6104,N_7545);
or U8957 (N_8957,N_7892,N_6775);
nand U8958 (N_8958,N_6774,N_7908);
and U8959 (N_8959,N_7445,N_7560);
nand U8960 (N_8960,N_7825,N_6710);
nand U8961 (N_8961,N_6476,N_7772);
nor U8962 (N_8962,N_7523,N_6998);
or U8963 (N_8963,N_6415,N_7667);
and U8964 (N_8964,N_7970,N_7822);
or U8965 (N_8965,N_6879,N_6968);
nor U8966 (N_8966,N_6915,N_6964);
nor U8967 (N_8967,N_6115,N_6315);
nand U8968 (N_8968,N_7679,N_7676);
xnor U8969 (N_8969,N_6240,N_6048);
and U8970 (N_8970,N_6734,N_7287);
nor U8971 (N_8971,N_7282,N_6930);
nand U8972 (N_8972,N_6537,N_7457);
nand U8973 (N_8973,N_6113,N_7954);
xnor U8974 (N_8974,N_7711,N_6843);
nor U8975 (N_8975,N_6664,N_7013);
nor U8976 (N_8976,N_7135,N_7278);
or U8977 (N_8977,N_7389,N_6559);
and U8978 (N_8978,N_6124,N_6841);
xor U8979 (N_8979,N_6148,N_6246);
and U8980 (N_8980,N_7617,N_7437);
xnor U8981 (N_8981,N_7045,N_7335);
nor U8982 (N_8982,N_6030,N_7417);
or U8983 (N_8983,N_7694,N_6744);
nor U8984 (N_8984,N_6574,N_6353);
nor U8985 (N_8985,N_7636,N_7700);
nand U8986 (N_8986,N_7154,N_6005);
xnor U8987 (N_8987,N_7867,N_6323);
xor U8988 (N_8988,N_6617,N_7987);
or U8989 (N_8989,N_7365,N_7950);
nor U8990 (N_8990,N_6709,N_7128);
and U8991 (N_8991,N_7727,N_7430);
nor U8992 (N_8992,N_6818,N_7495);
and U8993 (N_8993,N_6031,N_6504);
nor U8994 (N_8994,N_7565,N_6563);
or U8995 (N_8995,N_7167,N_7566);
nand U8996 (N_8996,N_7756,N_6743);
and U8997 (N_8997,N_6584,N_6096);
and U8998 (N_8998,N_7828,N_6530);
or U8999 (N_8999,N_6426,N_6937);
xor U9000 (N_9000,N_6090,N_7263);
or U9001 (N_9001,N_6526,N_7074);
and U9002 (N_9002,N_6575,N_7399);
and U9003 (N_9003,N_7488,N_6945);
xor U9004 (N_9004,N_7116,N_6469);
xor U9005 (N_9005,N_7378,N_7625);
nor U9006 (N_9006,N_7530,N_6398);
xor U9007 (N_9007,N_6224,N_6866);
nand U9008 (N_9008,N_7945,N_6903);
nor U9009 (N_9009,N_6461,N_7950);
xnor U9010 (N_9010,N_6824,N_6321);
xor U9011 (N_9011,N_6643,N_7702);
xnor U9012 (N_9012,N_7446,N_7360);
or U9013 (N_9013,N_6477,N_6209);
xor U9014 (N_9014,N_7654,N_6604);
nor U9015 (N_9015,N_6465,N_7540);
nor U9016 (N_9016,N_6421,N_7951);
xnor U9017 (N_9017,N_7297,N_6006);
and U9018 (N_9018,N_7217,N_7491);
or U9019 (N_9019,N_6847,N_7962);
nor U9020 (N_9020,N_6843,N_6432);
and U9021 (N_9021,N_6374,N_6490);
or U9022 (N_9022,N_7367,N_6578);
and U9023 (N_9023,N_6576,N_7546);
nor U9024 (N_9024,N_6609,N_7224);
or U9025 (N_9025,N_6250,N_6914);
and U9026 (N_9026,N_7120,N_6675);
or U9027 (N_9027,N_7450,N_7147);
or U9028 (N_9028,N_7125,N_6468);
and U9029 (N_9029,N_6046,N_7571);
or U9030 (N_9030,N_7899,N_6337);
and U9031 (N_9031,N_7825,N_7753);
nand U9032 (N_9032,N_6929,N_6064);
nand U9033 (N_9033,N_7347,N_7655);
and U9034 (N_9034,N_6529,N_6650);
and U9035 (N_9035,N_6109,N_7889);
nor U9036 (N_9036,N_7887,N_7921);
and U9037 (N_9037,N_7464,N_6198);
or U9038 (N_9038,N_7947,N_7854);
xor U9039 (N_9039,N_7075,N_6950);
nand U9040 (N_9040,N_6837,N_6339);
nand U9041 (N_9041,N_6140,N_7839);
and U9042 (N_9042,N_6674,N_6744);
nor U9043 (N_9043,N_7249,N_7182);
or U9044 (N_9044,N_7507,N_7856);
nor U9045 (N_9045,N_6549,N_7828);
or U9046 (N_9046,N_7526,N_6453);
or U9047 (N_9047,N_7022,N_7909);
nor U9048 (N_9048,N_7433,N_6958);
nand U9049 (N_9049,N_6921,N_6739);
nand U9050 (N_9050,N_6132,N_7183);
or U9051 (N_9051,N_6182,N_6313);
or U9052 (N_9052,N_7463,N_6208);
xnor U9053 (N_9053,N_6470,N_6207);
xor U9054 (N_9054,N_7100,N_6512);
or U9055 (N_9055,N_7706,N_7435);
or U9056 (N_9056,N_6708,N_7297);
xnor U9057 (N_9057,N_7789,N_7924);
and U9058 (N_9058,N_7548,N_6864);
xnor U9059 (N_9059,N_6713,N_7093);
or U9060 (N_9060,N_7749,N_7874);
nor U9061 (N_9061,N_6908,N_7150);
xnor U9062 (N_9062,N_7099,N_6106);
or U9063 (N_9063,N_6348,N_7220);
and U9064 (N_9064,N_6752,N_6248);
xnor U9065 (N_9065,N_7908,N_6357);
nand U9066 (N_9066,N_7685,N_6726);
or U9067 (N_9067,N_7302,N_6240);
xor U9068 (N_9068,N_7745,N_6240);
or U9069 (N_9069,N_7339,N_7091);
and U9070 (N_9070,N_7101,N_6823);
or U9071 (N_9071,N_7629,N_7491);
or U9072 (N_9072,N_7973,N_7721);
nand U9073 (N_9073,N_6205,N_7342);
nor U9074 (N_9074,N_6118,N_7894);
nand U9075 (N_9075,N_6489,N_7172);
or U9076 (N_9076,N_6595,N_6078);
and U9077 (N_9077,N_6097,N_6457);
nand U9078 (N_9078,N_7890,N_7818);
nor U9079 (N_9079,N_6179,N_7123);
nor U9080 (N_9080,N_6291,N_7118);
nand U9081 (N_9081,N_7351,N_6130);
nand U9082 (N_9082,N_7083,N_6383);
xor U9083 (N_9083,N_6409,N_6965);
nor U9084 (N_9084,N_6425,N_6393);
or U9085 (N_9085,N_6586,N_7744);
xnor U9086 (N_9086,N_7933,N_6722);
and U9087 (N_9087,N_7167,N_7999);
xor U9088 (N_9088,N_7729,N_6098);
xnor U9089 (N_9089,N_6216,N_7607);
or U9090 (N_9090,N_6601,N_6111);
xor U9091 (N_9091,N_7223,N_6672);
nor U9092 (N_9092,N_6416,N_6547);
nor U9093 (N_9093,N_6157,N_7912);
nor U9094 (N_9094,N_6055,N_6000);
xnor U9095 (N_9095,N_6595,N_6453);
and U9096 (N_9096,N_6443,N_6480);
nor U9097 (N_9097,N_7621,N_7415);
or U9098 (N_9098,N_6898,N_6002);
nor U9099 (N_9099,N_7072,N_6047);
and U9100 (N_9100,N_6636,N_7522);
or U9101 (N_9101,N_6586,N_7336);
or U9102 (N_9102,N_7457,N_6572);
xnor U9103 (N_9103,N_6819,N_6893);
and U9104 (N_9104,N_7481,N_7168);
nand U9105 (N_9105,N_7866,N_7450);
or U9106 (N_9106,N_6839,N_7924);
and U9107 (N_9107,N_7633,N_7410);
nor U9108 (N_9108,N_6810,N_6823);
nand U9109 (N_9109,N_6917,N_6276);
nand U9110 (N_9110,N_7444,N_6336);
or U9111 (N_9111,N_7871,N_6744);
nor U9112 (N_9112,N_6384,N_6084);
xnor U9113 (N_9113,N_7984,N_7657);
xor U9114 (N_9114,N_6860,N_6539);
and U9115 (N_9115,N_6585,N_6549);
nor U9116 (N_9116,N_7399,N_6083);
and U9117 (N_9117,N_6709,N_7185);
or U9118 (N_9118,N_6004,N_7351);
or U9119 (N_9119,N_6749,N_6284);
xor U9120 (N_9120,N_6962,N_6932);
nor U9121 (N_9121,N_6374,N_6732);
nor U9122 (N_9122,N_6746,N_6444);
or U9123 (N_9123,N_7800,N_6110);
nand U9124 (N_9124,N_6319,N_7546);
xnor U9125 (N_9125,N_7169,N_6894);
or U9126 (N_9126,N_7411,N_7338);
nor U9127 (N_9127,N_6817,N_6444);
and U9128 (N_9128,N_6704,N_6791);
nand U9129 (N_9129,N_7496,N_6021);
and U9130 (N_9130,N_6921,N_6725);
and U9131 (N_9131,N_6723,N_6592);
and U9132 (N_9132,N_6670,N_6298);
or U9133 (N_9133,N_7413,N_7114);
nor U9134 (N_9134,N_6129,N_6501);
or U9135 (N_9135,N_7142,N_6420);
or U9136 (N_9136,N_7077,N_6449);
xor U9137 (N_9137,N_7893,N_7270);
xor U9138 (N_9138,N_7645,N_7810);
or U9139 (N_9139,N_6970,N_6964);
and U9140 (N_9140,N_7670,N_7319);
nor U9141 (N_9141,N_7623,N_7442);
xor U9142 (N_9142,N_7494,N_6788);
and U9143 (N_9143,N_6787,N_6589);
xnor U9144 (N_9144,N_6107,N_7924);
nand U9145 (N_9145,N_7773,N_7021);
nand U9146 (N_9146,N_7689,N_7969);
nand U9147 (N_9147,N_6447,N_7621);
xnor U9148 (N_9148,N_7782,N_7039);
nor U9149 (N_9149,N_7092,N_6694);
and U9150 (N_9150,N_7878,N_7665);
nand U9151 (N_9151,N_7723,N_7009);
and U9152 (N_9152,N_7299,N_6544);
xor U9153 (N_9153,N_7715,N_6156);
and U9154 (N_9154,N_7259,N_7477);
nand U9155 (N_9155,N_6849,N_6685);
nor U9156 (N_9156,N_6449,N_7721);
or U9157 (N_9157,N_6862,N_7717);
and U9158 (N_9158,N_6224,N_6611);
or U9159 (N_9159,N_6158,N_7052);
nand U9160 (N_9160,N_7269,N_6571);
or U9161 (N_9161,N_6291,N_6336);
and U9162 (N_9162,N_6755,N_6943);
or U9163 (N_9163,N_7188,N_7461);
nand U9164 (N_9164,N_7149,N_7620);
and U9165 (N_9165,N_7693,N_6534);
and U9166 (N_9166,N_6193,N_6891);
xnor U9167 (N_9167,N_7303,N_7011);
nor U9168 (N_9168,N_7301,N_6709);
nand U9169 (N_9169,N_6845,N_7542);
xnor U9170 (N_9170,N_7521,N_6866);
nor U9171 (N_9171,N_7531,N_6634);
xnor U9172 (N_9172,N_7744,N_6769);
and U9173 (N_9173,N_7798,N_7836);
xor U9174 (N_9174,N_6644,N_7580);
nor U9175 (N_9175,N_7796,N_6436);
nand U9176 (N_9176,N_6443,N_7836);
and U9177 (N_9177,N_7992,N_6859);
xnor U9178 (N_9178,N_6242,N_6467);
or U9179 (N_9179,N_7134,N_7465);
nor U9180 (N_9180,N_6527,N_7089);
nand U9181 (N_9181,N_6100,N_7568);
nor U9182 (N_9182,N_7771,N_7495);
or U9183 (N_9183,N_6817,N_6853);
nand U9184 (N_9184,N_6944,N_6754);
nand U9185 (N_9185,N_6384,N_7328);
and U9186 (N_9186,N_7391,N_7795);
or U9187 (N_9187,N_7246,N_6032);
or U9188 (N_9188,N_6007,N_6574);
or U9189 (N_9189,N_7868,N_6466);
nand U9190 (N_9190,N_6568,N_7167);
xnor U9191 (N_9191,N_6366,N_7653);
nand U9192 (N_9192,N_6787,N_6844);
xnor U9193 (N_9193,N_7482,N_6907);
xnor U9194 (N_9194,N_6853,N_7297);
nand U9195 (N_9195,N_6021,N_6046);
xnor U9196 (N_9196,N_6027,N_6850);
xor U9197 (N_9197,N_7653,N_7453);
xnor U9198 (N_9198,N_6227,N_7162);
nand U9199 (N_9199,N_7102,N_7683);
or U9200 (N_9200,N_7327,N_6797);
nand U9201 (N_9201,N_6436,N_7559);
nor U9202 (N_9202,N_6595,N_6280);
nand U9203 (N_9203,N_6747,N_7905);
and U9204 (N_9204,N_7612,N_6997);
or U9205 (N_9205,N_7543,N_7141);
nor U9206 (N_9206,N_7788,N_7127);
xnor U9207 (N_9207,N_6938,N_6824);
or U9208 (N_9208,N_7700,N_6190);
xor U9209 (N_9209,N_7657,N_6593);
nor U9210 (N_9210,N_7749,N_6661);
and U9211 (N_9211,N_6783,N_7089);
xnor U9212 (N_9212,N_6510,N_6955);
and U9213 (N_9213,N_7657,N_7104);
nand U9214 (N_9214,N_6026,N_7519);
nor U9215 (N_9215,N_6245,N_7039);
and U9216 (N_9216,N_6264,N_6948);
and U9217 (N_9217,N_6445,N_7384);
or U9218 (N_9218,N_7514,N_6751);
or U9219 (N_9219,N_6618,N_7714);
nor U9220 (N_9220,N_7889,N_7547);
nor U9221 (N_9221,N_6452,N_7418);
xor U9222 (N_9222,N_6811,N_6678);
nor U9223 (N_9223,N_6188,N_7703);
xor U9224 (N_9224,N_7135,N_6142);
nand U9225 (N_9225,N_6977,N_7959);
nor U9226 (N_9226,N_6299,N_6560);
and U9227 (N_9227,N_6756,N_6291);
or U9228 (N_9228,N_7255,N_7195);
or U9229 (N_9229,N_6815,N_6211);
or U9230 (N_9230,N_7447,N_7268);
or U9231 (N_9231,N_6911,N_7095);
nand U9232 (N_9232,N_6540,N_6127);
nor U9233 (N_9233,N_6958,N_6707);
xor U9234 (N_9234,N_6506,N_7425);
or U9235 (N_9235,N_7379,N_7720);
or U9236 (N_9236,N_6399,N_7731);
nand U9237 (N_9237,N_6569,N_7564);
nand U9238 (N_9238,N_6157,N_7844);
or U9239 (N_9239,N_6715,N_6825);
or U9240 (N_9240,N_7689,N_7439);
nor U9241 (N_9241,N_7847,N_6512);
xnor U9242 (N_9242,N_7676,N_6689);
xor U9243 (N_9243,N_7486,N_6889);
nand U9244 (N_9244,N_6340,N_6018);
nor U9245 (N_9245,N_7767,N_7890);
xor U9246 (N_9246,N_6798,N_7933);
nand U9247 (N_9247,N_7435,N_6029);
or U9248 (N_9248,N_7252,N_6309);
xor U9249 (N_9249,N_6305,N_7981);
and U9250 (N_9250,N_7737,N_6613);
xnor U9251 (N_9251,N_6696,N_6220);
or U9252 (N_9252,N_7162,N_6407);
nor U9253 (N_9253,N_7566,N_7974);
nand U9254 (N_9254,N_7950,N_7607);
xnor U9255 (N_9255,N_6579,N_6163);
and U9256 (N_9256,N_7222,N_6212);
or U9257 (N_9257,N_7528,N_6860);
nand U9258 (N_9258,N_6527,N_6747);
nor U9259 (N_9259,N_7607,N_6506);
nor U9260 (N_9260,N_7563,N_7290);
nor U9261 (N_9261,N_6585,N_7849);
nor U9262 (N_9262,N_7350,N_6553);
xor U9263 (N_9263,N_6496,N_6828);
xor U9264 (N_9264,N_7191,N_6179);
nor U9265 (N_9265,N_7755,N_7468);
xor U9266 (N_9266,N_6127,N_6922);
xnor U9267 (N_9267,N_7585,N_6148);
or U9268 (N_9268,N_7164,N_6076);
nor U9269 (N_9269,N_6304,N_6645);
or U9270 (N_9270,N_7051,N_6304);
and U9271 (N_9271,N_7792,N_7852);
or U9272 (N_9272,N_6374,N_6495);
nor U9273 (N_9273,N_7082,N_6454);
xnor U9274 (N_9274,N_6002,N_6712);
xor U9275 (N_9275,N_7132,N_7514);
or U9276 (N_9276,N_7711,N_6531);
nor U9277 (N_9277,N_6655,N_7596);
xnor U9278 (N_9278,N_7484,N_7033);
xor U9279 (N_9279,N_6849,N_7164);
nor U9280 (N_9280,N_7776,N_7714);
and U9281 (N_9281,N_7943,N_7071);
nor U9282 (N_9282,N_7456,N_7916);
nand U9283 (N_9283,N_6254,N_6001);
nor U9284 (N_9284,N_6650,N_7492);
or U9285 (N_9285,N_6929,N_7849);
and U9286 (N_9286,N_6822,N_7466);
and U9287 (N_9287,N_6027,N_6593);
xor U9288 (N_9288,N_6678,N_7658);
xor U9289 (N_9289,N_6052,N_6894);
nor U9290 (N_9290,N_6751,N_6906);
xnor U9291 (N_9291,N_6647,N_7063);
nand U9292 (N_9292,N_7122,N_6007);
or U9293 (N_9293,N_7903,N_7834);
nand U9294 (N_9294,N_6084,N_6812);
and U9295 (N_9295,N_7303,N_6054);
and U9296 (N_9296,N_6290,N_7878);
nand U9297 (N_9297,N_7483,N_6419);
xor U9298 (N_9298,N_6685,N_6029);
or U9299 (N_9299,N_7898,N_6920);
nand U9300 (N_9300,N_7712,N_6651);
and U9301 (N_9301,N_7771,N_6753);
nand U9302 (N_9302,N_7627,N_6294);
nand U9303 (N_9303,N_7128,N_7710);
nor U9304 (N_9304,N_6109,N_7488);
or U9305 (N_9305,N_6637,N_7719);
xnor U9306 (N_9306,N_6646,N_6691);
xnor U9307 (N_9307,N_7480,N_6841);
nand U9308 (N_9308,N_6371,N_7870);
nand U9309 (N_9309,N_7528,N_7159);
nand U9310 (N_9310,N_6532,N_6000);
xor U9311 (N_9311,N_6398,N_7184);
xor U9312 (N_9312,N_6079,N_7176);
xnor U9313 (N_9313,N_6869,N_7638);
or U9314 (N_9314,N_7737,N_6194);
nand U9315 (N_9315,N_6230,N_6258);
or U9316 (N_9316,N_6910,N_7842);
and U9317 (N_9317,N_6282,N_7006);
nor U9318 (N_9318,N_6568,N_7806);
or U9319 (N_9319,N_6759,N_6015);
and U9320 (N_9320,N_6923,N_6015);
or U9321 (N_9321,N_7102,N_6002);
nand U9322 (N_9322,N_7689,N_6308);
and U9323 (N_9323,N_6857,N_7279);
nand U9324 (N_9324,N_6317,N_6978);
nand U9325 (N_9325,N_7254,N_6097);
or U9326 (N_9326,N_6011,N_7197);
or U9327 (N_9327,N_6089,N_7350);
xor U9328 (N_9328,N_6160,N_6225);
xnor U9329 (N_9329,N_6994,N_7359);
nor U9330 (N_9330,N_7618,N_6488);
nand U9331 (N_9331,N_7012,N_6696);
xor U9332 (N_9332,N_6818,N_6846);
and U9333 (N_9333,N_6116,N_6894);
nand U9334 (N_9334,N_6415,N_6383);
xor U9335 (N_9335,N_6945,N_6187);
nor U9336 (N_9336,N_7037,N_6542);
xnor U9337 (N_9337,N_7883,N_6107);
and U9338 (N_9338,N_7684,N_6648);
xnor U9339 (N_9339,N_6225,N_6421);
nand U9340 (N_9340,N_7652,N_7862);
nor U9341 (N_9341,N_6826,N_7427);
or U9342 (N_9342,N_7938,N_7016);
and U9343 (N_9343,N_7798,N_7767);
nor U9344 (N_9344,N_7623,N_7212);
xnor U9345 (N_9345,N_7912,N_6220);
or U9346 (N_9346,N_6501,N_6689);
and U9347 (N_9347,N_6001,N_7602);
and U9348 (N_9348,N_6289,N_6944);
or U9349 (N_9349,N_6867,N_6237);
nor U9350 (N_9350,N_6840,N_7858);
nor U9351 (N_9351,N_6182,N_6604);
nand U9352 (N_9352,N_7387,N_6671);
and U9353 (N_9353,N_6069,N_7977);
and U9354 (N_9354,N_7457,N_7035);
and U9355 (N_9355,N_6988,N_7276);
and U9356 (N_9356,N_6667,N_6871);
or U9357 (N_9357,N_7091,N_7718);
or U9358 (N_9358,N_7782,N_7686);
nor U9359 (N_9359,N_6989,N_6228);
xnor U9360 (N_9360,N_7561,N_6253);
and U9361 (N_9361,N_6950,N_6226);
and U9362 (N_9362,N_6634,N_6653);
nand U9363 (N_9363,N_6408,N_6534);
nor U9364 (N_9364,N_6563,N_6115);
or U9365 (N_9365,N_6879,N_7032);
nor U9366 (N_9366,N_7517,N_6304);
or U9367 (N_9367,N_7260,N_7551);
nor U9368 (N_9368,N_7250,N_6657);
and U9369 (N_9369,N_6429,N_7272);
nor U9370 (N_9370,N_7416,N_6088);
xnor U9371 (N_9371,N_6293,N_7683);
or U9372 (N_9372,N_6323,N_7583);
xnor U9373 (N_9373,N_6171,N_7231);
nor U9374 (N_9374,N_7450,N_7759);
nand U9375 (N_9375,N_6489,N_7236);
nor U9376 (N_9376,N_7860,N_7913);
or U9377 (N_9377,N_6113,N_7287);
nor U9378 (N_9378,N_7588,N_7679);
or U9379 (N_9379,N_7722,N_7485);
or U9380 (N_9380,N_7187,N_6542);
nor U9381 (N_9381,N_7568,N_7641);
and U9382 (N_9382,N_6989,N_6725);
nand U9383 (N_9383,N_6847,N_6477);
xor U9384 (N_9384,N_6421,N_7522);
nand U9385 (N_9385,N_6515,N_6355);
nor U9386 (N_9386,N_7640,N_6184);
nand U9387 (N_9387,N_6033,N_6542);
xnor U9388 (N_9388,N_6539,N_7237);
xor U9389 (N_9389,N_6482,N_6940);
nand U9390 (N_9390,N_7308,N_6914);
or U9391 (N_9391,N_6684,N_6083);
nor U9392 (N_9392,N_6033,N_6780);
nand U9393 (N_9393,N_6788,N_7491);
nand U9394 (N_9394,N_6593,N_7208);
or U9395 (N_9395,N_7280,N_7553);
nand U9396 (N_9396,N_7518,N_6441);
xor U9397 (N_9397,N_6072,N_6572);
or U9398 (N_9398,N_7940,N_7449);
nor U9399 (N_9399,N_6176,N_6599);
and U9400 (N_9400,N_6919,N_7880);
nand U9401 (N_9401,N_7993,N_7708);
xor U9402 (N_9402,N_7534,N_7760);
nand U9403 (N_9403,N_7768,N_7538);
and U9404 (N_9404,N_7727,N_7977);
and U9405 (N_9405,N_7189,N_7290);
xnor U9406 (N_9406,N_6190,N_7402);
or U9407 (N_9407,N_6508,N_7980);
xor U9408 (N_9408,N_7921,N_6302);
nand U9409 (N_9409,N_6758,N_7577);
nand U9410 (N_9410,N_7169,N_7932);
nor U9411 (N_9411,N_7365,N_6640);
xnor U9412 (N_9412,N_6564,N_7338);
xor U9413 (N_9413,N_7232,N_6211);
xor U9414 (N_9414,N_6518,N_7274);
or U9415 (N_9415,N_7082,N_6999);
and U9416 (N_9416,N_6373,N_6363);
and U9417 (N_9417,N_6092,N_7907);
nand U9418 (N_9418,N_7940,N_6013);
and U9419 (N_9419,N_6258,N_6401);
nor U9420 (N_9420,N_6529,N_7447);
nor U9421 (N_9421,N_6346,N_6113);
xor U9422 (N_9422,N_6843,N_6068);
and U9423 (N_9423,N_7022,N_7448);
nand U9424 (N_9424,N_7409,N_7246);
and U9425 (N_9425,N_6144,N_7264);
nor U9426 (N_9426,N_6125,N_7610);
or U9427 (N_9427,N_6902,N_6317);
nor U9428 (N_9428,N_6476,N_6583);
nand U9429 (N_9429,N_6962,N_7941);
nand U9430 (N_9430,N_7698,N_6555);
nor U9431 (N_9431,N_6810,N_7412);
nand U9432 (N_9432,N_7745,N_6559);
or U9433 (N_9433,N_6575,N_6284);
nor U9434 (N_9434,N_6681,N_7191);
and U9435 (N_9435,N_6860,N_7393);
or U9436 (N_9436,N_6196,N_7724);
and U9437 (N_9437,N_7161,N_7706);
xor U9438 (N_9438,N_6096,N_7685);
and U9439 (N_9439,N_6187,N_7364);
and U9440 (N_9440,N_6904,N_7180);
nor U9441 (N_9441,N_7769,N_6577);
nand U9442 (N_9442,N_6650,N_7973);
nor U9443 (N_9443,N_7687,N_6410);
and U9444 (N_9444,N_6464,N_6559);
xor U9445 (N_9445,N_7638,N_7231);
nor U9446 (N_9446,N_6735,N_6584);
xor U9447 (N_9447,N_6864,N_6604);
xnor U9448 (N_9448,N_6357,N_7322);
and U9449 (N_9449,N_7419,N_7931);
nor U9450 (N_9450,N_6334,N_6928);
or U9451 (N_9451,N_7688,N_6661);
nor U9452 (N_9452,N_6046,N_6671);
and U9453 (N_9453,N_6348,N_7428);
or U9454 (N_9454,N_6091,N_7497);
nor U9455 (N_9455,N_6194,N_6401);
and U9456 (N_9456,N_7470,N_7939);
nor U9457 (N_9457,N_6647,N_6813);
xor U9458 (N_9458,N_7981,N_6925);
nand U9459 (N_9459,N_6460,N_7971);
or U9460 (N_9460,N_7029,N_7767);
and U9461 (N_9461,N_6943,N_7934);
and U9462 (N_9462,N_6301,N_6350);
xor U9463 (N_9463,N_7440,N_7503);
nor U9464 (N_9464,N_7591,N_7644);
and U9465 (N_9465,N_6920,N_7011);
and U9466 (N_9466,N_7801,N_7879);
xor U9467 (N_9467,N_7277,N_6760);
or U9468 (N_9468,N_7394,N_6690);
xnor U9469 (N_9469,N_7100,N_6851);
or U9470 (N_9470,N_7004,N_7166);
and U9471 (N_9471,N_6909,N_7756);
nor U9472 (N_9472,N_6890,N_6409);
nand U9473 (N_9473,N_7363,N_6772);
nand U9474 (N_9474,N_6056,N_6943);
nand U9475 (N_9475,N_6795,N_6189);
and U9476 (N_9476,N_6982,N_7783);
xnor U9477 (N_9477,N_7418,N_6160);
or U9478 (N_9478,N_6712,N_7830);
and U9479 (N_9479,N_6706,N_7620);
and U9480 (N_9480,N_6141,N_7322);
nand U9481 (N_9481,N_7615,N_6901);
nor U9482 (N_9482,N_7070,N_7458);
and U9483 (N_9483,N_7699,N_7576);
or U9484 (N_9484,N_6503,N_6462);
and U9485 (N_9485,N_7278,N_7926);
and U9486 (N_9486,N_6207,N_7931);
nand U9487 (N_9487,N_7072,N_6902);
xnor U9488 (N_9488,N_6974,N_7375);
nand U9489 (N_9489,N_7512,N_7537);
nor U9490 (N_9490,N_7062,N_7515);
xor U9491 (N_9491,N_7679,N_6074);
or U9492 (N_9492,N_7144,N_7938);
nand U9493 (N_9493,N_7225,N_7849);
and U9494 (N_9494,N_7613,N_7968);
or U9495 (N_9495,N_6357,N_6946);
or U9496 (N_9496,N_6173,N_7930);
xnor U9497 (N_9497,N_6792,N_6109);
nor U9498 (N_9498,N_6940,N_7447);
nand U9499 (N_9499,N_6993,N_7199);
nand U9500 (N_9500,N_7628,N_7170);
nand U9501 (N_9501,N_6337,N_6806);
and U9502 (N_9502,N_6606,N_6070);
xnor U9503 (N_9503,N_7280,N_7253);
nand U9504 (N_9504,N_7580,N_6532);
nor U9505 (N_9505,N_7121,N_6231);
xnor U9506 (N_9506,N_7830,N_6699);
nor U9507 (N_9507,N_6451,N_6162);
or U9508 (N_9508,N_7324,N_7622);
nand U9509 (N_9509,N_6065,N_7241);
xor U9510 (N_9510,N_6085,N_6053);
and U9511 (N_9511,N_6981,N_6355);
and U9512 (N_9512,N_6927,N_6607);
and U9513 (N_9513,N_7031,N_7328);
or U9514 (N_9514,N_6805,N_7283);
nor U9515 (N_9515,N_6754,N_6539);
xnor U9516 (N_9516,N_7499,N_7740);
xor U9517 (N_9517,N_7326,N_7247);
and U9518 (N_9518,N_7916,N_7172);
or U9519 (N_9519,N_6030,N_6394);
or U9520 (N_9520,N_6311,N_7264);
xor U9521 (N_9521,N_6338,N_7570);
nand U9522 (N_9522,N_6914,N_7514);
nor U9523 (N_9523,N_7648,N_6787);
or U9524 (N_9524,N_6512,N_6813);
or U9525 (N_9525,N_7434,N_6014);
nor U9526 (N_9526,N_7349,N_7844);
nor U9527 (N_9527,N_6743,N_7725);
xor U9528 (N_9528,N_6911,N_7163);
nand U9529 (N_9529,N_7859,N_6783);
and U9530 (N_9530,N_7359,N_6985);
nor U9531 (N_9531,N_6322,N_6488);
nor U9532 (N_9532,N_6326,N_7280);
nand U9533 (N_9533,N_6613,N_7049);
or U9534 (N_9534,N_6186,N_6969);
nor U9535 (N_9535,N_7236,N_6259);
or U9536 (N_9536,N_7682,N_6363);
nand U9537 (N_9537,N_7059,N_6725);
and U9538 (N_9538,N_7114,N_6052);
nor U9539 (N_9539,N_7947,N_6710);
xor U9540 (N_9540,N_6697,N_7555);
or U9541 (N_9541,N_6587,N_6777);
nor U9542 (N_9542,N_7902,N_7873);
nand U9543 (N_9543,N_6143,N_6561);
nand U9544 (N_9544,N_6939,N_6810);
or U9545 (N_9545,N_7151,N_7207);
xor U9546 (N_9546,N_6593,N_7184);
nor U9547 (N_9547,N_6474,N_6657);
or U9548 (N_9548,N_7128,N_7465);
nand U9549 (N_9549,N_6092,N_7033);
xor U9550 (N_9550,N_7411,N_7686);
xnor U9551 (N_9551,N_6412,N_6641);
and U9552 (N_9552,N_6341,N_7962);
nand U9553 (N_9553,N_6558,N_7864);
or U9554 (N_9554,N_7361,N_6743);
and U9555 (N_9555,N_7427,N_7417);
nand U9556 (N_9556,N_7866,N_7392);
xnor U9557 (N_9557,N_6775,N_7464);
nor U9558 (N_9558,N_6791,N_6464);
xnor U9559 (N_9559,N_6136,N_6245);
or U9560 (N_9560,N_6217,N_7401);
or U9561 (N_9561,N_7020,N_7566);
xnor U9562 (N_9562,N_6673,N_7104);
xnor U9563 (N_9563,N_6003,N_7377);
and U9564 (N_9564,N_6315,N_6418);
or U9565 (N_9565,N_7968,N_6744);
and U9566 (N_9566,N_6430,N_6578);
xnor U9567 (N_9567,N_7411,N_6468);
nand U9568 (N_9568,N_6893,N_6033);
and U9569 (N_9569,N_6261,N_6065);
and U9570 (N_9570,N_6245,N_6347);
or U9571 (N_9571,N_7499,N_7625);
or U9572 (N_9572,N_7619,N_7024);
xor U9573 (N_9573,N_6127,N_6646);
or U9574 (N_9574,N_7393,N_7367);
xor U9575 (N_9575,N_6830,N_6747);
or U9576 (N_9576,N_6711,N_6459);
and U9577 (N_9577,N_6776,N_6262);
or U9578 (N_9578,N_7407,N_6724);
and U9579 (N_9579,N_7418,N_6541);
xnor U9580 (N_9580,N_6211,N_6415);
and U9581 (N_9581,N_6720,N_6891);
xnor U9582 (N_9582,N_6086,N_6591);
or U9583 (N_9583,N_6910,N_6526);
or U9584 (N_9584,N_6582,N_6419);
nand U9585 (N_9585,N_6437,N_7545);
or U9586 (N_9586,N_6984,N_6737);
or U9587 (N_9587,N_7180,N_7428);
or U9588 (N_9588,N_7046,N_7075);
and U9589 (N_9589,N_7092,N_6024);
and U9590 (N_9590,N_6083,N_6115);
or U9591 (N_9591,N_7246,N_6737);
and U9592 (N_9592,N_6975,N_6252);
or U9593 (N_9593,N_7049,N_7731);
or U9594 (N_9594,N_7329,N_7519);
and U9595 (N_9595,N_6551,N_7436);
and U9596 (N_9596,N_6650,N_6088);
xnor U9597 (N_9597,N_7590,N_6628);
and U9598 (N_9598,N_6065,N_6820);
nand U9599 (N_9599,N_7643,N_6733);
or U9600 (N_9600,N_6216,N_6392);
xor U9601 (N_9601,N_6012,N_7947);
xor U9602 (N_9602,N_6277,N_7488);
xor U9603 (N_9603,N_7476,N_6041);
and U9604 (N_9604,N_7534,N_7037);
nand U9605 (N_9605,N_7554,N_6818);
xnor U9606 (N_9606,N_7002,N_7969);
nand U9607 (N_9607,N_6377,N_6688);
and U9608 (N_9608,N_6230,N_6954);
xor U9609 (N_9609,N_6924,N_6507);
nor U9610 (N_9610,N_7973,N_7604);
or U9611 (N_9611,N_6270,N_7225);
or U9612 (N_9612,N_6740,N_6398);
and U9613 (N_9613,N_6247,N_7469);
nor U9614 (N_9614,N_6823,N_7844);
nand U9615 (N_9615,N_6489,N_6854);
nor U9616 (N_9616,N_7427,N_6576);
nor U9617 (N_9617,N_7392,N_7502);
nand U9618 (N_9618,N_6081,N_6653);
and U9619 (N_9619,N_7153,N_6916);
nand U9620 (N_9620,N_6859,N_7113);
or U9621 (N_9621,N_7290,N_7749);
and U9622 (N_9622,N_7445,N_7013);
nor U9623 (N_9623,N_6001,N_7069);
nor U9624 (N_9624,N_7926,N_6474);
and U9625 (N_9625,N_6223,N_7212);
or U9626 (N_9626,N_6939,N_7886);
nand U9627 (N_9627,N_7174,N_7818);
nor U9628 (N_9628,N_6914,N_6737);
nand U9629 (N_9629,N_6186,N_7122);
nand U9630 (N_9630,N_6448,N_6956);
nand U9631 (N_9631,N_7457,N_6221);
and U9632 (N_9632,N_6664,N_6058);
nor U9633 (N_9633,N_6906,N_6839);
or U9634 (N_9634,N_6870,N_6355);
xnor U9635 (N_9635,N_6104,N_7887);
nor U9636 (N_9636,N_7795,N_6088);
or U9637 (N_9637,N_7174,N_7564);
or U9638 (N_9638,N_6254,N_6675);
nand U9639 (N_9639,N_6449,N_6100);
and U9640 (N_9640,N_6450,N_7784);
nor U9641 (N_9641,N_7644,N_6787);
nor U9642 (N_9642,N_6861,N_7533);
xnor U9643 (N_9643,N_6596,N_7048);
nand U9644 (N_9644,N_7449,N_7635);
nand U9645 (N_9645,N_6788,N_6308);
nand U9646 (N_9646,N_7112,N_7016);
xnor U9647 (N_9647,N_7961,N_6126);
nand U9648 (N_9648,N_6218,N_7680);
nor U9649 (N_9649,N_7322,N_6609);
or U9650 (N_9650,N_6483,N_7017);
or U9651 (N_9651,N_7242,N_7331);
and U9652 (N_9652,N_6065,N_7973);
and U9653 (N_9653,N_6384,N_7921);
xor U9654 (N_9654,N_6457,N_7045);
nand U9655 (N_9655,N_6589,N_7812);
and U9656 (N_9656,N_6988,N_7804);
xor U9657 (N_9657,N_7471,N_6717);
or U9658 (N_9658,N_6208,N_6015);
or U9659 (N_9659,N_7404,N_6971);
and U9660 (N_9660,N_6147,N_7694);
xnor U9661 (N_9661,N_6889,N_7562);
nor U9662 (N_9662,N_6930,N_6456);
nor U9663 (N_9663,N_6181,N_6264);
nand U9664 (N_9664,N_7947,N_6850);
xnor U9665 (N_9665,N_6407,N_6406);
or U9666 (N_9666,N_7009,N_6618);
xnor U9667 (N_9667,N_7022,N_6795);
or U9668 (N_9668,N_7821,N_7344);
nor U9669 (N_9669,N_6890,N_7718);
nand U9670 (N_9670,N_6823,N_6525);
or U9671 (N_9671,N_6998,N_7781);
nand U9672 (N_9672,N_6189,N_7515);
xor U9673 (N_9673,N_7865,N_7399);
nand U9674 (N_9674,N_6789,N_6010);
nor U9675 (N_9675,N_7504,N_6494);
nand U9676 (N_9676,N_7808,N_7296);
and U9677 (N_9677,N_7928,N_7588);
nor U9678 (N_9678,N_6629,N_7668);
nor U9679 (N_9679,N_7366,N_7517);
nor U9680 (N_9680,N_7192,N_7011);
or U9681 (N_9681,N_6690,N_6639);
or U9682 (N_9682,N_7155,N_7811);
or U9683 (N_9683,N_6800,N_6471);
nor U9684 (N_9684,N_6383,N_6522);
and U9685 (N_9685,N_7288,N_6852);
and U9686 (N_9686,N_7866,N_7398);
and U9687 (N_9687,N_6765,N_6903);
or U9688 (N_9688,N_6351,N_6315);
or U9689 (N_9689,N_6446,N_6352);
nand U9690 (N_9690,N_7011,N_7016);
nor U9691 (N_9691,N_7595,N_7572);
or U9692 (N_9692,N_6389,N_6310);
xnor U9693 (N_9693,N_7112,N_7917);
nand U9694 (N_9694,N_7991,N_6650);
nor U9695 (N_9695,N_6198,N_7290);
xnor U9696 (N_9696,N_7782,N_6016);
xor U9697 (N_9697,N_6141,N_7870);
or U9698 (N_9698,N_7389,N_6995);
and U9699 (N_9699,N_7643,N_6129);
xnor U9700 (N_9700,N_6472,N_6925);
nand U9701 (N_9701,N_7080,N_6535);
nand U9702 (N_9702,N_7811,N_6011);
nor U9703 (N_9703,N_7045,N_7222);
and U9704 (N_9704,N_7869,N_7966);
nor U9705 (N_9705,N_6205,N_6497);
or U9706 (N_9706,N_6200,N_6202);
and U9707 (N_9707,N_7347,N_6772);
or U9708 (N_9708,N_6622,N_7199);
and U9709 (N_9709,N_7769,N_7400);
and U9710 (N_9710,N_7071,N_6359);
nor U9711 (N_9711,N_7857,N_6665);
nor U9712 (N_9712,N_7854,N_7979);
and U9713 (N_9713,N_6734,N_7778);
or U9714 (N_9714,N_6490,N_7803);
xor U9715 (N_9715,N_6714,N_7059);
or U9716 (N_9716,N_7969,N_6579);
and U9717 (N_9717,N_7150,N_7822);
or U9718 (N_9718,N_7703,N_7475);
and U9719 (N_9719,N_6385,N_7261);
nor U9720 (N_9720,N_7246,N_7563);
or U9721 (N_9721,N_7365,N_6450);
or U9722 (N_9722,N_6329,N_7249);
nor U9723 (N_9723,N_6933,N_6508);
nor U9724 (N_9724,N_7311,N_6836);
nand U9725 (N_9725,N_6405,N_6230);
nand U9726 (N_9726,N_7854,N_6557);
nand U9727 (N_9727,N_6081,N_6868);
nand U9728 (N_9728,N_6968,N_6898);
and U9729 (N_9729,N_7338,N_6808);
nor U9730 (N_9730,N_7658,N_7671);
and U9731 (N_9731,N_6485,N_6079);
nand U9732 (N_9732,N_7080,N_7543);
xnor U9733 (N_9733,N_6101,N_6475);
xnor U9734 (N_9734,N_6415,N_7061);
nand U9735 (N_9735,N_7771,N_6877);
nand U9736 (N_9736,N_7615,N_6849);
or U9737 (N_9737,N_7354,N_6705);
or U9738 (N_9738,N_7879,N_6089);
nand U9739 (N_9739,N_6998,N_6363);
and U9740 (N_9740,N_7600,N_7263);
nor U9741 (N_9741,N_6800,N_6565);
xor U9742 (N_9742,N_6529,N_6857);
or U9743 (N_9743,N_6666,N_7497);
and U9744 (N_9744,N_6311,N_7623);
nor U9745 (N_9745,N_6008,N_6426);
or U9746 (N_9746,N_6351,N_7854);
nand U9747 (N_9747,N_7103,N_7664);
nor U9748 (N_9748,N_6729,N_6440);
nand U9749 (N_9749,N_6921,N_6910);
and U9750 (N_9750,N_7168,N_6429);
or U9751 (N_9751,N_7023,N_6464);
nand U9752 (N_9752,N_7465,N_7752);
and U9753 (N_9753,N_6506,N_6984);
xnor U9754 (N_9754,N_7937,N_7315);
xnor U9755 (N_9755,N_7654,N_6269);
nor U9756 (N_9756,N_7116,N_7531);
nor U9757 (N_9757,N_7006,N_6381);
nor U9758 (N_9758,N_6425,N_7864);
and U9759 (N_9759,N_7338,N_6399);
xnor U9760 (N_9760,N_7559,N_7111);
and U9761 (N_9761,N_7198,N_6177);
and U9762 (N_9762,N_7521,N_7593);
or U9763 (N_9763,N_6506,N_7596);
nand U9764 (N_9764,N_7500,N_6976);
and U9765 (N_9765,N_7675,N_7107);
nor U9766 (N_9766,N_7819,N_6235);
or U9767 (N_9767,N_7787,N_6999);
xor U9768 (N_9768,N_7909,N_6728);
nor U9769 (N_9769,N_6752,N_6980);
xor U9770 (N_9770,N_6733,N_6834);
nor U9771 (N_9771,N_7710,N_6718);
or U9772 (N_9772,N_6121,N_6822);
or U9773 (N_9773,N_6644,N_6637);
xor U9774 (N_9774,N_6648,N_6821);
xnor U9775 (N_9775,N_6287,N_7997);
and U9776 (N_9776,N_6131,N_6775);
xor U9777 (N_9777,N_7092,N_7859);
and U9778 (N_9778,N_7606,N_7208);
nand U9779 (N_9779,N_6643,N_6623);
and U9780 (N_9780,N_6352,N_6469);
nor U9781 (N_9781,N_7748,N_6869);
and U9782 (N_9782,N_7901,N_7101);
or U9783 (N_9783,N_7745,N_6468);
nor U9784 (N_9784,N_6518,N_6223);
nor U9785 (N_9785,N_7874,N_6866);
and U9786 (N_9786,N_6878,N_6812);
nand U9787 (N_9787,N_7756,N_6715);
xnor U9788 (N_9788,N_6198,N_6687);
nand U9789 (N_9789,N_6548,N_6686);
and U9790 (N_9790,N_6246,N_6893);
and U9791 (N_9791,N_7471,N_7715);
nor U9792 (N_9792,N_7483,N_6856);
nor U9793 (N_9793,N_6020,N_6420);
or U9794 (N_9794,N_6188,N_7632);
and U9795 (N_9795,N_6085,N_7528);
or U9796 (N_9796,N_7551,N_6377);
or U9797 (N_9797,N_7893,N_7567);
xnor U9798 (N_9798,N_6161,N_6706);
or U9799 (N_9799,N_6446,N_6421);
nor U9800 (N_9800,N_7175,N_6696);
xnor U9801 (N_9801,N_6223,N_6779);
or U9802 (N_9802,N_6710,N_7203);
xnor U9803 (N_9803,N_6013,N_7760);
or U9804 (N_9804,N_6455,N_7358);
nand U9805 (N_9805,N_7664,N_6269);
and U9806 (N_9806,N_6539,N_6793);
nand U9807 (N_9807,N_7966,N_6581);
and U9808 (N_9808,N_7082,N_6512);
and U9809 (N_9809,N_7392,N_7268);
nand U9810 (N_9810,N_7779,N_6599);
xnor U9811 (N_9811,N_6997,N_6341);
xor U9812 (N_9812,N_6588,N_6949);
nand U9813 (N_9813,N_6244,N_7816);
or U9814 (N_9814,N_7677,N_7763);
nand U9815 (N_9815,N_7668,N_7429);
and U9816 (N_9816,N_7506,N_7028);
nor U9817 (N_9817,N_7484,N_6722);
and U9818 (N_9818,N_6787,N_6288);
xnor U9819 (N_9819,N_7216,N_7369);
nand U9820 (N_9820,N_7235,N_7459);
or U9821 (N_9821,N_6542,N_6419);
nor U9822 (N_9822,N_6359,N_7270);
nand U9823 (N_9823,N_6094,N_6517);
or U9824 (N_9824,N_7736,N_6470);
and U9825 (N_9825,N_6106,N_6419);
nor U9826 (N_9826,N_7218,N_7366);
and U9827 (N_9827,N_7818,N_7567);
and U9828 (N_9828,N_7892,N_6670);
nand U9829 (N_9829,N_6812,N_6533);
nor U9830 (N_9830,N_7081,N_7313);
and U9831 (N_9831,N_7077,N_6360);
or U9832 (N_9832,N_6213,N_6074);
and U9833 (N_9833,N_7332,N_6160);
nand U9834 (N_9834,N_7668,N_7414);
nor U9835 (N_9835,N_6270,N_6492);
xor U9836 (N_9836,N_6831,N_7401);
nand U9837 (N_9837,N_7948,N_7472);
nand U9838 (N_9838,N_6202,N_6161);
nor U9839 (N_9839,N_6205,N_7388);
nor U9840 (N_9840,N_7774,N_6541);
nand U9841 (N_9841,N_6706,N_6609);
xor U9842 (N_9842,N_7104,N_6608);
nor U9843 (N_9843,N_6609,N_6701);
xor U9844 (N_9844,N_7759,N_6705);
nand U9845 (N_9845,N_6557,N_7941);
nor U9846 (N_9846,N_7828,N_7320);
nor U9847 (N_9847,N_6135,N_7980);
and U9848 (N_9848,N_7897,N_6163);
or U9849 (N_9849,N_7373,N_7393);
or U9850 (N_9850,N_7629,N_7482);
nand U9851 (N_9851,N_7611,N_6915);
nand U9852 (N_9852,N_6434,N_6117);
nor U9853 (N_9853,N_7924,N_7557);
or U9854 (N_9854,N_6691,N_7975);
nor U9855 (N_9855,N_6940,N_6339);
xnor U9856 (N_9856,N_6052,N_6120);
and U9857 (N_9857,N_7144,N_7777);
xor U9858 (N_9858,N_6432,N_7921);
xnor U9859 (N_9859,N_7911,N_7900);
xor U9860 (N_9860,N_6423,N_7135);
and U9861 (N_9861,N_6193,N_7875);
nor U9862 (N_9862,N_6839,N_7546);
or U9863 (N_9863,N_7567,N_7121);
and U9864 (N_9864,N_6892,N_6069);
xor U9865 (N_9865,N_7734,N_6554);
or U9866 (N_9866,N_6306,N_7079);
xor U9867 (N_9867,N_6432,N_6593);
xnor U9868 (N_9868,N_7881,N_6620);
nor U9869 (N_9869,N_7003,N_6342);
xor U9870 (N_9870,N_7810,N_7554);
and U9871 (N_9871,N_7086,N_6563);
nand U9872 (N_9872,N_6206,N_6266);
or U9873 (N_9873,N_6092,N_7643);
or U9874 (N_9874,N_6730,N_6258);
and U9875 (N_9875,N_7655,N_7926);
nor U9876 (N_9876,N_7114,N_6823);
and U9877 (N_9877,N_7401,N_6042);
or U9878 (N_9878,N_6138,N_6954);
nor U9879 (N_9879,N_6848,N_7070);
and U9880 (N_9880,N_6838,N_6591);
nand U9881 (N_9881,N_7983,N_7461);
nand U9882 (N_9882,N_7895,N_7695);
nand U9883 (N_9883,N_6846,N_7979);
and U9884 (N_9884,N_6804,N_6077);
nand U9885 (N_9885,N_6747,N_7382);
or U9886 (N_9886,N_7851,N_7580);
and U9887 (N_9887,N_6901,N_7399);
nand U9888 (N_9888,N_7006,N_7861);
xnor U9889 (N_9889,N_7524,N_7260);
or U9890 (N_9890,N_6390,N_7586);
and U9891 (N_9891,N_7157,N_7700);
xnor U9892 (N_9892,N_7780,N_7963);
nor U9893 (N_9893,N_7341,N_7689);
and U9894 (N_9894,N_6208,N_6774);
nand U9895 (N_9895,N_6895,N_7268);
or U9896 (N_9896,N_6895,N_6942);
xnor U9897 (N_9897,N_7646,N_6005);
xor U9898 (N_9898,N_7972,N_7147);
nand U9899 (N_9899,N_6905,N_7431);
xnor U9900 (N_9900,N_7768,N_7906);
nand U9901 (N_9901,N_6705,N_7936);
nor U9902 (N_9902,N_7120,N_6312);
and U9903 (N_9903,N_7333,N_6591);
and U9904 (N_9904,N_7431,N_7636);
and U9905 (N_9905,N_6997,N_6927);
and U9906 (N_9906,N_6910,N_6780);
xnor U9907 (N_9907,N_7990,N_7040);
nand U9908 (N_9908,N_7934,N_6004);
xor U9909 (N_9909,N_6762,N_7494);
nand U9910 (N_9910,N_7161,N_7543);
or U9911 (N_9911,N_7089,N_6605);
nand U9912 (N_9912,N_6801,N_6639);
xor U9913 (N_9913,N_7165,N_6665);
nand U9914 (N_9914,N_7212,N_6762);
nand U9915 (N_9915,N_6739,N_7677);
or U9916 (N_9916,N_6447,N_6646);
nand U9917 (N_9917,N_6152,N_7004);
and U9918 (N_9918,N_6593,N_7161);
nand U9919 (N_9919,N_7289,N_7290);
xor U9920 (N_9920,N_7913,N_7988);
and U9921 (N_9921,N_6013,N_7811);
and U9922 (N_9922,N_7960,N_7493);
and U9923 (N_9923,N_6338,N_6027);
nand U9924 (N_9924,N_6872,N_7278);
or U9925 (N_9925,N_7966,N_6793);
xnor U9926 (N_9926,N_7610,N_6923);
or U9927 (N_9927,N_6693,N_7774);
or U9928 (N_9928,N_6723,N_6220);
nand U9929 (N_9929,N_7895,N_6921);
xnor U9930 (N_9930,N_6740,N_6320);
xor U9931 (N_9931,N_6408,N_7873);
nor U9932 (N_9932,N_6329,N_7911);
xnor U9933 (N_9933,N_7784,N_6819);
and U9934 (N_9934,N_6433,N_7242);
or U9935 (N_9935,N_6129,N_6782);
xnor U9936 (N_9936,N_6607,N_6894);
nand U9937 (N_9937,N_7636,N_7570);
nor U9938 (N_9938,N_7725,N_6611);
xnor U9939 (N_9939,N_6183,N_6592);
or U9940 (N_9940,N_6626,N_6008);
and U9941 (N_9941,N_7815,N_6609);
and U9942 (N_9942,N_6047,N_7721);
nor U9943 (N_9943,N_7141,N_6926);
nor U9944 (N_9944,N_6176,N_6989);
nand U9945 (N_9945,N_6319,N_7929);
and U9946 (N_9946,N_7597,N_7749);
xor U9947 (N_9947,N_6414,N_7810);
nor U9948 (N_9948,N_7296,N_6899);
nand U9949 (N_9949,N_6096,N_6420);
or U9950 (N_9950,N_7282,N_7582);
nor U9951 (N_9951,N_7908,N_6045);
nand U9952 (N_9952,N_7785,N_6985);
nor U9953 (N_9953,N_7340,N_6285);
xor U9954 (N_9954,N_7090,N_7511);
nor U9955 (N_9955,N_7250,N_7976);
xor U9956 (N_9956,N_6930,N_7513);
nand U9957 (N_9957,N_7770,N_7581);
or U9958 (N_9958,N_6673,N_7491);
nand U9959 (N_9959,N_7037,N_6116);
and U9960 (N_9960,N_7836,N_6856);
or U9961 (N_9961,N_7278,N_6940);
nor U9962 (N_9962,N_7798,N_6228);
nand U9963 (N_9963,N_6654,N_7799);
nor U9964 (N_9964,N_6987,N_6965);
xor U9965 (N_9965,N_7045,N_6285);
or U9966 (N_9966,N_6219,N_6602);
nor U9967 (N_9967,N_7762,N_7744);
xor U9968 (N_9968,N_7928,N_6789);
nor U9969 (N_9969,N_7712,N_6798);
or U9970 (N_9970,N_6559,N_6908);
or U9971 (N_9971,N_6992,N_6481);
or U9972 (N_9972,N_6772,N_6650);
xnor U9973 (N_9973,N_7776,N_7783);
or U9974 (N_9974,N_7297,N_7198);
or U9975 (N_9975,N_6873,N_7828);
or U9976 (N_9976,N_6362,N_7548);
nor U9977 (N_9977,N_7212,N_6866);
xnor U9978 (N_9978,N_6271,N_6439);
nor U9979 (N_9979,N_7475,N_7228);
nand U9980 (N_9980,N_6952,N_7291);
nand U9981 (N_9981,N_7446,N_6941);
nand U9982 (N_9982,N_7566,N_6996);
nand U9983 (N_9983,N_7539,N_7100);
nor U9984 (N_9984,N_6007,N_7408);
xnor U9985 (N_9985,N_6697,N_6678);
or U9986 (N_9986,N_7816,N_7886);
nor U9987 (N_9987,N_7707,N_6303);
nor U9988 (N_9988,N_7521,N_6243);
nor U9989 (N_9989,N_6254,N_7345);
nand U9990 (N_9990,N_6545,N_7951);
nor U9991 (N_9991,N_6912,N_7281);
nand U9992 (N_9992,N_7166,N_6727);
or U9993 (N_9993,N_6668,N_6037);
nor U9994 (N_9994,N_6649,N_6036);
xor U9995 (N_9995,N_7301,N_6038);
or U9996 (N_9996,N_6611,N_6836);
nor U9997 (N_9997,N_6828,N_6144);
nor U9998 (N_9998,N_7630,N_6829);
nand U9999 (N_9999,N_6132,N_6322);
nand U10000 (N_10000,N_8009,N_9794);
or U10001 (N_10001,N_9904,N_9239);
nor U10002 (N_10002,N_9583,N_9952);
nand U10003 (N_10003,N_9608,N_8852);
xnor U10004 (N_10004,N_9787,N_8329);
nor U10005 (N_10005,N_9784,N_8476);
xor U10006 (N_10006,N_9433,N_9716);
nor U10007 (N_10007,N_9225,N_8931);
nor U10008 (N_10008,N_9832,N_8529);
nand U10009 (N_10009,N_8877,N_9993);
or U10010 (N_10010,N_8681,N_9727);
and U10011 (N_10011,N_9493,N_8391);
nand U10012 (N_10012,N_8558,N_9294);
nor U10013 (N_10013,N_8628,N_9097);
and U10014 (N_10014,N_9461,N_8702);
or U10015 (N_10015,N_8651,N_9371);
or U10016 (N_10016,N_8661,N_9025);
nor U10017 (N_10017,N_9886,N_8217);
xor U10018 (N_10018,N_8600,N_9365);
nand U10019 (N_10019,N_9532,N_9694);
xor U10020 (N_10020,N_8381,N_8609);
and U10021 (N_10021,N_8924,N_9489);
nor U10022 (N_10022,N_9342,N_8131);
nand U10023 (N_10023,N_8906,N_9935);
xnor U10024 (N_10024,N_9723,N_9796);
and U10025 (N_10025,N_8575,N_8146);
nand U10026 (N_10026,N_9813,N_9776);
or U10027 (N_10027,N_9252,N_9878);
xnor U10028 (N_10028,N_8659,N_8492);
nand U10029 (N_10029,N_8481,N_8264);
and U10030 (N_10030,N_8098,N_8686);
xnor U10031 (N_10031,N_8197,N_8064);
xnor U10032 (N_10032,N_8000,N_9009);
and U10033 (N_10033,N_8074,N_8224);
or U10034 (N_10034,N_8284,N_8759);
and U10035 (N_10035,N_8996,N_9645);
and U10036 (N_10036,N_9159,N_8248);
xnor U10037 (N_10037,N_9254,N_8177);
xor U10038 (N_10038,N_9466,N_9057);
and U10039 (N_10039,N_8688,N_9803);
xor U10040 (N_10040,N_8103,N_8446);
nand U10041 (N_10041,N_9484,N_9315);
and U10042 (N_10042,N_9596,N_9859);
nand U10043 (N_10043,N_9641,N_8780);
nor U10044 (N_10044,N_8891,N_8901);
or U10045 (N_10045,N_9231,N_9205);
nand U10046 (N_10046,N_8701,N_8514);
nand U10047 (N_10047,N_9801,N_8049);
xor U10048 (N_10048,N_8505,N_9381);
nand U10049 (N_10049,N_8057,N_9293);
or U10050 (N_10050,N_9976,N_9635);
and U10051 (N_10051,N_9441,N_8148);
nand U10052 (N_10052,N_8301,N_9982);
and U10053 (N_10053,N_9033,N_8194);
and U10054 (N_10054,N_8537,N_9100);
nand U10055 (N_10055,N_8680,N_8771);
and U10056 (N_10056,N_8866,N_8497);
and U10057 (N_10057,N_9680,N_9606);
xnor U10058 (N_10058,N_9649,N_8261);
nor U10059 (N_10059,N_8305,N_9788);
and U10060 (N_10060,N_8174,N_9448);
nand U10061 (N_10061,N_9184,N_8119);
nand U10062 (N_10062,N_9196,N_9013);
or U10063 (N_10063,N_9705,N_8460);
and U10064 (N_10064,N_8795,N_8092);
nand U10065 (N_10065,N_9790,N_8489);
xor U10066 (N_10066,N_9800,N_8228);
nand U10067 (N_10067,N_9364,N_8640);
xor U10068 (N_10068,N_8854,N_8243);
xor U10069 (N_10069,N_9490,N_9944);
or U10070 (N_10070,N_8803,N_8849);
nor U10071 (N_10071,N_9912,N_9169);
nand U10072 (N_10072,N_9173,N_9749);
nand U10073 (N_10073,N_9158,N_9913);
and U10074 (N_10074,N_8533,N_8698);
nor U10075 (N_10075,N_8905,N_8732);
or U10076 (N_10076,N_9497,N_9517);
nand U10077 (N_10077,N_9191,N_8602);
and U10078 (N_10078,N_8495,N_9760);
xnor U10079 (N_10079,N_9568,N_9321);
nor U10080 (N_10080,N_8627,N_9619);
xnor U10081 (N_10081,N_9696,N_9729);
or U10082 (N_10082,N_9420,N_8766);
or U10083 (N_10083,N_9411,N_9856);
nor U10084 (N_10084,N_9594,N_8206);
xnor U10085 (N_10085,N_9947,N_9047);
or U10086 (N_10086,N_9609,N_8617);
xnor U10087 (N_10087,N_8531,N_8020);
nand U10088 (N_10088,N_8226,N_8626);
nand U10089 (N_10089,N_9921,N_9247);
nor U10090 (N_10090,N_9653,N_9302);
or U10091 (N_10091,N_9853,N_8090);
nand U10092 (N_10092,N_8504,N_8292);
nor U10093 (N_10093,N_8947,N_8536);
or U10094 (N_10094,N_8330,N_9133);
or U10095 (N_10095,N_9682,N_9602);
or U10096 (N_10096,N_8032,N_9094);
or U10097 (N_10097,N_8325,N_8080);
nand U10098 (N_10098,N_9015,N_8031);
nand U10099 (N_10099,N_8452,N_8973);
xnor U10100 (N_10100,N_8689,N_8653);
or U10101 (N_10101,N_8969,N_8585);
nor U10102 (N_10102,N_9277,N_9917);
or U10103 (N_10103,N_8298,N_9499);
or U10104 (N_10104,N_9415,N_8512);
nor U10105 (N_10105,N_8036,N_8503);
nand U10106 (N_10106,N_8511,N_9845);
and U10107 (N_10107,N_8500,N_8636);
and U10108 (N_10108,N_9745,N_8012);
nand U10109 (N_10109,N_9617,N_8915);
nand U10110 (N_10110,N_8844,N_9445);
nand U10111 (N_10111,N_9632,N_9377);
nand U10112 (N_10112,N_8084,N_8096);
or U10113 (N_10113,N_9345,N_8438);
nand U10114 (N_10114,N_9123,N_8925);
and U10115 (N_10115,N_9049,N_8216);
xnor U10116 (N_10116,N_8315,N_8233);
and U10117 (N_10117,N_9238,N_8610);
xor U10118 (N_10118,N_8061,N_8188);
nand U10119 (N_10119,N_8705,N_8142);
or U10120 (N_10120,N_8839,N_8480);
or U10121 (N_10121,N_9193,N_8379);
nand U10122 (N_10122,N_9915,N_9156);
or U10123 (N_10123,N_8250,N_8351);
nor U10124 (N_10124,N_9740,N_9018);
xor U10125 (N_10125,N_9126,N_9873);
or U10126 (N_10126,N_8453,N_8059);
or U10127 (N_10127,N_9422,N_9836);
xnor U10128 (N_10128,N_9551,N_9945);
and U10129 (N_10129,N_9750,N_8909);
and U10130 (N_10130,N_9770,N_9084);
or U10131 (N_10131,N_8373,N_9661);
nand U10132 (N_10132,N_9029,N_8355);
and U10133 (N_10133,N_8784,N_8730);
nor U10134 (N_10134,N_8644,N_9523);
nor U10135 (N_10135,N_9052,N_8521);
xnor U10136 (N_10136,N_8790,N_9809);
or U10137 (N_10137,N_8593,N_9303);
nor U10138 (N_10138,N_8836,N_8294);
nand U10139 (N_10139,N_8742,N_8265);
nand U10140 (N_10140,N_9147,N_9791);
nor U10141 (N_10141,N_9469,N_9000);
nand U10142 (N_10142,N_9533,N_9369);
xor U10143 (N_10143,N_9177,N_8941);
xnor U10144 (N_10144,N_8138,N_9937);
nor U10145 (N_10145,N_9736,N_9181);
nor U10146 (N_10146,N_8992,N_9704);
nand U10147 (N_10147,N_8756,N_8753);
xnor U10148 (N_10148,N_8578,N_9862);
nor U10149 (N_10149,N_9037,N_8683);
xor U10150 (N_10150,N_9567,N_8582);
nand U10151 (N_10151,N_8193,N_8339);
or U10152 (N_10152,N_8252,N_9578);
xnor U10153 (N_10153,N_9633,N_9462);
or U10154 (N_10154,N_9120,N_8477);
nand U10155 (N_10155,N_8372,N_9317);
xor U10156 (N_10156,N_9703,N_8458);
or U10157 (N_10157,N_8786,N_9706);
nor U10158 (N_10158,N_8011,N_9540);
and U10159 (N_10159,N_8955,N_9206);
xnor U10160 (N_10160,N_8450,N_9827);
or U10161 (N_10161,N_8898,N_9201);
and U10162 (N_10162,N_9604,N_8390);
xor U10163 (N_10163,N_8740,N_9848);
nor U10164 (N_10164,N_9419,N_8605);
and U10165 (N_10165,N_9136,N_8408);
xor U10166 (N_10166,N_9652,N_8868);
and U10167 (N_10167,N_8069,N_9591);
xnor U10168 (N_10168,N_8184,N_8806);
nor U10169 (N_10169,N_8833,N_9542);
or U10170 (N_10170,N_8321,N_8407);
xor U10171 (N_10171,N_8101,N_9061);
nor U10172 (N_10172,N_8162,N_8997);
or U10173 (N_10173,N_8869,N_9732);
nor U10174 (N_10174,N_9687,N_8630);
and U10175 (N_10175,N_8612,N_8451);
or U10176 (N_10176,N_9797,N_9688);
xor U10177 (N_10177,N_8758,N_8035);
and U10178 (N_10178,N_9036,N_8275);
nor U10179 (N_10179,N_9217,N_8274);
nand U10180 (N_10180,N_9629,N_9927);
and U10181 (N_10181,N_8879,N_8423);
nor U10182 (N_10182,N_9566,N_9424);
xor U10183 (N_10183,N_8914,N_9308);
and U10184 (N_10184,N_8562,N_9949);
nor U10185 (N_10185,N_8729,N_9785);
or U10186 (N_10186,N_8871,N_8970);
xor U10187 (N_10187,N_8728,N_8387);
xor U10188 (N_10188,N_8894,N_8136);
or U10189 (N_10189,N_9710,N_8318);
xor U10190 (N_10190,N_8362,N_8178);
and U10191 (N_10191,N_9051,N_9505);
xor U10192 (N_10192,N_9820,N_8870);
xor U10193 (N_10193,N_8077,N_9486);
or U10194 (N_10194,N_9011,N_8733);
nor U10195 (N_10195,N_8989,N_8073);
and U10196 (N_10196,N_9387,N_9228);
or U10197 (N_10197,N_9518,N_9581);
nor U10198 (N_10198,N_8980,N_9799);
or U10199 (N_10199,N_9874,N_9669);
xor U10200 (N_10200,N_8949,N_8889);
nor U10201 (N_10201,N_8144,N_8140);
nand U10202 (N_10202,N_9108,N_8694);
nand U10203 (N_10203,N_9202,N_9452);
and U10204 (N_10204,N_8246,N_9507);
xnor U10205 (N_10205,N_9409,N_8106);
nand U10206 (N_10206,N_9455,N_8864);
or U10207 (N_10207,N_8097,N_9375);
xor U10208 (N_10208,N_8621,N_9435);
nand U10209 (N_10209,N_9751,N_9292);
xor U10210 (N_10210,N_8436,N_8165);
xor U10211 (N_10211,N_9279,N_9816);
nor U10212 (N_10212,N_8191,N_9979);
and U10213 (N_10213,N_9022,N_8115);
xor U10214 (N_10214,N_8897,N_9597);
nor U10215 (N_10215,N_9739,N_8764);
xor U10216 (N_10216,N_8647,N_9166);
xnor U10217 (N_10217,N_8616,N_9906);
nand U10218 (N_10218,N_9837,N_8723);
or U10219 (N_10219,N_8555,N_8048);
nor U10220 (N_10220,N_8768,N_9464);
nand U10221 (N_10221,N_8703,N_8591);
and U10222 (N_10222,N_8545,N_9589);
or U10223 (N_10223,N_8385,N_9646);
nor U10224 (N_10224,N_9341,N_9271);
or U10225 (N_10225,N_9755,N_9062);
xor U10226 (N_10226,N_9686,N_9471);
and U10227 (N_10227,N_8026,N_8171);
nand U10228 (N_10228,N_8260,N_9351);
and U10229 (N_10229,N_9167,N_9953);
xnor U10230 (N_10230,N_8952,N_9130);
and U10231 (N_10231,N_8002,N_8066);
nor U10232 (N_10232,N_8649,N_9726);
xor U10233 (N_10233,N_9880,N_8722);
xnor U10234 (N_10234,N_8058,N_8067);
and U10235 (N_10235,N_8276,N_9242);
nor U10236 (N_10236,N_8513,N_9431);
and U10237 (N_10237,N_9907,N_8382);
or U10238 (N_10238,N_9195,N_8884);
xor U10239 (N_10239,N_9257,N_8123);
nand U10240 (N_10240,N_8961,N_8209);
or U10241 (N_10241,N_8946,N_9972);
nor U10242 (N_10242,N_9373,N_8682);
or U10243 (N_10243,N_9849,N_9519);
or U10244 (N_10244,N_9630,N_9223);
and U10245 (N_10245,N_9414,N_9512);
and U10246 (N_10246,N_9418,N_9870);
xnor U10247 (N_10247,N_8323,N_8834);
and U10248 (N_10248,N_9742,N_8147);
xor U10249 (N_10249,N_9931,N_8523);
xnor U10250 (N_10250,N_8781,N_9556);
xor U10251 (N_10251,N_9587,N_8203);
or U10252 (N_10252,N_8467,N_9086);
nor U10253 (N_10253,N_8639,N_8974);
nand U10254 (N_10254,N_8972,N_9973);
or U10255 (N_10255,N_9657,N_9383);
or U10256 (N_10256,N_8645,N_8375);
or U10257 (N_10257,N_8642,N_8071);
xnor U10258 (N_10258,N_8485,N_9155);
and U10259 (N_10259,N_8114,N_8517);
nand U10260 (N_10260,N_8724,N_8953);
and U10261 (N_10261,N_8402,N_8968);
nor U10262 (N_10262,N_8386,N_8300);
or U10263 (N_10263,N_8113,N_8629);
nor U10264 (N_10264,N_9258,N_8079);
nor U10265 (N_10265,N_8690,N_8003);
or U10266 (N_10266,N_8900,N_8872);
xor U10267 (N_10267,N_8230,N_8763);
or U10268 (N_10268,N_8283,N_9747);
or U10269 (N_10269,N_8404,N_8999);
nand U10270 (N_10270,N_9132,N_8320);
or U10271 (N_10271,N_8308,N_9525);
xnor U10272 (N_10272,N_8405,N_8775);
nand U10273 (N_10273,N_9528,N_9334);
xnor U10274 (N_10274,N_9808,N_8643);
xnor U10275 (N_10275,N_8401,N_9220);
or U10276 (N_10276,N_8739,N_9081);
or U10277 (N_10277,N_8396,N_9823);
and U10278 (N_10278,N_9554,N_8470);
nor U10279 (N_10279,N_8708,N_9187);
and U10280 (N_10280,N_9579,N_9361);
and U10281 (N_10281,N_8825,N_9693);
xor U10282 (N_10282,N_9040,N_8416);
and U10283 (N_10283,N_8544,N_9143);
xor U10284 (N_10284,N_8530,N_9001);
and U10285 (N_10285,N_9472,N_8371);
nor U10286 (N_10286,N_8977,N_8215);
nor U10287 (N_10287,N_9311,N_9316);
nor U10288 (N_10288,N_8161,N_9582);
xnor U10289 (N_10289,N_8338,N_8368);
xor U10290 (N_10290,N_9988,N_9203);
and U10291 (N_10291,N_8590,N_9936);
or U10292 (N_10292,N_8821,N_8021);
xnor U10293 (N_10293,N_8310,N_8772);
and U10294 (N_10294,N_9229,N_8851);
nor U10295 (N_10295,N_8176,N_9867);
or U10296 (N_10296,N_9875,N_8346);
and U10297 (N_10297,N_8041,N_8172);
nand U10298 (N_10298,N_8859,N_9970);
or U10299 (N_10299,N_9104,N_8285);
nor U10300 (N_10300,N_8774,N_9207);
xor U10301 (N_10301,N_8519,N_9208);
nor U10302 (N_10302,N_8637,N_8154);
or U10303 (N_10303,N_8887,N_9073);
nor U10304 (N_10304,N_9851,N_8822);
or U10305 (N_10305,N_8302,N_9610);
and U10306 (N_10306,N_9668,N_8410);
xnor U10307 (N_10307,N_9131,N_8873);
nor U10308 (N_10308,N_8374,N_8152);
xor U10309 (N_10309,N_8309,N_9508);
or U10310 (N_10310,N_8847,N_9349);
nand U10311 (N_10311,N_8076,N_9850);
nor U10312 (N_10312,N_8631,N_9707);
xnor U10313 (N_10313,N_9004,N_9529);
or U10314 (N_10314,N_8672,N_9288);
nand U10315 (N_10315,N_9103,N_8950);
and U10316 (N_10316,N_9889,N_9847);
and U10317 (N_10317,N_8473,N_9975);
nor U10318 (N_10318,N_9868,N_9457);
xor U10319 (N_10319,N_9607,N_8607);
nor U10320 (N_10320,N_8288,N_8799);
xor U10321 (N_10321,N_8322,N_8182);
xor U10322 (N_10322,N_9185,N_9614);
and U10323 (N_10323,N_9285,N_9593);
and U10324 (N_10324,N_9685,N_8155);
or U10325 (N_10325,N_9164,N_9830);
nor U10326 (N_10326,N_9453,N_9246);
nor U10327 (N_10327,N_9929,N_9183);
nor U10328 (N_10328,N_8549,N_8815);
nor U10329 (N_10329,N_9230,N_9775);
xor U10330 (N_10330,N_9658,N_9172);
and U10331 (N_10331,N_8581,N_9188);
or U10332 (N_10332,N_8269,N_9459);
nand U10333 (N_10333,N_9428,N_9374);
nand U10334 (N_10334,N_9140,N_9950);
nor U10335 (N_10335,N_8938,N_8001);
or U10336 (N_10336,N_9006,N_9838);
nor U10337 (N_10337,N_8911,N_8664);
nand U10338 (N_10338,N_8624,N_8056);
xor U10339 (N_10339,N_9503,N_9436);
or U10340 (N_10340,N_9672,N_9574);
and U10341 (N_10341,N_8807,N_8359);
and U10342 (N_10342,N_8124,N_9400);
nand U10343 (N_10343,N_9069,N_8366);
xor U10344 (N_10344,N_8565,N_9485);
and U10345 (N_10345,N_9746,N_9286);
nand U10346 (N_10346,N_9833,N_8944);
or U10347 (N_10347,N_8024,N_9628);
nor U10348 (N_10348,N_8055,N_8757);
and U10349 (N_10349,N_8561,N_8420);
nor U10350 (N_10350,N_8711,N_8595);
xnor U10351 (N_10351,N_9482,N_8455);
and U10352 (N_10352,N_9941,N_8456);
and U10353 (N_10353,N_9038,N_8546);
xor U10354 (N_10354,N_9779,N_9417);
nor U10355 (N_10355,N_8468,N_8223);
and U10356 (N_10356,N_9841,N_8658);
and U10357 (N_10357,N_8618,N_8717);
and U10358 (N_10358,N_9210,N_9538);
nand U10359 (N_10359,N_8232,N_8910);
nand U10360 (N_10360,N_9980,N_9249);
nand U10361 (N_10361,N_9437,N_9291);
nand U10362 (N_10362,N_9212,N_9267);
nand U10363 (N_10363,N_9079,N_9226);
and U10364 (N_10364,N_9721,N_9115);
nand U10365 (N_10365,N_8427,N_9692);
and U10366 (N_10366,N_8027,N_8479);
or U10367 (N_10367,N_9888,N_9082);
or U10368 (N_10368,N_8328,N_8376);
nor U10369 (N_10369,N_9216,N_8266);
nor U10370 (N_10370,N_9359,N_9048);
xnor U10371 (N_10371,N_9987,N_9541);
or U10372 (N_10372,N_9717,N_9449);
nand U10373 (N_10373,N_9480,N_9440);
and U10374 (N_10374,N_8334,N_8258);
or U10375 (N_10375,N_9698,N_9733);
nand U10376 (N_10376,N_8179,N_9899);
nand U10377 (N_10377,N_8981,N_9432);
and U10378 (N_10378,N_9378,N_9241);
and U10379 (N_10379,N_8107,N_9588);
or U10380 (N_10380,N_9251,N_8572);
nor U10381 (N_10381,N_8560,N_8463);
and U10382 (N_10382,N_9691,N_8615);
or U10383 (N_10383,N_8158,N_9034);
xnor U10384 (N_10384,N_9088,N_8008);
or U10385 (N_10385,N_9798,N_8710);
nor U10386 (N_10386,N_9531,N_8475);
xnor U10387 (N_10387,N_9676,N_8983);
nand U10388 (N_10388,N_8282,N_8262);
xor U10389 (N_10389,N_9909,N_8229);
xor U10390 (N_10390,N_8358,N_8291);
or U10391 (N_10391,N_9546,N_8242);
nor U10392 (N_10392,N_8670,N_9430);
or U10393 (N_10393,N_9180,N_9865);
nor U10394 (N_10394,N_9442,N_9110);
and U10395 (N_10395,N_9186,N_8608);
or U10396 (N_10396,N_9817,N_9930);
nand U10397 (N_10397,N_8222,N_9618);
nor U10398 (N_10398,N_9928,N_8133);
nand U10399 (N_10399,N_8982,N_9272);
xnor U10400 (N_10400,N_9340,N_8044);
xor U10401 (N_10401,N_8676,N_9117);
or U10402 (N_10402,N_9262,N_9215);
xor U10403 (N_10403,N_9537,N_9677);
xnor U10404 (N_10404,N_8586,N_8400);
nor U10405 (N_10405,N_8287,N_9268);
and U10406 (N_10406,N_9569,N_9160);
nand U10407 (N_10407,N_8445,N_8589);
and U10408 (N_10408,N_8743,N_8361);
xnor U10409 (N_10409,N_8802,N_9520);
nand U10410 (N_10410,N_9766,N_8860);
nor U10411 (N_10411,N_8395,N_9974);
or U10412 (N_10412,N_9883,N_9571);
or U10413 (N_10413,N_8959,N_9995);
and U10414 (N_10414,N_9762,N_9943);
or U10415 (N_10415,N_8614,N_8019);
nand U10416 (N_10416,N_9240,N_9500);
xnor U10417 (N_10417,N_9324,N_8139);
nand U10418 (N_10418,N_8432,N_8820);
nor U10419 (N_10419,N_8765,N_8352);
nor U10420 (N_10420,N_9450,N_9358);
or U10421 (N_10421,N_9095,N_8399);
or U10422 (N_10422,N_8199,N_9911);
xnor U10423 (N_10423,N_8932,N_9516);
nor U10424 (N_10424,N_9300,N_8838);
xnor U10425 (N_10425,N_9237,N_9664);
nor U10426 (N_10426,N_8313,N_8297);
or U10427 (N_10427,N_8028,N_8837);
xnor U10428 (N_10428,N_8662,N_8263);
nand U10429 (N_10429,N_8665,N_8515);
or U10430 (N_10430,N_8738,N_8335);
xnor U10431 (N_10431,N_8882,N_9942);
or U10432 (N_10432,N_8259,N_9218);
or U10433 (N_10433,N_8281,N_8207);
and U10434 (N_10434,N_9957,N_8472);
nand U10435 (N_10435,N_8016,N_9968);
or U10436 (N_10436,N_8340,N_9168);
nand U10437 (N_10437,N_9329,N_9125);
and U10438 (N_10438,N_8967,N_9319);
nand U10439 (N_10439,N_8566,N_8777);
nand U10440 (N_10440,N_9902,N_9603);
xnor U10441 (N_10441,N_9895,N_8474);
and U10442 (N_10442,N_8798,N_8563);
and U10443 (N_10443,N_8746,N_9368);
xnor U10444 (N_10444,N_9429,N_9498);
nor U10445 (N_10445,N_8443,N_9310);
and U10446 (N_10446,N_8135,N_9557);
and U10447 (N_10447,N_8137,N_8863);
and U10448 (N_10448,N_9028,N_9994);
nand U10449 (N_10449,N_9659,N_9406);
or U10450 (N_10450,N_9623,N_8579);
or U10451 (N_10451,N_8449,N_8018);
nand U10452 (N_10452,N_8062,N_8010);
and U10453 (N_10453,N_8792,N_8535);
xor U10454 (N_10454,N_9356,N_8173);
xnor U10455 (N_10455,N_8333,N_9697);
nor U10456 (N_10456,N_8788,N_9427);
or U10457 (N_10457,N_9376,N_9289);
xnor U10458 (N_10458,N_8760,N_9275);
and U10459 (N_10459,N_8988,N_8945);
xnor U10460 (N_10460,N_9007,N_8271);
and U10461 (N_10461,N_8697,N_8594);
nor U10462 (N_10462,N_8421,N_8160);
nand U10463 (N_10463,N_8934,N_8151);
xnor U10464 (N_10464,N_8735,N_9810);
xor U10465 (N_10465,N_9852,N_9107);
xnor U10466 (N_10466,N_8337,N_9807);
or U10467 (N_10467,N_8431,N_8380);
and U10468 (N_10468,N_9363,N_8826);
xor U10469 (N_10469,N_8070,N_9655);
and U10470 (N_10470,N_8181,N_9992);
and U10471 (N_10471,N_9743,N_9956);
or U10472 (N_10472,N_8095,N_9305);
xor U10473 (N_10473,N_8406,N_9621);
nand U10474 (N_10474,N_8773,N_9394);
xnor U10475 (N_10475,N_8039,N_9297);
and U10476 (N_10476,N_8611,N_8674);
and U10477 (N_10477,N_8800,N_8948);
and U10478 (N_10478,N_9922,N_8874);
or U10479 (N_10479,N_9559,N_8005);
nand U10480 (N_10480,N_9598,N_9331);
or U10481 (N_10481,N_9724,N_9266);
nand U10482 (N_10482,N_9078,N_8078);
nand U10483 (N_10483,N_9157,N_9021);
nand U10484 (N_10484,N_8324,N_9933);
xnor U10485 (N_10485,N_8065,N_9397);
nand U10486 (N_10486,N_8522,N_9565);
and U10487 (N_10487,N_8750,N_9413);
nand U10488 (N_10488,N_9304,N_9198);
xnor U10489 (N_10489,N_9054,N_8200);
and U10490 (N_10490,N_9651,N_9720);
and U10491 (N_10491,N_9666,N_8571);
xor U10492 (N_10492,N_9773,N_8237);
or U10493 (N_10493,N_9625,N_9410);
nand U10494 (N_10494,N_8116,N_9113);
and U10495 (N_10495,N_9058,N_9350);
and U10496 (N_10496,N_8706,N_8306);
nor U10497 (N_10497,N_8189,N_9134);
nand U10498 (N_10498,N_9347,N_8597);
nand U10499 (N_10499,N_9256,N_8539);
nand U10500 (N_10500,N_9446,N_8634);
xnor U10501 (N_10501,N_9020,N_9407);
nand U10502 (N_10502,N_8933,N_8086);
nand U10503 (N_10503,N_8397,N_8761);
xnor U10504 (N_10504,N_9802,N_9337);
nor U10505 (N_10505,N_9127,N_9227);
or U10506 (N_10506,N_8244,N_8118);
and U10507 (N_10507,N_9199,N_9575);
nor U10508 (N_10508,N_9932,N_9274);
nand U10509 (N_10509,N_9398,N_9026);
and U10510 (N_10510,N_9362,N_9154);
nand U10511 (N_10511,N_8141,N_9370);
or U10512 (N_10512,N_8129,N_8937);
and U10513 (N_10513,N_9738,N_8403);
or U10514 (N_10514,N_8417,N_9767);
nor U10515 (N_10515,N_8483,N_8211);
nand U10516 (N_10516,N_8030,N_8951);
xnor U10517 (N_10517,N_8164,N_9178);
nand U10518 (N_10518,N_9473,N_9884);
or U10519 (N_10519,N_9301,N_9416);
or U10520 (N_10520,N_8804,N_9744);
nor U10521 (N_10521,N_9355,N_9121);
or U10522 (N_10522,N_8344,N_8047);
nor U10523 (N_10523,N_9600,N_8559);
or U10524 (N_10524,N_9111,N_9615);
nor U10525 (N_10525,N_9096,N_9562);
xor U10526 (N_10526,N_9580,N_8442);
nand U10527 (N_10527,N_9162,N_9754);
or U10528 (N_10528,N_8940,N_8707);
xnor U10529 (N_10529,N_9515,N_9656);
nand U10530 (N_10530,N_8430,N_8731);
and U10531 (N_10531,N_9654,N_8893);
and U10532 (N_10532,N_8994,N_8130);
nand U10533 (N_10533,N_9234,N_9759);
and U10534 (N_10534,N_9914,N_9881);
xnor U10535 (N_10535,N_9761,N_8128);
or U10536 (N_10536,N_8506,N_9637);
nand U10537 (N_10537,N_8567,N_9639);
and U10538 (N_10538,N_8532,N_9966);
nand U10539 (N_10539,N_8890,N_8004);
nor U10540 (N_10540,N_8508,N_9024);
nand U10541 (N_10541,N_9741,N_9327);
nand U10542 (N_10542,N_9783,N_9248);
or U10543 (N_10543,N_9782,N_8527);
xor U10544 (N_10544,N_9576,N_9290);
and U10545 (N_10545,N_8409,N_8196);
nand U10546 (N_10546,N_9395,N_9483);
or U10547 (N_10547,N_9521,N_9900);
nand U10548 (N_10548,N_9535,N_9855);
xor U10549 (N_10549,N_9163,N_8633);
nand U10550 (N_10550,N_9866,N_8231);
or U10551 (N_10551,N_9320,N_9963);
or U10552 (N_10552,N_9718,N_8556);
xor U10553 (N_10553,N_9991,N_9959);
nor U10554 (N_10554,N_9998,N_9434);
nor U10555 (N_10555,N_9940,N_9366);
xor U10556 (N_10556,N_8726,N_9438);
or U10557 (N_10557,N_9592,N_8202);
or U10558 (N_10558,N_9488,N_9481);
xor U10559 (N_10559,N_9002,N_8394);
xor U10560 (N_10560,N_8520,N_8289);
nor U10561 (N_10561,N_9918,N_8493);
or U10562 (N_10562,N_9098,N_8022);
and U10563 (N_10563,N_8251,N_9897);
nor U10564 (N_10564,N_9971,N_8125);
and U10565 (N_10565,N_9792,N_8907);
or U10566 (N_10566,N_8635,N_9129);
nand U10567 (N_10567,N_9492,N_8797);
or U10568 (N_10568,N_9352,N_9209);
or U10569 (N_10569,N_8721,N_8214);
nand U10570 (N_10570,N_9077,N_8132);
or U10571 (N_10571,N_8525,N_8696);
or U10572 (N_10572,N_9030,N_8936);
nor U10573 (N_10573,N_8034,N_8169);
and U10574 (N_10574,N_8060,N_8687);
nor U10575 (N_10575,N_8678,N_8081);
and U10576 (N_10576,N_8964,N_9804);
nand U10577 (N_10577,N_8895,N_9699);
and U10578 (N_10578,N_9662,N_8083);
nor U10579 (N_10579,N_9824,N_9831);
and U10580 (N_10580,N_9451,N_9323);
or U10581 (N_10581,N_8239,N_9674);
xor U10582 (N_10582,N_8923,N_8916);
nor U10583 (N_10583,N_8577,N_9421);
or U10584 (N_10584,N_9343,N_9425);
nand U10585 (N_10585,N_9616,N_9843);
nand U10586 (N_10586,N_9601,N_9961);
nand U10587 (N_10587,N_8314,N_9224);
or U10588 (N_10588,N_8712,N_9695);
nor U10589 (N_10589,N_8878,N_9871);
nor U10590 (N_10590,N_9312,N_8652);
xnor U10591 (N_10591,N_8052,N_8279);
and U10592 (N_10592,N_8876,N_8979);
xnor U10593 (N_10593,N_8277,N_9118);
xnor U10594 (N_10594,N_9690,N_8935);
and U10595 (N_10595,N_9584,N_9644);
nor U10596 (N_10596,N_8411,N_8810);
nor U10597 (N_10597,N_9728,N_9105);
and U10598 (N_10598,N_9265,N_8551);
xor U10599 (N_10599,N_8720,N_9681);
xor U10600 (N_10600,N_9951,N_8675);
or U10601 (N_10601,N_8827,N_9017);
and U10602 (N_10602,N_8167,N_8855);
nand U10603 (N_10603,N_9506,N_9116);
xnor U10604 (N_10604,N_9526,N_8013);
or U10605 (N_10605,N_8596,N_8484);
nand U10606 (N_10606,N_8435,N_9314);
or U10607 (N_10607,N_9939,N_8332);
and U10608 (N_10608,N_9236,N_9905);
and U10609 (N_10609,N_8692,N_9821);
nor U10610 (N_10610,N_8718,N_9549);
xnor U10611 (N_10611,N_9467,N_8033);
and U10612 (N_10612,N_9825,N_8848);
or U10613 (N_10613,N_8091,N_8159);
or U10614 (N_10614,N_8714,N_8153);
nor U10615 (N_10615,N_9380,N_8111);
nand U10616 (N_10616,N_9715,N_8814);
and U10617 (N_10617,N_9269,N_8466);
and U10618 (N_10618,N_8312,N_9408);
or U10619 (N_10619,N_9065,N_8388);
nor U10620 (N_10620,N_9260,N_9829);
and U10621 (N_10621,N_9711,N_9175);
and U10622 (N_10622,N_9055,N_8755);
nor U10623 (N_10623,N_9955,N_8553);
nand U10624 (N_10624,N_8122,N_9553);
xnor U10625 (N_10625,N_9511,N_8029);
and U10626 (N_10626,N_8516,N_8927);
nand U10627 (N_10627,N_8747,N_9984);
xnor U10628 (N_10628,N_8304,N_8606);
xor U10629 (N_10629,N_8198,N_8220);
nand U10630 (N_10630,N_8441,N_8255);
or U10631 (N_10631,N_8121,N_8528);
and U10632 (N_10632,N_8347,N_8424);
and U10633 (N_10633,N_8867,N_9090);
and U10634 (N_10634,N_9650,N_9857);
nor U10635 (N_10635,N_9805,N_9080);
or U10636 (N_10636,N_9444,N_8037);
nor U10637 (N_10637,N_8748,N_8767);
xnor U10638 (N_10638,N_8235,N_8418);
and U10639 (N_10639,N_8384,N_9660);
xor U10640 (N_10640,N_8105,N_9572);
xor U10641 (N_10641,N_9385,N_9882);
nor U10642 (N_10642,N_9958,N_8749);
or U10643 (N_10643,N_8524,N_8054);
nand U10644 (N_10644,N_8234,N_8741);
xnor U10645 (N_10645,N_8419,N_8965);
and U10646 (N_10646,N_8770,N_9948);
and U10647 (N_10647,N_8236,N_9276);
nand U10648 (N_10648,N_8023,N_9670);
nor U10649 (N_10649,N_8326,N_8241);
nand U10650 (N_10650,N_9046,N_8225);
nor U10651 (N_10651,N_9780,N_9032);
nor U10652 (N_10652,N_8623,N_9771);
xor U10653 (N_10653,N_9713,N_9233);
xor U10654 (N_10654,N_9283,N_8085);
xor U10655 (N_10655,N_8902,N_8272);
nor U10656 (N_10656,N_9014,N_9834);
xnor U10657 (N_10657,N_9719,N_9977);
and U10658 (N_10658,N_8087,N_9093);
xnor U10659 (N_10659,N_9896,N_9259);
and U10660 (N_10660,N_8254,N_8862);
or U10661 (N_10661,N_8247,N_8638);
nor U10662 (N_10662,N_8912,N_8256);
and U10663 (N_10663,N_9068,N_9863);
xor U10664 (N_10664,N_8072,N_9643);
nand U10665 (N_10665,N_8883,N_8094);
nand U10666 (N_10666,N_8960,N_9357);
or U10667 (N_10667,N_8620,N_8482);
nor U10668 (N_10668,N_9039,N_8502);
xnor U10669 (N_10669,N_8580,N_8824);
xnor U10670 (N_10670,N_8045,N_8109);
and U10671 (N_10671,N_8754,N_8365);
nor U10672 (N_10672,N_9124,N_9031);
or U10673 (N_10673,N_8303,N_8956);
and U10674 (N_10674,N_9712,N_8360);
and U10675 (N_10675,N_8110,N_9468);
nand U10676 (N_10676,N_8853,N_8439);
nor U10677 (N_10677,N_8296,N_9510);
nor U10678 (N_10678,N_8604,N_8370);
nand U10679 (N_10679,N_8267,N_9089);
and U10680 (N_10680,N_8584,N_9182);
nor U10681 (N_10681,N_9527,N_8543);
and U10682 (N_10682,N_8677,N_8829);
nand U10683 (N_10683,N_9573,N_9338);
or U10684 (N_10684,N_9954,N_9112);
nor U10685 (N_10685,N_8538,N_8858);
nor U10686 (N_10686,N_8063,N_9035);
nor U10687 (N_10687,N_9978,N_8699);
and U10688 (N_10688,N_9737,N_9388);
xor U10689 (N_10689,N_9232,N_9545);
and U10690 (N_10690,N_8995,N_9908);
nand U10691 (N_10691,N_8112,N_9585);
nand U10692 (N_10692,N_8319,N_9076);
xor U10693 (N_10693,N_8903,N_8392);
nand U10694 (N_10694,N_9620,N_9964);
nor U10695 (N_10695,N_9854,N_8613);
xnor U10696 (N_10696,N_8212,N_9638);
or U10697 (N_10697,N_9458,N_9270);
nor U10698 (N_10698,N_8440,N_9923);
or U10699 (N_10699,N_8422,N_9530);
and U10700 (N_10700,N_8782,N_8278);
nand U10701 (N_10701,N_8857,N_9734);
and U10702 (N_10702,N_8679,N_8377);
and U10703 (N_10703,N_9135,N_9916);
nand U10704 (N_10704,N_8428,N_9764);
xnor U10705 (N_10705,N_9064,N_9335);
nand U10706 (N_10706,N_9826,N_8666);
and U10707 (N_10707,N_9642,N_9513);
and U10708 (N_10708,N_8488,N_8971);
and U10709 (N_10709,N_8715,N_8478);
xnor U10710 (N_10710,N_9967,N_9284);
or U10711 (N_10711,N_9273,N_8709);
and U10712 (N_10712,N_9748,N_8930);
and U10713 (N_10713,N_9811,N_8501);
xor U10714 (N_10714,N_8088,N_9091);
or U10715 (N_10715,N_8348,N_8598);
xor U10716 (N_10716,N_9085,N_9403);
and U10717 (N_10717,N_9893,N_9756);
or U10718 (N_10718,N_8356,N_9460);
xnor U10719 (N_10719,N_8447,N_9396);
or U10720 (N_10720,N_8491,N_8192);
or U10721 (N_10721,N_9752,N_8921);
nor U10722 (N_10722,N_8787,N_9960);
nand U10723 (N_10723,N_9986,N_8163);
nand U10724 (N_10724,N_8751,N_9211);
or U10725 (N_10725,N_9200,N_9479);
nor U10726 (N_10726,N_9555,N_8693);
and U10727 (N_10727,N_9287,N_9702);
nand U10728 (N_10728,N_9887,N_8783);
nor U10729 (N_10729,N_8471,N_9045);
or U10730 (N_10730,N_9426,N_8896);
xnor U10731 (N_10731,N_8357,N_9763);
and U10732 (N_10732,N_9539,N_8835);
and U10733 (N_10733,N_9477,N_9536);
xnor U10734 (N_10734,N_8166,N_8210);
nor U10735 (N_10735,N_9474,N_9612);
or U10736 (N_10736,N_9934,N_9812);
and U10737 (N_10737,N_9735,N_8454);
and U10738 (N_10738,N_8461,N_9969);
xnor U10739 (N_10739,N_8208,N_9814);
xnor U10740 (N_10740,N_8249,N_9890);
and U10741 (N_10741,N_8354,N_9326);
or U10742 (N_10742,N_9495,N_9903);
nand U10743 (N_10743,N_9353,N_8068);
and U10744 (N_10744,N_9876,N_8695);
nand U10745 (N_10745,N_9731,N_8962);
nand U10746 (N_10746,N_8632,N_8881);
or U10747 (N_10747,N_8785,N_9189);
and U10748 (N_10748,N_8227,N_8568);
nor U10749 (N_10749,N_8550,N_8816);
nor U10750 (N_10750,N_9558,N_9161);
xor U10751 (N_10751,N_9502,N_8987);
or U10752 (N_10752,N_8201,N_8998);
and U10753 (N_10753,N_8007,N_8654);
nand U10754 (N_10754,N_9332,N_8817);
nor U10755 (N_10755,N_9399,N_8540);
or U10756 (N_10756,N_9544,N_8669);
xor U10757 (N_10757,N_9390,N_8204);
nand U10758 (N_10758,N_8975,N_9280);
and U10759 (N_10759,N_8190,N_8526);
xnor U10760 (N_10760,N_9099,N_9348);
nand U10761 (N_10761,N_8592,N_8794);
nand U10762 (N_10762,N_8574,N_9074);
xor U10763 (N_10763,N_9213,N_9626);
nor U10764 (N_10764,N_9137,N_8587);
xnor U10765 (N_10765,N_8350,N_9869);
or U10766 (N_10766,N_9722,N_8976);
and U10767 (N_10767,N_9299,N_9543);
or U10768 (N_10768,N_8725,N_9547);
or U10769 (N_10769,N_8053,N_9153);
and U10770 (N_10770,N_8926,N_8552);
nor U10771 (N_10771,N_9152,N_9443);
or U10772 (N_10772,N_8727,N_9204);
nand U10773 (N_10773,N_9023,N_9296);
xor U10774 (N_10774,N_9222,N_9003);
xor U10775 (N_10775,N_9894,N_9561);
nor U10776 (N_10776,N_8993,N_9392);
and U10777 (N_10777,N_9372,N_9101);
and U10778 (N_10778,N_9412,N_9891);
and U10779 (N_10779,N_8861,N_9860);
xor U10780 (N_10780,N_9379,N_8510);
xnor U10781 (N_10781,N_8888,N_9769);
nand U10782 (N_10782,N_9524,N_9926);
xor U10783 (N_10783,N_8286,N_9786);
nor U10784 (N_10784,N_9885,N_8918);
and U10785 (N_10785,N_9063,N_8089);
nor U10786 (N_10786,N_9087,N_8547);
and U10787 (N_10787,N_9264,N_8108);
and U10788 (N_10788,N_9774,N_8331);
nand U10789 (N_10789,N_8917,N_8963);
nor U10790 (N_10790,N_9354,N_9640);
and U10791 (N_10791,N_9072,N_9534);
or U10792 (N_10792,N_9384,N_8745);
or U10793 (N_10793,N_8850,N_8904);
and U10794 (N_10794,N_9818,N_9806);
and U10795 (N_10795,N_8127,N_9892);
or U10796 (N_10796,N_9599,N_8541);
xnor U10797 (N_10797,N_9391,N_9605);
nor U10798 (N_10798,N_8908,N_9194);
and U10799 (N_10799,N_8880,N_9083);
nor U10800 (N_10800,N_9648,N_9261);
or U10801 (N_10801,N_8919,N_9631);
nand U10802 (N_10802,N_9689,N_8205);
and U10803 (N_10803,N_9560,N_9595);
and U10804 (N_10804,N_9282,N_8448);
and U10805 (N_10805,N_9781,N_9839);
or U10806 (N_10806,N_8762,N_8425);
nand U10807 (N_10807,N_9679,N_9577);
or U10808 (N_10808,N_9925,N_8175);
or U10809 (N_10809,N_9066,N_8498);
and U10810 (N_10810,N_9165,N_9684);
and U10811 (N_10811,N_9985,N_8769);
nand U10812 (N_10812,N_9119,N_9465);
or U10813 (N_10813,N_8099,N_9060);
nor U10814 (N_10814,N_9278,N_9487);
or U10815 (N_10815,N_8145,N_8886);
nand U10816 (N_10816,N_8238,N_8157);
nand U10817 (N_10817,N_8656,N_9245);
and U10818 (N_10818,N_9447,N_8776);
nand U10819 (N_10819,N_9142,N_9996);
nor U10820 (N_10820,N_8465,N_9564);
or U10821 (N_10821,N_9962,N_8809);
nand U10822 (N_10822,N_8818,N_8828);
nand U10823 (N_10823,N_8104,N_8426);
or U10824 (N_10824,N_9990,N_8856);
nor U10825 (N_10825,N_8496,N_8805);
and U10826 (N_10826,N_9636,N_9253);
nand U10827 (N_10827,N_8518,N_9709);
xnor U10828 (N_10828,N_8412,N_9012);
and U10829 (N_10829,N_8704,N_9404);
nor U10830 (N_10830,N_9439,N_8245);
or U10831 (N_10831,N_9092,N_9139);
nor U10832 (N_10832,N_8899,N_9330);
and U10833 (N_10833,N_9965,N_9346);
xor U10834 (N_10834,N_8156,N_8929);
nor U10835 (N_10835,N_8548,N_9019);
and U10836 (N_10836,N_9898,N_9145);
nand U10837 (N_10837,N_8343,N_9924);
nand U10838 (N_10838,N_9828,N_8170);
xnor U10839 (N_10839,N_9846,N_9586);
xnor U10840 (N_10840,N_9910,N_8736);
nand U10841 (N_10841,N_8991,N_8040);
xnor U10842 (N_10842,N_9613,N_8290);
and U10843 (N_10843,N_8389,N_8051);
and U10844 (N_10844,N_8311,N_8459);
nor U10845 (N_10845,N_8415,N_8414);
or U10846 (N_10846,N_8102,N_9861);
nor U10847 (N_10847,N_9344,N_9059);
and U10848 (N_10848,N_8832,N_8564);
or U10849 (N_10849,N_9753,N_8014);
nand U10850 (N_10850,N_9401,N_8469);
or U10851 (N_10851,N_9509,N_8588);
or U10852 (N_10852,N_8650,N_9514);
xnor U10853 (N_10853,N_8437,N_8734);
nor U10854 (N_10854,N_8187,N_9627);
nand U10855 (N_10855,N_9714,N_8444);
or U10856 (N_10856,N_9938,N_8646);
nand U10857 (N_10857,N_9456,N_8603);
or U10858 (N_10858,N_8793,N_9840);
or U10859 (N_10859,N_9322,N_8576);
and U10860 (N_10860,N_8316,N_9758);
nor U10861 (N_10861,N_8842,N_9701);
nor U10862 (N_10862,N_9730,N_8811);
nand U10863 (N_10863,N_9170,N_8378);
nor U10864 (N_10864,N_8043,N_9008);
xor U10865 (N_10865,N_9772,N_8213);
and U10866 (N_10866,N_8038,N_8601);
nor U10867 (N_10867,N_8943,N_8823);
nor U10868 (N_10868,N_8457,N_9795);
nor U10869 (N_10869,N_8942,N_8990);
xor U10870 (N_10870,N_9470,N_8293);
and U10871 (N_10871,N_9611,N_8509);
or U10872 (N_10872,N_9179,N_9501);
nor U10873 (N_10873,N_9041,N_9144);
nand U10874 (N_10874,N_9478,N_9491);
nor U10875 (N_10875,N_8685,N_8363);
or U10876 (N_10876,N_8486,N_9844);
or U10877 (N_10877,N_9067,N_9864);
nor U10878 (N_10878,N_8349,N_9250);
nor U10879 (N_10879,N_8042,N_8922);
and U10880 (N_10880,N_8660,N_8719);
xnor U10881 (N_10881,N_9815,N_8015);
nand U10882 (N_10882,N_8168,N_9570);
and U10883 (N_10883,N_8195,N_8892);
nor U10884 (N_10884,N_8622,N_9504);
nor U10885 (N_10885,N_9822,N_8143);
nor U10886 (N_10886,N_9777,N_8327);
and U10887 (N_10887,N_9789,N_9708);
nor U10888 (N_10888,N_8554,N_9765);
xnor U10889 (N_10889,N_9983,N_9056);
nand U10890 (N_10890,N_9109,N_8663);
and U10891 (N_10891,N_9042,N_8398);
and U10892 (N_10892,N_8180,N_8126);
and U10893 (N_10893,N_8100,N_8134);
xor U10894 (N_10894,N_9757,N_8986);
or U10895 (N_10895,N_8006,N_9454);
or U10896 (N_10896,N_9494,N_9336);
nor U10897 (N_10897,N_9190,N_8779);
nand U10898 (N_10898,N_9665,N_9700);
nand U10899 (N_10899,N_9872,N_9151);
nand U10900 (N_10900,N_9005,N_8840);
and U10901 (N_10901,N_9393,N_8534);
and U10902 (N_10902,N_9328,N_9171);
or U10903 (N_10903,N_8557,N_8737);
or U10904 (N_10904,N_9678,N_9333);
nand U10905 (N_10905,N_9138,N_8668);
or U10906 (N_10906,N_9141,N_9386);
or U10907 (N_10907,N_8583,N_8657);
xnor U10908 (N_10908,N_8845,N_8150);
nor U10909 (N_10909,N_9146,N_8684);
and U10910 (N_10910,N_9044,N_9920);
nor U10911 (N_10911,N_8353,N_8928);
and U10912 (N_10912,N_9405,N_8778);
xnor U10913 (N_10913,N_9306,N_8280);
nand U10914 (N_10914,N_9102,N_8490);
nor U10915 (N_10915,N_9221,N_8569);
and U10916 (N_10916,N_8093,N_8218);
nor U10917 (N_10917,N_9174,N_8494);
xor U10918 (N_10918,N_8542,N_8499);
xnor U10919 (N_10919,N_9475,N_8673);
xor U10920 (N_10920,N_8655,N_9819);
nand U10921 (N_10921,N_8383,N_8671);
xnor U10922 (N_10922,N_9075,N_8599);
and U10923 (N_10923,N_8939,N_9522);
or U10924 (N_10924,N_8017,N_8812);
nand U10925 (N_10925,N_9647,N_8185);
and U10926 (N_10926,N_8865,N_8984);
nor U10927 (N_10927,N_9877,N_9778);
nor U10928 (N_10928,N_8369,N_9027);
nor U10929 (N_10929,N_8713,N_9675);
and U10930 (N_10930,N_8985,N_9981);
and U10931 (N_10931,N_8619,N_9901);
and U10932 (N_10932,N_9106,N_9858);
and U10933 (N_10933,N_9309,N_8885);
xor U10934 (N_10934,N_9563,N_9835);
nor U10935 (N_10935,N_8050,N_9219);
nand U10936 (N_10936,N_8691,N_9122);
or U10937 (N_10937,N_9235,N_8667);
nor U10938 (N_10938,N_9382,N_9673);
nor U10939 (N_10939,N_8846,N_8841);
nand U10940 (N_10940,N_9496,N_8831);
and U10941 (N_10941,N_9768,N_8573);
and U10942 (N_10942,N_8958,N_9255);
nand U10943 (N_10943,N_9043,N_8830);
and U10944 (N_10944,N_8920,N_9671);
xnor U10945 (N_10945,N_9879,N_9243);
and U10946 (N_10946,N_8393,N_8744);
nand U10947 (N_10947,N_9476,N_9552);
xnor U10948 (N_10948,N_9550,N_8240);
or U10949 (N_10949,N_8434,N_9016);
nor U10950 (N_10950,N_9149,N_8341);
and U10951 (N_10951,N_9313,N_8957);
or U10952 (N_10952,N_9667,N_8433);
nand U10953 (N_10953,N_8978,N_8791);
or U10954 (N_10954,N_8082,N_9590);
and U10955 (N_10955,N_8149,N_8913);
xor U10956 (N_10956,N_8641,N_8813);
and U10957 (N_10957,N_9663,N_8336);
or U10958 (N_10958,N_8342,N_8317);
nor U10959 (N_10959,N_8367,N_9010);
and U10960 (N_10960,N_8257,N_9999);
or U10961 (N_10961,N_8966,N_8295);
nand U10962 (N_10962,N_9128,N_8796);
or U10963 (N_10963,N_8253,N_8843);
and U10964 (N_10964,N_8462,N_8046);
or U10965 (N_10965,N_9463,N_9402);
nor U10966 (N_10966,N_9389,N_8307);
nor U10967 (N_10967,N_8789,N_8487);
or U10968 (N_10968,N_8273,N_8716);
and U10969 (N_10969,N_9946,N_9307);
xnor U10970 (N_10970,N_8025,N_9997);
nand U10971 (N_10971,N_9214,N_9050);
nor U10972 (N_10972,N_9725,N_8268);
or U10973 (N_10973,N_9298,N_9148);
nand U10974 (N_10974,N_9622,N_9071);
and U10975 (N_10975,N_9295,N_8801);
or U10976 (N_10976,N_8183,N_8648);
and U10977 (N_10977,N_9624,N_8808);
or U10978 (N_10978,N_8875,N_8464);
nand U10979 (N_10979,N_9919,N_8270);
and U10980 (N_10980,N_9070,N_8954);
and U10981 (N_10981,N_9150,N_8429);
and U10982 (N_10982,N_9548,N_8625);
nor U10983 (N_10983,N_9367,N_8413);
nor U10984 (N_10984,N_9423,N_9114);
nand U10985 (N_10985,N_8819,N_8075);
or U10986 (N_10986,N_8752,N_9325);
or U10987 (N_10987,N_8507,N_8700);
xor U10988 (N_10988,N_9339,N_8120);
nor U10989 (N_10989,N_9634,N_9683);
nor U10990 (N_10990,N_8299,N_9176);
nand U10991 (N_10991,N_8221,N_9318);
nor U10992 (N_10992,N_8570,N_9360);
xnor U10993 (N_10993,N_8186,N_8345);
nor U10994 (N_10994,N_8219,N_8364);
nor U10995 (N_10995,N_9793,N_9244);
nand U10996 (N_10996,N_9989,N_8117);
nor U10997 (N_10997,N_9192,N_9281);
nor U10998 (N_10998,N_9263,N_9197);
or U10999 (N_10999,N_9053,N_9842);
nand U11000 (N_11000,N_9168,N_9785);
and U11001 (N_11001,N_8769,N_8952);
or U11002 (N_11002,N_9655,N_9174);
nand U11003 (N_11003,N_8820,N_9524);
nand U11004 (N_11004,N_8799,N_8801);
and U11005 (N_11005,N_8035,N_8678);
or U11006 (N_11006,N_8311,N_8585);
nand U11007 (N_11007,N_9553,N_8447);
nand U11008 (N_11008,N_9259,N_9386);
nor U11009 (N_11009,N_8217,N_9990);
or U11010 (N_11010,N_8921,N_9135);
and U11011 (N_11011,N_9828,N_8083);
and U11012 (N_11012,N_9082,N_9406);
xnor U11013 (N_11013,N_9487,N_8957);
nor U11014 (N_11014,N_8919,N_9766);
and U11015 (N_11015,N_8996,N_9353);
and U11016 (N_11016,N_9828,N_8009);
nand U11017 (N_11017,N_8398,N_9424);
or U11018 (N_11018,N_9759,N_9633);
or U11019 (N_11019,N_8330,N_8451);
nand U11020 (N_11020,N_9856,N_9425);
xnor U11021 (N_11021,N_9030,N_9938);
nor U11022 (N_11022,N_9416,N_8044);
nand U11023 (N_11023,N_8621,N_8681);
nor U11024 (N_11024,N_9102,N_9932);
and U11025 (N_11025,N_8259,N_9072);
xnor U11026 (N_11026,N_8341,N_9104);
nor U11027 (N_11027,N_8253,N_8555);
nor U11028 (N_11028,N_8390,N_9994);
xnor U11029 (N_11029,N_9820,N_8894);
and U11030 (N_11030,N_8078,N_8632);
and U11031 (N_11031,N_8083,N_8943);
and U11032 (N_11032,N_8504,N_8154);
nand U11033 (N_11033,N_8719,N_8847);
nand U11034 (N_11034,N_8693,N_9267);
nor U11035 (N_11035,N_9583,N_8714);
xnor U11036 (N_11036,N_8190,N_9555);
xnor U11037 (N_11037,N_9941,N_9177);
and U11038 (N_11038,N_9251,N_9331);
or U11039 (N_11039,N_8324,N_9957);
and U11040 (N_11040,N_9907,N_9949);
xnor U11041 (N_11041,N_9787,N_9271);
and U11042 (N_11042,N_8423,N_8656);
nor U11043 (N_11043,N_8419,N_8985);
xor U11044 (N_11044,N_9148,N_8375);
or U11045 (N_11045,N_9831,N_8597);
nand U11046 (N_11046,N_8969,N_8012);
xnor U11047 (N_11047,N_9493,N_9566);
nand U11048 (N_11048,N_8838,N_8325);
nor U11049 (N_11049,N_8202,N_9859);
and U11050 (N_11050,N_9787,N_9994);
xnor U11051 (N_11051,N_8922,N_9903);
xor U11052 (N_11052,N_8496,N_8790);
nor U11053 (N_11053,N_9291,N_8645);
xor U11054 (N_11054,N_9654,N_9901);
nand U11055 (N_11055,N_9295,N_9499);
nor U11056 (N_11056,N_9348,N_9919);
nand U11057 (N_11057,N_8621,N_9185);
or U11058 (N_11058,N_8680,N_8969);
xor U11059 (N_11059,N_8540,N_9546);
nor U11060 (N_11060,N_9043,N_8639);
xor U11061 (N_11061,N_8017,N_8273);
nor U11062 (N_11062,N_8357,N_9504);
and U11063 (N_11063,N_8347,N_9705);
xor U11064 (N_11064,N_9519,N_8706);
xnor U11065 (N_11065,N_9945,N_9147);
nand U11066 (N_11066,N_8326,N_9085);
and U11067 (N_11067,N_9126,N_8883);
nor U11068 (N_11068,N_8453,N_8020);
nor U11069 (N_11069,N_9481,N_9781);
xnor U11070 (N_11070,N_9365,N_9863);
nand U11071 (N_11071,N_8712,N_9921);
or U11072 (N_11072,N_8098,N_8175);
xnor U11073 (N_11073,N_9819,N_8489);
xor U11074 (N_11074,N_9358,N_8916);
and U11075 (N_11075,N_9136,N_8635);
xnor U11076 (N_11076,N_8353,N_9313);
xnor U11077 (N_11077,N_9013,N_9455);
or U11078 (N_11078,N_8267,N_9603);
or U11079 (N_11079,N_8396,N_8208);
xor U11080 (N_11080,N_8593,N_9847);
or U11081 (N_11081,N_8027,N_8384);
nand U11082 (N_11082,N_8353,N_9072);
nand U11083 (N_11083,N_8999,N_9392);
and U11084 (N_11084,N_8900,N_9598);
nor U11085 (N_11085,N_9603,N_8339);
and U11086 (N_11086,N_8889,N_9736);
xor U11087 (N_11087,N_9353,N_8428);
and U11088 (N_11088,N_8161,N_9017);
and U11089 (N_11089,N_9162,N_9308);
xor U11090 (N_11090,N_9761,N_9704);
or U11091 (N_11091,N_8865,N_8014);
or U11092 (N_11092,N_8126,N_8555);
nor U11093 (N_11093,N_8120,N_9875);
and U11094 (N_11094,N_9161,N_8196);
or U11095 (N_11095,N_8612,N_9498);
nor U11096 (N_11096,N_8087,N_8701);
or U11097 (N_11097,N_9671,N_9567);
or U11098 (N_11098,N_9041,N_8016);
nor U11099 (N_11099,N_8283,N_9875);
xor U11100 (N_11100,N_8676,N_8286);
nor U11101 (N_11101,N_9033,N_9441);
nand U11102 (N_11102,N_9432,N_8436);
and U11103 (N_11103,N_9324,N_8083);
and U11104 (N_11104,N_8274,N_8628);
xor U11105 (N_11105,N_8511,N_9075);
or U11106 (N_11106,N_8132,N_8501);
and U11107 (N_11107,N_9784,N_9770);
xor U11108 (N_11108,N_8749,N_9790);
and U11109 (N_11109,N_8325,N_8947);
or U11110 (N_11110,N_9967,N_8819);
xnor U11111 (N_11111,N_8127,N_9832);
nand U11112 (N_11112,N_9397,N_9038);
nand U11113 (N_11113,N_9516,N_9561);
xnor U11114 (N_11114,N_8578,N_9678);
xnor U11115 (N_11115,N_8460,N_8068);
nand U11116 (N_11116,N_9548,N_8057);
xor U11117 (N_11117,N_9691,N_9883);
xnor U11118 (N_11118,N_8089,N_8567);
nand U11119 (N_11119,N_8655,N_8200);
xnor U11120 (N_11120,N_8976,N_9213);
and U11121 (N_11121,N_8500,N_8945);
xnor U11122 (N_11122,N_8980,N_9147);
or U11123 (N_11123,N_9825,N_9307);
or U11124 (N_11124,N_8451,N_8270);
nand U11125 (N_11125,N_9901,N_8841);
and U11126 (N_11126,N_8785,N_9305);
nand U11127 (N_11127,N_8402,N_9801);
nand U11128 (N_11128,N_9497,N_9973);
nand U11129 (N_11129,N_9501,N_8163);
and U11130 (N_11130,N_8210,N_9292);
nor U11131 (N_11131,N_9701,N_9275);
or U11132 (N_11132,N_9594,N_8717);
and U11133 (N_11133,N_8216,N_9669);
nor U11134 (N_11134,N_9304,N_9238);
nor U11135 (N_11135,N_8007,N_9276);
and U11136 (N_11136,N_9629,N_8413);
nand U11137 (N_11137,N_8530,N_8131);
or U11138 (N_11138,N_8932,N_8514);
nand U11139 (N_11139,N_8583,N_8702);
nor U11140 (N_11140,N_9803,N_9810);
and U11141 (N_11141,N_8094,N_9217);
or U11142 (N_11142,N_9088,N_9318);
nor U11143 (N_11143,N_9778,N_8781);
nand U11144 (N_11144,N_9898,N_8370);
nor U11145 (N_11145,N_9375,N_8478);
nor U11146 (N_11146,N_9095,N_9724);
nor U11147 (N_11147,N_8225,N_9397);
and U11148 (N_11148,N_8552,N_8883);
or U11149 (N_11149,N_8677,N_8702);
xnor U11150 (N_11150,N_8744,N_8855);
xnor U11151 (N_11151,N_9399,N_9988);
nor U11152 (N_11152,N_9657,N_9750);
xor U11153 (N_11153,N_8132,N_9914);
or U11154 (N_11154,N_8594,N_8938);
or U11155 (N_11155,N_8678,N_8238);
or U11156 (N_11156,N_9765,N_8728);
nand U11157 (N_11157,N_8631,N_9536);
and U11158 (N_11158,N_8006,N_9536);
nand U11159 (N_11159,N_8751,N_9920);
and U11160 (N_11160,N_9455,N_9446);
and U11161 (N_11161,N_9844,N_9577);
nand U11162 (N_11162,N_8072,N_9202);
xnor U11163 (N_11163,N_9936,N_8702);
or U11164 (N_11164,N_9689,N_9079);
or U11165 (N_11165,N_8844,N_9240);
nand U11166 (N_11166,N_8452,N_8073);
xnor U11167 (N_11167,N_8864,N_9630);
nand U11168 (N_11168,N_8183,N_8788);
and U11169 (N_11169,N_8134,N_9794);
nor U11170 (N_11170,N_9077,N_9958);
or U11171 (N_11171,N_9369,N_9072);
nand U11172 (N_11172,N_9943,N_8958);
nand U11173 (N_11173,N_8973,N_8789);
nor U11174 (N_11174,N_9053,N_8373);
nand U11175 (N_11175,N_8370,N_8396);
or U11176 (N_11176,N_8912,N_9429);
or U11177 (N_11177,N_9355,N_8784);
nor U11178 (N_11178,N_9181,N_8719);
xnor U11179 (N_11179,N_8939,N_8161);
and U11180 (N_11180,N_8677,N_9810);
nand U11181 (N_11181,N_8633,N_9036);
nand U11182 (N_11182,N_8371,N_8695);
nand U11183 (N_11183,N_9256,N_9701);
or U11184 (N_11184,N_9198,N_9399);
nand U11185 (N_11185,N_9137,N_9070);
and U11186 (N_11186,N_9927,N_9864);
or U11187 (N_11187,N_8555,N_8200);
nor U11188 (N_11188,N_9902,N_9827);
nand U11189 (N_11189,N_8799,N_8691);
nor U11190 (N_11190,N_8403,N_9550);
xor U11191 (N_11191,N_9377,N_8123);
or U11192 (N_11192,N_9475,N_8384);
or U11193 (N_11193,N_8666,N_9907);
xnor U11194 (N_11194,N_9387,N_9891);
nor U11195 (N_11195,N_9969,N_8624);
nor U11196 (N_11196,N_8556,N_9873);
and U11197 (N_11197,N_9798,N_9663);
or U11198 (N_11198,N_9562,N_8008);
or U11199 (N_11199,N_8763,N_9616);
and U11200 (N_11200,N_8614,N_8950);
or U11201 (N_11201,N_9629,N_8120);
nor U11202 (N_11202,N_8671,N_9053);
xnor U11203 (N_11203,N_9527,N_9788);
nand U11204 (N_11204,N_9322,N_9811);
nand U11205 (N_11205,N_9328,N_9422);
nor U11206 (N_11206,N_9340,N_8876);
nor U11207 (N_11207,N_9479,N_9634);
nor U11208 (N_11208,N_8770,N_8992);
or U11209 (N_11209,N_8049,N_9336);
and U11210 (N_11210,N_8151,N_8749);
xnor U11211 (N_11211,N_8918,N_8493);
or U11212 (N_11212,N_8484,N_8464);
nor U11213 (N_11213,N_9020,N_9092);
and U11214 (N_11214,N_9325,N_9618);
xnor U11215 (N_11215,N_9708,N_8902);
xor U11216 (N_11216,N_9881,N_9364);
xor U11217 (N_11217,N_8145,N_9362);
or U11218 (N_11218,N_9949,N_9201);
xor U11219 (N_11219,N_8077,N_8232);
and U11220 (N_11220,N_8838,N_8110);
xor U11221 (N_11221,N_8025,N_9620);
xnor U11222 (N_11222,N_9566,N_8277);
nor U11223 (N_11223,N_8880,N_9222);
and U11224 (N_11224,N_9959,N_9673);
and U11225 (N_11225,N_8901,N_8808);
nand U11226 (N_11226,N_8716,N_9083);
xnor U11227 (N_11227,N_8160,N_9781);
or U11228 (N_11228,N_9047,N_8851);
and U11229 (N_11229,N_8377,N_9633);
xor U11230 (N_11230,N_8764,N_9259);
xor U11231 (N_11231,N_9700,N_9790);
and U11232 (N_11232,N_8008,N_8780);
or U11233 (N_11233,N_8039,N_9421);
nor U11234 (N_11234,N_8450,N_9267);
nor U11235 (N_11235,N_9375,N_8162);
nand U11236 (N_11236,N_9100,N_9813);
and U11237 (N_11237,N_9037,N_8894);
or U11238 (N_11238,N_9286,N_9354);
or U11239 (N_11239,N_8991,N_8709);
nor U11240 (N_11240,N_8373,N_8990);
nor U11241 (N_11241,N_8210,N_9033);
nand U11242 (N_11242,N_8104,N_8547);
and U11243 (N_11243,N_9373,N_8941);
nor U11244 (N_11244,N_9527,N_8997);
and U11245 (N_11245,N_8499,N_8187);
and U11246 (N_11246,N_8457,N_8242);
or U11247 (N_11247,N_8050,N_8484);
nor U11248 (N_11248,N_8301,N_8779);
nor U11249 (N_11249,N_9517,N_8285);
and U11250 (N_11250,N_9225,N_9851);
nor U11251 (N_11251,N_8552,N_8708);
xor U11252 (N_11252,N_8754,N_9277);
and U11253 (N_11253,N_9297,N_8686);
xor U11254 (N_11254,N_9833,N_9102);
nor U11255 (N_11255,N_9833,N_9287);
nor U11256 (N_11256,N_8803,N_8147);
or U11257 (N_11257,N_9336,N_8002);
nand U11258 (N_11258,N_8256,N_8359);
or U11259 (N_11259,N_8811,N_8939);
nor U11260 (N_11260,N_8013,N_8908);
nand U11261 (N_11261,N_8999,N_9363);
xnor U11262 (N_11262,N_8475,N_9514);
nor U11263 (N_11263,N_8570,N_9509);
and U11264 (N_11264,N_9817,N_9649);
nand U11265 (N_11265,N_8942,N_8462);
xnor U11266 (N_11266,N_9196,N_8154);
nand U11267 (N_11267,N_8949,N_8730);
and U11268 (N_11268,N_8380,N_9545);
xnor U11269 (N_11269,N_9413,N_8070);
and U11270 (N_11270,N_9750,N_8313);
nor U11271 (N_11271,N_8215,N_9305);
nor U11272 (N_11272,N_9311,N_8223);
and U11273 (N_11273,N_8021,N_9951);
nor U11274 (N_11274,N_9443,N_8161);
nor U11275 (N_11275,N_9390,N_9152);
nor U11276 (N_11276,N_8640,N_9219);
xor U11277 (N_11277,N_8055,N_8590);
and U11278 (N_11278,N_9815,N_9797);
or U11279 (N_11279,N_9398,N_9850);
nand U11280 (N_11280,N_8078,N_9453);
xnor U11281 (N_11281,N_9391,N_9342);
nand U11282 (N_11282,N_9900,N_9806);
xnor U11283 (N_11283,N_8504,N_9863);
nand U11284 (N_11284,N_9546,N_9430);
or U11285 (N_11285,N_9935,N_8847);
xor U11286 (N_11286,N_9114,N_9886);
nand U11287 (N_11287,N_8120,N_8523);
nor U11288 (N_11288,N_8286,N_9766);
or U11289 (N_11289,N_9339,N_8591);
or U11290 (N_11290,N_8904,N_8049);
nand U11291 (N_11291,N_8414,N_8837);
and U11292 (N_11292,N_9117,N_9620);
nand U11293 (N_11293,N_8740,N_9323);
nor U11294 (N_11294,N_8287,N_8398);
or U11295 (N_11295,N_9911,N_8379);
nor U11296 (N_11296,N_8018,N_9154);
and U11297 (N_11297,N_9761,N_9139);
and U11298 (N_11298,N_8587,N_8863);
or U11299 (N_11299,N_8891,N_9968);
xnor U11300 (N_11300,N_8159,N_9638);
nor U11301 (N_11301,N_8616,N_9568);
nor U11302 (N_11302,N_9589,N_9788);
xnor U11303 (N_11303,N_9354,N_8310);
nor U11304 (N_11304,N_8244,N_9910);
or U11305 (N_11305,N_9506,N_9516);
nand U11306 (N_11306,N_8442,N_8777);
or U11307 (N_11307,N_8788,N_8002);
xor U11308 (N_11308,N_9664,N_9076);
xnor U11309 (N_11309,N_8527,N_9272);
nand U11310 (N_11310,N_8744,N_9521);
nor U11311 (N_11311,N_8987,N_9332);
nor U11312 (N_11312,N_9769,N_8887);
nand U11313 (N_11313,N_9343,N_8998);
or U11314 (N_11314,N_9825,N_9872);
or U11315 (N_11315,N_8257,N_8438);
nor U11316 (N_11316,N_8922,N_9218);
or U11317 (N_11317,N_9473,N_9785);
nand U11318 (N_11318,N_8109,N_8495);
or U11319 (N_11319,N_9865,N_9338);
and U11320 (N_11320,N_9840,N_8086);
or U11321 (N_11321,N_9694,N_8491);
or U11322 (N_11322,N_8256,N_8110);
xnor U11323 (N_11323,N_9218,N_8145);
or U11324 (N_11324,N_8292,N_9679);
and U11325 (N_11325,N_8497,N_8103);
nand U11326 (N_11326,N_9159,N_9941);
nor U11327 (N_11327,N_8650,N_9961);
xor U11328 (N_11328,N_9230,N_9125);
and U11329 (N_11329,N_8992,N_8911);
or U11330 (N_11330,N_9067,N_8313);
or U11331 (N_11331,N_9528,N_8889);
and U11332 (N_11332,N_9488,N_9931);
nand U11333 (N_11333,N_9215,N_8947);
nor U11334 (N_11334,N_8008,N_9472);
nand U11335 (N_11335,N_9658,N_8354);
nor U11336 (N_11336,N_9248,N_9477);
and U11337 (N_11337,N_8267,N_9064);
xor U11338 (N_11338,N_8325,N_9929);
and U11339 (N_11339,N_9518,N_9588);
nand U11340 (N_11340,N_9966,N_9854);
nand U11341 (N_11341,N_8651,N_9040);
or U11342 (N_11342,N_8400,N_9030);
and U11343 (N_11343,N_9883,N_8627);
xor U11344 (N_11344,N_9161,N_9825);
or U11345 (N_11345,N_8685,N_8657);
or U11346 (N_11346,N_8601,N_8314);
and U11347 (N_11347,N_9403,N_9858);
or U11348 (N_11348,N_9241,N_8073);
and U11349 (N_11349,N_8082,N_8146);
and U11350 (N_11350,N_9810,N_9528);
xor U11351 (N_11351,N_8957,N_9378);
or U11352 (N_11352,N_8565,N_8139);
nand U11353 (N_11353,N_8491,N_9494);
xor U11354 (N_11354,N_9859,N_9693);
xor U11355 (N_11355,N_8763,N_9852);
nand U11356 (N_11356,N_9756,N_9899);
xnor U11357 (N_11357,N_8192,N_8917);
xnor U11358 (N_11358,N_8040,N_8113);
nor U11359 (N_11359,N_8082,N_8480);
nor U11360 (N_11360,N_8283,N_8528);
xnor U11361 (N_11361,N_8191,N_9725);
nand U11362 (N_11362,N_8581,N_8432);
nor U11363 (N_11363,N_9468,N_8051);
and U11364 (N_11364,N_9222,N_8009);
nand U11365 (N_11365,N_9014,N_9064);
or U11366 (N_11366,N_9562,N_8690);
xor U11367 (N_11367,N_8240,N_8193);
or U11368 (N_11368,N_9799,N_9278);
or U11369 (N_11369,N_8527,N_9788);
nand U11370 (N_11370,N_9197,N_8934);
and U11371 (N_11371,N_8413,N_9183);
nand U11372 (N_11372,N_9980,N_9939);
nand U11373 (N_11373,N_8231,N_8475);
xor U11374 (N_11374,N_8257,N_8516);
and U11375 (N_11375,N_9030,N_9953);
and U11376 (N_11376,N_8030,N_8172);
nor U11377 (N_11377,N_9501,N_8759);
and U11378 (N_11378,N_8476,N_8288);
nor U11379 (N_11379,N_9299,N_9346);
nor U11380 (N_11380,N_8685,N_8871);
nand U11381 (N_11381,N_9392,N_9288);
nor U11382 (N_11382,N_8855,N_8979);
xor U11383 (N_11383,N_8780,N_8611);
xnor U11384 (N_11384,N_9918,N_9569);
nand U11385 (N_11385,N_9689,N_8496);
and U11386 (N_11386,N_9289,N_9038);
nand U11387 (N_11387,N_8387,N_8145);
xor U11388 (N_11388,N_8636,N_8787);
nor U11389 (N_11389,N_8635,N_9359);
and U11390 (N_11390,N_8345,N_9522);
and U11391 (N_11391,N_9686,N_8565);
and U11392 (N_11392,N_9050,N_9889);
xor U11393 (N_11393,N_8100,N_8114);
nor U11394 (N_11394,N_9739,N_8385);
nand U11395 (N_11395,N_9032,N_8798);
and U11396 (N_11396,N_8453,N_8560);
nand U11397 (N_11397,N_9701,N_8315);
and U11398 (N_11398,N_8974,N_8593);
and U11399 (N_11399,N_9729,N_8129);
or U11400 (N_11400,N_9134,N_9612);
nand U11401 (N_11401,N_9525,N_8275);
nor U11402 (N_11402,N_9901,N_8722);
or U11403 (N_11403,N_9558,N_9480);
xnor U11404 (N_11404,N_8915,N_9489);
nand U11405 (N_11405,N_9464,N_9676);
xnor U11406 (N_11406,N_9911,N_8294);
nand U11407 (N_11407,N_8193,N_8495);
nor U11408 (N_11408,N_9504,N_8439);
xor U11409 (N_11409,N_8201,N_9199);
xnor U11410 (N_11410,N_8554,N_9505);
nor U11411 (N_11411,N_8071,N_9477);
xnor U11412 (N_11412,N_8258,N_8910);
nand U11413 (N_11413,N_9975,N_9776);
nor U11414 (N_11414,N_8343,N_8568);
and U11415 (N_11415,N_9176,N_9571);
and U11416 (N_11416,N_9410,N_9552);
nand U11417 (N_11417,N_9681,N_8295);
xnor U11418 (N_11418,N_9507,N_8461);
or U11419 (N_11419,N_9965,N_9166);
xnor U11420 (N_11420,N_9903,N_8726);
or U11421 (N_11421,N_9769,N_9026);
or U11422 (N_11422,N_8321,N_9758);
nand U11423 (N_11423,N_8714,N_9219);
and U11424 (N_11424,N_8564,N_8350);
xnor U11425 (N_11425,N_9277,N_9640);
xnor U11426 (N_11426,N_8694,N_9281);
nor U11427 (N_11427,N_8393,N_9161);
and U11428 (N_11428,N_8655,N_8580);
xnor U11429 (N_11429,N_8734,N_8388);
nor U11430 (N_11430,N_9698,N_8792);
nand U11431 (N_11431,N_8942,N_9135);
nor U11432 (N_11432,N_9381,N_9308);
xor U11433 (N_11433,N_8088,N_9567);
or U11434 (N_11434,N_9312,N_9567);
and U11435 (N_11435,N_9909,N_8195);
or U11436 (N_11436,N_9253,N_8651);
and U11437 (N_11437,N_9083,N_9697);
nand U11438 (N_11438,N_8722,N_8099);
xor U11439 (N_11439,N_9022,N_8769);
nor U11440 (N_11440,N_8301,N_8836);
nor U11441 (N_11441,N_8414,N_8560);
nor U11442 (N_11442,N_8046,N_9357);
nand U11443 (N_11443,N_9840,N_9614);
or U11444 (N_11444,N_8319,N_9371);
nor U11445 (N_11445,N_8182,N_8161);
nor U11446 (N_11446,N_8369,N_9120);
or U11447 (N_11447,N_9871,N_8632);
xnor U11448 (N_11448,N_9303,N_9719);
and U11449 (N_11449,N_8671,N_8260);
xnor U11450 (N_11450,N_8732,N_9937);
xnor U11451 (N_11451,N_9412,N_8303);
and U11452 (N_11452,N_8298,N_8035);
and U11453 (N_11453,N_8631,N_9643);
or U11454 (N_11454,N_8205,N_9838);
nand U11455 (N_11455,N_8994,N_8950);
nor U11456 (N_11456,N_9492,N_9313);
xor U11457 (N_11457,N_8711,N_9877);
nand U11458 (N_11458,N_9904,N_9686);
xor U11459 (N_11459,N_9614,N_8256);
and U11460 (N_11460,N_8621,N_9387);
and U11461 (N_11461,N_8417,N_8636);
nor U11462 (N_11462,N_8797,N_9769);
nor U11463 (N_11463,N_8329,N_9193);
or U11464 (N_11464,N_9807,N_9788);
nor U11465 (N_11465,N_9515,N_8650);
xor U11466 (N_11466,N_9159,N_9725);
nor U11467 (N_11467,N_9436,N_9722);
and U11468 (N_11468,N_8743,N_9895);
or U11469 (N_11469,N_8587,N_8160);
nand U11470 (N_11470,N_8655,N_9714);
or U11471 (N_11471,N_9016,N_9093);
nor U11472 (N_11472,N_8755,N_8664);
xor U11473 (N_11473,N_9286,N_9274);
xnor U11474 (N_11474,N_9743,N_9593);
xnor U11475 (N_11475,N_9845,N_9691);
or U11476 (N_11476,N_9189,N_9972);
or U11477 (N_11477,N_9587,N_8291);
xnor U11478 (N_11478,N_8044,N_9964);
nand U11479 (N_11479,N_9300,N_9556);
nor U11480 (N_11480,N_9347,N_8545);
nor U11481 (N_11481,N_9448,N_9998);
nand U11482 (N_11482,N_8992,N_8983);
nor U11483 (N_11483,N_8153,N_8097);
and U11484 (N_11484,N_8014,N_9023);
nor U11485 (N_11485,N_9692,N_9289);
xnor U11486 (N_11486,N_9885,N_8629);
or U11487 (N_11487,N_9199,N_9200);
nand U11488 (N_11488,N_8705,N_9840);
xnor U11489 (N_11489,N_9312,N_9331);
nand U11490 (N_11490,N_8728,N_9532);
and U11491 (N_11491,N_8373,N_9543);
nor U11492 (N_11492,N_8081,N_9563);
and U11493 (N_11493,N_8350,N_8381);
nor U11494 (N_11494,N_9288,N_9547);
nor U11495 (N_11495,N_9956,N_9634);
nand U11496 (N_11496,N_8279,N_9725);
nand U11497 (N_11497,N_8378,N_9380);
nor U11498 (N_11498,N_8764,N_8687);
or U11499 (N_11499,N_8614,N_8745);
nand U11500 (N_11500,N_9538,N_8592);
or U11501 (N_11501,N_8857,N_8257);
or U11502 (N_11502,N_9352,N_8641);
nor U11503 (N_11503,N_8479,N_8343);
xnor U11504 (N_11504,N_9637,N_8138);
nor U11505 (N_11505,N_8313,N_9127);
xnor U11506 (N_11506,N_8976,N_8019);
and U11507 (N_11507,N_9748,N_8764);
xnor U11508 (N_11508,N_8514,N_8505);
xnor U11509 (N_11509,N_9798,N_9719);
xor U11510 (N_11510,N_9940,N_9974);
or U11511 (N_11511,N_9242,N_8245);
or U11512 (N_11512,N_8506,N_8851);
and U11513 (N_11513,N_9022,N_8391);
xnor U11514 (N_11514,N_9332,N_8654);
xnor U11515 (N_11515,N_9985,N_9366);
or U11516 (N_11516,N_8941,N_9881);
and U11517 (N_11517,N_8655,N_9416);
nand U11518 (N_11518,N_8241,N_8256);
xnor U11519 (N_11519,N_8007,N_8254);
nor U11520 (N_11520,N_8086,N_9996);
nor U11521 (N_11521,N_9125,N_8201);
xor U11522 (N_11522,N_9723,N_9119);
nor U11523 (N_11523,N_9595,N_8934);
nand U11524 (N_11524,N_9285,N_8400);
xnor U11525 (N_11525,N_9954,N_8842);
xor U11526 (N_11526,N_8091,N_9324);
xnor U11527 (N_11527,N_8503,N_8673);
and U11528 (N_11528,N_8228,N_9346);
nor U11529 (N_11529,N_9936,N_8137);
or U11530 (N_11530,N_9891,N_9714);
xor U11531 (N_11531,N_9112,N_9947);
nand U11532 (N_11532,N_8261,N_8782);
and U11533 (N_11533,N_9636,N_8159);
and U11534 (N_11534,N_8090,N_9516);
and U11535 (N_11535,N_8580,N_9358);
nand U11536 (N_11536,N_8145,N_9723);
nand U11537 (N_11537,N_8164,N_9127);
or U11538 (N_11538,N_8837,N_9256);
and U11539 (N_11539,N_8935,N_9076);
xnor U11540 (N_11540,N_8755,N_9197);
nor U11541 (N_11541,N_8834,N_9658);
nor U11542 (N_11542,N_8626,N_8186);
and U11543 (N_11543,N_8586,N_8631);
nor U11544 (N_11544,N_8918,N_9261);
xor U11545 (N_11545,N_8980,N_9980);
xnor U11546 (N_11546,N_8701,N_8912);
nand U11547 (N_11547,N_9850,N_9827);
xor U11548 (N_11548,N_9965,N_9083);
nand U11549 (N_11549,N_8918,N_8225);
and U11550 (N_11550,N_9483,N_9576);
xor U11551 (N_11551,N_8691,N_8436);
and U11552 (N_11552,N_9362,N_9844);
and U11553 (N_11553,N_8625,N_8325);
nand U11554 (N_11554,N_8339,N_9221);
nor U11555 (N_11555,N_8040,N_8653);
xor U11556 (N_11556,N_8393,N_9748);
and U11557 (N_11557,N_8444,N_9701);
and U11558 (N_11558,N_9843,N_9395);
and U11559 (N_11559,N_9434,N_8494);
nor U11560 (N_11560,N_8124,N_9229);
or U11561 (N_11561,N_9593,N_9566);
nor U11562 (N_11562,N_9088,N_8629);
or U11563 (N_11563,N_9264,N_9312);
xor U11564 (N_11564,N_9204,N_8830);
xnor U11565 (N_11565,N_9970,N_9609);
and U11566 (N_11566,N_8438,N_8804);
xor U11567 (N_11567,N_9691,N_8719);
nor U11568 (N_11568,N_8001,N_8547);
nand U11569 (N_11569,N_8552,N_9803);
nand U11570 (N_11570,N_9371,N_8331);
xnor U11571 (N_11571,N_8887,N_9326);
nand U11572 (N_11572,N_9519,N_9237);
nand U11573 (N_11573,N_9100,N_9103);
and U11574 (N_11574,N_8520,N_8705);
or U11575 (N_11575,N_9169,N_8369);
xnor U11576 (N_11576,N_9065,N_9883);
or U11577 (N_11577,N_8697,N_9432);
or U11578 (N_11578,N_8886,N_9911);
or U11579 (N_11579,N_8125,N_8098);
nand U11580 (N_11580,N_9001,N_8929);
xor U11581 (N_11581,N_9223,N_8776);
nor U11582 (N_11582,N_8162,N_9644);
nand U11583 (N_11583,N_9201,N_8482);
nand U11584 (N_11584,N_8673,N_9245);
or U11585 (N_11585,N_8071,N_8108);
xnor U11586 (N_11586,N_9475,N_9840);
and U11587 (N_11587,N_8864,N_8282);
nor U11588 (N_11588,N_9643,N_9485);
nor U11589 (N_11589,N_8168,N_8247);
or U11590 (N_11590,N_9196,N_8467);
nand U11591 (N_11591,N_8571,N_9367);
nand U11592 (N_11592,N_8776,N_8285);
xnor U11593 (N_11593,N_8870,N_9586);
and U11594 (N_11594,N_8817,N_9985);
nor U11595 (N_11595,N_8757,N_8331);
or U11596 (N_11596,N_8353,N_9152);
nor U11597 (N_11597,N_8433,N_9475);
or U11598 (N_11598,N_8871,N_9467);
and U11599 (N_11599,N_9476,N_8422);
or U11600 (N_11600,N_9850,N_9134);
or U11601 (N_11601,N_9616,N_9798);
and U11602 (N_11602,N_8577,N_8975);
xnor U11603 (N_11603,N_8981,N_9385);
nand U11604 (N_11604,N_9518,N_9573);
nand U11605 (N_11605,N_9613,N_9539);
or U11606 (N_11606,N_8985,N_8718);
and U11607 (N_11607,N_9102,N_8617);
or U11608 (N_11608,N_8640,N_8804);
nand U11609 (N_11609,N_9576,N_9223);
or U11610 (N_11610,N_8327,N_8918);
or U11611 (N_11611,N_9969,N_9063);
or U11612 (N_11612,N_9065,N_9271);
nor U11613 (N_11613,N_9138,N_9455);
and U11614 (N_11614,N_8650,N_8060);
or U11615 (N_11615,N_8372,N_8360);
xnor U11616 (N_11616,N_8576,N_8605);
nand U11617 (N_11617,N_8007,N_8915);
and U11618 (N_11618,N_8353,N_9543);
nor U11619 (N_11619,N_9447,N_8616);
and U11620 (N_11620,N_9957,N_8261);
nor U11621 (N_11621,N_9105,N_8674);
nand U11622 (N_11622,N_9081,N_8850);
nand U11623 (N_11623,N_9782,N_9892);
xor U11624 (N_11624,N_8151,N_9547);
nor U11625 (N_11625,N_9968,N_8156);
or U11626 (N_11626,N_9789,N_9138);
xnor U11627 (N_11627,N_9596,N_8712);
xnor U11628 (N_11628,N_9659,N_9821);
nor U11629 (N_11629,N_8790,N_8635);
nand U11630 (N_11630,N_8544,N_9097);
and U11631 (N_11631,N_9255,N_9984);
and U11632 (N_11632,N_8216,N_8944);
xor U11633 (N_11633,N_8785,N_8218);
nor U11634 (N_11634,N_9256,N_9342);
nand U11635 (N_11635,N_8488,N_9003);
nand U11636 (N_11636,N_9815,N_9696);
xnor U11637 (N_11637,N_9405,N_8652);
or U11638 (N_11638,N_9203,N_8457);
nor U11639 (N_11639,N_8148,N_9239);
and U11640 (N_11640,N_9778,N_8581);
or U11641 (N_11641,N_8681,N_8187);
nor U11642 (N_11642,N_9679,N_8389);
xor U11643 (N_11643,N_8306,N_8434);
nor U11644 (N_11644,N_8862,N_9754);
or U11645 (N_11645,N_9489,N_9633);
xnor U11646 (N_11646,N_8505,N_9092);
nor U11647 (N_11647,N_8244,N_8003);
or U11648 (N_11648,N_9590,N_8859);
nor U11649 (N_11649,N_8921,N_9632);
nand U11650 (N_11650,N_9676,N_9097);
nand U11651 (N_11651,N_8344,N_9183);
and U11652 (N_11652,N_8123,N_9086);
and U11653 (N_11653,N_9255,N_9926);
and U11654 (N_11654,N_9440,N_9202);
xnor U11655 (N_11655,N_8432,N_9355);
xnor U11656 (N_11656,N_9386,N_8380);
or U11657 (N_11657,N_8502,N_8127);
nand U11658 (N_11658,N_8158,N_9882);
xor U11659 (N_11659,N_9376,N_8895);
or U11660 (N_11660,N_9290,N_8141);
or U11661 (N_11661,N_8092,N_9174);
or U11662 (N_11662,N_9601,N_9402);
or U11663 (N_11663,N_9910,N_9345);
nand U11664 (N_11664,N_9693,N_9931);
xnor U11665 (N_11665,N_8992,N_8440);
and U11666 (N_11666,N_8792,N_8425);
nor U11667 (N_11667,N_9884,N_8954);
nand U11668 (N_11668,N_8215,N_9849);
nor U11669 (N_11669,N_8747,N_8899);
and U11670 (N_11670,N_8479,N_8708);
nor U11671 (N_11671,N_9996,N_8180);
nand U11672 (N_11672,N_9378,N_9489);
or U11673 (N_11673,N_9184,N_9481);
xnor U11674 (N_11674,N_8834,N_9710);
or U11675 (N_11675,N_9762,N_9939);
and U11676 (N_11676,N_8974,N_8645);
and U11677 (N_11677,N_8993,N_9636);
or U11678 (N_11678,N_8739,N_8763);
xor U11679 (N_11679,N_9898,N_8448);
nor U11680 (N_11680,N_9401,N_8848);
or U11681 (N_11681,N_8292,N_8394);
xor U11682 (N_11682,N_8498,N_9091);
or U11683 (N_11683,N_9356,N_8004);
nor U11684 (N_11684,N_9710,N_9716);
nor U11685 (N_11685,N_8021,N_8251);
and U11686 (N_11686,N_9875,N_9305);
or U11687 (N_11687,N_9190,N_9545);
nand U11688 (N_11688,N_8739,N_8382);
nand U11689 (N_11689,N_8947,N_9531);
nor U11690 (N_11690,N_9501,N_9572);
or U11691 (N_11691,N_9867,N_9984);
nor U11692 (N_11692,N_9367,N_9591);
nand U11693 (N_11693,N_9761,N_9350);
nor U11694 (N_11694,N_9695,N_8968);
nor U11695 (N_11695,N_9349,N_8232);
xor U11696 (N_11696,N_9016,N_9886);
nor U11697 (N_11697,N_9638,N_8138);
or U11698 (N_11698,N_9321,N_9319);
xnor U11699 (N_11699,N_9736,N_9314);
nor U11700 (N_11700,N_8672,N_8404);
nor U11701 (N_11701,N_8461,N_9773);
xnor U11702 (N_11702,N_9035,N_9269);
or U11703 (N_11703,N_9333,N_8189);
nor U11704 (N_11704,N_9638,N_9755);
xor U11705 (N_11705,N_8442,N_9145);
nor U11706 (N_11706,N_9547,N_8970);
nand U11707 (N_11707,N_9981,N_9784);
nor U11708 (N_11708,N_8898,N_8890);
and U11709 (N_11709,N_8685,N_8938);
xor U11710 (N_11710,N_8661,N_8909);
xnor U11711 (N_11711,N_9969,N_9500);
nand U11712 (N_11712,N_9801,N_8368);
and U11713 (N_11713,N_9872,N_8063);
and U11714 (N_11714,N_9568,N_9834);
or U11715 (N_11715,N_9259,N_9142);
nor U11716 (N_11716,N_9399,N_9539);
xnor U11717 (N_11717,N_9515,N_8165);
nor U11718 (N_11718,N_9923,N_8045);
and U11719 (N_11719,N_9679,N_8272);
nor U11720 (N_11720,N_8188,N_9857);
xor U11721 (N_11721,N_9743,N_9941);
xor U11722 (N_11722,N_8778,N_8761);
or U11723 (N_11723,N_8090,N_9204);
and U11724 (N_11724,N_9759,N_9304);
xor U11725 (N_11725,N_8614,N_9510);
nor U11726 (N_11726,N_9590,N_8853);
nor U11727 (N_11727,N_9963,N_8351);
or U11728 (N_11728,N_9874,N_9168);
xnor U11729 (N_11729,N_8066,N_8105);
xor U11730 (N_11730,N_8399,N_9672);
and U11731 (N_11731,N_9098,N_8709);
nand U11732 (N_11732,N_9656,N_9355);
and U11733 (N_11733,N_8872,N_8771);
and U11734 (N_11734,N_9337,N_9825);
nand U11735 (N_11735,N_8654,N_9407);
xnor U11736 (N_11736,N_9459,N_9387);
nor U11737 (N_11737,N_8841,N_8024);
and U11738 (N_11738,N_8812,N_9338);
xnor U11739 (N_11739,N_8828,N_9165);
nand U11740 (N_11740,N_8173,N_8529);
nand U11741 (N_11741,N_9803,N_8144);
nand U11742 (N_11742,N_8752,N_8894);
nor U11743 (N_11743,N_8052,N_8525);
nor U11744 (N_11744,N_9862,N_8550);
xor U11745 (N_11745,N_8483,N_8284);
or U11746 (N_11746,N_9971,N_9249);
or U11747 (N_11747,N_9220,N_8528);
nand U11748 (N_11748,N_9103,N_8206);
or U11749 (N_11749,N_9678,N_8940);
nand U11750 (N_11750,N_8634,N_8068);
and U11751 (N_11751,N_9061,N_9947);
nand U11752 (N_11752,N_8649,N_8278);
nand U11753 (N_11753,N_9907,N_9459);
nand U11754 (N_11754,N_8139,N_9238);
nand U11755 (N_11755,N_8244,N_9453);
nand U11756 (N_11756,N_8013,N_8395);
nor U11757 (N_11757,N_8902,N_9476);
nor U11758 (N_11758,N_9941,N_8847);
or U11759 (N_11759,N_9381,N_8816);
xnor U11760 (N_11760,N_8012,N_9341);
nand U11761 (N_11761,N_8497,N_9026);
and U11762 (N_11762,N_9585,N_9964);
or U11763 (N_11763,N_8385,N_8462);
xnor U11764 (N_11764,N_8062,N_9476);
and U11765 (N_11765,N_9737,N_9325);
xor U11766 (N_11766,N_9732,N_8233);
xor U11767 (N_11767,N_8518,N_8865);
or U11768 (N_11768,N_9253,N_8460);
nand U11769 (N_11769,N_9946,N_8768);
or U11770 (N_11770,N_9808,N_8655);
xor U11771 (N_11771,N_9145,N_9991);
or U11772 (N_11772,N_9487,N_9614);
or U11773 (N_11773,N_9181,N_8359);
nand U11774 (N_11774,N_8639,N_8430);
nor U11775 (N_11775,N_8958,N_9847);
and U11776 (N_11776,N_8239,N_9033);
xor U11777 (N_11777,N_8758,N_8487);
xnor U11778 (N_11778,N_8205,N_8643);
nor U11779 (N_11779,N_9658,N_9199);
nor U11780 (N_11780,N_8891,N_8300);
nor U11781 (N_11781,N_9262,N_9737);
xor U11782 (N_11782,N_8048,N_9126);
and U11783 (N_11783,N_8195,N_9561);
xnor U11784 (N_11784,N_8213,N_9150);
nand U11785 (N_11785,N_8337,N_8108);
nor U11786 (N_11786,N_9854,N_9554);
or U11787 (N_11787,N_8445,N_8669);
nor U11788 (N_11788,N_8311,N_8536);
nor U11789 (N_11789,N_9670,N_8446);
xnor U11790 (N_11790,N_9900,N_9930);
xor U11791 (N_11791,N_8171,N_8302);
or U11792 (N_11792,N_8850,N_9475);
or U11793 (N_11793,N_9371,N_8676);
xor U11794 (N_11794,N_8491,N_8642);
nor U11795 (N_11795,N_8859,N_8879);
and U11796 (N_11796,N_9846,N_9351);
or U11797 (N_11797,N_9173,N_9371);
or U11798 (N_11798,N_9252,N_9057);
and U11799 (N_11799,N_8302,N_8055);
nand U11800 (N_11800,N_8849,N_9499);
nand U11801 (N_11801,N_8380,N_9749);
nor U11802 (N_11802,N_9065,N_9305);
nor U11803 (N_11803,N_9053,N_9756);
xnor U11804 (N_11804,N_9083,N_9107);
nor U11805 (N_11805,N_8021,N_9457);
nand U11806 (N_11806,N_9707,N_9883);
and U11807 (N_11807,N_8888,N_8847);
nand U11808 (N_11808,N_8106,N_8619);
nor U11809 (N_11809,N_9551,N_8204);
and U11810 (N_11810,N_9649,N_8848);
or U11811 (N_11811,N_9721,N_8261);
and U11812 (N_11812,N_9869,N_8057);
and U11813 (N_11813,N_8942,N_9513);
and U11814 (N_11814,N_9429,N_8893);
nor U11815 (N_11815,N_8866,N_9903);
nand U11816 (N_11816,N_8765,N_9896);
nand U11817 (N_11817,N_9214,N_9789);
or U11818 (N_11818,N_8383,N_9496);
and U11819 (N_11819,N_8820,N_8724);
or U11820 (N_11820,N_8764,N_8697);
xnor U11821 (N_11821,N_8057,N_9913);
or U11822 (N_11822,N_9540,N_8970);
nor U11823 (N_11823,N_9080,N_8261);
and U11824 (N_11824,N_8530,N_8730);
or U11825 (N_11825,N_8010,N_8755);
nand U11826 (N_11826,N_8292,N_9670);
nand U11827 (N_11827,N_9327,N_8398);
nor U11828 (N_11828,N_9640,N_8369);
xor U11829 (N_11829,N_9310,N_8759);
and U11830 (N_11830,N_9567,N_8943);
nand U11831 (N_11831,N_9264,N_9272);
xor U11832 (N_11832,N_8852,N_8637);
or U11833 (N_11833,N_8134,N_9731);
nor U11834 (N_11834,N_8457,N_8839);
and U11835 (N_11835,N_9777,N_9391);
and U11836 (N_11836,N_9701,N_9678);
or U11837 (N_11837,N_9826,N_9324);
xnor U11838 (N_11838,N_9951,N_9644);
nand U11839 (N_11839,N_8330,N_9444);
nor U11840 (N_11840,N_9817,N_9701);
nand U11841 (N_11841,N_9583,N_9466);
or U11842 (N_11842,N_8358,N_8632);
nor U11843 (N_11843,N_8340,N_9451);
and U11844 (N_11844,N_8717,N_8321);
nand U11845 (N_11845,N_9203,N_8164);
or U11846 (N_11846,N_8945,N_8594);
xnor U11847 (N_11847,N_8621,N_9359);
and U11848 (N_11848,N_8576,N_8052);
nand U11849 (N_11849,N_9366,N_8046);
xnor U11850 (N_11850,N_9426,N_9138);
nor U11851 (N_11851,N_9952,N_8803);
or U11852 (N_11852,N_8446,N_8353);
nor U11853 (N_11853,N_9733,N_9914);
or U11854 (N_11854,N_9459,N_8601);
or U11855 (N_11855,N_9488,N_9775);
or U11856 (N_11856,N_8912,N_9263);
xor U11857 (N_11857,N_8609,N_9042);
xnor U11858 (N_11858,N_9350,N_9628);
nand U11859 (N_11859,N_9724,N_8345);
nor U11860 (N_11860,N_9030,N_8661);
nand U11861 (N_11861,N_9339,N_8781);
nor U11862 (N_11862,N_8163,N_8276);
nand U11863 (N_11863,N_8769,N_8687);
or U11864 (N_11864,N_8478,N_9930);
nor U11865 (N_11865,N_9387,N_8509);
xnor U11866 (N_11866,N_8537,N_9138);
nor U11867 (N_11867,N_8713,N_8761);
nor U11868 (N_11868,N_8466,N_8114);
nand U11869 (N_11869,N_9229,N_9053);
nor U11870 (N_11870,N_9565,N_9690);
or U11871 (N_11871,N_9751,N_8799);
xor U11872 (N_11872,N_9110,N_8947);
and U11873 (N_11873,N_9335,N_9010);
and U11874 (N_11874,N_8849,N_9884);
nor U11875 (N_11875,N_9095,N_9345);
nand U11876 (N_11876,N_8248,N_9471);
nor U11877 (N_11877,N_9334,N_8671);
or U11878 (N_11878,N_8630,N_8301);
and U11879 (N_11879,N_9060,N_9479);
and U11880 (N_11880,N_8319,N_9134);
or U11881 (N_11881,N_8921,N_8311);
nand U11882 (N_11882,N_8650,N_8980);
nand U11883 (N_11883,N_8256,N_9107);
and U11884 (N_11884,N_9470,N_8215);
nand U11885 (N_11885,N_9417,N_8496);
nand U11886 (N_11886,N_8455,N_9242);
or U11887 (N_11887,N_9478,N_8446);
xor U11888 (N_11888,N_8997,N_9001);
xnor U11889 (N_11889,N_9435,N_8375);
xor U11890 (N_11890,N_8277,N_9045);
nand U11891 (N_11891,N_9279,N_9835);
nand U11892 (N_11892,N_8466,N_8041);
or U11893 (N_11893,N_9636,N_9399);
or U11894 (N_11894,N_9635,N_8836);
or U11895 (N_11895,N_8314,N_9035);
or U11896 (N_11896,N_8844,N_9563);
and U11897 (N_11897,N_9347,N_9434);
xnor U11898 (N_11898,N_8845,N_8696);
or U11899 (N_11899,N_9580,N_8357);
xor U11900 (N_11900,N_8885,N_8449);
and U11901 (N_11901,N_8098,N_9903);
xor U11902 (N_11902,N_9293,N_9911);
xnor U11903 (N_11903,N_8771,N_8429);
xnor U11904 (N_11904,N_9954,N_9730);
and U11905 (N_11905,N_9454,N_9240);
and U11906 (N_11906,N_8191,N_9145);
nor U11907 (N_11907,N_9498,N_9693);
nand U11908 (N_11908,N_9019,N_8203);
and U11909 (N_11909,N_8572,N_8200);
nand U11910 (N_11910,N_9400,N_8267);
and U11911 (N_11911,N_9084,N_8897);
nand U11912 (N_11912,N_8753,N_8005);
xor U11913 (N_11913,N_8973,N_8170);
and U11914 (N_11914,N_8844,N_9666);
or U11915 (N_11915,N_9228,N_9643);
and U11916 (N_11916,N_8220,N_8352);
nand U11917 (N_11917,N_8909,N_8106);
xnor U11918 (N_11918,N_9566,N_8197);
nand U11919 (N_11919,N_8295,N_9400);
xnor U11920 (N_11920,N_8112,N_8519);
or U11921 (N_11921,N_8066,N_8633);
nor U11922 (N_11922,N_8566,N_9412);
or U11923 (N_11923,N_9787,N_8842);
and U11924 (N_11924,N_8524,N_8658);
nor U11925 (N_11925,N_9153,N_8220);
nor U11926 (N_11926,N_8466,N_9587);
and U11927 (N_11927,N_9317,N_8641);
nor U11928 (N_11928,N_9469,N_8570);
and U11929 (N_11929,N_9168,N_8781);
or U11930 (N_11930,N_9609,N_8140);
xnor U11931 (N_11931,N_9054,N_8374);
xnor U11932 (N_11932,N_9890,N_8617);
and U11933 (N_11933,N_9261,N_8532);
xnor U11934 (N_11934,N_8824,N_8028);
or U11935 (N_11935,N_8900,N_8492);
nand U11936 (N_11936,N_8729,N_8803);
nand U11937 (N_11937,N_9026,N_9567);
nand U11938 (N_11938,N_8979,N_8431);
or U11939 (N_11939,N_9502,N_9752);
nor U11940 (N_11940,N_8336,N_9492);
nand U11941 (N_11941,N_9346,N_9343);
nand U11942 (N_11942,N_9635,N_9412);
or U11943 (N_11943,N_8101,N_9386);
and U11944 (N_11944,N_8671,N_9813);
xnor U11945 (N_11945,N_8335,N_8462);
or U11946 (N_11946,N_9416,N_8000);
and U11947 (N_11947,N_9272,N_8135);
nand U11948 (N_11948,N_9647,N_8291);
and U11949 (N_11949,N_8546,N_9444);
or U11950 (N_11950,N_8311,N_9129);
or U11951 (N_11951,N_9484,N_9451);
and U11952 (N_11952,N_8180,N_8882);
nand U11953 (N_11953,N_8512,N_8381);
and U11954 (N_11954,N_8386,N_8487);
nor U11955 (N_11955,N_8395,N_8267);
or U11956 (N_11956,N_8503,N_8359);
xnor U11957 (N_11957,N_9389,N_8964);
xnor U11958 (N_11958,N_8958,N_9836);
nand U11959 (N_11959,N_9839,N_9975);
xnor U11960 (N_11960,N_9049,N_8110);
xor U11961 (N_11961,N_9316,N_8827);
or U11962 (N_11962,N_9656,N_8800);
xor U11963 (N_11963,N_8845,N_8253);
nor U11964 (N_11964,N_9295,N_8132);
nor U11965 (N_11965,N_9276,N_9186);
nor U11966 (N_11966,N_8856,N_8252);
or U11967 (N_11967,N_8039,N_8458);
or U11968 (N_11968,N_9137,N_8798);
and U11969 (N_11969,N_9263,N_8306);
xor U11970 (N_11970,N_8622,N_8283);
nand U11971 (N_11971,N_8780,N_8142);
nand U11972 (N_11972,N_9646,N_8383);
and U11973 (N_11973,N_9323,N_9609);
or U11974 (N_11974,N_9144,N_9019);
and U11975 (N_11975,N_8593,N_9191);
nand U11976 (N_11976,N_8819,N_8461);
or U11977 (N_11977,N_9613,N_9056);
nand U11978 (N_11978,N_8961,N_8169);
nor U11979 (N_11979,N_9485,N_8924);
or U11980 (N_11980,N_9532,N_8009);
or U11981 (N_11981,N_8036,N_9871);
and U11982 (N_11982,N_8725,N_8931);
nand U11983 (N_11983,N_9803,N_9817);
nor U11984 (N_11984,N_9114,N_8083);
or U11985 (N_11985,N_8448,N_9320);
nand U11986 (N_11986,N_8552,N_9006);
xnor U11987 (N_11987,N_8530,N_9221);
xor U11988 (N_11988,N_8517,N_8486);
xor U11989 (N_11989,N_8264,N_8233);
nor U11990 (N_11990,N_9725,N_9019);
or U11991 (N_11991,N_9392,N_8564);
or U11992 (N_11992,N_9835,N_9029);
nor U11993 (N_11993,N_8563,N_9894);
nand U11994 (N_11994,N_8112,N_8348);
nand U11995 (N_11995,N_9409,N_9787);
or U11996 (N_11996,N_8957,N_9242);
nand U11997 (N_11997,N_9443,N_9386);
nor U11998 (N_11998,N_9495,N_9398);
and U11999 (N_11999,N_8345,N_9780);
nand U12000 (N_12000,N_11907,N_10507);
or U12001 (N_12001,N_11733,N_10462);
or U12002 (N_12002,N_10206,N_10993);
nand U12003 (N_12003,N_11843,N_10465);
xnor U12004 (N_12004,N_11928,N_11629);
xor U12005 (N_12005,N_10457,N_10094);
or U12006 (N_12006,N_10105,N_10558);
xnor U12007 (N_12007,N_10724,N_11701);
xnor U12008 (N_12008,N_10021,N_10381);
and U12009 (N_12009,N_10464,N_11477);
and U12010 (N_12010,N_10446,N_10124);
and U12011 (N_12011,N_10132,N_10324);
nor U12012 (N_12012,N_10005,N_10807);
xor U12013 (N_12013,N_10916,N_10732);
xnor U12014 (N_12014,N_11746,N_10871);
or U12015 (N_12015,N_11908,N_11302);
and U12016 (N_12016,N_11898,N_11094);
nor U12017 (N_12017,N_10991,N_11541);
or U12018 (N_12018,N_11974,N_10809);
xnor U12019 (N_12019,N_11820,N_10880);
and U12020 (N_12020,N_10628,N_11841);
xnor U12021 (N_12021,N_10263,N_11053);
or U12022 (N_12022,N_11529,N_10624);
or U12023 (N_12023,N_11487,N_11555);
xor U12024 (N_12024,N_10163,N_11805);
and U12025 (N_12025,N_11246,N_10606);
nand U12026 (N_12026,N_10625,N_11848);
or U12027 (N_12027,N_11750,N_10986);
nand U12028 (N_12028,N_10047,N_10503);
nand U12029 (N_12029,N_11222,N_11773);
nand U12030 (N_12030,N_10716,N_11622);
and U12031 (N_12031,N_11258,N_11400);
nor U12032 (N_12032,N_10221,N_11927);
or U12033 (N_12033,N_10403,N_10755);
nor U12034 (N_12034,N_11207,N_11424);
xor U12035 (N_12035,N_11786,N_10605);
nand U12036 (N_12036,N_10333,N_11602);
nand U12037 (N_12037,N_10265,N_11252);
xnor U12038 (N_12038,N_11531,N_11788);
xnor U12039 (N_12039,N_11236,N_10758);
or U12040 (N_12040,N_10033,N_10424);
xnor U12041 (N_12041,N_11539,N_11705);
or U12042 (N_12042,N_10839,N_10767);
and U12043 (N_12043,N_10795,N_11544);
or U12044 (N_12044,N_11017,N_11772);
nand U12045 (N_12045,N_11620,N_11725);
xnor U12046 (N_12046,N_10821,N_10996);
nor U12047 (N_12047,N_11552,N_11003);
nand U12048 (N_12048,N_11692,N_10869);
nand U12049 (N_12049,N_11727,N_11918);
nor U12050 (N_12050,N_10121,N_10523);
nor U12051 (N_12051,N_11914,N_10659);
and U12052 (N_12052,N_10228,N_10521);
xor U12053 (N_12053,N_10886,N_11981);
nand U12054 (N_12054,N_10301,N_11693);
and U12055 (N_12055,N_11376,N_11334);
xor U12056 (N_12056,N_11663,N_10579);
nor U12057 (N_12057,N_10917,N_10475);
xnor U12058 (N_12058,N_10452,N_11426);
and U12059 (N_12059,N_10385,N_11808);
xor U12060 (N_12060,N_11203,N_10212);
and U12061 (N_12061,N_11036,N_11512);
nor U12062 (N_12062,N_10834,N_10331);
nor U12063 (N_12063,N_10406,N_10812);
or U12064 (N_12064,N_11495,N_11975);
or U12065 (N_12065,N_11489,N_11888);
xnor U12066 (N_12066,N_10499,N_10925);
or U12067 (N_12067,N_11642,N_11110);
nor U12068 (N_12068,N_11174,N_10494);
or U12069 (N_12069,N_11357,N_10567);
or U12070 (N_12070,N_10610,N_10425);
nor U12071 (N_12071,N_11165,N_10972);
or U12072 (N_12072,N_11880,N_10289);
xor U12073 (N_12073,N_10750,N_11994);
nand U12074 (N_12074,N_10747,N_10438);
nand U12075 (N_12075,N_11086,N_11016);
nor U12076 (N_12076,N_10046,N_11675);
or U12077 (N_12077,N_10942,N_11151);
and U12078 (N_12078,N_10654,N_10007);
nand U12079 (N_12079,N_10737,N_11483);
and U12080 (N_12080,N_11121,N_10118);
nand U12081 (N_12081,N_10547,N_10820);
and U12082 (N_12082,N_10527,N_10687);
and U12083 (N_12083,N_10208,N_11149);
and U12084 (N_12084,N_11333,N_10211);
nand U12085 (N_12085,N_11083,N_10017);
nand U12086 (N_12086,N_10949,N_11319);
nand U12087 (N_12087,N_10231,N_11902);
nand U12088 (N_12088,N_11726,N_10634);
nor U12089 (N_12089,N_10364,N_11795);
nand U12090 (N_12090,N_11241,N_11300);
nand U12091 (N_12091,N_10893,N_10290);
and U12092 (N_12092,N_11837,N_11474);
and U12093 (N_12093,N_10116,N_11636);
xor U12094 (N_12094,N_10883,N_11396);
or U12095 (N_12095,N_10128,N_10770);
nand U12096 (N_12096,N_10690,N_11591);
xor U12097 (N_12097,N_10371,N_11811);
xor U12098 (N_12098,N_10775,N_10491);
or U12099 (N_12099,N_11368,N_10146);
nand U12100 (N_12100,N_10341,N_10517);
or U12101 (N_12101,N_10911,N_10298);
nor U12102 (N_12102,N_10978,N_11522);
xor U12103 (N_12103,N_10794,N_11467);
nand U12104 (N_12104,N_10431,N_11488);
nand U12105 (N_12105,N_10565,N_10485);
xor U12106 (N_12106,N_11815,N_11961);
nand U12107 (N_12107,N_10902,N_10885);
nor U12108 (N_12108,N_10343,N_10003);
or U12109 (N_12109,N_10010,N_11128);
and U12110 (N_12110,N_10781,N_10941);
and U12111 (N_12111,N_10751,N_11369);
xnor U12112 (N_12112,N_11669,N_10059);
nor U12113 (N_12113,N_10850,N_11690);
or U12114 (N_12114,N_11264,N_10651);
or U12115 (N_12115,N_11090,N_11910);
nor U12116 (N_12116,N_11077,N_10276);
and U12117 (N_12117,N_11113,N_11991);
and U12118 (N_12118,N_10546,N_10748);
or U12119 (N_12119,N_10102,N_11001);
and U12120 (N_12120,N_10673,N_11569);
nand U12121 (N_12121,N_10736,N_10246);
and U12122 (N_12122,N_11678,N_10185);
xnor U12123 (N_12123,N_10359,N_11890);
or U12124 (N_12124,N_10952,N_11243);
nor U12125 (N_12125,N_11188,N_10387);
and U12126 (N_12126,N_11519,N_11904);
and U12127 (N_12127,N_10209,N_10609);
nor U12128 (N_12128,N_10989,N_11406);
xnor U12129 (N_12129,N_11643,N_10603);
xnor U12130 (N_12130,N_10951,N_10488);
and U12131 (N_12131,N_10216,N_10837);
xnor U12132 (N_12132,N_11574,N_11760);
nand U12133 (N_12133,N_11419,N_10778);
and U12134 (N_12134,N_10137,N_10598);
nor U12135 (N_12135,N_10113,N_11123);
or U12136 (N_12136,N_10934,N_10159);
xnor U12137 (N_12137,N_10308,N_11307);
and U12138 (N_12138,N_11491,N_11784);
or U12139 (N_12139,N_11955,N_10374);
xnor U12140 (N_12140,N_10420,N_10715);
nor U12141 (N_12141,N_10513,N_11440);
xor U12142 (N_12142,N_10819,N_10486);
and U12143 (N_12143,N_11109,N_10316);
and U12144 (N_12144,N_10099,N_10366);
xor U12145 (N_12145,N_11015,N_10490);
or U12146 (N_12146,N_10427,N_10608);
xnor U12147 (N_12147,N_11422,N_10468);
or U12148 (N_12148,N_10518,N_10245);
and U12149 (N_12149,N_11193,N_10064);
and U12150 (N_12150,N_10484,N_11458);
xor U12151 (N_12151,N_10631,N_11482);
nor U12152 (N_12152,N_10461,N_11798);
nand U12153 (N_12153,N_10866,N_11685);
and U12154 (N_12154,N_10337,N_11562);
nand U12155 (N_12155,N_11377,N_10958);
or U12156 (N_12156,N_11176,N_11306);
or U12157 (N_12157,N_10740,N_11713);
nor U12158 (N_12158,N_10764,N_11381);
or U12159 (N_12159,N_11220,N_11271);
nand U12160 (N_12160,N_11660,N_10671);
or U12161 (N_12161,N_11657,N_11018);
or U12162 (N_12162,N_11803,N_11799);
and U12163 (N_12163,N_10140,N_11510);
nand U12164 (N_12164,N_10847,N_11765);
and U12165 (N_12165,N_11249,N_10145);
or U12166 (N_12166,N_10285,N_11796);
and U12167 (N_12167,N_10418,N_11136);
or U12168 (N_12168,N_10127,N_11409);
nor U12169 (N_12169,N_10342,N_10573);
nor U12170 (N_12170,N_11330,N_10432);
nor U12171 (N_12171,N_11164,N_10478);
nand U12172 (N_12172,N_11343,N_11738);
nor U12173 (N_12173,N_10087,N_10583);
nand U12174 (N_12174,N_10607,N_10796);
or U12175 (N_12175,N_11091,N_10858);
and U12176 (N_12176,N_11704,N_11610);
nor U12177 (N_12177,N_11038,N_10882);
xor U12178 (N_12178,N_11321,N_10260);
or U12179 (N_12179,N_11156,N_11431);
xnor U12180 (N_12180,N_10828,N_11792);
or U12181 (N_12181,N_10313,N_11163);
or U12182 (N_12182,N_11697,N_11944);
nand U12183 (N_12183,N_10063,N_11980);
nor U12184 (N_12184,N_10879,N_11049);
and U12185 (N_12185,N_11239,N_11534);
xor U12186 (N_12186,N_10372,N_11852);
xor U12187 (N_12187,N_11374,N_11118);
and U12188 (N_12188,N_11768,N_10469);
or U12189 (N_12189,N_10838,N_10562);
or U12190 (N_12190,N_11990,N_10509);
nand U12191 (N_12191,N_10780,N_11976);
and U12192 (N_12192,N_10162,N_10340);
or U12193 (N_12193,N_10901,N_11178);
and U12194 (N_12194,N_10470,N_11171);
xnor U12195 (N_12195,N_11635,N_10346);
nand U12196 (N_12196,N_11715,N_11004);
nand U12197 (N_12197,N_11948,N_11854);
nand U12198 (N_12198,N_11548,N_11402);
nand U12199 (N_12199,N_11836,N_10103);
nand U12200 (N_12200,N_10810,N_11702);
and U12201 (N_12201,N_10864,N_10237);
or U12202 (N_12202,N_10542,N_10540);
nand U12203 (N_12203,N_10918,N_10225);
or U12204 (N_12204,N_10709,N_11305);
xnor U12205 (N_12205,N_11470,N_10139);
nor U12206 (N_12206,N_11331,N_11199);
and U12207 (N_12207,N_11339,N_11162);
nand U12208 (N_12208,N_11835,N_10990);
nor U12209 (N_12209,N_10330,N_10173);
nand U12210 (N_12210,N_10066,N_10070);
xor U12211 (N_12211,N_10293,N_10122);
and U12212 (N_12212,N_10806,N_10629);
and U12213 (N_12213,N_11966,N_11380);
and U12214 (N_12214,N_10199,N_10440);
or U12215 (N_12215,N_11245,N_11443);
or U12216 (N_12216,N_11957,N_11652);
and U12217 (N_12217,N_11528,N_10197);
nor U12218 (N_12218,N_10296,N_11871);
or U12219 (N_12219,N_10480,N_10338);
or U12220 (N_12220,N_11045,N_10236);
and U12221 (N_12221,N_10247,N_11082);
or U12222 (N_12222,N_10600,N_10319);
and U12223 (N_12223,N_10620,N_10919);
nand U12224 (N_12224,N_11417,N_11352);
and U12225 (N_12225,N_11340,N_10528);
or U12226 (N_12226,N_11523,N_10531);
nor U12227 (N_12227,N_11168,N_10179);
xor U12228 (N_12228,N_10943,N_10114);
nand U12229 (N_12229,N_10912,N_10852);
nor U12230 (N_12230,N_10039,N_10450);
nand U12231 (N_12231,N_11979,N_11047);
nor U12232 (N_12232,N_11497,N_10404);
xor U12233 (N_12233,N_10594,N_11439);
or U12234 (N_12234,N_11362,N_10008);
and U12235 (N_12235,N_11219,N_10048);
nor U12236 (N_12236,N_10135,N_10648);
xnor U12237 (N_12237,N_10653,N_11311);
nand U12238 (N_12238,N_11614,N_11509);
and U12239 (N_12239,N_11063,N_10312);
and U12240 (N_12240,N_10699,N_10970);
nor U12241 (N_12241,N_11926,N_11596);
nand U12242 (N_12242,N_11297,N_11893);
nand U12243 (N_12243,N_11457,N_10138);
nand U12244 (N_12244,N_11612,N_11924);
and U12245 (N_12245,N_10933,N_11274);
xor U12246 (N_12246,N_11929,N_11679);
nor U12247 (N_12247,N_10756,N_11290);
or U12248 (N_12248,N_11378,N_11498);
and U12249 (N_12249,N_10092,N_11496);
xnor U12250 (N_12250,N_11185,N_11956);
nand U12251 (N_12251,N_10870,N_10028);
nand U12252 (N_12252,N_11338,N_10790);
nand U12253 (N_12253,N_11181,N_10449);
or U12254 (N_12254,N_11647,N_10924);
or U12255 (N_12255,N_10339,N_10156);
nand U12256 (N_12256,N_10906,N_10602);
nand U12257 (N_12257,N_11998,N_10823);
nor U12258 (N_12258,N_10123,N_11335);
and U12259 (N_12259,N_11283,N_10131);
xor U12260 (N_12260,N_10905,N_10353);
or U12261 (N_12261,N_10686,N_10347);
or U12262 (N_12262,N_11999,N_10550);
and U12263 (N_12263,N_10935,N_10031);
nor U12264 (N_12264,N_10076,N_10639);
and U12265 (N_12265,N_11205,N_11351);
nor U12266 (N_12266,N_11711,N_11767);
nand U12267 (N_12267,N_11588,N_10705);
or U12268 (N_12268,N_10940,N_10282);
xnor U12269 (N_12269,N_11317,N_10712);
nor U12270 (N_12270,N_11579,N_10900);
nand U12271 (N_12271,N_10155,N_10698);
and U12272 (N_12272,N_11279,N_11724);
and U12273 (N_12273,N_10963,N_10115);
or U12274 (N_12274,N_10956,N_10255);
or U12275 (N_12275,N_11664,N_11213);
nand U12276 (N_12276,N_11742,N_10323);
nand U12277 (N_12277,N_11587,N_10174);
and U12278 (N_12278,N_10741,N_10233);
xnor U12279 (N_12279,N_11833,N_10477);
xnor U12280 (N_12280,N_10899,N_10154);
nand U12281 (N_12281,N_10825,N_11446);
nand U12282 (N_12282,N_10520,N_11326);
nand U12283 (N_12283,N_10204,N_10969);
and U12284 (N_12284,N_11353,N_10412);
or U12285 (N_12285,N_11631,N_10896);
and U12286 (N_12286,N_10904,N_11556);
xor U12287 (N_12287,N_11229,N_11624);
or U12288 (N_12288,N_10694,N_11560);
xnor U12289 (N_12289,N_11609,N_11076);
xor U12290 (N_12290,N_11824,N_11584);
or U12291 (N_12291,N_11896,N_11081);
or U12292 (N_12292,N_10797,N_10081);
and U12293 (N_12293,N_11709,N_11885);
nor U12294 (N_12294,N_10168,N_10926);
nand U12295 (N_12295,N_10665,N_10352);
and U12296 (N_12296,N_11456,N_10393);
xor U12297 (N_12297,N_11138,N_11056);
or U12298 (N_12298,N_11722,N_11284);
and U12299 (N_12299,N_10130,N_10306);
xnor U12300 (N_12300,N_11859,N_10612);
nor U12301 (N_12301,N_11410,N_11397);
or U12302 (N_12302,N_10239,N_10095);
nor U12303 (N_12303,N_11559,N_11449);
nor U12304 (N_12304,N_11000,N_11484);
or U12305 (N_12305,N_10774,N_10459);
xnor U12306 (N_12306,N_11251,N_10026);
xnor U12307 (N_12307,N_11698,N_11242);
nor U12308 (N_12308,N_10368,N_11169);
or U12309 (N_12309,N_11743,N_11723);
and U12310 (N_12310,N_10569,N_10971);
or U12311 (N_12311,N_10332,N_11382);
or U12312 (N_12312,N_11364,N_10277);
and U12313 (N_12313,N_11348,N_11350);
nor U12314 (N_12314,N_10416,N_10844);
and U12315 (N_12315,N_10792,N_11987);
nor U12316 (N_12316,N_11891,N_11571);
nand U12317 (N_12317,N_10083,N_10647);
and U12318 (N_12318,N_11776,N_11206);
nor U12319 (N_12319,N_10541,N_10230);
xor U12320 (N_12320,N_10058,N_10545);
nand U12321 (N_12321,N_11684,N_10321);
nor U12322 (N_12322,N_10358,N_11448);
xnor U12323 (N_12323,N_10638,N_10614);
nand U12324 (N_12324,N_11389,N_11821);
nand U12325 (N_12325,N_11847,N_11375);
nand U12326 (N_12326,N_10077,N_11009);
or U12327 (N_12327,N_11810,N_11876);
xor U12328 (N_12328,N_11800,N_11184);
or U12329 (N_12329,N_11007,N_10800);
nand U12330 (N_12330,N_10143,N_10184);
or U12331 (N_12331,N_10281,N_10407);
nand U12332 (N_12332,N_11144,N_11195);
or U12333 (N_12333,N_11802,N_10336);
xnor U12334 (N_12334,N_10006,N_10254);
xor U12335 (N_12335,N_11593,N_11407);
or U12336 (N_12336,N_10695,N_11313);
xor U12337 (N_12337,N_11575,N_11041);
or U12338 (N_12338,N_10836,N_11517);
xnor U12339 (N_12339,N_11674,N_10738);
xnor U12340 (N_12340,N_10318,N_11740);
or U12341 (N_12341,N_10663,N_11565);
or U12342 (N_12342,N_10273,N_11347);
nor U12343 (N_12343,N_11813,N_10742);
xor U12344 (N_12344,N_11666,N_10240);
xor U12345 (N_12345,N_11756,N_11633);
and U12346 (N_12346,N_10746,N_10067);
or U12347 (N_12347,N_10129,N_10326);
or U12348 (N_12348,N_10670,N_11244);
xnor U12349 (N_12349,N_11526,N_11322);
nor U12350 (N_12350,N_10098,N_10965);
or U12351 (N_12351,N_11586,N_11842);
or U12352 (N_12352,N_10884,N_11710);
nand U12353 (N_12353,N_10061,N_10731);
xnor U12354 (N_12354,N_10030,N_11993);
or U12355 (N_12355,N_10717,N_11884);
nand U12356 (N_12356,N_10219,N_11233);
or U12357 (N_12357,N_10691,N_10708);
xor U12358 (N_12358,N_11754,N_11774);
or U12359 (N_12359,N_10198,N_11167);
xnor U12360 (N_12360,N_11900,N_11256);
and U12361 (N_12361,N_10314,N_10560);
xnor U12362 (N_12362,N_10682,N_10055);
or U12363 (N_12363,N_10250,N_10120);
xor U12364 (N_12364,N_11459,N_10726);
or U12365 (N_12365,N_11892,N_10530);
nor U12366 (N_12366,N_10481,N_11327);
nor U12367 (N_12367,N_11235,N_11114);
nor U12368 (N_12368,N_10053,N_11515);
xnor U12369 (N_12369,N_10291,N_11019);
nor U12370 (N_12370,N_11816,N_11255);
or U12371 (N_12371,N_10954,N_10423);
xnor U12372 (N_12372,N_11425,N_11518);
nor U12373 (N_12373,N_11051,N_11570);
nor U12374 (N_12374,N_11173,N_11438);
and U12375 (N_12375,N_11147,N_10824);
or U12376 (N_12376,N_11062,N_11861);
or U12377 (N_12377,N_11269,N_10596);
nand U12378 (N_12378,N_11014,N_11691);
xnor U12379 (N_12379,N_11455,N_11159);
or U12380 (N_12380,N_11897,N_10808);
nand U12381 (N_12381,N_10643,N_10946);
nand U12382 (N_12382,N_11260,N_10072);
and U12383 (N_12383,N_10591,N_11278);
xnor U12384 (N_12384,N_11328,N_10075);
or U12385 (N_12385,N_11514,N_11155);
nand U12386 (N_12386,N_11060,N_10455);
nor U12387 (N_12387,N_11970,N_11933);
xnor U12388 (N_12388,N_11111,N_10303);
or U12389 (N_12389,N_11959,N_10091);
or U12390 (N_12390,N_11716,N_11035);
and U12391 (N_12391,N_10966,N_10166);
xor U12392 (N_12392,N_11226,N_10840);
or U12393 (N_12393,N_10202,N_10657);
xnor U12394 (N_12394,N_10492,N_11877);
nor U12395 (N_12395,N_11404,N_10642);
nand U12396 (N_12396,N_10974,N_10718);
nor U12397 (N_12397,N_10959,N_10107);
xor U12398 (N_12398,N_10025,N_10369);
or U12399 (N_12399,N_11291,N_10370);
xnor U12400 (N_12400,N_10704,N_11216);
or U12401 (N_12401,N_10329,N_11059);
or U12402 (N_12402,N_11797,N_10586);
xor U12403 (N_12403,N_11578,N_11507);
or U12404 (N_12404,N_11782,N_10408);
nor U12405 (N_12405,N_10229,N_11680);
and U12406 (N_12406,N_10627,N_10292);
nand U12407 (N_12407,N_11465,N_10538);
or U12408 (N_12408,N_11124,N_10997);
and U12409 (N_12409,N_11865,N_10004);
nor U12410 (N_12410,N_11028,N_10011);
or U12411 (N_12411,N_10088,N_10473);
nand U12412 (N_12412,N_10217,N_10622);
nand U12413 (N_12413,N_11054,N_10190);
and U12414 (N_12414,N_11050,N_10533);
xnor U12415 (N_12415,N_10950,N_11794);
or U12416 (N_12416,N_11911,N_10035);
nand U12417 (N_12417,N_10681,N_11649);
xnor U12418 (N_12418,N_10637,N_11758);
xnor U12419 (N_12419,N_10344,N_10619);
xnor U12420 (N_12420,N_11237,N_11965);
xor U12421 (N_12421,N_10045,N_10975);
nand U12422 (N_12422,N_10655,N_10439);
xnor U12423 (N_12423,N_10793,N_11150);
or U12424 (N_12424,N_10382,N_10201);
and U12425 (N_12425,N_10071,N_11442);
nor U12426 (N_12426,N_11427,N_10315);
nand U12427 (N_12427,N_10034,N_10287);
or U12428 (N_12428,N_11479,N_11273);
or U12429 (N_12429,N_10413,N_10040);
or U12430 (N_12430,N_10234,N_11218);
and U12431 (N_12431,N_11345,N_11801);
xor U12432 (N_12432,N_10985,N_11366);
xor U12433 (N_12433,N_11096,N_11154);
and U12434 (N_12434,N_10428,N_10258);
nand U12435 (N_12435,N_10664,N_11566);
or U12436 (N_12436,N_10534,N_11550);
nand U12437 (N_12437,N_11535,N_11468);
xnor U12438 (N_12438,N_10914,N_11102);
xnor U12439 (N_12439,N_11394,N_11533);
or U12440 (N_12440,N_10522,N_11763);
xor U12441 (N_12441,N_10018,N_11950);
or U12442 (N_12442,N_10539,N_11197);
nor U12443 (N_12443,N_10264,N_11392);
or U12444 (N_12444,N_11573,N_10680);
or U12445 (N_12445,N_10041,N_10015);
or U12446 (N_12446,N_10307,N_10078);
nand U12447 (N_12447,N_11639,N_10749);
nand U12448 (N_12448,N_11887,N_11232);
and U12449 (N_12449,N_10335,N_10981);
xnor U12450 (N_12450,N_11851,N_10426);
nor U12451 (N_12451,N_11006,N_11099);
or U12452 (N_12452,N_11270,N_10769);
and U12453 (N_12453,N_10171,N_10766);
and U12454 (N_12454,N_10782,N_10020);
xor U12455 (N_12455,N_10409,N_10615);
nand U12456 (N_12456,N_11433,N_11623);
nand U12457 (N_12457,N_10430,N_10960);
and U12458 (N_12458,N_11002,N_11341);
nand U12459 (N_12459,N_11025,N_11324);
nor U12460 (N_12460,N_10036,N_10158);
nor U12461 (N_12461,N_11230,N_10529);
xnor U12462 (N_12462,N_11665,N_11714);
xor U12463 (N_12463,N_11505,N_11936);
xor U12464 (N_12464,N_10354,N_10037);
or U12465 (N_12465,N_10172,N_10592);
or U12466 (N_12466,N_11423,N_10841);
nor U12467 (N_12467,N_10253,N_10776);
nand U12468 (N_12468,N_10554,N_11770);
nor U12469 (N_12469,N_10096,N_10286);
and U12470 (N_12470,N_10570,N_10576);
nor U12471 (N_12471,N_11211,N_11694);
and U12472 (N_12472,N_10402,N_11026);
nor U12473 (N_12473,N_10553,N_10584);
or U12474 (N_12474,N_10843,N_10367);
xor U12475 (N_12475,N_11878,N_11747);
nand U12476 (N_12476,N_10693,N_11137);
nor U12477 (N_12477,N_11864,N_11160);
nand U12478 (N_12478,N_10415,N_10785);
or U12479 (N_12479,N_11011,N_10759);
nand U12480 (N_12480,N_10526,N_10181);
or U12481 (N_12481,N_10251,N_10524);
nor U12482 (N_12482,N_11329,N_10977);
and U12483 (N_12483,N_10144,N_10434);
xor U12484 (N_12484,N_10588,N_10112);
and U12485 (N_12485,N_10399,N_10669);
nor U12486 (N_12486,N_10725,N_10496);
or U12487 (N_12487,N_11215,N_11867);
xor U12488 (N_12488,N_10279,N_10396);
xnor U12489 (N_12489,N_11611,N_11689);
nand U12490 (N_12490,N_10684,N_11266);
or U12491 (N_12491,N_11478,N_10043);
and U12492 (N_12492,N_11536,N_10888);
nor U12493 (N_12493,N_10760,N_11092);
and U12494 (N_12494,N_11903,N_10753);
nor U12495 (N_12495,N_11506,N_10180);
xnor U12496 (N_12496,N_10556,N_10022);
and U12497 (N_12497,N_11065,N_11530);
nand U12498 (N_12498,N_11676,N_10915);
nor U12499 (N_12499,N_10557,N_10666);
and U12500 (N_12500,N_10762,N_10495);
or U12501 (N_12501,N_11916,N_11127);
nor U12502 (N_12502,N_11386,N_10019);
nor U12503 (N_12503,N_11720,N_10150);
and U12504 (N_12504,N_10995,N_11267);
xnor U12505 (N_12505,N_10310,N_10923);
xor U12506 (N_12506,N_10411,N_10325);
and U12507 (N_12507,N_11986,N_10597);
xor U12508 (N_12508,N_10689,N_10783);
or U12509 (N_12509,N_11601,N_11250);
nand U12510 (N_12510,N_11894,N_10988);
and U12511 (N_12511,N_10196,N_10833);
or U12512 (N_12512,N_11615,N_10791);
nand U12513 (N_12513,N_10079,N_11212);
nand U12514 (N_12514,N_11312,N_11132);
xor U12515 (N_12515,N_11415,N_10443);
nand U12516 (N_12516,N_10744,N_11503);
and U12517 (N_12517,N_11043,N_10897);
and U12518 (N_12518,N_11198,N_10062);
xor U12519 (N_12519,N_10397,N_11460);
or U12520 (N_12520,N_10288,N_11037);
xnor U12521 (N_12521,N_11502,N_11673);
and U12522 (N_12522,N_11921,N_11912);
and U12523 (N_12523,N_10051,N_11817);
nor U12524 (N_12524,N_10555,N_10679);
and U12525 (N_12525,N_11525,N_11413);
xor U12526 (N_12526,N_10873,N_11734);
xor U12527 (N_12527,N_10710,N_11134);
and U12528 (N_12528,N_11485,N_11027);
and U12529 (N_12529,N_11640,N_11175);
nor U12530 (N_12530,N_11071,N_10964);
xnor U12531 (N_12531,N_10765,N_11582);
and U12532 (N_12532,N_11695,N_11625);
nor U12533 (N_12533,N_10696,N_11787);
xor U12534 (N_12534,N_11293,N_10270);
or U12535 (N_12535,N_10500,N_10803);
nand U12536 (N_12536,N_10787,N_11728);
xor U12537 (N_12537,N_10014,N_11013);
nor U12538 (N_12538,N_11793,N_10012);
or U12539 (N_12539,N_10493,N_10616);
or U12540 (N_12540,N_10745,N_11712);
nor U12541 (N_12541,N_10857,N_10502);
or U12542 (N_12542,N_10463,N_10024);
or U12543 (N_12543,N_11745,N_11105);
or U12544 (N_12544,N_11729,N_11475);
xor U12545 (N_12545,N_10141,N_10535);
nand U12546 (N_12546,N_10516,N_10714);
nand U12547 (N_12547,N_10626,N_10829);
or U12548 (N_12548,N_10176,N_11558);
xnor U12549 (N_12549,N_10119,N_10514);
or U12550 (N_12550,N_11450,N_11672);
xnor U12551 (N_12551,N_10734,N_10227);
nand U12552 (N_12552,N_10133,N_10895);
xnor U12553 (N_12553,N_10830,N_11112);
xor U12554 (N_12554,N_11336,N_11846);
xnor U12555 (N_12555,N_10487,N_10471);
and U12556 (N_12556,N_11855,N_11637);
xnor U12557 (N_12557,N_11401,N_11234);
xnor U12558 (N_12558,N_11646,N_11466);
nand U12559 (N_12559,N_10375,N_10349);
or U12560 (N_12560,N_11671,N_11031);
or U12561 (N_12561,N_10948,N_11133);
nand U12562 (N_12562,N_10649,N_10903);
nor U12563 (N_12563,N_11656,N_10910);
xnor U12564 (N_12564,N_11945,N_11481);
and U12565 (N_12565,N_11863,N_11621);
and U12566 (N_12566,N_11995,N_10973);
or U12567 (N_12567,N_10853,N_10193);
or U12568 (N_12568,N_10242,N_11812);
xnor U12569 (N_12569,N_11057,N_11913);
and U12570 (N_12570,N_11769,N_11858);
and U12571 (N_12571,N_11304,N_11032);
and U12572 (N_12572,N_11934,N_11524);
xnor U12573 (N_12573,N_10856,N_11010);
nor U12574 (N_12574,N_11066,N_11542);
nand U12575 (N_12575,N_11078,N_11839);
or U12576 (N_12576,N_11598,N_11761);
or U12577 (N_12577,N_11882,N_11363);
nand U12578 (N_12578,N_10149,N_10675);
nor U12579 (N_12579,N_10692,N_10178);
nand U12580 (N_12580,N_10947,N_10599);
or U12581 (N_12581,N_11973,N_10378);
nand U12582 (N_12582,N_10786,N_11303);
xor U12583 (N_12583,N_10392,N_11783);
or U12584 (N_12584,N_10618,N_11655);
xnor U12585 (N_12585,N_10383,N_11288);
nor U12586 (N_12586,N_11116,N_11985);
and U12587 (N_12587,N_11906,N_10157);
and U12588 (N_12588,N_11832,N_10249);
nand U12589 (N_12589,N_11988,N_11780);
nand U12590 (N_12590,N_10278,N_11286);
nor U12591 (N_12591,N_11257,N_10822);
nand U12592 (N_12592,N_10422,N_10311);
or U12593 (N_12593,N_11930,N_10322);
or U12594 (N_12594,N_11192,N_11521);
or U12595 (N_12595,N_10865,N_11508);
nand U12596 (N_12596,N_10611,N_10357);
nor U12597 (N_12597,N_11073,N_11749);
nor U12598 (N_12598,N_10982,N_11757);
xnor U12599 (N_12599,N_10259,N_11277);
or U12600 (N_12600,N_11120,N_10688);
and U12601 (N_12601,N_11755,N_11472);
nand U12602 (N_12602,N_11971,N_11700);
xnor U12603 (N_12603,N_10581,N_11889);
xor U12604 (N_12604,N_10636,N_10142);
and U12605 (N_12605,N_11370,N_11922);
nand U12606 (N_12606,N_11046,N_10268);
nand U12607 (N_12607,N_11909,N_10804);
nor U12608 (N_12608,N_10050,N_10016);
or U12609 (N_12609,N_10685,N_11501);
nor U12610 (N_12610,N_11845,N_11289);
or U12611 (N_12611,N_11135,N_11748);
nor U12612 (N_12612,N_11968,N_10703);
and U12613 (N_12613,N_11282,N_10365);
nor U12614 (N_12614,N_10566,N_11564);
nor U12615 (N_12615,N_10187,N_11915);
or U12616 (N_12616,N_10454,N_10564);
and U12617 (N_12617,N_11670,N_10799);
nor U12618 (N_12618,N_10678,N_11068);
nand U12619 (N_12619,N_10645,N_10773);
nor U12620 (N_12620,N_11543,N_10571);
or U12621 (N_12621,N_11739,N_11084);
or U12622 (N_12622,N_10136,N_11608);
or U12623 (N_12623,N_10683,N_11964);
or U12624 (N_12624,N_10272,N_10779);
xnor U12625 (N_12625,N_11779,N_10768);
nand U12626 (N_12626,N_11735,N_11033);
nor U12627 (N_12627,N_10928,N_10656);
xnor U12628 (N_12628,N_11958,N_11653);
nor U12629 (N_12629,N_11553,N_11451);
nand U12630 (N_12630,N_11668,N_11183);
nand U12631 (N_12631,N_10676,N_10537);
xor U12632 (N_12632,N_10274,N_10177);
or U12633 (N_12633,N_11039,N_11141);
or U12634 (N_12634,N_10713,N_10658);
nand U12635 (N_12635,N_10401,N_10205);
and U12636 (N_12636,N_11471,N_11527);
or U12637 (N_12637,N_11405,N_11194);
nor U12638 (N_12638,N_11532,N_11823);
nor U12639 (N_12639,N_11603,N_11923);
nand U12640 (N_12640,N_10498,N_10891);
and U12641 (N_12641,N_11421,N_11034);
or U12642 (N_12642,N_10027,N_11358);
nand U12643 (N_12643,N_11581,N_10001);
or U12644 (N_12644,N_11721,N_11436);
xor U12645 (N_12645,N_11130,N_11079);
xor U12646 (N_12646,N_11179,N_10125);
nand U12647 (N_12647,N_10842,N_10892);
nand U12648 (N_12648,N_11022,N_10266);
nor U12649 (N_12649,N_10417,N_11590);
xnor U12650 (N_12650,N_11686,N_11414);
nand U12651 (N_12651,N_11791,N_10875);
nor U12652 (N_12652,N_10100,N_10572);
or U12653 (N_12653,N_10472,N_10504);
nor U12654 (N_12654,N_11115,N_10938);
and U12655 (N_12655,N_11337,N_10827);
and U12656 (N_12656,N_10299,N_11298);
nand U12657 (N_12657,N_11316,N_11997);
and U12658 (N_12658,N_10348,N_11828);
or U12659 (N_12659,N_11947,N_10927);
nor U12660 (N_12660,N_11771,N_11617);
nand U12661 (N_12661,N_11087,N_10727);
or U12662 (N_12662,N_11310,N_10976);
xor U12663 (N_12663,N_10735,N_10044);
and U12664 (N_12664,N_10574,N_10700);
and U12665 (N_12665,N_10932,N_10720);
nand U12666 (N_12666,N_11790,N_11872);
and U12667 (N_12667,N_11021,N_11919);
nand U12668 (N_12668,N_11085,N_10271);
xor U12669 (N_12669,N_11605,N_10860);
or U12670 (N_12670,N_11696,N_10309);
xnor U12671 (N_12671,N_11849,N_11398);
or U12672 (N_12672,N_11967,N_10214);
nand U12673 (N_12673,N_10613,N_10210);
xnor U12674 (N_12674,N_10816,N_10998);
and U12675 (N_12675,N_10235,N_10029);
xor U12676 (N_12676,N_11387,N_10363);
or U12677 (N_12677,N_11323,N_11868);
nand U12678 (N_12678,N_10419,N_11190);
and U12679 (N_12679,N_11182,N_11411);
nand U12680 (N_12680,N_11299,N_11604);
or U12681 (N_12681,N_10849,N_11391);
xnor U12682 (N_12682,N_10261,N_10512);
and U12683 (N_12683,N_10161,N_10057);
xor U12684 (N_12684,N_11379,N_11023);
nor U12685 (N_12685,N_10373,N_11953);
and U12686 (N_12686,N_11572,N_10552);
nor U12687 (N_12687,N_11634,N_10108);
xnor U12688 (N_12688,N_10984,N_10384);
and U12689 (N_12689,N_11759,N_11383);
nor U12690 (N_12690,N_10818,N_11403);
nand U12691 (N_12691,N_10621,N_10644);
nand U12692 (N_12692,N_11453,N_10243);
nor U12693 (N_12693,N_11650,N_11384);
and U12694 (N_12694,N_10929,N_11520);
nor U12695 (N_12695,N_11613,N_11157);
nand U12696 (N_12696,N_11822,N_10106);
and U12697 (N_12697,N_10361,N_11644);
or U12698 (N_12698,N_11180,N_11494);
or U12699 (N_12699,N_11870,N_11511);
xor U12700 (N_12700,N_11187,N_10525);
xor U12701 (N_12701,N_10536,N_10376);
nand U12702 (N_12702,N_11240,N_11984);
or U12703 (N_12703,N_10913,N_11315);
and U12704 (N_12704,N_10147,N_11231);
nand U12705 (N_12705,N_10511,N_10451);
xnor U12706 (N_12706,N_11408,N_11308);
xor U12707 (N_12707,N_11445,N_11831);
and U12708 (N_12708,N_10110,N_10994);
or U12709 (N_12709,N_11075,N_11486);
nor U12710 (N_12710,N_11883,N_10832);
or U12711 (N_12711,N_10453,N_11452);
xor U12712 (N_12712,N_10167,N_11365);
nand U12713 (N_12713,N_11873,N_11937);
nor U12714 (N_12714,N_11818,N_11641);
nand U12715 (N_12715,N_11344,N_11583);
nor U12716 (N_12716,N_10894,N_10962);
nor U12717 (N_12717,N_10668,N_11905);
or U12718 (N_12718,N_10248,N_11067);
nand U12719 (N_12719,N_10543,N_11191);
nand U12720 (N_12720,N_10169,N_11170);
or U12721 (N_12721,N_11461,N_11412);
nand U12722 (N_12722,N_10937,N_11549);
nand U12723 (N_12723,N_10456,N_11825);
nand U12724 (N_12724,N_10662,N_10788);
xnor U12725 (N_12725,N_11881,N_11717);
or U12726 (N_12726,N_10640,N_10082);
xor U12727 (N_12727,N_10661,N_11977);
nor U12728 (N_12728,N_10874,N_10414);
or U12729 (N_12729,N_10489,N_10930);
nor U12730 (N_12730,N_11008,N_10582);
and U12731 (N_12731,N_10815,N_11434);
and U12732 (N_12732,N_11309,N_10980);
and U12733 (N_12733,N_11221,N_11314);
or U12734 (N_12734,N_10561,N_11287);
xor U12735 (N_12735,N_10862,N_11557);
or U12736 (N_12736,N_11616,N_11618);
or U12737 (N_12737,N_11972,N_11932);
nor U12738 (N_12738,N_10890,N_10084);
and U12739 (N_12739,N_11804,N_11247);
and U12740 (N_12740,N_11044,N_10876);
nand U12741 (N_12741,N_11435,N_11119);
and U12742 (N_12742,N_11430,N_10304);
nor U12743 (N_12743,N_11632,N_10294);
nand U12744 (N_12744,N_10032,N_10429);
nor U12745 (N_12745,N_10109,N_10851);
or U12746 (N_12746,N_11599,N_10595);
nand U12747 (N_12747,N_11429,N_10267);
and U12748 (N_12748,N_11920,N_11983);
and U12749 (N_12749,N_10801,N_10548);
xor U12750 (N_12750,N_11857,N_10448);
and U12751 (N_12751,N_10232,N_11416);
xor U12752 (N_12752,N_11651,N_10878);
nor U12753 (N_12753,N_11703,N_11607);
xnor U12754 (N_12754,N_10283,N_11371);
nand U12755 (N_12755,N_10811,N_10126);
and U12756 (N_12756,N_11682,N_10093);
and U12757 (N_12757,N_11681,N_10967);
or U12758 (N_12758,N_10848,N_10953);
xnor U12759 (N_12759,N_10907,N_10317);
xor U12760 (N_12760,N_10042,N_11146);
nand U12761 (N_12761,N_10065,N_10936);
xor U12762 (N_12762,N_10667,N_11214);
nand U12763 (N_12763,N_10134,N_10761);
xnor U12764 (N_12764,N_10922,N_11577);
or U12765 (N_12765,N_11070,N_10200);
and U12766 (N_12766,N_11901,N_11751);
nand U12767 (N_12767,N_11960,N_10506);
nor U12768 (N_12768,N_10889,N_11766);
or U12769 (N_12769,N_10215,N_10722);
or U12770 (N_12770,N_10805,N_10784);
and U12771 (N_12771,N_10056,N_10887);
nand U12772 (N_12772,N_11838,N_10345);
xnor U12773 (N_12773,N_10183,N_10327);
nor U12774 (N_12774,N_10238,N_10908);
nor U12775 (N_12775,N_11730,N_10182);
xnor U12776 (N_12776,N_10575,N_11143);
or U12777 (N_12777,N_11706,N_10441);
nand U12778 (N_12778,N_11963,N_11263);
xor U12779 (N_12779,N_10593,N_10069);
nand U12780 (N_12780,N_11349,N_11117);
xnor U12781 (N_12781,N_11940,N_11208);
nor U12782 (N_12782,N_11129,N_11080);
or U12783 (N_12783,N_11055,N_10437);
and U12784 (N_12784,N_10074,N_11492);
xor U12785 (N_12785,N_11224,N_11592);
nor U12786 (N_12786,N_11103,N_10224);
and U12787 (N_12787,N_11029,N_11585);
nor U12788 (N_12788,N_11061,N_11597);
and U12789 (N_12789,N_11332,N_11546);
nor U12790 (N_12790,N_10945,N_11285);
xnor U12791 (N_12791,N_10148,N_11708);
nand U12792 (N_12792,N_10073,N_10466);
or U12793 (N_12793,N_10587,N_10931);
nand U12794 (N_12794,N_11879,N_11372);
xor U12795 (N_12795,N_11568,N_10442);
nand U12796 (N_12796,N_11874,N_10445);
xnor U12797 (N_12797,N_11789,N_10049);
or U12798 (N_12798,N_11125,N_10152);
or U12799 (N_12799,N_11687,N_11554);
xnor U12800 (N_12800,N_11454,N_10706);
and U12801 (N_12801,N_10983,N_11095);
nor U12802 (N_12802,N_11594,N_11654);
and U12803 (N_12803,N_11942,N_10719);
nand U12804 (N_12804,N_10400,N_11012);
xor U12805 (N_12805,N_11699,N_10476);
and U12806 (N_12806,N_11074,N_10577);
or U12807 (N_12807,N_11104,N_10702);
and U12808 (N_12808,N_10305,N_10111);
nand U12809 (N_12809,N_10729,N_10220);
or U12810 (N_12810,N_11661,N_11806);
nor U12811 (N_12811,N_11225,N_10754);
and U12812 (N_12812,N_11935,N_10859);
nor U12813 (N_12813,N_11158,N_10845);
or U12814 (N_12814,N_10877,N_10153);
nand U12815 (N_12815,N_11320,N_11238);
nand U12816 (N_12816,N_11020,N_11469);
and U12817 (N_12817,N_10777,N_11969);
or U12818 (N_12818,N_10585,N_10275);
nand U12819 (N_12819,N_10360,N_10389);
or U12820 (N_12820,N_10226,N_10854);
or U12821 (N_12821,N_11500,N_11040);
nor U12822 (N_12822,N_11606,N_11480);
nand U12823 (N_12823,N_10164,N_10672);
xnor U12824 (N_12824,N_10730,N_10391);
nand U12825 (N_12825,N_11551,N_10068);
or U12826 (N_12826,N_11301,N_11295);
or U12827 (N_12827,N_10898,N_11385);
nor U12828 (N_12828,N_10632,N_11248);
and U12829 (N_12829,N_11268,N_11938);
and U12830 (N_12830,N_10999,N_10652);
nand U12831 (N_12831,N_10117,N_10394);
nor U12832 (N_12832,N_11281,N_11819);
xor U12833 (N_12833,N_10435,N_10650);
and U12834 (N_12834,N_10590,N_11630);
and U12835 (N_12835,N_11659,N_11688);
nand U12836 (N_12836,N_11196,N_10257);
nand U12837 (N_12837,N_11658,N_10697);
or U12838 (N_12838,N_11860,N_11600);
nor U12839 (N_12839,N_11840,N_10549);
nor U12840 (N_12840,N_10817,N_11042);
nor U12841 (N_12841,N_11567,N_11954);
or U12842 (N_12842,N_10992,N_11048);
xor U12843 (N_12843,N_11106,N_10405);
nand U12844 (N_12844,N_11580,N_10189);
and U12845 (N_12845,N_10395,N_11189);
nor U12846 (N_12846,N_10356,N_11540);
nand U12847 (N_12847,N_10295,N_11373);
and U12848 (N_12848,N_11946,N_10002);
nor U12849 (N_12849,N_10252,N_10444);
nor U12850 (N_12850,N_10814,N_11996);
nand U12851 (N_12851,N_11276,N_10802);
or U12852 (N_12852,N_11209,N_10009);
xor U12853 (N_12853,N_11645,N_10551);
and U12854 (N_12854,N_10868,N_11775);
nand U12855 (N_12855,N_10510,N_11677);
or U12856 (N_12856,N_11829,N_10763);
or U12857 (N_12857,N_10013,N_10101);
xnor U12858 (N_12858,N_11093,N_10623);
xnor U12859 (N_12859,N_10458,N_10515);
nor U12860 (N_12860,N_10213,N_11499);
nand U12861 (N_12861,N_10955,N_11172);
and U12862 (N_12862,N_11844,N_10151);
nand U12863 (N_12863,N_10297,N_10563);
xor U12864 (N_12864,N_11473,N_10660);
nand U12865 (N_12865,N_11886,N_11830);
nand U12866 (N_12866,N_11166,N_11516);
nand U12867 (N_12867,N_11826,N_11367);
nand U12868 (N_12868,N_11753,N_10054);
and U12869 (N_12869,N_10244,N_10089);
xor U12870 (N_12870,N_11513,N_11741);
xor U12871 (N_12871,N_11762,N_10165);
nor U12872 (N_12872,N_11827,N_10379);
or U12873 (N_12873,N_10320,N_10987);
or U12874 (N_12874,N_10813,N_11627);
or U12875 (N_12875,N_11862,N_11275);
nand U12876 (N_12876,N_10380,N_11217);
nand U12877 (N_12877,N_11626,N_10961);
and U12878 (N_12878,N_11432,N_11294);
xnor U12879 (N_12879,N_11781,N_10831);
and U12880 (N_12880,N_11265,N_10421);
nor U12881 (N_12881,N_10505,N_10677);
nor U12882 (N_12882,N_11418,N_10957);
nor U12883 (N_12883,N_10728,N_10544);
xor U12884 (N_12884,N_11707,N_11122);
xnor U12885 (N_12885,N_10195,N_10223);
or U12886 (N_12886,N_10519,N_10433);
and U12887 (N_12887,N_10241,N_11949);
xor U12888 (N_12888,N_11978,N_11504);
nand U12889 (N_12889,N_10646,N_10362);
and U12890 (N_12890,N_10328,N_11732);
xor U12891 (N_12891,N_10532,N_11941);
nand U12892 (N_12892,N_11356,N_10207);
or U12893 (N_12893,N_10944,N_11777);
nand U12894 (N_12894,N_10867,N_11444);
nor U12895 (N_12895,N_10388,N_10772);
nor U12896 (N_12896,N_10863,N_10160);
nand U12897 (N_12897,N_11683,N_11145);
nor U12898 (N_12898,N_11476,N_10080);
nand U12899 (N_12899,N_10798,N_11490);
and U12900 (N_12900,N_11390,N_11619);
nand U12901 (N_12901,N_10467,N_10872);
nor U12902 (N_12902,N_10284,N_10855);
or U12903 (N_12903,N_11325,N_10630);
xnor U12904 (N_12904,N_11108,N_11088);
nand U12905 (N_12905,N_11869,N_10707);
or U12906 (N_12906,N_10604,N_11346);
xor U12907 (N_12907,N_10909,N_10826);
xor U12908 (N_12908,N_11201,N_11648);
xnor U12909 (N_12909,N_10633,N_10355);
nor U12910 (N_12910,N_11261,N_11850);
and U12911 (N_12911,N_10280,N_11428);
or U12912 (N_12912,N_11052,N_10191);
nand U12913 (N_12913,N_11202,N_10447);
and U12914 (N_12914,N_11853,N_10218);
or U12915 (N_12915,N_10921,N_11589);
or U12916 (N_12916,N_11097,N_11227);
nor U12917 (N_12917,N_11318,N_10192);
and U12918 (N_12918,N_10460,N_11161);
or U12919 (N_12919,N_11142,N_10635);
xnor U12920 (N_12920,N_10739,N_11951);
or U12921 (N_12921,N_10351,N_10771);
xor U12922 (N_12922,N_11856,N_10835);
or U12923 (N_12923,N_10170,N_11447);
or U12924 (N_12924,N_11005,N_10979);
nor U12925 (N_12925,N_10474,N_11139);
and U12926 (N_12926,N_11072,N_11200);
nand U12927 (N_12927,N_10479,N_10789);
and U12928 (N_12928,N_10436,N_11204);
and U12929 (N_12929,N_10377,N_10641);
or U12930 (N_12930,N_10262,N_10743);
nand U12931 (N_12931,N_10186,N_11210);
xor U12932 (N_12932,N_11807,N_11024);
and U12933 (N_12933,N_10086,N_11441);
nand U12934 (N_12934,N_11186,N_10222);
or U12935 (N_12935,N_11736,N_11254);
or U12936 (N_12936,N_11462,N_11939);
and U12937 (N_12937,N_11545,N_11809);
nand U12938 (N_12938,N_10300,N_11393);
nor U12939 (N_12939,N_10023,N_10617);
nand U12940 (N_12940,N_11576,N_11420);
or U12941 (N_12941,N_11280,N_11354);
nor U12942 (N_12942,N_10861,N_11638);
and U12943 (N_12943,N_11177,N_11259);
nand U12944 (N_12944,N_10386,N_10568);
nor U12945 (N_12945,N_11628,N_10674);
nand U12946 (N_12946,N_10508,N_10559);
and U12947 (N_12947,N_11262,N_10350);
nor U12948 (N_12948,N_11064,N_11223);
nor U12949 (N_12949,N_11359,N_11388);
xor U12950 (N_12950,N_10483,N_11785);
and U12951 (N_12951,N_11563,N_11538);
xnor U12952 (N_12952,N_10269,N_10390);
xor U12953 (N_12953,N_10052,N_11875);
nor U12954 (N_12954,N_11296,N_11464);
nor U12955 (N_12955,N_10085,N_11962);
nand U12956 (N_12956,N_11272,N_11152);
or U12957 (N_12957,N_10846,N_11355);
or U12958 (N_12958,N_10711,N_10881);
and U12959 (N_12959,N_10578,N_11719);
nor U12960 (N_12960,N_11126,N_10038);
and U12961 (N_12961,N_11253,N_11992);
nor U12962 (N_12962,N_10175,N_10482);
or U12963 (N_12963,N_11030,N_11148);
nand U12964 (N_12964,N_11899,N_11140);
and U12965 (N_12965,N_11925,N_10097);
xnor U12966 (N_12966,N_11752,N_11395);
nor U12967 (N_12967,N_11463,N_10920);
nor U12968 (N_12968,N_10589,N_10723);
nor U12969 (N_12969,N_11561,N_11595);
nor U12970 (N_12970,N_11737,N_10939);
nand U12971 (N_12971,N_10000,N_10256);
and U12972 (N_12972,N_11058,N_10752);
nor U12973 (N_12973,N_10601,N_11718);
and U12974 (N_12974,N_11228,N_11361);
or U12975 (N_12975,N_11744,N_11101);
nand U12976 (N_12976,N_10410,N_10701);
xor U12977 (N_12977,N_11814,N_11292);
and U12978 (N_12978,N_11931,N_10104);
nand U12979 (N_12979,N_10090,N_11089);
nand U12980 (N_12980,N_10497,N_10188);
nand U12981 (N_12981,N_10302,N_11360);
or U12982 (N_12982,N_10060,N_11100);
xor U12983 (N_12983,N_11943,N_11895);
and U12984 (N_12984,N_10733,N_10721);
and U12985 (N_12985,N_11866,N_10203);
xor U12986 (N_12986,N_11342,N_11537);
nor U12987 (N_12987,N_11731,N_11107);
nor U12988 (N_12988,N_11764,N_10194);
nor U12989 (N_12989,N_10501,N_11982);
xnor U12990 (N_12990,N_11778,N_11069);
nor U12991 (N_12991,N_11662,N_11952);
and U12992 (N_12992,N_10398,N_11667);
or U12993 (N_12993,N_11131,N_11493);
or U12994 (N_12994,N_10580,N_11917);
and U12995 (N_12995,N_10334,N_11989);
nand U12996 (N_12996,N_11547,N_11834);
or U12997 (N_12997,N_11399,N_11153);
and U12998 (N_12998,N_10757,N_11098);
xor U12999 (N_12999,N_10968,N_11437);
or U13000 (N_13000,N_10916,N_11369);
and U13001 (N_13001,N_11168,N_10964);
and U13002 (N_13002,N_11384,N_10530);
xnor U13003 (N_13003,N_10436,N_11827);
or U13004 (N_13004,N_10537,N_11616);
nor U13005 (N_13005,N_11649,N_11765);
xnor U13006 (N_13006,N_10206,N_10163);
and U13007 (N_13007,N_11343,N_10754);
nor U13008 (N_13008,N_10798,N_11097);
or U13009 (N_13009,N_11322,N_10055);
and U13010 (N_13010,N_10043,N_11037);
or U13011 (N_13011,N_11234,N_11634);
nand U13012 (N_13012,N_10727,N_11732);
and U13013 (N_13013,N_11598,N_11112);
and U13014 (N_13014,N_10196,N_10706);
or U13015 (N_13015,N_10824,N_10658);
or U13016 (N_13016,N_11056,N_11008);
nand U13017 (N_13017,N_10230,N_10154);
nor U13018 (N_13018,N_10602,N_11450);
and U13019 (N_13019,N_10646,N_10548);
nand U13020 (N_13020,N_10571,N_11018);
or U13021 (N_13021,N_11816,N_10237);
and U13022 (N_13022,N_11223,N_11680);
nand U13023 (N_13023,N_11600,N_11940);
nor U13024 (N_13024,N_11736,N_11401);
or U13025 (N_13025,N_10595,N_11415);
xor U13026 (N_13026,N_11576,N_10137);
nand U13027 (N_13027,N_11334,N_10285);
and U13028 (N_13028,N_10886,N_11764);
nor U13029 (N_13029,N_10274,N_11057);
nor U13030 (N_13030,N_11752,N_10611);
nand U13031 (N_13031,N_11736,N_10826);
xor U13032 (N_13032,N_11086,N_10535);
nand U13033 (N_13033,N_10682,N_11021);
and U13034 (N_13034,N_10648,N_10195);
nand U13035 (N_13035,N_10438,N_11985);
and U13036 (N_13036,N_10690,N_10000);
and U13037 (N_13037,N_10828,N_11789);
nor U13038 (N_13038,N_10140,N_10410);
nand U13039 (N_13039,N_10948,N_11299);
and U13040 (N_13040,N_11559,N_11279);
and U13041 (N_13041,N_10853,N_10418);
xor U13042 (N_13042,N_10856,N_11022);
nand U13043 (N_13043,N_11013,N_10252);
nand U13044 (N_13044,N_11677,N_11989);
xnor U13045 (N_13045,N_11714,N_10448);
nand U13046 (N_13046,N_11361,N_11723);
or U13047 (N_13047,N_11219,N_11170);
xor U13048 (N_13048,N_10132,N_10558);
xor U13049 (N_13049,N_10750,N_10219);
xor U13050 (N_13050,N_11489,N_11324);
or U13051 (N_13051,N_10226,N_10792);
nor U13052 (N_13052,N_10305,N_11108);
and U13053 (N_13053,N_10366,N_11600);
xor U13054 (N_13054,N_10558,N_10525);
and U13055 (N_13055,N_10446,N_11947);
or U13056 (N_13056,N_11024,N_11543);
xnor U13057 (N_13057,N_10098,N_10611);
nand U13058 (N_13058,N_11299,N_11201);
xnor U13059 (N_13059,N_10888,N_11908);
nand U13060 (N_13060,N_11750,N_10051);
and U13061 (N_13061,N_11880,N_11792);
xor U13062 (N_13062,N_11796,N_10003);
or U13063 (N_13063,N_11998,N_10145);
nor U13064 (N_13064,N_11281,N_10864);
and U13065 (N_13065,N_11659,N_11316);
xnor U13066 (N_13066,N_11076,N_10308);
or U13067 (N_13067,N_11775,N_10702);
nor U13068 (N_13068,N_11359,N_11834);
nand U13069 (N_13069,N_11722,N_10607);
nor U13070 (N_13070,N_11999,N_11980);
and U13071 (N_13071,N_11356,N_11304);
xor U13072 (N_13072,N_11048,N_11089);
nand U13073 (N_13073,N_10875,N_11859);
xor U13074 (N_13074,N_11172,N_10885);
nor U13075 (N_13075,N_11747,N_11871);
nor U13076 (N_13076,N_11664,N_11052);
and U13077 (N_13077,N_11741,N_11761);
nor U13078 (N_13078,N_11135,N_11025);
or U13079 (N_13079,N_10394,N_10483);
nor U13080 (N_13080,N_10356,N_10023);
and U13081 (N_13081,N_11945,N_11869);
or U13082 (N_13082,N_10527,N_11814);
xnor U13083 (N_13083,N_11836,N_10356);
xor U13084 (N_13084,N_10462,N_11127);
and U13085 (N_13085,N_11780,N_10639);
xnor U13086 (N_13086,N_11626,N_11115);
nand U13087 (N_13087,N_11003,N_10084);
xor U13088 (N_13088,N_11067,N_10649);
and U13089 (N_13089,N_10543,N_11574);
and U13090 (N_13090,N_11551,N_10052);
and U13091 (N_13091,N_10591,N_10871);
xnor U13092 (N_13092,N_11587,N_11935);
nand U13093 (N_13093,N_11946,N_11704);
xor U13094 (N_13094,N_11308,N_11104);
or U13095 (N_13095,N_11872,N_10867);
or U13096 (N_13096,N_10464,N_11615);
nand U13097 (N_13097,N_11706,N_10207);
or U13098 (N_13098,N_10035,N_11444);
xor U13099 (N_13099,N_10963,N_10892);
xor U13100 (N_13100,N_11251,N_10576);
or U13101 (N_13101,N_11323,N_11345);
or U13102 (N_13102,N_11151,N_10699);
or U13103 (N_13103,N_10292,N_11510);
or U13104 (N_13104,N_10789,N_10673);
or U13105 (N_13105,N_11419,N_11153);
nand U13106 (N_13106,N_11908,N_11636);
nand U13107 (N_13107,N_11408,N_10506);
xor U13108 (N_13108,N_10992,N_10279);
nand U13109 (N_13109,N_11241,N_11120);
and U13110 (N_13110,N_10312,N_10738);
xor U13111 (N_13111,N_10023,N_10050);
nor U13112 (N_13112,N_10705,N_11898);
or U13113 (N_13113,N_10130,N_11649);
and U13114 (N_13114,N_10663,N_11173);
nor U13115 (N_13115,N_10153,N_11407);
xnor U13116 (N_13116,N_11093,N_10517);
xnor U13117 (N_13117,N_10106,N_10464);
nor U13118 (N_13118,N_10775,N_10359);
nor U13119 (N_13119,N_11219,N_10924);
xor U13120 (N_13120,N_11578,N_11458);
nand U13121 (N_13121,N_10890,N_11045);
xor U13122 (N_13122,N_11261,N_10293);
and U13123 (N_13123,N_10260,N_10030);
or U13124 (N_13124,N_11631,N_11853);
nand U13125 (N_13125,N_11467,N_10034);
or U13126 (N_13126,N_10748,N_10815);
xor U13127 (N_13127,N_10695,N_10678);
xnor U13128 (N_13128,N_10224,N_11689);
nor U13129 (N_13129,N_10948,N_11973);
or U13130 (N_13130,N_11522,N_10397);
and U13131 (N_13131,N_10982,N_11350);
nand U13132 (N_13132,N_11948,N_10093);
and U13133 (N_13133,N_11550,N_11549);
xnor U13134 (N_13134,N_10036,N_10785);
xnor U13135 (N_13135,N_10223,N_10426);
xor U13136 (N_13136,N_10062,N_10160);
xnor U13137 (N_13137,N_11882,N_10119);
and U13138 (N_13138,N_10222,N_10128);
nand U13139 (N_13139,N_11293,N_10772);
xor U13140 (N_13140,N_11280,N_10010);
nand U13141 (N_13141,N_10167,N_11551);
nor U13142 (N_13142,N_10043,N_10210);
or U13143 (N_13143,N_11896,N_10125);
nor U13144 (N_13144,N_10301,N_11763);
nor U13145 (N_13145,N_11757,N_10935);
nor U13146 (N_13146,N_11289,N_10075);
and U13147 (N_13147,N_10605,N_11988);
nand U13148 (N_13148,N_10604,N_11718);
and U13149 (N_13149,N_10251,N_10837);
xnor U13150 (N_13150,N_10933,N_11916);
nand U13151 (N_13151,N_10755,N_11955);
or U13152 (N_13152,N_10764,N_11010);
and U13153 (N_13153,N_11482,N_10752);
xnor U13154 (N_13154,N_10839,N_11525);
nor U13155 (N_13155,N_10773,N_11735);
xor U13156 (N_13156,N_10051,N_10097);
xnor U13157 (N_13157,N_11979,N_10824);
nand U13158 (N_13158,N_10930,N_10749);
nand U13159 (N_13159,N_11002,N_11753);
nor U13160 (N_13160,N_10361,N_10723);
or U13161 (N_13161,N_10861,N_11035);
nor U13162 (N_13162,N_10870,N_10831);
nor U13163 (N_13163,N_11368,N_11099);
nor U13164 (N_13164,N_10289,N_11650);
nand U13165 (N_13165,N_11563,N_10655);
and U13166 (N_13166,N_11756,N_11062);
nand U13167 (N_13167,N_11588,N_11056);
xnor U13168 (N_13168,N_10435,N_10602);
nand U13169 (N_13169,N_11744,N_11652);
and U13170 (N_13170,N_10790,N_10663);
nor U13171 (N_13171,N_11571,N_11540);
xor U13172 (N_13172,N_10624,N_11376);
nand U13173 (N_13173,N_11104,N_11903);
nand U13174 (N_13174,N_10784,N_11527);
xnor U13175 (N_13175,N_10206,N_11722);
nor U13176 (N_13176,N_10766,N_10443);
nand U13177 (N_13177,N_11123,N_11921);
and U13178 (N_13178,N_10160,N_10903);
xor U13179 (N_13179,N_11072,N_10305);
nand U13180 (N_13180,N_10286,N_11200);
or U13181 (N_13181,N_11609,N_10156);
or U13182 (N_13182,N_10350,N_10212);
xnor U13183 (N_13183,N_11838,N_10962);
nand U13184 (N_13184,N_11786,N_10509);
nor U13185 (N_13185,N_11330,N_10871);
or U13186 (N_13186,N_11606,N_11674);
nor U13187 (N_13187,N_10740,N_11055);
xnor U13188 (N_13188,N_11217,N_11709);
nor U13189 (N_13189,N_11155,N_11114);
xnor U13190 (N_13190,N_10920,N_11284);
xor U13191 (N_13191,N_10138,N_11417);
xor U13192 (N_13192,N_10370,N_10884);
nor U13193 (N_13193,N_11589,N_10644);
nor U13194 (N_13194,N_10733,N_10169);
and U13195 (N_13195,N_10526,N_11842);
or U13196 (N_13196,N_10713,N_11320);
xnor U13197 (N_13197,N_11028,N_11667);
or U13198 (N_13198,N_10928,N_11145);
xor U13199 (N_13199,N_10556,N_10724);
xor U13200 (N_13200,N_10898,N_10129);
and U13201 (N_13201,N_11871,N_11814);
and U13202 (N_13202,N_11703,N_10225);
nand U13203 (N_13203,N_10159,N_11729);
nand U13204 (N_13204,N_10077,N_11626);
xnor U13205 (N_13205,N_10762,N_11944);
nor U13206 (N_13206,N_11865,N_10732);
nor U13207 (N_13207,N_11857,N_11406);
nor U13208 (N_13208,N_11048,N_10174);
nand U13209 (N_13209,N_11763,N_11083);
and U13210 (N_13210,N_11838,N_11070);
or U13211 (N_13211,N_10661,N_10902);
nor U13212 (N_13212,N_11346,N_11661);
or U13213 (N_13213,N_11426,N_10894);
and U13214 (N_13214,N_10387,N_11239);
nand U13215 (N_13215,N_10715,N_11800);
and U13216 (N_13216,N_10018,N_10518);
xnor U13217 (N_13217,N_10739,N_10403);
nand U13218 (N_13218,N_11105,N_11465);
xor U13219 (N_13219,N_10915,N_10031);
or U13220 (N_13220,N_10792,N_10151);
nand U13221 (N_13221,N_10423,N_10029);
or U13222 (N_13222,N_10826,N_10749);
nand U13223 (N_13223,N_11823,N_11459);
nor U13224 (N_13224,N_11720,N_11670);
xor U13225 (N_13225,N_11040,N_10871);
and U13226 (N_13226,N_11001,N_10920);
or U13227 (N_13227,N_11091,N_10919);
nor U13228 (N_13228,N_11192,N_11718);
xnor U13229 (N_13229,N_11156,N_10932);
and U13230 (N_13230,N_11613,N_10935);
nor U13231 (N_13231,N_11285,N_10710);
or U13232 (N_13232,N_10548,N_10048);
and U13233 (N_13233,N_10232,N_11513);
and U13234 (N_13234,N_10164,N_11931);
or U13235 (N_13235,N_10677,N_10496);
xnor U13236 (N_13236,N_10911,N_11240);
or U13237 (N_13237,N_10148,N_11609);
or U13238 (N_13238,N_11502,N_10692);
and U13239 (N_13239,N_11852,N_11145);
nor U13240 (N_13240,N_11078,N_10044);
nand U13241 (N_13241,N_11903,N_11835);
nor U13242 (N_13242,N_10348,N_11294);
or U13243 (N_13243,N_11127,N_11841);
nand U13244 (N_13244,N_11341,N_11172);
xnor U13245 (N_13245,N_10579,N_10428);
nand U13246 (N_13246,N_11778,N_10522);
xnor U13247 (N_13247,N_10688,N_11119);
nor U13248 (N_13248,N_10218,N_11257);
nand U13249 (N_13249,N_10586,N_11775);
nor U13250 (N_13250,N_11840,N_11367);
nor U13251 (N_13251,N_10117,N_11157);
or U13252 (N_13252,N_11104,N_10540);
xor U13253 (N_13253,N_11599,N_11520);
nand U13254 (N_13254,N_10512,N_11998);
and U13255 (N_13255,N_10847,N_10057);
and U13256 (N_13256,N_11846,N_10198);
nand U13257 (N_13257,N_10824,N_10237);
or U13258 (N_13258,N_10047,N_11809);
or U13259 (N_13259,N_11531,N_11039);
and U13260 (N_13260,N_11885,N_11004);
nand U13261 (N_13261,N_10776,N_11426);
nor U13262 (N_13262,N_11327,N_11118);
nor U13263 (N_13263,N_11007,N_11755);
or U13264 (N_13264,N_11487,N_10282);
xor U13265 (N_13265,N_11392,N_10065);
nor U13266 (N_13266,N_10906,N_11317);
xnor U13267 (N_13267,N_10510,N_10747);
and U13268 (N_13268,N_11137,N_11554);
and U13269 (N_13269,N_11083,N_10559);
or U13270 (N_13270,N_10694,N_11978);
nor U13271 (N_13271,N_11704,N_11223);
or U13272 (N_13272,N_10240,N_11357);
nand U13273 (N_13273,N_11134,N_11756);
nor U13274 (N_13274,N_11904,N_10138);
or U13275 (N_13275,N_10679,N_10506);
and U13276 (N_13276,N_11965,N_11931);
xor U13277 (N_13277,N_11659,N_10565);
nor U13278 (N_13278,N_10633,N_10021);
or U13279 (N_13279,N_10628,N_10329);
xor U13280 (N_13280,N_11692,N_11417);
and U13281 (N_13281,N_11406,N_10129);
nor U13282 (N_13282,N_10233,N_10318);
and U13283 (N_13283,N_11665,N_10197);
xor U13284 (N_13284,N_11144,N_11172);
nor U13285 (N_13285,N_10569,N_11976);
and U13286 (N_13286,N_11121,N_10872);
and U13287 (N_13287,N_11477,N_10729);
and U13288 (N_13288,N_11627,N_10099);
nor U13289 (N_13289,N_10354,N_11767);
nor U13290 (N_13290,N_11225,N_10463);
or U13291 (N_13291,N_10448,N_11523);
and U13292 (N_13292,N_10888,N_10132);
or U13293 (N_13293,N_10540,N_10071);
nor U13294 (N_13294,N_10439,N_11767);
nand U13295 (N_13295,N_11068,N_10536);
or U13296 (N_13296,N_11826,N_11119);
or U13297 (N_13297,N_10690,N_11180);
nor U13298 (N_13298,N_10480,N_11297);
xor U13299 (N_13299,N_10020,N_10132);
nor U13300 (N_13300,N_10283,N_10326);
and U13301 (N_13301,N_10065,N_11059);
or U13302 (N_13302,N_11580,N_11240);
nand U13303 (N_13303,N_11157,N_11211);
nor U13304 (N_13304,N_10241,N_10974);
or U13305 (N_13305,N_11296,N_11613);
and U13306 (N_13306,N_10661,N_10817);
nand U13307 (N_13307,N_10827,N_10651);
nor U13308 (N_13308,N_10657,N_10956);
nor U13309 (N_13309,N_11815,N_11036);
and U13310 (N_13310,N_11011,N_10636);
xor U13311 (N_13311,N_11959,N_11862);
nand U13312 (N_13312,N_11431,N_10095);
or U13313 (N_13313,N_10654,N_10370);
nand U13314 (N_13314,N_11588,N_10085);
xor U13315 (N_13315,N_10573,N_11471);
or U13316 (N_13316,N_10998,N_11634);
nor U13317 (N_13317,N_11588,N_11760);
nor U13318 (N_13318,N_10240,N_11577);
nor U13319 (N_13319,N_10674,N_10304);
nand U13320 (N_13320,N_11249,N_10938);
nor U13321 (N_13321,N_10469,N_10331);
nor U13322 (N_13322,N_10907,N_10084);
nor U13323 (N_13323,N_10438,N_10697);
xnor U13324 (N_13324,N_11514,N_11144);
xnor U13325 (N_13325,N_10026,N_11338);
or U13326 (N_13326,N_11325,N_10309);
and U13327 (N_13327,N_11558,N_10610);
xor U13328 (N_13328,N_10866,N_11314);
and U13329 (N_13329,N_10606,N_11475);
nor U13330 (N_13330,N_10397,N_11379);
and U13331 (N_13331,N_11481,N_11467);
nor U13332 (N_13332,N_11792,N_11744);
and U13333 (N_13333,N_11344,N_11039);
and U13334 (N_13334,N_11104,N_10265);
and U13335 (N_13335,N_11365,N_11876);
and U13336 (N_13336,N_10608,N_11446);
or U13337 (N_13337,N_11426,N_10739);
and U13338 (N_13338,N_11088,N_11145);
nor U13339 (N_13339,N_10509,N_11237);
and U13340 (N_13340,N_11925,N_11494);
xor U13341 (N_13341,N_11567,N_10945);
or U13342 (N_13342,N_10341,N_11519);
or U13343 (N_13343,N_11905,N_11384);
nor U13344 (N_13344,N_11636,N_10538);
or U13345 (N_13345,N_10776,N_10082);
and U13346 (N_13346,N_10332,N_11395);
nor U13347 (N_13347,N_11384,N_11061);
or U13348 (N_13348,N_10603,N_10681);
xnor U13349 (N_13349,N_11510,N_10890);
and U13350 (N_13350,N_11481,N_10591);
nor U13351 (N_13351,N_11547,N_11412);
nor U13352 (N_13352,N_10371,N_11929);
nand U13353 (N_13353,N_10272,N_10499);
nor U13354 (N_13354,N_11181,N_10540);
or U13355 (N_13355,N_11146,N_11500);
nand U13356 (N_13356,N_10230,N_11957);
xnor U13357 (N_13357,N_11857,N_10757);
nand U13358 (N_13358,N_11568,N_11810);
nor U13359 (N_13359,N_11864,N_11046);
nand U13360 (N_13360,N_10938,N_10997);
nand U13361 (N_13361,N_11785,N_10770);
or U13362 (N_13362,N_10794,N_10372);
xor U13363 (N_13363,N_11504,N_10780);
xnor U13364 (N_13364,N_11614,N_10605);
or U13365 (N_13365,N_11936,N_10053);
nor U13366 (N_13366,N_10770,N_10207);
nand U13367 (N_13367,N_10603,N_10552);
nand U13368 (N_13368,N_11844,N_10162);
nor U13369 (N_13369,N_11276,N_11651);
nor U13370 (N_13370,N_11343,N_11544);
or U13371 (N_13371,N_11811,N_10526);
xor U13372 (N_13372,N_11133,N_10159);
xnor U13373 (N_13373,N_11040,N_11804);
nor U13374 (N_13374,N_11665,N_10157);
and U13375 (N_13375,N_11193,N_10480);
and U13376 (N_13376,N_11399,N_11927);
or U13377 (N_13377,N_11798,N_10057);
or U13378 (N_13378,N_10826,N_10415);
nand U13379 (N_13379,N_10121,N_11032);
nor U13380 (N_13380,N_10212,N_11174);
and U13381 (N_13381,N_10459,N_11048);
xor U13382 (N_13382,N_11972,N_11978);
nand U13383 (N_13383,N_10838,N_10362);
or U13384 (N_13384,N_11817,N_11856);
nand U13385 (N_13385,N_10375,N_11450);
xor U13386 (N_13386,N_10036,N_11131);
xnor U13387 (N_13387,N_11103,N_10800);
nand U13388 (N_13388,N_10936,N_11202);
xnor U13389 (N_13389,N_10719,N_10206);
xor U13390 (N_13390,N_11006,N_10307);
xor U13391 (N_13391,N_11836,N_10067);
nor U13392 (N_13392,N_10504,N_10278);
nand U13393 (N_13393,N_10874,N_11209);
nand U13394 (N_13394,N_11043,N_11198);
or U13395 (N_13395,N_10795,N_11294);
or U13396 (N_13396,N_10677,N_10201);
nand U13397 (N_13397,N_11013,N_11995);
nand U13398 (N_13398,N_11911,N_11930);
nor U13399 (N_13399,N_10970,N_10644);
nand U13400 (N_13400,N_11069,N_10997);
xor U13401 (N_13401,N_11845,N_10987);
or U13402 (N_13402,N_11825,N_11761);
xor U13403 (N_13403,N_11599,N_10108);
xnor U13404 (N_13404,N_10494,N_11592);
or U13405 (N_13405,N_11794,N_10182);
nor U13406 (N_13406,N_11486,N_10443);
xnor U13407 (N_13407,N_11972,N_11810);
nand U13408 (N_13408,N_10802,N_10743);
or U13409 (N_13409,N_10313,N_10702);
xnor U13410 (N_13410,N_11475,N_11682);
and U13411 (N_13411,N_10344,N_10155);
nand U13412 (N_13412,N_10642,N_10563);
xnor U13413 (N_13413,N_10617,N_10649);
nand U13414 (N_13414,N_10382,N_10000);
or U13415 (N_13415,N_10475,N_10196);
and U13416 (N_13416,N_11729,N_10080);
nor U13417 (N_13417,N_11515,N_11017);
and U13418 (N_13418,N_10534,N_11110);
nor U13419 (N_13419,N_11424,N_11556);
nor U13420 (N_13420,N_11895,N_10810);
and U13421 (N_13421,N_11480,N_10121);
nand U13422 (N_13422,N_11758,N_11208);
or U13423 (N_13423,N_11384,N_10283);
nand U13424 (N_13424,N_10675,N_11053);
or U13425 (N_13425,N_11765,N_10604);
and U13426 (N_13426,N_10584,N_10094);
xnor U13427 (N_13427,N_10660,N_10790);
and U13428 (N_13428,N_10980,N_10258);
and U13429 (N_13429,N_10619,N_11148);
nand U13430 (N_13430,N_10959,N_10640);
and U13431 (N_13431,N_11229,N_10307);
nand U13432 (N_13432,N_10828,N_10710);
xor U13433 (N_13433,N_10206,N_11145);
nor U13434 (N_13434,N_11086,N_11430);
xnor U13435 (N_13435,N_10336,N_11924);
nand U13436 (N_13436,N_10609,N_11579);
nor U13437 (N_13437,N_11365,N_11154);
xor U13438 (N_13438,N_11811,N_11362);
xnor U13439 (N_13439,N_10028,N_11216);
xnor U13440 (N_13440,N_11115,N_10785);
xor U13441 (N_13441,N_10683,N_11965);
or U13442 (N_13442,N_11690,N_10838);
nand U13443 (N_13443,N_10527,N_11483);
nand U13444 (N_13444,N_11385,N_11267);
xnor U13445 (N_13445,N_10465,N_11580);
or U13446 (N_13446,N_11859,N_11714);
xnor U13447 (N_13447,N_10649,N_10830);
nor U13448 (N_13448,N_11291,N_11559);
and U13449 (N_13449,N_10726,N_11641);
and U13450 (N_13450,N_10212,N_11885);
xnor U13451 (N_13451,N_11418,N_10526);
xnor U13452 (N_13452,N_10563,N_11856);
xor U13453 (N_13453,N_10110,N_11762);
nand U13454 (N_13454,N_11700,N_10375);
and U13455 (N_13455,N_10766,N_11574);
and U13456 (N_13456,N_10713,N_11832);
and U13457 (N_13457,N_10638,N_11415);
xor U13458 (N_13458,N_11712,N_10996);
xnor U13459 (N_13459,N_10172,N_11700);
or U13460 (N_13460,N_10794,N_10039);
nand U13461 (N_13461,N_10889,N_11682);
xnor U13462 (N_13462,N_11270,N_11462);
or U13463 (N_13463,N_10232,N_10719);
xnor U13464 (N_13464,N_11966,N_11787);
nor U13465 (N_13465,N_10936,N_11137);
nand U13466 (N_13466,N_11263,N_10222);
nor U13467 (N_13467,N_10108,N_10540);
or U13468 (N_13468,N_11071,N_11347);
nor U13469 (N_13469,N_11560,N_10529);
nor U13470 (N_13470,N_11408,N_10427);
nand U13471 (N_13471,N_11167,N_10344);
xor U13472 (N_13472,N_11160,N_11208);
nand U13473 (N_13473,N_11163,N_11626);
nand U13474 (N_13474,N_11754,N_11738);
xor U13475 (N_13475,N_10885,N_10672);
and U13476 (N_13476,N_10157,N_10476);
nand U13477 (N_13477,N_10958,N_11138);
nand U13478 (N_13478,N_10965,N_10172);
nand U13479 (N_13479,N_11816,N_11751);
and U13480 (N_13480,N_10412,N_10299);
and U13481 (N_13481,N_11946,N_10455);
or U13482 (N_13482,N_10259,N_10215);
and U13483 (N_13483,N_11197,N_11493);
or U13484 (N_13484,N_11040,N_11233);
and U13485 (N_13485,N_10186,N_11647);
nor U13486 (N_13486,N_11103,N_10791);
and U13487 (N_13487,N_10038,N_11689);
nand U13488 (N_13488,N_10423,N_11397);
or U13489 (N_13489,N_10292,N_10398);
nor U13490 (N_13490,N_10573,N_10209);
nor U13491 (N_13491,N_10931,N_11944);
nor U13492 (N_13492,N_10954,N_10111);
and U13493 (N_13493,N_11004,N_10774);
and U13494 (N_13494,N_11413,N_10199);
nor U13495 (N_13495,N_11626,N_10540);
or U13496 (N_13496,N_11202,N_10405);
xor U13497 (N_13497,N_10751,N_11235);
xor U13498 (N_13498,N_11210,N_10806);
or U13499 (N_13499,N_11154,N_11648);
nor U13500 (N_13500,N_11057,N_10101);
and U13501 (N_13501,N_11602,N_10088);
and U13502 (N_13502,N_10589,N_11893);
and U13503 (N_13503,N_10164,N_11608);
and U13504 (N_13504,N_10432,N_11272);
nand U13505 (N_13505,N_10350,N_10199);
or U13506 (N_13506,N_10203,N_10540);
nand U13507 (N_13507,N_10759,N_11030);
xor U13508 (N_13508,N_10978,N_11866);
and U13509 (N_13509,N_11156,N_10903);
and U13510 (N_13510,N_11776,N_10746);
and U13511 (N_13511,N_10108,N_10200);
or U13512 (N_13512,N_11861,N_11196);
or U13513 (N_13513,N_11952,N_10900);
nand U13514 (N_13514,N_11682,N_10217);
and U13515 (N_13515,N_10666,N_10636);
or U13516 (N_13516,N_10319,N_10545);
and U13517 (N_13517,N_11882,N_11974);
nand U13518 (N_13518,N_10049,N_10895);
xnor U13519 (N_13519,N_11313,N_10024);
or U13520 (N_13520,N_11966,N_11631);
and U13521 (N_13521,N_10279,N_11696);
and U13522 (N_13522,N_11947,N_11593);
and U13523 (N_13523,N_11912,N_11859);
and U13524 (N_13524,N_10241,N_11252);
or U13525 (N_13525,N_11208,N_11223);
and U13526 (N_13526,N_10314,N_11838);
or U13527 (N_13527,N_11736,N_11576);
and U13528 (N_13528,N_11605,N_10100);
nor U13529 (N_13529,N_11490,N_11283);
or U13530 (N_13530,N_10247,N_10257);
and U13531 (N_13531,N_11525,N_10785);
and U13532 (N_13532,N_10605,N_10442);
xnor U13533 (N_13533,N_11191,N_11981);
xnor U13534 (N_13534,N_10055,N_10667);
xnor U13535 (N_13535,N_11579,N_10311);
xor U13536 (N_13536,N_10384,N_11154);
or U13537 (N_13537,N_10855,N_10856);
and U13538 (N_13538,N_11687,N_10157);
nand U13539 (N_13539,N_10695,N_11040);
nand U13540 (N_13540,N_10377,N_11791);
and U13541 (N_13541,N_10373,N_10277);
nand U13542 (N_13542,N_10000,N_10338);
nand U13543 (N_13543,N_11152,N_11582);
nand U13544 (N_13544,N_10686,N_11095);
nand U13545 (N_13545,N_10512,N_10488);
nand U13546 (N_13546,N_10560,N_11705);
nor U13547 (N_13547,N_11141,N_10734);
nor U13548 (N_13548,N_11284,N_11323);
nand U13549 (N_13549,N_11908,N_10674);
nand U13550 (N_13550,N_10965,N_11043);
or U13551 (N_13551,N_10104,N_10554);
nand U13552 (N_13552,N_11352,N_11852);
or U13553 (N_13553,N_10526,N_11574);
xor U13554 (N_13554,N_11447,N_10700);
nor U13555 (N_13555,N_11355,N_10910);
nand U13556 (N_13556,N_11819,N_10038);
and U13557 (N_13557,N_11869,N_11596);
xnor U13558 (N_13558,N_11374,N_10681);
nor U13559 (N_13559,N_10127,N_10919);
or U13560 (N_13560,N_11365,N_10474);
nor U13561 (N_13561,N_11022,N_10729);
or U13562 (N_13562,N_11548,N_11821);
and U13563 (N_13563,N_11199,N_10300);
or U13564 (N_13564,N_11606,N_11281);
xnor U13565 (N_13565,N_11280,N_11210);
xnor U13566 (N_13566,N_10264,N_10114);
nor U13567 (N_13567,N_10920,N_11131);
xor U13568 (N_13568,N_11186,N_10245);
and U13569 (N_13569,N_11762,N_10134);
or U13570 (N_13570,N_11317,N_11573);
or U13571 (N_13571,N_11313,N_10905);
or U13572 (N_13572,N_11502,N_10554);
or U13573 (N_13573,N_10088,N_11106);
nand U13574 (N_13574,N_11450,N_11618);
nand U13575 (N_13575,N_11186,N_11651);
and U13576 (N_13576,N_10178,N_11496);
nor U13577 (N_13577,N_11846,N_11174);
or U13578 (N_13578,N_11912,N_10665);
and U13579 (N_13579,N_11034,N_10097);
nor U13580 (N_13580,N_11412,N_11459);
nor U13581 (N_13581,N_11952,N_10178);
or U13582 (N_13582,N_10870,N_11976);
nor U13583 (N_13583,N_11477,N_11068);
and U13584 (N_13584,N_10635,N_10733);
nor U13585 (N_13585,N_11780,N_10581);
and U13586 (N_13586,N_10830,N_10158);
and U13587 (N_13587,N_11250,N_10505);
nor U13588 (N_13588,N_10763,N_11228);
or U13589 (N_13589,N_11789,N_10999);
nand U13590 (N_13590,N_11940,N_10507);
nand U13591 (N_13591,N_10729,N_11335);
nor U13592 (N_13592,N_10697,N_11027);
or U13593 (N_13593,N_11298,N_11168);
or U13594 (N_13594,N_11984,N_11503);
nand U13595 (N_13595,N_11545,N_10284);
nand U13596 (N_13596,N_10227,N_10726);
nand U13597 (N_13597,N_10596,N_11181);
and U13598 (N_13598,N_11088,N_11168);
nor U13599 (N_13599,N_11786,N_11112);
nand U13600 (N_13600,N_10665,N_10395);
nor U13601 (N_13601,N_10003,N_10160);
nand U13602 (N_13602,N_10843,N_10934);
and U13603 (N_13603,N_10716,N_10956);
nand U13604 (N_13604,N_11893,N_10610);
xnor U13605 (N_13605,N_11050,N_11309);
or U13606 (N_13606,N_10200,N_10189);
nand U13607 (N_13607,N_10769,N_11768);
or U13608 (N_13608,N_11680,N_11139);
nand U13609 (N_13609,N_11203,N_11550);
or U13610 (N_13610,N_11476,N_11199);
or U13611 (N_13611,N_10291,N_11400);
and U13612 (N_13612,N_11055,N_10168);
nand U13613 (N_13613,N_10495,N_11159);
nor U13614 (N_13614,N_11303,N_10260);
nand U13615 (N_13615,N_10267,N_10334);
nand U13616 (N_13616,N_10471,N_10140);
nor U13617 (N_13617,N_11809,N_11604);
xnor U13618 (N_13618,N_10321,N_10014);
or U13619 (N_13619,N_10390,N_10588);
or U13620 (N_13620,N_10539,N_11151);
nor U13621 (N_13621,N_10769,N_10633);
nand U13622 (N_13622,N_10662,N_11322);
nor U13623 (N_13623,N_10872,N_10067);
and U13624 (N_13624,N_11702,N_11595);
xnor U13625 (N_13625,N_10555,N_10749);
xor U13626 (N_13626,N_10154,N_10994);
xor U13627 (N_13627,N_11736,N_10752);
xor U13628 (N_13628,N_10776,N_11799);
xnor U13629 (N_13629,N_11199,N_11642);
xnor U13630 (N_13630,N_11839,N_10327);
nand U13631 (N_13631,N_10558,N_11743);
nor U13632 (N_13632,N_10524,N_11414);
xor U13633 (N_13633,N_11539,N_10454);
xor U13634 (N_13634,N_10623,N_10982);
xnor U13635 (N_13635,N_11842,N_11059);
nand U13636 (N_13636,N_11180,N_10560);
and U13637 (N_13637,N_10984,N_11249);
nand U13638 (N_13638,N_11033,N_11191);
or U13639 (N_13639,N_10595,N_11962);
and U13640 (N_13640,N_10309,N_10380);
nor U13641 (N_13641,N_11361,N_10466);
nand U13642 (N_13642,N_11780,N_10687);
nor U13643 (N_13643,N_10576,N_10297);
and U13644 (N_13644,N_10260,N_11995);
or U13645 (N_13645,N_11324,N_11340);
and U13646 (N_13646,N_10303,N_10217);
nor U13647 (N_13647,N_10951,N_10127);
and U13648 (N_13648,N_11175,N_10395);
nor U13649 (N_13649,N_10097,N_10953);
nand U13650 (N_13650,N_10948,N_11903);
nand U13651 (N_13651,N_11463,N_10005);
nand U13652 (N_13652,N_10218,N_11100);
nand U13653 (N_13653,N_10636,N_11973);
or U13654 (N_13654,N_11597,N_11269);
and U13655 (N_13655,N_11411,N_10920);
nand U13656 (N_13656,N_10193,N_10888);
xnor U13657 (N_13657,N_11921,N_10096);
nor U13658 (N_13658,N_11675,N_11695);
nor U13659 (N_13659,N_10138,N_10722);
and U13660 (N_13660,N_10950,N_11315);
or U13661 (N_13661,N_11105,N_10720);
nand U13662 (N_13662,N_10044,N_10105);
xor U13663 (N_13663,N_10321,N_10009);
xnor U13664 (N_13664,N_10615,N_10590);
and U13665 (N_13665,N_10009,N_10199);
or U13666 (N_13666,N_11281,N_10453);
and U13667 (N_13667,N_10942,N_11021);
and U13668 (N_13668,N_10086,N_10990);
and U13669 (N_13669,N_10881,N_10833);
or U13670 (N_13670,N_10763,N_10469);
nor U13671 (N_13671,N_10684,N_10976);
xor U13672 (N_13672,N_11828,N_10245);
xor U13673 (N_13673,N_10311,N_11430);
xnor U13674 (N_13674,N_11670,N_11566);
nand U13675 (N_13675,N_10122,N_11973);
nand U13676 (N_13676,N_11253,N_10437);
or U13677 (N_13677,N_11344,N_11119);
xor U13678 (N_13678,N_11400,N_10667);
or U13679 (N_13679,N_11535,N_11090);
xnor U13680 (N_13680,N_11255,N_10229);
nor U13681 (N_13681,N_10587,N_11395);
xnor U13682 (N_13682,N_11754,N_10772);
or U13683 (N_13683,N_11046,N_11699);
and U13684 (N_13684,N_11127,N_10822);
xnor U13685 (N_13685,N_10046,N_11453);
nand U13686 (N_13686,N_11579,N_10994);
nand U13687 (N_13687,N_10182,N_10300);
and U13688 (N_13688,N_11297,N_11016);
and U13689 (N_13689,N_11645,N_10277);
or U13690 (N_13690,N_11680,N_10772);
nand U13691 (N_13691,N_11648,N_11373);
or U13692 (N_13692,N_10489,N_10676);
and U13693 (N_13693,N_11460,N_10877);
nor U13694 (N_13694,N_11395,N_11721);
xor U13695 (N_13695,N_11294,N_11968);
xor U13696 (N_13696,N_11633,N_10133);
or U13697 (N_13697,N_11389,N_10410);
xnor U13698 (N_13698,N_11068,N_10925);
xnor U13699 (N_13699,N_11460,N_10283);
nor U13700 (N_13700,N_11908,N_11447);
or U13701 (N_13701,N_10717,N_11745);
nor U13702 (N_13702,N_11467,N_10353);
nand U13703 (N_13703,N_10447,N_10887);
nand U13704 (N_13704,N_11785,N_11847);
xor U13705 (N_13705,N_11977,N_11403);
or U13706 (N_13706,N_11236,N_11260);
nand U13707 (N_13707,N_10649,N_10942);
nor U13708 (N_13708,N_10259,N_11230);
nand U13709 (N_13709,N_10257,N_10190);
xor U13710 (N_13710,N_10796,N_10634);
or U13711 (N_13711,N_10864,N_10647);
and U13712 (N_13712,N_10711,N_10438);
nand U13713 (N_13713,N_10020,N_11992);
or U13714 (N_13714,N_11669,N_10813);
nor U13715 (N_13715,N_10030,N_10372);
xor U13716 (N_13716,N_11953,N_11815);
or U13717 (N_13717,N_11630,N_10172);
and U13718 (N_13718,N_10585,N_11451);
and U13719 (N_13719,N_10813,N_11153);
xor U13720 (N_13720,N_10658,N_10441);
nand U13721 (N_13721,N_11221,N_11016);
nor U13722 (N_13722,N_10604,N_10531);
nor U13723 (N_13723,N_11855,N_11754);
and U13724 (N_13724,N_11446,N_10267);
nand U13725 (N_13725,N_10624,N_10047);
nand U13726 (N_13726,N_11637,N_11181);
nor U13727 (N_13727,N_11352,N_11001);
or U13728 (N_13728,N_11180,N_10279);
nor U13729 (N_13729,N_10053,N_11413);
and U13730 (N_13730,N_10896,N_10579);
nor U13731 (N_13731,N_10188,N_11873);
nor U13732 (N_13732,N_10208,N_11984);
and U13733 (N_13733,N_10322,N_11312);
nor U13734 (N_13734,N_11948,N_11776);
nor U13735 (N_13735,N_11582,N_11153);
or U13736 (N_13736,N_10284,N_10513);
and U13737 (N_13737,N_10241,N_11360);
nand U13738 (N_13738,N_11233,N_10476);
and U13739 (N_13739,N_11728,N_11617);
xor U13740 (N_13740,N_11291,N_11103);
nand U13741 (N_13741,N_11749,N_11649);
and U13742 (N_13742,N_11445,N_11530);
nand U13743 (N_13743,N_10464,N_11107);
and U13744 (N_13744,N_11758,N_10294);
or U13745 (N_13745,N_11855,N_11385);
nand U13746 (N_13746,N_10582,N_11148);
nor U13747 (N_13747,N_10593,N_10470);
and U13748 (N_13748,N_10576,N_11061);
nor U13749 (N_13749,N_10214,N_10960);
xor U13750 (N_13750,N_10763,N_11321);
nand U13751 (N_13751,N_11486,N_11159);
nand U13752 (N_13752,N_10946,N_11950);
or U13753 (N_13753,N_10476,N_11109);
xnor U13754 (N_13754,N_10006,N_11620);
nor U13755 (N_13755,N_11388,N_11453);
or U13756 (N_13756,N_10147,N_10628);
nor U13757 (N_13757,N_11572,N_10201);
and U13758 (N_13758,N_10464,N_11097);
nor U13759 (N_13759,N_11369,N_10923);
or U13760 (N_13760,N_11004,N_10236);
and U13761 (N_13761,N_11025,N_10305);
or U13762 (N_13762,N_10704,N_10457);
nand U13763 (N_13763,N_10020,N_11790);
and U13764 (N_13764,N_11814,N_10505);
nor U13765 (N_13765,N_10615,N_11375);
and U13766 (N_13766,N_10074,N_11613);
xor U13767 (N_13767,N_10097,N_11447);
nor U13768 (N_13768,N_11307,N_11170);
nor U13769 (N_13769,N_10797,N_10376);
xor U13770 (N_13770,N_10286,N_10678);
and U13771 (N_13771,N_11365,N_11422);
or U13772 (N_13772,N_11767,N_11798);
nand U13773 (N_13773,N_10250,N_10195);
nor U13774 (N_13774,N_11230,N_10862);
nand U13775 (N_13775,N_10288,N_11215);
nand U13776 (N_13776,N_11195,N_11296);
nand U13777 (N_13777,N_10499,N_11917);
xor U13778 (N_13778,N_10718,N_10411);
nor U13779 (N_13779,N_11154,N_10498);
xor U13780 (N_13780,N_10458,N_11442);
nand U13781 (N_13781,N_11107,N_11188);
or U13782 (N_13782,N_11027,N_10233);
xor U13783 (N_13783,N_11463,N_11329);
nand U13784 (N_13784,N_11385,N_10353);
and U13785 (N_13785,N_10294,N_11244);
or U13786 (N_13786,N_11985,N_11692);
and U13787 (N_13787,N_10410,N_11525);
and U13788 (N_13788,N_10815,N_10878);
and U13789 (N_13789,N_10636,N_10499);
xor U13790 (N_13790,N_11335,N_11462);
nand U13791 (N_13791,N_10042,N_11032);
xor U13792 (N_13792,N_11622,N_11476);
nor U13793 (N_13793,N_10594,N_11552);
and U13794 (N_13794,N_11683,N_10571);
nor U13795 (N_13795,N_11876,N_11596);
or U13796 (N_13796,N_11179,N_11690);
xor U13797 (N_13797,N_10056,N_11369);
nand U13798 (N_13798,N_11042,N_11149);
or U13799 (N_13799,N_11333,N_10416);
nor U13800 (N_13800,N_10661,N_11370);
nand U13801 (N_13801,N_10452,N_10647);
nand U13802 (N_13802,N_10061,N_10318);
and U13803 (N_13803,N_10658,N_11737);
or U13804 (N_13804,N_10954,N_10979);
xor U13805 (N_13805,N_10809,N_10206);
or U13806 (N_13806,N_10726,N_10070);
and U13807 (N_13807,N_10703,N_11077);
nand U13808 (N_13808,N_10334,N_10404);
nand U13809 (N_13809,N_10974,N_10490);
nand U13810 (N_13810,N_10492,N_10889);
xnor U13811 (N_13811,N_10751,N_10748);
or U13812 (N_13812,N_10155,N_10208);
and U13813 (N_13813,N_10657,N_10003);
xnor U13814 (N_13814,N_11613,N_11964);
xnor U13815 (N_13815,N_10815,N_11837);
or U13816 (N_13816,N_10951,N_10173);
or U13817 (N_13817,N_10101,N_11492);
or U13818 (N_13818,N_10198,N_10823);
and U13819 (N_13819,N_11736,N_11919);
or U13820 (N_13820,N_11158,N_10842);
and U13821 (N_13821,N_11251,N_10513);
and U13822 (N_13822,N_11380,N_10717);
or U13823 (N_13823,N_11371,N_10285);
nand U13824 (N_13824,N_11688,N_11942);
nand U13825 (N_13825,N_11791,N_10938);
or U13826 (N_13826,N_11701,N_10659);
xor U13827 (N_13827,N_11502,N_10452);
and U13828 (N_13828,N_11604,N_11729);
nor U13829 (N_13829,N_11747,N_11173);
and U13830 (N_13830,N_11037,N_11575);
or U13831 (N_13831,N_10183,N_10268);
and U13832 (N_13832,N_10093,N_11360);
or U13833 (N_13833,N_11201,N_11908);
or U13834 (N_13834,N_10446,N_10319);
nand U13835 (N_13835,N_10087,N_10322);
xor U13836 (N_13836,N_10740,N_10202);
nor U13837 (N_13837,N_11770,N_10016);
nand U13838 (N_13838,N_10759,N_10381);
xnor U13839 (N_13839,N_11804,N_10335);
xnor U13840 (N_13840,N_10375,N_11616);
nand U13841 (N_13841,N_10695,N_10164);
nand U13842 (N_13842,N_10580,N_10792);
or U13843 (N_13843,N_11199,N_10941);
nor U13844 (N_13844,N_10835,N_10229);
or U13845 (N_13845,N_11006,N_10835);
or U13846 (N_13846,N_11809,N_11470);
nand U13847 (N_13847,N_11558,N_10479);
or U13848 (N_13848,N_11220,N_11611);
and U13849 (N_13849,N_10660,N_11967);
xnor U13850 (N_13850,N_10434,N_11984);
and U13851 (N_13851,N_10388,N_10171);
nand U13852 (N_13852,N_11609,N_11386);
or U13853 (N_13853,N_11000,N_10933);
or U13854 (N_13854,N_10402,N_11163);
nor U13855 (N_13855,N_10715,N_11293);
and U13856 (N_13856,N_11609,N_11248);
nand U13857 (N_13857,N_11848,N_10893);
nor U13858 (N_13858,N_11641,N_10671);
or U13859 (N_13859,N_11413,N_11859);
and U13860 (N_13860,N_10965,N_11324);
nor U13861 (N_13861,N_10712,N_11607);
and U13862 (N_13862,N_11823,N_10065);
xnor U13863 (N_13863,N_11438,N_10010);
or U13864 (N_13864,N_10521,N_10263);
and U13865 (N_13865,N_10903,N_11614);
nor U13866 (N_13866,N_10251,N_10239);
nand U13867 (N_13867,N_11311,N_10229);
nor U13868 (N_13868,N_11139,N_11475);
and U13869 (N_13869,N_11747,N_10212);
nand U13870 (N_13870,N_10364,N_10611);
xnor U13871 (N_13871,N_10516,N_10495);
and U13872 (N_13872,N_11919,N_10793);
nor U13873 (N_13873,N_11627,N_11688);
xor U13874 (N_13874,N_10844,N_11814);
nor U13875 (N_13875,N_10037,N_11749);
and U13876 (N_13876,N_10081,N_10706);
xor U13877 (N_13877,N_11014,N_10767);
or U13878 (N_13878,N_10276,N_10108);
and U13879 (N_13879,N_10297,N_10765);
nor U13880 (N_13880,N_10851,N_11446);
nor U13881 (N_13881,N_11442,N_10722);
nor U13882 (N_13882,N_10273,N_10327);
and U13883 (N_13883,N_11847,N_10381);
or U13884 (N_13884,N_11640,N_11267);
or U13885 (N_13885,N_10005,N_10007);
nand U13886 (N_13886,N_11124,N_10971);
xnor U13887 (N_13887,N_11372,N_11423);
or U13888 (N_13888,N_11244,N_11422);
xnor U13889 (N_13889,N_10847,N_11074);
nor U13890 (N_13890,N_11803,N_10202);
xnor U13891 (N_13891,N_11286,N_10256);
or U13892 (N_13892,N_10211,N_11055);
or U13893 (N_13893,N_11791,N_11523);
xor U13894 (N_13894,N_10901,N_10595);
or U13895 (N_13895,N_11984,N_10711);
xor U13896 (N_13896,N_10919,N_11699);
nand U13897 (N_13897,N_10373,N_11580);
xnor U13898 (N_13898,N_10899,N_10631);
xor U13899 (N_13899,N_11828,N_10974);
or U13900 (N_13900,N_10115,N_10540);
nand U13901 (N_13901,N_11031,N_11532);
and U13902 (N_13902,N_10085,N_11432);
nand U13903 (N_13903,N_10260,N_11938);
xor U13904 (N_13904,N_11076,N_11126);
nand U13905 (N_13905,N_10603,N_11216);
and U13906 (N_13906,N_11497,N_11593);
or U13907 (N_13907,N_10683,N_11334);
xor U13908 (N_13908,N_10500,N_10428);
or U13909 (N_13909,N_11718,N_11277);
or U13910 (N_13910,N_11003,N_10169);
and U13911 (N_13911,N_10258,N_11837);
nand U13912 (N_13912,N_10523,N_11361);
xnor U13913 (N_13913,N_11894,N_10168);
nor U13914 (N_13914,N_11229,N_11763);
nor U13915 (N_13915,N_11510,N_11485);
xor U13916 (N_13916,N_10296,N_11635);
nand U13917 (N_13917,N_11978,N_11417);
xnor U13918 (N_13918,N_11656,N_11128);
and U13919 (N_13919,N_11054,N_10527);
and U13920 (N_13920,N_10298,N_11287);
nor U13921 (N_13921,N_11276,N_10402);
xnor U13922 (N_13922,N_10273,N_11800);
nor U13923 (N_13923,N_11183,N_10667);
nand U13924 (N_13924,N_10086,N_10217);
nand U13925 (N_13925,N_10196,N_11775);
nor U13926 (N_13926,N_10227,N_10051);
and U13927 (N_13927,N_10721,N_11672);
nor U13928 (N_13928,N_10321,N_11536);
xnor U13929 (N_13929,N_11399,N_11609);
or U13930 (N_13930,N_11764,N_11194);
and U13931 (N_13931,N_11413,N_10252);
or U13932 (N_13932,N_11281,N_10477);
nand U13933 (N_13933,N_10663,N_11664);
xnor U13934 (N_13934,N_10141,N_11917);
nor U13935 (N_13935,N_11634,N_11623);
and U13936 (N_13936,N_10222,N_11730);
and U13937 (N_13937,N_10658,N_11261);
and U13938 (N_13938,N_10016,N_10699);
and U13939 (N_13939,N_10955,N_10676);
or U13940 (N_13940,N_11935,N_10116);
xnor U13941 (N_13941,N_11849,N_10739);
nand U13942 (N_13942,N_11595,N_10841);
xor U13943 (N_13943,N_10621,N_10516);
or U13944 (N_13944,N_10649,N_11055);
or U13945 (N_13945,N_11616,N_10223);
or U13946 (N_13946,N_10218,N_10350);
nand U13947 (N_13947,N_11201,N_11092);
nand U13948 (N_13948,N_10741,N_10851);
nor U13949 (N_13949,N_10309,N_11932);
xnor U13950 (N_13950,N_10944,N_11085);
nand U13951 (N_13951,N_10632,N_10950);
and U13952 (N_13952,N_10211,N_10717);
nand U13953 (N_13953,N_11130,N_10225);
nor U13954 (N_13954,N_11061,N_10764);
nor U13955 (N_13955,N_11433,N_10267);
xnor U13956 (N_13956,N_11696,N_11281);
and U13957 (N_13957,N_10525,N_10817);
nand U13958 (N_13958,N_11874,N_11627);
and U13959 (N_13959,N_10863,N_11273);
and U13960 (N_13960,N_11519,N_10484);
xor U13961 (N_13961,N_11070,N_11062);
xnor U13962 (N_13962,N_11855,N_11400);
nand U13963 (N_13963,N_11609,N_10090);
or U13964 (N_13964,N_11408,N_11765);
nor U13965 (N_13965,N_10760,N_11785);
xnor U13966 (N_13966,N_10215,N_10218);
and U13967 (N_13967,N_10571,N_10676);
nor U13968 (N_13968,N_10226,N_10221);
or U13969 (N_13969,N_11285,N_11748);
nand U13970 (N_13970,N_11687,N_10606);
and U13971 (N_13971,N_10936,N_10561);
or U13972 (N_13972,N_11757,N_10680);
nand U13973 (N_13973,N_11630,N_10521);
nand U13974 (N_13974,N_10062,N_11355);
nand U13975 (N_13975,N_10800,N_11950);
or U13976 (N_13976,N_11607,N_11156);
xnor U13977 (N_13977,N_11892,N_10197);
and U13978 (N_13978,N_10889,N_10368);
nand U13979 (N_13979,N_10118,N_11578);
or U13980 (N_13980,N_11431,N_11470);
or U13981 (N_13981,N_11553,N_10394);
nand U13982 (N_13982,N_11499,N_10188);
xor U13983 (N_13983,N_11167,N_10216);
nor U13984 (N_13984,N_10447,N_11876);
nor U13985 (N_13985,N_10915,N_11384);
or U13986 (N_13986,N_11757,N_10507);
nand U13987 (N_13987,N_11727,N_10874);
nor U13988 (N_13988,N_11167,N_11513);
nor U13989 (N_13989,N_10784,N_10887);
xnor U13990 (N_13990,N_10811,N_10808);
nand U13991 (N_13991,N_10688,N_11584);
nor U13992 (N_13992,N_10977,N_11763);
and U13993 (N_13993,N_11334,N_10634);
or U13994 (N_13994,N_11046,N_10585);
nor U13995 (N_13995,N_10041,N_11188);
and U13996 (N_13996,N_11197,N_11209);
xor U13997 (N_13997,N_10659,N_11346);
nor U13998 (N_13998,N_11931,N_11620);
or U13999 (N_13999,N_11850,N_10720);
nand U14000 (N_14000,N_13892,N_12554);
nor U14001 (N_14001,N_12144,N_12056);
nor U14002 (N_14002,N_13218,N_12289);
or U14003 (N_14003,N_12116,N_12307);
nor U14004 (N_14004,N_13247,N_13314);
xnor U14005 (N_14005,N_12372,N_12716);
nor U14006 (N_14006,N_12294,N_13684);
nand U14007 (N_14007,N_12113,N_12445);
nor U14008 (N_14008,N_12215,N_13301);
nor U14009 (N_14009,N_12744,N_13741);
nand U14010 (N_14010,N_12933,N_13309);
or U14011 (N_14011,N_12172,N_12351);
nor U14012 (N_14012,N_13780,N_13115);
or U14013 (N_14013,N_13402,N_12325);
nand U14014 (N_14014,N_13491,N_13912);
or U14015 (N_14015,N_13215,N_13047);
nand U14016 (N_14016,N_13583,N_12597);
nor U14017 (N_14017,N_12395,N_13384);
nand U14018 (N_14018,N_12474,N_12441);
xor U14019 (N_14019,N_12678,N_13669);
nand U14020 (N_14020,N_12064,N_13101);
nor U14021 (N_14021,N_12671,N_13067);
xor U14022 (N_14022,N_12539,N_13295);
or U14023 (N_14023,N_12838,N_13578);
nand U14024 (N_14024,N_13958,N_13721);
xnor U14025 (N_14025,N_12428,N_12324);
and U14026 (N_14026,N_12538,N_12879);
nand U14027 (N_14027,N_12305,N_13222);
nand U14028 (N_14028,N_12035,N_12287);
and U14029 (N_14029,N_12656,N_13725);
nand U14030 (N_14030,N_13106,N_13522);
or U14031 (N_14031,N_12313,N_12051);
or U14032 (N_14032,N_13670,N_12980);
and U14033 (N_14033,N_12537,N_12640);
nor U14034 (N_14034,N_12530,N_12863);
and U14035 (N_14035,N_13330,N_12764);
nand U14036 (N_14036,N_13265,N_13751);
and U14037 (N_14037,N_13060,N_13050);
nor U14038 (N_14038,N_13974,N_12438);
nand U14039 (N_14039,N_12948,N_12277);
or U14040 (N_14040,N_13278,N_13369);
xor U14041 (N_14041,N_13723,N_12881);
nor U14042 (N_14042,N_12623,N_13023);
nor U14043 (N_14043,N_13039,N_13948);
xor U14044 (N_14044,N_12505,N_13297);
or U14045 (N_14045,N_12252,N_12932);
xnor U14046 (N_14046,N_13924,N_12513);
xor U14047 (N_14047,N_13416,N_12664);
nand U14048 (N_14048,N_13173,N_13848);
nand U14049 (N_14049,N_13382,N_13433);
xnor U14050 (N_14050,N_13421,N_12048);
or U14051 (N_14051,N_13586,N_13826);
nand U14052 (N_14052,N_13000,N_12194);
or U14053 (N_14053,N_12379,N_13443);
and U14054 (N_14054,N_13571,N_13731);
nor U14055 (N_14055,N_13786,N_12464);
xnor U14056 (N_14056,N_13652,N_12675);
nor U14057 (N_14057,N_13619,N_12618);
xor U14058 (N_14058,N_12951,N_13146);
and U14059 (N_14059,N_13064,N_12390);
xor U14060 (N_14060,N_13094,N_13355);
and U14061 (N_14061,N_13037,N_12126);
or U14062 (N_14062,N_13160,N_13843);
or U14063 (N_14063,N_13654,N_12407);
or U14064 (N_14064,N_13679,N_13362);
xnor U14065 (N_14065,N_13955,N_12225);
xor U14066 (N_14066,N_13434,N_12136);
or U14067 (N_14067,N_12741,N_13941);
nor U14068 (N_14068,N_12058,N_13150);
or U14069 (N_14069,N_13995,N_13557);
nand U14070 (N_14070,N_12853,N_13807);
or U14071 (N_14071,N_12631,N_12532);
nor U14072 (N_14072,N_12080,N_12192);
xnor U14073 (N_14073,N_13599,N_13641);
nor U14074 (N_14074,N_13242,N_12386);
or U14075 (N_14075,N_12273,N_13745);
nor U14076 (N_14076,N_13354,N_13001);
nand U14077 (N_14077,N_12179,N_13187);
and U14078 (N_14078,N_13076,N_12643);
nand U14079 (N_14079,N_13097,N_12016);
nand U14080 (N_14080,N_13823,N_13083);
nor U14081 (N_14081,N_13701,N_12270);
and U14082 (N_14082,N_13482,N_13926);
xor U14083 (N_14083,N_12278,N_13556);
or U14084 (N_14084,N_13647,N_12998);
nand U14085 (N_14085,N_12074,N_12087);
nor U14086 (N_14086,N_13987,N_12706);
nand U14087 (N_14087,N_13748,N_13660);
xnor U14088 (N_14088,N_13612,N_13928);
nor U14089 (N_14089,N_12828,N_13322);
nand U14090 (N_14090,N_12495,N_13841);
or U14091 (N_14091,N_13026,N_12686);
xnor U14092 (N_14092,N_12490,N_13051);
nand U14093 (N_14093,N_12806,N_13874);
nor U14094 (N_14094,N_13320,N_13676);
nor U14095 (N_14095,N_13850,N_12634);
nor U14096 (N_14096,N_12920,N_12430);
nand U14097 (N_14097,N_13856,N_13582);
nand U14098 (N_14098,N_12272,N_13473);
or U14099 (N_14099,N_13165,N_12213);
and U14100 (N_14100,N_12384,N_13161);
nor U14101 (N_14101,N_13639,N_13925);
nand U14102 (N_14102,N_13842,N_12545);
and U14103 (N_14103,N_12067,N_13738);
and U14104 (N_14104,N_12024,N_13609);
nand U14105 (N_14105,N_13481,N_13153);
nand U14106 (N_14106,N_12284,N_12915);
nand U14107 (N_14107,N_12349,N_12825);
nand U14108 (N_14108,N_13517,N_13539);
nor U14109 (N_14109,N_13552,N_13216);
nor U14110 (N_14110,N_13888,N_12504);
or U14111 (N_14111,N_13922,N_13290);
and U14112 (N_14112,N_13866,N_13159);
nand U14113 (N_14113,N_12711,N_12492);
and U14114 (N_14114,N_12217,N_12800);
xor U14115 (N_14115,N_12072,N_13274);
or U14116 (N_14116,N_12952,N_13492);
xor U14117 (N_14117,N_12109,N_12301);
xor U14118 (N_14118,N_13066,N_13464);
and U14119 (N_14119,N_13107,N_13595);
xor U14120 (N_14120,N_12171,N_13308);
and U14121 (N_14121,N_13919,N_12917);
nand U14122 (N_14122,N_12224,N_13622);
and U14123 (N_14123,N_12698,N_12275);
and U14124 (N_14124,N_13770,N_12979);
nor U14125 (N_14125,N_13028,N_13704);
xor U14126 (N_14126,N_13547,N_13880);
nor U14127 (N_14127,N_12646,N_13335);
or U14128 (N_14128,N_13437,N_12615);
xnor U14129 (N_14129,N_13559,N_12935);
xnor U14130 (N_14130,N_12282,N_12667);
xor U14131 (N_14131,N_13813,N_12086);
and U14132 (N_14132,N_12121,N_12839);
or U14133 (N_14133,N_12996,N_12626);
or U14134 (N_14134,N_12169,N_12997);
nand U14135 (N_14135,N_12266,N_13577);
and U14136 (N_14136,N_13913,N_13267);
nand U14137 (N_14137,N_13456,N_12326);
nor U14138 (N_14138,N_13317,N_12883);
and U14139 (N_14139,N_13135,N_12066);
nor U14140 (N_14140,N_13631,N_12258);
or U14141 (N_14141,N_13575,N_12712);
and U14142 (N_14142,N_13773,N_12900);
and U14143 (N_14143,N_12693,N_12755);
or U14144 (N_14144,N_13605,N_13239);
nand U14145 (N_14145,N_13960,N_12143);
nand U14146 (N_14146,N_13746,N_12250);
and U14147 (N_14147,N_13411,N_12904);
xor U14148 (N_14148,N_12279,N_12207);
nand U14149 (N_14149,N_13111,N_12784);
nor U14150 (N_14150,N_13872,N_12185);
xnor U14151 (N_14151,N_12364,N_13142);
or U14152 (N_14152,N_12589,N_13640);
and U14153 (N_14153,N_13678,N_13246);
nor U14154 (N_14154,N_12059,N_12098);
and U14155 (N_14155,N_13140,N_12469);
nor U14156 (N_14156,N_13334,N_12713);
xnor U14157 (N_14157,N_13794,N_13085);
nor U14158 (N_14158,N_13742,N_12359);
nand U14159 (N_14159,N_13304,N_13348);
nor U14160 (N_14160,N_12888,N_12235);
nor U14161 (N_14161,N_12833,N_12902);
xor U14162 (N_14162,N_13923,N_12370);
nand U14163 (N_14163,N_12999,N_13326);
and U14164 (N_14164,N_13835,N_13381);
nand U14165 (N_14165,N_12354,N_12831);
nand U14166 (N_14166,N_12117,N_12984);
nor U14167 (N_14167,N_12779,N_12847);
xnor U14168 (N_14168,N_12174,N_12329);
nor U14169 (N_14169,N_12673,N_12052);
and U14170 (N_14170,N_12734,N_12965);
or U14171 (N_14171,N_13477,N_12756);
nand U14172 (N_14172,N_13680,N_13367);
nand U14173 (N_14173,N_12899,N_12429);
or U14174 (N_14174,N_13011,N_12840);
nor U14175 (N_14175,N_13779,N_12531);
nand U14176 (N_14176,N_13091,N_13021);
and U14177 (N_14177,N_12890,N_12118);
nor U14178 (N_14178,N_13105,N_12160);
or U14179 (N_14179,N_13180,N_13031);
or U14180 (N_14180,N_13802,N_13396);
or U14181 (N_14181,N_13346,N_13128);
nor U14182 (N_14182,N_12168,N_13642);
nand U14183 (N_14183,N_12022,N_13302);
nand U14184 (N_14184,N_13656,N_12241);
or U14185 (N_14185,N_12083,N_13811);
nor U14186 (N_14186,N_13080,N_12070);
and U14187 (N_14187,N_13019,N_12233);
nor U14188 (N_14188,N_13071,N_13562);
xnor U14189 (N_14189,N_12491,N_13401);
nand U14190 (N_14190,N_12891,N_13414);
and U14191 (N_14191,N_13675,N_12494);
or U14192 (N_14192,N_13756,N_13903);
and U14193 (N_14193,N_12226,N_12849);
nand U14194 (N_14194,N_12222,N_12789);
nand U14195 (N_14195,N_13906,N_12201);
or U14196 (N_14196,N_13250,N_12295);
and U14197 (N_14197,N_13988,N_13226);
nand U14198 (N_14198,N_12700,N_12245);
or U14199 (N_14199,N_12666,N_12916);
or U14200 (N_14200,N_12230,N_13677);
nor U14201 (N_14201,N_12662,N_13757);
nor U14202 (N_14202,N_12209,N_13891);
xor U14203 (N_14203,N_13580,N_13363);
or U14204 (N_14204,N_13487,N_13079);
nor U14205 (N_14205,N_12042,N_12312);
xnor U14206 (N_14206,N_12660,N_13234);
or U14207 (N_14207,N_12894,N_13938);
nor U14208 (N_14208,N_12971,N_12846);
and U14209 (N_14209,N_13428,N_13446);
nand U14210 (N_14210,N_12843,N_12638);
or U14211 (N_14211,N_13978,N_12315);
or U14212 (N_14212,N_13409,N_13137);
and U14213 (N_14213,N_12078,N_13185);
nand U14214 (N_14214,N_13495,N_12410);
nand U14215 (N_14215,N_12556,N_13935);
xor U14216 (N_14216,N_12454,N_13531);
and U14217 (N_14217,N_13964,N_13708);
nor U14218 (N_14218,N_13496,N_12013);
xnor U14219 (N_14219,N_13035,N_13550);
nand U14220 (N_14220,N_13342,N_12540);
and U14221 (N_14221,N_13962,N_12647);
or U14222 (N_14222,N_12760,N_13846);
nor U14223 (N_14223,N_13236,N_12196);
xnor U14224 (N_14224,N_12269,N_13458);
xnor U14225 (N_14225,N_12715,N_13244);
nor U14226 (N_14226,N_12925,N_12330);
nor U14227 (N_14227,N_12957,N_13114);
nor U14228 (N_14228,N_12114,N_12021);
nand U14229 (N_14229,N_12824,N_12674);
nor U14230 (N_14230,N_12767,N_12534);
nor U14231 (N_14231,N_13287,N_12099);
or U14232 (N_14232,N_13034,N_13003);
nor U14233 (N_14233,N_13178,N_13144);
nor U14234 (N_14234,N_12865,N_12757);
nand U14235 (N_14235,N_13420,N_13068);
nand U14236 (N_14236,N_12104,N_12140);
and U14237 (N_14237,N_12544,N_12122);
nand U14238 (N_14238,N_13908,N_13617);
and U14239 (N_14239,N_12095,N_12772);
or U14240 (N_14240,N_13388,N_12229);
xor U14241 (N_14241,N_13682,N_12029);
or U14242 (N_14242,N_13610,N_12054);
nor U14243 (N_14243,N_13074,N_12376);
or U14244 (N_14244,N_12723,N_13829);
xnor U14245 (N_14245,N_12399,N_13310);
xnor U14246 (N_14246,N_13073,N_13484);
and U14247 (N_14247,N_13805,N_13549);
nor U14248 (N_14248,N_12096,N_12014);
or U14249 (N_14249,N_13368,N_12347);
xnor U14250 (N_14250,N_13498,N_12341);
xor U14251 (N_14251,N_13306,N_12960);
nor U14252 (N_14252,N_12954,N_13095);
nor U14253 (N_14253,N_12285,N_13327);
and U14254 (N_14254,N_12550,N_12733);
and U14255 (N_14255,N_13257,N_12392);
and U14256 (N_14256,N_12249,N_12721);
or U14257 (N_14257,N_13545,N_13002);
and U14258 (N_14258,N_13581,N_13737);
xor U14259 (N_14259,N_12406,N_12802);
nand U14260 (N_14260,N_12906,N_12856);
nor U14261 (N_14261,N_13956,N_12928);
or U14262 (N_14262,N_13351,N_12963);
nand U14263 (N_14263,N_13664,N_12026);
xor U14264 (N_14264,N_12696,N_12703);
nor U14265 (N_14265,N_13331,N_12527);
nor U14266 (N_14266,N_12821,N_12683);
or U14267 (N_14267,N_13593,N_12497);
nor U14268 (N_14268,N_12896,N_12761);
nand U14269 (N_14269,N_12573,N_12893);
nand U14270 (N_14270,N_12027,N_12866);
nand U14271 (N_14271,N_13120,N_12579);
nand U14272 (N_14272,N_13657,N_13385);
xor U14273 (N_14273,N_12649,N_13131);
nor U14274 (N_14274,N_12553,N_13378);
nor U14275 (N_14275,N_12552,N_12763);
and U14276 (N_14276,N_13585,N_12815);
or U14277 (N_14277,N_13777,N_12134);
or U14278 (N_14278,N_12138,N_13788);
nand U14279 (N_14279,N_13429,N_12751);
or U14280 (N_14280,N_13809,N_13984);
and U14281 (N_14281,N_13444,N_13782);
nor U14282 (N_14282,N_12509,N_13801);
or U14283 (N_14283,N_12841,N_13190);
and U14284 (N_14284,N_12559,N_12938);
xor U14285 (N_14285,N_12470,N_12293);
nand U14286 (N_14286,N_12510,N_13199);
nand U14287 (N_14287,N_12868,N_12154);
and U14288 (N_14288,N_13567,N_12318);
and U14289 (N_14289,N_12017,N_13920);
or U14290 (N_14290,N_13873,N_13383);
and U14291 (N_14291,N_12988,N_13232);
and U14292 (N_14292,N_13439,N_12768);
or U14293 (N_14293,N_13449,N_13992);
and U14294 (N_14294,N_13712,N_13077);
nand U14295 (N_14295,N_12818,N_13293);
or U14296 (N_14296,N_12989,N_13424);
nand U14297 (N_14297,N_12378,N_13589);
nand U14298 (N_14298,N_12486,N_13405);
or U14299 (N_14299,N_13831,N_12685);
nor U14300 (N_14300,N_12858,N_12561);
xnor U14301 (N_14301,N_13740,N_13694);
nand U14302 (N_14302,N_13103,N_12010);
nand U14303 (N_14303,N_13529,N_13436);
xor U14304 (N_14304,N_12898,N_13207);
nand U14305 (N_14305,N_12236,N_12271);
nand U14306 (N_14306,N_13253,N_12323);
and U14307 (N_14307,N_13551,N_13685);
xnor U14308 (N_14308,N_12738,N_13288);
xor U14309 (N_14309,N_13453,N_13600);
xor U14310 (N_14310,N_12343,N_13102);
nor U14311 (N_14311,N_13006,N_13084);
nand U14312 (N_14312,N_13790,N_12165);
or U14313 (N_14313,N_13905,N_12472);
nand U14314 (N_14314,N_13722,N_13460);
xnor U14315 (N_14315,N_13629,N_13849);
and U14316 (N_14316,N_12131,N_13425);
nor U14317 (N_14317,N_13658,N_13315);
nor U14318 (N_14318,N_13300,N_13432);
nor U14319 (N_14319,N_12197,N_12254);
xor U14320 (N_14320,N_13057,N_12216);
nand U14321 (N_14321,N_13294,N_12298);
nand U14322 (N_14322,N_12947,N_12874);
or U14323 (N_14323,N_13882,N_13154);
and U14324 (N_14324,N_12692,N_13603);
xor U14325 (N_14325,N_13747,N_12344);
nand U14326 (N_14326,N_13686,N_13463);
nor U14327 (N_14327,N_13223,N_13230);
xnor U14328 (N_14328,N_13263,N_12882);
nor U14329 (N_14329,N_12003,N_13720);
nand U14330 (N_14330,N_13797,N_12419);
nor U14331 (N_14331,N_13010,N_12599);
nand U14332 (N_14332,N_13999,N_13323);
nor U14333 (N_14333,N_13467,N_13096);
and U14334 (N_14334,N_12455,N_13784);
or U14335 (N_14335,N_12220,N_12986);
and U14336 (N_14336,N_13285,N_12268);
nand U14337 (N_14337,N_12875,N_13252);
or U14338 (N_14338,N_12246,N_13918);
and U14339 (N_14339,N_13847,N_13134);
nand U14340 (N_14340,N_12210,N_12519);
nor U14341 (N_14341,N_12465,N_13177);
nor U14342 (N_14342,N_12542,N_12630);
or U14343 (N_14343,N_12089,N_13181);
or U14344 (N_14344,N_13466,N_12422);
or U14345 (N_14345,N_12961,N_13715);
or U14346 (N_14346,N_12237,N_12115);
nand U14347 (N_14347,N_13220,N_12672);
xor U14348 (N_14348,N_12091,N_13778);
xor U14349 (N_14349,N_12357,N_13868);
nand U14350 (N_14350,N_13447,N_13957);
nor U14351 (N_14351,N_13005,N_12790);
nand U14352 (N_14352,N_12857,N_13927);
nor U14353 (N_14353,N_12191,N_13167);
and U14354 (N_14354,N_12476,N_13441);
and U14355 (N_14355,N_12619,N_13902);
and U14356 (N_14356,N_12990,N_13804);
nor U14357 (N_14357,N_12020,N_12062);
and U14358 (N_14358,N_12684,N_12468);
and U14359 (N_14359,N_13865,N_13755);
nor U14360 (N_14360,N_13929,N_12974);
and U14361 (N_14361,N_12887,N_12467);
or U14362 (N_14362,N_13387,N_13053);
xor U14363 (N_14363,N_12132,N_12023);
xnor U14364 (N_14364,N_12608,N_13705);
nor U14365 (N_14365,N_13611,N_13130);
or U14366 (N_14366,N_12565,N_12823);
or U14367 (N_14367,N_12025,N_12926);
nand U14368 (N_14368,N_13587,N_13148);
xnor U14369 (N_14369,N_12931,N_13337);
xor U14370 (N_14370,N_13238,N_12255);
xor U14371 (N_14371,N_12358,N_12423);
xnor U14372 (N_14372,N_12367,N_13196);
nand U14373 (N_14373,N_12817,N_12369);
nor U14374 (N_14374,N_13340,N_12940);
and U14375 (N_14375,N_12570,N_13022);
nand U14376 (N_14376,N_12500,N_12304);
and U14377 (N_14377,N_12004,N_12077);
and U14378 (N_14378,N_12777,N_12133);
or U14379 (N_14379,N_13931,N_13833);
nor U14380 (N_14380,N_13404,N_12718);
nand U14381 (N_14381,N_12600,N_13965);
nand U14382 (N_14382,N_12097,N_13266);
and U14383 (N_14383,N_12264,N_13151);
xor U14384 (N_14384,N_12611,N_12598);
xnor U14385 (N_14385,N_12409,N_12652);
and U14386 (N_14386,N_13681,N_13270);
or U14387 (N_14387,N_12995,N_13949);
nand U14388 (N_14388,N_12199,N_13769);
and U14389 (N_14389,N_13659,N_12927);
xnor U14390 (N_14390,N_13109,N_13934);
nor U14391 (N_14391,N_13976,N_12012);
nand U14392 (N_14392,N_12176,N_13776);
xor U14393 (N_14393,N_12994,N_13372);
and U14394 (N_14394,N_12234,N_12411);
xor U14395 (N_14395,N_12642,N_12198);
nor U14396 (N_14396,N_12944,N_13243);
and U14397 (N_14397,N_13697,N_13889);
or U14398 (N_14398,N_13235,N_13799);
nand U14399 (N_14399,N_13344,N_12895);
xnor U14400 (N_14400,N_13158,N_12415);
xor U14401 (N_14401,N_13009,N_12039);
and U14402 (N_14402,N_12516,N_12381);
or U14403 (N_14403,N_13004,N_12690);
xor U14404 (N_14404,N_13325,N_13395);
or U14405 (N_14405,N_13281,N_13933);
or U14406 (N_14406,N_13982,N_13370);
nand U14407 (N_14407,N_13486,N_12725);
and U14408 (N_14408,N_12005,N_13568);
or U14409 (N_14409,N_12501,N_13426);
xnor U14410 (N_14410,N_12568,N_13818);
nand U14411 (N_14411,N_13695,N_13289);
and U14412 (N_14412,N_13968,N_13621);
nand U14413 (N_14413,N_12854,N_12212);
xor U14414 (N_14414,N_13648,N_12475);
nor U14415 (N_14415,N_12443,N_13358);
or U14416 (N_14416,N_13909,N_13885);
nand U14417 (N_14417,N_13798,N_13018);
or U14418 (N_14418,N_12396,N_12752);
nand U14419 (N_14419,N_12582,N_13427);
xnor U14420 (N_14420,N_12383,N_13620);
xor U14421 (N_14421,N_12111,N_13566);
nor U14422 (N_14422,N_13832,N_13890);
nand U14423 (N_14423,N_13979,N_12480);
nor U14424 (N_14424,N_12334,N_12651);
nor U14425 (N_14425,N_13376,N_12801);
and U14426 (N_14426,N_13089,N_13570);
xor U14427 (N_14427,N_12253,N_12574);
xnor U14428 (N_14428,N_12248,N_12170);
or U14429 (N_14429,N_12414,N_12417);
or U14430 (N_14430,N_13635,N_12361);
and U14431 (N_14431,N_13380,N_13534);
xnor U14432 (N_14432,N_13069,N_12541);
nor U14433 (N_14433,N_13020,N_13328);
xor U14434 (N_14434,N_12560,N_12496);
nor U14435 (N_14435,N_13126,N_13350);
xnor U14436 (N_14436,N_12549,N_12232);
xnor U14437 (N_14437,N_13646,N_12622);
or U14438 (N_14438,N_13584,N_13508);
nor U14439 (N_14439,N_13506,N_13863);
and U14440 (N_14440,N_13468,N_12112);
nor U14441 (N_14441,N_12930,N_13391);
xor U14442 (N_14442,N_12444,N_13942);
nor U14443 (N_14443,N_12202,N_13186);
or U14444 (N_14444,N_12884,N_12949);
and U14445 (N_14445,N_13632,N_12695);
nor U14446 (N_14446,N_12106,N_12807);
or U14447 (N_14447,N_13707,N_12180);
nand U14448 (N_14448,N_13643,N_13081);
xor U14449 (N_14449,N_13781,N_12082);
nand U14450 (N_14450,N_13046,N_12985);
and U14451 (N_14451,N_13078,N_12593);
or U14452 (N_14452,N_13900,N_13717);
or U14453 (N_14453,N_13027,N_13633);
and U14454 (N_14454,N_12290,N_12507);
nand U14455 (N_14455,N_12719,N_12867);
nor U14456 (N_14456,N_12694,N_12466);
xnor U14457 (N_14457,N_13744,N_12736);
and U14458 (N_14458,N_12488,N_12645);
nor U14459 (N_14459,N_13406,N_13822);
and U14460 (N_14460,N_12300,N_13854);
nor U14461 (N_14461,N_13129,N_12546);
nor U14462 (N_14462,N_12173,N_13538);
and U14463 (N_14463,N_12870,N_13113);
and U14464 (N_14464,N_12969,N_12418);
xnor U14465 (N_14465,N_13602,N_12748);
xnor U14466 (N_14466,N_13674,N_13700);
or U14467 (N_14467,N_12592,N_13961);
nor U14468 (N_14468,N_12148,N_13087);
nor U14469 (N_14469,N_13937,N_12363);
and U14470 (N_14470,N_12605,N_12810);
nor U14471 (N_14471,N_13993,N_12781);
and U14472 (N_14472,N_13554,N_13896);
xnor U14473 (N_14473,N_13510,N_13591);
xnor U14474 (N_14474,N_13911,N_13616);
and U14475 (N_14475,N_12071,N_12730);
nor U14476 (N_14476,N_12548,N_12088);
nand U14477 (N_14477,N_13282,N_13791);
and U14478 (N_14478,N_13512,N_13398);
nand U14479 (N_14479,N_12337,N_13785);
nand U14480 (N_14480,N_13973,N_13361);
nor U14481 (N_14481,N_12448,N_13763);
nand U14482 (N_14482,N_12911,N_12613);
nor U14483 (N_14483,N_13830,N_13431);
nor U14484 (N_14484,N_13504,N_13663);
nand U14485 (N_14485,N_12322,N_12040);
xor U14486 (N_14486,N_13172,N_13219);
and U14487 (N_14487,N_12090,N_12518);
nor U14488 (N_14488,N_12795,N_12243);
and U14489 (N_14489,N_13224,N_12769);
xnor U14490 (N_14490,N_12065,N_13795);
nor U14491 (N_14491,N_13975,N_13284);
nand U14492 (N_14492,N_13542,N_13500);
nor U14493 (N_14493,N_12657,N_12805);
nor U14494 (N_14494,N_13838,N_12528);
nor U14495 (N_14495,N_12621,N_13099);
nor U14496 (N_14496,N_13417,N_13688);
nand U14497 (N_14497,N_13377,N_12835);
xnor U14498 (N_14498,N_13479,N_13360);
nor U14499 (N_14499,N_12680,N_12166);
nand U14500 (N_14500,N_12231,N_12585);
xnor U14501 (N_14501,N_12950,N_13227);
nor U14502 (N_14502,N_13897,N_12914);
xor U14503 (N_14503,N_13469,N_12976);
and U14504 (N_14504,N_12130,N_13726);
or U14505 (N_14505,N_12362,N_12595);
xnor U14506 (N_14506,N_12333,N_12446);
nor U14507 (N_14507,N_13191,N_13536);
nor U14508 (N_14508,N_13043,N_13606);
nand U14509 (N_14509,N_12859,N_12830);
or U14510 (N_14510,N_12778,N_13604);
nor U14511 (N_14511,N_13374,N_13225);
and U14512 (N_14512,N_13025,N_12829);
or U14513 (N_14513,N_13193,N_13171);
or U14514 (N_14514,N_12567,N_12814);
or U14515 (N_14515,N_12918,N_12729);
xnor U14516 (N_14516,N_13261,N_13319);
or U14517 (N_14517,N_13530,N_13162);
xnor U14518 (N_14518,N_12221,N_12263);
xor U14519 (N_14519,N_12002,N_13352);
nand U14520 (N_14520,N_12261,N_13108);
and U14521 (N_14521,N_12485,N_12970);
nor U14522 (N_14522,N_12754,N_12602);
and U14523 (N_14523,N_12483,N_13208);
nand U14524 (N_14524,N_12412,N_12331);
nand U14525 (N_14525,N_13662,N_12584);
nand U14526 (N_14526,N_12762,N_12204);
xor U14527 (N_14527,N_12163,N_13553);
or U14528 (N_14528,N_12257,N_12208);
xor U14529 (N_14529,N_12811,N_13163);
xor U14530 (N_14530,N_12937,N_13119);
nand U14531 (N_14531,N_13470,N_12770);
and U14532 (N_14532,N_13012,N_12434);
nor U14533 (N_14533,N_12691,N_12400);
nand U14534 (N_14534,N_12151,N_12791);
and U14535 (N_14535,N_13977,N_13438);
nand U14536 (N_14536,N_12792,N_13630);
xor U14537 (N_14537,N_12705,N_13292);
nand U14538 (N_14538,N_13264,N_13524);
and U14539 (N_14539,N_12687,N_12129);
and U14540 (N_14540,N_12377,N_12031);
nand U14541 (N_14541,N_12008,N_12119);
xor U14542 (N_14542,N_12648,N_13655);
nand U14543 (N_14543,N_12603,N_13296);
nor U14544 (N_14544,N_12627,N_13932);
nand U14545 (N_14545,N_12872,N_13014);
nand U14546 (N_14546,N_13572,N_12819);
and U14547 (N_14547,N_12590,N_13910);
or U14548 (N_14548,N_13514,N_13251);
xnor U14549 (N_14549,N_13200,N_12663);
xor U14550 (N_14550,N_13279,N_12826);
or U14551 (N_14551,N_12808,N_13944);
nand U14552 (N_14552,N_13750,N_13418);
xnor U14553 (N_14553,N_13347,N_13859);
xnor U14554 (N_14554,N_12569,N_13951);
nand U14555 (N_14555,N_12028,N_13869);
nor U14556 (N_14556,N_13070,N_13543);
and U14557 (N_14557,N_12260,N_12743);
nand U14558 (N_14558,N_12668,N_12387);
and U14559 (N_14559,N_13893,N_13526);
nor U14560 (N_14560,N_13164,N_12836);
or U14561 (N_14561,N_12676,N_12520);
nor U14562 (N_14562,N_13573,N_12426);
and U14563 (N_14563,N_13170,N_12750);
and U14564 (N_14564,N_12084,N_12616);
or U14565 (N_14565,N_13359,N_13898);
and U14566 (N_14566,N_13939,N_12845);
and U14567 (N_14567,N_13861,N_13489);
or U14568 (N_14568,N_13752,N_13179);
nand U14569 (N_14569,N_12793,N_13967);
nor U14570 (N_14570,N_12759,N_12972);
and U14571 (N_14571,N_13558,N_13714);
nor U14572 (N_14572,N_13201,N_12809);
nor U14573 (N_14573,N_13241,N_13249);
xnor U14574 (N_14574,N_13313,N_13415);
or U14575 (N_14575,N_12624,N_13561);
nor U14576 (N_14576,N_13189,N_12975);
and U14577 (N_14577,N_12205,N_12368);
nor U14578 (N_14578,N_12787,N_12371);
nand U14579 (N_14579,N_13963,N_12463);
nor U14580 (N_14580,N_13272,N_13936);
nor U14581 (N_14581,N_13299,N_13412);
xnor U14582 (N_14582,N_13753,N_13277);
nor U14583 (N_14583,N_13775,N_13403);
xnor U14584 (N_14584,N_12742,N_13845);
or U14585 (N_14585,N_12327,N_13623);
or U14586 (N_14586,N_12350,N_13445);
xor U14587 (N_14587,N_12447,N_13981);
nor U14588 (N_14588,N_13462,N_12484);
nor U14589 (N_14589,N_12162,N_12036);
nor U14590 (N_14590,N_12296,N_12922);
xor U14591 (N_14591,N_13886,N_12566);
nand U14592 (N_14592,N_12709,N_13423);
nor U14593 (N_14593,N_12735,N_12482);
and U14594 (N_14594,N_13548,N_13182);
and U14595 (N_14595,N_13132,N_13810);
or U14596 (N_14596,N_12717,N_13271);
and U14597 (N_14597,N_13455,N_12697);
and U14598 (N_14598,N_13564,N_13152);
xor U14599 (N_14599,N_13059,N_13389);
and U14600 (N_14600,N_13597,N_13860);
nand U14601 (N_14601,N_12873,N_12966);
nand U14602 (N_14602,N_12732,N_13055);
xnor U14603 (N_14603,N_13197,N_13240);
nand U14604 (N_14604,N_13221,N_13749);
or U14605 (N_14605,N_12720,N_12228);
nand U14606 (N_14606,N_13793,N_12489);
nor U14607 (N_14607,N_13138,N_13194);
nor U14608 (N_14608,N_12594,N_13036);
xnor U14609 (N_14609,N_13666,N_12726);
xor U14610 (N_14610,N_12728,N_13590);
nor U14611 (N_14611,N_13237,N_12432);
and U14612 (N_14612,N_13147,N_13817);
xnor U14613 (N_14613,N_13739,N_12308);
nor U14614 (N_14614,N_13341,N_12385);
and U14615 (N_14615,N_12178,N_12661);
or U14616 (N_14616,N_13947,N_12079);
and U14617 (N_14617,N_12547,N_12473);
xnor U14618 (N_14618,N_12905,N_13175);
xnor U14619 (N_14619,N_12788,N_12158);
and U14620 (N_14620,N_12451,N_12749);
or U14621 (N_14621,N_13090,N_13032);
nand U14622 (N_14622,N_13422,N_13318);
and U14623 (N_14623,N_12044,N_13513);
and U14624 (N_14624,N_12146,N_12105);
or U14625 (N_14625,N_12576,N_12394);
nor U14626 (N_14626,N_13116,N_13228);
nand U14627 (N_14627,N_13048,N_12650);
nor U14628 (N_14628,N_13184,N_13870);
xnor U14629 (N_14629,N_12218,N_13718);
and U14630 (N_14630,N_12514,N_13231);
xor U14631 (N_14631,N_12011,N_12993);
xnor U14632 (N_14632,N_12633,N_12773);
and U14633 (N_14633,N_12001,N_12745);
nand U14634 (N_14634,N_13806,N_13719);
or U14635 (N_14635,N_12992,N_12424);
nor U14636 (N_14636,N_13592,N_12124);
nand U14637 (N_14637,N_12654,N_12903);
xor U14638 (N_14638,N_12375,N_12515);
nor U14639 (N_14639,N_12125,N_13895);
xnor U14640 (N_14640,N_12045,N_12460);
and U14641 (N_14641,N_12127,N_13772);
nand U14642 (N_14642,N_13195,N_13448);
nand U14643 (N_14643,N_13525,N_13565);
nor U14644 (N_14644,N_12702,N_13511);
nor U14645 (N_14645,N_12562,N_13483);
nand U14646 (N_14646,N_13803,N_13209);
nor U14647 (N_14647,N_13198,N_13373);
nand U14648 (N_14648,N_12727,N_13356);
xnor U14649 (N_14649,N_12033,N_12320);
nor U14650 (N_14650,N_13442,N_13598);
or U14651 (N_14651,N_13515,N_13307);
and U14652 (N_14652,N_12159,N_13672);
xnor U14653 (N_14653,N_12848,N_12731);
xnor U14654 (N_14654,N_13729,N_12481);
and U14655 (N_14655,N_12366,N_12345);
xnor U14656 (N_14656,N_13728,N_13054);
nand U14657 (N_14657,N_12037,N_13357);
xnor U14658 (N_14658,N_12107,N_13435);
or U14659 (N_14659,N_12991,N_12389);
xnor U14660 (N_14660,N_12797,N_12506);
xnor U14661 (N_14661,N_12110,N_13969);
nand U14662 (N_14662,N_13767,N_13879);
and U14663 (N_14663,N_13555,N_13754);
and U14664 (N_14664,N_12397,N_12775);
and U14665 (N_14665,N_12572,N_13907);
and U14666 (N_14666,N_12223,N_12211);
or U14667 (N_14667,N_12499,N_12786);
and U14668 (N_14668,N_12046,N_12018);
nor U14669 (N_14669,N_13488,N_13413);
xnor U14670 (N_14670,N_13634,N_12827);
or U14671 (N_14671,N_13275,N_12536);
nand U14672 (N_14672,N_13858,N_13497);
nor U14673 (N_14673,N_13716,N_12043);
nand U14674 (N_14674,N_13139,N_12958);
nor U14675 (N_14675,N_12128,N_12292);
nand U14676 (N_14676,N_12297,N_13176);
nand U14677 (N_14677,N_12457,N_12404);
xor U14678 (N_14678,N_12227,N_13451);
and U14679 (N_14679,N_13210,N_13789);
xor U14680 (N_14680,N_13528,N_12139);
nor U14681 (N_14681,N_12183,N_13454);
and U14682 (N_14682,N_13349,N_13110);
or U14683 (N_14683,N_13256,N_12588);
or U14684 (N_14684,N_12244,N_12689);
nor U14685 (N_14685,N_13112,N_12393);
nor U14686 (N_14686,N_13324,N_13093);
and U14687 (N_14687,N_12929,N_13864);
and U14688 (N_14688,N_13502,N_12063);
nand U14689 (N_14689,N_12799,N_13156);
or U14690 (N_14690,N_13338,N_12653);
nor U14691 (N_14691,N_12606,N_13771);
nand U14692 (N_14692,N_12936,N_13945);
or U14693 (N_14693,N_12195,N_12655);
or U14694 (N_14694,N_12521,N_12612);
xor U14695 (N_14695,N_12206,N_12425);
nand U14696 (N_14696,N_12526,N_12316);
and U14697 (N_14697,N_12604,N_13624);
or U14698 (N_14698,N_13914,N_12120);
or U14699 (N_14699,N_13472,N_12459);
or U14700 (N_14700,N_12512,N_12941);
and U14701 (N_14701,N_12053,N_12487);
and U14702 (N_14702,N_13291,N_12822);
and U14703 (N_14703,N_12785,N_13269);
nor U14704 (N_14704,N_12529,N_12753);
xnor U14705 (N_14705,N_12746,N_12659);
xnor U14706 (N_14706,N_13576,N_12878);
xnor U14707 (N_14707,N_12511,N_13206);
xnor U14708 (N_14708,N_12641,N_12291);
nor U14709 (N_14709,N_13485,N_13397);
or U14710 (N_14710,N_12834,N_13671);
nor U14711 (N_14711,N_12092,N_13650);
or U14712 (N_14712,N_12167,N_12880);
and U14713 (N_14713,N_13509,N_12498);
nand U14714 (N_14714,N_12276,N_13364);
and U14715 (N_14715,N_12360,N_12150);
xnor U14716 (N_14716,N_12203,N_12247);
nor U14717 (N_14717,N_13143,N_12682);
nand U14718 (N_14718,N_12701,N_13997);
and U14719 (N_14719,N_12259,N_13063);
xnor U14720 (N_14720,N_12288,N_13820);
and U14721 (N_14721,N_13613,N_12714);
nor U14722 (N_14722,N_12871,N_12478);
nor U14723 (N_14723,N_12555,N_13013);
and U14724 (N_14724,N_12141,N_12877);
or U14725 (N_14725,N_12658,N_13127);
xor U14726 (N_14726,N_12335,N_12193);
nand U14727 (N_14727,N_12471,N_13038);
nand U14728 (N_14728,N_12314,N_13499);
nand U14729 (N_14729,N_13703,N_13980);
nor U14730 (N_14730,N_12189,N_12239);
or U14731 (N_14731,N_13916,N_13877);
or U14732 (N_14732,N_13041,N_12299);
nand U14733 (N_14733,N_13202,N_13878);
nor U14734 (N_14734,N_12103,N_12461);
nand U14735 (N_14735,N_13440,N_12061);
or U14736 (N_14736,N_13168,N_12435);
nor U14737 (N_14737,N_13494,N_13419);
and U14738 (N_14738,N_13518,N_13007);
xor U14739 (N_14739,N_13996,N_12380);
or U14740 (N_14740,N_12851,N_13574);
or U14741 (N_14741,N_13711,N_12523);
xor U14742 (N_14742,N_13298,N_13516);
or U14743 (N_14743,N_13594,N_12265);
nand U14744 (N_14744,N_13761,N_12776);
xor U14745 (N_14745,N_13088,N_12632);
nand U14746 (N_14746,N_13033,N_12946);
and U14747 (N_14747,N_13649,N_12722);
nor U14748 (N_14748,N_13691,N_13092);
nor U14749 (N_14749,N_13736,N_13533);
or U14750 (N_14750,N_12453,N_12339);
xor U14751 (N_14751,N_12458,N_12421);
nor U14752 (N_14752,N_12581,N_12864);
xor U14753 (N_14753,N_12182,N_13311);
nor U14754 (N_14754,N_12620,N_13614);
and U14755 (N_14755,N_12525,N_12644);
nor U14756 (N_14756,N_13329,N_13212);
xor U14757 (N_14757,N_13008,N_13459);
nor U14758 (N_14758,N_12405,N_12628);
xnor U14759 (N_14759,N_13268,N_12820);
or U14760 (N_14760,N_13262,N_13734);
nor U14761 (N_14761,N_13871,N_12517);
and U14762 (N_14762,N_12665,N_13123);
nor U14763 (N_14763,N_12850,N_13812);
and U14764 (N_14764,N_13312,N_12310);
and U14765 (N_14765,N_12869,N_12558);
nand U14766 (N_14766,N_13527,N_13476);
nor U14767 (N_14767,N_13490,N_13827);
xnor U14768 (N_14768,N_13505,N_12796);
nand U14769 (N_14769,N_13392,N_13052);
nand U14770 (N_14770,N_13800,N_13765);
or U14771 (N_14771,N_13930,N_13857);
nor U14772 (N_14772,N_12968,N_13332);
nor U14773 (N_14773,N_12766,N_12533);
and U14774 (N_14774,N_13203,N_13045);
xor U14775 (N_14775,N_12075,N_13917);
xnor U14776 (N_14776,N_13217,N_12340);
xnor U14777 (N_14777,N_13122,N_12431);
xor U14778 (N_14778,N_13970,N_13946);
nand U14779 (N_14779,N_13713,N_13321);
or U14780 (N_14780,N_13082,N_12420);
and U14781 (N_14781,N_13875,N_13544);
and U14782 (N_14782,N_12041,N_13661);
and U14783 (N_14783,N_13345,N_12267);
nor U14784 (N_14784,N_12242,N_12909);
or U14785 (N_14785,N_12617,N_13276);
and U14786 (N_14786,N_13764,N_13901);
or U14787 (N_14787,N_12073,N_13836);
nor U14788 (N_14788,N_13638,N_12317);
or U14789 (N_14789,N_12953,N_12747);
or U14790 (N_14790,N_12281,N_13702);
nor U14791 (N_14791,N_13626,N_13952);
nand U14792 (N_14792,N_12782,N_13408);
nand U14793 (N_14793,N_12681,N_13710);
xnor U14794 (N_14794,N_12955,N_12256);
xor U14795 (N_14795,N_12081,N_13665);
and U14796 (N_14796,N_13365,N_13213);
or U14797 (N_14797,N_12401,N_13056);
and U14798 (N_14798,N_13174,N_13166);
nor U14799 (N_14799,N_12508,N_13667);
and U14800 (N_14800,N_13316,N_13787);
and U14801 (N_14801,N_13400,N_12123);
xnor U14802 (N_14802,N_13233,N_13303);
or U14803 (N_14803,N_13410,N_12076);
or U14804 (N_14804,N_13867,N_13696);
and U14805 (N_14805,N_13735,N_12152);
and U14806 (N_14806,N_12983,N_13254);
nand U14807 (N_14807,N_13839,N_13730);
or U14808 (N_14808,N_12765,N_13636);
nor U14809 (N_14809,N_12034,N_12571);
xor U14810 (N_14810,N_13971,N_12861);
and U14811 (N_14811,N_13608,N_13283);
nand U14812 (N_14812,N_13117,N_13625);
and U14813 (N_14813,N_13471,N_13687);
xnor U14814 (N_14814,N_13255,N_13371);
xnor U14815 (N_14815,N_12336,N_12897);
nor U14816 (N_14816,N_12901,N_12200);
and U14817 (N_14817,N_12440,N_12382);
nand U14818 (N_14818,N_13887,N_13693);
nand U14819 (N_14819,N_12408,N_12427);
nand U14820 (N_14820,N_12452,N_12610);
and U14821 (N_14821,N_12780,N_13724);
or U14822 (N_14822,N_12462,N_12503);
or U14823 (N_14823,N_12055,N_12240);
nor U14824 (N_14824,N_12000,N_13683);
xor U14825 (N_14825,N_12798,N_13851);
or U14826 (N_14826,N_12145,N_13940);
nand U14827 (N_14827,N_13532,N_12707);
nand U14828 (N_14828,N_13991,N_12577);
and U14829 (N_14829,N_12844,N_12050);
or U14830 (N_14830,N_13024,N_12962);
nor U14831 (N_14831,N_13783,N_13336);
or U14832 (N_14832,N_13596,N_12049);
and U14833 (N_14833,N_13651,N_13169);
or U14834 (N_14834,N_12964,N_13192);
and U14835 (N_14835,N_12038,N_13044);
or U14836 (N_14836,N_12181,N_12032);
nor U14837 (N_14837,N_13894,N_13017);
xnor U14838 (N_14838,N_13615,N_12156);
nand U14839 (N_14839,N_12551,N_12439);
or U14840 (N_14840,N_13759,N_12302);
nor U14841 (N_14841,N_13042,N_13136);
xor U14842 (N_14842,N_12635,N_12101);
nand U14843 (N_14843,N_13689,N_12587);
and U14844 (N_14844,N_12108,N_12596);
xnor U14845 (N_14845,N_12710,N_12945);
nand U14846 (N_14846,N_13493,N_13125);
and U14847 (N_14847,N_12135,N_12524);
and U14848 (N_14848,N_12456,N_12601);
and U14849 (N_14849,N_13985,N_13983);
xnor U14850 (N_14850,N_12934,N_13204);
xor U14851 (N_14851,N_13855,N_13452);
or U14852 (N_14852,N_13816,N_13461);
nor U14853 (N_14853,N_12625,N_13998);
or U14854 (N_14854,N_12283,N_13673);
nor U14855 (N_14855,N_13732,N_12982);
nor U14856 (N_14856,N_12771,N_12398);
nor U14857 (N_14857,N_12977,N_13862);
nand U14858 (N_14858,N_13072,N_13774);
nor U14859 (N_14859,N_13853,N_13229);
and U14860 (N_14860,N_12332,N_12575);
nor U14861 (N_14861,N_13540,N_12812);
and U14862 (N_14862,N_12591,N_12939);
and U14863 (N_14863,N_13698,N_12837);
and U14864 (N_14864,N_12724,N_13628);
or U14865 (N_14865,N_12137,N_13286);
nand U14866 (N_14866,N_13478,N_13519);
nor U14867 (N_14867,N_12813,N_12391);
nor U14868 (N_14868,N_12153,N_12885);
nand U14869 (N_14869,N_12892,N_12522);
nand U14870 (N_14870,N_13637,N_12388);
or U14871 (N_14871,N_13884,N_12923);
and U14872 (N_14872,N_13366,N_13104);
xnor U14873 (N_14873,N_13758,N_13155);
nand U14874 (N_14874,N_13118,N_12477);
xnor U14875 (N_14875,N_13465,N_13133);
and U14876 (N_14876,N_13333,N_13474);
nor U14877 (N_14877,N_12669,N_12774);
nand U14878 (N_14878,N_12670,N_13211);
or U14879 (N_14879,N_12739,N_13768);
nor U14880 (N_14880,N_13145,N_13535);
xnor U14881 (N_14881,N_12794,N_12373);
nor U14882 (N_14882,N_13921,N_13407);
nor U14883 (N_14883,N_13259,N_12704);
xor U14884 (N_14884,N_12543,N_13706);
nand U14885 (N_14885,N_12636,N_12069);
or U14886 (N_14886,N_12353,N_13943);
nand U14887 (N_14887,N_13990,N_12093);
xor U14888 (N_14888,N_12803,N_13075);
xor U14889 (N_14889,N_12009,N_13375);
nand U14890 (N_14890,N_12238,N_12679);
or U14891 (N_14891,N_12987,N_13507);
xnor U14892 (N_14892,N_12629,N_13188);
nor U14893 (N_14893,N_12973,N_12913);
and U14894 (N_14894,N_13339,N_12437);
or U14895 (N_14895,N_12175,N_12564);
nand U14896 (N_14896,N_13260,N_12047);
and U14897 (N_14897,N_13379,N_12502);
nand U14898 (N_14898,N_13305,N_12100);
xnor U14899 (N_14899,N_12924,N_12433);
nand U14900 (N_14900,N_12060,N_12563);
or U14901 (N_14901,N_13430,N_13501);
or U14902 (N_14902,N_13709,N_13692);
or U14903 (N_14903,N_13699,N_13098);
and U14904 (N_14904,N_13792,N_12311);
nand U14905 (N_14905,N_12177,N_13399);
or U14906 (N_14906,N_12586,N_12374);
or U14907 (N_14907,N_13743,N_13954);
xnor U14908 (N_14908,N_13814,N_13994);
or U14909 (N_14909,N_12493,N_13618);
nand U14910 (N_14910,N_13953,N_13457);
nand U14911 (N_14911,N_13966,N_13245);
xor U14912 (N_14912,N_12142,N_13834);
and U14913 (N_14913,N_13450,N_13824);
xor U14914 (N_14914,N_13523,N_12967);
and U14915 (N_14915,N_12910,N_13899);
nand U14916 (N_14916,N_12855,N_12186);
nand U14917 (N_14917,N_13588,N_12912);
and U14918 (N_14918,N_12006,N_13214);
nand U14919 (N_14919,N_12155,N_13016);
nor U14920 (N_14920,N_13503,N_12449);
nor U14921 (N_14921,N_13541,N_12580);
and U14922 (N_14922,N_13915,N_13986);
xor U14923 (N_14923,N_13644,N_13904);
xnor U14924 (N_14924,N_13086,N_12309);
and U14925 (N_14925,N_12328,N_12981);
xnor U14926 (N_14926,N_12286,N_13537);
nand U14927 (N_14927,N_12842,N_13645);
xor U14928 (N_14928,N_12740,N_12614);
and U14929 (N_14929,N_13825,N_12306);
or U14930 (N_14930,N_13563,N_12413);
nor U14931 (N_14931,N_12860,N_13762);
nor U14932 (N_14932,N_13579,N_13157);
nor U14933 (N_14933,N_12251,N_12149);
nor U14934 (N_14934,N_13844,N_12365);
or U14935 (N_14935,N_12677,N_13840);
nor U14936 (N_14936,N_13015,N_12639);
xor U14937 (N_14937,N_12959,N_13121);
and U14938 (N_14938,N_12783,N_13546);
or U14939 (N_14939,N_12164,N_12355);
nand U14940 (N_14940,N_13727,N_13815);
nand U14941 (N_14941,N_13607,N_12348);
nand U14942 (N_14942,N_12147,N_13653);
or U14943 (N_14943,N_13280,N_12030);
and U14944 (N_14944,N_12876,N_13393);
nor U14945 (N_14945,N_12708,N_12436);
or U14946 (N_14946,N_13248,N_12886);
nor U14947 (N_14947,N_13183,N_13821);
nor U14948 (N_14948,N_13141,N_12403);
and U14949 (N_14949,N_12479,N_12889);
and U14950 (N_14950,N_13959,N_12578);
or U14951 (N_14951,N_13569,N_12535);
nand U14952 (N_14952,N_13601,N_12737);
and U14953 (N_14953,N_13394,N_12102);
nor U14954 (N_14954,N_13668,N_13796);
nand U14955 (N_14955,N_13475,N_13353);
or U14956 (N_14956,N_12346,N_12758);
xnor U14957 (N_14957,N_13029,N_13560);
and U14958 (N_14958,N_13690,N_12402);
xnor U14959 (N_14959,N_13390,N_12921);
and U14960 (N_14960,N_13040,N_12416);
xnor U14961 (N_14961,N_13480,N_13520);
nand U14962 (N_14962,N_12852,N_12450);
nor U14963 (N_14963,N_12356,N_13883);
xnor U14964 (N_14964,N_12442,N_12262);
nand U14965 (N_14965,N_13627,N_12007);
or U14966 (N_14966,N_12187,N_12352);
nor U14967 (N_14967,N_12321,N_12274);
nor U14968 (N_14968,N_12068,N_13828);
nand U14969 (N_14969,N_12184,N_12907);
or U14970 (N_14970,N_12607,N_13386);
nand U14971 (N_14971,N_13100,N_12085);
or U14972 (N_14972,N_13273,N_13837);
nor U14973 (N_14973,N_13989,N_12609);
and U14974 (N_14974,N_13521,N_13258);
nor U14975 (N_14975,N_12157,N_13049);
and U14976 (N_14976,N_13343,N_12816);
or U14977 (N_14977,N_12637,N_12094);
and U14978 (N_14978,N_13760,N_13058);
or U14979 (N_14979,N_12688,N_12832);
nor U14980 (N_14980,N_12699,N_12919);
nor U14981 (N_14981,N_13124,N_12057);
xor U14982 (N_14982,N_13808,N_13733);
nor U14983 (N_14983,N_12019,N_12342);
nor U14984 (N_14984,N_13819,N_12338);
nor U14985 (N_14985,N_12214,N_13972);
and U14986 (N_14986,N_13881,N_12015);
nand U14987 (N_14987,N_12943,N_12908);
or U14988 (N_14988,N_13149,N_12188);
or U14989 (N_14989,N_13852,N_12219);
nor U14990 (N_14990,N_12190,N_13950);
and U14991 (N_14991,N_12862,N_12583);
nand U14992 (N_14992,N_13030,N_13876);
and U14993 (N_14993,N_12942,N_13766);
and U14994 (N_14994,N_12280,N_13205);
or U14995 (N_14995,N_12804,N_13061);
nand U14996 (N_14996,N_12956,N_12161);
xnor U14997 (N_14997,N_12319,N_12978);
or U14998 (N_14998,N_12303,N_13065);
xnor U14999 (N_14999,N_12557,N_13062);
xnor U15000 (N_15000,N_12614,N_13605);
and U15001 (N_15001,N_12728,N_13446);
nand U15002 (N_15002,N_12653,N_13623);
or U15003 (N_15003,N_13707,N_12890);
or U15004 (N_15004,N_12498,N_13490);
nand U15005 (N_15005,N_12787,N_13751);
nor U15006 (N_15006,N_12825,N_13628);
and U15007 (N_15007,N_13007,N_12685);
nand U15008 (N_15008,N_12848,N_12262);
xor U15009 (N_15009,N_12605,N_13106);
nand U15010 (N_15010,N_12513,N_13190);
nor U15011 (N_15011,N_13409,N_12529);
xor U15012 (N_15012,N_13783,N_13769);
or U15013 (N_15013,N_13844,N_12125);
nand U15014 (N_15014,N_13901,N_13223);
nand U15015 (N_15015,N_13474,N_12954);
and U15016 (N_15016,N_13215,N_13804);
xor U15017 (N_15017,N_13982,N_12825);
xnor U15018 (N_15018,N_13832,N_13284);
nor U15019 (N_15019,N_12930,N_12889);
and U15020 (N_15020,N_13446,N_12799);
nand U15021 (N_15021,N_13968,N_12067);
or U15022 (N_15022,N_12378,N_13248);
or U15023 (N_15023,N_13007,N_12880);
or U15024 (N_15024,N_13623,N_12897);
nor U15025 (N_15025,N_12355,N_13847);
xor U15026 (N_15026,N_12561,N_12172);
or U15027 (N_15027,N_13544,N_13183);
nor U15028 (N_15028,N_12163,N_12265);
nand U15029 (N_15029,N_13924,N_12162);
nor U15030 (N_15030,N_12954,N_12704);
nor U15031 (N_15031,N_13959,N_13789);
xnor U15032 (N_15032,N_13368,N_12327);
and U15033 (N_15033,N_13968,N_13310);
nor U15034 (N_15034,N_13911,N_12522);
or U15035 (N_15035,N_13217,N_12011);
nor U15036 (N_15036,N_12923,N_12534);
nor U15037 (N_15037,N_13439,N_12422);
nand U15038 (N_15038,N_13943,N_13309);
nand U15039 (N_15039,N_13401,N_12346);
or U15040 (N_15040,N_13602,N_13296);
nand U15041 (N_15041,N_12231,N_12760);
or U15042 (N_15042,N_13672,N_13791);
or U15043 (N_15043,N_13944,N_13365);
or U15044 (N_15044,N_12049,N_12894);
nand U15045 (N_15045,N_12998,N_12820);
or U15046 (N_15046,N_12188,N_13322);
nand U15047 (N_15047,N_13965,N_13414);
xnor U15048 (N_15048,N_13008,N_12915);
and U15049 (N_15049,N_12485,N_13981);
xnor U15050 (N_15050,N_13867,N_13853);
or U15051 (N_15051,N_12603,N_12895);
xnor U15052 (N_15052,N_13058,N_12511);
and U15053 (N_15053,N_12347,N_13436);
nand U15054 (N_15054,N_12801,N_13372);
and U15055 (N_15055,N_13912,N_13267);
and U15056 (N_15056,N_13056,N_12369);
nor U15057 (N_15057,N_13261,N_13189);
nor U15058 (N_15058,N_12486,N_13028);
xnor U15059 (N_15059,N_13511,N_13386);
nand U15060 (N_15060,N_12709,N_13706);
and U15061 (N_15061,N_12936,N_13401);
xor U15062 (N_15062,N_13168,N_13021);
xnor U15063 (N_15063,N_12484,N_12078);
nand U15064 (N_15064,N_12215,N_12148);
xor U15065 (N_15065,N_12076,N_13087);
nor U15066 (N_15066,N_12342,N_13484);
and U15067 (N_15067,N_12873,N_12000);
or U15068 (N_15068,N_13742,N_12726);
nand U15069 (N_15069,N_12827,N_12921);
xnor U15070 (N_15070,N_13874,N_13279);
xnor U15071 (N_15071,N_13523,N_13527);
or U15072 (N_15072,N_13628,N_13933);
xor U15073 (N_15073,N_12301,N_12220);
xnor U15074 (N_15074,N_12518,N_12447);
nor U15075 (N_15075,N_13375,N_13191);
nor U15076 (N_15076,N_12516,N_12577);
xnor U15077 (N_15077,N_13757,N_13314);
nor U15078 (N_15078,N_13102,N_13513);
and U15079 (N_15079,N_12180,N_13231);
nand U15080 (N_15080,N_12473,N_12125);
and U15081 (N_15081,N_12148,N_13300);
or U15082 (N_15082,N_13231,N_12213);
nand U15083 (N_15083,N_13505,N_12656);
nand U15084 (N_15084,N_13789,N_13014);
and U15085 (N_15085,N_12883,N_12107);
and U15086 (N_15086,N_13346,N_13676);
nand U15087 (N_15087,N_12612,N_13516);
nand U15088 (N_15088,N_12246,N_12048);
nor U15089 (N_15089,N_13227,N_12164);
nand U15090 (N_15090,N_13639,N_12660);
xor U15091 (N_15091,N_12967,N_12621);
or U15092 (N_15092,N_13696,N_13448);
and U15093 (N_15093,N_12289,N_12881);
or U15094 (N_15094,N_12065,N_13392);
and U15095 (N_15095,N_13074,N_12031);
nand U15096 (N_15096,N_13356,N_12931);
or U15097 (N_15097,N_13405,N_13367);
or U15098 (N_15098,N_12141,N_13480);
nor U15099 (N_15099,N_12020,N_12112);
or U15100 (N_15100,N_13516,N_12233);
xnor U15101 (N_15101,N_13529,N_12145);
nand U15102 (N_15102,N_13987,N_13902);
nor U15103 (N_15103,N_12149,N_13886);
or U15104 (N_15104,N_12506,N_13485);
or U15105 (N_15105,N_12989,N_13330);
nor U15106 (N_15106,N_12878,N_13804);
nor U15107 (N_15107,N_13633,N_13367);
xor U15108 (N_15108,N_13211,N_13884);
or U15109 (N_15109,N_12645,N_12945);
or U15110 (N_15110,N_13495,N_12720);
nand U15111 (N_15111,N_13071,N_13956);
xor U15112 (N_15112,N_12250,N_12332);
nand U15113 (N_15113,N_13547,N_12706);
nand U15114 (N_15114,N_12656,N_12736);
nand U15115 (N_15115,N_13152,N_13234);
nand U15116 (N_15116,N_12609,N_13182);
nor U15117 (N_15117,N_12240,N_13869);
nand U15118 (N_15118,N_13842,N_12278);
and U15119 (N_15119,N_13655,N_13052);
nor U15120 (N_15120,N_12380,N_13593);
nor U15121 (N_15121,N_12253,N_12546);
nand U15122 (N_15122,N_13809,N_12313);
nor U15123 (N_15123,N_12114,N_13102);
nand U15124 (N_15124,N_12174,N_13607);
and U15125 (N_15125,N_13898,N_13004);
xor U15126 (N_15126,N_12198,N_12582);
xnor U15127 (N_15127,N_12309,N_13220);
or U15128 (N_15128,N_12691,N_12044);
and U15129 (N_15129,N_12339,N_13318);
or U15130 (N_15130,N_13922,N_13001);
nand U15131 (N_15131,N_13288,N_12513);
or U15132 (N_15132,N_13109,N_13952);
and U15133 (N_15133,N_13370,N_13857);
nand U15134 (N_15134,N_12631,N_13161);
or U15135 (N_15135,N_12273,N_12560);
or U15136 (N_15136,N_13155,N_12856);
xor U15137 (N_15137,N_13538,N_12440);
nand U15138 (N_15138,N_12467,N_13947);
and U15139 (N_15139,N_12907,N_13427);
and U15140 (N_15140,N_12649,N_13198);
nand U15141 (N_15141,N_12035,N_12263);
and U15142 (N_15142,N_12172,N_13553);
or U15143 (N_15143,N_13144,N_12993);
and U15144 (N_15144,N_13942,N_12823);
nand U15145 (N_15145,N_12638,N_13173);
or U15146 (N_15146,N_13837,N_12370);
nor U15147 (N_15147,N_13071,N_12057);
nor U15148 (N_15148,N_13008,N_12134);
and U15149 (N_15149,N_12841,N_12838);
or U15150 (N_15150,N_12076,N_13050);
and U15151 (N_15151,N_13169,N_13271);
xnor U15152 (N_15152,N_12352,N_13761);
nor U15153 (N_15153,N_12469,N_13600);
nand U15154 (N_15154,N_12243,N_13776);
nor U15155 (N_15155,N_12561,N_12612);
nor U15156 (N_15156,N_13852,N_12002);
or U15157 (N_15157,N_13665,N_12299);
or U15158 (N_15158,N_13726,N_13783);
xor U15159 (N_15159,N_12320,N_12020);
nor U15160 (N_15160,N_12677,N_12220);
xor U15161 (N_15161,N_13112,N_13864);
nand U15162 (N_15162,N_12960,N_12929);
and U15163 (N_15163,N_13761,N_13858);
nor U15164 (N_15164,N_12553,N_13721);
xor U15165 (N_15165,N_13006,N_12513);
nor U15166 (N_15166,N_13997,N_12305);
nand U15167 (N_15167,N_12756,N_13869);
or U15168 (N_15168,N_12315,N_13539);
nand U15169 (N_15169,N_13007,N_13344);
nand U15170 (N_15170,N_12335,N_12967);
and U15171 (N_15171,N_13545,N_12932);
or U15172 (N_15172,N_12732,N_12434);
or U15173 (N_15173,N_12030,N_12359);
nand U15174 (N_15174,N_13493,N_12398);
and U15175 (N_15175,N_12793,N_12621);
and U15176 (N_15176,N_12127,N_12940);
or U15177 (N_15177,N_12843,N_13345);
xnor U15178 (N_15178,N_13190,N_12729);
nand U15179 (N_15179,N_12347,N_13662);
nor U15180 (N_15180,N_12292,N_13260);
nand U15181 (N_15181,N_12832,N_13240);
or U15182 (N_15182,N_12937,N_13743);
nand U15183 (N_15183,N_13836,N_12907);
and U15184 (N_15184,N_12552,N_12423);
nor U15185 (N_15185,N_12229,N_12588);
xor U15186 (N_15186,N_12711,N_13602);
and U15187 (N_15187,N_13472,N_12635);
and U15188 (N_15188,N_12014,N_12530);
nor U15189 (N_15189,N_13277,N_12070);
nand U15190 (N_15190,N_12730,N_13049);
xnor U15191 (N_15191,N_12994,N_12527);
or U15192 (N_15192,N_12952,N_13080);
or U15193 (N_15193,N_13662,N_12192);
nand U15194 (N_15194,N_12003,N_13088);
or U15195 (N_15195,N_13652,N_13437);
nor U15196 (N_15196,N_13234,N_12438);
or U15197 (N_15197,N_13334,N_12249);
xnor U15198 (N_15198,N_12290,N_12098);
nand U15199 (N_15199,N_12101,N_12311);
nand U15200 (N_15200,N_12634,N_13241);
xnor U15201 (N_15201,N_13462,N_13234);
xnor U15202 (N_15202,N_12494,N_12787);
or U15203 (N_15203,N_12783,N_12890);
or U15204 (N_15204,N_13539,N_12022);
or U15205 (N_15205,N_13525,N_13965);
nor U15206 (N_15206,N_12540,N_13167);
or U15207 (N_15207,N_12358,N_12893);
or U15208 (N_15208,N_13454,N_13173);
and U15209 (N_15209,N_12855,N_12798);
or U15210 (N_15210,N_13203,N_12717);
xnor U15211 (N_15211,N_13091,N_13979);
nor U15212 (N_15212,N_12550,N_12818);
nand U15213 (N_15213,N_13818,N_13113);
xnor U15214 (N_15214,N_12083,N_12830);
or U15215 (N_15215,N_13061,N_13484);
or U15216 (N_15216,N_12081,N_13635);
xnor U15217 (N_15217,N_13206,N_12531);
or U15218 (N_15218,N_12391,N_12494);
xnor U15219 (N_15219,N_12275,N_12740);
and U15220 (N_15220,N_12235,N_13064);
xor U15221 (N_15221,N_12515,N_13796);
or U15222 (N_15222,N_12084,N_12789);
or U15223 (N_15223,N_13680,N_12517);
or U15224 (N_15224,N_13131,N_12746);
nand U15225 (N_15225,N_13757,N_12398);
or U15226 (N_15226,N_12654,N_13691);
or U15227 (N_15227,N_13840,N_12758);
and U15228 (N_15228,N_12169,N_12318);
or U15229 (N_15229,N_12269,N_13801);
nand U15230 (N_15230,N_12166,N_13282);
or U15231 (N_15231,N_12893,N_13825);
or U15232 (N_15232,N_13341,N_13065);
or U15233 (N_15233,N_13391,N_12431);
nor U15234 (N_15234,N_12630,N_13167);
nor U15235 (N_15235,N_13486,N_13727);
nand U15236 (N_15236,N_13110,N_12498);
nor U15237 (N_15237,N_13772,N_12321);
nand U15238 (N_15238,N_12716,N_13274);
nand U15239 (N_15239,N_13165,N_13100);
and U15240 (N_15240,N_12658,N_12238);
and U15241 (N_15241,N_13468,N_13443);
nor U15242 (N_15242,N_13460,N_13128);
nor U15243 (N_15243,N_12596,N_13669);
and U15244 (N_15244,N_13458,N_13091);
xnor U15245 (N_15245,N_13669,N_12038);
xnor U15246 (N_15246,N_13719,N_13392);
nand U15247 (N_15247,N_13986,N_13702);
nor U15248 (N_15248,N_12187,N_12449);
or U15249 (N_15249,N_12577,N_13176);
nor U15250 (N_15250,N_13230,N_13102);
xor U15251 (N_15251,N_12726,N_12822);
nor U15252 (N_15252,N_12410,N_13771);
xnor U15253 (N_15253,N_12761,N_13252);
nand U15254 (N_15254,N_13608,N_13634);
or U15255 (N_15255,N_12652,N_13294);
xnor U15256 (N_15256,N_12603,N_12599);
nand U15257 (N_15257,N_12366,N_13373);
nand U15258 (N_15258,N_13805,N_12255);
or U15259 (N_15259,N_12497,N_13248);
xor U15260 (N_15260,N_12104,N_13996);
nor U15261 (N_15261,N_12086,N_13066);
or U15262 (N_15262,N_13693,N_13088);
xnor U15263 (N_15263,N_12192,N_12190);
nand U15264 (N_15264,N_12406,N_13438);
nand U15265 (N_15265,N_13925,N_13579);
xnor U15266 (N_15266,N_13462,N_13493);
or U15267 (N_15267,N_12567,N_12491);
or U15268 (N_15268,N_12887,N_13120);
and U15269 (N_15269,N_12165,N_12206);
or U15270 (N_15270,N_13626,N_13003);
xor U15271 (N_15271,N_12751,N_13349);
nand U15272 (N_15272,N_13964,N_13617);
nor U15273 (N_15273,N_13803,N_12738);
nor U15274 (N_15274,N_13421,N_13772);
nand U15275 (N_15275,N_12671,N_13272);
or U15276 (N_15276,N_13463,N_13959);
xnor U15277 (N_15277,N_12042,N_12130);
nand U15278 (N_15278,N_13948,N_13525);
nand U15279 (N_15279,N_13454,N_12965);
nand U15280 (N_15280,N_12714,N_12512);
nand U15281 (N_15281,N_12818,N_12507);
or U15282 (N_15282,N_13698,N_12880);
nand U15283 (N_15283,N_13749,N_12281);
nand U15284 (N_15284,N_12137,N_12125);
or U15285 (N_15285,N_12007,N_12637);
and U15286 (N_15286,N_13066,N_12168);
nor U15287 (N_15287,N_13313,N_12351);
and U15288 (N_15288,N_13017,N_13528);
nor U15289 (N_15289,N_12490,N_13554);
xnor U15290 (N_15290,N_12093,N_12150);
nand U15291 (N_15291,N_12701,N_12988);
xor U15292 (N_15292,N_12779,N_12686);
nor U15293 (N_15293,N_13689,N_13275);
or U15294 (N_15294,N_12987,N_12237);
nand U15295 (N_15295,N_13543,N_13587);
nand U15296 (N_15296,N_13596,N_13246);
nand U15297 (N_15297,N_12327,N_13835);
nand U15298 (N_15298,N_12610,N_12368);
xnor U15299 (N_15299,N_12682,N_13924);
or U15300 (N_15300,N_12771,N_13526);
or U15301 (N_15301,N_12739,N_12655);
and U15302 (N_15302,N_13703,N_12027);
nor U15303 (N_15303,N_13663,N_12266);
nand U15304 (N_15304,N_13055,N_12278);
xor U15305 (N_15305,N_12654,N_12593);
nand U15306 (N_15306,N_12871,N_12067);
nor U15307 (N_15307,N_13754,N_13072);
nor U15308 (N_15308,N_13183,N_12475);
xnor U15309 (N_15309,N_13630,N_12855);
xnor U15310 (N_15310,N_12347,N_12063);
and U15311 (N_15311,N_12884,N_13058);
nor U15312 (N_15312,N_13684,N_13611);
nand U15313 (N_15313,N_12041,N_12396);
nand U15314 (N_15314,N_12200,N_13689);
nor U15315 (N_15315,N_12790,N_13833);
nor U15316 (N_15316,N_12475,N_13459);
nand U15317 (N_15317,N_13935,N_13675);
xnor U15318 (N_15318,N_13306,N_13214);
xnor U15319 (N_15319,N_12587,N_13220);
nand U15320 (N_15320,N_13234,N_12982);
or U15321 (N_15321,N_13815,N_12988);
or U15322 (N_15322,N_13499,N_13403);
nand U15323 (N_15323,N_12302,N_12163);
and U15324 (N_15324,N_13172,N_12954);
nand U15325 (N_15325,N_13543,N_12410);
nor U15326 (N_15326,N_12265,N_12903);
nor U15327 (N_15327,N_13711,N_12942);
xor U15328 (N_15328,N_13100,N_13356);
or U15329 (N_15329,N_13230,N_13831);
or U15330 (N_15330,N_12105,N_12371);
or U15331 (N_15331,N_12854,N_12419);
or U15332 (N_15332,N_13972,N_12958);
and U15333 (N_15333,N_12955,N_12092);
xnor U15334 (N_15334,N_13284,N_12727);
nand U15335 (N_15335,N_13828,N_12217);
or U15336 (N_15336,N_12698,N_13297);
xnor U15337 (N_15337,N_13566,N_12485);
nor U15338 (N_15338,N_13757,N_12435);
and U15339 (N_15339,N_12396,N_13948);
nor U15340 (N_15340,N_12594,N_12791);
or U15341 (N_15341,N_12147,N_13815);
and U15342 (N_15342,N_12757,N_13912);
xnor U15343 (N_15343,N_13824,N_12011);
nor U15344 (N_15344,N_12053,N_12052);
nor U15345 (N_15345,N_12960,N_12601);
xor U15346 (N_15346,N_13202,N_13920);
and U15347 (N_15347,N_12285,N_13507);
xnor U15348 (N_15348,N_12950,N_12292);
or U15349 (N_15349,N_12758,N_13613);
xor U15350 (N_15350,N_13857,N_13865);
nand U15351 (N_15351,N_12026,N_12055);
and U15352 (N_15352,N_13620,N_12697);
xor U15353 (N_15353,N_12854,N_13076);
nand U15354 (N_15354,N_12123,N_12431);
and U15355 (N_15355,N_13674,N_12746);
nand U15356 (N_15356,N_13580,N_12068);
xor U15357 (N_15357,N_13450,N_12083);
xnor U15358 (N_15358,N_12842,N_12655);
nor U15359 (N_15359,N_13957,N_12664);
or U15360 (N_15360,N_13441,N_12811);
nor U15361 (N_15361,N_12886,N_12236);
nor U15362 (N_15362,N_12456,N_13009);
xnor U15363 (N_15363,N_12788,N_12916);
nand U15364 (N_15364,N_13075,N_12218);
xor U15365 (N_15365,N_12052,N_12427);
xor U15366 (N_15366,N_12174,N_13810);
or U15367 (N_15367,N_13489,N_13215);
nand U15368 (N_15368,N_13677,N_13270);
nand U15369 (N_15369,N_12263,N_12680);
and U15370 (N_15370,N_13690,N_12275);
xor U15371 (N_15371,N_12353,N_13536);
and U15372 (N_15372,N_12948,N_12436);
xnor U15373 (N_15373,N_12674,N_13664);
or U15374 (N_15374,N_13497,N_13064);
nor U15375 (N_15375,N_12437,N_12066);
and U15376 (N_15376,N_13308,N_12900);
xnor U15377 (N_15377,N_12955,N_13822);
nand U15378 (N_15378,N_12044,N_12887);
and U15379 (N_15379,N_12258,N_12321);
nand U15380 (N_15380,N_12587,N_13595);
nand U15381 (N_15381,N_13519,N_12800);
or U15382 (N_15382,N_13498,N_13178);
and U15383 (N_15383,N_13880,N_12569);
nand U15384 (N_15384,N_12665,N_12778);
nor U15385 (N_15385,N_13139,N_13731);
xnor U15386 (N_15386,N_12699,N_13001);
or U15387 (N_15387,N_12643,N_12264);
or U15388 (N_15388,N_13393,N_12142);
nand U15389 (N_15389,N_12747,N_12138);
nand U15390 (N_15390,N_12820,N_12498);
or U15391 (N_15391,N_13184,N_13955);
nand U15392 (N_15392,N_12601,N_12835);
nor U15393 (N_15393,N_12747,N_13250);
nand U15394 (N_15394,N_13128,N_13822);
and U15395 (N_15395,N_13818,N_12157);
or U15396 (N_15396,N_12229,N_13717);
and U15397 (N_15397,N_12565,N_12611);
and U15398 (N_15398,N_12758,N_13556);
or U15399 (N_15399,N_13557,N_13348);
and U15400 (N_15400,N_13724,N_13635);
nor U15401 (N_15401,N_12881,N_13729);
nand U15402 (N_15402,N_12123,N_12998);
xor U15403 (N_15403,N_13427,N_13608);
nor U15404 (N_15404,N_13493,N_13414);
nor U15405 (N_15405,N_12369,N_12973);
or U15406 (N_15406,N_13681,N_13763);
nand U15407 (N_15407,N_13488,N_13117);
nor U15408 (N_15408,N_12481,N_12725);
nand U15409 (N_15409,N_12582,N_13071);
nand U15410 (N_15410,N_12235,N_12257);
nand U15411 (N_15411,N_13761,N_13242);
nor U15412 (N_15412,N_12032,N_12731);
and U15413 (N_15413,N_12411,N_12929);
xnor U15414 (N_15414,N_13417,N_12355);
and U15415 (N_15415,N_12919,N_13297);
or U15416 (N_15416,N_12167,N_12960);
nor U15417 (N_15417,N_13497,N_13294);
xnor U15418 (N_15418,N_13859,N_13129);
or U15419 (N_15419,N_13715,N_13557);
nor U15420 (N_15420,N_12573,N_12642);
nor U15421 (N_15421,N_12205,N_13298);
or U15422 (N_15422,N_12781,N_13742);
or U15423 (N_15423,N_13968,N_12173);
xor U15424 (N_15424,N_13229,N_12027);
xor U15425 (N_15425,N_13140,N_12703);
and U15426 (N_15426,N_13674,N_13438);
or U15427 (N_15427,N_12310,N_12359);
or U15428 (N_15428,N_13127,N_12935);
nor U15429 (N_15429,N_12365,N_13362);
xnor U15430 (N_15430,N_13126,N_12266);
nand U15431 (N_15431,N_13260,N_12402);
or U15432 (N_15432,N_12617,N_12773);
nor U15433 (N_15433,N_13088,N_12779);
and U15434 (N_15434,N_12809,N_12557);
nor U15435 (N_15435,N_13945,N_12813);
nor U15436 (N_15436,N_13738,N_12986);
nor U15437 (N_15437,N_13292,N_13153);
and U15438 (N_15438,N_12970,N_12957);
nor U15439 (N_15439,N_12877,N_12532);
or U15440 (N_15440,N_13843,N_12622);
xnor U15441 (N_15441,N_13599,N_12554);
nand U15442 (N_15442,N_13149,N_13305);
nor U15443 (N_15443,N_12143,N_13545);
xor U15444 (N_15444,N_12317,N_13114);
and U15445 (N_15445,N_12602,N_13510);
xnor U15446 (N_15446,N_12383,N_13975);
nand U15447 (N_15447,N_12185,N_12373);
nand U15448 (N_15448,N_13042,N_13725);
xor U15449 (N_15449,N_13409,N_12397);
nor U15450 (N_15450,N_12958,N_13747);
nor U15451 (N_15451,N_13664,N_12910);
xnor U15452 (N_15452,N_13271,N_13919);
nor U15453 (N_15453,N_12893,N_13611);
and U15454 (N_15454,N_13268,N_13370);
nand U15455 (N_15455,N_13069,N_12826);
and U15456 (N_15456,N_13704,N_13922);
nor U15457 (N_15457,N_13025,N_13110);
nand U15458 (N_15458,N_13413,N_12959);
or U15459 (N_15459,N_13986,N_12149);
nand U15460 (N_15460,N_12372,N_13083);
nor U15461 (N_15461,N_13184,N_13734);
xnor U15462 (N_15462,N_13197,N_13128);
xor U15463 (N_15463,N_13021,N_13058);
nor U15464 (N_15464,N_13956,N_13064);
xnor U15465 (N_15465,N_13505,N_13995);
nand U15466 (N_15466,N_12939,N_12089);
and U15467 (N_15467,N_12027,N_13475);
nor U15468 (N_15468,N_12242,N_13932);
or U15469 (N_15469,N_12741,N_12303);
nor U15470 (N_15470,N_13623,N_12806);
or U15471 (N_15471,N_12644,N_12770);
nor U15472 (N_15472,N_12418,N_13258);
nand U15473 (N_15473,N_13281,N_13059);
nor U15474 (N_15474,N_13778,N_12006);
nand U15475 (N_15475,N_12241,N_12704);
nand U15476 (N_15476,N_12748,N_13425);
or U15477 (N_15477,N_13925,N_13360);
or U15478 (N_15478,N_12354,N_12390);
nand U15479 (N_15479,N_13511,N_12753);
nor U15480 (N_15480,N_12013,N_13835);
and U15481 (N_15481,N_12318,N_12316);
nand U15482 (N_15482,N_13397,N_13799);
and U15483 (N_15483,N_12915,N_12269);
nand U15484 (N_15484,N_13401,N_12388);
nor U15485 (N_15485,N_12412,N_12989);
or U15486 (N_15486,N_12098,N_13899);
nor U15487 (N_15487,N_13258,N_13949);
and U15488 (N_15488,N_13817,N_12454);
xor U15489 (N_15489,N_13174,N_12384);
or U15490 (N_15490,N_12431,N_12882);
nand U15491 (N_15491,N_13653,N_12358);
nand U15492 (N_15492,N_12642,N_13296);
nor U15493 (N_15493,N_13149,N_12443);
xor U15494 (N_15494,N_12388,N_12985);
xor U15495 (N_15495,N_12327,N_12886);
nor U15496 (N_15496,N_13440,N_12080);
nor U15497 (N_15497,N_12223,N_13153);
or U15498 (N_15498,N_12079,N_12592);
or U15499 (N_15499,N_12447,N_12865);
and U15500 (N_15500,N_13304,N_13417);
nor U15501 (N_15501,N_13536,N_12667);
nand U15502 (N_15502,N_13960,N_12911);
or U15503 (N_15503,N_12022,N_12729);
nor U15504 (N_15504,N_12208,N_12090);
or U15505 (N_15505,N_13246,N_13884);
xor U15506 (N_15506,N_12830,N_12325);
or U15507 (N_15507,N_13785,N_12322);
or U15508 (N_15508,N_12204,N_13098);
xnor U15509 (N_15509,N_12506,N_13305);
and U15510 (N_15510,N_12708,N_12438);
xor U15511 (N_15511,N_12204,N_13875);
nand U15512 (N_15512,N_12275,N_13418);
or U15513 (N_15513,N_13698,N_12410);
xor U15514 (N_15514,N_12795,N_12884);
xor U15515 (N_15515,N_12433,N_12933);
xor U15516 (N_15516,N_12131,N_12133);
or U15517 (N_15517,N_12552,N_13750);
nor U15518 (N_15518,N_13214,N_12720);
nor U15519 (N_15519,N_12113,N_13776);
and U15520 (N_15520,N_12703,N_12971);
xor U15521 (N_15521,N_13231,N_13065);
xnor U15522 (N_15522,N_13718,N_12861);
xnor U15523 (N_15523,N_13826,N_13482);
xor U15524 (N_15524,N_13688,N_13889);
nor U15525 (N_15525,N_13372,N_13738);
nor U15526 (N_15526,N_13366,N_12688);
nand U15527 (N_15527,N_12123,N_13166);
nor U15528 (N_15528,N_13623,N_12790);
nand U15529 (N_15529,N_13916,N_12473);
nor U15530 (N_15530,N_12990,N_12122);
nand U15531 (N_15531,N_12003,N_12542);
xor U15532 (N_15532,N_13891,N_13822);
nand U15533 (N_15533,N_12020,N_13133);
xnor U15534 (N_15534,N_13001,N_13014);
nand U15535 (N_15535,N_12139,N_13538);
nand U15536 (N_15536,N_13352,N_12289);
nand U15537 (N_15537,N_12754,N_12701);
nand U15538 (N_15538,N_13384,N_12094);
xor U15539 (N_15539,N_12378,N_12216);
or U15540 (N_15540,N_12542,N_13891);
nor U15541 (N_15541,N_13515,N_12966);
and U15542 (N_15542,N_13662,N_13755);
or U15543 (N_15543,N_12565,N_13151);
or U15544 (N_15544,N_13233,N_13057);
nand U15545 (N_15545,N_12920,N_12510);
and U15546 (N_15546,N_13756,N_12972);
or U15547 (N_15547,N_13574,N_12206);
nor U15548 (N_15548,N_12938,N_13677);
nand U15549 (N_15549,N_13398,N_13932);
nand U15550 (N_15550,N_13820,N_13179);
xor U15551 (N_15551,N_12602,N_13568);
nor U15552 (N_15552,N_12924,N_12384);
nand U15553 (N_15553,N_12476,N_12783);
or U15554 (N_15554,N_12788,N_13081);
nand U15555 (N_15555,N_13722,N_13941);
and U15556 (N_15556,N_13944,N_12331);
xor U15557 (N_15557,N_13207,N_12337);
and U15558 (N_15558,N_13402,N_13189);
nand U15559 (N_15559,N_12422,N_12789);
xnor U15560 (N_15560,N_12873,N_12748);
nand U15561 (N_15561,N_13000,N_13490);
nand U15562 (N_15562,N_12866,N_12330);
nand U15563 (N_15563,N_12878,N_13355);
xor U15564 (N_15564,N_13974,N_13577);
and U15565 (N_15565,N_12890,N_12101);
or U15566 (N_15566,N_13229,N_13800);
or U15567 (N_15567,N_12930,N_13697);
and U15568 (N_15568,N_12231,N_12247);
xnor U15569 (N_15569,N_13513,N_12841);
nor U15570 (N_15570,N_13847,N_13129);
nand U15571 (N_15571,N_12909,N_13923);
nand U15572 (N_15572,N_13063,N_13206);
and U15573 (N_15573,N_13191,N_12161);
xor U15574 (N_15574,N_12720,N_12220);
or U15575 (N_15575,N_13909,N_13396);
nand U15576 (N_15576,N_12533,N_13234);
xor U15577 (N_15577,N_12836,N_12665);
or U15578 (N_15578,N_12412,N_13485);
and U15579 (N_15579,N_13493,N_13392);
nand U15580 (N_15580,N_13665,N_13032);
nor U15581 (N_15581,N_12131,N_12978);
nor U15582 (N_15582,N_12593,N_13161);
nor U15583 (N_15583,N_13261,N_13079);
and U15584 (N_15584,N_12123,N_13742);
or U15585 (N_15585,N_13103,N_13344);
nor U15586 (N_15586,N_13385,N_12841);
xor U15587 (N_15587,N_13871,N_13897);
xor U15588 (N_15588,N_12411,N_13439);
nor U15589 (N_15589,N_13628,N_12411);
or U15590 (N_15590,N_12378,N_12210);
and U15591 (N_15591,N_13062,N_12624);
nor U15592 (N_15592,N_12090,N_12222);
or U15593 (N_15593,N_12798,N_13314);
xor U15594 (N_15594,N_12275,N_12652);
nand U15595 (N_15595,N_12229,N_12330);
or U15596 (N_15596,N_13373,N_13316);
nor U15597 (N_15597,N_13875,N_13932);
and U15598 (N_15598,N_13268,N_13154);
and U15599 (N_15599,N_13823,N_12612);
nor U15600 (N_15600,N_13129,N_12064);
and U15601 (N_15601,N_13438,N_12454);
nor U15602 (N_15602,N_13347,N_13878);
or U15603 (N_15603,N_13401,N_12232);
and U15604 (N_15604,N_12666,N_13418);
nand U15605 (N_15605,N_13512,N_13846);
nand U15606 (N_15606,N_13854,N_13517);
xor U15607 (N_15607,N_12225,N_12110);
nor U15608 (N_15608,N_13014,N_12067);
or U15609 (N_15609,N_13288,N_13667);
and U15610 (N_15610,N_12160,N_13017);
and U15611 (N_15611,N_13998,N_13479);
and U15612 (N_15612,N_12794,N_12633);
or U15613 (N_15613,N_12838,N_12753);
nor U15614 (N_15614,N_13170,N_13272);
nand U15615 (N_15615,N_13786,N_12141);
nor U15616 (N_15616,N_12391,N_13695);
and U15617 (N_15617,N_12956,N_13832);
or U15618 (N_15618,N_13187,N_12326);
nand U15619 (N_15619,N_12130,N_12513);
nand U15620 (N_15620,N_12689,N_12526);
nor U15621 (N_15621,N_13823,N_12718);
nor U15622 (N_15622,N_13322,N_13213);
nand U15623 (N_15623,N_12435,N_12497);
or U15624 (N_15624,N_12883,N_13587);
nor U15625 (N_15625,N_12058,N_12248);
or U15626 (N_15626,N_12666,N_12312);
nand U15627 (N_15627,N_13322,N_12494);
and U15628 (N_15628,N_12528,N_13055);
and U15629 (N_15629,N_12183,N_13277);
nor U15630 (N_15630,N_12134,N_12928);
and U15631 (N_15631,N_13145,N_13660);
or U15632 (N_15632,N_12045,N_12636);
xor U15633 (N_15633,N_12811,N_12479);
nand U15634 (N_15634,N_12270,N_12073);
nor U15635 (N_15635,N_12163,N_12592);
nand U15636 (N_15636,N_13468,N_13543);
nor U15637 (N_15637,N_13632,N_13661);
nand U15638 (N_15638,N_12315,N_12383);
nor U15639 (N_15639,N_13357,N_12106);
or U15640 (N_15640,N_12247,N_12775);
and U15641 (N_15641,N_12060,N_12727);
nor U15642 (N_15642,N_13604,N_13306);
nor U15643 (N_15643,N_12678,N_12024);
xnor U15644 (N_15644,N_12896,N_13791);
and U15645 (N_15645,N_13488,N_12491);
nand U15646 (N_15646,N_13487,N_12328);
nand U15647 (N_15647,N_13621,N_13900);
or U15648 (N_15648,N_13773,N_13218);
and U15649 (N_15649,N_12291,N_13482);
and U15650 (N_15650,N_13981,N_12259);
and U15651 (N_15651,N_12661,N_12292);
nor U15652 (N_15652,N_12532,N_13234);
nor U15653 (N_15653,N_12060,N_13370);
nor U15654 (N_15654,N_12023,N_13246);
nand U15655 (N_15655,N_13981,N_13319);
and U15656 (N_15656,N_12686,N_12143);
or U15657 (N_15657,N_12805,N_13453);
and U15658 (N_15658,N_12906,N_12040);
nand U15659 (N_15659,N_13688,N_12903);
xnor U15660 (N_15660,N_13981,N_12613);
and U15661 (N_15661,N_12594,N_13788);
and U15662 (N_15662,N_12321,N_12080);
nor U15663 (N_15663,N_12450,N_12587);
nand U15664 (N_15664,N_13767,N_12121);
and U15665 (N_15665,N_12372,N_13024);
or U15666 (N_15666,N_12758,N_12316);
and U15667 (N_15667,N_12172,N_13170);
nand U15668 (N_15668,N_12713,N_13347);
xor U15669 (N_15669,N_13680,N_12948);
nor U15670 (N_15670,N_13652,N_12857);
xor U15671 (N_15671,N_13468,N_12481);
and U15672 (N_15672,N_12724,N_12155);
nand U15673 (N_15673,N_13335,N_12622);
xnor U15674 (N_15674,N_12839,N_12688);
and U15675 (N_15675,N_12385,N_12871);
and U15676 (N_15676,N_13295,N_13960);
or U15677 (N_15677,N_13534,N_12746);
and U15678 (N_15678,N_13900,N_12059);
nor U15679 (N_15679,N_13854,N_13104);
and U15680 (N_15680,N_13132,N_13883);
nand U15681 (N_15681,N_13095,N_12649);
and U15682 (N_15682,N_13356,N_12895);
or U15683 (N_15683,N_13055,N_12767);
xnor U15684 (N_15684,N_12426,N_13937);
nand U15685 (N_15685,N_12258,N_13624);
nor U15686 (N_15686,N_13726,N_13060);
nand U15687 (N_15687,N_12344,N_13742);
or U15688 (N_15688,N_13722,N_12928);
and U15689 (N_15689,N_12214,N_12978);
or U15690 (N_15690,N_12354,N_12667);
nor U15691 (N_15691,N_13241,N_12564);
nand U15692 (N_15692,N_13630,N_12135);
and U15693 (N_15693,N_12778,N_13395);
and U15694 (N_15694,N_13763,N_13931);
nor U15695 (N_15695,N_12819,N_13058);
xor U15696 (N_15696,N_12404,N_13186);
nand U15697 (N_15697,N_13091,N_12682);
nor U15698 (N_15698,N_12434,N_13072);
and U15699 (N_15699,N_13792,N_12879);
nand U15700 (N_15700,N_12523,N_12807);
and U15701 (N_15701,N_13405,N_13791);
xor U15702 (N_15702,N_12734,N_13796);
or U15703 (N_15703,N_12480,N_12567);
nand U15704 (N_15704,N_12368,N_12190);
and U15705 (N_15705,N_12922,N_13753);
nor U15706 (N_15706,N_13999,N_12425);
xor U15707 (N_15707,N_13513,N_12237);
or U15708 (N_15708,N_12858,N_12758);
nand U15709 (N_15709,N_12017,N_12633);
nor U15710 (N_15710,N_13939,N_12463);
or U15711 (N_15711,N_12985,N_12074);
nand U15712 (N_15712,N_12528,N_13663);
or U15713 (N_15713,N_13528,N_13156);
and U15714 (N_15714,N_12989,N_13255);
and U15715 (N_15715,N_13001,N_12210);
xor U15716 (N_15716,N_12113,N_13287);
and U15717 (N_15717,N_13483,N_12201);
nor U15718 (N_15718,N_12833,N_13694);
and U15719 (N_15719,N_13468,N_12030);
and U15720 (N_15720,N_12248,N_12334);
nand U15721 (N_15721,N_13127,N_13051);
nand U15722 (N_15722,N_12227,N_12808);
or U15723 (N_15723,N_12285,N_12136);
and U15724 (N_15724,N_12311,N_12485);
or U15725 (N_15725,N_12504,N_12338);
and U15726 (N_15726,N_13404,N_13807);
and U15727 (N_15727,N_13013,N_13556);
nor U15728 (N_15728,N_13321,N_12248);
xor U15729 (N_15729,N_12421,N_12367);
nand U15730 (N_15730,N_12318,N_13564);
nand U15731 (N_15731,N_13831,N_13706);
and U15732 (N_15732,N_12629,N_13888);
and U15733 (N_15733,N_12999,N_12412);
and U15734 (N_15734,N_12204,N_12405);
xor U15735 (N_15735,N_13929,N_13172);
nand U15736 (N_15736,N_12390,N_12400);
or U15737 (N_15737,N_13665,N_13281);
nor U15738 (N_15738,N_12761,N_12317);
xor U15739 (N_15739,N_13555,N_12702);
and U15740 (N_15740,N_13929,N_12613);
and U15741 (N_15741,N_12704,N_13027);
and U15742 (N_15742,N_13476,N_13534);
or U15743 (N_15743,N_13314,N_12568);
and U15744 (N_15744,N_12350,N_13003);
or U15745 (N_15745,N_13049,N_13146);
and U15746 (N_15746,N_13315,N_12237);
xor U15747 (N_15747,N_12517,N_12690);
and U15748 (N_15748,N_12151,N_13570);
and U15749 (N_15749,N_12883,N_12584);
nor U15750 (N_15750,N_13753,N_12164);
nor U15751 (N_15751,N_12885,N_12348);
nand U15752 (N_15752,N_13188,N_12097);
nor U15753 (N_15753,N_12295,N_12995);
and U15754 (N_15754,N_13709,N_12099);
xnor U15755 (N_15755,N_13362,N_12986);
and U15756 (N_15756,N_13526,N_12325);
nor U15757 (N_15757,N_12279,N_12851);
nor U15758 (N_15758,N_12831,N_12805);
nor U15759 (N_15759,N_12776,N_12854);
nor U15760 (N_15760,N_12316,N_13985);
or U15761 (N_15761,N_13337,N_12767);
or U15762 (N_15762,N_13752,N_12333);
or U15763 (N_15763,N_12091,N_13992);
or U15764 (N_15764,N_13112,N_12727);
nor U15765 (N_15765,N_12860,N_13532);
nand U15766 (N_15766,N_12372,N_13351);
or U15767 (N_15767,N_13103,N_12914);
nand U15768 (N_15768,N_12858,N_12277);
nand U15769 (N_15769,N_13488,N_13536);
and U15770 (N_15770,N_12895,N_13666);
nand U15771 (N_15771,N_13944,N_13924);
and U15772 (N_15772,N_12158,N_12805);
nor U15773 (N_15773,N_12949,N_12586);
and U15774 (N_15774,N_12228,N_13217);
xor U15775 (N_15775,N_12150,N_12577);
or U15776 (N_15776,N_13193,N_12444);
xor U15777 (N_15777,N_13458,N_12327);
xor U15778 (N_15778,N_12758,N_12715);
nand U15779 (N_15779,N_12235,N_12955);
and U15780 (N_15780,N_13335,N_13809);
xnor U15781 (N_15781,N_13668,N_12123);
xor U15782 (N_15782,N_13928,N_13072);
and U15783 (N_15783,N_13455,N_13861);
nor U15784 (N_15784,N_12111,N_13815);
xnor U15785 (N_15785,N_12080,N_12863);
or U15786 (N_15786,N_13181,N_12252);
xor U15787 (N_15787,N_12574,N_13416);
nor U15788 (N_15788,N_12241,N_13138);
xnor U15789 (N_15789,N_13387,N_12315);
xnor U15790 (N_15790,N_12091,N_12960);
and U15791 (N_15791,N_12352,N_12445);
nor U15792 (N_15792,N_12089,N_13900);
nand U15793 (N_15793,N_12733,N_13665);
or U15794 (N_15794,N_13901,N_12378);
nor U15795 (N_15795,N_13415,N_13970);
and U15796 (N_15796,N_12224,N_13917);
xor U15797 (N_15797,N_13326,N_12791);
or U15798 (N_15798,N_12505,N_12146);
and U15799 (N_15799,N_12016,N_12338);
or U15800 (N_15800,N_12574,N_12857);
or U15801 (N_15801,N_13526,N_13824);
xnor U15802 (N_15802,N_12817,N_13990);
and U15803 (N_15803,N_12192,N_13852);
and U15804 (N_15804,N_12581,N_13578);
nand U15805 (N_15805,N_13204,N_12112);
xnor U15806 (N_15806,N_13757,N_13536);
or U15807 (N_15807,N_13247,N_12004);
nor U15808 (N_15808,N_13757,N_12213);
xor U15809 (N_15809,N_13550,N_12013);
and U15810 (N_15810,N_13870,N_12974);
nor U15811 (N_15811,N_13742,N_13882);
or U15812 (N_15812,N_13057,N_13772);
nor U15813 (N_15813,N_12775,N_12440);
nor U15814 (N_15814,N_13976,N_12317);
nor U15815 (N_15815,N_13194,N_12644);
xnor U15816 (N_15816,N_13015,N_12248);
and U15817 (N_15817,N_13968,N_13571);
nand U15818 (N_15818,N_12395,N_12022);
xor U15819 (N_15819,N_13368,N_12302);
or U15820 (N_15820,N_13660,N_12552);
and U15821 (N_15821,N_12229,N_12247);
xnor U15822 (N_15822,N_13875,N_12911);
nor U15823 (N_15823,N_13926,N_13415);
and U15824 (N_15824,N_12596,N_12677);
and U15825 (N_15825,N_12043,N_12125);
and U15826 (N_15826,N_12726,N_12772);
or U15827 (N_15827,N_12730,N_13535);
and U15828 (N_15828,N_12502,N_12624);
or U15829 (N_15829,N_13444,N_12463);
nor U15830 (N_15830,N_12724,N_13578);
or U15831 (N_15831,N_13550,N_12674);
xnor U15832 (N_15832,N_13765,N_12855);
xnor U15833 (N_15833,N_13277,N_12822);
xnor U15834 (N_15834,N_13894,N_13696);
or U15835 (N_15835,N_13168,N_13243);
or U15836 (N_15836,N_13853,N_13899);
and U15837 (N_15837,N_13952,N_12657);
nand U15838 (N_15838,N_13068,N_13178);
and U15839 (N_15839,N_12001,N_12181);
nand U15840 (N_15840,N_13049,N_12781);
nor U15841 (N_15841,N_12690,N_13029);
or U15842 (N_15842,N_13037,N_12687);
xnor U15843 (N_15843,N_12742,N_13579);
nor U15844 (N_15844,N_12458,N_13101);
nand U15845 (N_15845,N_13095,N_12617);
nor U15846 (N_15846,N_13928,N_13159);
or U15847 (N_15847,N_13615,N_12293);
nand U15848 (N_15848,N_13805,N_13988);
nor U15849 (N_15849,N_13354,N_13443);
nand U15850 (N_15850,N_13946,N_12549);
and U15851 (N_15851,N_12619,N_12834);
and U15852 (N_15852,N_13083,N_12033);
nand U15853 (N_15853,N_12571,N_12006);
nand U15854 (N_15854,N_12387,N_12248);
nor U15855 (N_15855,N_12922,N_13534);
nand U15856 (N_15856,N_13427,N_12111);
xor U15857 (N_15857,N_12293,N_13451);
nor U15858 (N_15858,N_13618,N_13757);
xnor U15859 (N_15859,N_12025,N_12079);
and U15860 (N_15860,N_12526,N_12680);
xnor U15861 (N_15861,N_13763,N_13425);
xor U15862 (N_15862,N_12884,N_12872);
or U15863 (N_15863,N_13035,N_12216);
nor U15864 (N_15864,N_13176,N_13330);
nor U15865 (N_15865,N_13959,N_12211);
xor U15866 (N_15866,N_13184,N_13342);
nand U15867 (N_15867,N_13799,N_13811);
xor U15868 (N_15868,N_13938,N_12651);
nor U15869 (N_15869,N_13772,N_13453);
or U15870 (N_15870,N_12678,N_13632);
xnor U15871 (N_15871,N_13047,N_13735);
nand U15872 (N_15872,N_12669,N_12082);
or U15873 (N_15873,N_13523,N_13673);
and U15874 (N_15874,N_12771,N_12453);
nand U15875 (N_15875,N_13105,N_12680);
nand U15876 (N_15876,N_13080,N_12897);
nand U15877 (N_15877,N_13630,N_13179);
nand U15878 (N_15878,N_13933,N_13423);
or U15879 (N_15879,N_12767,N_12617);
and U15880 (N_15880,N_12379,N_13806);
xor U15881 (N_15881,N_13088,N_13368);
nand U15882 (N_15882,N_12994,N_12698);
xor U15883 (N_15883,N_13976,N_12101);
and U15884 (N_15884,N_12273,N_13517);
and U15885 (N_15885,N_13865,N_13908);
or U15886 (N_15886,N_12551,N_13810);
nor U15887 (N_15887,N_13209,N_13049);
and U15888 (N_15888,N_12882,N_12433);
xnor U15889 (N_15889,N_13940,N_12745);
nand U15890 (N_15890,N_12534,N_13961);
or U15891 (N_15891,N_13603,N_13161);
and U15892 (N_15892,N_12794,N_13942);
nand U15893 (N_15893,N_12443,N_12331);
xnor U15894 (N_15894,N_13704,N_13176);
nor U15895 (N_15895,N_12675,N_13634);
nor U15896 (N_15896,N_12232,N_13698);
nand U15897 (N_15897,N_13808,N_12896);
and U15898 (N_15898,N_12575,N_12288);
nand U15899 (N_15899,N_13670,N_12277);
nor U15900 (N_15900,N_13371,N_13400);
nor U15901 (N_15901,N_12764,N_12395);
and U15902 (N_15902,N_13047,N_12405);
nand U15903 (N_15903,N_13798,N_12432);
and U15904 (N_15904,N_12207,N_12675);
or U15905 (N_15905,N_12044,N_13306);
xor U15906 (N_15906,N_12900,N_13417);
xor U15907 (N_15907,N_12652,N_12799);
xnor U15908 (N_15908,N_12672,N_13264);
nand U15909 (N_15909,N_12603,N_13124);
nor U15910 (N_15910,N_12114,N_13840);
or U15911 (N_15911,N_13997,N_12375);
and U15912 (N_15912,N_12634,N_12891);
and U15913 (N_15913,N_12095,N_12879);
and U15914 (N_15914,N_12997,N_13767);
or U15915 (N_15915,N_12479,N_13688);
nand U15916 (N_15916,N_13755,N_12315);
and U15917 (N_15917,N_13005,N_12582);
and U15918 (N_15918,N_13097,N_12423);
or U15919 (N_15919,N_12198,N_13888);
nand U15920 (N_15920,N_13538,N_13193);
xor U15921 (N_15921,N_13149,N_12194);
nand U15922 (N_15922,N_12520,N_12390);
nand U15923 (N_15923,N_12986,N_13281);
nand U15924 (N_15924,N_13932,N_12322);
xnor U15925 (N_15925,N_12633,N_13794);
or U15926 (N_15926,N_12151,N_13421);
nor U15927 (N_15927,N_13786,N_13934);
or U15928 (N_15928,N_13060,N_13485);
or U15929 (N_15929,N_13905,N_13944);
nor U15930 (N_15930,N_12993,N_13694);
xor U15931 (N_15931,N_13976,N_13441);
and U15932 (N_15932,N_12720,N_12848);
nor U15933 (N_15933,N_12420,N_12237);
or U15934 (N_15934,N_13508,N_13476);
or U15935 (N_15935,N_12718,N_13822);
nand U15936 (N_15936,N_12354,N_12981);
nor U15937 (N_15937,N_12757,N_13240);
or U15938 (N_15938,N_12401,N_12612);
xnor U15939 (N_15939,N_13221,N_12701);
nor U15940 (N_15940,N_12297,N_12748);
and U15941 (N_15941,N_12750,N_12906);
nor U15942 (N_15942,N_12397,N_13194);
nand U15943 (N_15943,N_12627,N_13963);
xnor U15944 (N_15944,N_12940,N_12863);
xnor U15945 (N_15945,N_13018,N_13147);
or U15946 (N_15946,N_13913,N_13864);
nand U15947 (N_15947,N_12761,N_13718);
or U15948 (N_15948,N_13661,N_13518);
or U15949 (N_15949,N_13059,N_12792);
and U15950 (N_15950,N_13540,N_13394);
or U15951 (N_15951,N_13345,N_12196);
xor U15952 (N_15952,N_12981,N_12675);
nor U15953 (N_15953,N_13317,N_13468);
or U15954 (N_15954,N_13267,N_12775);
nor U15955 (N_15955,N_12507,N_13142);
nand U15956 (N_15956,N_13552,N_12720);
nand U15957 (N_15957,N_13170,N_12429);
nor U15958 (N_15958,N_13978,N_12212);
nor U15959 (N_15959,N_13587,N_13171);
and U15960 (N_15960,N_12565,N_12644);
nor U15961 (N_15961,N_12863,N_12409);
nand U15962 (N_15962,N_13070,N_12683);
or U15963 (N_15963,N_13416,N_12453);
nor U15964 (N_15964,N_12839,N_12482);
nand U15965 (N_15965,N_13140,N_13207);
and U15966 (N_15966,N_13226,N_13731);
and U15967 (N_15967,N_13677,N_12632);
nor U15968 (N_15968,N_12000,N_13823);
nand U15969 (N_15969,N_12396,N_12890);
nand U15970 (N_15970,N_12380,N_13953);
or U15971 (N_15971,N_12127,N_12578);
or U15972 (N_15972,N_13524,N_12252);
nor U15973 (N_15973,N_13765,N_12303);
nand U15974 (N_15974,N_13199,N_13848);
and U15975 (N_15975,N_12211,N_13238);
nor U15976 (N_15976,N_12036,N_12728);
or U15977 (N_15977,N_13974,N_12943);
and U15978 (N_15978,N_13977,N_12137);
or U15979 (N_15979,N_12241,N_13953);
and U15980 (N_15980,N_13058,N_13322);
xnor U15981 (N_15981,N_13185,N_13779);
xnor U15982 (N_15982,N_13764,N_12905);
nand U15983 (N_15983,N_12116,N_12343);
nand U15984 (N_15984,N_12406,N_13492);
and U15985 (N_15985,N_13931,N_13990);
and U15986 (N_15986,N_12487,N_12935);
or U15987 (N_15987,N_12309,N_13958);
xnor U15988 (N_15988,N_12883,N_13921);
nand U15989 (N_15989,N_13482,N_12421);
or U15990 (N_15990,N_12171,N_13968);
nor U15991 (N_15991,N_13471,N_12688);
xor U15992 (N_15992,N_12608,N_13975);
nand U15993 (N_15993,N_13343,N_12114);
and U15994 (N_15994,N_13240,N_13236);
or U15995 (N_15995,N_13120,N_13897);
xnor U15996 (N_15996,N_12408,N_12945);
and U15997 (N_15997,N_12630,N_13504);
and U15998 (N_15998,N_13282,N_12876);
and U15999 (N_15999,N_12372,N_12310);
or U16000 (N_16000,N_15714,N_15004);
nand U16001 (N_16001,N_15921,N_15616);
nor U16002 (N_16002,N_14878,N_14388);
nand U16003 (N_16003,N_14830,N_14521);
and U16004 (N_16004,N_14938,N_14644);
nand U16005 (N_16005,N_15148,N_14279);
nand U16006 (N_16006,N_14249,N_15003);
nor U16007 (N_16007,N_14678,N_15890);
nand U16008 (N_16008,N_15316,N_14760);
or U16009 (N_16009,N_15906,N_14578);
or U16010 (N_16010,N_14560,N_14164);
xor U16011 (N_16011,N_14302,N_15822);
or U16012 (N_16012,N_15733,N_15274);
nor U16013 (N_16013,N_14787,N_15839);
nor U16014 (N_16014,N_14334,N_14987);
xnor U16015 (N_16015,N_14937,N_14055);
nor U16016 (N_16016,N_14538,N_15641);
or U16017 (N_16017,N_14196,N_15734);
xnor U16018 (N_16018,N_15294,N_15408);
or U16019 (N_16019,N_14243,N_15767);
nor U16020 (N_16020,N_14321,N_14180);
or U16021 (N_16021,N_14147,N_15521);
or U16022 (N_16022,N_15805,N_14033);
nand U16023 (N_16023,N_15357,N_15529);
and U16024 (N_16024,N_14237,N_15830);
xnor U16025 (N_16025,N_14096,N_15423);
or U16026 (N_16026,N_15668,N_15639);
nor U16027 (N_16027,N_14006,N_14268);
or U16028 (N_16028,N_15171,N_14218);
nor U16029 (N_16029,N_14295,N_14308);
nor U16030 (N_16030,N_15591,N_14959);
and U16031 (N_16031,N_14517,N_14478);
xnor U16032 (N_16032,N_14684,N_14383);
and U16033 (N_16033,N_14296,N_15306);
or U16034 (N_16034,N_15178,N_14299);
xor U16035 (N_16035,N_14715,N_14463);
or U16036 (N_16036,N_15273,N_15942);
nand U16037 (N_16037,N_15211,N_15541);
nor U16038 (N_16038,N_14105,N_14947);
or U16039 (N_16039,N_14322,N_15223);
or U16040 (N_16040,N_14373,N_15311);
nand U16041 (N_16041,N_15926,N_15015);
nand U16042 (N_16042,N_15469,N_15545);
xor U16043 (N_16043,N_14624,N_14184);
or U16044 (N_16044,N_14451,N_14958);
and U16045 (N_16045,N_15585,N_14936);
xnor U16046 (N_16046,N_14364,N_15018);
or U16047 (N_16047,N_15910,N_14877);
xnor U16048 (N_16048,N_14792,N_14523);
nand U16049 (N_16049,N_14604,N_14272);
or U16050 (N_16050,N_14428,N_14193);
nor U16051 (N_16051,N_14933,N_14356);
nor U16052 (N_16052,N_14113,N_15950);
nand U16053 (N_16053,N_14853,N_15508);
or U16054 (N_16054,N_14257,N_15676);
nand U16055 (N_16055,N_15502,N_15744);
nand U16056 (N_16056,N_14053,N_14719);
or U16057 (N_16057,N_14355,N_15012);
and U16058 (N_16058,N_15621,N_15738);
nand U16059 (N_16059,N_14532,N_14271);
and U16060 (N_16060,N_14856,N_15033);
or U16061 (N_16061,N_14941,N_15620);
or U16062 (N_16062,N_14804,N_14969);
xor U16063 (N_16063,N_14814,N_15882);
and U16064 (N_16064,N_15358,N_15479);
nor U16065 (N_16065,N_14325,N_14574);
nand U16066 (N_16066,N_15888,N_15704);
xnor U16067 (N_16067,N_15658,N_14262);
xnor U16068 (N_16068,N_15883,N_15908);
nor U16069 (N_16069,N_14362,N_15737);
or U16070 (N_16070,N_14723,N_14945);
and U16071 (N_16071,N_14313,N_15577);
and U16072 (N_16072,N_14772,N_14155);
nand U16073 (N_16073,N_15808,N_15542);
and U16074 (N_16074,N_15602,N_15762);
nand U16075 (N_16075,N_14991,N_14960);
or U16076 (N_16076,N_14426,N_15899);
nor U16077 (N_16077,N_14064,N_15555);
and U16078 (N_16078,N_15080,N_15525);
xnor U16079 (N_16079,N_15834,N_15247);
or U16080 (N_16080,N_14192,N_15538);
xnor U16081 (N_16081,N_15665,N_14570);
nor U16082 (N_16082,N_15261,N_14444);
nor U16083 (N_16083,N_14095,N_15967);
nand U16084 (N_16084,N_15982,N_14032);
nand U16085 (N_16085,N_14762,N_15023);
nor U16086 (N_16086,N_14505,N_15308);
or U16087 (N_16087,N_15233,N_14892);
nor U16088 (N_16088,N_14816,N_14396);
xnor U16089 (N_16089,N_14351,N_14569);
or U16090 (N_16090,N_14980,N_14459);
nor U16091 (N_16091,N_14031,N_14627);
xnor U16092 (N_16092,N_15813,N_15975);
or U16093 (N_16093,N_14763,N_14482);
and U16094 (N_16094,N_15586,N_15401);
or U16095 (N_16095,N_15672,N_14412);
nand U16096 (N_16096,N_14861,N_14005);
or U16097 (N_16097,N_15007,N_15800);
nor U16098 (N_16098,N_15544,N_15938);
xor U16099 (N_16099,N_14658,N_14087);
and U16100 (N_16100,N_14042,N_15703);
xnor U16101 (N_16101,N_15041,N_14316);
and U16102 (N_16102,N_15299,N_14258);
nor U16103 (N_16103,N_15466,N_14798);
nor U16104 (N_16104,N_14977,N_15600);
and U16105 (N_16105,N_14379,N_14725);
and U16106 (N_16106,N_15103,N_15318);
xnor U16107 (N_16107,N_14222,N_14978);
and U16108 (N_16108,N_14007,N_14124);
and U16109 (N_16109,N_15979,N_14994);
or U16110 (N_16110,N_14278,N_14617);
and U16111 (N_16111,N_15201,N_15472);
nor U16112 (N_16112,N_14674,N_15240);
nor U16113 (N_16113,N_15107,N_15901);
xor U16114 (N_16114,N_14669,N_14546);
nand U16115 (N_16115,N_15780,N_15660);
and U16116 (N_16116,N_15409,N_14215);
and U16117 (N_16117,N_15608,N_14447);
xnor U16118 (N_16118,N_14750,N_15393);
xnor U16119 (N_16119,N_14034,N_15073);
and U16120 (N_16120,N_15783,N_14956);
or U16121 (N_16121,N_14389,N_15597);
and U16122 (N_16122,N_14305,N_14718);
nor U16123 (N_16123,N_14866,N_15289);
and U16124 (N_16124,N_15701,N_15027);
or U16125 (N_16125,N_15098,N_15729);
xor U16126 (N_16126,N_14742,N_15803);
nor U16127 (N_16127,N_14775,N_14415);
or U16128 (N_16128,N_14509,N_14361);
and U16129 (N_16129,N_15396,N_15659);
xnor U16130 (N_16130,N_14626,N_14204);
nand U16131 (N_16131,N_15527,N_14484);
nor U16132 (N_16132,N_15885,N_15269);
and U16133 (N_16133,N_15799,N_15109);
xor U16134 (N_16134,N_14199,N_15452);
xnor U16135 (N_16135,N_14900,N_15941);
or U16136 (N_16136,N_14741,N_14551);
nand U16137 (N_16137,N_15194,N_14073);
nand U16138 (N_16138,N_14635,N_15925);
or U16139 (N_16139,N_14771,N_14822);
or U16140 (N_16140,N_14177,N_15939);
and U16141 (N_16141,N_14848,N_15374);
xor U16142 (N_16142,N_14476,N_15126);
or U16143 (N_16143,N_14288,N_14090);
xor U16144 (N_16144,N_14659,N_15909);
nand U16145 (N_16145,N_14185,N_14015);
nor U16146 (N_16146,N_15314,N_15997);
and U16147 (N_16147,N_15112,N_15656);
or U16148 (N_16148,N_15039,N_15286);
and U16149 (N_16149,N_15042,N_15715);
and U16150 (N_16150,N_15111,N_14721);
nand U16151 (N_16151,N_15961,N_14815);
nand U16152 (N_16152,N_14306,N_15172);
nor U16153 (N_16153,N_15420,N_14191);
nand U16154 (N_16154,N_14094,N_15203);
nor U16155 (N_16155,N_14246,N_14609);
and U16156 (N_16156,N_15528,N_15446);
and U16157 (N_16157,N_15645,N_15598);
nor U16158 (N_16158,N_15560,N_14284);
nand U16159 (N_16159,N_14360,N_14893);
nor U16160 (N_16160,N_15666,N_15089);
nand U16161 (N_16161,N_14217,N_15323);
nor U16162 (N_16162,N_14520,N_14758);
or U16163 (N_16163,N_14023,N_14581);
and U16164 (N_16164,N_15313,N_14270);
nand U16165 (N_16165,N_14216,N_14126);
nor U16166 (N_16166,N_15413,N_15363);
nor U16167 (N_16167,N_15492,N_14886);
nand U16168 (N_16168,N_15731,N_14359);
and U16169 (N_16169,N_14766,N_15977);
nand U16170 (N_16170,N_14871,N_15465);
nand U16171 (N_16171,N_15152,N_15784);
xnor U16172 (N_16172,N_14746,N_14139);
nand U16173 (N_16173,N_15721,N_14151);
nor U16174 (N_16174,N_15991,N_14595);
xnor U16175 (N_16175,N_15488,N_14533);
or U16176 (N_16176,N_14357,N_14138);
nor U16177 (N_16177,N_14697,N_15139);
nor U16178 (N_16178,N_15736,N_15030);
nand U16179 (N_16179,N_15853,N_14944);
and U16180 (N_16180,N_15697,N_15686);
xor U16181 (N_16181,N_14130,N_14870);
xnor U16182 (N_16182,N_15695,N_14738);
nand U16183 (N_16183,N_15692,N_14590);
nand U16184 (N_16184,N_14748,N_15275);
xor U16185 (N_16185,N_15722,N_15394);
nand U16186 (N_16186,N_14386,N_14835);
nand U16187 (N_16187,N_15464,N_15128);
xnor U16188 (N_16188,N_14169,N_15045);
nor U16189 (N_16189,N_15747,N_15937);
xnor U16190 (N_16190,N_14083,N_14253);
and U16191 (N_16191,N_14238,N_15779);
xor U16192 (N_16192,N_15589,N_14039);
xor U16193 (N_16193,N_14283,N_14873);
nand U16194 (N_16194,N_14461,N_15129);
and U16195 (N_16195,N_14239,N_14143);
or U16196 (N_16196,N_14384,N_14672);
or U16197 (N_16197,N_14205,N_15617);
xnor U16198 (N_16198,N_15566,N_14378);
xnor U16199 (N_16199,N_15752,N_14012);
xnor U16200 (N_16200,N_14410,N_15681);
or U16201 (N_16201,N_15168,N_14917);
and U16202 (N_16202,N_15213,N_15436);
xor U16203 (N_16203,N_15142,N_14442);
nand U16204 (N_16204,N_15376,N_15724);
nand U16205 (N_16205,N_14225,N_15696);
xnor U16206 (N_16206,N_15110,N_15327);
or U16207 (N_16207,N_14099,N_14558);
nand U16208 (N_16208,N_15694,N_15445);
and U16209 (N_16209,N_15680,N_15758);
nand U16210 (N_16210,N_15305,N_14694);
or U16211 (N_16211,N_15797,N_15386);
nand U16212 (N_16212,N_14739,N_15537);
nor U16213 (N_16213,N_14207,N_14179);
xor U16214 (N_16214,N_14078,N_15993);
nor U16215 (N_16215,N_15079,N_15087);
and U16216 (N_16216,N_14240,N_14770);
nor U16217 (N_16217,N_14988,N_14267);
xor U16218 (N_16218,N_14491,N_15169);
or U16219 (N_16219,N_14757,N_15193);
xnor U16220 (N_16220,N_14690,N_15594);
xor U16221 (N_16221,N_14662,N_14740);
nand U16222 (N_16222,N_14864,N_14883);
nand U16223 (N_16223,N_15075,N_15331);
nor U16224 (N_16224,N_14525,N_15569);
xor U16225 (N_16225,N_15343,N_15412);
nor U16226 (N_16226,N_15277,N_14918);
nor U16227 (N_16227,N_14640,N_15795);
xor U16228 (N_16228,N_14693,N_15051);
or U16229 (N_16229,N_14990,N_14997);
xnor U16230 (N_16230,N_14705,N_15263);
and U16231 (N_16231,N_14160,N_14788);
and U16232 (N_16232,N_15490,N_15264);
or U16233 (N_16233,N_14342,N_14122);
nand U16234 (N_16234,N_15920,N_14374);
xor U16235 (N_16235,N_15625,N_14377);
nor U16236 (N_16236,N_15916,N_14608);
xnor U16237 (N_16237,N_14454,N_15468);
xnor U16238 (N_16238,N_14148,N_14874);
and U16239 (N_16239,N_15857,N_15028);
nor U16240 (N_16240,N_15157,N_14860);
xnor U16241 (N_16241,N_15335,N_14294);
nor U16242 (N_16242,N_14343,N_14974);
nand U16243 (N_16243,N_14691,N_14636);
and U16244 (N_16244,N_14200,N_15367);
or U16245 (N_16245,N_15898,N_15040);
xnor U16246 (N_16246,N_14231,N_14493);
and U16247 (N_16247,N_14811,N_15825);
or U16248 (N_16248,N_14655,N_15361);
nand U16249 (N_16249,N_14565,N_15174);
and U16250 (N_16250,N_15236,N_15842);
nand U16251 (N_16251,N_14474,N_15212);
xor U16252 (N_16252,N_14735,N_14405);
or U16253 (N_16253,N_14001,N_15760);
nor U16254 (N_16254,N_15310,N_15994);
or U16255 (N_16255,N_15662,N_14119);
or U16256 (N_16256,N_15140,N_15561);
xor U16257 (N_16257,N_14080,N_15647);
nand U16258 (N_16258,N_14260,N_14875);
or U16259 (N_16259,N_14986,N_15824);
nand U16260 (N_16260,N_15485,N_15547);
nor U16261 (N_16261,N_15443,N_14531);
nor U16262 (N_16262,N_15471,N_15333);
nand U16263 (N_16263,N_15428,N_15162);
and U16264 (N_16264,N_15410,N_14473);
nand U16265 (N_16265,N_15631,N_15949);
nor U16266 (N_16266,N_15417,N_14108);
xnor U16267 (N_16267,N_14904,N_14110);
nor U16268 (N_16268,N_14320,N_14086);
xnor U16269 (N_16269,N_15802,N_15447);
or U16270 (N_16270,N_15437,N_15182);
xor U16271 (N_16271,N_14752,N_15362);
nand U16272 (N_16272,N_15011,N_14776);
xnor U16273 (N_16273,N_15919,N_14082);
xor U16274 (N_16274,N_14929,N_15959);
xor U16275 (N_16275,N_14477,N_14230);
and U16276 (N_16276,N_14008,N_15978);
nor U16277 (N_16277,N_15536,N_14851);
nand U16278 (N_16278,N_14518,N_14181);
nand U16279 (N_16279,N_14708,N_14158);
xor U16280 (N_16280,N_14176,N_14406);
nor U16281 (N_16281,N_14663,N_14390);
xor U16282 (N_16282,N_14401,N_14354);
nor U16283 (N_16283,N_15849,N_14488);
and U16284 (N_16284,N_15295,N_14371);
or U16285 (N_16285,N_15225,N_15347);
nand U16286 (N_16286,N_15392,N_14779);
nand U16287 (N_16287,N_15014,N_14527);
and U16288 (N_16288,N_15422,N_14004);
nor U16289 (N_16289,N_14955,N_15285);
xnor U16290 (N_16290,N_15298,N_14823);
or U16291 (N_16291,N_14832,N_14729);
or U16292 (N_16292,N_14954,N_15134);
and U16293 (N_16293,N_15083,N_15583);
or U16294 (N_16294,N_14736,N_14774);
nor U16295 (N_16295,N_15161,N_15553);
nand U16296 (N_16296,N_14035,N_14842);
nand U16297 (N_16297,N_15205,N_15596);
and U16298 (N_16298,N_14685,N_14701);
and U16299 (N_16299,N_14496,N_14345);
nand U16300 (N_16300,N_15491,N_15814);
xor U16301 (N_16301,N_15595,N_14602);
or U16302 (N_16302,N_14137,N_14768);
nor U16303 (N_16303,N_14112,N_14976);
nand U16304 (N_16304,N_15054,N_15221);
xor U16305 (N_16305,N_15685,N_15067);
and U16306 (N_16306,N_15931,N_14865);
nand U16307 (N_16307,N_14710,N_14962);
nor U16308 (N_16308,N_14797,N_14510);
nor U16309 (N_16309,N_15850,N_14166);
xor U16310 (N_16310,N_14136,N_14791);
and U16311 (N_16311,N_14924,N_15877);
and U16312 (N_16312,N_14419,N_14472);
or U16313 (N_16313,N_15532,N_15719);
xnor U16314 (N_16314,N_14530,N_14628);
xor U16315 (N_16315,N_15986,N_15682);
nor U16316 (N_16316,N_15293,N_15727);
or U16317 (N_16317,N_14908,N_15001);
and U16318 (N_16318,N_15276,N_14844);
and U16319 (N_16319,N_15930,N_14186);
and U16320 (N_16320,N_15244,N_14115);
and U16321 (N_16321,N_14499,N_14275);
or U16322 (N_16322,N_15699,N_15884);
and U16323 (N_16323,N_15563,N_15279);
or U16324 (N_16324,N_14065,N_14117);
xnor U16325 (N_16325,N_14582,N_15953);
xor U16326 (N_16326,N_15257,N_15047);
or U16327 (N_16327,N_14907,N_14328);
nand U16328 (N_16328,N_15593,N_14985);
nand U16329 (N_16329,N_15092,N_14059);
xor U16330 (N_16330,N_14913,N_14704);
xnor U16331 (N_16331,N_14414,N_14161);
and U16332 (N_16332,N_15066,N_14408);
and U16333 (N_16333,N_15763,N_14398);
and U16334 (N_16334,N_15995,N_15969);
nor U16335 (N_16335,N_14665,N_14413);
or U16336 (N_16336,N_15120,N_15281);
xor U16337 (N_16337,N_14107,N_15966);
or U16338 (N_16338,N_15539,N_15440);
or U16339 (N_16339,N_14048,N_14555);
or U16340 (N_16340,N_14188,N_14026);
or U16341 (N_16341,N_14319,N_15267);
and U16342 (N_16342,N_14011,N_14021);
and U16343 (N_16343,N_14514,N_15749);
nand U16344 (N_16344,N_15913,N_14625);
nor U16345 (N_16345,N_15858,N_15534);
and U16346 (N_16346,N_15973,N_14132);
nor U16347 (N_16347,N_15618,N_15998);
nor U16348 (N_16348,N_14038,N_15280);
nand U16349 (N_16349,N_15136,N_15520);
nor U16350 (N_16350,N_15227,N_15869);
and U16351 (N_16351,N_14706,N_15143);
xnor U16352 (N_16352,N_15068,N_15106);
nand U16353 (N_16353,N_15249,N_14897);
xnor U16354 (N_16354,N_15892,N_15670);
xor U16355 (N_16355,N_14072,N_14067);
xor U16356 (N_16356,N_14599,N_14054);
or U16357 (N_16357,N_15228,N_14661);
nand U16358 (N_16358,N_14149,N_15202);
xor U16359 (N_16359,N_15020,N_15826);
or U16360 (N_16360,N_14572,N_15439);
xor U16361 (N_16361,N_15823,N_14651);
nor U16362 (N_16362,N_14524,N_15918);
or U16363 (N_16363,N_15632,N_14452);
xor U16364 (N_16364,N_15131,N_14767);
nand U16365 (N_16365,N_14887,N_14490);
nand U16366 (N_16366,N_15852,N_15756);
xor U16367 (N_16367,N_14819,N_14261);
nor U16368 (N_16368,N_14097,N_15819);
xor U16369 (N_16369,N_14195,N_14712);
and U16370 (N_16370,N_14547,N_15829);
or U16371 (N_16371,N_14403,N_15968);
nand U16372 (N_16372,N_15880,N_15981);
nand U16373 (N_16373,N_14671,N_15706);
nand U16374 (N_16374,N_15815,N_15354);
or U16375 (N_16375,N_15832,N_15377);
nand U16376 (N_16376,N_14407,N_15667);
xnor U16377 (N_16377,N_15511,N_14202);
xnor U16378 (N_16378,N_15496,N_14562);
and U16379 (N_16379,N_15187,N_14732);
nor U16380 (N_16380,N_15514,N_15630);
and U16381 (N_16381,N_15848,N_15444);
nor U16382 (N_16382,N_15008,N_15914);
and U16383 (N_16383,N_14743,N_14443);
nor U16384 (N_16384,N_15955,N_15652);
nor U16385 (N_16385,N_15772,N_15766);
or U16386 (N_16386,N_14198,N_15024);
nor U16387 (N_16387,N_15530,N_15506);
nor U16388 (N_16388,N_15441,N_15663);
nor U16389 (N_16389,N_14129,N_15765);
nor U16390 (N_16390,N_14382,N_15932);
or U16391 (N_16391,N_14022,N_15096);
nand U16392 (N_16392,N_14504,N_15972);
nor U16393 (N_16393,N_15946,N_14948);
nand U16394 (N_16394,N_15130,N_15404);
nor U16395 (N_16395,N_15700,N_14047);
nor U16396 (N_16396,N_14508,N_15348);
xnor U16397 (N_16397,N_15455,N_14849);
or U16398 (N_16398,N_15461,N_14714);
xor U16399 (N_16399,N_14074,N_15456);
and U16400 (N_16400,N_14939,N_15940);
and U16401 (N_16401,N_15009,N_15642);
nand U16402 (N_16402,N_14722,N_14943);
xor U16403 (N_16403,N_15117,N_15382);
nor U16404 (N_16404,N_14553,N_15032);
or U16405 (N_16405,N_14344,N_15330);
xnor U16406 (N_16406,N_14648,N_15251);
and U16407 (N_16407,N_14675,N_14615);
nand U16408 (N_16408,N_15372,N_14290);
and U16409 (N_16409,N_14392,N_14713);
xnor U16410 (N_16410,N_14983,N_14556);
nor U16411 (N_16411,N_15716,N_15720);
xnor U16412 (N_16412,N_15114,N_15248);
xnor U16413 (N_16413,N_15405,N_14445);
nand U16414 (N_16414,N_15801,N_14934);
or U16415 (N_16415,N_15757,N_15873);
nor U16416 (N_16416,N_14037,N_15153);
nor U16417 (N_16417,N_15198,N_14695);
nand U16418 (N_16418,N_14836,N_14286);
xnor U16419 (N_16419,N_15889,N_15718);
and U16420 (N_16420,N_14820,N_15743);
nor U16421 (N_16421,N_14906,N_15183);
xnor U16422 (N_16422,N_15933,N_14120);
and U16423 (N_16423,N_15498,N_14228);
xor U16424 (N_16424,N_14497,N_15118);
nor U16425 (N_16425,N_15990,N_15470);
or U16426 (N_16426,N_14810,N_14650);
nand U16427 (N_16427,N_15518,N_15352);
nand U16428 (N_16428,N_14336,N_14716);
nor U16429 (N_16429,N_15788,N_15231);
or U16430 (N_16430,N_14058,N_15149);
and U16431 (N_16431,N_15533,N_15615);
or U16432 (N_16432,N_15384,N_14821);
xnor U16433 (N_16433,N_15613,N_15069);
xnor U16434 (N_16434,N_14773,N_15375);
nor U16435 (N_16435,N_15071,N_15606);
nand U16436 (N_16436,N_14614,N_14995);
nor U16437 (N_16437,N_14114,N_15291);
xnor U16438 (N_16438,N_14480,N_15368);
xnor U16439 (N_16439,N_15200,N_15513);
xnor U16440 (N_16440,N_14220,N_15093);
and U16441 (N_16441,N_14764,N_14061);
nor U16442 (N_16442,N_14536,N_15403);
nor U16443 (N_16443,N_15216,N_15454);
or U16444 (N_16444,N_15411,N_15322);
or U16445 (N_16445,N_15255,N_14922);
nor U16446 (N_16446,N_15947,N_15176);
nand U16447 (N_16447,N_14737,N_14855);
and U16448 (N_16448,N_15026,N_15693);
nand U16449 (N_16449,N_14146,N_14395);
or U16450 (N_16450,N_15859,N_14528);
xor U16451 (N_16451,N_15122,N_15177);
xor U16452 (N_16452,N_14173,N_14834);
xor U16453 (N_16453,N_14479,N_15035);
xnor U16454 (N_16454,N_15371,N_14352);
or U16455 (N_16455,N_14300,N_14009);
xnor U16456 (N_16456,N_14068,N_15841);
or U16457 (N_16457,N_14545,N_14639);
or U16458 (N_16458,N_14422,N_15378);
nand U16459 (N_16459,N_14437,N_14197);
xor U16460 (N_16460,N_15059,N_14802);
nor U16461 (N_16461,N_14676,N_14077);
xor U16462 (N_16462,N_14104,N_15369);
or U16463 (N_16463,N_14881,N_15381);
nor U16464 (N_16464,N_15416,N_14968);
nand U16465 (N_16465,N_14254,N_14470);
or U16466 (N_16466,N_14448,N_14541);
xnor U16467 (N_16467,N_15688,N_15207);
or U16468 (N_16468,N_15397,N_15086);
or U16469 (N_16469,N_15056,N_14502);
nand U16470 (N_16470,N_14794,N_15817);
and U16471 (N_16471,N_14466,N_14965);
and U16472 (N_16472,N_14232,N_14433);
xor U16473 (N_16473,N_15980,N_14707);
and U16474 (N_16474,N_15713,N_14621);
nand U16475 (N_16475,N_14411,N_14882);
xnor U16476 (N_16476,N_14311,N_15076);
nor U16477 (N_16477,N_14367,N_14337);
or U16478 (N_16478,N_15818,N_14890);
xnor U16479 (N_16479,N_15791,N_14332);
and U16480 (N_16480,N_14668,N_15809);
or U16481 (N_16481,N_14098,N_15006);
xnor U16482 (N_16482,N_14044,N_15170);
and U16483 (N_16483,N_14314,N_14996);
and U16484 (N_16484,N_14309,N_15677);
and U16485 (N_16485,N_14927,N_15442);
and U16486 (N_16486,N_15655,N_14630);
xnor U16487 (N_16487,N_15970,N_14397);
nand U16488 (N_16488,N_14214,N_15246);
nor U16489 (N_16489,N_14673,N_15774);
nor U16490 (N_16490,N_14588,N_14326);
and U16491 (N_16491,N_15104,N_14157);
or U16492 (N_16492,N_15907,N_15876);
or U16493 (N_16493,N_15296,N_15781);
or U16494 (N_16494,N_14229,N_14394);
xor U16495 (N_16495,N_14002,N_14273);
and U16496 (N_16496,N_14828,N_14656);
or U16497 (N_16497,N_14550,N_15186);
nor U16498 (N_16498,N_14600,N_15345);
and U16499 (N_16499,N_15543,N_14711);
xnor U16500 (N_16500,N_14580,N_14421);
nand U16501 (N_16501,N_14807,N_15215);
xnor U16502 (N_16502,N_14134,N_15552);
xor U16503 (N_16503,N_14167,N_14869);
nand U16504 (N_16504,N_14304,N_14833);
nor U16505 (N_16505,N_14812,N_15497);
xor U16506 (N_16506,N_14040,N_15373);
xnor U16507 (N_16507,N_14680,N_14487);
xnor U16508 (N_16508,N_14456,N_14436);
xnor U16509 (N_16509,N_15708,N_15489);
xnor U16510 (N_16510,N_15151,N_14111);
xor U16511 (N_16511,N_14057,N_15429);
xor U16512 (N_16512,N_14501,N_14076);
nand U16513 (N_16513,N_15951,N_14341);
and U16514 (N_16514,N_15522,N_14781);
nor U16515 (N_16515,N_15964,N_14298);
xor U16516 (N_16516,N_15851,N_14331);
or U16517 (N_16517,N_14416,N_15156);
or U16518 (N_16518,N_15878,N_14393);
or U16519 (N_16519,N_15806,N_15433);
and U16520 (N_16520,N_14862,N_14809);
nand U16521 (N_16521,N_15861,N_15337);
and U16522 (N_16522,N_14857,N_14380);
nor U16523 (N_16523,N_15634,N_14863);
or U16524 (N_16524,N_15678,N_15773);
or U16525 (N_16525,N_14156,N_14803);
and U16526 (N_16526,N_15046,N_15792);
or U16527 (N_16527,N_14686,N_15601);
xor U16528 (N_16528,N_15633,N_15192);
nor U16529 (N_16529,N_14879,N_15989);
nor U16530 (N_16530,N_15728,N_15328);
nand U16531 (N_16531,N_15965,N_15711);
xnor U16532 (N_16532,N_14552,N_15575);
and U16533 (N_16533,N_14079,N_14404);
or U16534 (N_16534,N_14175,N_14102);
or U16535 (N_16535,N_15874,N_15865);
and U16536 (N_16536,N_14657,N_14277);
nand U16537 (N_16537,N_14365,N_14660);
and U16538 (N_16538,N_15432,N_14966);
or U16539 (N_16539,N_15983,N_14567);
and U16540 (N_16540,N_14535,N_15188);
and U16541 (N_16541,N_15984,N_15796);
xor U16542 (N_16542,N_15732,N_15204);
and U16543 (N_16543,N_14561,N_14616);
or U16544 (N_16544,N_15088,N_15777);
nor U16545 (N_16545,N_14914,N_15317);
nand U16546 (N_16546,N_15385,N_15121);
nand U16547 (N_16547,N_14912,N_15838);
nand U16548 (N_16548,N_15426,N_15599);
and U16549 (N_16549,N_14542,N_15266);
nand U16550 (N_16550,N_14841,N_15021);
nand U16551 (N_16551,N_15265,N_15000);
nor U16552 (N_16552,N_14301,N_15929);
or U16553 (N_16553,N_15319,N_15956);
xor U16554 (N_16554,N_15301,N_15388);
or U16555 (N_16555,N_14465,N_15565);
or U16556 (N_16556,N_15759,N_15741);
or U16557 (N_16557,N_14084,N_14586);
nand U16558 (N_16558,N_15283,N_15292);
or U16559 (N_16559,N_14679,N_14441);
nand U16560 (N_16560,N_15451,N_15414);
nor U16561 (N_16561,N_14297,N_14251);
or U16562 (N_16562,N_15340,N_15559);
nand U16563 (N_16563,N_14940,N_14210);
xnor U16564 (N_16564,N_15060,N_14338);
nand U16565 (N_16565,N_15610,N_14646);
xor U16566 (N_16566,N_15935,N_14370);
nor U16567 (N_16567,N_14431,N_15493);
nand U16568 (N_16568,N_14733,N_15504);
and U16569 (N_16569,N_14500,N_14664);
nand U16570 (N_16570,N_15748,N_15936);
nor U16571 (N_16571,N_14385,N_14818);
nor U16572 (N_16572,N_14381,N_14653);
nand U16573 (N_16573,N_14557,N_14790);
or U16574 (N_16574,N_15501,N_14622);
and U16575 (N_16575,N_15769,N_15359);
nand U16576 (N_16576,N_15312,N_15891);
xnor U16577 (N_16577,N_15754,N_14896);
and U16578 (N_16578,N_15840,N_14285);
and U16579 (N_16579,N_15144,N_15903);
xnor U16580 (N_16580,N_14189,N_15029);
and U16581 (N_16581,N_14756,N_14434);
nand U16582 (N_16582,N_15258,N_14566);
xor U16583 (N_16583,N_15836,N_14596);
nor U16584 (N_16584,N_14970,N_15971);
xnor U16585 (N_16585,N_14152,N_15460);
nand U16586 (N_16586,N_14963,N_14513);
and U16587 (N_16587,N_14610,N_15090);
nor U16588 (N_16588,N_15572,N_14647);
or U16589 (N_16589,N_15590,N_14209);
nor U16590 (N_16590,N_15671,N_15775);
nor U16591 (N_16591,N_14455,N_14088);
nand U16592 (N_16592,N_15108,N_15478);
or U16593 (N_16593,N_15821,N_14953);
nor U16594 (N_16594,N_14182,N_15674);
or U16595 (N_16595,N_15637,N_15091);
and U16596 (N_16596,N_15896,N_15095);
or U16597 (N_16597,N_14420,N_15210);
and U16598 (N_16598,N_14638,N_14276);
nand U16599 (N_16599,N_14492,N_15482);
xor U16600 (N_16600,N_14427,N_14506);
or U16601 (N_16601,N_15627,N_14683);
or U16602 (N_16602,N_14526,N_15958);
nand U16603 (N_16603,N_15094,N_14241);
nor U16604 (N_16604,N_14689,N_15048);
xor U16605 (N_16605,N_14916,N_15058);
nand U16606 (N_16606,N_14901,N_14312);
and U16607 (N_16607,N_14245,N_14839);
nand U16608 (N_16608,N_14495,N_15395);
nor U16609 (N_16609,N_14754,N_15626);
nand U16610 (N_16610,N_14142,N_14363);
nand U16611 (N_16611,N_15418,N_14010);
or U16612 (N_16612,N_14793,N_15034);
nor U16613 (N_16613,N_15776,N_15790);
nand U16614 (N_16614,N_15239,N_14335);
or U16615 (N_16615,N_15243,N_15218);
nand U16616 (N_16616,N_14795,N_15019);
and U16617 (N_16617,N_14247,N_14358);
xnor U16618 (N_16618,N_15505,N_14464);
nand U16619 (N_16619,N_14928,N_14439);
nand U16620 (N_16620,N_15831,N_15044);
nor U16621 (N_16621,N_14013,N_14637);
and U16622 (N_16622,N_14806,N_15229);
nor U16623 (N_16623,N_15370,N_14100);
or U16624 (N_16624,N_15897,N_15163);
xnor U16625 (N_16625,N_15584,N_15871);
or U16626 (N_16626,N_14446,N_15189);
nand U16627 (N_16627,N_15224,N_15167);
or U16628 (N_16628,N_14717,N_14785);
nand U16629 (N_16629,N_15175,N_14603);
and U16630 (N_16630,N_15499,N_15619);
xnor U16631 (N_16631,N_14618,N_14872);
nand U16632 (N_16632,N_15341,N_14141);
and U16633 (N_16633,N_14453,N_14782);
nor U16634 (N_16634,N_15687,N_15875);
xnor U16635 (N_16635,N_15057,N_14549);
nor U16636 (N_16636,N_15985,N_15567);
and U16637 (N_16637,N_14071,N_15082);
or U16638 (N_16638,N_14999,N_14745);
xnor U16639 (N_16639,N_15794,N_15603);
nand U16640 (N_16640,N_14780,N_15250);
or U16641 (N_16641,N_14631,N_15562);
xor U16642 (N_16642,N_15811,N_14993);
or U16643 (N_16643,N_15992,N_14085);
or U16644 (N_16644,N_15915,N_14469);
nor U16645 (N_16645,N_15582,N_14777);
nor U16646 (N_16646,N_15070,N_15558);
nor U16647 (N_16647,N_14190,N_14967);
nand U16648 (N_16648,N_14903,N_15957);
or U16649 (N_16649,N_14449,N_14584);
nor U16650 (N_16650,N_15158,N_15576);
and U16651 (N_16651,N_14327,N_15463);
xnor U16652 (N_16652,N_14534,N_15166);
nor U16653 (N_16653,N_14919,N_14417);
nand U16654 (N_16654,N_15726,N_14548);
or U16655 (N_16655,N_15827,N_14784);
xor U16656 (N_16656,N_14154,N_15155);
xor U16657 (N_16657,N_14069,N_14981);
or U16658 (N_16658,N_14537,N_15612);
or U16659 (N_16659,N_14778,N_14529);
nor U16660 (N_16660,N_14244,N_14127);
and U16661 (N_16661,N_15181,N_15270);
nand U16662 (N_16662,N_15526,N_14516);
and U16663 (N_16663,N_15587,N_15487);
xnor U16664 (N_16664,N_15074,N_14891);
or U16665 (N_16665,N_15016,N_15866);
nand U16666 (N_16666,N_15649,N_14366);
and U16667 (N_16667,N_14387,N_15307);
or U16668 (N_16668,N_14457,N_14063);
nor U16669 (N_16669,N_15654,N_15462);
or U16670 (N_16670,N_15551,N_15364);
nor U16671 (N_16671,N_14025,N_15988);
xnor U16672 (N_16672,N_14540,N_14643);
xnor U16673 (N_16673,N_15164,N_15862);
or U16674 (N_16674,N_15053,N_14347);
and U16675 (N_16675,N_15657,N_15304);
and U16676 (N_16676,N_15450,N_15770);
xor U16677 (N_16677,N_15100,N_14350);
and U16678 (N_16678,N_14611,N_15287);
nand U16679 (N_16679,N_14573,N_15467);
nand U16680 (N_16680,N_15816,N_14168);
nand U16681 (N_16681,N_15868,N_15554);
xor U16682 (N_16682,N_15365,N_14753);
nand U16683 (N_16683,N_15510,N_15116);
nand U16684 (N_16684,N_14642,N_14315);
or U16685 (N_16685,N_14755,N_14221);
or U16686 (N_16686,N_14589,N_14046);
and U16687 (N_16687,N_14435,N_14623);
and U16688 (N_16688,N_14587,N_14020);
and U16689 (N_16689,N_15415,N_14730);
and U16690 (N_16690,N_14165,N_14989);
nand U16691 (N_16691,N_15355,N_14749);
nor U16692 (N_16692,N_14799,N_15260);
nand U16693 (N_16693,N_14952,N_14888);
nand U16694 (N_16694,N_15383,N_15419);
xor U16695 (N_16695,N_15288,N_14424);
and U16696 (N_16696,N_15324,N_15844);
nor U16697 (N_16697,N_15923,N_14645);
nand U16698 (N_16698,N_15350,N_15425);
nor U16699 (N_16699,N_14266,N_15302);
and U16700 (N_16700,N_14789,N_15278);
and U16701 (N_16701,N_15256,N_15448);
and U16702 (N_16702,N_14174,N_15135);
or U16703 (N_16703,N_14605,N_14670);
and U16704 (N_16704,N_15389,N_15325);
nor U16705 (N_16705,N_15119,N_15237);
and U16706 (N_16706,N_14219,N_15179);
nor U16707 (N_16707,N_15651,N_14579);
or U16708 (N_16708,N_14349,N_14607);
xor U16709 (N_16709,N_14957,N_15475);
or U16710 (N_16710,N_15253,N_15854);
nand U16711 (N_16711,N_15962,N_15424);
nor U16712 (N_16712,N_15105,N_14682);
xor U16713 (N_16713,N_14423,N_15614);
nand U16714 (N_16714,N_14583,N_14353);
xnor U16715 (N_16715,N_14041,N_14052);
or U16716 (N_16716,N_15191,N_15945);
nand U16717 (N_16717,N_14979,N_14880);
nand U16718 (N_16718,N_15458,N_14485);
nand U16719 (N_16719,N_14018,N_14858);
or U16720 (N_16720,N_15740,N_14850);
nor U16721 (N_16721,N_15764,N_14187);
nor U16722 (N_16722,N_14131,N_14992);
nand U16723 (N_16723,N_15507,N_15531);
nor U16724 (N_16724,N_15833,N_14728);
and U16725 (N_16725,N_14634,N_14961);
nand U16726 (N_16726,N_15588,N_14667);
nor U16727 (N_16727,N_14211,N_14571);
nor U16728 (N_16728,N_14091,N_15739);
and U16729 (N_16729,N_15477,N_15241);
nor U16730 (N_16730,N_14734,N_15623);
nor U16731 (N_16731,N_14905,N_14418);
or U16732 (N_16732,N_14703,N_15629);
xor U16733 (N_16733,N_15689,N_14089);
xnor U16734 (N_16734,N_14075,N_14236);
nand U16735 (N_16735,N_15101,N_15010);
and U16736 (N_16736,N_15607,N_14677);
or U16737 (N_16737,N_15987,N_14688);
and U16738 (N_16738,N_14935,N_14081);
or U16739 (N_16739,N_14761,N_14543);
nand U16740 (N_16740,N_15217,N_14150);
nand U16741 (N_16741,N_15761,N_15535);
or U16742 (N_16742,N_14515,N_15895);
and U16743 (N_16743,N_14593,N_15702);
nand U16744 (N_16744,N_15725,N_14003);
xor U16745 (N_16745,N_14498,N_15043);
or U16746 (N_16746,N_14594,N_14696);
and U16747 (N_16747,N_14121,N_14213);
xnor U16748 (N_16748,N_14183,N_14840);
nor U16749 (N_16749,N_14103,N_15782);
or U16750 (N_16750,N_15334,N_15353);
or U16751 (N_16751,N_15902,N_14931);
or U16752 (N_16752,N_15160,N_14591);
nor U16753 (N_16753,N_14925,N_14265);
and U16754 (N_16754,N_15391,N_15480);
xor U16755 (N_16755,N_15449,N_15592);
or U16756 (N_16756,N_15390,N_15102);
nor U16757 (N_16757,N_15081,N_14829);
or U16758 (N_16758,N_15709,N_14923);
nor U16759 (N_16759,N_15481,N_15342);
and U16760 (N_16760,N_15234,N_15315);
xnor U16761 (N_16761,N_14606,N_15282);
xnor U16762 (N_16762,N_14727,N_15879);
and U16763 (N_16763,N_14281,N_15579);
xor U16764 (N_16764,N_14751,N_14264);
and U16765 (N_16765,N_15646,N_15500);
and U16766 (N_16766,N_15664,N_14425);
or U16767 (N_16767,N_14471,N_14369);
xnor U16768 (N_16768,N_14932,N_14287);
nor U16769 (N_16769,N_14062,N_15271);
nor U16770 (N_16770,N_15690,N_15976);
nand U16771 (N_16771,N_15300,N_15077);
or U16772 (N_16772,N_14876,N_15556);
or U16773 (N_16773,N_15828,N_14223);
or U16774 (N_16774,N_14116,N_14726);
or U16775 (N_16775,N_15745,N_14269);
nor U16776 (N_16776,N_15820,N_14926);
nand U16777 (N_16777,N_15398,N_15065);
nor U16778 (N_16778,N_15113,N_14178);
and U16779 (N_16779,N_14585,N_14340);
and U16780 (N_16780,N_14093,N_15887);
or U16781 (N_16781,N_15948,N_14894);
xor U16782 (N_16782,N_15434,N_15356);
or U16783 (N_16783,N_14597,N_15768);
or U16784 (N_16784,N_15934,N_14837);
and U16785 (N_16785,N_15924,N_14769);
and U16786 (N_16786,N_14280,N_14051);
nand U16787 (N_16787,N_15999,N_15038);
nand U16788 (N_16788,N_14028,N_14024);
xnor U16789 (N_16789,N_15943,N_15845);
nor U16790 (N_16790,N_15219,N_15421);
nand U16791 (N_16791,N_14400,N_14303);
or U16792 (N_16792,N_14709,N_14133);
and U16793 (N_16793,N_15127,N_14845);
and U16794 (N_16794,N_14291,N_14125);
or U16795 (N_16795,N_15366,N_15855);
xnor U16796 (N_16796,N_15185,N_14563);
and U16797 (N_16797,N_15184,N_14234);
and U16798 (N_16798,N_15332,N_14971);
or U16799 (N_16799,N_14666,N_15459);
xnor U16800 (N_16800,N_14826,N_15125);
or U16801 (N_16801,N_14274,N_14731);
and U16802 (N_16802,N_15062,N_15611);
nand U16803 (N_16803,N_14786,N_14838);
and U16804 (N_16804,N_15512,N_14263);
or U16805 (N_16805,N_15326,N_15960);
xor U16806 (N_16806,N_15870,N_14014);
nand U16807 (N_16807,N_15837,N_15195);
or U16808 (N_16808,N_14203,N_15133);
nand U16809 (N_16809,N_14641,N_15351);
and U16810 (N_16810,N_14045,N_15474);
xor U16811 (N_16811,N_15735,N_14118);
xnor U16812 (N_16812,N_14512,N_15846);
or U16813 (N_16813,N_14376,N_14511);
or U16814 (N_16814,N_14212,N_15379);
or U16815 (N_16815,N_15078,N_14507);
or U16816 (N_16816,N_14019,N_15519);
and U16817 (N_16817,N_15843,N_15123);
xnor U16818 (N_16818,N_15049,N_15580);
nor U16819 (N_16819,N_14889,N_14503);
xor U16820 (N_16820,N_14206,N_14592);
nor U16821 (N_16821,N_14483,N_15675);
and U16822 (N_16822,N_14317,N_14092);
xnor U16823 (N_16823,N_15180,N_15771);
and U16824 (N_16824,N_15785,N_14577);
nand U16825 (N_16825,N_15571,N_15025);
or U16826 (N_16826,N_15321,N_15476);
nand U16827 (N_16827,N_14050,N_14171);
xnor U16828 (N_16828,N_15214,N_15329);
or U16829 (N_16829,N_15473,N_15640);
nand U16830 (N_16830,N_14747,N_15564);
nor U16831 (N_16831,N_15886,N_15628);
xnor U16832 (N_16832,N_15807,N_15402);
or U16833 (N_16833,N_14293,N_14432);
nand U16834 (N_16834,N_15917,N_15206);
or U16835 (N_16835,N_15549,N_15427);
nand U16836 (N_16836,N_15712,N_14796);
xnor U16837 (N_16837,N_15284,N_14964);
xnor U16838 (N_16838,N_15578,N_15272);
xor U16839 (N_16839,N_15636,N_14066);
and U16840 (N_16840,N_15573,N_15309);
nor U16841 (N_16841,N_15900,N_14681);
nand U16842 (N_16842,N_14982,N_15483);
xnor U16843 (N_16843,N_14462,N_14915);
nand U16844 (N_16844,N_15196,N_14885);
nand U16845 (N_16845,N_14998,N_14475);
nand U16846 (N_16846,N_14884,N_14030);
nand U16847 (N_16847,N_14481,N_14468);
and U16848 (N_16848,N_15050,N_15635);
xnor U16849 (N_16849,N_15523,N_14902);
nor U16850 (N_16850,N_14951,N_14700);
xnor U16851 (N_16851,N_14930,N_14194);
nor U16852 (N_16852,N_14942,N_15810);
or U16853 (N_16853,N_15604,N_14486);
nor U16854 (N_16854,N_15540,N_14601);
nand U16855 (N_16855,N_14765,N_14330);
xor U16856 (N_16856,N_14973,N_15648);
and U16857 (N_16857,N_14652,N_15515);
nor U16858 (N_16858,N_14895,N_15339);
xor U16859 (N_16859,N_14522,N_14460);
nand U16860 (N_16860,N_14619,N_14430);
or U16861 (N_16861,N_15005,N_15864);
and U16862 (N_16862,N_14946,N_14162);
nor U16863 (N_16863,N_15036,N_15746);
nand U16864 (N_16864,N_14256,N_15638);
nor U16865 (N_16865,N_15723,N_15173);
xnor U16866 (N_16866,N_15550,N_15052);
xor U16867 (N_16867,N_15683,N_15254);
nor U16868 (N_16868,N_14827,N_14554);
and U16869 (N_16869,N_15669,N_14153);
or U16870 (N_16870,N_14720,N_15856);
or U16871 (N_16871,N_14898,N_14613);
xor U16872 (N_16872,N_14144,N_14984);
and U16873 (N_16873,N_14049,N_15320);
nand U16874 (N_16874,N_14450,N_15208);
and U16875 (N_16875,N_14519,N_15303);
nor U16876 (N_16876,N_14783,N_15145);
xor U16877 (N_16877,N_15431,N_14235);
nor U16878 (N_16878,N_14744,N_14226);
nor U16879 (N_16879,N_14252,N_15904);
and U16880 (N_16880,N_14224,N_14805);
xnor U16881 (N_16881,N_14318,N_14950);
nand U16882 (N_16882,N_15653,N_15055);
nor U16883 (N_16883,N_15037,N_14016);
nand U16884 (N_16884,N_15238,N_14201);
and U16885 (N_16885,N_15730,N_15974);
nand U16886 (N_16886,N_15605,N_15624);
nor U16887 (N_16887,N_15812,N_14544);
nor U16888 (N_16888,N_15644,N_15742);
nand U16889 (N_16889,N_14629,N_15268);
xor U16890 (N_16890,N_14036,N_15691);
nand U16891 (N_16891,N_14867,N_14843);
or U16892 (N_16892,N_14698,N_14489);
nor U16893 (N_16893,N_15661,N_15905);
or U16894 (N_16894,N_14724,N_14060);
nor U16895 (N_16895,N_15022,N_15717);
xor U16896 (N_16896,N_14825,N_15778);
or U16897 (N_16897,N_15486,N_14140);
nand U16898 (N_16898,N_15072,N_14846);
and U16899 (N_16899,N_15574,N_15509);
xor U16900 (N_16900,N_14163,N_15235);
nand U16901 (N_16901,N_15996,N_14831);
and U16902 (N_16902,N_14307,N_14282);
xor U16903 (N_16903,N_14043,N_15013);
nor U16904 (N_16904,N_14128,N_15400);
nand U16905 (N_16905,N_14633,N_14109);
and U16906 (N_16906,N_14975,N_15753);
and U16907 (N_16907,N_15643,N_15798);
xnor U16908 (N_16908,N_15146,N_15548);
and U16909 (N_16909,N_14292,N_14559);
nand U16910 (N_16910,N_14372,N_14911);
xnor U16911 (N_16911,N_14494,N_15380);
nor U16912 (N_16912,N_15457,N_15349);
nand U16913 (N_16913,N_15159,N_14248);
nand U16914 (N_16914,N_15755,N_14242);
nor U16915 (N_16915,N_15115,N_15399);
or U16916 (N_16916,N_14612,N_15230);
xnor U16917 (N_16917,N_15085,N_14654);
xnor U16918 (N_16918,N_14145,N_15707);
or U16919 (N_16919,N_14135,N_14568);
or U16920 (N_16920,N_15787,N_14467);
and U16921 (N_16921,N_15705,N_14692);
and U16922 (N_16922,N_14333,N_15099);
nand U16923 (N_16923,N_14106,N_15097);
and U16924 (N_16924,N_14620,N_14699);
or U16925 (N_16925,N_15503,N_15259);
xnor U16926 (N_16926,N_14575,N_15952);
xor U16927 (N_16927,N_15138,N_15245);
xnor U16928 (N_16928,N_15252,N_14310);
nor U16929 (N_16929,N_14170,N_15137);
nand U16930 (N_16930,N_14817,N_14056);
or U16931 (N_16931,N_14346,N_15872);
xor U16932 (N_16932,N_14972,N_15609);
nor U16933 (N_16933,N_14399,N_14391);
nor U16934 (N_16934,N_14259,N_15453);
xor U16935 (N_16935,N_15804,N_14458);
and U16936 (N_16936,N_15710,N_14233);
or U16937 (N_16937,N_14921,N_15406);
nor U16938 (N_16938,N_14440,N_15494);
nand U16939 (N_16939,N_15061,N_14899);
nor U16940 (N_16940,N_15209,N_15894);
and U16941 (N_16941,N_15338,N_15154);
nand U16942 (N_16942,N_14029,N_15570);
nand U16943 (N_16943,N_14429,N_15017);
and U16944 (N_16944,N_15673,N_14027);
or U16945 (N_16945,N_15963,N_15495);
xor U16946 (N_16946,N_14123,N_14868);
nor U16947 (N_16947,N_15484,N_14687);
nand U16948 (N_16948,N_15297,N_15911);
or U16949 (N_16949,N_15622,N_14324);
xnor U16950 (N_16950,N_15360,N_15881);
xor U16951 (N_16951,N_15084,N_15242);
nand U16952 (N_16952,N_14070,N_15222);
or U16953 (N_16953,N_14375,N_15698);
nand U16954 (N_16954,N_15435,N_14564);
nor U16955 (N_16955,N_15262,N_15165);
nand U16956 (N_16956,N_15793,N_14909);
xnor U16957 (N_16957,N_15860,N_14255);
and U16958 (N_16958,N_14539,N_14632);
or U16959 (N_16959,N_15557,N_14172);
nand U16960 (N_16960,N_15430,N_15002);
nor U16961 (N_16961,N_15954,N_15346);
and U16962 (N_16962,N_15064,N_15517);
nor U16963 (N_16963,N_15581,N_14598);
or U16964 (N_16964,N_15031,N_15928);
nand U16965 (N_16965,N_15751,N_14808);
or U16966 (N_16966,N_15344,N_15232);
and U16967 (N_16967,N_14859,N_15922);
or U16968 (N_16968,N_15438,N_15132);
xnor U16969 (N_16969,N_15226,N_15524);
nor U16970 (N_16970,N_15190,N_15516);
or U16971 (N_16971,N_15893,N_15407);
or U16972 (N_16972,N_14649,N_14910);
or U16973 (N_16973,N_15336,N_14854);
and U16974 (N_16974,N_14402,N_14702);
and U16975 (N_16975,N_14813,N_14289);
xnor U16976 (N_16976,N_14847,N_14368);
xnor U16977 (N_16977,N_15546,N_15750);
and U16978 (N_16978,N_14101,N_14949);
xor U16979 (N_16979,N_15863,N_15387);
xor U16980 (N_16980,N_14759,N_14348);
xnor U16981 (N_16981,N_15568,N_15650);
xnor U16982 (N_16982,N_14801,N_15679);
nand U16983 (N_16983,N_14208,N_15290);
and U16984 (N_16984,N_14000,N_15789);
xnor U16985 (N_16985,N_15124,N_15835);
and U16986 (N_16986,N_15927,N_15141);
nand U16987 (N_16987,N_14824,N_15867);
xor U16988 (N_16988,N_15912,N_14409);
and U16989 (N_16989,N_14250,N_14323);
nand U16990 (N_16990,N_15197,N_14852);
or U16991 (N_16991,N_15684,N_14227);
or U16992 (N_16992,N_14017,N_15786);
or U16993 (N_16993,N_14800,N_15847);
and U16994 (N_16994,N_14438,N_15220);
nand U16995 (N_16995,N_14159,N_14576);
xor U16996 (N_16996,N_15150,N_15944);
nor U16997 (N_16997,N_14920,N_15063);
nor U16998 (N_16998,N_15147,N_14339);
and U16999 (N_16999,N_14329,N_15199);
nand U17000 (N_17000,N_15768,N_15886);
or U17001 (N_17001,N_15134,N_14542);
nor U17002 (N_17002,N_15067,N_15090);
or U17003 (N_17003,N_15639,N_14811);
nor U17004 (N_17004,N_14447,N_15830);
or U17005 (N_17005,N_15824,N_14484);
nand U17006 (N_17006,N_14976,N_14496);
xor U17007 (N_17007,N_14315,N_14716);
xor U17008 (N_17008,N_14792,N_14210);
or U17009 (N_17009,N_15243,N_14392);
nor U17010 (N_17010,N_15504,N_15934);
xnor U17011 (N_17011,N_14122,N_14388);
nand U17012 (N_17012,N_14817,N_15912);
or U17013 (N_17013,N_14860,N_14605);
nor U17014 (N_17014,N_15526,N_14776);
nor U17015 (N_17015,N_14718,N_14863);
and U17016 (N_17016,N_14795,N_15219);
and U17017 (N_17017,N_14496,N_15411);
and U17018 (N_17018,N_14056,N_14323);
xnor U17019 (N_17019,N_14728,N_15160);
or U17020 (N_17020,N_14821,N_15565);
or U17021 (N_17021,N_15981,N_15947);
nand U17022 (N_17022,N_15057,N_14282);
or U17023 (N_17023,N_14771,N_14500);
and U17024 (N_17024,N_14653,N_14132);
xnor U17025 (N_17025,N_14047,N_15000);
and U17026 (N_17026,N_14129,N_15119);
and U17027 (N_17027,N_15990,N_15918);
nor U17028 (N_17028,N_15518,N_15263);
or U17029 (N_17029,N_14395,N_14758);
nor U17030 (N_17030,N_15751,N_14035);
xnor U17031 (N_17031,N_14963,N_15115);
nand U17032 (N_17032,N_15038,N_14211);
nand U17033 (N_17033,N_15099,N_15782);
and U17034 (N_17034,N_15583,N_14661);
or U17035 (N_17035,N_14040,N_15075);
or U17036 (N_17036,N_14745,N_15671);
xnor U17037 (N_17037,N_15650,N_14751);
or U17038 (N_17038,N_14490,N_15792);
nand U17039 (N_17039,N_14364,N_15269);
or U17040 (N_17040,N_15112,N_15784);
and U17041 (N_17041,N_15109,N_14903);
nand U17042 (N_17042,N_15972,N_15372);
and U17043 (N_17043,N_15057,N_14760);
or U17044 (N_17044,N_14513,N_14458);
or U17045 (N_17045,N_15081,N_15571);
nor U17046 (N_17046,N_14118,N_14690);
xnor U17047 (N_17047,N_15331,N_15002);
and U17048 (N_17048,N_14528,N_15760);
nor U17049 (N_17049,N_15861,N_14423);
nor U17050 (N_17050,N_15265,N_14453);
and U17051 (N_17051,N_14385,N_15495);
and U17052 (N_17052,N_15028,N_14237);
and U17053 (N_17053,N_14521,N_15124);
or U17054 (N_17054,N_14504,N_15971);
xor U17055 (N_17055,N_14365,N_14128);
or U17056 (N_17056,N_14810,N_15407);
or U17057 (N_17057,N_14455,N_15903);
nor U17058 (N_17058,N_15456,N_15563);
and U17059 (N_17059,N_15794,N_14914);
nand U17060 (N_17060,N_14781,N_15141);
xor U17061 (N_17061,N_15118,N_14698);
or U17062 (N_17062,N_14172,N_15729);
or U17063 (N_17063,N_14780,N_14776);
nand U17064 (N_17064,N_15023,N_15979);
or U17065 (N_17065,N_15413,N_15080);
nand U17066 (N_17066,N_14941,N_15677);
and U17067 (N_17067,N_15064,N_14781);
nor U17068 (N_17068,N_14191,N_15630);
nand U17069 (N_17069,N_15746,N_14251);
xor U17070 (N_17070,N_15278,N_15025);
xnor U17071 (N_17071,N_15806,N_14233);
nand U17072 (N_17072,N_14503,N_15551);
or U17073 (N_17073,N_15424,N_14795);
nor U17074 (N_17074,N_14093,N_14981);
nor U17075 (N_17075,N_14087,N_14954);
nand U17076 (N_17076,N_14610,N_15690);
and U17077 (N_17077,N_14828,N_14885);
nand U17078 (N_17078,N_15504,N_15369);
nand U17079 (N_17079,N_14867,N_15908);
or U17080 (N_17080,N_14476,N_15276);
nor U17081 (N_17081,N_14722,N_15032);
xnor U17082 (N_17082,N_14133,N_15757);
nand U17083 (N_17083,N_15191,N_15075);
xnor U17084 (N_17084,N_15245,N_14027);
nand U17085 (N_17085,N_15044,N_14896);
nand U17086 (N_17086,N_15693,N_14250);
or U17087 (N_17087,N_15259,N_14549);
nor U17088 (N_17088,N_15914,N_15896);
or U17089 (N_17089,N_14745,N_14815);
nor U17090 (N_17090,N_15266,N_14414);
or U17091 (N_17091,N_15674,N_14172);
xnor U17092 (N_17092,N_15683,N_15410);
nand U17093 (N_17093,N_15264,N_15244);
or U17094 (N_17094,N_15164,N_14837);
nand U17095 (N_17095,N_15715,N_15929);
nand U17096 (N_17096,N_15628,N_15793);
nor U17097 (N_17097,N_14934,N_15286);
nor U17098 (N_17098,N_14011,N_14556);
and U17099 (N_17099,N_15045,N_15267);
xnor U17100 (N_17100,N_15413,N_15852);
nand U17101 (N_17101,N_15538,N_15271);
or U17102 (N_17102,N_15438,N_15465);
and U17103 (N_17103,N_14516,N_14610);
nand U17104 (N_17104,N_14033,N_14532);
xnor U17105 (N_17105,N_14515,N_14882);
and U17106 (N_17106,N_15776,N_15899);
or U17107 (N_17107,N_15648,N_14498);
nor U17108 (N_17108,N_15484,N_14247);
and U17109 (N_17109,N_14865,N_14124);
nor U17110 (N_17110,N_14863,N_14368);
xor U17111 (N_17111,N_15086,N_14060);
or U17112 (N_17112,N_15566,N_15544);
nand U17113 (N_17113,N_15670,N_14690);
xnor U17114 (N_17114,N_15601,N_14659);
and U17115 (N_17115,N_15074,N_15095);
nand U17116 (N_17116,N_15447,N_14088);
or U17117 (N_17117,N_15905,N_14059);
xor U17118 (N_17118,N_14832,N_14335);
and U17119 (N_17119,N_15110,N_15283);
and U17120 (N_17120,N_14359,N_14413);
nand U17121 (N_17121,N_15463,N_14799);
nand U17122 (N_17122,N_15238,N_14470);
or U17123 (N_17123,N_14135,N_14919);
nand U17124 (N_17124,N_15205,N_14861);
xor U17125 (N_17125,N_14619,N_15685);
and U17126 (N_17126,N_15814,N_15976);
nand U17127 (N_17127,N_14155,N_14682);
and U17128 (N_17128,N_14699,N_14341);
nand U17129 (N_17129,N_14921,N_14386);
or U17130 (N_17130,N_14924,N_14443);
or U17131 (N_17131,N_14438,N_14654);
or U17132 (N_17132,N_14255,N_15888);
or U17133 (N_17133,N_14852,N_14590);
xnor U17134 (N_17134,N_14195,N_15986);
and U17135 (N_17135,N_15107,N_14432);
or U17136 (N_17136,N_15894,N_15380);
nor U17137 (N_17137,N_15865,N_15277);
nand U17138 (N_17138,N_14969,N_14438);
and U17139 (N_17139,N_15261,N_15207);
and U17140 (N_17140,N_15400,N_15345);
nor U17141 (N_17141,N_14465,N_14925);
or U17142 (N_17142,N_14789,N_14444);
xor U17143 (N_17143,N_14129,N_15121);
and U17144 (N_17144,N_15876,N_15015);
or U17145 (N_17145,N_14635,N_14333);
and U17146 (N_17146,N_14074,N_15924);
and U17147 (N_17147,N_15034,N_14954);
and U17148 (N_17148,N_14142,N_14750);
nor U17149 (N_17149,N_15153,N_15746);
or U17150 (N_17150,N_15923,N_15574);
nand U17151 (N_17151,N_15929,N_14154);
or U17152 (N_17152,N_14377,N_14645);
xor U17153 (N_17153,N_15527,N_14910);
nand U17154 (N_17154,N_15102,N_15515);
or U17155 (N_17155,N_14310,N_15198);
nand U17156 (N_17156,N_15785,N_14035);
nand U17157 (N_17157,N_14688,N_14201);
or U17158 (N_17158,N_15552,N_15946);
or U17159 (N_17159,N_15920,N_14134);
xnor U17160 (N_17160,N_15278,N_15427);
nand U17161 (N_17161,N_15112,N_14148);
or U17162 (N_17162,N_14216,N_14597);
nand U17163 (N_17163,N_14854,N_15691);
or U17164 (N_17164,N_14983,N_14960);
and U17165 (N_17165,N_15570,N_15335);
and U17166 (N_17166,N_15272,N_15922);
xnor U17167 (N_17167,N_15387,N_14555);
nand U17168 (N_17168,N_14668,N_14280);
xnor U17169 (N_17169,N_15756,N_15733);
and U17170 (N_17170,N_15596,N_14553);
or U17171 (N_17171,N_14026,N_14871);
nand U17172 (N_17172,N_14176,N_14803);
xnor U17173 (N_17173,N_15400,N_15382);
and U17174 (N_17174,N_15902,N_14843);
xnor U17175 (N_17175,N_15040,N_15855);
and U17176 (N_17176,N_15678,N_14999);
nor U17177 (N_17177,N_15795,N_14218);
nand U17178 (N_17178,N_15684,N_15821);
nor U17179 (N_17179,N_14856,N_14535);
nor U17180 (N_17180,N_14006,N_14369);
nand U17181 (N_17181,N_14617,N_15260);
or U17182 (N_17182,N_14397,N_14921);
xor U17183 (N_17183,N_14805,N_14756);
nor U17184 (N_17184,N_14990,N_14060);
or U17185 (N_17185,N_14137,N_15471);
and U17186 (N_17186,N_15312,N_15470);
nor U17187 (N_17187,N_14721,N_14768);
xor U17188 (N_17188,N_14444,N_15682);
and U17189 (N_17189,N_15710,N_14415);
or U17190 (N_17190,N_14938,N_15331);
and U17191 (N_17191,N_15383,N_15672);
nand U17192 (N_17192,N_14433,N_14599);
or U17193 (N_17193,N_14844,N_14329);
and U17194 (N_17194,N_14509,N_14649);
and U17195 (N_17195,N_15614,N_14498);
nand U17196 (N_17196,N_15884,N_15418);
xor U17197 (N_17197,N_15821,N_15955);
or U17198 (N_17198,N_14306,N_15144);
nor U17199 (N_17199,N_14615,N_15820);
xor U17200 (N_17200,N_15507,N_14805);
nor U17201 (N_17201,N_14394,N_15284);
or U17202 (N_17202,N_15454,N_14096);
and U17203 (N_17203,N_14374,N_14980);
or U17204 (N_17204,N_14973,N_15235);
and U17205 (N_17205,N_14170,N_15116);
or U17206 (N_17206,N_14902,N_15713);
nand U17207 (N_17207,N_14528,N_14895);
nand U17208 (N_17208,N_14012,N_15985);
xor U17209 (N_17209,N_15020,N_14545);
nand U17210 (N_17210,N_15365,N_15395);
nand U17211 (N_17211,N_15364,N_14930);
xor U17212 (N_17212,N_15566,N_14530);
nand U17213 (N_17213,N_14962,N_14273);
nor U17214 (N_17214,N_15429,N_14266);
nand U17215 (N_17215,N_14398,N_14765);
xor U17216 (N_17216,N_14060,N_15659);
nor U17217 (N_17217,N_15845,N_14820);
nand U17218 (N_17218,N_15312,N_15023);
xor U17219 (N_17219,N_14036,N_14402);
or U17220 (N_17220,N_15060,N_15594);
and U17221 (N_17221,N_14153,N_15052);
and U17222 (N_17222,N_14507,N_15496);
and U17223 (N_17223,N_15775,N_15308);
nor U17224 (N_17224,N_15278,N_14046);
xnor U17225 (N_17225,N_14721,N_14320);
nor U17226 (N_17226,N_15873,N_15779);
or U17227 (N_17227,N_15372,N_14806);
xnor U17228 (N_17228,N_14223,N_14771);
and U17229 (N_17229,N_15799,N_14165);
nand U17230 (N_17230,N_15425,N_14678);
and U17231 (N_17231,N_14147,N_14202);
nand U17232 (N_17232,N_15339,N_14020);
nand U17233 (N_17233,N_14394,N_14523);
nand U17234 (N_17234,N_14357,N_14791);
or U17235 (N_17235,N_15922,N_15656);
or U17236 (N_17236,N_15655,N_15061);
nor U17237 (N_17237,N_14606,N_14696);
and U17238 (N_17238,N_15305,N_14802);
nand U17239 (N_17239,N_15177,N_14907);
nand U17240 (N_17240,N_14758,N_15564);
and U17241 (N_17241,N_15449,N_15189);
and U17242 (N_17242,N_15140,N_14374);
xor U17243 (N_17243,N_15502,N_14902);
and U17244 (N_17244,N_14321,N_14473);
or U17245 (N_17245,N_15336,N_15917);
xnor U17246 (N_17246,N_14374,N_14604);
and U17247 (N_17247,N_14644,N_14589);
and U17248 (N_17248,N_15418,N_14735);
nand U17249 (N_17249,N_14222,N_15706);
or U17250 (N_17250,N_15471,N_15389);
nor U17251 (N_17251,N_14380,N_15807);
xor U17252 (N_17252,N_14385,N_15233);
nor U17253 (N_17253,N_14378,N_14220);
xnor U17254 (N_17254,N_14400,N_15066);
xor U17255 (N_17255,N_14299,N_14826);
and U17256 (N_17256,N_15653,N_15340);
nor U17257 (N_17257,N_14429,N_15064);
nor U17258 (N_17258,N_15732,N_14583);
or U17259 (N_17259,N_14322,N_14821);
nor U17260 (N_17260,N_14944,N_14743);
xnor U17261 (N_17261,N_15836,N_14935);
and U17262 (N_17262,N_14523,N_14388);
nor U17263 (N_17263,N_14457,N_14978);
and U17264 (N_17264,N_14437,N_15944);
and U17265 (N_17265,N_15700,N_14791);
nor U17266 (N_17266,N_14854,N_15230);
xor U17267 (N_17267,N_14929,N_14905);
nand U17268 (N_17268,N_15630,N_15994);
and U17269 (N_17269,N_15327,N_14938);
and U17270 (N_17270,N_15147,N_15815);
nand U17271 (N_17271,N_14895,N_14514);
xor U17272 (N_17272,N_15952,N_14060);
nor U17273 (N_17273,N_15131,N_15468);
or U17274 (N_17274,N_14097,N_14684);
nand U17275 (N_17275,N_14298,N_14649);
or U17276 (N_17276,N_15803,N_15203);
xnor U17277 (N_17277,N_14912,N_14086);
xnor U17278 (N_17278,N_15534,N_14281);
xnor U17279 (N_17279,N_14328,N_15333);
nand U17280 (N_17280,N_15760,N_15168);
or U17281 (N_17281,N_15525,N_14163);
and U17282 (N_17282,N_14840,N_14582);
nand U17283 (N_17283,N_14942,N_15997);
nor U17284 (N_17284,N_14461,N_14403);
or U17285 (N_17285,N_14444,N_14998);
or U17286 (N_17286,N_14730,N_15455);
nand U17287 (N_17287,N_14467,N_14553);
nor U17288 (N_17288,N_15747,N_14105);
xnor U17289 (N_17289,N_15378,N_15197);
or U17290 (N_17290,N_15335,N_15839);
nor U17291 (N_17291,N_15804,N_14124);
xnor U17292 (N_17292,N_14227,N_14504);
nand U17293 (N_17293,N_15184,N_14515);
or U17294 (N_17294,N_15488,N_14076);
nor U17295 (N_17295,N_14061,N_14737);
or U17296 (N_17296,N_15883,N_15080);
nand U17297 (N_17297,N_15240,N_14914);
and U17298 (N_17298,N_14125,N_14166);
nor U17299 (N_17299,N_15547,N_15469);
and U17300 (N_17300,N_15683,N_15833);
nor U17301 (N_17301,N_14842,N_15378);
xor U17302 (N_17302,N_14015,N_14477);
and U17303 (N_17303,N_15666,N_15306);
nor U17304 (N_17304,N_15532,N_14601);
nand U17305 (N_17305,N_15618,N_14691);
nand U17306 (N_17306,N_14900,N_14990);
nand U17307 (N_17307,N_15884,N_15105);
or U17308 (N_17308,N_14036,N_14410);
nand U17309 (N_17309,N_14106,N_14014);
xor U17310 (N_17310,N_15134,N_15606);
xor U17311 (N_17311,N_15490,N_14581);
xor U17312 (N_17312,N_14634,N_15599);
nand U17313 (N_17313,N_15518,N_15563);
nor U17314 (N_17314,N_15512,N_14400);
nor U17315 (N_17315,N_14518,N_14419);
nand U17316 (N_17316,N_14500,N_14203);
nand U17317 (N_17317,N_15002,N_15463);
nor U17318 (N_17318,N_15558,N_14931);
nor U17319 (N_17319,N_14604,N_14749);
nand U17320 (N_17320,N_14546,N_14972);
nor U17321 (N_17321,N_15892,N_15564);
and U17322 (N_17322,N_15391,N_14747);
or U17323 (N_17323,N_15466,N_15116);
and U17324 (N_17324,N_15132,N_14922);
or U17325 (N_17325,N_15606,N_14188);
nand U17326 (N_17326,N_15301,N_14771);
or U17327 (N_17327,N_14197,N_15547);
nor U17328 (N_17328,N_14859,N_14395);
xnor U17329 (N_17329,N_14861,N_14787);
nand U17330 (N_17330,N_14226,N_15834);
nand U17331 (N_17331,N_15010,N_14731);
xor U17332 (N_17332,N_14647,N_15322);
nand U17333 (N_17333,N_14412,N_15960);
nand U17334 (N_17334,N_15940,N_14988);
nand U17335 (N_17335,N_15027,N_15245);
nor U17336 (N_17336,N_14763,N_14520);
or U17337 (N_17337,N_15301,N_14487);
xnor U17338 (N_17338,N_15815,N_14792);
nand U17339 (N_17339,N_14127,N_14691);
or U17340 (N_17340,N_14563,N_14572);
xnor U17341 (N_17341,N_14233,N_15503);
nor U17342 (N_17342,N_14732,N_15912);
nor U17343 (N_17343,N_15147,N_15481);
nand U17344 (N_17344,N_15902,N_14404);
nor U17345 (N_17345,N_14697,N_15153);
nor U17346 (N_17346,N_14639,N_15339);
nor U17347 (N_17347,N_15612,N_15052);
nor U17348 (N_17348,N_15431,N_14766);
nand U17349 (N_17349,N_15423,N_14048);
or U17350 (N_17350,N_14433,N_15965);
xnor U17351 (N_17351,N_14511,N_15971);
or U17352 (N_17352,N_15294,N_14557);
nor U17353 (N_17353,N_15501,N_15744);
xnor U17354 (N_17354,N_15060,N_15111);
or U17355 (N_17355,N_15557,N_15426);
and U17356 (N_17356,N_15737,N_15036);
xnor U17357 (N_17357,N_15079,N_14711);
or U17358 (N_17358,N_14668,N_14159);
nand U17359 (N_17359,N_15847,N_14358);
or U17360 (N_17360,N_14786,N_14804);
xnor U17361 (N_17361,N_15421,N_14929);
or U17362 (N_17362,N_14760,N_14813);
nand U17363 (N_17363,N_14350,N_14620);
and U17364 (N_17364,N_14960,N_15142);
xnor U17365 (N_17365,N_14562,N_15886);
or U17366 (N_17366,N_14406,N_15734);
and U17367 (N_17367,N_14087,N_15868);
nand U17368 (N_17368,N_15475,N_14508);
or U17369 (N_17369,N_14326,N_15000);
nand U17370 (N_17370,N_15940,N_15639);
nor U17371 (N_17371,N_15067,N_14258);
nand U17372 (N_17372,N_15317,N_15055);
nand U17373 (N_17373,N_14887,N_15807);
or U17374 (N_17374,N_15003,N_15659);
or U17375 (N_17375,N_14518,N_14583);
nand U17376 (N_17376,N_15142,N_14183);
and U17377 (N_17377,N_15737,N_14255);
and U17378 (N_17378,N_15484,N_14182);
or U17379 (N_17379,N_15604,N_15134);
xnor U17380 (N_17380,N_15035,N_14645);
nand U17381 (N_17381,N_14723,N_15403);
and U17382 (N_17382,N_14147,N_14004);
and U17383 (N_17383,N_14350,N_14824);
or U17384 (N_17384,N_14580,N_15923);
xor U17385 (N_17385,N_14843,N_15612);
nor U17386 (N_17386,N_15571,N_14553);
or U17387 (N_17387,N_15366,N_14407);
nand U17388 (N_17388,N_14417,N_14176);
and U17389 (N_17389,N_14888,N_15113);
and U17390 (N_17390,N_14309,N_15586);
nand U17391 (N_17391,N_14319,N_15147);
xnor U17392 (N_17392,N_15938,N_14259);
and U17393 (N_17393,N_14374,N_14051);
or U17394 (N_17394,N_14863,N_15052);
nand U17395 (N_17395,N_15405,N_15437);
xor U17396 (N_17396,N_14790,N_14088);
xor U17397 (N_17397,N_14159,N_14561);
nand U17398 (N_17398,N_15886,N_14295);
nor U17399 (N_17399,N_14029,N_14287);
nand U17400 (N_17400,N_15427,N_14832);
and U17401 (N_17401,N_14483,N_14676);
or U17402 (N_17402,N_15204,N_15797);
nor U17403 (N_17403,N_15863,N_14389);
and U17404 (N_17404,N_14510,N_14671);
or U17405 (N_17405,N_15064,N_14002);
nor U17406 (N_17406,N_14245,N_14090);
or U17407 (N_17407,N_15593,N_14821);
or U17408 (N_17408,N_15982,N_14925);
or U17409 (N_17409,N_14043,N_14446);
xnor U17410 (N_17410,N_15017,N_14266);
nand U17411 (N_17411,N_14755,N_15426);
nor U17412 (N_17412,N_15297,N_14683);
nand U17413 (N_17413,N_14335,N_14523);
or U17414 (N_17414,N_15341,N_15095);
nand U17415 (N_17415,N_15987,N_15690);
xor U17416 (N_17416,N_15400,N_14301);
nand U17417 (N_17417,N_14670,N_14277);
xor U17418 (N_17418,N_14867,N_15232);
xnor U17419 (N_17419,N_14054,N_14911);
nand U17420 (N_17420,N_14478,N_14252);
or U17421 (N_17421,N_15532,N_15974);
and U17422 (N_17422,N_15111,N_14386);
or U17423 (N_17423,N_14488,N_15185);
xor U17424 (N_17424,N_15048,N_14716);
or U17425 (N_17425,N_14009,N_14203);
or U17426 (N_17426,N_14279,N_15271);
xnor U17427 (N_17427,N_14629,N_14524);
and U17428 (N_17428,N_15702,N_14955);
and U17429 (N_17429,N_14766,N_15039);
nor U17430 (N_17430,N_14834,N_15884);
nand U17431 (N_17431,N_15499,N_15550);
nand U17432 (N_17432,N_15821,N_15978);
xor U17433 (N_17433,N_15058,N_15503);
xnor U17434 (N_17434,N_15781,N_15946);
or U17435 (N_17435,N_14764,N_15987);
nand U17436 (N_17436,N_14143,N_14921);
xor U17437 (N_17437,N_15285,N_14859);
nand U17438 (N_17438,N_14012,N_15434);
nor U17439 (N_17439,N_14799,N_15939);
xor U17440 (N_17440,N_15092,N_15872);
nor U17441 (N_17441,N_15742,N_14036);
nand U17442 (N_17442,N_14702,N_14565);
or U17443 (N_17443,N_15410,N_14622);
nand U17444 (N_17444,N_14988,N_14725);
and U17445 (N_17445,N_14235,N_15676);
nand U17446 (N_17446,N_14670,N_15041);
xor U17447 (N_17447,N_14361,N_14622);
xor U17448 (N_17448,N_15399,N_14162);
or U17449 (N_17449,N_14794,N_14050);
nor U17450 (N_17450,N_15099,N_14911);
nor U17451 (N_17451,N_15149,N_15673);
xor U17452 (N_17452,N_15259,N_14510);
and U17453 (N_17453,N_14631,N_14973);
and U17454 (N_17454,N_15624,N_15922);
xnor U17455 (N_17455,N_14319,N_14864);
nand U17456 (N_17456,N_14843,N_15424);
or U17457 (N_17457,N_15510,N_15461);
nor U17458 (N_17458,N_14197,N_15070);
and U17459 (N_17459,N_15917,N_15087);
xnor U17460 (N_17460,N_14784,N_14484);
xor U17461 (N_17461,N_15346,N_14234);
nand U17462 (N_17462,N_15728,N_14669);
or U17463 (N_17463,N_15909,N_15279);
or U17464 (N_17464,N_14666,N_14564);
and U17465 (N_17465,N_14546,N_14732);
nand U17466 (N_17466,N_15126,N_14362);
and U17467 (N_17467,N_14780,N_15462);
and U17468 (N_17468,N_14998,N_14551);
nand U17469 (N_17469,N_15248,N_15671);
and U17470 (N_17470,N_14221,N_14313);
nor U17471 (N_17471,N_15248,N_15933);
or U17472 (N_17472,N_14519,N_15898);
or U17473 (N_17473,N_15138,N_15404);
or U17474 (N_17474,N_15097,N_15790);
or U17475 (N_17475,N_14658,N_15330);
or U17476 (N_17476,N_14270,N_15092);
xnor U17477 (N_17477,N_14705,N_14863);
xnor U17478 (N_17478,N_15045,N_15078);
nand U17479 (N_17479,N_14943,N_14937);
nor U17480 (N_17480,N_15028,N_15216);
xor U17481 (N_17481,N_15288,N_15125);
nand U17482 (N_17482,N_14237,N_15256);
or U17483 (N_17483,N_15727,N_15945);
nand U17484 (N_17484,N_15981,N_14509);
nand U17485 (N_17485,N_14085,N_15778);
nor U17486 (N_17486,N_14187,N_15355);
nor U17487 (N_17487,N_15662,N_14500);
nand U17488 (N_17488,N_14209,N_14697);
or U17489 (N_17489,N_14386,N_14719);
and U17490 (N_17490,N_15022,N_14919);
nor U17491 (N_17491,N_14453,N_14053);
nor U17492 (N_17492,N_15199,N_14050);
xor U17493 (N_17493,N_14421,N_15711);
or U17494 (N_17494,N_15901,N_15759);
nor U17495 (N_17495,N_14251,N_14835);
nor U17496 (N_17496,N_15283,N_14405);
nand U17497 (N_17497,N_14416,N_14338);
or U17498 (N_17498,N_15126,N_15137);
xor U17499 (N_17499,N_15463,N_15833);
nand U17500 (N_17500,N_14069,N_15165);
nand U17501 (N_17501,N_15466,N_15800);
and U17502 (N_17502,N_14848,N_15660);
and U17503 (N_17503,N_14304,N_14851);
and U17504 (N_17504,N_15626,N_14609);
nand U17505 (N_17505,N_14072,N_15526);
nand U17506 (N_17506,N_15732,N_14766);
xor U17507 (N_17507,N_14948,N_14339);
nand U17508 (N_17508,N_14925,N_14753);
and U17509 (N_17509,N_14795,N_15485);
xnor U17510 (N_17510,N_14214,N_14161);
nor U17511 (N_17511,N_15685,N_14142);
or U17512 (N_17512,N_15327,N_14509);
or U17513 (N_17513,N_15338,N_15636);
xnor U17514 (N_17514,N_15756,N_14015);
or U17515 (N_17515,N_15391,N_15821);
nand U17516 (N_17516,N_14715,N_15315);
nor U17517 (N_17517,N_15004,N_14719);
and U17518 (N_17518,N_14329,N_14593);
xnor U17519 (N_17519,N_15019,N_14764);
xor U17520 (N_17520,N_15965,N_14964);
nor U17521 (N_17521,N_15411,N_15346);
and U17522 (N_17522,N_14907,N_15672);
nor U17523 (N_17523,N_15649,N_15026);
or U17524 (N_17524,N_14648,N_15421);
nand U17525 (N_17525,N_15493,N_14522);
xnor U17526 (N_17526,N_15423,N_15769);
nor U17527 (N_17527,N_15037,N_14182);
nand U17528 (N_17528,N_15289,N_14524);
and U17529 (N_17529,N_15842,N_14545);
nand U17530 (N_17530,N_14756,N_14990);
xnor U17531 (N_17531,N_14758,N_14876);
xor U17532 (N_17532,N_14455,N_14452);
xnor U17533 (N_17533,N_15062,N_15888);
nor U17534 (N_17534,N_14277,N_14053);
xor U17535 (N_17535,N_14240,N_15295);
and U17536 (N_17536,N_15583,N_14607);
nor U17537 (N_17537,N_14897,N_14138);
xnor U17538 (N_17538,N_14723,N_14146);
and U17539 (N_17539,N_14466,N_15189);
xor U17540 (N_17540,N_14743,N_15969);
and U17541 (N_17541,N_14775,N_15330);
xnor U17542 (N_17542,N_15612,N_14898);
and U17543 (N_17543,N_15484,N_15597);
and U17544 (N_17544,N_15342,N_15897);
or U17545 (N_17545,N_15569,N_15749);
nand U17546 (N_17546,N_15119,N_15274);
nor U17547 (N_17547,N_15713,N_15522);
and U17548 (N_17548,N_14156,N_15655);
nand U17549 (N_17549,N_14348,N_15370);
or U17550 (N_17550,N_15022,N_14893);
xor U17551 (N_17551,N_15935,N_14969);
xnor U17552 (N_17552,N_14910,N_15877);
nor U17553 (N_17553,N_14205,N_15235);
and U17554 (N_17554,N_15180,N_14548);
or U17555 (N_17555,N_14590,N_14377);
nor U17556 (N_17556,N_15804,N_15316);
nor U17557 (N_17557,N_14350,N_14924);
nor U17558 (N_17558,N_14638,N_15603);
nand U17559 (N_17559,N_14988,N_14996);
nand U17560 (N_17560,N_14971,N_14203);
nor U17561 (N_17561,N_14550,N_15676);
and U17562 (N_17562,N_14788,N_14192);
or U17563 (N_17563,N_15158,N_14830);
nor U17564 (N_17564,N_15951,N_15741);
nand U17565 (N_17565,N_14086,N_14183);
or U17566 (N_17566,N_15443,N_15788);
nand U17567 (N_17567,N_14592,N_15232);
or U17568 (N_17568,N_15907,N_14551);
and U17569 (N_17569,N_14227,N_14524);
nor U17570 (N_17570,N_15831,N_14643);
or U17571 (N_17571,N_15958,N_15479);
xor U17572 (N_17572,N_14290,N_15006);
or U17573 (N_17573,N_14524,N_15679);
nand U17574 (N_17574,N_15464,N_15919);
and U17575 (N_17575,N_14579,N_14809);
nand U17576 (N_17576,N_15002,N_14818);
xor U17577 (N_17577,N_15430,N_14983);
xnor U17578 (N_17578,N_14316,N_15786);
xnor U17579 (N_17579,N_14038,N_15377);
nand U17580 (N_17580,N_14293,N_14778);
or U17581 (N_17581,N_14534,N_14790);
xor U17582 (N_17582,N_15562,N_15916);
and U17583 (N_17583,N_15065,N_15017);
and U17584 (N_17584,N_15530,N_15216);
and U17585 (N_17585,N_15023,N_15622);
xnor U17586 (N_17586,N_15924,N_14376);
xnor U17587 (N_17587,N_14910,N_14523);
xor U17588 (N_17588,N_14447,N_15851);
nand U17589 (N_17589,N_15711,N_15177);
nand U17590 (N_17590,N_15060,N_14478);
xor U17591 (N_17591,N_14798,N_15948);
nor U17592 (N_17592,N_15968,N_14240);
xnor U17593 (N_17593,N_14929,N_15196);
and U17594 (N_17594,N_15652,N_14377);
xor U17595 (N_17595,N_15527,N_15668);
and U17596 (N_17596,N_15068,N_15276);
and U17597 (N_17597,N_14199,N_15977);
and U17598 (N_17598,N_14229,N_15841);
nand U17599 (N_17599,N_15101,N_14791);
or U17600 (N_17600,N_14378,N_15897);
xnor U17601 (N_17601,N_15101,N_15988);
or U17602 (N_17602,N_14779,N_14802);
nand U17603 (N_17603,N_14767,N_14206);
xor U17604 (N_17604,N_15812,N_15196);
nor U17605 (N_17605,N_15611,N_14929);
nor U17606 (N_17606,N_14740,N_14964);
xor U17607 (N_17607,N_15071,N_15800);
and U17608 (N_17608,N_15247,N_15331);
xnor U17609 (N_17609,N_14419,N_14631);
nor U17610 (N_17610,N_15799,N_15098);
xor U17611 (N_17611,N_15728,N_15507);
and U17612 (N_17612,N_15111,N_14344);
nand U17613 (N_17613,N_14344,N_14153);
nor U17614 (N_17614,N_14480,N_15509);
nor U17615 (N_17615,N_14318,N_14130);
nor U17616 (N_17616,N_14606,N_15276);
and U17617 (N_17617,N_14555,N_14150);
and U17618 (N_17618,N_15740,N_15663);
nand U17619 (N_17619,N_14280,N_15912);
or U17620 (N_17620,N_14118,N_15182);
xor U17621 (N_17621,N_15999,N_14451);
nand U17622 (N_17622,N_14988,N_15490);
and U17623 (N_17623,N_14902,N_15153);
nand U17624 (N_17624,N_15619,N_14416);
or U17625 (N_17625,N_14388,N_15577);
nand U17626 (N_17626,N_15324,N_14658);
nand U17627 (N_17627,N_14786,N_15676);
or U17628 (N_17628,N_14964,N_14876);
or U17629 (N_17629,N_14937,N_14970);
nor U17630 (N_17630,N_15501,N_14053);
nor U17631 (N_17631,N_14856,N_15109);
nor U17632 (N_17632,N_15297,N_15614);
or U17633 (N_17633,N_14014,N_15783);
or U17634 (N_17634,N_14429,N_14500);
and U17635 (N_17635,N_15345,N_15354);
xor U17636 (N_17636,N_15538,N_15509);
and U17637 (N_17637,N_15618,N_15934);
nor U17638 (N_17638,N_15241,N_15181);
xor U17639 (N_17639,N_15783,N_15606);
nand U17640 (N_17640,N_15426,N_15019);
and U17641 (N_17641,N_14227,N_15981);
and U17642 (N_17642,N_15276,N_14110);
nor U17643 (N_17643,N_14153,N_15832);
xor U17644 (N_17644,N_15942,N_15182);
xor U17645 (N_17645,N_15014,N_14363);
xor U17646 (N_17646,N_14954,N_14502);
and U17647 (N_17647,N_14240,N_15175);
xnor U17648 (N_17648,N_15373,N_14361);
nor U17649 (N_17649,N_15409,N_15853);
and U17650 (N_17650,N_15235,N_15412);
nand U17651 (N_17651,N_15641,N_15914);
nor U17652 (N_17652,N_15382,N_14497);
or U17653 (N_17653,N_14668,N_15388);
nand U17654 (N_17654,N_14436,N_15283);
xnor U17655 (N_17655,N_14377,N_15989);
and U17656 (N_17656,N_14668,N_14579);
nand U17657 (N_17657,N_14910,N_15092);
and U17658 (N_17658,N_14089,N_14035);
nor U17659 (N_17659,N_14901,N_14292);
nor U17660 (N_17660,N_15255,N_14208);
or U17661 (N_17661,N_15587,N_15614);
or U17662 (N_17662,N_15244,N_14619);
or U17663 (N_17663,N_15656,N_15652);
nand U17664 (N_17664,N_15334,N_15042);
and U17665 (N_17665,N_15736,N_14256);
and U17666 (N_17666,N_14268,N_15175);
and U17667 (N_17667,N_15359,N_14715);
and U17668 (N_17668,N_15531,N_14186);
nand U17669 (N_17669,N_15480,N_15055);
nand U17670 (N_17670,N_15154,N_14639);
xnor U17671 (N_17671,N_15337,N_15301);
and U17672 (N_17672,N_14775,N_15185);
and U17673 (N_17673,N_15021,N_14163);
or U17674 (N_17674,N_14136,N_14924);
or U17675 (N_17675,N_14075,N_14210);
and U17676 (N_17676,N_14979,N_14190);
or U17677 (N_17677,N_15928,N_15825);
xor U17678 (N_17678,N_15721,N_15714);
xor U17679 (N_17679,N_15866,N_14822);
nor U17680 (N_17680,N_15876,N_14768);
xor U17681 (N_17681,N_14939,N_14779);
or U17682 (N_17682,N_15363,N_14864);
xnor U17683 (N_17683,N_14092,N_14796);
xor U17684 (N_17684,N_14059,N_15727);
xnor U17685 (N_17685,N_15840,N_15220);
xor U17686 (N_17686,N_14993,N_14699);
xor U17687 (N_17687,N_15544,N_14822);
nand U17688 (N_17688,N_14733,N_14230);
and U17689 (N_17689,N_14270,N_15513);
nor U17690 (N_17690,N_15103,N_14472);
nand U17691 (N_17691,N_15269,N_15176);
and U17692 (N_17692,N_15519,N_15712);
xnor U17693 (N_17693,N_15728,N_15279);
xor U17694 (N_17694,N_14455,N_15642);
nor U17695 (N_17695,N_14559,N_14242);
and U17696 (N_17696,N_15038,N_15767);
nand U17697 (N_17697,N_15447,N_15900);
nor U17698 (N_17698,N_15129,N_15935);
nor U17699 (N_17699,N_15478,N_14837);
nor U17700 (N_17700,N_14470,N_15642);
or U17701 (N_17701,N_14879,N_15477);
nor U17702 (N_17702,N_15192,N_14196);
nand U17703 (N_17703,N_15175,N_15955);
nor U17704 (N_17704,N_14206,N_15753);
nor U17705 (N_17705,N_15083,N_14284);
or U17706 (N_17706,N_14182,N_15144);
nand U17707 (N_17707,N_15842,N_15137);
and U17708 (N_17708,N_15568,N_15139);
and U17709 (N_17709,N_15579,N_15090);
and U17710 (N_17710,N_14877,N_15641);
xnor U17711 (N_17711,N_15404,N_15466);
nand U17712 (N_17712,N_15485,N_15752);
and U17713 (N_17713,N_15018,N_15784);
or U17714 (N_17714,N_14298,N_14149);
or U17715 (N_17715,N_15614,N_14980);
nor U17716 (N_17716,N_15001,N_15256);
nand U17717 (N_17717,N_14878,N_14844);
or U17718 (N_17718,N_15461,N_14760);
nand U17719 (N_17719,N_14737,N_14664);
or U17720 (N_17720,N_15305,N_14305);
xnor U17721 (N_17721,N_15125,N_14783);
nor U17722 (N_17722,N_15454,N_15239);
nor U17723 (N_17723,N_15254,N_14636);
nand U17724 (N_17724,N_15385,N_14053);
xor U17725 (N_17725,N_15936,N_14906);
and U17726 (N_17726,N_15545,N_15728);
nand U17727 (N_17727,N_14013,N_14038);
xor U17728 (N_17728,N_14900,N_15446);
nor U17729 (N_17729,N_14760,N_15571);
xor U17730 (N_17730,N_14004,N_14746);
nor U17731 (N_17731,N_14675,N_15064);
nor U17732 (N_17732,N_14161,N_14429);
and U17733 (N_17733,N_15983,N_15008);
or U17734 (N_17734,N_15308,N_14441);
nor U17735 (N_17735,N_15747,N_15037);
or U17736 (N_17736,N_15560,N_14021);
nor U17737 (N_17737,N_14726,N_15748);
xor U17738 (N_17738,N_14949,N_15881);
and U17739 (N_17739,N_14887,N_15518);
and U17740 (N_17740,N_14918,N_14451);
and U17741 (N_17741,N_14674,N_14876);
nor U17742 (N_17742,N_15087,N_14476);
nor U17743 (N_17743,N_14760,N_15747);
nor U17744 (N_17744,N_14564,N_15376);
and U17745 (N_17745,N_15420,N_15215);
nand U17746 (N_17746,N_14490,N_15603);
nor U17747 (N_17747,N_14143,N_15488);
and U17748 (N_17748,N_14424,N_15556);
or U17749 (N_17749,N_15773,N_15195);
xnor U17750 (N_17750,N_14640,N_14509);
or U17751 (N_17751,N_15864,N_14354);
or U17752 (N_17752,N_15983,N_14471);
nand U17753 (N_17753,N_15129,N_15379);
and U17754 (N_17754,N_14218,N_14916);
and U17755 (N_17755,N_15867,N_14971);
xnor U17756 (N_17756,N_15359,N_14378);
nand U17757 (N_17757,N_15808,N_15185);
nand U17758 (N_17758,N_14762,N_14159);
xor U17759 (N_17759,N_15898,N_15807);
and U17760 (N_17760,N_14704,N_15616);
nand U17761 (N_17761,N_15178,N_14278);
xnor U17762 (N_17762,N_14228,N_14789);
or U17763 (N_17763,N_14087,N_14767);
nor U17764 (N_17764,N_15710,N_15862);
nor U17765 (N_17765,N_15768,N_14587);
xor U17766 (N_17766,N_14188,N_15118);
and U17767 (N_17767,N_14415,N_14810);
and U17768 (N_17768,N_15445,N_14285);
nand U17769 (N_17769,N_15298,N_14122);
nand U17770 (N_17770,N_15730,N_15741);
xnor U17771 (N_17771,N_14129,N_15412);
nand U17772 (N_17772,N_15283,N_14662);
and U17773 (N_17773,N_15958,N_15583);
or U17774 (N_17774,N_15988,N_14936);
nand U17775 (N_17775,N_15391,N_14958);
and U17776 (N_17776,N_14648,N_15653);
nor U17777 (N_17777,N_14130,N_15478);
and U17778 (N_17778,N_15490,N_14917);
xor U17779 (N_17779,N_15581,N_14508);
xnor U17780 (N_17780,N_15559,N_14381);
nand U17781 (N_17781,N_14556,N_14544);
and U17782 (N_17782,N_14385,N_15177);
and U17783 (N_17783,N_14478,N_14366);
nor U17784 (N_17784,N_15427,N_14733);
xor U17785 (N_17785,N_14757,N_15307);
nand U17786 (N_17786,N_14328,N_14991);
and U17787 (N_17787,N_14351,N_15168);
and U17788 (N_17788,N_15518,N_15924);
nor U17789 (N_17789,N_15616,N_14325);
xor U17790 (N_17790,N_15453,N_14721);
or U17791 (N_17791,N_15441,N_14890);
or U17792 (N_17792,N_14860,N_14126);
nand U17793 (N_17793,N_15580,N_15664);
nand U17794 (N_17794,N_14181,N_15933);
xnor U17795 (N_17795,N_14089,N_15469);
or U17796 (N_17796,N_14958,N_15508);
or U17797 (N_17797,N_15909,N_15549);
xor U17798 (N_17798,N_15825,N_14765);
nand U17799 (N_17799,N_15198,N_15933);
or U17800 (N_17800,N_15214,N_15077);
nor U17801 (N_17801,N_15860,N_15382);
or U17802 (N_17802,N_14624,N_15763);
xor U17803 (N_17803,N_14849,N_14869);
xnor U17804 (N_17804,N_14101,N_15012);
or U17805 (N_17805,N_14577,N_15749);
xnor U17806 (N_17806,N_15028,N_14381);
or U17807 (N_17807,N_15196,N_15503);
xnor U17808 (N_17808,N_14591,N_15331);
and U17809 (N_17809,N_14680,N_15828);
xnor U17810 (N_17810,N_15528,N_15809);
or U17811 (N_17811,N_15384,N_15289);
nor U17812 (N_17812,N_14823,N_15290);
or U17813 (N_17813,N_14532,N_15946);
and U17814 (N_17814,N_14492,N_14091);
and U17815 (N_17815,N_15909,N_14670);
and U17816 (N_17816,N_14584,N_14751);
or U17817 (N_17817,N_14178,N_15107);
nor U17818 (N_17818,N_14095,N_15691);
and U17819 (N_17819,N_15973,N_15581);
nand U17820 (N_17820,N_14527,N_14479);
nor U17821 (N_17821,N_14292,N_15408);
or U17822 (N_17822,N_14287,N_14128);
nor U17823 (N_17823,N_15995,N_15313);
and U17824 (N_17824,N_14063,N_15767);
nor U17825 (N_17825,N_14720,N_15294);
or U17826 (N_17826,N_14224,N_15564);
nor U17827 (N_17827,N_14421,N_14470);
nand U17828 (N_17828,N_14981,N_14005);
nand U17829 (N_17829,N_14698,N_14799);
nand U17830 (N_17830,N_15413,N_14139);
nor U17831 (N_17831,N_15456,N_14383);
or U17832 (N_17832,N_14653,N_15061);
nor U17833 (N_17833,N_15771,N_14508);
and U17834 (N_17834,N_15485,N_15098);
nand U17835 (N_17835,N_15832,N_15488);
nand U17836 (N_17836,N_14278,N_14346);
nor U17837 (N_17837,N_14191,N_15586);
and U17838 (N_17838,N_14676,N_14089);
or U17839 (N_17839,N_14899,N_14854);
or U17840 (N_17840,N_14946,N_15541);
and U17841 (N_17841,N_14093,N_15022);
xnor U17842 (N_17842,N_14682,N_14398);
or U17843 (N_17843,N_15408,N_15836);
and U17844 (N_17844,N_14823,N_15363);
and U17845 (N_17845,N_14941,N_15611);
nor U17846 (N_17846,N_15464,N_15812);
nor U17847 (N_17847,N_14675,N_15821);
xor U17848 (N_17848,N_15125,N_15469);
xor U17849 (N_17849,N_15799,N_14386);
nand U17850 (N_17850,N_15730,N_15908);
nor U17851 (N_17851,N_14391,N_15343);
and U17852 (N_17852,N_14365,N_15220);
nor U17853 (N_17853,N_14146,N_14582);
nand U17854 (N_17854,N_15269,N_15156);
nor U17855 (N_17855,N_15764,N_14150);
nand U17856 (N_17856,N_14801,N_14326);
xor U17857 (N_17857,N_14847,N_14897);
or U17858 (N_17858,N_15582,N_15665);
and U17859 (N_17859,N_14151,N_15691);
and U17860 (N_17860,N_15415,N_15798);
nand U17861 (N_17861,N_15690,N_15810);
and U17862 (N_17862,N_15909,N_15478);
nand U17863 (N_17863,N_15234,N_15348);
nor U17864 (N_17864,N_14948,N_15199);
and U17865 (N_17865,N_14916,N_15845);
nand U17866 (N_17866,N_14262,N_14942);
xor U17867 (N_17867,N_14271,N_14632);
and U17868 (N_17868,N_15071,N_15094);
nand U17869 (N_17869,N_14258,N_15213);
or U17870 (N_17870,N_15373,N_15930);
and U17871 (N_17871,N_15280,N_14239);
or U17872 (N_17872,N_15607,N_15140);
and U17873 (N_17873,N_15359,N_14954);
xor U17874 (N_17874,N_14251,N_14791);
and U17875 (N_17875,N_15181,N_14946);
nand U17876 (N_17876,N_14920,N_14622);
and U17877 (N_17877,N_14755,N_15398);
nor U17878 (N_17878,N_14681,N_15028);
nor U17879 (N_17879,N_15883,N_14917);
or U17880 (N_17880,N_15789,N_15458);
and U17881 (N_17881,N_15026,N_14980);
nor U17882 (N_17882,N_14282,N_14708);
xor U17883 (N_17883,N_14203,N_15580);
or U17884 (N_17884,N_15009,N_15077);
nor U17885 (N_17885,N_15998,N_15293);
nand U17886 (N_17886,N_15398,N_14390);
or U17887 (N_17887,N_14247,N_14022);
xor U17888 (N_17888,N_15795,N_14885);
nand U17889 (N_17889,N_14460,N_15041);
or U17890 (N_17890,N_15668,N_15122);
or U17891 (N_17891,N_15578,N_14534);
or U17892 (N_17892,N_15159,N_14757);
or U17893 (N_17893,N_14432,N_15853);
nor U17894 (N_17894,N_14766,N_15129);
nand U17895 (N_17895,N_15328,N_15640);
and U17896 (N_17896,N_15100,N_15602);
and U17897 (N_17897,N_14342,N_15517);
xnor U17898 (N_17898,N_14618,N_14998);
xnor U17899 (N_17899,N_15491,N_14722);
and U17900 (N_17900,N_14627,N_15274);
and U17901 (N_17901,N_15266,N_14486);
nand U17902 (N_17902,N_14994,N_14518);
and U17903 (N_17903,N_15624,N_15265);
xor U17904 (N_17904,N_15981,N_15674);
or U17905 (N_17905,N_15761,N_14020);
xor U17906 (N_17906,N_15855,N_15565);
or U17907 (N_17907,N_15044,N_15335);
nand U17908 (N_17908,N_14913,N_15542);
nand U17909 (N_17909,N_14549,N_15627);
or U17910 (N_17910,N_15946,N_14719);
xor U17911 (N_17911,N_14955,N_14833);
xor U17912 (N_17912,N_14008,N_15927);
nor U17913 (N_17913,N_14321,N_15124);
xor U17914 (N_17914,N_14880,N_14130);
nand U17915 (N_17915,N_15826,N_14023);
nand U17916 (N_17916,N_14447,N_14703);
nor U17917 (N_17917,N_14901,N_15780);
and U17918 (N_17918,N_15428,N_15274);
nor U17919 (N_17919,N_15810,N_14384);
xnor U17920 (N_17920,N_15655,N_14512);
xnor U17921 (N_17921,N_14080,N_14382);
nand U17922 (N_17922,N_14466,N_15611);
xnor U17923 (N_17923,N_15552,N_14371);
nor U17924 (N_17924,N_14073,N_14841);
and U17925 (N_17925,N_14540,N_14917);
and U17926 (N_17926,N_14886,N_14018);
or U17927 (N_17927,N_14879,N_14822);
or U17928 (N_17928,N_14043,N_15108);
xnor U17929 (N_17929,N_15554,N_14540);
xor U17930 (N_17930,N_15758,N_14763);
nand U17931 (N_17931,N_15522,N_15975);
or U17932 (N_17932,N_15387,N_14500);
nor U17933 (N_17933,N_14551,N_14575);
xnor U17934 (N_17934,N_15235,N_14901);
or U17935 (N_17935,N_14495,N_15835);
xnor U17936 (N_17936,N_15284,N_15903);
and U17937 (N_17937,N_14372,N_14943);
and U17938 (N_17938,N_14466,N_15771);
and U17939 (N_17939,N_15210,N_14635);
nand U17940 (N_17940,N_15995,N_14041);
xor U17941 (N_17941,N_15717,N_14150);
or U17942 (N_17942,N_15277,N_15978);
nand U17943 (N_17943,N_14955,N_14315);
nand U17944 (N_17944,N_14320,N_15816);
and U17945 (N_17945,N_14071,N_14612);
or U17946 (N_17946,N_14490,N_15659);
nand U17947 (N_17947,N_14376,N_15340);
or U17948 (N_17948,N_15447,N_14375);
or U17949 (N_17949,N_15869,N_14953);
xnor U17950 (N_17950,N_14402,N_15218);
nand U17951 (N_17951,N_15914,N_14611);
and U17952 (N_17952,N_14482,N_14667);
nor U17953 (N_17953,N_14106,N_14203);
nor U17954 (N_17954,N_14715,N_15629);
and U17955 (N_17955,N_15258,N_15912);
xor U17956 (N_17956,N_14101,N_15585);
nand U17957 (N_17957,N_14875,N_14799);
nor U17958 (N_17958,N_14404,N_15814);
nor U17959 (N_17959,N_15786,N_14663);
nand U17960 (N_17960,N_15232,N_14263);
and U17961 (N_17961,N_14862,N_14904);
and U17962 (N_17962,N_15001,N_14856);
nor U17963 (N_17963,N_15716,N_14108);
xnor U17964 (N_17964,N_15525,N_15839);
and U17965 (N_17965,N_15338,N_14515);
or U17966 (N_17966,N_14399,N_15171);
nor U17967 (N_17967,N_14792,N_15387);
and U17968 (N_17968,N_14377,N_14977);
or U17969 (N_17969,N_14530,N_15804);
xor U17970 (N_17970,N_15158,N_14290);
and U17971 (N_17971,N_15859,N_14131);
nor U17972 (N_17972,N_14437,N_14346);
or U17973 (N_17973,N_15996,N_14658);
and U17974 (N_17974,N_15667,N_14780);
nand U17975 (N_17975,N_15953,N_15464);
and U17976 (N_17976,N_15568,N_14154);
xnor U17977 (N_17977,N_15410,N_14288);
nand U17978 (N_17978,N_15379,N_15438);
xor U17979 (N_17979,N_14283,N_14081);
or U17980 (N_17980,N_15264,N_14629);
nor U17981 (N_17981,N_15845,N_15467);
or U17982 (N_17982,N_14797,N_15431);
nor U17983 (N_17983,N_14865,N_14295);
nor U17984 (N_17984,N_15762,N_14368);
xor U17985 (N_17985,N_14505,N_15713);
xnor U17986 (N_17986,N_14071,N_15601);
nor U17987 (N_17987,N_15998,N_15620);
and U17988 (N_17988,N_15587,N_15799);
xnor U17989 (N_17989,N_15832,N_15391);
nand U17990 (N_17990,N_14018,N_14424);
nor U17991 (N_17991,N_15011,N_14188);
xnor U17992 (N_17992,N_14269,N_15987);
nand U17993 (N_17993,N_14994,N_14707);
nor U17994 (N_17994,N_14046,N_14621);
or U17995 (N_17995,N_15955,N_14971);
and U17996 (N_17996,N_15167,N_14247);
xnor U17997 (N_17997,N_15999,N_15346);
nand U17998 (N_17998,N_15894,N_15202);
nand U17999 (N_17999,N_14271,N_15779);
or U18000 (N_18000,N_17754,N_17422);
xnor U18001 (N_18001,N_16221,N_16673);
xnor U18002 (N_18002,N_16217,N_17606);
and U18003 (N_18003,N_16632,N_16480);
nand U18004 (N_18004,N_16824,N_17161);
nor U18005 (N_18005,N_16404,N_16297);
or U18006 (N_18006,N_17016,N_16934);
xnor U18007 (N_18007,N_16285,N_16823);
or U18008 (N_18008,N_16324,N_16128);
and U18009 (N_18009,N_17572,N_16112);
nor U18010 (N_18010,N_16138,N_16422);
and U18011 (N_18011,N_17830,N_17586);
or U18012 (N_18012,N_16930,N_16062);
xor U18013 (N_18013,N_17323,N_16765);
or U18014 (N_18014,N_16931,N_16603);
xnor U18015 (N_18015,N_16838,N_16118);
xnor U18016 (N_18016,N_17827,N_16518);
or U18017 (N_18017,N_16047,N_16644);
or U18018 (N_18018,N_16107,N_16362);
nand U18019 (N_18019,N_16883,N_16859);
and U18020 (N_18020,N_17976,N_16901);
and U18021 (N_18021,N_16148,N_16431);
nand U18022 (N_18022,N_16952,N_17130);
nor U18023 (N_18023,N_17887,N_17461);
nor U18024 (N_18024,N_17185,N_17256);
nor U18025 (N_18025,N_16638,N_16448);
and U18026 (N_18026,N_17675,N_16831);
nor U18027 (N_18027,N_17479,N_16164);
nand U18028 (N_18028,N_17408,N_17287);
and U18029 (N_18029,N_16271,N_16872);
xor U18030 (N_18030,N_17707,N_17747);
or U18031 (N_18031,N_16977,N_16668);
nand U18032 (N_18032,N_16794,N_17162);
nor U18033 (N_18033,N_17147,N_17796);
nor U18034 (N_18034,N_16911,N_17312);
or U18035 (N_18035,N_16007,N_16861);
nor U18036 (N_18036,N_17493,N_17954);
and U18037 (N_18037,N_16569,N_17849);
nand U18038 (N_18038,N_17218,N_17184);
nor U18039 (N_18039,N_16142,N_17038);
or U18040 (N_18040,N_17496,N_17415);
or U18041 (N_18041,N_17427,N_17335);
nor U18042 (N_18042,N_17180,N_16230);
or U18043 (N_18043,N_16447,N_16593);
nor U18044 (N_18044,N_17265,N_16833);
nand U18045 (N_18045,N_16388,N_16174);
or U18046 (N_18046,N_16200,N_17610);
xor U18047 (N_18047,N_17376,N_16209);
and U18048 (N_18048,N_16167,N_16568);
nand U18049 (N_18049,N_16249,N_17640);
and U18050 (N_18050,N_16320,N_16332);
nand U18051 (N_18051,N_17968,N_16845);
and U18052 (N_18052,N_16081,N_17979);
nand U18053 (N_18053,N_16565,N_16598);
or U18054 (N_18054,N_17800,N_17398);
nand U18055 (N_18055,N_16897,N_16982);
and U18056 (N_18056,N_17739,N_16359);
nand U18057 (N_18057,N_17146,N_17542);
or U18058 (N_18058,N_16922,N_17786);
and U18059 (N_18059,N_16312,N_16319);
and U18060 (N_18060,N_16670,N_17907);
nand U18061 (N_18061,N_17230,N_16772);
nor U18062 (N_18062,N_16775,N_16905);
xnor U18063 (N_18063,N_17115,N_16000);
nor U18064 (N_18064,N_16067,N_17011);
or U18065 (N_18065,N_17641,N_17351);
and U18066 (N_18066,N_16528,N_16640);
and U18067 (N_18067,N_16292,N_16269);
and U18068 (N_18068,N_16354,N_16178);
xnor U18069 (N_18069,N_17083,N_17137);
nand U18070 (N_18070,N_17985,N_16099);
nand U18071 (N_18071,N_16659,N_17839);
or U18072 (N_18072,N_17724,N_17876);
xor U18073 (N_18073,N_17387,N_16994);
and U18074 (N_18074,N_17391,N_17223);
nand U18075 (N_18075,N_16223,N_16427);
nor U18076 (N_18076,N_16170,N_17898);
or U18077 (N_18077,N_16773,N_17144);
nor U18078 (N_18078,N_17611,N_17533);
or U18079 (N_18079,N_16596,N_16222);
nand U18080 (N_18080,N_17128,N_17091);
nor U18081 (N_18081,N_17352,N_16790);
nor U18082 (N_18082,N_17731,N_16401);
xnor U18083 (N_18083,N_16914,N_17506);
or U18084 (N_18084,N_16061,N_17660);
xnor U18085 (N_18085,N_17220,N_16253);
xnor U18086 (N_18086,N_17740,N_16954);
xor U18087 (N_18087,N_17695,N_16296);
nand U18088 (N_18088,N_16323,N_17282);
nand U18089 (N_18089,N_17395,N_16821);
or U18090 (N_18090,N_16495,N_17487);
xor U18091 (N_18091,N_17164,N_17439);
nor U18092 (N_18092,N_16122,N_16692);
nor U18093 (N_18093,N_16349,N_16988);
or U18094 (N_18094,N_17274,N_16117);
xnor U18095 (N_18095,N_16642,N_17713);
xor U18096 (N_18096,N_16127,N_16155);
or U18097 (N_18097,N_17622,N_16396);
or U18098 (N_18098,N_17916,N_16798);
xor U18099 (N_18099,N_16442,N_17237);
and U18100 (N_18100,N_16793,N_16357);
or U18101 (N_18101,N_16889,N_17944);
nand U18102 (N_18102,N_17716,N_17929);
and U18103 (N_18103,N_17776,N_16559);
xor U18104 (N_18104,N_16120,N_16944);
or U18105 (N_18105,N_17581,N_16239);
nand U18106 (N_18106,N_16909,N_17447);
nor U18107 (N_18107,N_17712,N_17911);
or U18108 (N_18108,N_16947,N_16393);
and U18109 (N_18109,N_17790,N_17890);
nor U18110 (N_18110,N_17076,N_16094);
or U18111 (N_18111,N_17688,N_17885);
xnor U18112 (N_18112,N_16441,N_17328);
and U18113 (N_18113,N_16262,N_16325);
and U18114 (N_18114,N_17116,N_16915);
nor U18115 (N_18115,N_16871,N_16599);
nor U18116 (N_18116,N_16158,N_17406);
and U18117 (N_18117,N_17700,N_17933);
or U18118 (N_18118,N_16465,N_16408);
and U18119 (N_18119,N_17206,N_16055);
and U18120 (N_18120,N_17359,N_16274);
nor U18121 (N_18121,N_16488,N_17058);
or U18122 (N_18122,N_17743,N_17329);
nand U18123 (N_18123,N_16027,N_16916);
and U18124 (N_18124,N_16433,N_16159);
nor U18125 (N_18125,N_17863,N_16413);
and U18126 (N_18126,N_16753,N_17131);
xor U18127 (N_18127,N_16343,N_16968);
xor U18128 (N_18128,N_16926,N_17270);
nor U18129 (N_18129,N_16643,N_16355);
xnor U18130 (N_18130,N_17880,N_17216);
xor U18131 (N_18131,N_16966,N_16581);
or U18132 (N_18132,N_17803,N_17215);
nor U18133 (N_18133,N_16813,N_17523);
nand U18134 (N_18134,N_17267,N_17041);
and U18135 (N_18135,N_16378,N_16661);
xor U18136 (N_18136,N_17819,N_17612);
nand U18137 (N_18137,N_16161,N_17782);
and U18138 (N_18138,N_16140,N_17926);
nor U18139 (N_18139,N_17298,N_17574);
or U18140 (N_18140,N_16571,N_17313);
or U18141 (N_18141,N_17124,N_17970);
nand U18142 (N_18142,N_16678,N_16676);
nand U18143 (N_18143,N_17242,N_17756);
nor U18144 (N_18144,N_17748,N_16685);
and U18145 (N_18145,N_16414,N_17588);
and U18146 (N_18146,N_16929,N_16848);
and U18147 (N_18147,N_17494,N_17928);
and U18148 (N_18148,N_16636,N_17526);
and U18149 (N_18149,N_16626,N_16902);
or U18150 (N_18150,N_17524,N_16760);
nor U18151 (N_18151,N_16549,N_16483);
xor U18152 (N_18152,N_17073,N_17818);
nor U18153 (N_18153,N_16031,N_17381);
nand U18154 (N_18154,N_16407,N_16814);
nor U18155 (N_18155,N_17857,N_17904);
nand U18156 (N_18156,N_17209,N_16123);
nor U18157 (N_18157,N_17889,N_17311);
xor U18158 (N_18158,N_16226,N_17132);
and U18159 (N_18159,N_16147,N_17993);
nand U18160 (N_18160,N_16696,N_16650);
and U18161 (N_18161,N_16469,N_17227);
and U18162 (N_18162,N_16308,N_17405);
nand U18163 (N_18163,N_17178,N_17915);
nor U18164 (N_18164,N_16432,N_16026);
xnor U18165 (N_18165,N_16220,N_16175);
nor U18166 (N_18166,N_16801,N_16564);
nand U18167 (N_18167,N_17771,N_16639);
or U18168 (N_18168,N_17251,N_16208);
or U18169 (N_18169,N_16656,N_17390);
and U18170 (N_18170,N_16374,N_16307);
nand U18171 (N_18171,N_16411,N_16029);
and U18172 (N_18172,N_17593,N_16205);
xnor U18173 (N_18173,N_17648,N_16115);
nor U18174 (N_18174,N_16959,N_16416);
and U18175 (N_18175,N_16674,N_17262);
and U18176 (N_18176,N_17983,N_17175);
nand U18177 (N_18177,N_17231,N_16256);
or U18178 (N_18178,N_17193,N_17589);
nor U18179 (N_18179,N_16820,N_17561);
and U18180 (N_18180,N_17763,N_16265);
and U18181 (N_18181,N_16494,N_17651);
xnor U18182 (N_18182,N_17015,N_16045);
xor U18183 (N_18183,N_17285,N_16754);
nor U18184 (N_18184,N_17597,N_17860);
nor U18185 (N_18185,N_17444,N_16286);
nand U18186 (N_18186,N_16702,N_17821);
and U18187 (N_18187,N_17169,N_16936);
nand U18188 (N_18188,N_16863,N_16006);
xnor U18189 (N_18189,N_17728,N_17718);
xor U18190 (N_18190,N_16880,N_17343);
nand U18191 (N_18191,N_16574,N_17618);
or U18192 (N_18192,N_17276,N_16669);
nand U18193 (N_18193,N_17601,N_17383);
xnor U18194 (N_18194,N_17198,N_17917);
or U18195 (N_18195,N_16383,N_17752);
nand U18196 (N_18196,N_16489,N_17170);
nand U18197 (N_18197,N_16651,N_17999);
and U18198 (N_18198,N_16671,N_17708);
and U18199 (N_18199,N_16195,N_17665);
xor U18200 (N_18200,N_17243,N_17201);
xor U18201 (N_18201,N_16553,N_16129);
nor U18202 (N_18202,N_16971,N_16338);
nor U18203 (N_18203,N_17955,N_16799);
nand U18204 (N_18204,N_17317,N_17684);
nand U18205 (N_18205,N_17195,N_16181);
nand U18206 (N_18206,N_17431,N_16939);
and U18207 (N_18207,N_17802,N_16160);
nor U18208 (N_18208,N_16254,N_16508);
and U18209 (N_18209,N_17501,N_17682);
xnor U18210 (N_18210,N_17527,N_16498);
and U18211 (N_18211,N_17678,N_16995);
nor U18212 (N_18212,N_16940,N_16403);
or U18213 (N_18213,N_17275,N_16400);
nand U18214 (N_18214,N_17505,N_16417);
nor U18215 (N_18215,N_17445,N_17967);
nor U18216 (N_18216,N_17241,N_17585);
nor U18217 (N_18217,N_17071,N_16248);
nand U18218 (N_18218,N_17417,N_17845);
nor U18219 (N_18219,N_17510,N_17530);
nand U18220 (N_18220,N_16758,N_17280);
nor U18221 (N_18221,N_16686,N_17554);
or U18222 (N_18222,N_17779,N_16885);
or U18223 (N_18223,N_16237,N_16154);
xnor U18224 (N_18224,N_17326,N_16548);
nor U18225 (N_18225,N_17875,N_16879);
nor U18226 (N_18226,N_17564,N_17174);
and U18227 (N_18227,N_17172,N_17511);
nor U18228 (N_18228,N_16665,N_17308);
or U18229 (N_18229,N_17772,N_16247);
nand U18230 (N_18230,N_16996,N_16965);
xnor U18231 (N_18231,N_16743,N_17987);
xnor U18232 (N_18232,N_16795,N_17454);
nor U18233 (N_18233,N_17951,N_17353);
nand U18234 (N_18234,N_16828,N_17134);
xnor U18235 (N_18235,N_16884,N_17703);
and U18236 (N_18236,N_17701,N_16337);
xor U18237 (N_18237,N_17532,N_17438);
and U18238 (N_18238,N_17872,N_17182);
or U18239 (N_18239,N_16989,N_16313);
and U18240 (N_18240,N_17153,N_17563);
nand U18241 (N_18241,N_16196,N_17942);
nand U18242 (N_18242,N_16891,N_16013);
nand U18243 (N_18243,N_16835,N_16532);
and U18244 (N_18244,N_16960,N_17903);
xnor U18245 (N_18245,N_17222,N_16451);
and U18246 (N_18246,N_17067,N_17957);
or U18247 (N_18247,N_16452,N_16784);
nand U18248 (N_18248,N_16005,N_16750);
nor U18249 (N_18249,N_16377,N_17052);
nand U18250 (N_18250,N_17043,N_17960);
or U18251 (N_18251,N_17859,N_17964);
and U18252 (N_18252,N_17809,N_16928);
or U18253 (N_18253,N_16725,N_16172);
nor U18254 (N_18254,N_16973,N_16764);
and U18255 (N_18255,N_16728,N_16143);
and U18256 (N_18256,N_16097,N_16156);
xnor U18257 (N_18257,N_16935,N_16091);
or U18258 (N_18258,N_17635,N_17503);
xor U18259 (N_18259,N_17314,N_17252);
nor U18260 (N_18260,N_16276,N_17344);
nand U18261 (N_18261,N_16198,N_16070);
xnor U18262 (N_18262,N_17507,N_16846);
and U18263 (N_18263,N_16920,N_17232);
and U18264 (N_18264,N_17111,N_17316);
xor U18265 (N_18265,N_17699,N_17927);
nand U18266 (N_18266,N_16851,N_16368);
or U18267 (N_18267,N_16924,N_16938);
and U18268 (N_18268,N_17744,N_17742);
nor U18269 (N_18269,N_16141,N_16534);
or U18270 (N_18270,N_17722,N_17571);
nor U18271 (N_18271,N_16487,N_16679);
nand U18272 (N_18272,N_16723,N_17977);
xor U18273 (N_18273,N_17047,N_16106);
nor U18274 (N_18274,N_17902,N_16149);
or U18275 (N_18275,N_17407,N_17514);
nand U18276 (N_18276,N_16941,N_16539);
and U18277 (N_18277,N_16242,N_17517);
xnor U18278 (N_18278,N_16504,N_17781);
xor U18279 (N_18279,N_17304,N_17382);
xor U18280 (N_18280,N_17664,N_17477);
nor U18281 (N_18281,N_16583,N_16856);
or U18282 (N_18282,N_16311,N_17009);
or U18283 (N_18283,N_16364,N_16521);
nor U18284 (N_18284,N_16506,N_17372);
xor U18285 (N_18285,N_17804,N_16300);
and U18286 (N_18286,N_17485,N_16500);
and U18287 (N_18287,N_17632,N_17306);
nor U18288 (N_18288,N_16346,N_17458);
nand U18289 (N_18289,N_17050,N_16322);
nand U18290 (N_18290,N_17394,N_17065);
or U18291 (N_18291,N_17261,N_16152);
xor U18292 (N_18292,N_17211,N_16998);
nand U18293 (N_18293,N_17366,N_16682);
nand U18294 (N_18294,N_16225,N_16216);
and U18295 (N_18295,N_17339,N_17495);
or U18296 (N_18296,N_16474,N_16387);
xor U18297 (N_18297,N_16918,N_16082);
or U18298 (N_18298,N_17758,N_16526);
xor U18299 (N_18299,N_16184,N_16363);
nor U18300 (N_18300,N_16955,N_16369);
or U18301 (N_18301,N_17026,N_16683);
xnor U18302 (N_18302,N_16654,N_16601);
nor U18303 (N_18303,N_17663,N_17441);
and U18304 (N_18304,N_17246,N_16752);
xnor U18305 (N_18305,N_16471,N_17850);
xor U18306 (N_18306,N_16365,N_17555);
nor U18307 (N_18307,N_16490,N_17649);
nand U18308 (N_18308,N_16294,N_16252);
or U18309 (N_18309,N_17093,N_17012);
nand U18310 (N_18310,N_17921,N_17300);
xnor U18311 (N_18311,N_17738,N_16672);
and U18312 (N_18312,N_17433,N_17403);
and U18313 (N_18313,N_16418,N_16986);
nand U18314 (N_18314,N_16980,N_17624);
or U18315 (N_18315,N_16781,N_16439);
nand U18316 (N_18316,N_16729,N_16903);
nor U18317 (N_18317,N_16745,N_16537);
or U18318 (N_18318,N_17551,N_16270);
or U18319 (N_18319,N_16116,N_16942);
nor U18320 (N_18320,N_16190,N_17055);
nand U18321 (N_18321,N_17842,N_16361);
nor U18322 (N_18322,N_16660,N_17825);
and U18323 (N_18323,N_17698,N_17320);
nor U18324 (N_18324,N_17614,N_16822);
and U18325 (N_18325,N_16957,N_16817);
and U18326 (N_18326,N_16295,N_16710);
and U18327 (N_18327,N_17709,N_16623);
xor U18328 (N_18328,N_16095,N_17913);
nor U18329 (N_18329,N_17751,N_17787);
nor U18330 (N_18330,N_17806,N_17187);
nand U18331 (N_18331,N_16321,N_16481);
and U18332 (N_18332,N_16063,N_16092);
and U18333 (N_18333,N_16479,N_17392);
nand U18334 (N_18334,N_17687,N_16653);
or U18335 (N_18335,N_16386,N_16853);
nand U18336 (N_18336,N_17254,N_16932);
nor U18337 (N_18337,N_16572,N_17181);
nor U18338 (N_18338,N_16328,N_16808);
or U18339 (N_18339,N_17521,N_16628);
and U18340 (N_18340,N_16203,N_17662);
nand U18341 (N_18341,N_16749,N_17646);
or U18342 (N_18342,N_16280,N_17443);
xor U18343 (N_18343,N_17998,N_16619);
or U18344 (N_18344,N_16782,N_16701);
and U18345 (N_18345,N_17375,N_17452);
and U18346 (N_18346,N_16570,N_17798);
and U18347 (N_18347,N_17948,N_17402);
nor U18348 (N_18348,N_16740,N_16815);
xor U18349 (N_18349,N_17021,N_16284);
nand U18350 (N_18350,N_17310,N_17036);
or U18351 (N_18351,N_17024,N_16087);
and U18352 (N_18352,N_17152,N_17122);
or U18353 (N_18353,N_16255,N_17656);
nand U18354 (N_18354,N_16961,N_17129);
nor U18355 (N_18355,N_16019,N_17749);
or U18356 (N_18356,N_17468,N_16768);
and U18357 (N_18357,N_16096,N_16896);
or U18358 (N_18358,N_16228,N_16282);
xnor U18359 (N_18359,N_17690,N_16552);
or U18360 (N_18360,N_17284,N_17360);
xnor U18361 (N_18361,N_17925,N_17389);
or U18362 (N_18362,N_17342,N_16792);
nand U18363 (N_18363,N_16541,N_17941);
or U18364 (N_18364,N_17730,N_17264);
and U18365 (N_18365,N_16895,N_16073);
or U18366 (N_18366,N_17637,N_17318);
nand U18367 (N_18367,N_17448,N_16529);
nor U18368 (N_18368,N_17856,N_17064);
nor U18369 (N_18369,N_17886,N_16204);
xnor U18370 (N_18370,N_17239,N_16951);
xnor U18371 (N_18371,N_17943,N_17042);
and U18372 (N_18372,N_17221,N_17636);
and U18373 (N_18373,N_16925,N_17667);
nand U18374 (N_18374,N_17573,N_17238);
and U18375 (N_18375,N_17105,N_17409);
nor U18376 (N_18376,N_16259,N_17789);
or U18377 (N_18377,N_16150,N_17714);
nor U18378 (N_18378,N_16563,N_17101);
or U18379 (N_18379,N_16366,N_16192);
nand U18380 (N_18380,N_17281,N_17732);
xor U18381 (N_18381,N_17775,N_16064);
xor U18382 (N_18382,N_17661,N_17460);
nor U18383 (N_18383,N_16756,N_16733);
or U18384 (N_18384,N_16796,N_16803);
and U18385 (N_18385,N_16969,N_16069);
xor U18386 (N_18386,N_17644,N_17783);
or U18387 (N_18387,N_16949,N_17531);
nand U18388 (N_18388,N_17504,N_16218);
xnor U18389 (N_18389,N_16809,N_16477);
nor U18390 (N_18390,N_17676,N_16011);
or U18391 (N_18391,N_16125,N_16778);
nand U18392 (N_18392,N_17340,N_17720);
or U18393 (N_18393,N_16514,N_17746);
or U18394 (N_18394,N_17007,N_16340);
nor U18395 (N_18395,N_17719,N_17568);
xnor U18396 (N_18396,N_16587,N_17399);
nand U18397 (N_18397,N_16136,N_16327);
nor U18398 (N_18398,N_16139,N_16179);
or U18399 (N_18399,N_17697,N_17575);
nor U18400 (N_18400,N_17871,N_16970);
nand U18401 (N_18401,N_16577,N_16862);
xor U18402 (N_18402,N_17186,N_16375);
xnor U18403 (N_18403,N_16899,N_16409);
xnor U18404 (N_18404,N_17145,N_17435);
or U18405 (N_18405,N_17140,N_16014);
or U18406 (N_18406,N_16397,N_17814);
or U18407 (N_18407,N_16726,N_17240);
and U18408 (N_18408,N_17081,N_17671);
xor U18409 (N_18409,N_16472,N_16215);
and U18410 (N_18410,N_16588,N_16687);
or U18411 (N_18411,N_17048,N_16789);
xnor U18412 (N_18412,N_16907,N_17099);
and U18413 (N_18413,N_16032,N_16350);
or U18414 (N_18414,N_17537,N_17436);
xnor U18415 (N_18415,N_17710,N_17670);
and U18416 (N_18416,N_16573,N_16306);
or U18417 (N_18417,N_17705,N_17768);
or U18418 (N_18418,N_16410,N_16492);
or U18419 (N_18419,N_16075,N_16034);
nand U18420 (N_18420,N_17033,N_17423);
or U18421 (N_18421,N_17778,N_16585);
or U18422 (N_18422,N_16449,N_16493);
nor U18423 (N_18423,N_17715,N_17725);
xor U18424 (N_18424,N_17547,N_17834);
nor U18425 (N_18425,N_16721,N_17484);
nand U18426 (N_18426,N_16381,N_17465);
or U18427 (N_18427,N_16243,N_16836);
nand U18428 (N_18428,N_16310,N_17330);
xor U18429 (N_18429,N_16993,N_17008);
nand U18430 (N_18430,N_17400,N_16617);
or U18431 (N_18431,N_16841,N_16134);
nand U18432 (N_18432,N_17290,N_16810);
and U18433 (N_18433,N_16315,N_16520);
nand U18434 (N_18434,N_16478,N_17031);
nor U18435 (N_18435,N_16456,N_16657);
or U18436 (N_18436,N_17257,N_16591);
and U18437 (N_18437,N_16036,N_16645);
xnor U18438 (N_18438,N_17397,N_17357);
and U18439 (N_18439,N_16157,N_16893);
and U18440 (N_18440,N_17693,N_16335);
or U18441 (N_18441,N_17418,N_17668);
nor U18442 (N_18442,N_16051,N_16834);
xnor U18443 (N_18443,N_17371,N_17605);
nor U18444 (N_18444,N_17475,N_17190);
nand U18445 (N_18445,N_17023,N_16077);
or U18446 (N_18446,N_17226,N_17986);
or U18447 (N_18447,N_17463,N_17565);
nor U18448 (N_18448,N_16625,N_17673);
or U18449 (N_18449,N_16385,N_17761);
xor U18450 (N_18450,N_16987,N_16206);
and U18451 (N_18451,N_17385,N_16110);
xor U18452 (N_18452,N_16207,N_16405);
and U18453 (N_18453,N_16180,N_17380);
or U18454 (N_18454,N_17529,N_16246);
nand U18455 (N_18455,N_17577,N_17723);
nand U18456 (N_18456,N_17269,N_16886);
and U18457 (N_18457,N_17032,N_16499);
or U18458 (N_18458,N_16807,N_16830);
xnor U18459 (N_18459,N_16104,N_16611);
nand U18460 (N_18460,N_16904,N_16839);
xor U18461 (N_18461,N_16059,N_16043);
nand U18462 (N_18462,N_17643,N_17522);
nand U18463 (N_18463,N_16038,N_17367);
or U18464 (N_18464,N_16309,N_16468);
and U18465 (N_18465,N_16878,N_16704);
and U18466 (N_18466,N_16089,N_17658);
or U18467 (N_18467,N_17583,N_16712);
or U18468 (N_18468,N_16797,N_17931);
xor U18469 (N_18469,N_16751,N_16551);
nor U18470 (N_18470,N_16616,N_16658);
nand U18471 (N_18471,N_16937,N_17356);
xor U18472 (N_18472,N_17920,N_16316);
or U18473 (N_18473,N_17733,N_17793);
or U18474 (N_18474,N_17347,N_17923);
xnor U18475 (N_18475,N_17613,N_16523);
and U18476 (N_18476,N_17579,N_16948);
xor U18477 (N_18477,N_17070,N_16126);
xnor U18478 (N_18478,N_17674,N_16166);
nand U18479 (N_18479,N_17333,N_17509);
nand U18480 (N_18480,N_17604,N_17046);
nor U18481 (N_18481,N_16395,N_16887);
and U18482 (N_18482,N_17324,N_16984);
and U18483 (N_18483,N_17841,N_16037);
or U18484 (N_18484,N_16461,N_17498);
or U18485 (N_18485,N_16805,N_16114);
and U18486 (N_18486,N_16348,N_16336);
and U18487 (N_18487,N_16339,N_17069);
xnor U18488 (N_18488,N_16974,N_16762);
nor U18489 (N_18489,N_17666,N_17840);
nor U18490 (N_18490,N_17214,N_17272);
nor U18491 (N_18491,N_16575,N_16964);
xor U18492 (N_18492,N_17429,N_17141);
nor U18493 (N_18493,N_17212,N_17411);
and U18494 (N_18494,N_17266,N_16426);
or U18495 (N_18495,N_16633,N_16722);
or U18496 (N_18496,N_16389,N_16202);
xnor U18497 (N_18497,N_17259,N_17106);
and U18498 (N_18498,N_16544,N_16496);
xnor U18499 (N_18499,N_16419,N_16858);
nand U18500 (N_18500,N_17654,N_17810);
xnor U18501 (N_18501,N_17535,N_16579);
and U18502 (N_18502,N_16074,N_17826);
nor U18503 (N_18503,N_17813,N_16716);
nand U18504 (N_18504,N_16849,N_17692);
or U18505 (N_18505,N_16763,N_17278);
nor U18506 (N_18506,N_17027,N_16662);
xnor U18507 (N_18507,N_17118,N_17039);
nand U18508 (N_18508,N_16266,N_17168);
nand U18509 (N_18509,N_16646,N_16124);
or U18510 (N_18510,N_16399,N_16076);
nand U18511 (N_18511,N_17621,N_16236);
or U18512 (N_18512,N_16690,N_17176);
or U18513 (N_18513,N_17994,N_17541);
or U18514 (N_18514,N_17286,N_17303);
xor U18515 (N_18515,N_16463,N_17735);
xnor U18516 (N_18516,N_16080,N_16227);
or U18517 (N_18517,N_17133,N_16829);
and U18518 (N_18518,N_17325,N_16894);
or U18519 (N_18519,N_16664,N_17861);
nor U18520 (N_18520,N_16101,N_16511);
xor U18521 (N_18521,N_17766,N_16454);
nor U18522 (N_18522,N_16111,N_16542);
nand U18523 (N_18523,N_17358,N_16543);
nand U18524 (N_18524,N_16761,N_16201);
or U18525 (N_18525,N_16912,N_16732);
xnor U18526 (N_18526,N_17154,N_16770);
xor U18527 (N_18527,N_17745,N_17457);
or U18528 (N_18528,N_17808,N_16450);
and U18529 (N_18529,N_17388,N_17361);
nand U18530 (N_18530,N_16545,N_17835);
or U18531 (N_18531,N_17580,N_16991);
and U18532 (N_18532,N_16371,N_16981);
xor U18533 (N_18533,N_16380,N_17001);
or U18534 (N_18534,N_16739,N_17877);
and U18535 (N_18535,N_17811,N_17179);
and U18536 (N_18536,N_17874,N_16283);
and U18537 (N_18537,N_17301,N_16415);
nor U18538 (N_18538,N_16457,N_16058);
nand U18539 (N_18539,N_17940,N_16039);
and U18540 (N_18540,N_17896,N_16695);
xnor U18541 (N_18541,N_16428,N_16609);
nor U18542 (N_18542,N_17481,N_17852);
nor U18543 (N_18543,N_16906,N_16304);
nor U18544 (N_18544,N_16597,N_17946);
xnor U18545 (N_18545,N_17053,N_17696);
or U18546 (N_18546,N_16533,N_16176);
nand U18547 (N_18547,N_17785,N_16742);
nor U18548 (N_18548,N_16017,N_17249);
xnor U18549 (N_18549,N_16210,N_16557);
nand U18550 (N_18550,N_17114,N_16021);
or U18551 (N_18551,N_16056,N_17138);
nor U18552 (N_18552,N_16898,N_17848);
or U18553 (N_18553,N_17953,N_16244);
or U18554 (N_18554,N_17978,N_16708);
nand U18555 (N_18555,N_16524,N_17686);
nor U18556 (N_18556,N_17726,N_16908);
nand U18557 (N_18557,N_17868,N_17255);
and U18558 (N_18558,N_17126,N_17924);
nand U18559 (N_18559,N_17553,N_17098);
and U18560 (N_18560,N_16566,N_17334);
nand U18561 (N_18561,N_17906,N_16622);
nand U18562 (N_18562,N_17283,N_17515);
or U18563 (N_18563,N_16020,N_16466);
xor U18564 (N_18564,N_16183,N_17655);
and U18565 (N_18565,N_17121,N_16877);
or U18566 (N_18566,N_17685,N_16185);
xnor U18567 (N_18567,N_16135,N_16607);
nor U18568 (N_18568,N_17453,N_17512);
nor U18569 (N_18569,N_17905,N_16287);
or U18570 (N_18570,N_17559,N_16855);
xnor U18571 (N_18571,N_16165,N_16440);
nand U18572 (N_18572,N_16113,N_17045);
nand U18573 (N_18573,N_17348,N_17909);
xnor U18574 (N_18574,N_17566,N_17207);
nor U18575 (N_18575,N_16301,N_16655);
nand U18576 (N_18576,N_16001,N_17097);
xnor U18577 (N_18577,N_16978,N_17100);
nand U18578 (N_18578,N_16714,N_17480);
xnor U18579 (N_18579,N_16538,N_17600);
xor U18580 (N_18580,N_17037,N_17828);
xor U18581 (N_18581,N_16923,N_17689);
nor U18582 (N_18582,N_16505,N_17812);
nor U18583 (N_18583,N_16594,N_16791);
or U18584 (N_18584,N_16718,N_16187);
xor U18585 (N_18585,N_16681,N_17820);
nand U18586 (N_18586,N_16602,N_17057);
nor U18587 (N_18587,N_16351,N_16015);
nand U18588 (N_18588,N_17767,N_16547);
or U18589 (N_18589,N_17975,N_16689);
xor U18590 (N_18590,N_17202,N_17142);
nor U18591 (N_18591,N_16736,N_17591);
or U18592 (N_18592,N_17474,N_17950);
and U18593 (N_18593,N_17379,N_16612);
nand U18594 (N_18594,N_16608,N_16724);
xnor U18595 (N_18595,N_16291,N_16331);
nand U18596 (N_18596,N_16869,N_17570);
nand U18597 (N_18597,N_17442,N_17592);
and U18598 (N_18598,N_17608,N_16913);
xnor U18599 (N_18599,N_16093,N_17233);
nor U18600 (N_18600,N_17888,N_16535);
nor U18601 (N_18601,N_16840,N_17365);
nor U18602 (N_18602,N_17792,N_17426);
nor U18603 (N_18603,N_16299,N_16360);
nand U18604 (N_18604,N_16108,N_16832);
or U18605 (N_18605,N_16525,N_17853);
nor U18606 (N_18606,N_17245,N_17963);
or U18607 (N_18607,N_17197,N_16590);
xnor U18608 (N_18608,N_17005,N_16334);
and U18609 (N_18609,N_17502,N_16509);
or U18610 (N_18610,N_17838,N_17516);
xor U18611 (N_18611,N_17125,N_16145);
nor U18612 (N_18612,N_16876,N_16584);
nor U18613 (N_18613,N_16010,N_16470);
nor U18614 (N_18614,N_16589,N_16691);
nor U18615 (N_18615,N_16434,N_17539);
or U18616 (N_18616,N_16921,N_17492);
nand U18617 (N_18617,N_16648,N_17321);
and U18618 (N_18618,N_16016,N_17755);
xnor U18619 (N_18619,N_16279,N_17336);
and U18620 (N_18620,N_16376,N_16329);
nor U18621 (N_18621,N_17870,N_17645);
nand U18622 (N_18622,N_16464,N_17794);
nor U18623 (N_18623,N_16049,N_17638);
and U18624 (N_18624,N_17331,N_16144);
and U18625 (N_18625,N_17077,N_17250);
or U18626 (N_18626,N_16515,N_17603);
xor U18627 (N_18627,N_17225,N_17862);
nand U18628 (N_18628,N_17119,N_16600);
or U18629 (N_18629,N_17159,N_17247);
or U18630 (N_18630,N_17120,N_17364);
nor U18631 (N_18631,N_16437,N_17582);
nand U18632 (N_18632,N_16629,N_17054);
xor U18633 (N_18633,N_17939,N_17002);
and U18634 (N_18634,N_16162,N_16857);
and U18635 (N_18635,N_16224,N_16663);
and U18636 (N_18636,N_17969,N_16777);
or U18637 (N_18637,N_16219,N_17882);
and U18638 (N_18638,N_16755,N_17590);
nand U18639 (N_18639,N_16444,N_17292);
and U18640 (N_18640,N_17945,N_17470);
xnor U18641 (N_18641,N_16546,N_16238);
and U18642 (N_18642,N_17235,N_17596);
nor U18643 (N_18643,N_17151,N_17892);
nand U18644 (N_18644,N_17337,N_16890);
and U18645 (N_18645,N_17958,N_17996);
xor U18646 (N_18646,N_16802,N_17647);
xor U18647 (N_18647,N_16819,N_16173);
nand U18648 (N_18648,N_16231,N_16052);
nand U18649 (N_18649,N_16002,N_17534);
or U18650 (N_18650,N_16028,N_16462);
nand U18651 (N_18651,N_16406,N_17386);
or U18652 (N_18652,N_16030,N_16476);
or U18653 (N_18653,N_17630,N_17873);
xor U18654 (N_18654,N_16497,N_17369);
and U18655 (N_18655,N_17991,N_16040);
nand U18656 (N_18656,N_16084,N_16715);
nor U18657 (N_18657,N_16424,N_17625);
nor U18658 (N_18658,N_17962,N_17901);
and U18659 (N_18659,N_16873,N_16975);
nand U18660 (N_18660,N_17595,N_16212);
and U18661 (N_18661,N_16555,N_17213);
or U18662 (N_18662,N_16519,N_17377);
and U18663 (N_18663,N_17727,N_16267);
nor U18664 (N_18664,N_17679,N_16098);
xnor U18665 (N_18665,N_17653,N_17824);
nand U18666 (N_18666,N_17628,N_17865);
nand U18667 (N_18667,N_17432,N_17160);
nand U18668 (N_18668,N_17472,N_17777);
nor U18669 (N_18669,N_16009,N_16131);
xnor U18670 (N_18670,N_17157,N_16429);
and U18671 (N_18671,N_17711,N_16384);
nand U18672 (N_18672,N_16303,N_16649);
nand U18673 (N_18673,N_16044,N_16576);
nand U18674 (N_18674,N_17341,N_16867);
or U18675 (N_18675,N_16618,N_17897);
nor U18676 (N_18676,N_17992,N_16605);
nor U18677 (N_18677,N_17434,N_17062);
or U18678 (N_18678,N_16927,N_16956);
or U18679 (N_18679,N_16090,N_17883);
and U18680 (N_18680,N_17412,N_16558);
nor U18681 (N_18681,N_16567,N_17639);
and U18682 (N_18682,N_16503,N_17919);
nand U18683 (N_18683,N_16731,N_16445);
and U18684 (N_18684,N_16394,N_16847);
nor U18685 (N_18685,N_16048,N_17843);
and U18686 (N_18686,N_16680,N_17764);
nand U18687 (N_18687,N_17520,N_16086);
and U18688 (N_18688,N_16620,N_17210);
and U18689 (N_18689,N_17188,N_16866);
or U18690 (N_18690,N_16945,N_16453);
xnor U18691 (N_18691,N_17866,N_17332);
or U18692 (N_18692,N_16967,N_16874);
nand U18693 (N_18693,N_17349,N_17629);
nand U18694 (N_18694,N_17801,N_16352);
and U18695 (N_18695,N_17576,N_17891);
and U18696 (N_18696,N_16741,N_16278);
or U18697 (N_18697,N_17881,N_16314);
nand U18698 (N_18698,N_16345,N_17224);
nor U18699 (N_18699,N_16711,N_16233);
and U18700 (N_18700,N_17519,N_16137);
or U18701 (N_18701,N_16194,N_17499);
xnor U18702 (N_18702,N_17918,N_16467);
nor U18703 (N_18703,N_17374,N_17378);
nor U18704 (N_18704,N_17569,N_17363);
nor U18705 (N_18705,N_16675,N_17833);
nand U18706 (N_18706,N_16392,N_17288);
nor U18707 (N_18707,N_17816,N_16510);
nor U18708 (N_18708,N_17416,N_17525);
nor U18709 (N_18709,N_17619,N_17309);
xnor U18710 (N_18710,N_16774,N_17095);
and U18711 (N_18711,N_16344,N_17704);
nor U18712 (N_18712,N_16720,N_17127);
nand U18713 (N_18713,N_16151,N_17074);
and U18714 (N_18714,N_16746,N_16263);
nand U18715 (N_18715,N_16358,N_17988);
xor U18716 (N_18716,N_16264,N_17769);
and U18717 (N_18717,N_16412,N_16677);
and U18718 (N_18718,N_17107,N_17229);
nor U18719 (N_18719,N_16769,N_16826);
xor U18720 (N_18720,N_17289,N_17959);
and U18721 (N_18721,N_17846,N_17900);
nor U18722 (N_18722,N_17599,N_16540);
nand U18723 (N_18723,N_17681,N_17459);
nor U18724 (N_18724,N_17158,N_17717);
nor U18725 (N_18725,N_16372,N_17741);
and U18726 (N_18726,N_16455,N_17914);
nand U18727 (N_18727,N_16103,N_16485);
and U18728 (N_18728,N_17844,N_16554);
xnor U18729 (N_18729,N_17557,N_16257);
or U18730 (N_18730,N_17087,N_16910);
or U18731 (N_18731,N_16776,N_17189);
nor U18732 (N_18732,N_16946,N_16888);
xor U18733 (N_18733,N_17263,N_16171);
nor U18734 (N_18734,N_17543,N_17061);
and U18735 (N_18735,N_17112,N_17770);
or U18736 (N_18736,N_16460,N_16717);
nand U18737 (N_18737,N_17205,N_16963);
nor U18738 (N_18738,N_16958,N_17236);
xor U18739 (N_18739,N_16634,N_16102);
nand U18740 (N_18740,N_17762,N_17702);
or U18741 (N_18741,N_16105,N_16513);
or U18742 (N_18742,N_16582,N_17410);
nand U18743 (N_18743,N_16277,N_17302);
nand U18744 (N_18744,N_16816,N_16647);
or U18745 (N_18745,N_17832,N_17598);
and U18746 (N_18746,N_16624,N_16703);
nand U18747 (N_18747,N_16766,N_17109);
xor U18748 (N_18748,N_17997,N_16050);
nor U18749 (N_18749,N_17419,N_16688);
and U18750 (N_18750,N_16827,N_17373);
nor U18751 (N_18751,N_16900,N_17338);
and U18752 (N_18752,N_16606,N_16119);
nor U18753 (N_18753,N_16512,N_17260);
xor U18754 (N_18754,N_16943,N_17949);
and U18755 (N_18755,N_17393,N_17019);
xor U18756 (N_18756,N_16719,N_17113);
xnor U18757 (N_18757,N_16023,N_16459);
nand U18758 (N_18758,N_17307,N_16260);
nand U18759 (N_18759,N_16561,N_16748);
nor U18760 (N_18760,N_16421,N_17268);
or U18761 (N_18761,N_17089,N_17401);
nor U18762 (N_18762,N_17947,N_17760);
and U18763 (N_18763,N_17200,N_16516);
and U18764 (N_18764,N_17044,N_17831);
nor U18765 (N_18765,N_17063,N_17578);
nand U18766 (N_18766,N_16522,N_17878);
xnor U18767 (N_18767,N_16812,N_16273);
and U18768 (N_18768,N_17010,N_16199);
xnor U18769 (N_18769,N_16843,N_16281);
xor U18770 (N_18770,N_17020,N_16517);
and U18771 (N_18771,N_17642,N_17362);
and U18772 (N_18772,N_16735,N_17014);
xor U18773 (N_18773,N_17110,N_16842);
nand U18774 (N_18774,N_17025,N_17980);
and U18775 (N_18775,N_17817,N_17084);
nor U18776 (N_18776,N_17930,N_16613);
nand U18777 (N_18777,N_17615,N_16035);
or U18778 (N_18778,N_17757,N_16088);
xor U18779 (N_18779,N_17490,N_17837);
and U18780 (N_18780,N_17258,N_16788);
xnor U18781 (N_18781,N_16825,N_16953);
and U18782 (N_18782,N_16785,N_16697);
and U18783 (N_18783,N_16771,N_16560);
nor U18784 (N_18784,N_17867,N_17545);
nand U18785 (N_18785,N_17550,N_17478);
and U18786 (N_18786,N_17973,N_17773);
or U18787 (N_18787,N_17094,N_16353);
and U18788 (N_18788,N_16302,N_16425);
nand U18789 (N_18789,N_17096,N_16163);
nor U18790 (N_18790,N_17079,N_17895);
and U18791 (N_18791,N_17694,N_17148);
nand U18792 (N_18792,N_16046,N_17086);
nor U18793 (N_18793,N_17879,N_17305);
and U18794 (N_18794,N_16527,N_17440);
nor U18795 (N_18795,N_17910,N_16610);
nand U18796 (N_18796,N_16290,N_17234);
and U18797 (N_18797,N_17368,N_17823);
xor U18798 (N_18798,N_17404,N_17556);
nand U18799 (N_18799,N_16153,N_17609);
or U18800 (N_18800,N_17623,N_16177);
nor U18801 (N_18801,N_17006,N_17464);
xor U18802 (N_18802,N_16706,N_16229);
nor U18803 (N_18803,N_16446,N_16018);
nand U18804 (N_18804,N_17346,N_16767);
xor U18805 (N_18805,N_17981,N_16390);
xor U18806 (N_18806,N_16458,N_17594);
nor U18807 (N_18807,N_17734,N_16933);
nand U18808 (N_18808,N_17354,N_17104);
and U18809 (N_18809,N_17414,N_16684);
nand U18810 (N_18810,N_16757,N_17136);
nand U18811 (N_18811,N_16250,N_16193);
nor U18812 (N_18812,N_16592,N_16004);
nor U18813 (N_18813,N_17279,N_16844);
nand U18814 (N_18814,N_17446,N_16232);
nor U18815 (N_18815,N_16298,N_16759);
or U18816 (N_18816,N_16042,N_16085);
nand U18817 (N_18817,N_17028,N_16235);
and U18818 (N_18818,N_16025,N_17488);
or U18819 (N_18819,N_16983,N_16882);
or U18820 (N_18820,N_17466,N_17683);
nand U18821 (N_18821,N_16734,N_16066);
nand U18822 (N_18822,N_16491,N_16875);
and U18823 (N_18823,N_17691,N_16241);
nand U18824 (N_18824,N_17791,N_17156);
and U18825 (N_18825,N_17072,N_17103);
xnor U18826 (N_18826,N_17018,N_16261);
xor U18827 (N_18827,N_16443,N_17774);
nand U18828 (N_18828,N_17204,N_17173);
nor U18829 (N_18829,N_17822,N_17003);
xnor U18830 (N_18830,N_17899,N_17538);
nand U18831 (N_18831,N_16293,N_17370);
xor U18832 (N_18832,N_17759,N_16627);
nand U18833 (N_18833,N_17469,N_16083);
nor U18834 (N_18834,N_17430,N_16595);
xor U18835 (N_18835,N_17327,N_16738);
or U18836 (N_18836,N_16109,N_17194);
nor U18837 (N_18837,N_17296,N_16436);
and U18838 (N_18838,N_16999,N_16041);
nor U18839 (N_18839,N_16747,N_17143);
nand U18840 (N_18840,N_17497,N_17489);
nor U18841 (N_18841,N_17248,N_17167);
nor U18842 (N_18842,N_17421,N_17199);
or U18843 (N_18843,N_17851,N_17171);
and U18844 (N_18844,N_17088,N_17467);
nor U18845 (N_18845,N_17912,N_16211);
nor U18846 (N_18846,N_17135,N_17546);
xnor U18847 (N_18847,N_16186,N_17737);
or U18848 (N_18848,N_16475,N_17652);
or U18849 (N_18849,N_17922,N_17587);
xnor U18850 (N_18850,N_16837,N_17750);
nand U18851 (N_18851,N_16614,N_16486);
and U18852 (N_18852,N_16972,N_16652);
and U18853 (N_18853,N_17558,N_17163);
xnor U18854 (N_18854,N_17449,N_16985);
xor U18855 (N_18855,N_17995,N_16060);
xor U18856 (N_18856,N_16191,N_16079);
xnor U18857 (N_18857,N_16367,N_16919);
nor U18858 (N_18858,N_16197,N_16033);
nor U18859 (N_18859,N_16054,N_16700);
or U18860 (N_18860,N_16188,N_17277);
and U18861 (N_18861,N_17068,N_17149);
xor U18862 (N_18862,N_16402,N_17150);
xor U18863 (N_18863,N_16121,N_16022);
or U18864 (N_18864,N_16860,N_17669);
nor U18865 (N_18865,N_16787,N_16550);
and U18866 (N_18866,N_17617,N_17029);
nor U18867 (N_18867,N_17117,N_16979);
nor U18868 (N_18868,N_16289,N_17540);
nor U18869 (N_18869,N_17092,N_17294);
and U18870 (N_18870,N_17765,N_16008);
or U18871 (N_18871,N_16382,N_16420);
or U18872 (N_18872,N_17355,N_17548);
or U18873 (N_18873,N_16892,N_17956);
nand U18874 (N_18874,N_17966,N_17864);
nor U18875 (N_18875,N_17706,N_16868);
nand U18876 (N_18876,N_16288,N_17253);
nand U18877 (N_18877,N_17934,N_17322);
or U18878 (N_18878,N_17022,N_17319);
xor U18879 (N_18879,N_16068,N_17345);
and U18880 (N_18880,N_16341,N_16251);
nor U18881 (N_18881,N_16641,N_16169);
xnor U18882 (N_18882,N_17729,N_17971);
nand U18883 (N_18883,N_16737,N_17560);
nor U18884 (N_18884,N_17482,N_16182);
and U18885 (N_18885,N_16637,N_16012);
and U18886 (N_18886,N_17894,N_16630);
or U18887 (N_18887,N_16272,N_17196);
and U18888 (N_18888,N_16694,N_16024);
nand U18889 (N_18889,N_17295,N_17244);
xnor U18890 (N_18890,N_17034,N_16330);
nor U18891 (N_18891,N_16635,N_16850);
nand U18892 (N_18892,N_17858,N_17471);
and U18893 (N_18893,N_17425,N_16240);
nor U18894 (N_18894,N_16473,N_16990);
nand U18895 (N_18895,N_16053,N_16130);
nand U18896 (N_18896,N_17299,N_17473);
or U18897 (N_18897,N_16536,N_17562);
nor U18898 (N_18898,N_17051,N_17155);
nor U18899 (N_18899,N_17080,N_16870);
or U18900 (N_18900,N_16744,N_16502);
xnor U18901 (N_18901,N_17056,N_17004);
nand U18902 (N_18902,N_17291,N_17483);
and U18903 (N_18903,N_17932,N_17797);
nand U18904 (N_18904,N_16707,N_16333);
or U18905 (N_18905,N_17315,N_17753);
and U18906 (N_18906,N_17680,N_17208);
and U18907 (N_18907,N_17082,N_16482);
nor U18908 (N_18908,N_16530,N_17528);
and U18909 (N_18909,N_16356,N_17035);
nand U18910 (N_18910,N_16234,N_16727);
nor U18911 (N_18911,N_17451,N_16709);
or U18912 (N_18912,N_17090,N_16818);
xnor U18913 (N_18913,N_17982,N_16072);
nor U18914 (N_18914,N_16373,N_17102);
nand U18915 (N_18915,N_16531,N_16992);
nor U18916 (N_18916,N_17549,N_16786);
and U18917 (N_18917,N_17784,N_16370);
nor U18918 (N_18918,N_16800,N_17544);
or U18919 (N_18919,N_17552,N_17536);
xor U18920 (N_18920,N_17633,N_17203);
xor U18921 (N_18921,N_16950,N_16705);
nor U18922 (N_18922,N_17486,N_16507);
xor U18923 (N_18923,N_16057,N_16811);
and U18924 (N_18924,N_17965,N_17139);
xor U18925 (N_18925,N_16423,N_16501);
and U18926 (N_18926,N_17059,N_16730);
nand U18927 (N_18927,N_17795,N_17780);
xor U18928 (N_18928,N_17938,N_17108);
or U18929 (N_18929,N_17984,N_16326);
nor U18930 (N_18930,N_16586,N_17078);
or U18931 (N_18931,N_16783,N_17166);
and U18932 (N_18932,N_17736,N_17500);
and U18933 (N_18933,N_16347,N_17672);
and U18934 (N_18934,N_17807,N_17066);
xnor U18935 (N_18935,N_17677,N_17413);
xor U18936 (N_18936,N_16667,N_16997);
nand U18937 (N_18937,N_16484,N_17075);
and U18938 (N_18938,N_17424,N_17491);
and U18939 (N_18939,N_17450,N_16071);
xor U18940 (N_18940,N_16698,N_17123);
nand U18941 (N_18941,N_16780,N_17060);
nor U18942 (N_18942,N_17836,N_17085);
xnor U18943 (N_18943,N_16003,N_16168);
xor U18944 (N_18944,N_17462,N_16604);
and U18945 (N_18945,N_16864,N_17476);
and U18946 (N_18946,N_16317,N_16779);
nand U18947 (N_18947,N_17165,N_16556);
and U18948 (N_18948,N_16854,N_16962);
xnor U18949 (N_18949,N_17952,N_16133);
or U18950 (N_18950,N_16578,N_17567);
nor U18951 (N_18951,N_17293,N_16976);
nor U18952 (N_18952,N_16065,N_17192);
nand U18953 (N_18953,N_17049,N_17815);
nor U18954 (N_18954,N_16318,N_17508);
xnor U18955 (N_18955,N_16214,N_16305);
and U18956 (N_18956,N_17384,N_16189);
nor U18957 (N_18957,N_16275,N_17228);
nor U18958 (N_18958,N_16398,N_16435);
or U18959 (N_18959,N_17437,N_16146);
nand U18960 (N_18960,N_17030,N_16666);
xor U18961 (N_18961,N_16100,N_17602);
and U18962 (N_18962,N_16430,N_16379);
or U18963 (N_18963,N_17961,N_16438);
nand U18964 (N_18964,N_17854,N_17273);
nand U18965 (N_18965,N_17847,N_17456);
and U18966 (N_18966,N_17518,N_17908);
xnor U18967 (N_18967,N_17607,N_17396);
and U18968 (N_18968,N_17297,N_16881);
nor U18969 (N_18969,N_16562,N_17935);
and U18970 (N_18970,N_17626,N_16804);
xnor U18971 (N_18971,N_16917,N_17799);
nand U18972 (N_18972,N_17788,N_16391);
and U18973 (N_18973,N_17869,N_17631);
nand U18974 (N_18974,N_17990,N_16693);
or U18975 (N_18975,N_17989,N_16245);
and U18976 (N_18976,N_17271,N_17616);
nor U18977 (N_18977,N_17350,N_16865);
xnor U18978 (N_18978,N_16631,N_17893);
nand U18979 (N_18979,N_16132,N_17829);
and U18980 (N_18980,N_16342,N_16268);
xnor U18981 (N_18981,N_17936,N_17650);
or U18982 (N_18982,N_17013,N_17627);
nor U18983 (N_18983,N_16852,N_17183);
and U18984 (N_18984,N_17017,N_16580);
xnor U18985 (N_18985,N_17420,N_17455);
or U18986 (N_18986,N_16213,N_17657);
or U18987 (N_18987,N_17620,N_17177);
nand U18988 (N_18988,N_17219,N_17000);
or U18989 (N_18989,N_17805,N_17884);
nor U18990 (N_18990,N_16258,N_17217);
and U18991 (N_18991,N_17974,N_17659);
nor U18992 (N_18992,N_17191,N_16713);
xnor U18993 (N_18993,N_17634,N_16699);
or U18994 (N_18994,N_16806,N_17855);
or U18995 (N_18995,N_17937,N_17584);
xnor U18996 (N_18996,N_17513,N_16615);
nor U18997 (N_18997,N_17428,N_17721);
or U18998 (N_18998,N_16621,N_17972);
xnor U18999 (N_18999,N_16078,N_17040);
nand U19000 (N_19000,N_17615,N_17878);
or U19001 (N_19001,N_16297,N_16652);
xnor U19002 (N_19002,N_17553,N_17656);
nor U19003 (N_19003,N_16889,N_17684);
and U19004 (N_19004,N_16402,N_17129);
xnor U19005 (N_19005,N_17641,N_16063);
or U19006 (N_19006,N_17829,N_16021);
nor U19007 (N_19007,N_16187,N_17280);
and U19008 (N_19008,N_17767,N_17036);
nand U19009 (N_19009,N_17087,N_16002);
xor U19010 (N_19010,N_17432,N_17598);
nand U19011 (N_19011,N_17792,N_16906);
or U19012 (N_19012,N_17593,N_16007);
or U19013 (N_19013,N_16600,N_17919);
nor U19014 (N_19014,N_16665,N_17035);
xnor U19015 (N_19015,N_16385,N_17876);
nand U19016 (N_19016,N_17187,N_17976);
nor U19017 (N_19017,N_17062,N_17499);
and U19018 (N_19018,N_17951,N_17580);
and U19019 (N_19019,N_17878,N_17084);
nand U19020 (N_19020,N_17663,N_17730);
nand U19021 (N_19021,N_16662,N_17102);
or U19022 (N_19022,N_17348,N_16322);
nor U19023 (N_19023,N_16956,N_16400);
and U19024 (N_19024,N_16617,N_16373);
and U19025 (N_19025,N_17843,N_16840);
nor U19026 (N_19026,N_16834,N_16703);
nand U19027 (N_19027,N_16824,N_17134);
or U19028 (N_19028,N_17167,N_16105);
or U19029 (N_19029,N_16858,N_17202);
nand U19030 (N_19030,N_17959,N_16480);
xnor U19031 (N_19031,N_16939,N_16846);
or U19032 (N_19032,N_17116,N_17986);
and U19033 (N_19033,N_17276,N_17930);
and U19034 (N_19034,N_17082,N_17970);
or U19035 (N_19035,N_16114,N_17938);
xor U19036 (N_19036,N_17708,N_17713);
and U19037 (N_19037,N_17886,N_17873);
or U19038 (N_19038,N_16012,N_17489);
nand U19039 (N_19039,N_16096,N_16357);
and U19040 (N_19040,N_17657,N_16862);
and U19041 (N_19041,N_16345,N_17194);
and U19042 (N_19042,N_16078,N_17346);
and U19043 (N_19043,N_17843,N_17946);
nand U19044 (N_19044,N_16973,N_16250);
nor U19045 (N_19045,N_17670,N_17620);
nor U19046 (N_19046,N_16479,N_17446);
nor U19047 (N_19047,N_17615,N_17971);
nor U19048 (N_19048,N_17827,N_17057);
nand U19049 (N_19049,N_16773,N_17764);
and U19050 (N_19050,N_17079,N_17537);
nand U19051 (N_19051,N_17864,N_17340);
and U19052 (N_19052,N_17119,N_16344);
or U19053 (N_19053,N_16631,N_16897);
and U19054 (N_19054,N_17083,N_16370);
and U19055 (N_19055,N_16089,N_16429);
or U19056 (N_19056,N_16541,N_17995);
or U19057 (N_19057,N_16329,N_17872);
or U19058 (N_19058,N_16217,N_16254);
xnor U19059 (N_19059,N_17742,N_16137);
xnor U19060 (N_19060,N_16506,N_16520);
nand U19061 (N_19061,N_16968,N_17150);
and U19062 (N_19062,N_16201,N_16625);
xnor U19063 (N_19063,N_16966,N_16424);
xnor U19064 (N_19064,N_16249,N_17988);
or U19065 (N_19065,N_16938,N_17916);
or U19066 (N_19066,N_16158,N_17967);
nand U19067 (N_19067,N_16698,N_17735);
and U19068 (N_19068,N_17174,N_17935);
or U19069 (N_19069,N_17087,N_16459);
nor U19070 (N_19070,N_17895,N_17304);
or U19071 (N_19071,N_16585,N_16381);
xor U19072 (N_19072,N_16789,N_17286);
nand U19073 (N_19073,N_17534,N_17909);
xor U19074 (N_19074,N_16810,N_17843);
nand U19075 (N_19075,N_17636,N_16258);
xor U19076 (N_19076,N_17895,N_16748);
xnor U19077 (N_19077,N_16380,N_16095);
and U19078 (N_19078,N_16529,N_17873);
xor U19079 (N_19079,N_16646,N_16984);
and U19080 (N_19080,N_17706,N_17713);
nor U19081 (N_19081,N_17133,N_17764);
xor U19082 (N_19082,N_16322,N_17014);
or U19083 (N_19083,N_16286,N_17206);
nand U19084 (N_19084,N_17584,N_17819);
nand U19085 (N_19085,N_16449,N_17918);
nor U19086 (N_19086,N_17277,N_17185);
and U19087 (N_19087,N_17809,N_16635);
or U19088 (N_19088,N_17494,N_17624);
xor U19089 (N_19089,N_16762,N_17168);
or U19090 (N_19090,N_17078,N_17464);
or U19091 (N_19091,N_16157,N_16312);
nand U19092 (N_19092,N_16642,N_17284);
or U19093 (N_19093,N_17999,N_16031);
nand U19094 (N_19094,N_16192,N_16706);
and U19095 (N_19095,N_17036,N_16041);
xor U19096 (N_19096,N_16821,N_16359);
nor U19097 (N_19097,N_17707,N_17206);
xnor U19098 (N_19098,N_16633,N_16981);
nor U19099 (N_19099,N_16679,N_17523);
and U19100 (N_19100,N_16732,N_16950);
nor U19101 (N_19101,N_16464,N_17804);
and U19102 (N_19102,N_17352,N_17250);
or U19103 (N_19103,N_16279,N_16632);
or U19104 (N_19104,N_16786,N_17441);
nand U19105 (N_19105,N_16273,N_16827);
and U19106 (N_19106,N_17107,N_17597);
xnor U19107 (N_19107,N_16524,N_17983);
or U19108 (N_19108,N_16907,N_16550);
xnor U19109 (N_19109,N_16876,N_16916);
xor U19110 (N_19110,N_17966,N_17215);
and U19111 (N_19111,N_16898,N_16275);
xnor U19112 (N_19112,N_16716,N_16056);
and U19113 (N_19113,N_16961,N_17724);
nor U19114 (N_19114,N_16835,N_16941);
nand U19115 (N_19115,N_16271,N_17724);
and U19116 (N_19116,N_17558,N_17060);
xnor U19117 (N_19117,N_17157,N_16774);
and U19118 (N_19118,N_16994,N_17721);
or U19119 (N_19119,N_16628,N_17683);
nand U19120 (N_19120,N_16139,N_17436);
nor U19121 (N_19121,N_16602,N_16292);
or U19122 (N_19122,N_16881,N_17969);
nor U19123 (N_19123,N_17772,N_16523);
xor U19124 (N_19124,N_16797,N_17244);
and U19125 (N_19125,N_17447,N_17736);
xnor U19126 (N_19126,N_17210,N_16684);
nand U19127 (N_19127,N_17153,N_17963);
xnor U19128 (N_19128,N_16705,N_17324);
nor U19129 (N_19129,N_17658,N_17748);
nand U19130 (N_19130,N_17116,N_16843);
nand U19131 (N_19131,N_17427,N_17089);
or U19132 (N_19132,N_17990,N_17154);
xor U19133 (N_19133,N_16063,N_16850);
nor U19134 (N_19134,N_17576,N_17354);
or U19135 (N_19135,N_17198,N_16350);
nor U19136 (N_19136,N_16490,N_17733);
xnor U19137 (N_19137,N_17153,N_17981);
and U19138 (N_19138,N_16427,N_17183);
nor U19139 (N_19139,N_16478,N_17966);
or U19140 (N_19140,N_16907,N_17048);
nor U19141 (N_19141,N_16283,N_17980);
and U19142 (N_19142,N_16192,N_16520);
and U19143 (N_19143,N_17003,N_17001);
nor U19144 (N_19144,N_17860,N_16814);
and U19145 (N_19145,N_16906,N_16871);
and U19146 (N_19146,N_17529,N_17161);
xnor U19147 (N_19147,N_16206,N_17413);
nand U19148 (N_19148,N_17356,N_17451);
nand U19149 (N_19149,N_17593,N_17445);
or U19150 (N_19150,N_17534,N_17391);
nor U19151 (N_19151,N_16925,N_16993);
and U19152 (N_19152,N_16336,N_17296);
nand U19153 (N_19153,N_17774,N_17928);
and U19154 (N_19154,N_16987,N_16841);
xor U19155 (N_19155,N_17604,N_17627);
nand U19156 (N_19156,N_17017,N_17575);
or U19157 (N_19157,N_17564,N_16483);
and U19158 (N_19158,N_17253,N_16905);
nor U19159 (N_19159,N_17650,N_16950);
nand U19160 (N_19160,N_16457,N_16514);
nand U19161 (N_19161,N_16668,N_16145);
nor U19162 (N_19162,N_16615,N_17938);
nor U19163 (N_19163,N_17190,N_17937);
nor U19164 (N_19164,N_17126,N_16246);
xor U19165 (N_19165,N_16280,N_17553);
and U19166 (N_19166,N_17479,N_16884);
nor U19167 (N_19167,N_17358,N_17999);
and U19168 (N_19168,N_17190,N_17706);
nor U19169 (N_19169,N_17160,N_17568);
or U19170 (N_19170,N_16521,N_16792);
nand U19171 (N_19171,N_17843,N_17884);
nor U19172 (N_19172,N_17564,N_16837);
xor U19173 (N_19173,N_17187,N_17278);
nand U19174 (N_19174,N_17193,N_17988);
and U19175 (N_19175,N_16051,N_16797);
xnor U19176 (N_19176,N_16155,N_16041);
nor U19177 (N_19177,N_17959,N_17437);
xnor U19178 (N_19178,N_16888,N_17165);
and U19179 (N_19179,N_17884,N_17707);
or U19180 (N_19180,N_16042,N_17274);
or U19181 (N_19181,N_17348,N_17566);
or U19182 (N_19182,N_16221,N_17977);
xnor U19183 (N_19183,N_17651,N_17174);
nand U19184 (N_19184,N_17650,N_17350);
or U19185 (N_19185,N_16779,N_17621);
and U19186 (N_19186,N_16749,N_16347);
and U19187 (N_19187,N_17470,N_16270);
xnor U19188 (N_19188,N_17963,N_16523);
xnor U19189 (N_19189,N_16546,N_17921);
and U19190 (N_19190,N_16519,N_16870);
nor U19191 (N_19191,N_16817,N_16803);
and U19192 (N_19192,N_16166,N_17819);
and U19193 (N_19193,N_16312,N_17454);
nand U19194 (N_19194,N_17544,N_17084);
and U19195 (N_19195,N_17931,N_17904);
nor U19196 (N_19196,N_17856,N_16926);
and U19197 (N_19197,N_17466,N_17317);
nand U19198 (N_19198,N_17175,N_17407);
xnor U19199 (N_19199,N_16273,N_16102);
nand U19200 (N_19200,N_17455,N_16982);
and U19201 (N_19201,N_17764,N_16915);
xnor U19202 (N_19202,N_17217,N_16220);
and U19203 (N_19203,N_17727,N_17617);
xor U19204 (N_19204,N_17245,N_17890);
and U19205 (N_19205,N_16590,N_17649);
or U19206 (N_19206,N_17879,N_16188);
nand U19207 (N_19207,N_17571,N_17962);
xor U19208 (N_19208,N_17879,N_16434);
and U19209 (N_19209,N_17895,N_17818);
or U19210 (N_19210,N_17084,N_16940);
and U19211 (N_19211,N_17305,N_17509);
and U19212 (N_19212,N_16582,N_17695);
and U19213 (N_19213,N_17910,N_17037);
or U19214 (N_19214,N_16670,N_16343);
nor U19215 (N_19215,N_16600,N_16350);
and U19216 (N_19216,N_16308,N_16411);
nand U19217 (N_19217,N_17758,N_16456);
and U19218 (N_19218,N_17123,N_16162);
and U19219 (N_19219,N_17398,N_17721);
nand U19220 (N_19220,N_16260,N_17034);
or U19221 (N_19221,N_17941,N_16786);
nor U19222 (N_19222,N_17269,N_16452);
xnor U19223 (N_19223,N_17679,N_16474);
or U19224 (N_19224,N_17516,N_16213);
nand U19225 (N_19225,N_17317,N_17404);
and U19226 (N_19226,N_16770,N_17662);
and U19227 (N_19227,N_16909,N_17059);
or U19228 (N_19228,N_17812,N_16076);
nand U19229 (N_19229,N_16364,N_16678);
xnor U19230 (N_19230,N_17989,N_17880);
and U19231 (N_19231,N_16862,N_17801);
and U19232 (N_19232,N_17471,N_17211);
and U19233 (N_19233,N_17179,N_16931);
or U19234 (N_19234,N_17714,N_17082);
nor U19235 (N_19235,N_17799,N_16946);
xnor U19236 (N_19236,N_17418,N_17043);
or U19237 (N_19237,N_17423,N_16809);
xnor U19238 (N_19238,N_16896,N_17434);
and U19239 (N_19239,N_17077,N_17343);
xnor U19240 (N_19240,N_17739,N_16610);
nand U19241 (N_19241,N_16966,N_17309);
and U19242 (N_19242,N_16155,N_16270);
and U19243 (N_19243,N_16606,N_16908);
or U19244 (N_19244,N_16167,N_17250);
nand U19245 (N_19245,N_17866,N_17251);
nor U19246 (N_19246,N_17172,N_16386);
nor U19247 (N_19247,N_16944,N_17122);
or U19248 (N_19248,N_17450,N_16941);
and U19249 (N_19249,N_17951,N_16453);
nand U19250 (N_19250,N_17135,N_17039);
nor U19251 (N_19251,N_16767,N_16331);
nor U19252 (N_19252,N_17637,N_17653);
xor U19253 (N_19253,N_17102,N_17850);
or U19254 (N_19254,N_16239,N_17311);
or U19255 (N_19255,N_16098,N_17304);
nor U19256 (N_19256,N_16429,N_16096);
and U19257 (N_19257,N_17685,N_17778);
and U19258 (N_19258,N_16397,N_16922);
or U19259 (N_19259,N_16864,N_16631);
and U19260 (N_19260,N_17903,N_16862);
or U19261 (N_19261,N_16869,N_17511);
or U19262 (N_19262,N_16230,N_16012);
nand U19263 (N_19263,N_16872,N_16020);
nor U19264 (N_19264,N_16949,N_16606);
nor U19265 (N_19265,N_17200,N_17712);
or U19266 (N_19266,N_16334,N_16708);
or U19267 (N_19267,N_17780,N_17039);
or U19268 (N_19268,N_16127,N_16418);
xnor U19269 (N_19269,N_17545,N_17979);
and U19270 (N_19270,N_16378,N_17397);
and U19271 (N_19271,N_17672,N_17803);
xnor U19272 (N_19272,N_17793,N_17783);
or U19273 (N_19273,N_16186,N_17524);
xnor U19274 (N_19274,N_16911,N_17320);
nor U19275 (N_19275,N_16445,N_16797);
nor U19276 (N_19276,N_17203,N_16051);
or U19277 (N_19277,N_17825,N_17640);
nor U19278 (N_19278,N_17963,N_17044);
nor U19279 (N_19279,N_17283,N_16117);
and U19280 (N_19280,N_16415,N_17476);
nand U19281 (N_19281,N_17059,N_17109);
or U19282 (N_19282,N_17145,N_16630);
nand U19283 (N_19283,N_16904,N_16697);
nor U19284 (N_19284,N_16508,N_16606);
nand U19285 (N_19285,N_16434,N_16164);
nor U19286 (N_19286,N_16955,N_17139);
nand U19287 (N_19287,N_16241,N_17221);
nor U19288 (N_19288,N_17148,N_16850);
or U19289 (N_19289,N_16952,N_17629);
and U19290 (N_19290,N_16362,N_16035);
nand U19291 (N_19291,N_17837,N_17025);
xnor U19292 (N_19292,N_16112,N_17847);
xor U19293 (N_19293,N_16707,N_16088);
nand U19294 (N_19294,N_16083,N_16027);
nand U19295 (N_19295,N_17681,N_16823);
nand U19296 (N_19296,N_17671,N_16741);
and U19297 (N_19297,N_17237,N_17088);
or U19298 (N_19298,N_16780,N_17987);
nand U19299 (N_19299,N_16194,N_17851);
and U19300 (N_19300,N_17635,N_17156);
xnor U19301 (N_19301,N_16615,N_17055);
or U19302 (N_19302,N_17309,N_16503);
xnor U19303 (N_19303,N_16547,N_16469);
and U19304 (N_19304,N_16956,N_17393);
and U19305 (N_19305,N_16731,N_16409);
nand U19306 (N_19306,N_17463,N_17716);
nor U19307 (N_19307,N_16862,N_17016);
and U19308 (N_19308,N_17845,N_16212);
and U19309 (N_19309,N_17269,N_17679);
or U19310 (N_19310,N_17745,N_16818);
and U19311 (N_19311,N_17916,N_17439);
xnor U19312 (N_19312,N_17344,N_16384);
xnor U19313 (N_19313,N_17724,N_16451);
nand U19314 (N_19314,N_16933,N_16156);
nor U19315 (N_19315,N_16874,N_17722);
and U19316 (N_19316,N_16078,N_16828);
and U19317 (N_19317,N_17299,N_16620);
or U19318 (N_19318,N_17082,N_16903);
or U19319 (N_19319,N_17276,N_17539);
and U19320 (N_19320,N_17743,N_16927);
or U19321 (N_19321,N_16025,N_16668);
nand U19322 (N_19322,N_16522,N_16806);
nor U19323 (N_19323,N_17528,N_17314);
or U19324 (N_19324,N_16572,N_16334);
nor U19325 (N_19325,N_16611,N_16766);
and U19326 (N_19326,N_17311,N_17664);
or U19327 (N_19327,N_16500,N_16666);
xnor U19328 (N_19328,N_16565,N_17574);
and U19329 (N_19329,N_16185,N_16665);
and U19330 (N_19330,N_16904,N_16253);
or U19331 (N_19331,N_17651,N_16870);
or U19332 (N_19332,N_17939,N_17170);
nand U19333 (N_19333,N_17493,N_16262);
or U19334 (N_19334,N_16805,N_16711);
nor U19335 (N_19335,N_16961,N_16299);
nor U19336 (N_19336,N_17316,N_17526);
nor U19337 (N_19337,N_16907,N_16173);
nor U19338 (N_19338,N_16734,N_16426);
and U19339 (N_19339,N_16622,N_17174);
and U19340 (N_19340,N_16599,N_16937);
xor U19341 (N_19341,N_17478,N_17720);
xnor U19342 (N_19342,N_17074,N_16179);
nand U19343 (N_19343,N_17733,N_17636);
nand U19344 (N_19344,N_16265,N_17201);
nor U19345 (N_19345,N_16940,N_16630);
xnor U19346 (N_19346,N_17838,N_17645);
nor U19347 (N_19347,N_16173,N_17869);
nor U19348 (N_19348,N_16977,N_17459);
and U19349 (N_19349,N_16881,N_16097);
nand U19350 (N_19350,N_17484,N_17194);
xnor U19351 (N_19351,N_16518,N_16574);
or U19352 (N_19352,N_17981,N_17711);
and U19353 (N_19353,N_17082,N_17769);
nand U19354 (N_19354,N_17774,N_17006);
nor U19355 (N_19355,N_16159,N_17218);
nand U19356 (N_19356,N_16856,N_16429);
nand U19357 (N_19357,N_16093,N_17014);
xor U19358 (N_19358,N_16739,N_16419);
xor U19359 (N_19359,N_16204,N_16806);
xor U19360 (N_19360,N_16619,N_17941);
or U19361 (N_19361,N_17576,N_17097);
xor U19362 (N_19362,N_16996,N_16666);
xor U19363 (N_19363,N_16607,N_17031);
nand U19364 (N_19364,N_16391,N_17387);
nor U19365 (N_19365,N_17244,N_16936);
nor U19366 (N_19366,N_16642,N_16608);
nor U19367 (N_19367,N_16869,N_17745);
or U19368 (N_19368,N_17012,N_17690);
or U19369 (N_19369,N_16578,N_17816);
or U19370 (N_19370,N_16123,N_17763);
nand U19371 (N_19371,N_17041,N_17206);
nand U19372 (N_19372,N_17068,N_16523);
or U19373 (N_19373,N_17165,N_17598);
nor U19374 (N_19374,N_17848,N_16923);
xnor U19375 (N_19375,N_17333,N_16606);
or U19376 (N_19376,N_16113,N_17462);
and U19377 (N_19377,N_16278,N_17892);
and U19378 (N_19378,N_17111,N_16993);
xnor U19379 (N_19379,N_16344,N_17893);
or U19380 (N_19380,N_16262,N_16744);
or U19381 (N_19381,N_17555,N_16627);
nor U19382 (N_19382,N_16094,N_17692);
or U19383 (N_19383,N_17374,N_17483);
or U19384 (N_19384,N_17027,N_17743);
or U19385 (N_19385,N_16341,N_16019);
or U19386 (N_19386,N_16690,N_16387);
nand U19387 (N_19387,N_17614,N_16421);
and U19388 (N_19388,N_16070,N_17655);
or U19389 (N_19389,N_17160,N_16420);
and U19390 (N_19390,N_16474,N_17750);
xnor U19391 (N_19391,N_16022,N_16054);
nand U19392 (N_19392,N_17887,N_16345);
nand U19393 (N_19393,N_16452,N_16509);
and U19394 (N_19394,N_17064,N_17374);
xnor U19395 (N_19395,N_17966,N_16939);
xnor U19396 (N_19396,N_17480,N_16457);
and U19397 (N_19397,N_16810,N_16140);
and U19398 (N_19398,N_16895,N_16016);
and U19399 (N_19399,N_17039,N_17093);
and U19400 (N_19400,N_16519,N_17995);
nor U19401 (N_19401,N_17084,N_16693);
nor U19402 (N_19402,N_16667,N_16498);
and U19403 (N_19403,N_16392,N_17881);
and U19404 (N_19404,N_17209,N_17993);
nor U19405 (N_19405,N_16926,N_17942);
or U19406 (N_19406,N_16484,N_16245);
xnor U19407 (N_19407,N_17203,N_17173);
xor U19408 (N_19408,N_16223,N_16459);
and U19409 (N_19409,N_16146,N_17732);
and U19410 (N_19410,N_16068,N_16186);
and U19411 (N_19411,N_17437,N_17182);
nor U19412 (N_19412,N_17668,N_17886);
nand U19413 (N_19413,N_17283,N_16248);
nor U19414 (N_19414,N_16967,N_17825);
and U19415 (N_19415,N_16616,N_16662);
nand U19416 (N_19416,N_16409,N_17395);
or U19417 (N_19417,N_16154,N_16405);
nand U19418 (N_19418,N_17555,N_16923);
nand U19419 (N_19419,N_17961,N_17429);
and U19420 (N_19420,N_17799,N_17388);
nor U19421 (N_19421,N_17145,N_17200);
or U19422 (N_19422,N_16641,N_17388);
nand U19423 (N_19423,N_17252,N_17607);
and U19424 (N_19424,N_16148,N_16714);
nor U19425 (N_19425,N_16834,N_17643);
nand U19426 (N_19426,N_17672,N_17086);
or U19427 (N_19427,N_17622,N_17566);
or U19428 (N_19428,N_17943,N_16955);
or U19429 (N_19429,N_16708,N_16185);
nor U19430 (N_19430,N_16555,N_17357);
and U19431 (N_19431,N_16574,N_17866);
nand U19432 (N_19432,N_16551,N_17289);
nand U19433 (N_19433,N_17982,N_16158);
xor U19434 (N_19434,N_17588,N_17641);
nand U19435 (N_19435,N_16247,N_16444);
xor U19436 (N_19436,N_17618,N_16459);
nand U19437 (N_19437,N_17159,N_17381);
or U19438 (N_19438,N_17633,N_16129);
or U19439 (N_19439,N_16266,N_17741);
nand U19440 (N_19440,N_17902,N_16205);
nand U19441 (N_19441,N_16114,N_17204);
xor U19442 (N_19442,N_16921,N_17302);
and U19443 (N_19443,N_17006,N_17715);
xnor U19444 (N_19444,N_16731,N_16624);
nor U19445 (N_19445,N_17093,N_17178);
and U19446 (N_19446,N_17292,N_16979);
nor U19447 (N_19447,N_16228,N_16520);
nor U19448 (N_19448,N_17969,N_17625);
or U19449 (N_19449,N_17706,N_17819);
or U19450 (N_19450,N_17988,N_16356);
and U19451 (N_19451,N_17199,N_16304);
nand U19452 (N_19452,N_17474,N_16215);
or U19453 (N_19453,N_16932,N_17716);
and U19454 (N_19454,N_16889,N_16073);
nor U19455 (N_19455,N_16935,N_17535);
xnor U19456 (N_19456,N_17101,N_17258);
and U19457 (N_19457,N_17738,N_16263);
nand U19458 (N_19458,N_16420,N_17455);
nand U19459 (N_19459,N_17273,N_17938);
nand U19460 (N_19460,N_16287,N_17786);
or U19461 (N_19461,N_16496,N_16310);
nand U19462 (N_19462,N_17341,N_17567);
xnor U19463 (N_19463,N_17475,N_17053);
nor U19464 (N_19464,N_16963,N_16909);
xnor U19465 (N_19465,N_17816,N_16400);
or U19466 (N_19466,N_16428,N_16944);
or U19467 (N_19467,N_17466,N_17998);
nand U19468 (N_19468,N_16726,N_16774);
xnor U19469 (N_19469,N_17682,N_17349);
and U19470 (N_19470,N_16466,N_16217);
and U19471 (N_19471,N_17661,N_17138);
and U19472 (N_19472,N_17166,N_16064);
xor U19473 (N_19473,N_16603,N_17221);
or U19474 (N_19474,N_17393,N_16159);
nor U19475 (N_19475,N_17265,N_16367);
and U19476 (N_19476,N_17423,N_16567);
and U19477 (N_19477,N_16468,N_17470);
nand U19478 (N_19478,N_17948,N_16615);
xnor U19479 (N_19479,N_17872,N_17224);
nand U19480 (N_19480,N_17930,N_17580);
nand U19481 (N_19481,N_17563,N_16423);
nand U19482 (N_19482,N_16537,N_17230);
xor U19483 (N_19483,N_17498,N_16622);
nand U19484 (N_19484,N_16657,N_17225);
nor U19485 (N_19485,N_16754,N_16682);
nor U19486 (N_19486,N_16710,N_17842);
xor U19487 (N_19487,N_16041,N_16700);
xnor U19488 (N_19488,N_16005,N_17194);
or U19489 (N_19489,N_17808,N_17509);
xnor U19490 (N_19490,N_17274,N_16297);
or U19491 (N_19491,N_17875,N_16481);
nand U19492 (N_19492,N_16077,N_16277);
and U19493 (N_19493,N_16703,N_17195);
xnor U19494 (N_19494,N_16253,N_16441);
and U19495 (N_19495,N_17841,N_16217);
xor U19496 (N_19496,N_17968,N_17834);
or U19497 (N_19497,N_16162,N_16632);
or U19498 (N_19498,N_17840,N_17907);
nand U19499 (N_19499,N_16661,N_17229);
and U19500 (N_19500,N_17649,N_16264);
nor U19501 (N_19501,N_16243,N_17409);
nor U19502 (N_19502,N_16737,N_17842);
nand U19503 (N_19503,N_17790,N_17541);
xor U19504 (N_19504,N_17263,N_16823);
nand U19505 (N_19505,N_17784,N_16468);
xor U19506 (N_19506,N_16291,N_17946);
or U19507 (N_19507,N_16436,N_16332);
nor U19508 (N_19508,N_16823,N_16962);
nor U19509 (N_19509,N_16434,N_17391);
and U19510 (N_19510,N_16118,N_16841);
and U19511 (N_19511,N_16772,N_17626);
or U19512 (N_19512,N_16341,N_17385);
and U19513 (N_19513,N_16608,N_17819);
nand U19514 (N_19514,N_17051,N_16711);
xor U19515 (N_19515,N_16680,N_16179);
and U19516 (N_19516,N_16774,N_17551);
nand U19517 (N_19517,N_16866,N_17269);
nor U19518 (N_19518,N_16499,N_17871);
xnor U19519 (N_19519,N_17200,N_16880);
nor U19520 (N_19520,N_16394,N_16832);
or U19521 (N_19521,N_16420,N_17781);
or U19522 (N_19522,N_16195,N_16726);
xnor U19523 (N_19523,N_16347,N_17436);
nand U19524 (N_19524,N_17991,N_17586);
or U19525 (N_19525,N_16725,N_16275);
nand U19526 (N_19526,N_16087,N_16220);
nor U19527 (N_19527,N_16118,N_17251);
nand U19528 (N_19528,N_16795,N_17143);
nand U19529 (N_19529,N_16803,N_17808);
xor U19530 (N_19530,N_17485,N_17974);
or U19531 (N_19531,N_16970,N_16203);
or U19532 (N_19532,N_16072,N_17335);
or U19533 (N_19533,N_16618,N_17491);
nor U19534 (N_19534,N_16678,N_17442);
and U19535 (N_19535,N_16569,N_17424);
or U19536 (N_19536,N_17420,N_17089);
and U19537 (N_19537,N_16482,N_17438);
nor U19538 (N_19538,N_17579,N_17721);
or U19539 (N_19539,N_17360,N_16341);
and U19540 (N_19540,N_16864,N_16897);
nor U19541 (N_19541,N_17758,N_17494);
or U19542 (N_19542,N_16968,N_17923);
xnor U19543 (N_19543,N_17104,N_16580);
nor U19544 (N_19544,N_17876,N_17610);
nor U19545 (N_19545,N_16092,N_17077);
and U19546 (N_19546,N_17406,N_16033);
nor U19547 (N_19547,N_17576,N_17256);
and U19548 (N_19548,N_16295,N_16720);
nor U19549 (N_19549,N_17184,N_17826);
or U19550 (N_19550,N_16176,N_17186);
xnor U19551 (N_19551,N_17257,N_16941);
xnor U19552 (N_19552,N_16792,N_17986);
xor U19553 (N_19553,N_16485,N_17156);
nor U19554 (N_19554,N_17125,N_17776);
xor U19555 (N_19555,N_17454,N_16320);
nand U19556 (N_19556,N_16570,N_17388);
nor U19557 (N_19557,N_17554,N_17794);
nor U19558 (N_19558,N_17429,N_17726);
or U19559 (N_19559,N_16324,N_16296);
and U19560 (N_19560,N_16969,N_16118);
xnor U19561 (N_19561,N_17741,N_17426);
or U19562 (N_19562,N_17593,N_16492);
nand U19563 (N_19563,N_17547,N_17172);
nand U19564 (N_19564,N_17623,N_16861);
and U19565 (N_19565,N_16748,N_16374);
and U19566 (N_19566,N_17312,N_17422);
nand U19567 (N_19567,N_16586,N_16175);
or U19568 (N_19568,N_17426,N_16143);
nor U19569 (N_19569,N_16241,N_17816);
nand U19570 (N_19570,N_16903,N_17927);
nand U19571 (N_19571,N_17429,N_16370);
nor U19572 (N_19572,N_17987,N_16745);
nor U19573 (N_19573,N_16960,N_17098);
or U19574 (N_19574,N_17841,N_16932);
and U19575 (N_19575,N_17532,N_17273);
nor U19576 (N_19576,N_17912,N_16213);
nor U19577 (N_19577,N_17236,N_17776);
or U19578 (N_19578,N_16574,N_17118);
xnor U19579 (N_19579,N_16129,N_17485);
nand U19580 (N_19580,N_17743,N_17738);
nand U19581 (N_19581,N_17432,N_16173);
and U19582 (N_19582,N_17605,N_17515);
xor U19583 (N_19583,N_17390,N_17955);
or U19584 (N_19584,N_17639,N_16261);
nand U19585 (N_19585,N_16997,N_16434);
nor U19586 (N_19586,N_16537,N_16327);
and U19587 (N_19587,N_17489,N_17885);
and U19588 (N_19588,N_16420,N_16544);
xnor U19589 (N_19589,N_16131,N_16925);
and U19590 (N_19590,N_17334,N_17077);
nor U19591 (N_19591,N_17968,N_17298);
nor U19592 (N_19592,N_17697,N_16603);
nand U19593 (N_19593,N_16541,N_17537);
or U19594 (N_19594,N_16896,N_17980);
xnor U19595 (N_19595,N_16117,N_17083);
and U19596 (N_19596,N_16495,N_16150);
and U19597 (N_19597,N_16675,N_16562);
xnor U19598 (N_19598,N_16050,N_16447);
nand U19599 (N_19599,N_16546,N_16626);
nand U19600 (N_19600,N_16486,N_17124);
and U19601 (N_19601,N_16804,N_17140);
xnor U19602 (N_19602,N_17566,N_16759);
or U19603 (N_19603,N_17878,N_17154);
nand U19604 (N_19604,N_16030,N_17773);
nor U19605 (N_19605,N_17788,N_16794);
and U19606 (N_19606,N_17956,N_16288);
nand U19607 (N_19607,N_17706,N_17877);
nand U19608 (N_19608,N_17041,N_17720);
nor U19609 (N_19609,N_16145,N_16665);
xnor U19610 (N_19610,N_17989,N_17469);
or U19611 (N_19611,N_17406,N_17358);
and U19612 (N_19612,N_17407,N_17279);
nand U19613 (N_19613,N_17536,N_17581);
or U19614 (N_19614,N_16212,N_16362);
or U19615 (N_19615,N_17618,N_17652);
and U19616 (N_19616,N_17401,N_16109);
nor U19617 (N_19617,N_16263,N_17519);
or U19618 (N_19618,N_17101,N_16751);
or U19619 (N_19619,N_16322,N_17224);
or U19620 (N_19620,N_16335,N_16976);
or U19621 (N_19621,N_17024,N_17334);
or U19622 (N_19622,N_17413,N_16036);
or U19623 (N_19623,N_16438,N_16063);
and U19624 (N_19624,N_16316,N_16526);
and U19625 (N_19625,N_16045,N_16255);
and U19626 (N_19626,N_16436,N_17395);
xor U19627 (N_19627,N_16656,N_17376);
xnor U19628 (N_19628,N_17746,N_16075);
and U19629 (N_19629,N_17570,N_17407);
or U19630 (N_19630,N_17699,N_16940);
and U19631 (N_19631,N_16366,N_16634);
xnor U19632 (N_19632,N_16761,N_17195);
and U19633 (N_19633,N_17866,N_17388);
xnor U19634 (N_19634,N_16194,N_16802);
nor U19635 (N_19635,N_17703,N_17422);
and U19636 (N_19636,N_17378,N_17244);
nand U19637 (N_19637,N_16120,N_17369);
xnor U19638 (N_19638,N_16701,N_16374);
nor U19639 (N_19639,N_16111,N_16881);
nor U19640 (N_19640,N_16598,N_16926);
xor U19641 (N_19641,N_16273,N_17507);
xnor U19642 (N_19642,N_16467,N_16319);
or U19643 (N_19643,N_17827,N_17654);
and U19644 (N_19644,N_16356,N_17342);
and U19645 (N_19645,N_17976,N_16961);
or U19646 (N_19646,N_16327,N_16829);
nand U19647 (N_19647,N_16217,N_16575);
nand U19648 (N_19648,N_17038,N_17968);
nor U19649 (N_19649,N_16758,N_17970);
xnor U19650 (N_19650,N_17442,N_17410);
and U19651 (N_19651,N_17604,N_16223);
xnor U19652 (N_19652,N_17355,N_17517);
nor U19653 (N_19653,N_17060,N_16681);
and U19654 (N_19654,N_16645,N_16176);
xor U19655 (N_19655,N_16227,N_17902);
xnor U19656 (N_19656,N_16128,N_17605);
xor U19657 (N_19657,N_17399,N_16231);
nor U19658 (N_19658,N_16216,N_16646);
and U19659 (N_19659,N_17490,N_17533);
xnor U19660 (N_19660,N_17263,N_17143);
nor U19661 (N_19661,N_17641,N_17853);
or U19662 (N_19662,N_16252,N_16088);
or U19663 (N_19663,N_17628,N_16021);
nor U19664 (N_19664,N_16551,N_17603);
xnor U19665 (N_19665,N_16191,N_16820);
nand U19666 (N_19666,N_17055,N_16046);
and U19667 (N_19667,N_17417,N_16231);
and U19668 (N_19668,N_17973,N_17922);
xnor U19669 (N_19669,N_17024,N_16815);
xnor U19670 (N_19670,N_16477,N_16517);
nand U19671 (N_19671,N_16286,N_17898);
or U19672 (N_19672,N_17126,N_17816);
nor U19673 (N_19673,N_17330,N_16559);
nor U19674 (N_19674,N_17005,N_17152);
nand U19675 (N_19675,N_16616,N_16583);
nand U19676 (N_19676,N_17419,N_16356);
nor U19677 (N_19677,N_17694,N_17735);
xnor U19678 (N_19678,N_16974,N_16861);
or U19679 (N_19679,N_17937,N_16899);
or U19680 (N_19680,N_17924,N_17787);
nand U19681 (N_19681,N_17079,N_17183);
or U19682 (N_19682,N_16219,N_16903);
and U19683 (N_19683,N_16120,N_16060);
nand U19684 (N_19684,N_16648,N_16566);
xnor U19685 (N_19685,N_16862,N_16799);
or U19686 (N_19686,N_17548,N_16859);
nand U19687 (N_19687,N_17784,N_17378);
xnor U19688 (N_19688,N_17333,N_16309);
or U19689 (N_19689,N_17816,N_16885);
or U19690 (N_19690,N_16197,N_17392);
nand U19691 (N_19691,N_17970,N_16525);
nor U19692 (N_19692,N_17803,N_16203);
xnor U19693 (N_19693,N_17287,N_16702);
and U19694 (N_19694,N_17022,N_16248);
nand U19695 (N_19695,N_16027,N_17666);
and U19696 (N_19696,N_17970,N_17629);
nor U19697 (N_19697,N_16049,N_16925);
nand U19698 (N_19698,N_17161,N_17194);
nand U19699 (N_19699,N_16111,N_17457);
nand U19700 (N_19700,N_17982,N_16378);
nand U19701 (N_19701,N_16690,N_16722);
nor U19702 (N_19702,N_17058,N_17266);
or U19703 (N_19703,N_17594,N_16160);
and U19704 (N_19704,N_17711,N_17669);
and U19705 (N_19705,N_16891,N_16274);
xnor U19706 (N_19706,N_17012,N_16002);
nor U19707 (N_19707,N_17596,N_16751);
or U19708 (N_19708,N_16246,N_17731);
nand U19709 (N_19709,N_16675,N_16412);
xnor U19710 (N_19710,N_17507,N_16681);
nand U19711 (N_19711,N_17566,N_17854);
xor U19712 (N_19712,N_16839,N_17838);
nand U19713 (N_19713,N_16686,N_17559);
or U19714 (N_19714,N_17600,N_17256);
and U19715 (N_19715,N_16495,N_17758);
xor U19716 (N_19716,N_16714,N_17610);
xnor U19717 (N_19717,N_16253,N_16388);
and U19718 (N_19718,N_17316,N_17309);
nand U19719 (N_19719,N_17803,N_16320);
xnor U19720 (N_19720,N_16291,N_17587);
nor U19721 (N_19721,N_17916,N_16081);
nand U19722 (N_19722,N_17624,N_16685);
nor U19723 (N_19723,N_16280,N_16922);
or U19724 (N_19724,N_17979,N_17711);
nor U19725 (N_19725,N_17257,N_17283);
or U19726 (N_19726,N_16520,N_16023);
nand U19727 (N_19727,N_17641,N_17075);
and U19728 (N_19728,N_16882,N_17930);
nand U19729 (N_19729,N_17656,N_16863);
and U19730 (N_19730,N_16727,N_16105);
and U19731 (N_19731,N_17813,N_17343);
xnor U19732 (N_19732,N_17348,N_17246);
nand U19733 (N_19733,N_17478,N_16794);
or U19734 (N_19734,N_16129,N_17908);
nor U19735 (N_19735,N_17920,N_17680);
nand U19736 (N_19736,N_17559,N_16952);
and U19737 (N_19737,N_16193,N_17413);
or U19738 (N_19738,N_17577,N_16711);
nor U19739 (N_19739,N_17671,N_16261);
and U19740 (N_19740,N_17926,N_16375);
and U19741 (N_19741,N_17939,N_16666);
nor U19742 (N_19742,N_17889,N_17924);
nand U19743 (N_19743,N_16384,N_17723);
xor U19744 (N_19744,N_16799,N_17371);
nand U19745 (N_19745,N_16708,N_16913);
xor U19746 (N_19746,N_17323,N_16574);
and U19747 (N_19747,N_17918,N_17968);
and U19748 (N_19748,N_17543,N_16542);
nor U19749 (N_19749,N_17674,N_17738);
nand U19750 (N_19750,N_16303,N_17761);
xnor U19751 (N_19751,N_16789,N_17988);
xnor U19752 (N_19752,N_17789,N_16935);
nor U19753 (N_19753,N_17587,N_16124);
and U19754 (N_19754,N_17637,N_17175);
and U19755 (N_19755,N_16336,N_17745);
nor U19756 (N_19756,N_17768,N_17836);
or U19757 (N_19757,N_17309,N_17131);
and U19758 (N_19758,N_17912,N_17966);
xor U19759 (N_19759,N_16540,N_16944);
xnor U19760 (N_19760,N_17568,N_17547);
xor U19761 (N_19761,N_16410,N_16368);
xor U19762 (N_19762,N_16174,N_16543);
nand U19763 (N_19763,N_16194,N_17165);
nor U19764 (N_19764,N_16590,N_16577);
nor U19765 (N_19765,N_16015,N_17038);
nand U19766 (N_19766,N_16245,N_17131);
or U19767 (N_19767,N_16452,N_16665);
xor U19768 (N_19768,N_17625,N_17421);
or U19769 (N_19769,N_16835,N_16962);
xor U19770 (N_19770,N_16131,N_16962);
and U19771 (N_19771,N_16713,N_17898);
xnor U19772 (N_19772,N_17416,N_16552);
nor U19773 (N_19773,N_17413,N_16784);
nand U19774 (N_19774,N_16126,N_17082);
xnor U19775 (N_19775,N_17471,N_17221);
xor U19776 (N_19776,N_17571,N_16892);
nor U19777 (N_19777,N_17237,N_17923);
and U19778 (N_19778,N_16108,N_17448);
xnor U19779 (N_19779,N_17985,N_16604);
or U19780 (N_19780,N_17804,N_17176);
and U19781 (N_19781,N_16375,N_16200);
nor U19782 (N_19782,N_17390,N_17393);
xor U19783 (N_19783,N_16140,N_17443);
nor U19784 (N_19784,N_16264,N_16649);
or U19785 (N_19785,N_16948,N_17302);
or U19786 (N_19786,N_17114,N_16808);
and U19787 (N_19787,N_16977,N_16720);
or U19788 (N_19788,N_16085,N_16694);
nand U19789 (N_19789,N_17457,N_17699);
nand U19790 (N_19790,N_16351,N_17686);
and U19791 (N_19791,N_16240,N_16336);
or U19792 (N_19792,N_17391,N_17325);
or U19793 (N_19793,N_16705,N_16377);
xnor U19794 (N_19794,N_17983,N_16635);
xor U19795 (N_19795,N_17507,N_17376);
or U19796 (N_19796,N_17871,N_16422);
nand U19797 (N_19797,N_16974,N_17923);
nand U19798 (N_19798,N_16136,N_16106);
nand U19799 (N_19799,N_17721,N_16449);
nand U19800 (N_19800,N_17273,N_16797);
nand U19801 (N_19801,N_17985,N_17730);
nor U19802 (N_19802,N_17868,N_16810);
and U19803 (N_19803,N_16442,N_17104);
xor U19804 (N_19804,N_17210,N_17074);
nor U19805 (N_19805,N_16529,N_17480);
nor U19806 (N_19806,N_16989,N_16072);
xor U19807 (N_19807,N_16653,N_17673);
xor U19808 (N_19808,N_16831,N_16304);
nand U19809 (N_19809,N_17300,N_16099);
nand U19810 (N_19810,N_16158,N_16058);
nand U19811 (N_19811,N_17568,N_17257);
nor U19812 (N_19812,N_17376,N_16895);
nor U19813 (N_19813,N_16113,N_16449);
nor U19814 (N_19814,N_17060,N_17435);
xor U19815 (N_19815,N_16191,N_17055);
and U19816 (N_19816,N_16650,N_16482);
or U19817 (N_19817,N_16612,N_17830);
nand U19818 (N_19818,N_16041,N_17162);
and U19819 (N_19819,N_16185,N_17432);
or U19820 (N_19820,N_16574,N_17651);
nor U19821 (N_19821,N_17597,N_17803);
or U19822 (N_19822,N_17166,N_16419);
and U19823 (N_19823,N_17824,N_16628);
and U19824 (N_19824,N_17521,N_16090);
nand U19825 (N_19825,N_17252,N_17957);
nor U19826 (N_19826,N_16018,N_17335);
xor U19827 (N_19827,N_16220,N_17143);
and U19828 (N_19828,N_16350,N_17042);
xor U19829 (N_19829,N_16226,N_16921);
nand U19830 (N_19830,N_17832,N_17509);
and U19831 (N_19831,N_17653,N_16249);
nand U19832 (N_19832,N_16984,N_17841);
xor U19833 (N_19833,N_16592,N_17950);
nand U19834 (N_19834,N_16445,N_17376);
or U19835 (N_19835,N_17437,N_17410);
and U19836 (N_19836,N_17461,N_17735);
nand U19837 (N_19837,N_17323,N_16533);
nor U19838 (N_19838,N_17216,N_16078);
or U19839 (N_19839,N_16531,N_17977);
nor U19840 (N_19840,N_16390,N_16023);
nor U19841 (N_19841,N_16379,N_16276);
and U19842 (N_19842,N_16394,N_16303);
nand U19843 (N_19843,N_16370,N_17187);
xor U19844 (N_19844,N_17182,N_16392);
nor U19845 (N_19845,N_17577,N_17203);
nor U19846 (N_19846,N_17083,N_16161);
nand U19847 (N_19847,N_16896,N_17498);
and U19848 (N_19848,N_16461,N_17571);
and U19849 (N_19849,N_16409,N_16768);
or U19850 (N_19850,N_16933,N_17780);
or U19851 (N_19851,N_17081,N_16544);
xnor U19852 (N_19852,N_16364,N_17442);
and U19853 (N_19853,N_17381,N_17195);
xnor U19854 (N_19854,N_17927,N_16631);
nand U19855 (N_19855,N_17770,N_16617);
or U19856 (N_19856,N_17356,N_16854);
nor U19857 (N_19857,N_16321,N_17683);
and U19858 (N_19858,N_16250,N_17983);
or U19859 (N_19859,N_17871,N_17472);
or U19860 (N_19860,N_17307,N_16979);
xnor U19861 (N_19861,N_16988,N_17320);
nand U19862 (N_19862,N_17005,N_16237);
xor U19863 (N_19863,N_17296,N_17907);
or U19864 (N_19864,N_16758,N_17849);
xnor U19865 (N_19865,N_16036,N_17287);
and U19866 (N_19866,N_16357,N_17988);
and U19867 (N_19867,N_17610,N_16892);
nor U19868 (N_19868,N_16072,N_17609);
nand U19869 (N_19869,N_17911,N_17011);
xor U19870 (N_19870,N_17188,N_16451);
or U19871 (N_19871,N_17908,N_17233);
nor U19872 (N_19872,N_17103,N_16119);
xnor U19873 (N_19873,N_17560,N_17824);
and U19874 (N_19874,N_17385,N_17583);
xor U19875 (N_19875,N_17272,N_16470);
or U19876 (N_19876,N_17936,N_16773);
and U19877 (N_19877,N_17750,N_16633);
or U19878 (N_19878,N_17312,N_17878);
or U19879 (N_19879,N_17151,N_16841);
nand U19880 (N_19880,N_17268,N_17389);
nand U19881 (N_19881,N_16455,N_17715);
nor U19882 (N_19882,N_16914,N_17587);
and U19883 (N_19883,N_16081,N_17904);
or U19884 (N_19884,N_16048,N_17445);
nor U19885 (N_19885,N_16993,N_16384);
or U19886 (N_19886,N_16920,N_17347);
nor U19887 (N_19887,N_16981,N_16617);
nand U19888 (N_19888,N_16654,N_17483);
and U19889 (N_19889,N_17286,N_17019);
nand U19890 (N_19890,N_16603,N_16569);
nor U19891 (N_19891,N_17065,N_17649);
xnor U19892 (N_19892,N_17687,N_16274);
and U19893 (N_19893,N_16839,N_17551);
and U19894 (N_19894,N_17323,N_17217);
or U19895 (N_19895,N_16196,N_17292);
nor U19896 (N_19896,N_16255,N_16612);
nand U19897 (N_19897,N_17241,N_16644);
xnor U19898 (N_19898,N_16415,N_16887);
or U19899 (N_19899,N_17689,N_17964);
nor U19900 (N_19900,N_16955,N_16080);
nor U19901 (N_19901,N_16554,N_16782);
or U19902 (N_19902,N_16577,N_17894);
or U19903 (N_19903,N_17242,N_16237);
and U19904 (N_19904,N_17273,N_17138);
xor U19905 (N_19905,N_16095,N_16255);
nand U19906 (N_19906,N_16118,N_16747);
or U19907 (N_19907,N_16906,N_16626);
and U19908 (N_19908,N_16116,N_17233);
or U19909 (N_19909,N_17212,N_17867);
or U19910 (N_19910,N_16753,N_17177);
nand U19911 (N_19911,N_17996,N_17981);
and U19912 (N_19912,N_17675,N_16640);
nand U19913 (N_19913,N_16864,N_17353);
nand U19914 (N_19914,N_16912,N_16102);
nand U19915 (N_19915,N_16581,N_16023);
xnor U19916 (N_19916,N_16899,N_17550);
xor U19917 (N_19917,N_17395,N_17056);
xnor U19918 (N_19918,N_17079,N_17327);
nand U19919 (N_19919,N_17313,N_16981);
nand U19920 (N_19920,N_17106,N_17683);
nor U19921 (N_19921,N_16659,N_17971);
nand U19922 (N_19922,N_16642,N_16043);
or U19923 (N_19923,N_16297,N_17636);
or U19924 (N_19924,N_16376,N_17876);
and U19925 (N_19925,N_16705,N_16488);
or U19926 (N_19926,N_16163,N_17326);
and U19927 (N_19927,N_16579,N_16226);
nor U19928 (N_19928,N_17169,N_17197);
or U19929 (N_19929,N_16898,N_16096);
or U19930 (N_19930,N_17166,N_17714);
xnor U19931 (N_19931,N_16695,N_16254);
xnor U19932 (N_19932,N_17768,N_17799);
and U19933 (N_19933,N_17901,N_16677);
or U19934 (N_19934,N_16817,N_16077);
or U19935 (N_19935,N_17127,N_17034);
xor U19936 (N_19936,N_17054,N_16136);
and U19937 (N_19937,N_17472,N_17655);
nand U19938 (N_19938,N_16690,N_16688);
nor U19939 (N_19939,N_16225,N_16502);
or U19940 (N_19940,N_17588,N_16288);
and U19941 (N_19941,N_16572,N_17271);
xnor U19942 (N_19942,N_16393,N_16382);
and U19943 (N_19943,N_16390,N_17553);
nor U19944 (N_19944,N_16064,N_17456);
xor U19945 (N_19945,N_16009,N_17719);
and U19946 (N_19946,N_17511,N_17672);
and U19947 (N_19947,N_17705,N_17536);
xor U19948 (N_19948,N_16537,N_17332);
nand U19949 (N_19949,N_17566,N_17555);
or U19950 (N_19950,N_17286,N_16371);
and U19951 (N_19951,N_16117,N_17830);
and U19952 (N_19952,N_16316,N_16121);
nand U19953 (N_19953,N_17634,N_16916);
or U19954 (N_19954,N_16112,N_16682);
and U19955 (N_19955,N_17732,N_17818);
or U19956 (N_19956,N_16906,N_16913);
xor U19957 (N_19957,N_16357,N_17664);
nand U19958 (N_19958,N_17096,N_17087);
and U19959 (N_19959,N_17247,N_17100);
nand U19960 (N_19960,N_16511,N_17991);
nand U19961 (N_19961,N_17014,N_16955);
and U19962 (N_19962,N_16688,N_17466);
or U19963 (N_19963,N_17731,N_16535);
or U19964 (N_19964,N_17417,N_17186);
or U19965 (N_19965,N_16154,N_17048);
nand U19966 (N_19966,N_17312,N_16625);
and U19967 (N_19967,N_16048,N_16040);
nand U19968 (N_19968,N_17289,N_17942);
nand U19969 (N_19969,N_16254,N_17001);
and U19970 (N_19970,N_16648,N_17128);
nand U19971 (N_19971,N_16734,N_16193);
nand U19972 (N_19972,N_17131,N_17827);
xnor U19973 (N_19973,N_16764,N_17065);
or U19974 (N_19974,N_17405,N_16000);
xor U19975 (N_19975,N_17863,N_16160);
or U19976 (N_19976,N_17499,N_16978);
and U19977 (N_19977,N_16786,N_17192);
or U19978 (N_19978,N_16026,N_17090);
and U19979 (N_19979,N_16947,N_17440);
nand U19980 (N_19980,N_17613,N_17644);
or U19981 (N_19981,N_16019,N_16141);
xor U19982 (N_19982,N_16249,N_16233);
xor U19983 (N_19983,N_17874,N_16316);
or U19984 (N_19984,N_16335,N_17673);
and U19985 (N_19985,N_17630,N_17407);
and U19986 (N_19986,N_17091,N_16592);
nor U19987 (N_19987,N_17910,N_16986);
nor U19988 (N_19988,N_16378,N_16078);
or U19989 (N_19989,N_16015,N_16311);
and U19990 (N_19990,N_17328,N_16305);
xnor U19991 (N_19991,N_16072,N_16435);
and U19992 (N_19992,N_17368,N_17574);
nor U19993 (N_19993,N_16192,N_16269);
xnor U19994 (N_19994,N_16624,N_17027);
or U19995 (N_19995,N_17041,N_16544);
nor U19996 (N_19996,N_16307,N_17077);
or U19997 (N_19997,N_16151,N_17424);
xnor U19998 (N_19998,N_16614,N_17994);
and U19999 (N_19999,N_16472,N_17919);
and U20000 (N_20000,N_18403,N_19821);
and U20001 (N_20001,N_18228,N_18157);
or U20002 (N_20002,N_19776,N_18912);
and U20003 (N_20003,N_19659,N_18033);
nand U20004 (N_20004,N_19143,N_18560);
xnor U20005 (N_20005,N_19059,N_18981);
nor U20006 (N_20006,N_19699,N_18372);
or U20007 (N_20007,N_19483,N_18668);
nand U20008 (N_20008,N_19184,N_19089);
or U20009 (N_20009,N_19269,N_18716);
and U20010 (N_20010,N_18522,N_18278);
or U20011 (N_20011,N_19218,N_18335);
nor U20012 (N_20012,N_19547,N_18294);
nand U20013 (N_20013,N_19477,N_18987);
or U20014 (N_20014,N_18221,N_19883);
or U20015 (N_20015,N_19681,N_18212);
nand U20016 (N_20016,N_18949,N_19401);
or U20017 (N_20017,N_18737,N_18176);
nor U20018 (N_20018,N_18217,N_19408);
nand U20019 (N_20019,N_19562,N_19406);
nand U20020 (N_20020,N_19279,N_18154);
nand U20021 (N_20021,N_19370,N_19651);
and U20022 (N_20022,N_18750,N_19083);
xor U20023 (N_20023,N_18236,N_18696);
nand U20024 (N_20024,N_18068,N_18362);
nor U20025 (N_20025,N_19325,N_19809);
nand U20026 (N_20026,N_19904,N_18563);
nand U20027 (N_20027,N_18506,N_19466);
xnor U20028 (N_20028,N_19860,N_18349);
nor U20029 (N_20029,N_18074,N_19046);
and U20030 (N_20030,N_19637,N_18614);
nand U20031 (N_20031,N_18100,N_19430);
and U20032 (N_20032,N_19747,N_19315);
xor U20033 (N_20033,N_18173,N_19373);
and U20034 (N_20034,N_18960,N_19800);
nor U20035 (N_20035,N_19073,N_18183);
nor U20036 (N_20036,N_18689,N_18321);
or U20037 (N_20037,N_18865,N_19364);
nand U20038 (N_20038,N_19443,N_18768);
nor U20039 (N_20039,N_18876,N_18771);
xnor U20040 (N_20040,N_19144,N_19485);
nor U20041 (N_20041,N_19645,N_18914);
and U20042 (N_20042,N_18685,N_19070);
or U20043 (N_20043,N_19424,N_19103);
xor U20044 (N_20044,N_19623,N_18859);
or U20045 (N_20045,N_18772,N_19224);
nand U20046 (N_20046,N_19322,N_18093);
or U20047 (N_20047,N_19422,N_18007);
and U20048 (N_20048,N_18323,N_19022);
xor U20049 (N_20049,N_18240,N_19689);
xnor U20050 (N_20050,N_18924,N_19423);
xnor U20051 (N_20051,N_18761,N_19425);
or U20052 (N_20052,N_18995,N_18430);
and U20053 (N_20053,N_19036,N_18940);
xor U20054 (N_20054,N_18029,N_19270);
or U20055 (N_20055,N_19072,N_19014);
or U20056 (N_20056,N_19565,N_18137);
nand U20057 (N_20057,N_19569,N_19152);
xnor U20058 (N_20058,N_19729,N_18518);
xor U20059 (N_20059,N_18302,N_19034);
and U20060 (N_20060,N_18637,N_19688);
or U20061 (N_20061,N_19399,N_18624);
or U20062 (N_20062,N_19716,N_19625);
and U20063 (N_20063,N_19824,N_19174);
nor U20064 (N_20064,N_19635,N_19508);
or U20065 (N_20065,N_18097,N_18079);
xnor U20066 (N_20066,N_18818,N_18308);
xnor U20067 (N_20067,N_18794,N_18680);
or U20068 (N_20068,N_18164,N_19177);
nor U20069 (N_20069,N_18819,N_19518);
and U20070 (N_20070,N_18799,N_18941);
nor U20071 (N_20071,N_19323,N_19032);
xnor U20072 (N_20072,N_19332,N_18424);
xnor U20073 (N_20073,N_18992,N_18836);
and U20074 (N_20074,N_18516,N_19135);
nor U20075 (N_20075,N_19116,N_18063);
or U20076 (N_20076,N_18036,N_19522);
nor U20077 (N_20077,N_18891,N_19390);
xnor U20078 (N_20078,N_18918,N_18070);
and U20079 (N_20079,N_18852,N_19428);
and U20080 (N_20080,N_19722,N_19843);
and U20081 (N_20081,N_19634,N_18042);
and U20082 (N_20082,N_18666,N_19272);
or U20083 (N_20083,N_19544,N_19138);
nor U20084 (N_20084,N_19222,N_19000);
nor U20085 (N_20085,N_18131,N_19762);
or U20086 (N_20086,N_19245,N_18965);
nand U20087 (N_20087,N_18444,N_19249);
xor U20088 (N_20088,N_18883,N_18727);
or U20089 (N_20089,N_19969,N_18448);
or U20090 (N_20090,N_18001,N_18863);
and U20091 (N_20091,N_19229,N_19437);
nand U20092 (N_20092,N_18931,N_19538);
and U20093 (N_20093,N_19705,N_18290);
or U20094 (N_20094,N_18222,N_19853);
nand U20095 (N_20095,N_19171,N_18710);
nand U20096 (N_20096,N_19781,N_19801);
xnor U20097 (N_20097,N_18408,N_18796);
and U20098 (N_20098,N_19080,N_18648);
nor U20099 (N_20099,N_19713,N_19134);
nor U20100 (N_20100,N_19907,N_19025);
nor U20101 (N_20101,N_19449,N_19403);
nor U20102 (N_20102,N_19182,N_18967);
nor U20103 (N_20103,N_19890,N_19361);
nor U20104 (N_20104,N_19710,N_18583);
nand U20105 (N_20105,N_18571,N_19368);
or U20106 (N_20106,N_18250,N_18446);
or U20107 (N_20107,N_19301,N_19504);
or U20108 (N_20108,N_18485,N_19395);
and U20109 (N_20109,N_18982,N_19393);
or U20110 (N_20110,N_18005,N_18520);
nor U20111 (N_20111,N_19082,N_18358);
and U20112 (N_20112,N_19844,N_18229);
xnor U20113 (N_20113,N_18718,N_19923);
or U20114 (N_20114,N_18249,N_18721);
or U20115 (N_20115,N_18986,N_19299);
and U20116 (N_20116,N_18880,N_19755);
and U20117 (N_20117,N_18199,N_19136);
and U20118 (N_20118,N_19398,N_19760);
or U20119 (N_20119,N_18990,N_19058);
xnor U20120 (N_20120,N_18385,N_18821);
nor U20121 (N_20121,N_18925,N_18251);
xnor U20122 (N_20122,N_19978,N_18704);
xor U20123 (N_20123,N_18023,N_19763);
nor U20124 (N_20124,N_18656,N_19313);
and U20125 (N_20125,N_19510,N_19856);
or U20126 (N_20126,N_18676,N_18850);
nor U20127 (N_20127,N_19546,N_18628);
and U20128 (N_20128,N_19861,N_19181);
nor U20129 (N_20129,N_19663,N_19740);
nand U20130 (N_20130,N_18782,N_19436);
or U20131 (N_20131,N_19010,N_18609);
xnor U20132 (N_20132,N_18592,N_19811);
nand U20133 (N_20133,N_18846,N_19990);
nor U20134 (N_20134,N_18622,N_19905);
and U20135 (N_20135,N_18184,N_19750);
nand U20136 (N_20136,N_18418,N_18928);
and U20137 (N_20137,N_19605,N_19071);
xor U20138 (N_20138,N_18998,N_19570);
or U20139 (N_20139,N_18599,N_19029);
nand U20140 (N_20140,N_18428,N_19870);
or U20141 (N_20141,N_19916,N_18177);
xnor U20142 (N_20142,N_18921,N_18031);
and U20143 (N_20143,N_19372,N_19385);
xnor U20144 (N_20144,N_19284,N_18617);
and U20145 (N_20145,N_19668,N_19382);
xnor U20146 (N_20146,N_18829,N_18345);
and U20147 (N_20147,N_18875,N_19557);
xnor U20148 (N_20148,N_19780,N_18463);
xnor U20149 (N_20149,N_18565,N_19197);
and U20150 (N_20150,N_19551,N_19097);
or U20151 (N_20151,N_19859,N_18310);
xnor U20152 (N_20152,N_18155,N_18165);
xor U20153 (N_20153,N_19037,N_18387);
and U20154 (N_20154,N_18320,N_19392);
and U20155 (N_20155,N_18101,N_18125);
xor U20156 (N_20156,N_19283,N_19078);
and U20157 (N_20157,N_18793,N_19992);
nand U20158 (N_20158,N_18313,N_19964);
or U20159 (N_20159,N_18469,N_19489);
xnor U20160 (N_20160,N_19888,N_18889);
and U20161 (N_20161,N_19559,N_19951);
and U20162 (N_20162,N_19342,N_19060);
xor U20163 (N_20163,N_19974,N_19153);
or U20164 (N_20164,N_19933,N_19062);
nor U20165 (N_20165,N_18851,N_18582);
and U20166 (N_20166,N_19556,N_19784);
nand U20167 (N_20167,N_19604,N_18479);
xor U20168 (N_20168,N_18646,N_19040);
nand U20169 (N_20169,N_19259,N_19051);
xor U20170 (N_20170,N_19291,N_18726);
xnor U20171 (N_20171,N_19346,N_18091);
nor U20172 (N_20172,N_18466,N_18871);
and U20173 (N_20173,N_18415,N_18351);
or U20174 (N_20174,N_19640,N_19327);
and U20175 (N_20175,N_18114,N_18507);
or U20176 (N_20176,N_19852,N_18433);
nor U20177 (N_20177,N_18650,N_18086);
nor U20178 (N_20178,N_19910,N_18795);
or U20179 (N_20179,N_18574,N_18511);
nor U20180 (N_20180,N_19986,N_19665);
nand U20181 (N_20181,N_18293,N_18645);
or U20182 (N_20182,N_18807,N_18247);
or U20183 (N_20183,N_18939,N_19490);
and U20184 (N_20184,N_19267,N_19217);
xnor U20185 (N_20185,N_18398,N_18275);
nand U20186 (N_20186,N_18567,N_19312);
xnor U20187 (N_20187,N_19446,N_19410);
nand U20188 (N_20188,N_19384,N_19375);
nor U20189 (N_20189,N_19758,N_18907);
nor U20190 (N_20190,N_19199,N_18585);
or U20191 (N_20191,N_19955,N_19934);
or U20192 (N_20192,N_19244,N_18206);
and U20193 (N_20193,N_19525,N_19421);
nand U20194 (N_20194,N_18025,N_19351);
and U20195 (N_20195,N_18179,N_18800);
and U20196 (N_20196,N_18739,N_18575);
or U20197 (N_20197,N_19028,N_18550);
nor U20198 (N_20198,N_18041,N_19488);
nor U20199 (N_20199,N_19769,N_18473);
xnor U20200 (N_20200,N_19118,N_19087);
nor U20201 (N_20201,N_18942,N_18845);
and U20202 (N_20202,N_18627,N_18066);
and U20203 (N_20203,N_19167,N_18734);
nor U20204 (N_20204,N_18088,N_18935);
nand U20205 (N_20205,N_18665,N_19629);
and U20206 (N_20206,N_19338,N_19761);
nand U20207 (N_20207,N_19328,N_18442);
or U20208 (N_20208,N_19924,N_18970);
nand U20209 (N_20209,N_18766,N_18438);
nand U20210 (N_20210,N_18738,N_19670);
nand U20211 (N_20211,N_19193,N_19413);
and U20212 (N_20212,N_18352,N_19994);
or U20213 (N_20213,N_19287,N_19516);
nor U20214 (N_20214,N_18467,N_18080);
or U20215 (N_20215,N_18555,N_19814);
or U20216 (N_20216,N_19976,N_18306);
nor U20217 (N_20217,N_19273,N_18156);
nor U20218 (N_20218,N_19369,N_19254);
nand U20219 (N_20219,N_18162,N_18402);
nand U20220 (N_20220,N_19336,N_18653);
nor U20221 (N_20221,N_18966,N_18143);
and U20222 (N_20222,N_18754,N_18030);
and U20223 (N_20223,N_19013,N_19977);
or U20224 (N_20224,N_18194,N_19360);
xor U20225 (N_20225,N_19643,N_18363);
xnor U20226 (N_20226,N_18246,N_18964);
and U20227 (N_20227,N_18498,N_18253);
or U20228 (N_20228,N_18142,N_19748);
xor U20229 (N_20229,N_18644,N_19444);
nand U20230 (N_20230,N_19157,N_19628);
and U20231 (N_20231,N_18693,N_19210);
nand U20232 (N_20232,N_19685,N_19148);
nand U20233 (N_20233,N_19632,N_18762);
or U20234 (N_20234,N_18632,N_19906);
nand U20235 (N_20235,N_18626,N_18468);
or U20236 (N_20236,N_19447,N_18943);
nor U20237 (N_20237,N_19137,N_18910);
or U20238 (N_20238,N_19965,N_18531);
nor U20239 (N_20239,N_18878,N_18200);
or U20240 (N_20240,N_19952,N_19595);
xor U20241 (N_20241,N_18434,N_19469);
or U20242 (N_20242,N_18346,N_18312);
xor U20243 (N_20243,N_18135,N_19110);
nand U20244 (N_20244,N_18396,N_18404);
and U20245 (N_20245,N_18751,N_19894);
xor U20246 (N_20246,N_19439,N_18535);
xor U20247 (N_20247,N_18687,N_18725);
xnor U20248 (N_20248,N_18407,N_19517);
xnor U20249 (N_20249,N_19956,N_18440);
nor U20250 (N_20250,N_18778,N_19828);
nor U20251 (N_20251,N_18746,N_18413);
or U20252 (N_20252,N_19711,N_19818);
nand U20253 (N_20253,N_19168,N_18860);
nand U20254 (N_20254,N_18115,N_19592);
xnor U20255 (N_20255,N_18549,N_19129);
and U20256 (N_20256,N_19063,N_19460);
and U20257 (N_20257,N_18929,N_18003);
xor U20258 (N_20258,N_19467,N_19105);
and U20259 (N_20259,N_18411,N_19065);
xor U20260 (N_20260,N_19094,N_18075);
and U20261 (N_20261,N_18060,N_19731);
or U20262 (N_20262,N_19260,N_19702);
xor U20263 (N_20263,N_18309,N_19473);
xnor U20264 (N_20264,N_19768,N_19957);
nor U20265 (N_20265,N_18455,N_18061);
and U20266 (N_20266,N_19201,N_18338);
and U20267 (N_20267,N_19339,N_19194);
and U20268 (N_20268,N_19414,N_19854);
or U20269 (N_20269,N_18368,N_19441);
xnor U20270 (N_20270,N_18618,N_18077);
xnor U20271 (N_20271,N_18374,N_18108);
and U20272 (N_20272,N_18777,N_18561);
nor U20273 (N_20273,N_19119,N_18615);
nor U20274 (N_20274,N_19012,N_19827);
and U20275 (N_20275,N_19999,N_19819);
xnor U20276 (N_20276,N_18745,N_18420);
nor U20277 (N_20277,N_19367,N_19603);
and U20278 (N_20278,N_18926,N_18528);
and U20279 (N_20279,N_19618,N_18279);
nand U20280 (N_20280,N_18529,N_18515);
xnor U20281 (N_20281,N_19812,N_18607);
or U20282 (N_20282,N_19732,N_18414);
nand U20283 (N_20283,N_19198,N_18056);
xor U20284 (N_20284,N_19541,N_19838);
or U20285 (N_20285,N_19627,N_19093);
xor U20286 (N_20286,N_18841,N_18775);
nand U20287 (N_20287,N_18215,N_18705);
xnor U20288 (N_20288,N_19112,N_19695);
nand U20289 (N_20289,N_18767,N_18877);
xor U20290 (N_20290,N_18011,N_19100);
nand U20291 (N_20291,N_19672,N_19589);
or U20292 (N_20292,N_18994,N_18603);
or U20293 (N_20293,N_19727,N_18616);
or U20294 (N_20294,N_19462,N_19175);
xor U20295 (N_20295,N_18825,N_18936);
xnor U20296 (N_20296,N_18867,N_19052);
and U20297 (N_20297,N_18714,N_18741);
nor U20298 (N_20298,N_19962,N_18629);
nand U20299 (N_20299,N_19615,N_18219);
nor U20300 (N_20300,N_19825,N_19054);
xnor U20301 (N_20301,N_19246,N_19793);
xnor U20302 (N_20302,N_18698,N_18728);
nor U20303 (N_20303,N_18623,N_18755);
xor U20304 (N_20304,N_19350,N_18381);
or U20305 (N_20305,N_18923,N_18817);
and U20306 (N_20306,N_19880,N_19026);
and U20307 (N_20307,N_18132,N_18786);
xor U20308 (N_20308,N_19730,N_19009);
and U20309 (N_20309,N_19739,N_18748);
xor U20310 (N_20310,N_18113,N_18858);
xor U20311 (N_20311,N_18127,N_18933);
and U20312 (N_20312,N_19912,N_19720);
or U20313 (N_20313,N_19987,N_18499);
or U20314 (N_20314,N_18158,N_19832);
xor U20315 (N_20315,N_18214,N_18071);
nor U20316 (N_20316,N_18930,N_19409);
and U20317 (N_20317,N_18613,N_18546);
xnor U20318 (N_20318,N_18882,N_19988);
nand U20319 (N_20319,N_19836,N_19981);
xnor U20320 (N_20320,N_19804,N_19024);
xor U20321 (N_20321,N_19400,N_18961);
and U20322 (N_20322,N_19268,N_19434);
xor U20323 (N_20323,N_18684,N_18733);
xnor U20324 (N_20324,N_18392,N_19122);
xnor U20325 (N_20325,N_19719,N_18758);
or U20326 (N_20326,N_19234,N_18118);
and U20327 (N_20327,N_18286,N_18631);
xnor U20328 (N_20328,N_18067,N_19867);
or U20329 (N_20329,N_19172,N_18090);
nor U20330 (N_20330,N_19653,N_19305);
nor U20331 (N_20331,N_18979,N_19366);
or U20332 (N_20332,N_18443,N_18129);
nor U20333 (N_20333,N_19225,N_19757);
and U20334 (N_20334,N_18119,N_18210);
or U20335 (N_20335,N_18674,N_18806);
nand U20336 (N_20336,N_18897,N_19468);
nand U20337 (N_20337,N_19124,N_19155);
nor U20338 (N_20338,N_18740,N_19391);
or U20339 (N_20339,N_18364,N_19285);
nor U20340 (N_20340,N_18519,N_18743);
xor U20341 (N_20341,N_19333,N_18901);
or U20342 (N_20342,N_19524,N_18054);
xor U20343 (N_20343,N_19652,N_18465);
nand U20344 (N_20344,N_18419,N_18834);
xnor U20345 (N_20345,N_19113,N_19030);
or U20346 (N_20346,N_19514,N_19458);
xor U20347 (N_20347,N_19253,N_18259);
and U20348 (N_20348,N_19146,N_19806);
or U20349 (N_20349,N_19214,N_18647);
and U20350 (N_20350,N_18804,N_18837);
xnor U20351 (N_20351,N_18216,N_19318);
or U20352 (N_20352,N_19127,N_19908);
nor U20353 (N_20353,N_18780,N_19042);
nand U20354 (N_20354,N_18749,N_18999);
and U20355 (N_20355,N_19344,N_19297);
nor U20356 (N_20356,N_18815,N_19501);
nor U20357 (N_20357,N_19728,N_18873);
and U20358 (N_20358,N_19335,N_19789);
or U20359 (N_20359,N_19884,N_18577);
nand U20360 (N_20360,N_18756,N_19102);
nand U20361 (N_20361,N_19221,N_19035);
xnor U20362 (N_20362,N_19376,N_19178);
or U20363 (N_20363,N_19076,N_19831);
or U20364 (N_20364,N_18094,N_18327);
nand U20365 (N_20365,N_18630,N_18572);
xnor U20366 (N_20366,N_19919,N_18483);
and U20367 (N_20367,N_19091,N_19461);
and U20368 (N_20368,N_18654,N_18120);
nor U20369 (N_20369,N_19170,N_19998);
and U20370 (N_20370,N_18678,N_18608);
nor U20371 (N_20371,N_18445,N_19950);
xnor U20372 (N_20372,N_18611,N_18089);
or U20373 (N_20373,N_18224,N_19989);
nand U20374 (N_20374,N_19031,N_19185);
and U20375 (N_20375,N_19250,N_18134);
nor U20376 (N_20376,N_19017,N_18272);
nand U20377 (N_20377,N_19191,N_18649);
nor U20378 (N_20378,N_19359,N_18002);
nor U20379 (N_20379,N_18126,N_19238);
nor U20380 (N_20380,N_18972,N_19872);
or U20381 (N_20381,N_19106,N_18497);
nor U20382 (N_20382,N_18573,N_19474);
xnor U20383 (N_20383,N_19785,N_18081);
xor U20384 (N_20384,N_19188,N_19644);
or U20385 (N_20385,N_18014,N_18591);
and U20386 (N_20386,N_18879,N_19145);
nor U20387 (N_20387,N_18422,N_19111);
nand U20388 (N_20388,N_18706,N_19797);
nand U20389 (N_20389,N_19650,N_19515);
nand U20390 (N_20390,N_18038,N_18416);
and U20391 (N_20391,N_18285,N_19209);
xor U20392 (N_20392,N_18301,N_18894);
and U20393 (N_20393,N_19521,N_18536);
xnor U20394 (N_20394,N_19180,N_19189);
and U20395 (N_20395,N_18092,N_19638);
nor U20396 (N_20396,N_18270,N_19823);
nor U20397 (N_20397,N_18412,N_19495);
nand U20398 (N_20398,N_19979,N_19614);
or U20399 (N_20399,N_18854,N_19163);
xor U20400 (N_20400,N_19343,N_18139);
or U20401 (N_20401,N_18744,N_19107);
and U20402 (N_20402,N_19772,N_19737);
or U20403 (N_20403,N_18830,N_18307);
and U20404 (N_20404,N_19481,N_18956);
and U20405 (N_20405,N_18017,N_18384);
xnor U20406 (N_20406,N_19531,N_19995);
nand U20407 (N_20407,N_18087,N_19271);
nand U20408 (N_20408,N_19736,N_18811);
xor U20409 (N_20409,N_19708,N_18357);
or U20410 (N_20410,N_19085,N_18579);
nor U20411 (N_20411,N_18322,N_19928);
or U20412 (N_20412,N_18759,N_18542);
and U20413 (N_20413,N_19889,N_19543);
and U20414 (N_20414,N_18109,N_18848);
and U20415 (N_20415,N_19104,N_19656);
or U20416 (N_20416,N_18258,N_18742);
or U20417 (N_20417,N_19735,N_18723);
xor U20418 (N_20418,N_18525,N_18110);
or U20419 (N_20419,N_19915,N_19165);
nand U20420 (N_20420,N_18035,N_19050);
nor U20421 (N_20421,N_19620,N_19892);
nand U20422 (N_20422,N_19683,N_19230);
nand U20423 (N_20423,N_18791,N_18513);
xnor U20424 (N_20424,N_19457,N_18547);
nor U20425 (N_20425,N_18973,N_19971);
nor U20426 (N_20426,N_18694,N_19298);
or U20427 (N_20427,N_19223,N_18356);
and U20428 (N_20428,N_19537,N_19139);
nand U20429 (N_20429,N_19341,N_19834);
nor U20430 (N_20430,N_18261,N_18810);
nand U20431 (N_20431,N_18371,N_18269);
or U20432 (N_20432,N_19863,N_19275);
nor U20433 (N_20433,N_19169,N_18974);
xor U20434 (N_20434,N_18190,N_19897);
and U20435 (N_20435,N_19611,N_19573);
or U20436 (N_20436,N_19725,N_18043);
nor U20437 (N_20437,N_18789,N_18152);
or U20438 (N_20438,N_19162,N_19622);
xnor U20439 (N_20439,N_19926,N_18764);
and U20440 (N_20440,N_18069,N_18773);
and U20441 (N_20441,N_18566,N_18559);
and U20442 (N_20442,N_18785,N_19004);
xnor U20443 (N_20443,N_18470,N_19802);
xnor U20444 (N_20444,N_19120,N_19787);
nor U20445 (N_20445,N_19452,N_18451);
and U20446 (N_20446,N_19079,N_19936);
and U20447 (N_20447,N_19451,N_18605);
xor U20448 (N_20448,N_19677,N_19433);
or U20449 (N_20449,N_18803,N_19426);
nand U20450 (N_20450,N_18695,N_19349);
nor U20451 (N_20451,N_18452,N_19745);
nor U20452 (N_20452,N_18776,N_19011);
or U20453 (N_20453,N_18441,N_19554);
xnor U20454 (N_20454,N_18328,N_18911);
nand U20455 (N_20455,N_19237,N_19846);
nand U20456 (N_20456,N_18193,N_18736);
and U20457 (N_20457,N_18098,N_18373);
xnor U20458 (N_20458,N_18458,N_19128);
nor U20459 (N_20459,N_18257,N_18857);
and U20460 (N_20460,N_19532,N_19602);
or U20461 (N_20461,N_18082,N_18957);
and U20462 (N_20462,N_18288,N_18341);
nor U20463 (N_20463,N_19081,N_18149);
or U20464 (N_20464,N_19816,N_19764);
xor U20465 (N_20465,N_19302,N_19893);
xnor U20466 (N_20466,N_19156,N_18204);
and U20467 (N_20467,N_18150,N_19450);
and U20468 (N_20468,N_18205,N_18289);
and U20469 (N_20469,N_19953,N_18378);
or U20470 (N_20470,N_19161,N_18581);
and U20471 (N_20471,N_18317,N_18227);
xor U20472 (N_20472,N_18480,N_18798);
or U20473 (N_20473,N_18874,N_18501);
or U20474 (N_20474,N_18065,N_19631);
nor U20475 (N_20475,N_18096,N_18051);
or U20476 (N_20476,N_18523,N_19712);
nor U20477 (N_20477,N_18192,N_18032);
nand U20478 (N_20478,N_18638,N_19154);
nand U20479 (N_20479,N_19311,N_19598);
nand U20480 (N_20480,N_19130,N_18147);
nand U20481 (N_20481,N_19389,N_19558);
nand U20482 (N_20482,N_18008,N_19326);
nor U20483 (N_20483,N_19205,N_18866);
and U20484 (N_20484,N_18625,N_19179);
nand U20485 (N_20485,N_19920,N_19057);
and U20486 (N_20486,N_19258,N_19362);
or U20487 (N_20487,N_18870,N_18655);
nand U20488 (N_20488,N_18887,N_19519);
xor U20489 (N_20489,N_19574,N_18765);
and U20490 (N_20490,N_18606,N_18849);
nand U20491 (N_20491,N_18658,N_19803);
xnor U20492 (N_20492,N_18230,N_19619);
or U20493 (N_20493,N_19718,N_19572);
and U20494 (N_20494,N_18046,N_18006);
or U20495 (N_20495,N_19061,N_18636);
nor U20496 (N_20496,N_18460,N_18673);
nand U20497 (N_20497,N_19123,N_19997);
xor U20498 (N_20498,N_18937,N_18012);
xor U20499 (N_20499,N_19542,N_18602);
xor U20500 (N_20500,N_19575,N_18146);
xnor U20501 (N_20501,N_19251,N_18209);
or U20502 (N_20502,N_19503,N_19109);
nor U20503 (N_20503,N_19734,N_18720);
nor U20504 (N_20504,N_18273,N_19835);
or U20505 (N_20505,N_18620,N_18872);
or U20506 (N_20506,N_19512,N_18487);
and U20507 (N_20507,N_19243,N_18331);
xnor U20508 (N_20508,N_18196,N_18541);
or U20509 (N_20509,N_19241,N_19585);
xnor U20510 (N_20510,N_18037,N_19917);
and U20511 (N_20511,N_19227,N_18753);
nand U20512 (N_20512,N_19680,N_18332);
nor U20513 (N_20513,N_18099,N_19767);
and U20514 (N_20514,N_18840,N_18556);
or U20515 (N_20515,N_18153,N_18292);
or U20516 (N_20516,N_18593,N_18144);
and U20517 (N_20517,N_18844,N_18314);
nand U20518 (N_20518,N_19868,N_18504);
nor U20519 (N_20519,N_19263,N_18138);
nor U20520 (N_20520,N_19088,N_18256);
nor U20521 (N_20521,N_18781,N_19190);
nand U20522 (N_20522,N_18174,N_18564);
xor U20523 (N_20523,N_18985,N_18393);
or U20524 (N_20524,N_19334,N_18300);
nand U20525 (N_20525,N_18554,N_19496);
or U20526 (N_20526,N_19647,N_19788);
nor U20527 (N_20527,N_18505,N_18447);
nand U20528 (N_20528,N_18968,N_18178);
xnor U20529 (N_20529,N_18816,N_19690);
and U20530 (N_20530,N_19983,N_18832);
and U20531 (N_20531,N_19958,N_19470);
xor U20532 (N_20532,N_19829,N_19943);
and U20533 (N_20533,N_19371,N_18000);
or U20534 (N_20534,N_19239,N_19493);
xnor U20535 (N_20535,N_19675,N_18130);
or U20536 (N_20536,N_19945,N_19453);
xnor U20537 (N_20537,N_19706,N_18195);
nor U20538 (N_20538,N_18427,N_19386);
and U20539 (N_20539,N_19862,N_19813);
and U20540 (N_20540,N_18978,N_18048);
nand U20541 (N_20541,N_18348,N_18218);
xor U20542 (N_20542,N_19662,N_18596);
or U20543 (N_20543,N_19590,N_18808);
and U20544 (N_20544,N_18477,N_19412);
and U20545 (N_20545,N_18024,N_18397);
or U20546 (N_20546,N_19023,N_19633);
and U20547 (N_20547,N_19869,N_19095);
nand U20548 (N_20548,N_18034,N_18388);
nor U20549 (N_20549,N_19513,N_18682);
xnor U20550 (N_20550,N_19126,N_19837);
xor U20551 (N_20551,N_19090,N_18220);
nor U20552 (N_20552,N_19497,N_18018);
or U20553 (N_20553,N_19377,N_19968);
xor U20554 (N_20554,N_19545,N_18813);
xnor U20555 (N_20555,N_18589,N_18234);
nor U20556 (N_20556,N_19117,N_19655);
or U20557 (N_20557,N_19183,N_18161);
and U20558 (N_20558,N_18769,N_19125);
or U20559 (N_20559,N_18337,N_19387);
xnor U20560 (N_20560,N_19577,N_19511);
and U20561 (N_20561,N_19815,N_18026);
or U20562 (N_20562,N_19141,N_19555);
nor U20563 (N_20563,N_19612,N_18494);
xnor U20564 (N_20564,N_18400,N_19865);
and U20565 (N_20565,N_18692,N_19654);
and U20566 (N_20566,N_18989,N_19966);
and U20567 (N_20567,N_19388,N_18537);
xnor U20568 (N_20568,N_18920,N_18580);
xnor U20569 (N_20569,N_18717,N_19252);
or U20570 (N_20570,N_18040,N_18826);
xor U20571 (N_20571,N_19563,N_18963);
nand U20572 (N_20572,N_19552,N_18802);
nand U20573 (N_20573,N_18324,N_18333);
nand U20574 (N_20574,N_19247,N_19895);
nor U20575 (N_20575,N_19586,N_19084);
xor U20576 (N_20576,N_19658,N_18595);
xor U20577 (N_20577,N_19526,N_19584);
and U20578 (N_20578,N_19753,N_18410);
nor U20579 (N_20579,N_19848,N_18252);
and U20580 (N_20580,N_18670,N_19459);
and U20581 (N_20581,N_18634,N_18488);
nor U20582 (N_20582,N_18284,N_18896);
or U20583 (N_20583,N_18828,N_18553);
or U20584 (N_20584,N_19363,N_18232);
nor U20585 (N_20585,N_18481,N_19355);
and U20586 (N_20586,N_18326,N_18083);
xor U20587 (N_20587,N_19972,N_19864);
or U20588 (N_20588,N_19231,N_18588);
or U20589 (N_20589,N_19448,N_18122);
xnor U20590 (N_20590,N_18980,N_19944);
xnor U20591 (N_20591,N_18235,N_19845);
or U20592 (N_20592,N_19160,N_19576);
or U20593 (N_20593,N_18962,N_18991);
nand U20594 (N_20594,N_18783,N_19808);
xnor U20595 (N_20595,N_18475,N_18248);
xnor U20596 (N_20596,N_18202,N_18484);
and U20597 (N_20597,N_18171,N_18927);
nand U20598 (N_20598,N_19970,N_18702);
xor U20599 (N_20599,N_19075,N_18291);
nor U20600 (N_20600,N_18339,N_18457);
xnor U20601 (N_20601,N_18534,N_19098);
and U20602 (N_20602,N_18639,N_18262);
or U20603 (N_20603,N_19693,N_18955);
xnor U20604 (N_20604,N_19927,N_18208);
nor U20605 (N_20605,N_19020,N_18735);
nor U20606 (N_20606,N_18170,N_18482);
or U20607 (N_20607,N_18827,N_18187);
nor U20608 (N_20608,N_18779,N_19418);
xor U20609 (N_20609,N_18568,N_19568);
nor U20610 (N_20610,N_19186,N_19173);
or U20611 (N_20611,N_18185,N_19949);
xor U20612 (N_20612,N_18908,N_18053);
nand U20613 (N_20613,N_19932,N_19946);
nand U20614 (N_20614,N_19530,N_18242);
nand U20615 (N_20615,N_18760,N_19219);
nor U20616 (N_20616,N_18558,N_19262);
xor U20617 (N_20617,N_19296,N_18426);
nand U20618 (N_20618,N_18975,N_19901);
xnor U20619 (N_20619,N_19475,N_18027);
or U20620 (N_20620,N_18983,N_18502);
nor U20621 (N_20621,N_19996,N_18377);
nand U20622 (N_20622,N_19016,N_18833);
and U20623 (N_20623,N_19528,N_19794);
or U20624 (N_20624,N_19044,N_19855);
nor U20625 (N_20625,N_18425,N_18524);
nand U20626 (N_20626,N_19242,N_19707);
xnor U20627 (N_20627,N_18226,N_18050);
and U20628 (N_20628,N_18952,N_19696);
nor U20629 (N_20629,N_18462,N_19232);
nor U20630 (N_20630,N_18948,N_19778);
nand U20631 (N_20631,N_18280,N_19005);
nor U20632 (N_20632,N_19921,N_18500);
or U20633 (N_20633,N_19858,N_18432);
or U20634 (N_20634,N_19484,N_18359);
nand U20635 (N_20635,N_18121,N_19203);
and U20636 (N_20636,N_19935,N_19041);
xnor U20637 (N_20637,N_18683,N_19857);
and U20638 (N_20638,N_18197,N_19841);
and U20639 (N_20639,N_18538,N_19150);
nand U20640 (N_20640,N_19435,N_18072);
nand U20641 (N_20641,N_18619,N_19621);
or U20642 (N_20642,N_18112,N_19746);
nor U20643 (N_20643,N_18757,N_19348);
or U20644 (N_20644,N_18971,N_19008);
and U20645 (N_20645,N_18584,N_19506);
xnor U20646 (N_20646,N_19931,N_18657);
nand U20647 (N_20647,N_19903,N_18533);
or U20648 (N_20648,N_18188,N_18732);
nor U20649 (N_20649,N_19669,N_19340);
nor U20650 (N_20650,N_19293,N_19397);
xnor U20651 (N_20651,N_19356,N_18045);
or U20652 (N_20652,N_19648,N_18490);
xor U20653 (N_20653,N_19074,N_18375);
or U20654 (N_20654,N_19015,N_18835);
nor U20655 (N_20655,N_19599,N_19626);
or U20656 (N_20656,N_18491,N_19320);
and U20657 (N_20657,N_18340,N_19396);
or U20658 (N_20658,N_18283,N_19849);
and U20659 (N_20659,N_18478,N_18905);
and U20660 (N_20660,N_19294,N_18842);
xnor U20661 (N_20661,N_19608,N_18211);
xnor U20662 (N_20662,N_19310,N_18182);
xor U20663 (N_20663,N_19779,N_18298);
and U20664 (N_20664,N_18633,N_18166);
nor U20665 (N_20665,N_18287,N_19357);
and U20666 (N_20666,N_19600,N_19265);
nor U20667 (N_20667,N_18839,N_18159);
or U20668 (N_20668,N_19973,N_19993);
and U20669 (N_20669,N_19791,N_18225);
or U20670 (N_20670,N_18361,N_19723);
xnor U20671 (N_20671,N_18449,N_18913);
nor U20672 (N_20672,N_18347,N_18268);
nand U20673 (N_20673,N_19101,N_19001);
nand U20674 (N_20674,N_18365,N_19206);
and U20675 (N_20675,N_18496,N_19984);
or U20676 (N_20676,N_19582,N_18945);
nand U20677 (N_20677,N_19578,N_19442);
and U20678 (N_20678,N_19405,N_18436);
and U20679 (N_20679,N_18953,N_18010);
nor U20680 (N_20680,N_19717,N_18435);
nor U20681 (N_20681,N_19140,N_18472);
and U20682 (N_20682,N_19257,N_19879);
nor U20683 (N_20683,N_19630,N_19187);
nor U20684 (N_20684,N_18635,N_18073);
xor U20685 (N_20685,N_19492,N_18198);
or U20686 (N_20686,N_18919,N_18747);
and U20687 (N_20687,N_19749,N_19248);
xor U20688 (N_20688,N_19876,N_18175);
and U20689 (N_20689,N_19799,N_18474);
and U20690 (N_20690,N_18344,N_18015);
and U20691 (N_20691,N_19472,N_18906);
xnor U20692 (N_20692,N_18057,N_19282);
nand U20693 (N_20693,N_19208,N_18612);
nor U20694 (N_20694,N_18020,N_19131);
and U20695 (N_20695,N_18587,N_18895);
or U20696 (N_20696,N_18104,N_19233);
nor U20697 (N_20697,N_19642,N_19866);
xnor U20698 (N_20698,N_18540,N_18763);
nor U20699 (N_20699,N_18677,N_18409);
and U20700 (N_20700,N_18389,N_18801);
xnor U20701 (N_20701,N_19507,N_18898);
nand U20702 (N_20702,N_19709,N_19309);
or U20703 (N_20703,N_18201,N_19420);
nor U20704 (N_20704,N_19985,N_18471);
nand U20705 (N_20705,N_19899,N_18296);
or U20706 (N_20706,N_19404,N_18281);
nor U20707 (N_20707,N_19679,N_18124);
and U20708 (N_20708,N_18370,N_18932);
nand U20709 (N_20709,N_18260,N_19704);
or U20710 (N_20710,N_18594,N_18604);
nor U20711 (N_20711,N_19115,N_18831);
or U20712 (N_20712,N_18076,N_18105);
or U20713 (N_20713,N_18578,N_18893);
and U20714 (N_20714,N_19752,N_18318);
and U20715 (N_20715,N_19830,N_19596);
xnor U20716 (N_20716,N_19549,N_19261);
nor U20717 (N_20717,N_18688,N_19292);
xnor U20718 (N_20718,N_18059,N_18640);
nor U20719 (N_20719,N_18111,N_19820);
xnor U20720 (N_20720,N_19851,N_19805);
nand U20721 (N_20721,N_18686,N_19609);
nor U20722 (N_20722,N_19280,N_18797);
or U20723 (N_20723,N_19840,N_18885);
xor U20724 (N_20724,N_18790,N_19303);
nand U20725 (N_20725,N_19942,N_18557);
nand U20726 (N_20726,N_19833,N_18315);
or U20727 (N_20727,N_18731,N_18492);
nand U20728 (N_20728,N_19038,N_18266);
nand U20729 (N_20729,N_19960,N_19345);
or U20730 (N_20730,N_18820,N_18903);
or U20731 (N_20731,N_19795,N_19068);
xor U20732 (N_20732,N_19697,N_19765);
nand U20733 (N_20733,N_19429,N_19207);
or U20734 (N_20734,N_19255,N_18303);
nand U20735 (N_20735,N_18047,N_19166);
nand U20736 (N_20736,N_19533,N_19810);
xor U20737 (N_20737,N_19317,N_18886);
or U20738 (N_20738,N_19053,N_18947);
or U20739 (N_20739,N_19613,N_18598);
nor U20740 (N_20740,N_18944,N_18590);
nor U20741 (N_20741,N_18391,N_18988);
nand U20742 (N_20742,N_18661,N_18597);
xor U20743 (N_20743,N_18276,N_18548);
nor U20744 (N_20744,N_18814,N_18774);
or U20745 (N_20745,N_18509,N_19295);
or U20746 (N_20746,N_18610,N_19694);
nor U20747 (N_20747,N_18824,N_18517);
or U20748 (N_20748,N_18148,N_19216);
nor U20749 (N_20749,N_18297,N_18532);
xor U20750 (N_20750,N_18450,N_18976);
nand U20751 (N_20751,N_18600,N_18669);
and U20752 (N_20752,N_19159,N_19056);
nand U20753 (N_20753,N_19529,N_19039);
xnor U20754 (N_20754,N_18729,N_18938);
xnor U20755 (N_20755,N_19667,N_19527);
xnor U20756 (N_20756,N_19211,N_19077);
and U20757 (N_20757,N_19266,N_19579);
and U20758 (N_20758,N_19817,N_18495);
nor U20759 (N_20759,N_18330,N_19478);
nor U20760 (N_20760,N_19324,N_19882);
nand U20761 (N_20761,N_18350,N_18353);
nor U20762 (N_20762,N_18213,N_19560);
nand U20763 (N_20763,N_19196,N_18243);
xor U20764 (N_20764,N_19381,N_18641);
nand U20765 (N_20765,N_19922,N_19479);
or U20766 (N_20766,N_18299,N_18454);
nand U20767 (N_20767,N_18103,N_19641);
xnor U20768 (N_20768,N_18643,N_18453);
nand U20769 (N_20769,N_18543,N_18044);
or U20770 (N_20770,N_19192,N_18151);
xnor U20771 (N_20771,N_19455,N_18334);
and U20772 (N_20772,N_18551,N_19948);
nand U20773 (N_20773,N_19939,N_19874);
nor U20774 (N_20774,N_19402,N_18231);
xor U20775 (N_20775,N_19947,N_19002);
nand U20776 (N_20776,N_19505,N_18847);
and U20777 (N_20777,N_19593,N_18163);
nor U20778 (N_20778,N_18951,N_18853);
nand U20779 (N_20779,N_18651,N_19967);
xor U20780 (N_20780,N_18690,N_19963);
xor U20781 (N_20781,N_19277,N_19314);
and U20782 (N_20782,N_18431,N_19606);
and U20783 (N_20783,N_19132,N_19536);
nor U20784 (N_20784,N_19509,N_18405);
and U20785 (N_20785,N_19407,N_19463);
nand U20786 (N_20786,N_19380,N_19798);
and U20787 (N_20787,N_18255,N_19347);
nand U20788 (N_20788,N_19610,N_19617);
or U20789 (N_20789,N_18868,N_19742);
nand U20790 (N_20790,N_19358,N_19726);
nand U20791 (N_20791,N_19733,N_19286);
xnor U20792 (N_20792,N_18085,N_18141);
or U20793 (N_20793,N_19047,N_18984);
and U20794 (N_20794,N_19133,N_18660);
nand U20795 (N_20795,N_18207,N_19204);
xor U20796 (N_20796,N_18019,N_18245);
and U20797 (N_20797,N_19096,N_19316);
or U20798 (N_20798,N_18304,N_18884);
or U20799 (N_20799,N_19431,N_19548);
and U20800 (N_20800,N_18316,N_18784);
nor U20801 (N_20801,N_18679,N_19069);
and U20802 (N_20802,N_19796,N_19891);
or U20803 (N_20803,N_18691,N_18787);
or U20804 (N_20804,N_18642,N_18267);
or U20805 (N_20805,N_18521,N_19321);
xnor U20806 (N_20806,N_19195,N_18459);
xor U20807 (N_20807,N_19108,N_19938);
nand U20808 (N_20808,N_18812,N_19487);
and U20809 (N_20809,N_18752,N_19902);
xnor U20810 (N_20810,N_19773,N_19411);
xnor U20811 (N_20811,N_18792,N_19975);
nand U20812 (N_20812,N_19415,N_18864);
and U20813 (N_20813,N_18102,N_19226);
and U20814 (N_20814,N_19553,N_19419);
nor U20815 (N_20815,N_18423,N_19826);
nor U20816 (N_20816,N_19822,N_18601);
xnor U20817 (N_20817,N_18123,N_19043);
xnor U20818 (N_20818,N_18064,N_18394);
nand U20819 (N_20819,N_19842,N_19639);
nand U20820 (N_20820,N_18544,N_19147);
nor U20821 (N_20821,N_18013,N_19580);
or U20822 (N_20822,N_18133,N_19306);
nor U20823 (N_20823,N_18539,N_18049);
nand U20824 (N_20824,N_18039,N_18770);
nand U20825 (N_20825,N_18168,N_19686);
nand U20826 (N_20826,N_18172,N_19770);
xor U20827 (N_20827,N_19900,N_18569);
nand U20828 (N_20828,N_19535,N_19278);
or U20829 (N_20829,N_19687,N_19086);
nand U20830 (N_20830,N_18379,N_18917);
nand U20831 (N_20831,N_18711,N_19588);
nand U20832 (N_20832,N_18274,N_19571);
nor U20833 (N_20833,N_18805,N_18508);
or U20834 (N_20834,N_18700,N_18708);
nand U20835 (N_20835,N_18390,N_19871);
nand U20836 (N_20836,N_19352,N_19929);
xor U20837 (N_20837,N_19700,N_19873);
nor U20838 (N_20838,N_19587,N_18241);
and U20839 (N_20839,N_18576,N_19616);
or U20840 (N_20840,N_19033,N_18203);
nand U20841 (N_20841,N_19520,N_18552);
nor U20842 (N_20842,N_18916,N_19583);
or U20843 (N_20843,N_18239,N_18900);
nor U20844 (N_20844,N_18545,N_19276);
and U20845 (N_20845,N_18652,N_19982);
nor U20846 (N_20846,N_18254,N_18437);
and U20847 (N_20847,N_18709,N_19839);
xnor U20848 (N_20848,N_18809,N_19440);
nor U20849 (N_20849,N_18672,N_19741);
or U20850 (N_20850,N_19480,N_18662);
nand U20851 (N_20851,N_18305,N_18169);
or U20852 (N_20852,N_19176,N_18186);
or U20853 (N_20853,N_19427,N_19561);
or U20854 (N_20854,N_19236,N_18263);
and U20855 (N_20855,N_19692,N_19540);
nor U20856 (N_20856,N_18295,N_19498);
and U20857 (N_20857,N_19682,N_19482);
nor U20858 (N_20858,N_18354,N_19212);
nand U20859 (N_20859,N_19471,N_18401);
or U20860 (N_20860,N_19877,N_19698);
xor U20861 (N_20861,N_18095,N_18360);
and U20862 (N_20862,N_18325,N_18715);
or U20863 (N_20863,N_19067,N_19782);
or U20864 (N_20864,N_19790,N_19240);
xnor U20865 (N_20865,N_19290,N_19142);
and U20866 (N_20866,N_19624,N_19918);
or U20867 (N_20867,N_19766,N_18712);
nor U20868 (N_20868,N_19792,N_18659);
and U20869 (N_20869,N_19567,N_18167);
xnor U20870 (N_20870,N_19164,N_19445);
and U20871 (N_20871,N_19980,N_18855);
or U20872 (N_20872,N_18869,N_18503);
and U20873 (N_20873,N_18862,N_19289);
or U20874 (N_20874,N_19055,N_18028);
or U20875 (N_20875,N_18719,N_18265);
and U20876 (N_20876,N_19564,N_18062);
xnor U20877 (N_20877,N_18526,N_18996);
nor U20878 (N_20878,N_18888,N_19416);
nand U20879 (N_20879,N_18180,N_19941);
xor U20880 (N_20880,N_19213,N_19594);
nor U20881 (N_20881,N_18476,N_19394);
xor U20882 (N_20882,N_19300,N_19158);
and U20883 (N_20883,N_19274,N_18140);
or U20884 (N_20884,N_19019,N_19465);
nand U20885 (N_20885,N_19003,N_18663);
xor U20886 (N_20886,N_18376,N_19691);
nand U20887 (N_20887,N_18084,N_18586);
nor U20888 (N_20888,N_19724,N_18058);
and U20889 (N_20889,N_18892,N_18856);
and U20890 (N_20890,N_19783,N_18128);
or U20891 (N_20891,N_18319,N_18380);
and U20892 (N_20892,N_19591,N_18514);
and U20893 (N_20893,N_18993,N_18342);
and U20894 (N_20894,N_18527,N_19661);
and U20895 (N_20895,N_18881,N_19319);
and U20896 (N_20896,N_18699,N_18950);
or U20897 (N_20897,N_19581,N_19601);
or U20898 (N_20898,N_18367,N_19887);
nand U20899 (N_20899,N_18160,N_19771);
nor U20900 (N_20900,N_19383,N_18117);
nand U20901 (N_20901,N_19714,N_18311);
or U20902 (N_20902,N_18004,N_19454);
nand U20903 (N_20903,N_19353,N_19754);
and U20904 (N_20904,N_19066,N_18277);
nor U20905 (N_20905,N_19913,N_19738);
or U20906 (N_20906,N_19337,N_18675);
or U20907 (N_20907,N_19775,N_19914);
xor U20908 (N_20908,N_18562,N_19256);
and U20909 (N_20909,N_19886,N_18055);
xnor U20910 (N_20910,N_18343,N_19417);
nor U20911 (N_20911,N_18386,N_19307);
or U20912 (N_20912,N_19756,N_19308);
xor U20913 (N_20913,N_18366,N_19850);
nor U20914 (N_20914,N_18954,N_18016);
and U20915 (N_20915,N_19744,N_18621);
xnor U20916 (N_20916,N_19200,N_18822);
nand U20917 (N_20917,N_19331,N_18456);
or U20918 (N_20918,N_18664,N_19499);
and U20919 (N_20919,N_18461,N_18264);
nand U20920 (N_20920,N_18904,N_19715);
xnor U20921 (N_20921,N_18282,N_19786);
nand U20922 (N_20922,N_19374,N_19961);
nor U20923 (N_20923,N_19676,N_18701);
or U20924 (N_20924,N_18922,N_19751);
or U20925 (N_20925,N_18021,N_19151);
xor U20926 (N_20926,N_19432,N_19878);
nor U20927 (N_20927,N_19534,N_19777);
xnor U20928 (N_20928,N_19491,N_19959);
nor U20929 (N_20929,N_19678,N_19486);
nand U20930 (N_20930,N_18399,N_18429);
or U20931 (N_20931,N_19896,N_18843);
nor U20932 (N_20932,N_18336,N_18934);
and U20933 (N_20933,N_19566,N_18145);
nor U20934 (N_20934,N_18724,N_19149);
or U20935 (N_20935,N_19875,N_18489);
xnor U20936 (N_20936,N_19006,N_18510);
xor U20937 (N_20937,N_18369,N_19666);
nand U20938 (N_20938,N_19881,N_18707);
nor U20939 (N_20939,N_19329,N_18493);
or U20940 (N_20940,N_18237,N_19684);
nor U20941 (N_20941,N_18486,N_19049);
nand U20942 (N_20942,N_18106,N_18383);
nand U20943 (N_20943,N_19494,N_18570);
and U20944 (N_20944,N_19847,N_18009);
xor U20945 (N_20945,N_19048,N_19220);
and U20946 (N_20946,N_18421,N_19438);
and U20947 (N_20947,N_18899,N_19092);
nor U20948 (N_20948,N_19228,N_18512);
xnor U20949 (N_20949,N_18902,N_19550);
or U20950 (N_20950,N_19660,N_18530);
nand U20951 (N_20951,N_19064,N_18946);
nor U20952 (N_20952,N_19940,N_18997);
nor U20953 (N_20953,N_19909,N_19930);
or U20954 (N_20954,N_19476,N_18838);
or U20955 (N_20955,N_18909,N_18890);
and U20956 (N_20956,N_19937,N_19264);
or U20957 (N_20957,N_19027,N_19330);
nor U20958 (N_20958,N_18395,N_18191);
or U20959 (N_20959,N_18713,N_19121);
or U20960 (N_20960,N_18116,N_19202);
nand U20961 (N_20961,N_19807,N_19657);
nand U20962 (N_20962,N_18681,N_19281);
nor U20963 (N_20963,N_18722,N_18022);
nor U20964 (N_20964,N_19215,N_19500);
xor U20965 (N_20965,N_19898,N_19597);
or U20966 (N_20966,N_19885,N_18382);
xnor U20967 (N_20967,N_18977,N_19235);
and U20968 (N_20968,N_18730,N_18969);
nand U20969 (N_20969,N_19354,N_19099);
and U20970 (N_20970,N_19456,N_18703);
nand U20971 (N_20971,N_19991,N_18107);
nor U20972 (N_20972,N_18915,N_19007);
xnor U20973 (N_20973,N_19664,N_18223);
nand U20974 (N_20974,N_19721,N_19646);
nand U20975 (N_20975,N_18355,N_18959);
xnor U20976 (N_20976,N_19671,N_19523);
and U20977 (N_20977,N_19674,N_18233);
nand U20978 (N_20978,N_19954,N_19288);
nand U20979 (N_20979,N_19701,N_19673);
xnor U20980 (N_20980,N_19649,N_19703);
and U20981 (N_20981,N_18861,N_19636);
or U20982 (N_20982,N_19114,N_18181);
nor U20983 (N_20983,N_19925,N_19539);
nor U20984 (N_20984,N_18238,N_18958);
xor U20985 (N_20985,N_18189,N_18329);
nand U20986 (N_20986,N_18439,N_18697);
nor U20987 (N_20987,N_19759,N_18671);
nor U20988 (N_20988,N_19502,N_19021);
or U20989 (N_20989,N_19743,N_19365);
xor U20990 (N_20990,N_18078,N_19607);
nand U20991 (N_20991,N_18244,N_18667);
nand U20992 (N_20992,N_18823,N_18788);
or U20993 (N_20993,N_18136,N_19911);
xnor U20994 (N_20994,N_18417,N_19304);
nand U20995 (N_20995,N_19379,N_19464);
xor U20996 (N_20996,N_19018,N_19774);
xor U20997 (N_20997,N_18464,N_18052);
nand U20998 (N_20998,N_18406,N_19378);
nor U20999 (N_20999,N_18271,N_19045);
nand U21000 (N_21000,N_19612,N_19362);
and U21001 (N_21001,N_19179,N_19681);
nand U21002 (N_21002,N_19298,N_19552);
or U21003 (N_21003,N_19371,N_18349);
and U21004 (N_21004,N_19714,N_18233);
nor U21005 (N_21005,N_19835,N_19190);
and U21006 (N_21006,N_19034,N_18031);
and U21007 (N_21007,N_19679,N_19417);
nor U21008 (N_21008,N_18270,N_18806);
or U21009 (N_21009,N_19437,N_19418);
xnor U21010 (N_21010,N_19832,N_19625);
xnor U21011 (N_21011,N_19080,N_18244);
nor U21012 (N_21012,N_18510,N_19575);
and U21013 (N_21013,N_18852,N_18726);
nor U21014 (N_21014,N_18064,N_18063);
xor U21015 (N_21015,N_19140,N_18853);
nand U21016 (N_21016,N_19279,N_19792);
nand U21017 (N_21017,N_19620,N_18127);
or U21018 (N_21018,N_18624,N_18755);
nor U21019 (N_21019,N_18836,N_18692);
nand U21020 (N_21020,N_19950,N_19986);
nor U21021 (N_21021,N_19029,N_18880);
or U21022 (N_21022,N_19931,N_18044);
xor U21023 (N_21023,N_18837,N_18662);
nor U21024 (N_21024,N_18140,N_18564);
or U21025 (N_21025,N_19660,N_18199);
or U21026 (N_21026,N_19755,N_19764);
and U21027 (N_21027,N_18966,N_19881);
or U21028 (N_21028,N_18458,N_19751);
and U21029 (N_21029,N_18481,N_19246);
nand U21030 (N_21030,N_18825,N_19367);
and U21031 (N_21031,N_19104,N_18810);
nor U21032 (N_21032,N_18763,N_18660);
nor U21033 (N_21033,N_18943,N_19782);
nand U21034 (N_21034,N_19912,N_18361);
or U21035 (N_21035,N_19250,N_18930);
nor U21036 (N_21036,N_19607,N_19526);
and U21037 (N_21037,N_18419,N_19126);
nand U21038 (N_21038,N_19535,N_18414);
nand U21039 (N_21039,N_18758,N_19199);
nand U21040 (N_21040,N_18882,N_19646);
nand U21041 (N_21041,N_18791,N_19055);
and U21042 (N_21042,N_19945,N_19820);
or U21043 (N_21043,N_18133,N_18753);
xor U21044 (N_21044,N_19344,N_19361);
and U21045 (N_21045,N_19755,N_18749);
nor U21046 (N_21046,N_18446,N_19716);
nand U21047 (N_21047,N_19961,N_18006);
xnor U21048 (N_21048,N_19086,N_19720);
nand U21049 (N_21049,N_19792,N_19984);
and U21050 (N_21050,N_19716,N_18009);
nand U21051 (N_21051,N_19318,N_19478);
nor U21052 (N_21052,N_18248,N_19498);
or U21053 (N_21053,N_19731,N_18789);
and U21054 (N_21054,N_18576,N_18472);
nand U21055 (N_21055,N_18112,N_18651);
or U21056 (N_21056,N_19246,N_18149);
nor U21057 (N_21057,N_18376,N_18862);
xor U21058 (N_21058,N_18097,N_18651);
nand U21059 (N_21059,N_19873,N_19433);
xor U21060 (N_21060,N_18250,N_19333);
nor U21061 (N_21061,N_18469,N_18626);
and U21062 (N_21062,N_18185,N_19602);
nor U21063 (N_21063,N_18787,N_18729);
nand U21064 (N_21064,N_18587,N_19315);
nand U21065 (N_21065,N_19851,N_18894);
and U21066 (N_21066,N_19011,N_18823);
nand U21067 (N_21067,N_18579,N_19174);
and U21068 (N_21068,N_19071,N_19453);
or U21069 (N_21069,N_18402,N_19794);
and U21070 (N_21070,N_18237,N_18151);
xnor U21071 (N_21071,N_18057,N_19353);
and U21072 (N_21072,N_18355,N_19515);
xor U21073 (N_21073,N_19124,N_19854);
nor U21074 (N_21074,N_19981,N_18783);
nor U21075 (N_21075,N_19985,N_19396);
and U21076 (N_21076,N_19173,N_18249);
xor U21077 (N_21077,N_18381,N_19236);
and U21078 (N_21078,N_18690,N_19485);
or U21079 (N_21079,N_19109,N_18817);
and U21080 (N_21080,N_19287,N_19150);
and U21081 (N_21081,N_18077,N_18050);
xnor U21082 (N_21082,N_18479,N_19147);
xnor U21083 (N_21083,N_19948,N_19555);
and U21084 (N_21084,N_19356,N_19929);
nor U21085 (N_21085,N_18566,N_19437);
nand U21086 (N_21086,N_18454,N_19868);
or U21087 (N_21087,N_18909,N_18221);
nand U21088 (N_21088,N_19600,N_18739);
xnor U21089 (N_21089,N_18398,N_19391);
or U21090 (N_21090,N_19753,N_18804);
and U21091 (N_21091,N_19018,N_18358);
xnor U21092 (N_21092,N_19091,N_18257);
xor U21093 (N_21093,N_19757,N_18913);
xnor U21094 (N_21094,N_19204,N_19175);
and U21095 (N_21095,N_19118,N_19375);
xnor U21096 (N_21096,N_18961,N_19086);
nand U21097 (N_21097,N_19000,N_18020);
xor U21098 (N_21098,N_19510,N_19277);
nand U21099 (N_21099,N_19439,N_18680);
nand U21100 (N_21100,N_18646,N_19728);
or U21101 (N_21101,N_18954,N_19368);
and U21102 (N_21102,N_19926,N_18820);
and U21103 (N_21103,N_19577,N_19156);
xnor U21104 (N_21104,N_18475,N_18067);
or U21105 (N_21105,N_18507,N_19885);
or U21106 (N_21106,N_18889,N_18780);
nand U21107 (N_21107,N_18384,N_18935);
xnor U21108 (N_21108,N_19993,N_19703);
nor U21109 (N_21109,N_19102,N_18135);
nor U21110 (N_21110,N_19922,N_19359);
or U21111 (N_21111,N_18592,N_18695);
and U21112 (N_21112,N_19757,N_18536);
or U21113 (N_21113,N_19911,N_19185);
xor U21114 (N_21114,N_19723,N_19080);
or U21115 (N_21115,N_18671,N_19536);
nand U21116 (N_21116,N_19760,N_18271);
nor U21117 (N_21117,N_18668,N_18807);
and U21118 (N_21118,N_19790,N_19112);
or U21119 (N_21119,N_19451,N_18338);
or U21120 (N_21120,N_19155,N_18526);
or U21121 (N_21121,N_19742,N_19347);
xor U21122 (N_21122,N_19495,N_18844);
and U21123 (N_21123,N_19638,N_19207);
nor U21124 (N_21124,N_18141,N_19598);
nand U21125 (N_21125,N_18113,N_18706);
and U21126 (N_21126,N_19221,N_18374);
nand U21127 (N_21127,N_18208,N_18257);
xnor U21128 (N_21128,N_19951,N_18890);
and U21129 (N_21129,N_19822,N_18033);
xor U21130 (N_21130,N_19877,N_19478);
or U21131 (N_21131,N_19110,N_19593);
nor U21132 (N_21132,N_19904,N_19802);
and U21133 (N_21133,N_19524,N_18217);
nor U21134 (N_21134,N_18702,N_18226);
or U21135 (N_21135,N_18420,N_18494);
or U21136 (N_21136,N_18752,N_19945);
nand U21137 (N_21137,N_18157,N_19333);
or U21138 (N_21138,N_18478,N_18257);
xor U21139 (N_21139,N_18750,N_18616);
nor U21140 (N_21140,N_19906,N_18855);
and U21141 (N_21141,N_18656,N_18951);
xnor U21142 (N_21142,N_18778,N_19844);
or U21143 (N_21143,N_18965,N_19739);
or U21144 (N_21144,N_18881,N_19989);
nor U21145 (N_21145,N_19485,N_18763);
and U21146 (N_21146,N_19228,N_19109);
xor U21147 (N_21147,N_19828,N_19571);
xnor U21148 (N_21148,N_18424,N_18290);
and U21149 (N_21149,N_19689,N_18597);
nor U21150 (N_21150,N_19793,N_19268);
nand U21151 (N_21151,N_19548,N_19580);
xnor U21152 (N_21152,N_18546,N_19821);
nand U21153 (N_21153,N_18548,N_19014);
xor U21154 (N_21154,N_18735,N_19110);
and U21155 (N_21155,N_19270,N_19293);
xnor U21156 (N_21156,N_18985,N_19363);
nand U21157 (N_21157,N_19836,N_19809);
or U21158 (N_21158,N_18450,N_18908);
xnor U21159 (N_21159,N_18546,N_19461);
nand U21160 (N_21160,N_19802,N_19126);
and U21161 (N_21161,N_18222,N_18691);
nand U21162 (N_21162,N_19111,N_18667);
nor U21163 (N_21163,N_19869,N_19917);
nand U21164 (N_21164,N_19629,N_18482);
xnor U21165 (N_21165,N_18240,N_18292);
nand U21166 (N_21166,N_18059,N_18491);
xnor U21167 (N_21167,N_19319,N_19178);
xor U21168 (N_21168,N_18264,N_18012);
and U21169 (N_21169,N_19791,N_19829);
xnor U21170 (N_21170,N_19586,N_18574);
or U21171 (N_21171,N_18472,N_18894);
or U21172 (N_21172,N_19830,N_19710);
and U21173 (N_21173,N_18071,N_18495);
and U21174 (N_21174,N_19444,N_18760);
and U21175 (N_21175,N_18038,N_19256);
xor U21176 (N_21176,N_18035,N_19691);
and U21177 (N_21177,N_18749,N_19883);
nor U21178 (N_21178,N_19366,N_19893);
nor U21179 (N_21179,N_19498,N_19270);
nand U21180 (N_21180,N_19968,N_19282);
and U21181 (N_21181,N_19532,N_18965);
xor U21182 (N_21182,N_19589,N_19559);
nand U21183 (N_21183,N_19692,N_19355);
or U21184 (N_21184,N_18961,N_18740);
or U21185 (N_21185,N_18736,N_18768);
xor U21186 (N_21186,N_19231,N_18485);
nand U21187 (N_21187,N_18575,N_19522);
and U21188 (N_21188,N_19073,N_19781);
nor U21189 (N_21189,N_18808,N_18706);
xor U21190 (N_21190,N_19755,N_18033);
or U21191 (N_21191,N_19001,N_19436);
and U21192 (N_21192,N_19938,N_19262);
nand U21193 (N_21193,N_19190,N_19078);
and U21194 (N_21194,N_19404,N_18458);
nor U21195 (N_21195,N_19854,N_19585);
and U21196 (N_21196,N_19908,N_18596);
xnor U21197 (N_21197,N_18446,N_19452);
nand U21198 (N_21198,N_19784,N_19379);
xnor U21199 (N_21199,N_18432,N_18078);
and U21200 (N_21200,N_18547,N_18865);
or U21201 (N_21201,N_18852,N_18633);
nor U21202 (N_21202,N_18305,N_19276);
and U21203 (N_21203,N_18115,N_19715);
nand U21204 (N_21204,N_19686,N_19999);
xor U21205 (N_21205,N_18104,N_18614);
nand U21206 (N_21206,N_19467,N_18328);
xor U21207 (N_21207,N_19857,N_18193);
or U21208 (N_21208,N_18949,N_18567);
nand U21209 (N_21209,N_18374,N_19971);
nor U21210 (N_21210,N_19469,N_19521);
or U21211 (N_21211,N_18694,N_18151);
nor U21212 (N_21212,N_19907,N_19402);
xnor U21213 (N_21213,N_19796,N_19327);
nand U21214 (N_21214,N_18634,N_19436);
nand U21215 (N_21215,N_18728,N_19956);
nor U21216 (N_21216,N_19240,N_19671);
or U21217 (N_21217,N_18149,N_18478);
or U21218 (N_21218,N_18512,N_18950);
nor U21219 (N_21219,N_19112,N_19570);
or U21220 (N_21220,N_18544,N_18912);
and U21221 (N_21221,N_18897,N_18834);
xnor U21222 (N_21222,N_18527,N_19775);
nor U21223 (N_21223,N_18218,N_18773);
nand U21224 (N_21224,N_18507,N_19702);
nor U21225 (N_21225,N_19533,N_19832);
nand U21226 (N_21226,N_19229,N_19964);
nor U21227 (N_21227,N_19348,N_18531);
nand U21228 (N_21228,N_18466,N_18276);
nand U21229 (N_21229,N_18310,N_18932);
nand U21230 (N_21230,N_19192,N_18847);
nor U21231 (N_21231,N_19882,N_19092);
nor U21232 (N_21232,N_18699,N_18338);
and U21233 (N_21233,N_19431,N_18165);
and U21234 (N_21234,N_19023,N_18406);
nand U21235 (N_21235,N_19766,N_19788);
or U21236 (N_21236,N_19869,N_18015);
or U21237 (N_21237,N_18769,N_18780);
xnor U21238 (N_21238,N_19676,N_18841);
and U21239 (N_21239,N_18613,N_18745);
or U21240 (N_21240,N_19081,N_19979);
xnor U21241 (N_21241,N_18099,N_18163);
nand U21242 (N_21242,N_19343,N_18036);
nor U21243 (N_21243,N_18554,N_18043);
or U21244 (N_21244,N_18537,N_19138);
and U21245 (N_21245,N_18420,N_18053);
and U21246 (N_21246,N_18724,N_19169);
nand U21247 (N_21247,N_18320,N_19152);
and U21248 (N_21248,N_18581,N_19470);
and U21249 (N_21249,N_18803,N_18942);
nand U21250 (N_21250,N_19657,N_19088);
nand U21251 (N_21251,N_18917,N_18260);
or U21252 (N_21252,N_19932,N_18694);
nor U21253 (N_21253,N_19580,N_18282);
and U21254 (N_21254,N_18102,N_19319);
nor U21255 (N_21255,N_18240,N_18044);
xor U21256 (N_21256,N_19873,N_18899);
nor U21257 (N_21257,N_19282,N_18490);
and U21258 (N_21258,N_19880,N_19983);
nand U21259 (N_21259,N_18560,N_19006);
nor U21260 (N_21260,N_19627,N_19952);
or U21261 (N_21261,N_18069,N_18169);
or U21262 (N_21262,N_19460,N_19832);
nand U21263 (N_21263,N_18164,N_18132);
nor U21264 (N_21264,N_19384,N_19347);
nor U21265 (N_21265,N_18700,N_18452);
xor U21266 (N_21266,N_19940,N_18803);
nor U21267 (N_21267,N_19999,N_18314);
nand U21268 (N_21268,N_18492,N_18275);
or U21269 (N_21269,N_18089,N_18105);
and U21270 (N_21270,N_18193,N_18035);
nor U21271 (N_21271,N_18074,N_19149);
nand U21272 (N_21272,N_19455,N_19019);
xnor U21273 (N_21273,N_18279,N_18408);
nor U21274 (N_21274,N_19419,N_18433);
nand U21275 (N_21275,N_19947,N_18115);
and U21276 (N_21276,N_19401,N_19051);
nor U21277 (N_21277,N_19678,N_19919);
or U21278 (N_21278,N_19086,N_19148);
nor U21279 (N_21279,N_19956,N_19218);
and U21280 (N_21280,N_18968,N_18536);
or U21281 (N_21281,N_18205,N_19412);
xnor U21282 (N_21282,N_19991,N_19337);
or U21283 (N_21283,N_19487,N_19687);
and U21284 (N_21284,N_18918,N_19054);
xor U21285 (N_21285,N_19809,N_19546);
nor U21286 (N_21286,N_18597,N_19965);
or U21287 (N_21287,N_18424,N_19526);
and U21288 (N_21288,N_19153,N_19106);
or U21289 (N_21289,N_18350,N_18014);
and U21290 (N_21290,N_18866,N_18634);
or U21291 (N_21291,N_19007,N_18994);
nand U21292 (N_21292,N_18361,N_19892);
or U21293 (N_21293,N_19722,N_18923);
xor U21294 (N_21294,N_18790,N_18807);
nor U21295 (N_21295,N_19108,N_19433);
or U21296 (N_21296,N_18464,N_19540);
xnor U21297 (N_21297,N_18818,N_19890);
nor U21298 (N_21298,N_19796,N_19264);
and U21299 (N_21299,N_18889,N_19217);
nand U21300 (N_21300,N_18066,N_18799);
and U21301 (N_21301,N_18062,N_18069);
xnor U21302 (N_21302,N_18669,N_18980);
and U21303 (N_21303,N_18903,N_19985);
and U21304 (N_21304,N_18764,N_19649);
or U21305 (N_21305,N_18102,N_19474);
xor U21306 (N_21306,N_19680,N_18022);
or U21307 (N_21307,N_18978,N_19572);
and U21308 (N_21308,N_19810,N_19545);
nor U21309 (N_21309,N_19246,N_19472);
xnor U21310 (N_21310,N_18396,N_19047);
nand U21311 (N_21311,N_18727,N_19306);
nand U21312 (N_21312,N_18359,N_18168);
xnor U21313 (N_21313,N_19356,N_19277);
xnor U21314 (N_21314,N_18086,N_18527);
nor U21315 (N_21315,N_18283,N_19518);
nand U21316 (N_21316,N_18880,N_18366);
nor U21317 (N_21317,N_18692,N_18650);
nand U21318 (N_21318,N_19810,N_19910);
and U21319 (N_21319,N_19030,N_19790);
nand U21320 (N_21320,N_19173,N_19250);
nor U21321 (N_21321,N_18899,N_18760);
xnor U21322 (N_21322,N_19106,N_18295);
nand U21323 (N_21323,N_19681,N_19630);
or U21324 (N_21324,N_18827,N_18648);
nand U21325 (N_21325,N_18324,N_19597);
and U21326 (N_21326,N_18575,N_18174);
xnor U21327 (N_21327,N_18460,N_19765);
nor U21328 (N_21328,N_19498,N_19016);
and U21329 (N_21329,N_18600,N_18241);
and U21330 (N_21330,N_18782,N_18759);
xnor U21331 (N_21331,N_18024,N_19398);
nor U21332 (N_21332,N_19022,N_18225);
nor U21333 (N_21333,N_19300,N_18448);
nor U21334 (N_21334,N_18884,N_19494);
nor U21335 (N_21335,N_19959,N_18287);
and U21336 (N_21336,N_19137,N_18971);
nor U21337 (N_21337,N_19936,N_19053);
nand U21338 (N_21338,N_18382,N_19205);
or U21339 (N_21339,N_19272,N_19648);
and U21340 (N_21340,N_19595,N_18313);
and U21341 (N_21341,N_19751,N_19573);
or U21342 (N_21342,N_19362,N_19241);
or U21343 (N_21343,N_18635,N_19368);
nand U21344 (N_21344,N_18166,N_19548);
nand U21345 (N_21345,N_18711,N_18305);
nand U21346 (N_21346,N_18079,N_19878);
and U21347 (N_21347,N_18905,N_19883);
xnor U21348 (N_21348,N_18178,N_19582);
nand U21349 (N_21349,N_19012,N_19274);
nor U21350 (N_21350,N_19851,N_18131);
xnor U21351 (N_21351,N_19838,N_18560);
xor U21352 (N_21352,N_19704,N_18199);
nor U21353 (N_21353,N_19280,N_18978);
or U21354 (N_21354,N_19290,N_19648);
nor U21355 (N_21355,N_19621,N_18896);
and U21356 (N_21356,N_19299,N_18389);
nor U21357 (N_21357,N_18738,N_18369);
nor U21358 (N_21358,N_19546,N_19970);
nor U21359 (N_21359,N_19845,N_19784);
nand U21360 (N_21360,N_18383,N_19440);
and U21361 (N_21361,N_19553,N_19204);
or U21362 (N_21362,N_18799,N_19800);
or U21363 (N_21363,N_19491,N_18979);
xnor U21364 (N_21364,N_18122,N_18594);
nor U21365 (N_21365,N_18894,N_19623);
nor U21366 (N_21366,N_19577,N_19821);
nand U21367 (N_21367,N_19644,N_18065);
and U21368 (N_21368,N_19367,N_18028);
nor U21369 (N_21369,N_19022,N_18431);
nand U21370 (N_21370,N_19516,N_18381);
xor U21371 (N_21371,N_19276,N_19928);
nor U21372 (N_21372,N_19038,N_18929);
and U21373 (N_21373,N_18589,N_18994);
and U21374 (N_21374,N_19394,N_19374);
nor U21375 (N_21375,N_18005,N_19369);
and U21376 (N_21376,N_19007,N_18443);
nand U21377 (N_21377,N_18168,N_18607);
nor U21378 (N_21378,N_18496,N_18607);
and U21379 (N_21379,N_18514,N_18820);
or U21380 (N_21380,N_18829,N_19679);
nand U21381 (N_21381,N_18993,N_18322);
xnor U21382 (N_21382,N_18548,N_19407);
nand U21383 (N_21383,N_19078,N_19262);
nand U21384 (N_21384,N_18577,N_18494);
nand U21385 (N_21385,N_19536,N_19103);
or U21386 (N_21386,N_18863,N_18674);
xor U21387 (N_21387,N_19517,N_19482);
nor U21388 (N_21388,N_18334,N_18329);
xor U21389 (N_21389,N_19716,N_19619);
xnor U21390 (N_21390,N_18896,N_18427);
nand U21391 (N_21391,N_19697,N_18792);
and U21392 (N_21392,N_19228,N_18768);
xnor U21393 (N_21393,N_18783,N_18925);
nand U21394 (N_21394,N_18479,N_19762);
nor U21395 (N_21395,N_19943,N_18666);
xor U21396 (N_21396,N_19808,N_19403);
or U21397 (N_21397,N_18977,N_19497);
or U21398 (N_21398,N_18587,N_18317);
nand U21399 (N_21399,N_18948,N_19862);
and U21400 (N_21400,N_18824,N_18905);
or U21401 (N_21401,N_18588,N_18690);
nand U21402 (N_21402,N_18347,N_18407);
nand U21403 (N_21403,N_19567,N_19666);
nor U21404 (N_21404,N_18220,N_18945);
and U21405 (N_21405,N_18161,N_19327);
or U21406 (N_21406,N_19113,N_18342);
or U21407 (N_21407,N_19080,N_18836);
nor U21408 (N_21408,N_19818,N_18467);
nor U21409 (N_21409,N_19199,N_19784);
nand U21410 (N_21410,N_18046,N_18268);
nor U21411 (N_21411,N_18652,N_18285);
xor U21412 (N_21412,N_19554,N_19598);
and U21413 (N_21413,N_19579,N_18537);
nand U21414 (N_21414,N_19064,N_19330);
nor U21415 (N_21415,N_19567,N_18717);
nand U21416 (N_21416,N_19408,N_18509);
nand U21417 (N_21417,N_19095,N_19401);
or U21418 (N_21418,N_19989,N_18498);
xor U21419 (N_21419,N_19878,N_18478);
xor U21420 (N_21420,N_19609,N_18894);
nor U21421 (N_21421,N_18097,N_18853);
or U21422 (N_21422,N_19733,N_18847);
xor U21423 (N_21423,N_18166,N_19240);
nor U21424 (N_21424,N_18870,N_18500);
xor U21425 (N_21425,N_18460,N_19161);
or U21426 (N_21426,N_18781,N_18445);
and U21427 (N_21427,N_19134,N_19265);
or U21428 (N_21428,N_18686,N_18583);
nand U21429 (N_21429,N_18612,N_18275);
nor U21430 (N_21430,N_18477,N_18311);
xor U21431 (N_21431,N_18080,N_18239);
nand U21432 (N_21432,N_19232,N_19360);
nor U21433 (N_21433,N_18381,N_18560);
and U21434 (N_21434,N_18519,N_18602);
and U21435 (N_21435,N_18514,N_18417);
and U21436 (N_21436,N_18806,N_19633);
xnor U21437 (N_21437,N_18207,N_19514);
or U21438 (N_21438,N_18699,N_18284);
and U21439 (N_21439,N_19698,N_18400);
and U21440 (N_21440,N_19213,N_19499);
and U21441 (N_21441,N_19349,N_19509);
nor U21442 (N_21442,N_19461,N_19595);
nand U21443 (N_21443,N_19487,N_19209);
nor U21444 (N_21444,N_18222,N_18814);
and U21445 (N_21445,N_18930,N_19682);
and U21446 (N_21446,N_18016,N_18655);
xor U21447 (N_21447,N_18522,N_18271);
and U21448 (N_21448,N_19775,N_19744);
or U21449 (N_21449,N_18458,N_19831);
xnor U21450 (N_21450,N_19446,N_18231);
xnor U21451 (N_21451,N_18543,N_19309);
and U21452 (N_21452,N_18778,N_19327);
nand U21453 (N_21453,N_19474,N_18751);
xor U21454 (N_21454,N_18751,N_18634);
nand U21455 (N_21455,N_18872,N_19201);
or U21456 (N_21456,N_19440,N_18199);
nor U21457 (N_21457,N_19322,N_18526);
nand U21458 (N_21458,N_19049,N_18035);
nand U21459 (N_21459,N_19794,N_19576);
xor U21460 (N_21460,N_19338,N_18647);
or U21461 (N_21461,N_19521,N_18724);
or U21462 (N_21462,N_18677,N_18294);
or U21463 (N_21463,N_19091,N_18542);
and U21464 (N_21464,N_18810,N_19283);
nor U21465 (N_21465,N_19412,N_19442);
xnor U21466 (N_21466,N_19380,N_18111);
nand U21467 (N_21467,N_18793,N_19246);
or U21468 (N_21468,N_18764,N_19247);
nor U21469 (N_21469,N_18838,N_19915);
and U21470 (N_21470,N_18113,N_18301);
xnor U21471 (N_21471,N_19469,N_19383);
nor U21472 (N_21472,N_18760,N_19869);
nand U21473 (N_21473,N_19131,N_19183);
and U21474 (N_21474,N_19207,N_18193);
nor U21475 (N_21475,N_18393,N_19267);
or U21476 (N_21476,N_19077,N_19794);
xor U21477 (N_21477,N_19988,N_19828);
nand U21478 (N_21478,N_19342,N_19377);
or U21479 (N_21479,N_19482,N_18642);
and U21480 (N_21480,N_19485,N_18536);
xnor U21481 (N_21481,N_19189,N_19385);
nor U21482 (N_21482,N_18428,N_18969);
nor U21483 (N_21483,N_19913,N_19280);
nor U21484 (N_21484,N_18267,N_18456);
xnor U21485 (N_21485,N_19305,N_18518);
nand U21486 (N_21486,N_18629,N_19326);
or U21487 (N_21487,N_18154,N_19810);
xnor U21488 (N_21488,N_18048,N_18406);
xor U21489 (N_21489,N_18179,N_18889);
or U21490 (N_21490,N_19218,N_18924);
or U21491 (N_21491,N_18739,N_18257);
or U21492 (N_21492,N_19109,N_19243);
xnor U21493 (N_21493,N_18386,N_18415);
or U21494 (N_21494,N_18708,N_18110);
or U21495 (N_21495,N_19681,N_19182);
or U21496 (N_21496,N_19079,N_19497);
xor U21497 (N_21497,N_19081,N_18558);
and U21498 (N_21498,N_19158,N_19274);
nand U21499 (N_21499,N_19845,N_19219);
nand U21500 (N_21500,N_19249,N_18973);
xnor U21501 (N_21501,N_19800,N_18801);
xnor U21502 (N_21502,N_19257,N_19645);
or U21503 (N_21503,N_19338,N_18012);
or U21504 (N_21504,N_19278,N_19964);
and U21505 (N_21505,N_18500,N_18839);
xor U21506 (N_21506,N_18430,N_19213);
nor U21507 (N_21507,N_19449,N_19740);
xor U21508 (N_21508,N_18191,N_19990);
nand U21509 (N_21509,N_19881,N_18704);
xor U21510 (N_21510,N_18368,N_19656);
or U21511 (N_21511,N_19902,N_19777);
or U21512 (N_21512,N_19155,N_18263);
xor U21513 (N_21513,N_18208,N_18372);
nand U21514 (N_21514,N_18500,N_18178);
and U21515 (N_21515,N_18048,N_18199);
nand U21516 (N_21516,N_18434,N_19823);
or U21517 (N_21517,N_19478,N_19139);
nor U21518 (N_21518,N_18177,N_18692);
xor U21519 (N_21519,N_19768,N_18973);
nand U21520 (N_21520,N_19032,N_18997);
nand U21521 (N_21521,N_19750,N_19229);
nor U21522 (N_21522,N_19214,N_19911);
or U21523 (N_21523,N_18983,N_18149);
nand U21524 (N_21524,N_19189,N_18436);
xor U21525 (N_21525,N_18061,N_18161);
and U21526 (N_21526,N_18593,N_18636);
and U21527 (N_21527,N_18846,N_18669);
nand U21528 (N_21528,N_19130,N_19113);
xnor U21529 (N_21529,N_19390,N_18139);
nor U21530 (N_21530,N_18698,N_18258);
or U21531 (N_21531,N_18119,N_19426);
or U21532 (N_21532,N_19817,N_19109);
nand U21533 (N_21533,N_19270,N_19631);
nor U21534 (N_21534,N_19952,N_18641);
nor U21535 (N_21535,N_19879,N_18489);
nor U21536 (N_21536,N_19844,N_19201);
xnor U21537 (N_21537,N_18074,N_18272);
xor U21538 (N_21538,N_19412,N_18440);
and U21539 (N_21539,N_18745,N_19467);
and U21540 (N_21540,N_19172,N_18366);
and U21541 (N_21541,N_18442,N_18062);
nand U21542 (N_21542,N_18416,N_18661);
and U21543 (N_21543,N_18340,N_18434);
nand U21544 (N_21544,N_18114,N_18816);
xnor U21545 (N_21545,N_18168,N_19435);
nand U21546 (N_21546,N_19290,N_18648);
xor U21547 (N_21547,N_19039,N_18239);
nand U21548 (N_21548,N_18026,N_18469);
nor U21549 (N_21549,N_19547,N_19342);
xnor U21550 (N_21550,N_18685,N_19960);
or U21551 (N_21551,N_18898,N_18543);
or U21552 (N_21552,N_19792,N_19825);
xnor U21553 (N_21553,N_19833,N_19267);
or U21554 (N_21554,N_18184,N_19128);
xor U21555 (N_21555,N_18921,N_18092);
nand U21556 (N_21556,N_18794,N_19752);
and U21557 (N_21557,N_18420,N_18958);
nand U21558 (N_21558,N_18013,N_19577);
or U21559 (N_21559,N_18441,N_19106);
xnor U21560 (N_21560,N_19170,N_19384);
and U21561 (N_21561,N_18949,N_19251);
and U21562 (N_21562,N_18314,N_19178);
or U21563 (N_21563,N_18962,N_19513);
xor U21564 (N_21564,N_19752,N_18237);
and U21565 (N_21565,N_19968,N_19768);
or U21566 (N_21566,N_18923,N_18247);
xnor U21567 (N_21567,N_18415,N_19050);
xor U21568 (N_21568,N_18954,N_19262);
and U21569 (N_21569,N_18426,N_18008);
nor U21570 (N_21570,N_19767,N_18347);
nor U21571 (N_21571,N_19512,N_18360);
nor U21572 (N_21572,N_19591,N_18302);
xor U21573 (N_21573,N_18503,N_19513);
xor U21574 (N_21574,N_18152,N_18452);
nor U21575 (N_21575,N_18543,N_19506);
nor U21576 (N_21576,N_18505,N_19676);
nand U21577 (N_21577,N_18984,N_18219);
nand U21578 (N_21578,N_18004,N_18692);
nor U21579 (N_21579,N_18988,N_19126);
and U21580 (N_21580,N_19805,N_19353);
xor U21581 (N_21581,N_18883,N_18254);
nor U21582 (N_21582,N_18484,N_18281);
or U21583 (N_21583,N_18151,N_19818);
nor U21584 (N_21584,N_18043,N_18516);
xor U21585 (N_21585,N_19006,N_18497);
nor U21586 (N_21586,N_19630,N_19249);
nand U21587 (N_21587,N_18517,N_19139);
and U21588 (N_21588,N_19066,N_19412);
nor U21589 (N_21589,N_19842,N_18850);
nor U21590 (N_21590,N_18386,N_19354);
or U21591 (N_21591,N_18875,N_19822);
xnor U21592 (N_21592,N_19425,N_18863);
xor U21593 (N_21593,N_18703,N_18446);
or U21594 (N_21594,N_19684,N_18340);
or U21595 (N_21595,N_18321,N_18875);
nand U21596 (N_21596,N_18155,N_18053);
nor U21597 (N_21597,N_18793,N_19960);
or U21598 (N_21598,N_18437,N_19100);
or U21599 (N_21599,N_19991,N_19256);
nand U21600 (N_21600,N_19420,N_19403);
nor U21601 (N_21601,N_18913,N_18865);
or U21602 (N_21602,N_19405,N_18071);
nand U21603 (N_21603,N_19159,N_18205);
or U21604 (N_21604,N_18834,N_19908);
or U21605 (N_21605,N_19027,N_19467);
nor U21606 (N_21606,N_19891,N_18355);
or U21607 (N_21607,N_18314,N_19752);
nand U21608 (N_21608,N_18261,N_18722);
or U21609 (N_21609,N_19870,N_19519);
xnor U21610 (N_21610,N_18821,N_19939);
nor U21611 (N_21611,N_18192,N_18401);
nand U21612 (N_21612,N_18628,N_18789);
or U21613 (N_21613,N_18362,N_19280);
or U21614 (N_21614,N_18853,N_18232);
and U21615 (N_21615,N_19136,N_18147);
nor U21616 (N_21616,N_19340,N_18242);
nand U21617 (N_21617,N_19862,N_19859);
nand U21618 (N_21618,N_19979,N_18179);
nor U21619 (N_21619,N_18783,N_19574);
and U21620 (N_21620,N_18325,N_18012);
nand U21621 (N_21621,N_18837,N_18962);
and U21622 (N_21622,N_18088,N_19344);
nor U21623 (N_21623,N_19855,N_19020);
and U21624 (N_21624,N_19717,N_19810);
or U21625 (N_21625,N_19813,N_18646);
or U21626 (N_21626,N_19798,N_19824);
and U21627 (N_21627,N_19517,N_18375);
nand U21628 (N_21628,N_18010,N_19646);
or U21629 (N_21629,N_19838,N_19655);
and U21630 (N_21630,N_18143,N_18633);
or U21631 (N_21631,N_18652,N_19489);
nor U21632 (N_21632,N_18302,N_18167);
nor U21633 (N_21633,N_19117,N_18517);
and U21634 (N_21634,N_18097,N_18089);
and U21635 (N_21635,N_18430,N_19272);
nor U21636 (N_21636,N_19232,N_18646);
or U21637 (N_21637,N_19714,N_19398);
or U21638 (N_21638,N_18107,N_18014);
and U21639 (N_21639,N_19505,N_18846);
xor U21640 (N_21640,N_19749,N_19746);
nand U21641 (N_21641,N_19565,N_18528);
nor U21642 (N_21642,N_18601,N_19220);
nor U21643 (N_21643,N_18335,N_18308);
xnor U21644 (N_21644,N_18021,N_18257);
and U21645 (N_21645,N_18631,N_18714);
or U21646 (N_21646,N_19549,N_19278);
nor U21647 (N_21647,N_18503,N_18144);
and U21648 (N_21648,N_18106,N_18679);
nor U21649 (N_21649,N_18002,N_18676);
xor U21650 (N_21650,N_18142,N_19037);
xnor U21651 (N_21651,N_18187,N_19128);
and U21652 (N_21652,N_19105,N_18672);
and U21653 (N_21653,N_18177,N_18089);
xor U21654 (N_21654,N_19599,N_19082);
and U21655 (N_21655,N_18159,N_19197);
xor U21656 (N_21656,N_18423,N_19683);
and U21657 (N_21657,N_19248,N_18477);
nor U21658 (N_21658,N_18453,N_18068);
nand U21659 (N_21659,N_19501,N_18300);
nor U21660 (N_21660,N_18090,N_18650);
xnor U21661 (N_21661,N_18641,N_19868);
or U21662 (N_21662,N_19922,N_18398);
or U21663 (N_21663,N_19787,N_18718);
or U21664 (N_21664,N_18829,N_19709);
nand U21665 (N_21665,N_18254,N_19859);
and U21666 (N_21666,N_19526,N_18621);
nor U21667 (N_21667,N_19439,N_19090);
nand U21668 (N_21668,N_19396,N_19302);
nor U21669 (N_21669,N_19819,N_19661);
or U21670 (N_21670,N_19565,N_19879);
and U21671 (N_21671,N_19060,N_19934);
and U21672 (N_21672,N_18675,N_18146);
nor U21673 (N_21673,N_18222,N_19200);
xnor U21674 (N_21674,N_18793,N_18882);
or U21675 (N_21675,N_18631,N_18842);
or U21676 (N_21676,N_19055,N_19715);
and U21677 (N_21677,N_19645,N_18517);
or U21678 (N_21678,N_18263,N_19728);
xnor U21679 (N_21679,N_19901,N_19641);
xor U21680 (N_21680,N_19136,N_19926);
xor U21681 (N_21681,N_18284,N_18748);
nor U21682 (N_21682,N_19303,N_19613);
nand U21683 (N_21683,N_18675,N_19526);
and U21684 (N_21684,N_18388,N_19624);
xor U21685 (N_21685,N_18773,N_18287);
nor U21686 (N_21686,N_19538,N_19750);
xnor U21687 (N_21687,N_19181,N_18554);
and U21688 (N_21688,N_18713,N_18745);
nor U21689 (N_21689,N_19324,N_18954);
or U21690 (N_21690,N_19825,N_18303);
or U21691 (N_21691,N_19498,N_18911);
nor U21692 (N_21692,N_19625,N_19599);
and U21693 (N_21693,N_19096,N_18895);
nand U21694 (N_21694,N_19133,N_18291);
nand U21695 (N_21695,N_18764,N_18314);
xnor U21696 (N_21696,N_19046,N_19066);
nand U21697 (N_21697,N_19773,N_19461);
xor U21698 (N_21698,N_19812,N_18675);
xnor U21699 (N_21699,N_18917,N_18707);
nor U21700 (N_21700,N_18236,N_19220);
xnor U21701 (N_21701,N_19770,N_18977);
or U21702 (N_21702,N_19367,N_18925);
nand U21703 (N_21703,N_19099,N_19151);
nor U21704 (N_21704,N_19850,N_18699);
nand U21705 (N_21705,N_18365,N_19647);
nand U21706 (N_21706,N_18523,N_19443);
or U21707 (N_21707,N_18217,N_18928);
xnor U21708 (N_21708,N_19131,N_19251);
and U21709 (N_21709,N_19350,N_19463);
and U21710 (N_21710,N_19204,N_19659);
nand U21711 (N_21711,N_19913,N_19646);
nor U21712 (N_21712,N_19573,N_18009);
xnor U21713 (N_21713,N_19509,N_18524);
nor U21714 (N_21714,N_18161,N_18579);
or U21715 (N_21715,N_19514,N_18062);
or U21716 (N_21716,N_18188,N_19537);
xor U21717 (N_21717,N_19399,N_18910);
nand U21718 (N_21718,N_18615,N_18920);
or U21719 (N_21719,N_19116,N_18458);
nand U21720 (N_21720,N_18594,N_19867);
nand U21721 (N_21721,N_18866,N_18905);
xnor U21722 (N_21722,N_18920,N_18422);
or U21723 (N_21723,N_19105,N_19642);
and U21724 (N_21724,N_19621,N_19628);
and U21725 (N_21725,N_18433,N_18256);
xnor U21726 (N_21726,N_19629,N_19662);
nor U21727 (N_21727,N_19682,N_18380);
xor U21728 (N_21728,N_19672,N_18190);
and U21729 (N_21729,N_19587,N_18374);
nand U21730 (N_21730,N_18212,N_18004);
and U21731 (N_21731,N_18068,N_19344);
and U21732 (N_21732,N_19777,N_19658);
nand U21733 (N_21733,N_18342,N_18815);
xnor U21734 (N_21734,N_18684,N_19341);
xnor U21735 (N_21735,N_18271,N_18209);
and U21736 (N_21736,N_18310,N_18832);
nand U21737 (N_21737,N_18301,N_18139);
nor U21738 (N_21738,N_18907,N_19007);
xor U21739 (N_21739,N_19498,N_18759);
nand U21740 (N_21740,N_18528,N_18998);
or U21741 (N_21741,N_18110,N_19292);
xor U21742 (N_21742,N_19591,N_18969);
or U21743 (N_21743,N_18665,N_18580);
nand U21744 (N_21744,N_19045,N_18989);
and U21745 (N_21745,N_19492,N_19630);
and U21746 (N_21746,N_19133,N_19175);
nand U21747 (N_21747,N_18905,N_18793);
xnor U21748 (N_21748,N_18802,N_18582);
or U21749 (N_21749,N_19020,N_18963);
nor U21750 (N_21750,N_18586,N_19497);
nor U21751 (N_21751,N_19279,N_19401);
xnor U21752 (N_21752,N_18317,N_18947);
or U21753 (N_21753,N_19156,N_18299);
or U21754 (N_21754,N_18403,N_19398);
or U21755 (N_21755,N_18573,N_19301);
nor U21756 (N_21756,N_19815,N_19663);
xor U21757 (N_21757,N_19201,N_18568);
nor U21758 (N_21758,N_18709,N_19711);
xnor U21759 (N_21759,N_19430,N_18787);
nand U21760 (N_21760,N_18764,N_19806);
nand U21761 (N_21761,N_18684,N_19307);
nor U21762 (N_21762,N_19723,N_18584);
nand U21763 (N_21763,N_19614,N_18318);
xor U21764 (N_21764,N_18173,N_19700);
nor U21765 (N_21765,N_19581,N_18089);
nand U21766 (N_21766,N_18536,N_18432);
xnor U21767 (N_21767,N_19358,N_18438);
or U21768 (N_21768,N_18244,N_18463);
nor U21769 (N_21769,N_18595,N_18969);
and U21770 (N_21770,N_18030,N_18436);
and U21771 (N_21771,N_19421,N_19022);
or U21772 (N_21772,N_18361,N_18414);
xor U21773 (N_21773,N_19334,N_19475);
nor U21774 (N_21774,N_18465,N_19172);
or U21775 (N_21775,N_19358,N_18450);
nand U21776 (N_21776,N_18211,N_18472);
and U21777 (N_21777,N_18767,N_18066);
nor U21778 (N_21778,N_18218,N_19893);
nor U21779 (N_21779,N_19539,N_18790);
nor U21780 (N_21780,N_18785,N_18546);
xor U21781 (N_21781,N_18931,N_19573);
xnor U21782 (N_21782,N_19208,N_18506);
or U21783 (N_21783,N_18813,N_18299);
nor U21784 (N_21784,N_18541,N_19694);
nor U21785 (N_21785,N_18315,N_19648);
and U21786 (N_21786,N_18651,N_19467);
and U21787 (N_21787,N_18349,N_18873);
or U21788 (N_21788,N_18547,N_19134);
xnor U21789 (N_21789,N_18035,N_19770);
and U21790 (N_21790,N_19006,N_19290);
xnor U21791 (N_21791,N_19268,N_18726);
nor U21792 (N_21792,N_18361,N_18755);
or U21793 (N_21793,N_18999,N_18491);
or U21794 (N_21794,N_19049,N_19188);
nor U21795 (N_21795,N_18289,N_18123);
nand U21796 (N_21796,N_19189,N_18310);
or U21797 (N_21797,N_18381,N_19571);
and U21798 (N_21798,N_19671,N_18809);
or U21799 (N_21799,N_19988,N_18156);
xor U21800 (N_21800,N_18243,N_19624);
or U21801 (N_21801,N_19019,N_18923);
nand U21802 (N_21802,N_19848,N_18423);
nand U21803 (N_21803,N_18052,N_18711);
or U21804 (N_21804,N_19541,N_19936);
nand U21805 (N_21805,N_19431,N_19881);
and U21806 (N_21806,N_19633,N_18234);
and U21807 (N_21807,N_19888,N_18232);
xor U21808 (N_21808,N_18242,N_19146);
and U21809 (N_21809,N_19297,N_19309);
nor U21810 (N_21810,N_18696,N_19655);
or U21811 (N_21811,N_18779,N_18418);
or U21812 (N_21812,N_19704,N_19590);
nand U21813 (N_21813,N_19874,N_19219);
nor U21814 (N_21814,N_18236,N_18701);
and U21815 (N_21815,N_19241,N_19376);
xnor U21816 (N_21816,N_19545,N_18964);
nor U21817 (N_21817,N_18712,N_19209);
nand U21818 (N_21818,N_18184,N_19470);
nor U21819 (N_21819,N_19277,N_19710);
nand U21820 (N_21820,N_19567,N_18258);
nor U21821 (N_21821,N_19713,N_18517);
xor U21822 (N_21822,N_19699,N_18081);
or U21823 (N_21823,N_19311,N_19774);
or U21824 (N_21824,N_18584,N_18285);
and U21825 (N_21825,N_19882,N_19238);
and U21826 (N_21826,N_19389,N_19122);
and U21827 (N_21827,N_18490,N_18548);
nand U21828 (N_21828,N_19459,N_18712);
or U21829 (N_21829,N_18271,N_19515);
or U21830 (N_21830,N_18917,N_19392);
and U21831 (N_21831,N_18466,N_19803);
nand U21832 (N_21832,N_19775,N_18556);
and U21833 (N_21833,N_18687,N_19638);
xnor U21834 (N_21834,N_19639,N_19079);
nor U21835 (N_21835,N_18215,N_19820);
nor U21836 (N_21836,N_18562,N_19123);
and U21837 (N_21837,N_18139,N_18496);
and U21838 (N_21838,N_19069,N_18483);
nand U21839 (N_21839,N_18277,N_18473);
xor U21840 (N_21840,N_18966,N_19946);
and U21841 (N_21841,N_18319,N_19415);
nand U21842 (N_21842,N_18419,N_19597);
and U21843 (N_21843,N_19461,N_19348);
xor U21844 (N_21844,N_19613,N_18757);
nand U21845 (N_21845,N_18599,N_18559);
or U21846 (N_21846,N_19494,N_19572);
nor U21847 (N_21847,N_18197,N_18141);
nor U21848 (N_21848,N_19860,N_19905);
or U21849 (N_21849,N_18276,N_19434);
and U21850 (N_21850,N_19389,N_18435);
or U21851 (N_21851,N_18273,N_19722);
nand U21852 (N_21852,N_19101,N_18342);
xor U21853 (N_21853,N_19355,N_18564);
nor U21854 (N_21854,N_19311,N_18841);
nand U21855 (N_21855,N_18593,N_18809);
nand U21856 (N_21856,N_19409,N_19089);
xor U21857 (N_21857,N_19192,N_18087);
and U21858 (N_21858,N_19139,N_19111);
nor U21859 (N_21859,N_18390,N_18516);
xor U21860 (N_21860,N_19690,N_18268);
and U21861 (N_21861,N_19676,N_18163);
or U21862 (N_21862,N_18877,N_19333);
or U21863 (N_21863,N_19566,N_18573);
xor U21864 (N_21864,N_19127,N_19970);
nand U21865 (N_21865,N_19243,N_18514);
and U21866 (N_21866,N_19667,N_18484);
or U21867 (N_21867,N_19281,N_19886);
or U21868 (N_21868,N_18193,N_19674);
and U21869 (N_21869,N_18541,N_18119);
xor U21870 (N_21870,N_18603,N_18956);
nor U21871 (N_21871,N_19741,N_18665);
and U21872 (N_21872,N_19060,N_18464);
or U21873 (N_21873,N_18488,N_18892);
xnor U21874 (N_21874,N_19333,N_19737);
xnor U21875 (N_21875,N_19207,N_18590);
nor U21876 (N_21876,N_19232,N_18491);
xor U21877 (N_21877,N_18542,N_19786);
or U21878 (N_21878,N_18992,N_19327);
xnor U21879 (N_21879,N_18224,N_18597);
xnor U21880 (N_21880,N_19673,N_18218);
or U21881 (N_21881,N_19189,N_18811);
nand U21882 (N_21882,N_19253,N_19476);
nor U21883 (N_21883,N_18518,N_18394);
and U21884 (N_21884,N_18520,N_18084);
nand U21885 (N_21885,N_18393,N_18113);
nor U21886 (N_21886,N_19639,N_18548);
and U21887 (N_21887,N_19186,N_19842);
or U21888 (N_21888,N_19826,N_19066);
and U21889 (N_21889,N_19191,N_19379);
nor U21890 (N_21890,N_18763,N_19897);
nand U21891 (N_21891,N_19720,N_18689);
and U21892 (N_21892,N_18331,N_18437);
and U21893 (N_21893,N_19777,N_18503);
nand U21894 (N_21894,N_19159,N_19763);
nand U21895 (N_21895,N_18217,N_18391);
nor U21896 (N_21896,N_19630,N_19774);
and U21897 (N_21897,N_18273,N_19616);
xor U21898 (N_21898,N_18870,N_19998);
xor U21899 (N_21899,N_19886,N_19312);
or U21900 (N_21900,N_19636,N_19732);
nand U21901 (N_21901,N_18235,N_19245);
nor U21902 (N_21902,N_19369,N_18164);
and U21903 (N_21903,N_18219,N_18538);
or U21904 (N_21904,N_18644,N_18442);
nor U21905 (N_21905,N_19365,N_18549);
nor U21906 (N_21906,N_19775,N_19027);
xor U21907 (N_21907,N_19155,N_18389);
xor U21908 (N_21908,N_19954,N_19983);
and U21909 (N_21909,N_19801,N_18821);
or U21910 (N_21910,N_19253,N_19776);
nand U21911 (N_21911,N_18531,N_19036);
xnor U21912 (N_21912,N_18173,N_18146);
nor U21913 (N_21913,N_18515,N_19230);
or U21914 (N_21914,N_18859,N_19721);
xnor U21915 (N_21915,N_18891,N_18971);
or U21916 (N_21916,N_19840,N_18228);
and U21917 (N_21917,N_19110,N_19768);
or U21918 (N_21918,N_18726,N_19753);
or U21919 (N_21919,N_18859,N_19512);
or U21920 (N_21920,N_18193,N_18593);
or U21921 (N_21921,N_18630,N_19141);
xor U21922 (N_21922,N_19342,N_19518);
and U21923 (N_21923,N_19558,N_18504);
xor U21924 (N_21924,N_18645,N_19775);
xnor U21925 (N_21925,N_19755,N_18856);
or U21926 (N_21926,N_18333,N_19118);
or U21927 (N_21927,N_19780,N_19310);
nor U21928 (N_21928,N_19542,N_19814);
nor U21929 (N_21929,N_18538,N_19085);
xor U21930 (N_21930,N_18443,N_18948);
or U21931 (N_21931,N_18436,N_19857);
or U21932 (N_21932,N_19135,N_18492);
or U21933 (N_21933,N_18468,N_19029);
nor U21934 (N_21934,N_18698,N_18935);
and U21935 (N_21935,N_18697,N_18146);
and U21936 (N_21936,N_18820,N_18594);
nand U21937 (N_21937,N_19863,N_18376);
xnor U21938 (N_21938,N_19644,N_18996);
or U21939 (N_21939,N_19500,N_18901);
and U21940 (N_21940,N_19447,N_19897);
and U21941 (N_21941,N_18084,N_18210);
nand U21942 (N_21942,N_19390,N_19027);
and U21943 (N_21943,N_18278,N_18321);
or U21944 (N_21944,N_18251,N_19001);
or U21945 (N_21945,N_19246,N_19910);
and U21946 (N_21946,N_19212,N_19257);
and U21947 (N_21947,N_18119,N_18272);
or U21948 (N_21948,N_19016,N_19805);
xor U21949 (N_21949,N_18251,N_18688);
nand U21950 (N_21950,N_18128,N_19735);
and U21951 (N_21951,N_18607,N_18997);
nor U21952 (N_21952,N_19143,N_18931);
nand U21953 (N_21953,N_18707,N_18222);
or U21954 (N_21954,N_19032,N_19784);
and U21955 (N_21955,N_18358,N_18692);
xor U21956 (N_21956,N_19675,N_18548);
and U21957 (N_21957,N_19265,N_18329);
xor U21958 (N_21958,N_18506,N_19734);
nand U21959 (N_21959,N_19733,N_18576);
nand U21960 (N_21960,N_18745,N_19275);
nand U21961 (N_21961,N_18216,N_19492);
nor U21962 (N_21962,N_19550,N_19768);
or U21963 (N_21963,N_18347,N_18564);
nor U21964 (N_21964,N_18587,N_18829);
xnor U21965 (N_21965,N_18246,N_19766);
nand U21966 (N_21966,N_18882,N_19745);
nand U21967 (N_21967,N_18930,N_19698);
nor U21968 (N_21968,N_19166,N_19125);
and U21969 (N_21969,N_19639,N_19065);
xor U21970 (N_21970,N_18350,N_18551);
or U21971 (N_21971,N_18751,N_18328);
and U21972 (N_21972,N_18140,N_18816);
xor U21973 (N_21973,N_19738,N_18740);
or U21974 (N_21974,N_18708,N_18054);
and U21975 (N_21975,N_19767,N_19336);
or U21976 (N_21976,N_19224,N_19726);
xor U21977 (N_21977,N_18470,N_19180);
and U21978 (N_21978,N_18683,N_19771);
xnor U21979 (N_21979,N_18415,N_19805);
and U21980 (N_21980,N_18640,N_19631);
xnor U21981 (N_21981,N_18039,N_19343);
nor U21982 (N_21982,N_18379,N_18979);
or U21983 (N_21983,N_19572,N_18996);
and U21984 (N_21984,N_18977,N_19922);
and U21985 (N_21985,N_18749,N_18944);
or U21986 (N_21986,N_19404,N_18835);
and U21987 (N_21987,N_18648,N_19003);
and U21988 (N_21988,N_18020,N_19816);
nor U21989 (N_21989,N_18792,N_19496);
and U21990 (N_21990,N_19101,N_19124);
nor U21991 (N_21991,N_18043,N_18016);
and U21992 (N_21992,N_19023,N_18167);
xnor U21993 (N_21993,N_19473,N_18888);
and U21994 (N_21994,N_19755,N_18823);
and U21995 (N_21995,N_19763,N_18499);
nand U21996 (N_21996,N_19148,N_18194);
nor U21997 (N_21997,N_19518,N_18296);
or U21998 (N_21998,N_19617,N_18629);
nand U21999 (N_21999,N_19898,N_19792);
nor U22000 (N_22000,N_20156,N_20003);
nor U22001 (N_22001,N_21945,N_21674);
and U22002 (N_22002,N_21242,N_21308);
or U22003 (N_22003,N_20699,N_21552);
or U22004 (N_22004,N_21558,N_20237);
or U22005 (N_22005,N_21883,N_20157);
and U22006 (N_22006,N_21388,N_21973);
nand U22007 (N_22007,N_20682,N_21857);
xnor U22008 (N_22008,N_20327,N_20059);
or U22009 (N_22009,N_20804,N_20436);
nand U22010 (N_22010,N_21757,N_20358);
nand U22011 (N_22011,N_21174,N_20026);
nor U22012 (N_22012,N_21090,N_20692);
nand U22013 (N_22013,N_21790,N_20365);
nor U22014 (N_22014,N_21358,N_20143);
xor U22015 (N_22015,N_20398,N_21393);
xor U22016 (N_22016,N_21766,N_21208);
and U22017 (N_22017,N_21931,N_20546);
xor U22018 (N_22018,N_20153,N_21296);
and U22019 (N_22019,N_21075,N_21853);
and U22020 (N_22020,N_21877,N_20636);
nor U22021 (N_22021,N_21613,N_20789);
or U22022 (N_22022,N_20185,N_21259);
nand U22023 (N_22023,N_20161,N_21038);
xor U22024 (N_22024,N_20674,N_20407);
xnor U22025 (N_22025,N_20272,N_21708);
nor U22026 (N_22026,N_21738,N_20426);
xor U22027 (N_22027,N_21053,N_21061);
nand U22028 (N_22028,N_21521,N_21999);
and U22029 (N_22029,N_21850,N_20085);
xor U22030 (N_22030,N_21445,N_20454);
and U22031 (N_22031,N_21142,N_21278);
and U22032 (N_22032,N_21171,N_21050);
or U22033 (N_22033,N_20459,N_20802);
nor U22034 (N_22034,N_21466,N_21702);
nor U22035 (N_22035,N_21018,N_20395);
and U22036 (N_22036,N_20173,N_21123);
or U22037 (N_22037,N_20368,N_21873);
xnor U22038 (N_22038,N_20463,N_21730);
or U22039 (N_22039,N_21482,N_20400);
nor U22040 (N_22040,N_21305,N_20431);
xnor U22041 (N_22041,N_20736,N_21763);
and U22042 (N_22042,N_21728,N_21668);
xnor U22043 (N_22043,N_20066,N_21011);
and U22044 (N_22044,N_21603,N_20107);
xnor U22045 (N_22045,N_20844,N_20671);
nor U22046 (N_22046,N_21656,N_21488);
nand U22047 (N_22047,N_21524,N_20110);
xor U22048 (N_22048,N_21864,N_20855);
or U22049 (N_22049,N_21186,N_21337);
xor U22050 (N_22050,N_20825,N_21933);
or U22051 (N_22051,N_21303,N_20527);
nand U22052 (N_22052,N_21349,N_20791);
nor U22053 (N_22053,N_20016,N_21441);
nor U22054 (N_22054,N_21426,N_20680);
nor U22055 (N_22055,N_21593,N_20442);
nand U22056 (N_22056,N_21254,N_21910);
nor U22057 (N_22057,N_20679,N_21246);
nor U22058 (N_22058,N_20572,N_20010);
nand U22059 (N_22059,N_20921,N_20158);
xor U22060 (N_22060,N_21887,N_20332);
xnor U22061 (N_22061,N_21882,N_20561);
nand U22062 (N_22062,N_21116,N_21487);
xor U22063 (N_22063,N_21102,N_21602);
or U22064 (N_22064,N_21250,N_20299);
and U22065 (N_22065,N_21084,N_21163);
xnor U22066 (N_22066,N_20351,N_21806);
nor U22067 (N_22067,N_20824,N_20735);
nand U22068 (N_22068,N_20579,N_21884);
xnor U22069 (N_22069,N_20468,N_21583);
and U22070 (N_22070,N_21671,N_20520);
nand U22071 (N_22071,N_21016,N_20606);
nand U22072 (N_22072,N_20275,N_21943);
xor U22073 (N_22073,N_21282,N_20260);
nand U22074 (N_22074,N_20754,N_21865);
nand U22075 (N_22075,N_20257,N_21506);
nand U22076 (N_22076,N_20709,N_20451);
xor U22077 (N_22077,N_21988,N_20730);
or U22078 (N_22078,N_20329,N_20382);
xor U22079 (N_22079,N_21907,N_21258);
nor U22080 (N_22080,N_20044,N_20467);
nor U22081 (N_22081,N_21664,N_20386);
nand U22082 (N_22082,N_21356,N_21399);
xor U22083 (N_22083,N_21146,N_21332);
and U22084 (N_22084,N_21585,N_21136);
and U22085 (N_22085,N_21972,N_21576);
xor U22086 (N_22086,N_20650,N_21727);
nor U22087 (N_22087,N_21161,N_20174);
or U22088 (N_22088,N_21484,N_21214);
nor U22089 (N_22089,N_21295,N_21808);
nand U22090 (N_22090,N_21469,N_21577);
nand U22091 (N_22091,N_21098,N_20806);
nand U22092 (N_22092,N_21540,N_21454);
xnor U22093 (N_22093,N_21798,N_21395);
xor U22094 (N_22094,N_21192,N_20387);
nand U22095 (N_22095,N_20183,N_20485);
nand U22096 (N_22096,N_21625,N_20539);
and U22097 (N_22097,N_20502,N_21516);
and U22098 (N_22098,N_20195,N_21162);
xor U22099 (N_22099,N_21754,N_21858);
nor U22100 (N_22100,N_20793,N_20437);
xnor U22101 (N_22101,N_20392,N_21252);
nor U22102 (N_22102,N_21211,N_21485);
xor U22103 (N_22103,N_21587,N_21543);
nor U22104 (N_22104,N_20181,N_20489);
xor U22105 (N_22105,N_21304,N_21379);
xor U22106 (N_22106,N_21334,N_21039);
or U22107 (N_22107,N_21059,N_20859);
nand U22108 (N_22108,N_21057,N_20111);
and U22109 (N_22109,N_21078,N_20402);
nor U22110 (N_22110,N_20975,N_21222);
or U22111 (N_22111,N_21753,N_20960);
nor U22112 (N_22112,N_20141,N_20390);
nand U22113 (N_22113,N_21658,N_21081);
or U22114 (N_22114,N_20642,N_20277);
nand U22115 (N_22115,N_20620,N_20089);
xor U22116 (N_22116,N_21971,N_21660);
xnor U22117 (N_22117,N_21031,N_21932);
nand U22118 (N_22118,N_20987,N_20867);
or U22119 (N_22119,N_20509,N_21443);
and U22120 (N_22120,N_20039,N_21079);
nor U22121 (N_22121,N_21329,N_20959);
nor U22122 (N_22122,N_21709,N_21848);
nand U22123 (N_22123,N_20775,N_21501);
nand U22124 (N_22124,N_21912,N_20949);
and U22125 (N_22125,N_21239,N_20799);
or U22126 (N_22126,N_21604,N_21825);
nor U22127 (N_22127,N_20635,N_21111);
or U22128 (N_22128,N_20826,N_21650);
nor U22129 (N_22129,N_21828,N_20250);
xnor U22130 (N_22130,N_20380,N_20823);
or U22131 (N_22131,N_20067,N_20136);
or U22132 (N_22132,N_21970,N_21006);
nand U22133 (N_22133,N_21721,N_20862);
xnor U22134 (N_22134,N_21427,N_20225);
xnor U22135 (N_22135,N_20715,N_20388);
xnor U22136 (N_22136,N_21251,N_20100);
nor U22137 (N_22137,N_20711,N_21983);
nor U22138 (N_22138,N_20201,N_21527);
nor U22139 (N_22139,N_21740,N_21977);
or U22140 (N_22140,N_20683,N_21622);
or U22141 (N_22141,N_21396,N_21037);
nand U22142 (N_22142,N_21535,N_21009);
nor U22143 (N_22143,N_21835,N_21237);
or U22144 (N_22144,N_21467,N_21082);
xnor U22145 (N_22145,N_20062,N_21867);
and U22146 (N_22146,N_21475,N_21385);
nand U22147 (N_22147,N_21590,N_21107);
xnor U22148 (N_22148,N_21348,N_20223);
nor U22149 (N_22149,N_20588,N_21989);
nand U22150 (N_22150,N_21741,N_21698);
nor U22151 (N_22151,N_20849,N_20995);
nor U22152 (N_22152,N_21408,N_21387);
nand U22153 (N_22153,N_21160,N_21816);
and U22154 (N_22154,N_20491,N_20764);
and U22155 (N_22155,N_20373,N_21263);
nand U22156 (N_22156,N_20098,N_21398);
xor U22157 (N_22157,N_20685,N_21908);
and U22158 (N_22158,N_21094,N_20877);
nand U22159 (N_22159,N_20105,N_20902);
nor U22160 (N_22160,N_21541,N_20193);
and U22161 (N_22161,N_21335,N_21126);
nor U22162 (N_22162,N_20318,N_20757);
and U22163 (N_22163,N_21209,N_21518);
xnor U22164 (N_22164,N_21834,N_21324);
nand U22165 (N_22165,N_20421,N_21369);
xnor U22166 (N_22166,N_20404,N_20099);
xnor U22167 (N_22167,N_21394,N_21444);
or U22168 (N_22168,N_21961,N_20627);
nand U22169 (N_22169,N_21364,N_20352);
nand U22170 (N_22170,N_20645,N_21270);
or U22171 (N_22171,N_20314,N_21409);
nand U22172 (N_22172,N_20551,N_20203);
or U22173 (N_22173,N_21986,N_21173);
nand U22174 (N_22174,N_20535,N_21720);
xor U22175 (N_22175,N_21878,N_21913);
nand U22176 (N_22176,N_20837,N_21810);
nor U22177 (N_22177,N_20768,N_20623);
or U22178 (N_22178,N_20629,N_21784);
or U22179 (N_22179,N_21235,N_21830);
xnor U22180 (N_22180,N_20394,N_20084);
and U22181 (N_22181,N_21472,N_21776);
and U22182 (N_22182,N_20909,N_21620);
xnor U22183 (N_22183,N_20043,N_21391);
nand U22184 (N_22184,N_21683,N_20166);
xnor U22185 (N_22185,N_21956,N_20154);
and U22186 (N_22186,N_21115,N_21134);
xor U22187 (N_22187,N_20544,N_20922);
xnor U22188 (N_22188,N_21580,N_20022);
or U22189 (N_22189,N_21119,N_20274);
and U22190 (N_22190,N_21814,N_21731);
or U22191 (N_22191,N_21184,N_20967);
and U22192 (N_22192,N_21657,N_21206);
and U22193 (N_22193,N_20749,N_20704);
xnor U22194 (N_22194,N_20870,N_20585);
or U22195 (N_22195,N_20772,N_20052);
xor U22196 (N_22196,N_20427,N_20236);
xnor U22197 (N_22197,N_20461,N_20769);
and U22198 (N_22198,N_21791,N_20821);
xor U22199 (N_22199,N_20777,N_21240);
nand U22200 (N_22200,N_20140,N_20372);
and U22201 (N_22201,N_21568,N_21693);
xor U22202 (N_22202,N_21299,N_20742);
xnor U22203 (N_22203,N_21440,N_21419);
xor U22204 (N_22204,N_20654,N_20978);
xor U22205 (N_22205,N_20233,N_20340);
xor U22206 (N_22206,N_21339,N_20335);
nand U22207 (N_22207,N_20522,N_20345);
xnor U22208 (N_22208,N_20077,N_21153);
nor U22209 (N_22209,N_20302,N_20384);
and U22210 (N_22210,N_21829,N_20121);
or U22211 (N_22211,N_20559,N_20560);
nand U22212 (N_22212,N_21981,N_21546);
nor U22213 (N_22213,N_20591,N_20076);
xor U22214 (N_22214,N_20162,N_21759);
or U22215 (N_22215,N_20895,N_20308);
xor U22216 (N_22216,N_20653,N_20350);
or U22217 (N_22217,N_21191,N_21694);
nand U22218 (N_22218,N_20150,N_21000);
nor U22219 (N_22219,N_20168,N_20907);
and U22220 (N_22220,N_21906,N_21143);
xor U22221 (N_22221,N_21779,N_21096);
nand U22222 (N_22222,N_21975,N_20297);
or U22223 (N_22223,N_20095,N_20752);
or U22224 (N_22224,N_20771,N_21493);
or U22225 (N_22225,N_20048,N_20575);
or U22226 (N_22226,N_20523,N_21570);
xnor U22227 (N_22227,N_21056,N_20836);
nand U22228 (N_22228,N_20720,N_21085);
and U22229 (N_22229,N_20011,N_21236);
and U22230 (N_22230,N_20230,N_21941);
nand U22231 (N_22231,N_21462,N_21370);
xnor U22232 (N_22232,N_21726,N_21782);
xor U22233 (N_22233,N_20131,N_20189);
or U22234 (N_22234,N_21780,N_20124);
nor U22235 (N_22235,N_21330,N_20547);
or U22236 (N_22236,N_21068,N_20578);
nand U22237 (N_22237,N_21225,N_20473);
and U22238 (N_22238,N_21434,N_21148);
xnor U22239 (N_22239,N_20840,N_21948);
or U22240 (N_22240,N_20795,N_20197);
and U22241 (N_22241,N_20882,N_20893);
nor U22242 (N_22242,N_20482,N_20422);
and U22243 (N_22243,N_21639,N_20073);
nor U22244 (N_22244,N_21967,N_21804);
xnor U22245 (N_22245,N_21241,N_21596);
xnor U22246 (N_22246,N_21080,N_20945);
and U22247 (N_22247,N_21903,N_21281);
xor U22248 (N_22248,N_21993,N_20601);
nor U22249 (N_22249,N_20714,N_20819);
xnor U22250 (N_22250,N_21612,N_20514);
or U22251 (N_22251,N_21478,N_21937);
nand U22252 (N_22252,N_21248,N_20060);
xor U22253 (N_22253,N_20243,N_20611);
xor U22254 (N_22254,N_21313,N_20313);
xnor U22255 (N_22255,N_20206,N_21991);
nand U22256 (N_22256,N_21083,N_20460);
and U22257 (N_22257,N_21752,N_20342);
or U22258 (N_22258,N_20758,N_20955);
nand U22259 (N_22259,N_21035,N_21003);
nor U22260 (N_22260,N_21794,N_20854);
nand U22261 (N_22261,N_21405,N_21761);
and U22262 (N_22262,N_20188,N_21522);
nand U22263 (N_22263,N_20139,N_20526);
nand U22264 (N_22264,N_21483,N_20018);
or U22265 (N_22265,N_20109,N_21023);
and U22266 (N_22266,N_21044,N_21925);
nand U22267 (N_22267,N_20869,N_21336);
and U22268 (N_22268,N_20924,N_21923);
xor U22269 (N_22269,N_20550,N_21821);
xnor U22270 (N_22270,N_20448,N_20160);
nor U22271 (N_22271,N_21697,N_20790);
and U22272 (N_22272,N_21769,N_20604);
nor U22273 (N_22273,N_20232,N_20622);
and U22274 (N_22274,N_21508,N_20739);
xor U22275 (N_22275,N_20567,N_21957);
nand U22276 (N_22276,N_20020,N_20224);
or U22277 (N_22277,N_20807,N_20965);
or U22278 (N_22278,N_21692,N_20737);
or U22279 (N_22279,N_20626,N_21382);
and U22280 (N_22280,N_20839,N_21895);
and U22281 (N_22281,N_20766,N_21617);
or U22282 (N_22282,N_21187,N_21953);
xor U22283 (N_22283,N_20226,N_20215);
or U22284 (N_22284,N_20943,N_20132);
or U22285 (N_22285,N_21344,N_20857);
xor U22286 (N_22286,N_21876,N_21285);
or U22287 (N_22287,N_21271,N_20419);
xor U22288 (N_22288,N_21450,N_20322);
nand U22289 (N_22289,N_20244,N_21954);
or U22290 (N_22290,N_21582,N_20525);
nand U22291 (N_22291,N_21047,N_20499);
nand U22292 (N_22292,N_20242,N_21188);
or U22293 (N_22293,N_20930,N_21432);
or U22294 (N_22294,N_20190,N_21700);
and U22295 (N_22295,N_20487,N_21890);
xor U22296 (N_22296,N_21520,N_20667);
nand U22297 (N_22297,N_21340,N_20847);
or U22298 (N_22298,N_20283,N_21742);
or U22299 (N_22299,N_21673,N_21392);
or U22300 (N_22300,N_20135,N_20029);
or U22301 (N_22301,N_21465,N_20383);
or U22302 (N_22302,N_21154,N_21390);
nand U22303 (N_22303,N_20898,N_21586);
and U22304 (N_22304,N_20753,N_21066);
or U22305 (N_22305,N_21510,N_20471);
nand U22306 (N_22306,N_20655,N_20581);
and U22307 (N_22307,N_21537,N_20106);
and U22308 (N_22308,N_20050,N_21049);
and U22309 (N_22309,N_21204,N_21809);
nand U22310 (N_22310,N_21891,N_21566);
and U22311 (N_22311,N_20164,N_21966);
and U22312 (N_22312,N_21223,N_20903);
nor U22313 (N_22313,N_20759,N_20198);
xor U22314 (N_22314,N_20926,N_21133);
xor U22315 (N_22315,N_21261,N_20298);
and U22316 (N_22316,N_21940,N_20021);
xor U22317 (N_22317,N_20894,N_21029);
xnor U22318 (N_22318,N_21463,N_20023);
xor U22319 (N_22319,N_21026,N_21797);
nand U22320 (N_22320,N_21114,N_20090);
xnor U22321 (N_22321,N_20458,N_20745);
xnor U22322 (N_22322,N_20008,N_21578);
xor U22323 (N_22323,N_20968,N_21178);
nand U22324 (N_22324,N_21514,N_20505);
or U22325 (N_22325,N_21077,N_20800);
nor U22326 (N_22326,N_20670,N_21213);
or U22327 (N_22327,N_21157,N_20536);
and U22328 (N_22328,N_21929,N_20783);
xor U22329 (N_22329,N_21205,N_20068);
nor U22330 (N_22330,N_20963,N_21447);
xnor U22331 (N_22331,N_21328,N_20796);
nor U22332 (N_22332,N_20493,N_21982);
nand U22333 (N_22333,N_21269,N_20541);
nor U22334 (N_22334,N_21479,N_21938);
xor U22335 (N_22335,N_21198,N_21277);
xor U22336 (N_22336,N_20177,N_21476);
nand U22337 (N_22337,N_20217,N_20456);
nand U22338 (N_22338,N_21888,N_21451);
xor U22339 (N_22339,N_20058,N_20979);
or U22340 (N_22340,N_21918,N_20644);
nor U22341 (N_22341,N_21418,N_21431);
xnor U22342 (N_22342,N_20005,N_21125);
xor U22343 (N_22343,N_21641,N_21800);
or U22344 (N_22344,N_20831,N_20580);
and U22345 (N_22345,N_21718,N_21151);
nand U22346 (N_22346,N_20480,N_20608);
nand U22347 (N_22347,N_20009,N_20891);
and U22348 (N_22348,N_20982,N_21733);
nand U22349 (N_22349,N_20897,N_20876);
and U22350 (N_22350,N_20321,N_20797);
xnor U22351 (N_22351,N_21960,N_20359);
nand U22352 (N_22352,N_21453,N_20123);
nor U22353 (N_22353,N_21342,N_20637);
nand U22354 (N_22354,N_20534,N_20142);
nand U22355 (N_22355,N_20037,N_20904);
or U22356 (N_22356,N_21074,N_21714);
xor U22357 (N_22357,N_20810,N_20208);
nand U22358 (N_22358,N_21103,N_21930);
or U22359 (N_22359,N_20348,N_21155);
and U22360 (N_22360,N_21856,N_21783);
xnor U22361 (N_22361,N_21224,N_21293);
xnor U22362 (N_22362,N_20378,N_20441);
nand U22363 (N_22363,N_20994,N_20952);
and U22364 (N_22364,N_20330,N_21219);
nor U22365 (N_22365,N_21531,N_20634);
nor U22366 (N_22366,N_20196,N_20271);
or U22367 (N_22367,N_21437,N_21542);
xnor U22368 (N_22368,N_21158,N_20721);
nor U22369 (N_22369,N_21316,N_20293);
and U22370 (N_22370,N_20070,N_21439);
xnor U22371 (N_22371,N_21500,N_21456);
xor U22372 (N_22372,N_21286,N_21351);
or U22373 (N_22373,N_20915,N_20492);
and U22374 (N_22374,N_20770,N_21924);
or U22375 (N_22375,N_21199,N_21958);
or U22376 (N_22376,N_20652,N_20477);
nand U22377 (N_22377,N_20621,N_21353);
xor U22378 (N_22378,N_21633,N_20657);
nand U22379 (N_22379,N_21807,N_20285);
nor U22380 (N_22380,N_21631,N_20780);
nand U22381 (N_22381,N_21257,N_21599);
nand U22382 (N_22382,N_21024,N_20033);
nand U22383 (N_22383,N_20125,N_20956);
and U22384 (N_22384,N_20462,N_20908);
xnor U22385 (N_22385,N_21609,N_21109);
or U22386 (N_22386,N_20532,N_20628);
nor U22387 (N_22387,N_21879,N_21365);
or U22388 (N_22388,N_20693,N_21900);
or U22389 (N_22389,N_21113,N_21283);
nand U22390 (N_22390,N_21127,N_21238);
and U22391 (N_22391,N_20087,N_21584);
xnor U22392 (N_22392,N_21574,N_21554);
nand U22393 (N_22393,N_20815,N_21400);
nand U22394 (N_22394,N_21383,N_20114);
or U22395 (N_22395,N_21167,N_20262);
or U22396 (N_22396,N_20379,N_20705);
and U22397 (N_22397,N_21985,N_21415);
nand U22398 (N_22398,N_21688,N_21628);
nor U22399 (N_22399,N_20694,N_20178);
or U22400 (N_22400,N_20740,N_20363);
nor U22401 (N_22401,N_20713,N_21289);
xnor U22402 (N_22402,N_20192,N_20906);
xnor U22403 (N_22403,N_20981,N_20747);
or U22404 (N_22404,N_20962,N_21859);
or U22405 (N_22405,N_21140,N_20868);
nor U22406 (N_22406,N_20172,N_20457);
nor U22407 (N_22407,N_20469,N_20453);
nand U22408 (N_22408,N_20937,N_20612);
or U22409 (N_22409,N_21818,N_21666);
xnor U22410 (N_22410,N_21013,N_20354);
nand U22411 (N_22411,N_21298,N_20884);
nand U22412 (N_22412,N_20942,N_21755);
nand U22413 (N_22413,N_20417,N_20498);
xnor U22414 (N_22414,N_21927,N_21823);
or U22415 (N_22415,N_21706,N_21597);
nand U22416 (N_22416,N_20179,N_20883);
xor U22417 (N_22417,N_21108,N_20167);
or U22418 (N_22418,N_21870,N_21185);
nand U22419 (N_22419,N_20725,N_21831);
nor U22420 (N_22420,N_21914,N_21359);
nand U22421 (N_22421,N_20258,N_20304);
nand U22422 (N_22422,N_21065,N_20415);
and U22423 (N_22423,N_20370,N_21667);
or U22424 (N_22424,N_21149,N_20896);
xor U22425 (N_22425,N_20091,N_20675);
xor U22426 (N_22426,N_20701,N_21840);
nor U22427 (N_22427,N_21600,N_21626);
nand U22428 (N_22428,N_20845,N_20678);
or U22429 (N_22429,N_20278,N_20557);
and U22430 (N_22430,N_20863,N_20901);
or U22431 (N_22431,N_21615,N_20432);
nor U22432 (N_22432,N_20695,N_20205);
xnor U22433 (N_22433,N_20133,N_21320);
nor U22434 (N_22434,N_20743,N_21314);
xor U22435 (N_22435,N_20887,N_21538);
and U22436 (N_22436,N_21575,N_21773);
nand U22437 (N_22437,N_20873,N_21743);
nand U22438 (N_22438,N_20101,N_21820);
nor U22439 (N_22439,N_21020,N_21486);
nor U22440 (N_22440,N_21539,N_21976);
and U22441 (N_22441,N_20801,N_20853);
nor U22442 (N_22442,N_21423,N_21051);
nor U22443 (N_22443,N_21560,N_21179);
or U22444 (N_22444,N_20054,N_20182);
and U22445 (N_22445,N_20838,N_20081);
and U22446 (N_22446,N_20497,N_21473);
xor U22447 (N_22447,N_21710,N_21815);
xnor U22448 (N_22448,N_20813,N_21963);
nor U22449 (N_22449,N_20885,N_21892);
nand U22450 (N_22450,N_21150,N_21934);
nand U22451 (N_22451,N_20306,N_21010);
nor U22452 (N_22452,N_21417,N_20986);
nor U22453 (N_22453,N_20778,N_21768);
or U22454 (N_22454,N_21354,N_20938);
and U22455 (N_22455,N_21407,N_20706);
nand U22456 (N_22456,N_20990,N_20104);
xnor U22457 (N_22457,N_20346,N_21045);
xor U22458 (N_22458,N_20276,N_21095);
xnor U22459 (N_22459,N_20216,N_21572);
xnor U22460 (N_22460,N_21772,N_21321);
and U22461 (N_22461,N_20376,N_20564);
xor U22462 (N_22462,N_20864,N_20718);
xor U22463 (N_22463,N_20587,N_20273);
nor U22464 (N_22464,N_21571,N_21406);
nor U22465 (N_22465,N_20061,N_20138);
nor U22466 (N_22466,N_20647,N_20966);
and U22467 (N_22467,N_20065,N_21646);
nand U22468 (N_22468,N_20001,N_20703);
or U22469 (N_22469,N_20843,N_20055);
nand U22470 (N_22470,N_20096,N_21632);
xor U22471 (N_22471,N_20122,N_21141);
and U22472 (N_22472,N_20528,N_20638);
nor U22473 (N_22473,N_20936,N_20447);
nor U22474 (N_22474,N_21515,N_21621);
and U22475 (N_22475,N_20576,N_21070);
nor U22476 (N_22476,N_21787,N_21361);
and U22477 (N_22477,N_21635,N_21803);
or U22478 (N_22478,N_21306,N_20063);
and U22479 (N_22479,N_21156,N_20204);
nor U22480 (N_22480,N_21644,N_20786);
xnor U22481 (N_22481,N_21413,N_20006);
nand U22482 (N_22482,N_20295,N_21421);
or U22483 (N_22483,N_21676,N_20219);
xnor U22484 (N_22484,N_20696,N_21300);
nand U22485 (N_22485,N_21360,N_20391);
nand U22486 (N_22486,N_20964,N_20300);
and U22487 (N_22487,N_21771,N_20586);
xor U22488 (N_22488,N_21629,N_20552);
nand U22489 (N_22489,N_20303,N_21682);
nor U22490 (N_22490,N_20374,N_20364);
xnor U22491 (N_22491,N_21058,N_20128);
xnor U22492 (N_22492,N_20229,N_20200);
nor U22493 (N_22493,N_21132,N_21091);
nand U22494 (N_22494,N_21684,N_21747);
or U22495 (N_22495,N_20078,N_21100);
or U22496 (N_22496,N_20779,N_20592);
nor U22497 (N_22497,N_21736,N_20971);
xnor U22498 (N_22498,N_21655,N_20305);
or U22499 (N_22499,N_21494,N_21651);
nand U22500 (N_22500,N_20251,N_20597);
nand U22501 (N_22501,N_21512,N_21373);
xor U22502 (N_22502,N_21661,N_21962);
or U22503 (N_22503,N_20890,N_20631);
xor U22504 (N_22504,N_21433,N_20056);
nor U22505 (N_22505,N_21331,N_20733);
nor U22506 (N_22506,N_20717,N_21659);
nand U22507 (N_22507,N_21926,N_21588);
or U22508 (N_22508,N_21430,N_21177);
xor U22509 (N_22509,N_20151,N_21420);
and U22510 (N_22510,N_20481,N_20723);
and U22511 (N_22511,N_21221,N_21904);
and U22512 (N_22512,N_21275,N_21844);
nor U22513 (N_22513,N_21063,N_20999);
nor U22514 (N_22514,N_21886,N_21627);
nor U22515 (N_22515,N_21279,N_21869);
nand U22516 (N_22516,N_20785,N_20088);
and U22517 (N_22517,N_20231,N_20538);
xnor U22518 (N_22518,N_20648,N_20049);
nor U22519 (N_22519,N_21922,N_20317);
or U22520 (N_22520,N_20989,N_21448);
nor U22521 (N_22521,N_21267,N_20549);
nand U22522 (N_22522,N_20941,N_21072);
and U22523 (N_22523,N_20603,N_21121);
and U22524 (N_22524,N_20543,N_20763);
and U22525 (N_22525,N_20152,N_21595);
or U22526 (N_22526,N_21866,N_20669);
nand U22527 (N_22527,N_20012,N_21170);
nand U22528 (N_22528,N_20841,N_21101);
nor U22529 (N_22529,N_21618,N_21376);
nand U22530 (N_22530,N_21847,N_20338);
xnor U22531 (N_22531,N_20661,N_21680);
nor U22532 (N_22532,N_21591,N_21117);
nand U22533 (N_22533,N_21827,N_20495);
xnor U22534 (N_22534,N_21229,N_20518);
and U22535 (N_22535,N_21984,N_21226);
nand U22536 (N_22536,N_21725,N_21435);
or U22537 (N_22537,N_20512,N_21611);
nor U22538 (N_22538,N_20577,N_20007);
and U22539 (N_22539,N_21284,N_20240);
nand U22540 (N_22540,N_20470,N_21881);
nor U22541 (N_22541,N_21813,N_20159);
and U22542 (N_22542,N_21380,N_20666);
nor U22543 (N_22543,N_21503,N_20291);
or U22544 (N_22544,N_21481,N_21686);
nor U22545 (N_22545,N_21675,N_20418);
or U22546 (N_22546,N_20676,N_21135);
xnor U22547 (N_22547,N_21168,N_21545);
nand U22548 (N_22548,N_21811,N_20599);
xor U22549 (N_22549,N_21549,N_21965);
and U22550 (N_22550,N_21734,N_21110);
nor U22551 (N_22551,N_21422,N_20687);
xor U22552 (N_22552,N_20665,N_21210);
nor U22553 (N_22553,N_20214,N_20976);
or U22554 (N_22554,N_20811,N_21942);
or U22555 (N_22555,N_20476,N_21172);
and U22556 (N_22556,N_20326,N_21490);
or U22557 (N_22557,N_20255,N_21849);
nand U22558 (N_22558,N_20598,N_20356);
nor U22559 (N_22559,N_21297,N_20985);
and U22560 (N_22560,N_20324,N_21468);
and U22561 (N_22561,N_20566,N_21950);
and U22562 (N_22562,N_21785,N_21607);
xnor U22563 (N_22563,N_21530,N_20732);
xnor U22564 (N_22564,N_20494,N_20483);
nor U22565 (N_22565,N_21505,N_21598);
nor U22566 (N_22566,N_20958,N_21233);
xnor U22567 (N_22567,N_20040,N_21323);
nor U22568 (N_22568,N_20583,N_20213);
nor U22569 (N_22569,N_21002,N_20531);
nor U22570 (N_22570,N_20988,N_21147);
and U22571 (N_22571,N_20212,N_21145);
or U22572 (N_22572,N_20690,N_20716);
or U22573 (N_22573,N_20919,N_20776);
xor U22574 (N_22574,N_21601,N_20728);
and U22575 (N_22575,N_21137,N_21525);
nor U22576 (N_22576,N_20513,N_21196);
nor U22577 (N_22577,N_20842,N_21624);
nand U22578 (N_22578,N_21290,N_20424);
xor U22579 (N_22579,N_21302,N_20148);
nand U22580 (N_22580,N_20472,N_20746);
xor U22581 (N_22581,N_20609,N_20034);
xor U22582 (N_22582,N_20659,N_20944);
or U22583 (N_22583,N_21777,N_20917);
or U22584 (N_22584,N_20227,N_21397);
xor U22585 (N_22585,N_21449,N_21307);
or U22586 (N_22586,N_21724,N_20031);
and U22587 (N_22587,N_21436,N_21836);
and U22588 (N_22588,N_21799,N_20038);
xor U22589 (N_22589,N_21088,N_21169);
and U22590 (N_22590,N_21648,N_21826);
xnor U22591 (N_22591,N_21845,N_20207);
xnor U22592 (N_22592,N_20662,N_21750);
and U22593 (N_22593,N_21581,N_21935);
nand U22594 (N_22594,N_21737,N_20571);
and U22595 (N_22595,N_21062,N_20474);
xor U22596 (N_22596,N_20465,N_21459);
or U22597 (N_22597,N_21645,N_21843);
and U22598 (N_22598,N_21868,N_21623);
xnor U22599 (N_22599,N_21854,N_21189);
nor U22600 (N_22600,N_20478,N_21384);
nand U22601 (N_22601,N_20729,N_20438);
or U22602 (N_22602,N_20507,N_20970);
nor U22603 (N_22603,N_21751,N_21244);
nor U22604 (N_22604,N_20036,N_21775);
and U22605 (N_22605,N_20787,N_20041);
nor U22606 (N_22606,N_20961,N_20475);
xnor U22607 (N_22607,N_21862,N_21120);
and U22608 (N_22608,N_21695,N_20002);
and U22609 (N_22609,N_21573,N_20865);
or U22610 (N_22610,N_21092,N_21401);
and U22611 (N_22611,N_20339,N_21054);
or U22612 (N_22612,N_21492,N_21871);
and U22613 (N_22613,N_20792,N_20946);
nor U22614 (N_22614,N_20024,N_20397);
nor U22615 (N_22615,N_21041,N_21634);
and U22616 (N_22616,N_20816,N_21841);
and U22617 (N_22617,N_20490,N_20102);
and U22618 (N_22618,N_20722,N_21822);
nor U22619 (N_22619,N_21928,N_20614);
xor U22620 (N_22620,N_21786,N_20245);
nor U22621 (N_22621,N_21386,N_20886);
nand U22622 (N_22622,N_21067,N_21939);
and U22623 (N_22623,N_20881,N_21979);
or U22624 (N_22624,N_20929,N_20656);
nand U22625 (N_22625,N_21052,N_21357);
or U22626 (N_22626,N_20312,N_20069);
or U22627 (N_22627,N_20878,N_21203);
xnor U22628 (N_22628,N_21951,N_20115);
nor U22629 (N_22629,N_20149,N_20280);
nor U22630 (N_22630,N_21760,N_21696);
or U22631 (N_22631,N_20905,N_21231);
and U22632 (N_22632,N_20145,N_21322);
and U22633 (N_22633,N_21266,N_21969);
and U22634 (N_22634,N_21319,N_21216);
nand U22635 (N_22635,N_20093,N_21442);
and U22636 (N_22636,N_21381,N_21491);
and U22637 (N_22637,N_20569,N_21498);
and U22638 (N_22638,N_20632,N_21677);
or U22639 (N_22639,N_20684,N_21812);
or U22640 (N_22640,N_21457,N_21046);
nor U22641 (N_22641,N_21218,N_20466);
nor U22642 (N_22642,N_20934,N_20035);
or U22643 (N_22643,N_21128,N_20134);
xnor U22644 (N_22644,N_20209,N_21681);
nor U22645 (N_22645,N_21990,N_21273);
xnor U22646 (N_22646,N_20146,N_21069);
xnor U22647 (N_22647,N_21669,N_21249);
nor U22648 (N_22648,N_21129,N_20017);
or U22649 (N_22649,N_20916,N_20912);
xnor U22650 (N_22650,N_21679,N_20186);
xor U22651 (N_22651,N_21544,N_20355);
nand U22652 (N_22652,N_20450,N_21017);
xnor U22653 (N_22653,N_21902,N_20334);
nor U22654 (N_22654,N_21183,N_20127);
nor U22655 (N_22655,N_21905,N_20913);
nand U22656 (N_22656,N_21312,N_20914);
or U22657 (N_22657,N_21723,N_21301);
nor U22658 (N_22658,N_21643,N_20923);
nand U22659 (N_22659,N_20554,N_21346);
nor U22660 (N_22660,N_20596,N_20664);
or U22661 (N_22661,N_21614,N_21735);
xnor U22662 (N_22662,N_21412,N_21202);
or U22663 (N_22663,N_20047,N_20389);
nand U22664 (N_22664,N_20371,N_20582);
nor U22665 (N_22665,N_20311,N_20267);
xnor U22666 (N_22666,N_20403,N_21247);
xnor U22667 (N_22667,N_20727,N_20349);
nor U22668 (N_22668,N_20516,N_21758);
nand U22669 (N_22669,N_20284,N_21701);
nand U22670 (N_22670,N_20741,N_20220);
nand U22671 (N_22671,N_21819,N_20032);
nor U22672 (N_22672,N_21517,N_20155);
nor U22673 (N_22673,N_20856,N_21536);
or U22674 (N_22674,N_21377,N_20997);
nand U22675 (N_22675,N_21610,N_21368);
xor U22676 (N_22676,N_20630,N_20430);
xor U22677 (N_22677,N_21374,N_21916);
or U22678 (N_22678,N_21424,N_20118);
and U22679 (N_22679,N_20042,N_21036);
and U22680 (N_22680,N_21042,N_20092);
or U22681 (N_22681,N_21529,N_20082);
and U22682 (N_22682,N_21774,N_20782);
xnor U22683 (N_22683,N_20889,N_21974);
nor U22684 (N_22684,N_21182,N_20202);
nand U22685 (N_22685,N_21996,N_21138);
nand U22686 (N_22686,N_20555,N_21144);
and U22687 (N_22687,N_20950,N_21446);
or U22688 (N_22688,N_20337,N_20542);
and U22689 (N_22689,N_20911,N_20064);
nand U22690 (N_22690,N_21678,N_20445);
and U22691 (N_22691,N_21294,N_21105);
nor U22692 (N_22692,N_20697,N_21555);
nand U22693 (N_22693,N_21458,N_20639);
nand U22694 (N_22694,N_20615,N_21118);
nand U22695 (N_22695,N_20500,N_20871);
nand U22696 (N_22696,N_21589,N_20595);
and U22697 (N_22697,N_21713,N_20194);
or U22698 (N_22698,N_20176,N_20320);
nand U22699 (N_22699,N_21647,N_21352);
or U22700 (N_22700,N_21460,N_21152);
nor U22701 (N_22701,N_21946,N_20892);
or U22702 (N_22702,N_21253,N_21287);
nor U22703 (N_22703,N_20028,N_21792);
and U22704 (N_22704,N_21228,N_21499);
nand U22705 (N_22705,N_21732,N_20030);
xnor U22706 (N_22706,N_20852,N_20731);
or U22707 (N_22707,N_20708,N_20187);
and U22708 (N_22708,N_20094,N_21672);
or U22709 (N_22709,N_20910,N_20616);
or U22710 (N_22710,N_20279,N_21086);
and U22711 (N_22711,N_21936,N_20822);
nand U22712 (N_22712,N_21980,N_21043);
or U22713 (N_22713,N_21994,N_21665);
or U22714 (N_22714,N_20984,N_20548);
and U22715 (N_22715,N_20640,N_20120);
nor U22716 (N_22716,N_20429,N_21343);
nor U22717 (N_22717,N_20116,N_20444);
nor U22718 (N_22718,N_21076,N_20443);
or U22719 (N_22719,N_20874,N_20211);
xor U22720 (N_22720,N_20519,N_21461);
or U22721 (N_22721,N_21832,N_20751);
nand U22722 (N_22722,N_21032,N_21744);
and U22723 (N_22723,N_20744,N_20169);
nor U22724 (N_22724,N_21001,N_20850);
xnor U22725 (N_22725,N_21662,N_21642);
or U22726 (N_22726,N_20301,N_20767);
and U22727 (N_22727,N_20574,N_21212);
and U22728 (N_22728,N_20180,N_20137);
nand U22729 (N_22729,N_21764,N_20649);
or U22730 (N_22730,N_20126,N_20353);
xnor U22731 (N_22731,N_20170,N_20307);
and U22732 (N_22732,N_21839,N_20996);
and U22733 (N_22733,N_21532,N_20805);
and U22734 (N_22734,N_21788,N_20761);
or U22735 (N_22735,N_21889,N_20399);
nand U22736 (N_22736,N_21875,N_20688);
nor U22737 (N_22737,N_20261,N_20700);
xor U22738 (N_22738,N_21716,N_20511);
and U22739 (N_22739,N_21861,N_21122);
xnor U22740 (N_22740,N_20310,N_21207);
xnor U22741 (N_22741,N_20951,N_21619);
nand U22742 (N_22742,N_20256,N_21562);
nand U22743 (N_22743,N_21901,N_20097);
nor U22744 (N_22744,N_21838,N_21739);
nor U22745 (N_22745,N_21230,N_21232);
xnor U22746 (N_22746,N_21033,N_21860);
nand U22747 (N_22747,N_20624,N_21347);
or U22748 (N_22748,N_21874,N_20607);
and U22749 (N_22749,N_20677,N_21048);
or U22750 (N_22750,N_21034,N_21704);
or U22751 (N_22751,N_20248,N_21345);
nand U22752 (N_22752,N_20673,N_20879);
and U22753 (N_22753,N_21378,N_21749);
xor U22754 (N_22754,N_21745,N_21471);
xnor U22755 (N_22755,N_20130,N_20375);
nand U22756 (N_22756,N_20660,N_20774);
xor U22757 (N_22757,N_20933,N_21567);
or U22758 (N_22758,N_20719,N_20414);
nor U22759 (N_22759,N_21638,N_20698);
nand U22760 (N_22760,N_20977,N_21019);
or U22761 (N_22761,N_21317,N_21215);
xor U22762 (N_22762,N_20218,N_20423);
nand U22763 (N_22763,N_21523,N_21637);
nand U22764 (N_22764,N_20858,N_20292);
nand U22765 (N_22765,N_21689,N_20972);
and U22766 (N_22766,N_21592,N_20268);
or U22767 (N_22767,N_20144,N_21507);
or U22768 (N_22768,N_20163,N_20835);
xor U22769 (N_22769,N_21550,N_20440);
nor U22770 (N_22770,N_21880,N_21608);
or U22771 (N_22771,N_20119,N_20633);
nand U22772 (N_22772,N_21630,N_21362);
nand U22773 (N_22773,N_21579,N_21403);
nor U22774 (N_22774,N_21652,N_20803);
or U22775 (N_22775,N_21130,N_20726);
nand U22776 (N_22776,N_21028,N_20920);
xnor U22777 (N_22777,N_20086,N_20568);
xnor U22778 (N_22778,N_20584,N_20529);
nor U22779 (N_22779,N_21687,N_20439);
nor U22780 (N_22780,N_20221,N_21919);
nand U22781 (N_22781,N_20738,N_21526);
nand U22782 (N_22782,N_20957,N_21564);
xor U22783 (N_22783,N_21756,N_21561);
and U22784 (N_22784,N_21949,N_20504);
or U22785 (N_22785,N_21021,N_21717);
or U22786 (N_22786,N_21649,N_20344);
nor U22787 (N_22787,N_20108,N_20563);
nor U22788 (N_22788,N_21004,N_20724);
nand U22789 (N_22789,N_20408,N_20517);
nor U22790 (N_22790,N_21060,N_21389);
or U22791 (N_22791,N_21605,N_21557);
nor U22792 (N_22792,N_20861,N_21606);
and U22793 (N_22793,N_20464,N_20872);
xnor U22794 (N_22794,N_20927,N_20080);
nand U22795 (N_22795,N_20613,N_20593);
xor U22796 (N_22796,N_21309,N_20866);
and U22797 (N_22797,N_21234,N_21594);
xnor U22798 (N_22798,N_20848,N_21653);
nand U22799 (N_22799,N_20594,N_20406);
nand U22800 (N_22800,N_20413,N_21318);
nor U22801 (N_22801,N_21998,N_20000);
xor U22802 (N_22802,N_21333,N_20393);
nand U22803 (N_22803,N_21707,N_20983);
or U22804 (N_22804,N_20366,N_21165);
and U22805 (N_22805,N_21089,N_20357);
nor U22806 (N_22806,N_20270,N_20045);
nand U22807 (N_22807,N_20798,N_21371);
xnor U22808 (N_22808,N_21995,N_20973);
nand U22809 (N_22809,N_21064,N_21987);
or U22810 (N_22810,N_21268,N_20057);
xnor U22811 (N_22811,N_20812,N_20832);
and U22812 (N_22812,N_20998,N_20515);
or U22813 (N_22813,N_21781,N_21762);
nand U22814 (N_22814,N_21012,N_20817);
xnor U22815 (N_22815,N_20479,N_21513);
xnor U22816 (N_22816,N_20452,N_20411);
nand U22817 (N_22817,N_20296,N_21636);
nor U22818 (N_22818,N_21220,N_20537);
nand U22819 (N_22819,N_21872,N_21898);
nand U22820 (N_22820,N_21640,N_20888);
or U22821 (N_22821,N_20416,N_21801);
nand U22822 (N_22822,N_21007,N_21480);
or U22823 (N_22823,N_20410,N_21851);
nand U22824 (N_22824,N_20425,N_21952);
nor U22825 (N_22825,N_21670,N_20361);
xor U22826 (N_22826,N_20288,N_20691);
or U22827 (N_22827,N_21326,N_20259);
nand U22828 (N_22828,N_21920,N_20191);
and U22829 (N_22829,N_20241,N_21944);
and U22830 (N_22830,N_20282,N_21181);
and U22831 (N_22831,N_21855,N_20993);
or U22832 (N_22832,N_20939,N_21616);
and U22833 (N_22833,N_20980,N_21842);
nor U22834 (N_22834,N_20820,N_21200);
xnor U22835 (N_22835,N_21425,N_20809);
and U22836 (N_22836,N_20239,N_20074);
nor U22837 (N_22837,N_20756,N_20651);
or U22838 (N_22838,N_21367,N_20600);
or U22839 (N_22839,N_20004,N_21350);
or U22840 (N_22840,N_20053,N_21087);
or U22841 (N_22841,N_21719,N_20249);
xnor U22842 (N_22842,N_20947,N_21428);
or U22843 (N_22843,N_20333,N_20362);
nand U22844 (N_22844,N_20343,N_21276);
xor U22845 (N_22845,N_21917,N_20412);
xnor U22846 (N_22846,N_21533,N_20238);
nand U22847 (N_22847,N_20014,N_21795);
nand U22848 (N_22848,N_21180,N_21553);
xnor U22849 (N_22849,N_21404,N_20784);
or U22850 (N_22850,N_20046,N_21166);
or U22851 (N_22851,N_20287,N_20590);
nor U22852 (N_22852,N_21528,N_20829);
or U22853 (N_22853,N_21292,N_21947);
and U22854 (N_22854,N_21915,N_21502);
xor U22855 (N_22855,N_20325,N_20420);
nor U22856 (N_22856,N_20940,N_20508);
nor U22857 (N_22857,N_20625,N_21227);
or U22858 (N_22858,N_21414,N_20501);
xor U22859 (N_22859,N_20875,N_20264);
xor U22860 (N_22860,N_20668,N_20619);
or U22861 (N_22861,N_21534,N_21470);
and U22862 (N_22862,N_21338,N_21194);
or U22863 (N_22863,N_21112,N_20446);
and U22864 (N_22864,N_21909,N_20788);
and U22865 (N_22865,N_21093,N_20210);
or U22866 (N_22866,N_20860,N_20707);
nand U22867 (N_22867,N_20954,N_20013);
nor U22868 (N_22868,N_20689,N_21703);
and U22869 (N_22869,N_20702,N_21563);
xor U22870 (N_22870,N_20103,N_21722);
nand U22871 (N_22871,N_21372,N_20079);
and U22872 (N_22872,N_21992,N_21654);
or U22873 (N_22873,N_20405,N_21547);
nor U22874 (N_22874,N_21691,N_21159);
and U22875 (N_22875,N_20396,N_21489);
and U22876 (N_22876,N_20449,N_20377);
or U22877 (N_22877,N_20834,N_20524);
xnor U22878 (N_22878,N_21824,N_20175);
nor U22879 (N_22879,N_20969,N_20019);
nand U22880 (N_22880,N_21715,N_21921);
xnor U22881 (N_22881,N_20316,N_21201);
xor U22882 (N_22882,N_21008,N_20589);
nand U22883 (N_22883,N_21164,N_21509);
nor U22884 (N_22884,N_21748,N_20234);
and U22885 (N_22885,N_20071,N_21355);
nand U22886 (N_22886,N_21893,N_21729);
or U22887 (N_22887,N_20755,N_21071);
and U22888 (N_22888,N_20428,N_20570);
xor U22889 (N_22889,N_20113,N_21429);
nor U22890 (N_22890,N_20540,N_20672);
or U22891 (N_22891,N_20556,N_20199);
nor U22892 (N_22892,N_21894,N_21341);
or U22893 (N_22893,N_21896,N_21375);
xor U22894 (N_22894,N_20331,N_21022);
nor U22895 (N_22895,N_20252,N_20827);
or U22896 (N_22896,N_20488,N_21770);
nand U22897 (N_22897,N_21245,N_21464);
nand U22898 (N_22898,N_20506,N_21195);
or U22899 (N_22899,N_21124,N_20605);
and U22900 (N_22900,N_21497,N_20748);
xor U22901 (N_22901,N_20558,N_20992);
xnor U22902 (N_22902,N_21978,N_21217);
or U22903 (N_22903,N_20286,N_21288);
xor U22904 (N_22904,N_20269,N_21025);
nor U22905 (N_22905,N_20360,N_20794);
or U22906 (N_22906,N_21559,N_20027);
nand U22907 (N_22907,N_20341,N_20294);
nand U22908 (N_22908,N_20991,N_20369);
xnor U22909 (N_22909,N_21504,N_21176);
and U22910 (N_22910,N_21262,N_21833);
nor U22911 (N_22911,N_21015,N_20503);
and U22912 (N_22912,N_20265,N_20833);
nor U22913 (N_22913,N_20562,N_20266);
nand U22914 (N_22914,N_20434,N_20228);
nand U22915 (N_22915,N_20484,N_20610);
or U22916 (N_22916,N_21363,N_20773);
nor U22917 (N_22917,N_20347,N_21455);
and U22918 (N_22918,N_21197,N_20328);
xor U22919 (N_22919,N_21899,N_21027);
or U22920 (N_22920,N_20051,N_20602);
xnor U22921 (N_22921,N_20401,N_20025);
xor U22922 (N_22922,N_20072,N_21073);
nand U22923 (N_22923,N_21327,N_20409);
or U22924 (N_22924,N_20385,N_21416);
nand U22925 (N_22925,N_21699,N_20734);
nand U22926 (N_22926,N_21256,N_21569);
and U22927 (N_22927,N_20381,N_20928);
xor U22928 (N_22928,N_20246,N_20846);
or U22929 (N_22929,N_21968,N_21055);
nand U22930 (N_22930,N_21310,N_20573);
nand U22931 (N_22931,N_20935,N_20762);
nor U22932 (N_22932,N_20117,N_20455);
nand U22933 (N_22933,N_21325,N_20323);
xnor U22934 (N_22934,N_21495,N_20880);
or U22935 (N_22935,N_21911,N_21030);
nor U22936 (N_22936,N_21260,N_21767);
xor U22937 (N_22937,N_21778,N_21014);
nor U22938 (N_22938,N_21846,N_21955);
xor U22939 (N_22939,N_20932,N_21097);
xor U22940 (N_22940,N_20765,N_21104);
and U22941 (N_22941,N_20281,N_20974);
and U22942 (N_22942,N_21863,N_21897);
nor U22943 (N_22943,N_21291,N_20814);
and U22944 (N_22944,N_20710,N_21272);
or U22945 (N_22945,N_21793,N_20129);
and U22946 (N_22946,N_20712,N_20112);
xor U22947 (N_22947,N_21274,N_20948);
and U22948 (N_22948,N_21315,N_21511);
xnor U22949 (N_22949,N_20486,N_20553);
nor U22950 (N_22950,N_21099,N_20900);
nor U22951 (N_22951,N_21193,N_20899);
nor U22952 (N_22952,N_21040,N_21265);
xor U22953 (N_22953,N_21474,N_20222);
nand U22954 (N_22954,N_21802,N_20818);
and U22955 (N_22955,N_21705,N_21438);
xnor U22956 (N_22956,N_20319,N_20435);
or U22957 (N_22957,N_20617,N_21837);
and U22958 (N_22958,N_21556,N_20184);
nor U22959 (N_22959,N_21964,N_20953);
or U22960 (N_22960,N_20235,N_21519);
or U22961 (N_22961,N_21410,N_20171);
and U22962 (N_22962,N_20496,N_20289);
and U22963 (N_22963,N_21746,N_21690);
nor U22964 (N_22964,N_21411,N_20247);
and U22965 (N_22965,N_20618,N_20433);
nand U22966 (N_22966,N_20336,N_21280);
or U22967 (N_22967,N_20686,N_21264);
nand U22968 (N_22968,N_20830,N_21496);
nor U22969 (N_22969,N_21565,N_20533);
nand U22970 (N_22970,N_20165,N_21817);
and U22971 (N_22971,N_21663,N_20681);
xnor U22972 (N_22972,N_20545,N_21190);
nand U22973 (N_22973,N_20663,N_20918);
and U22974 (N_22974,N_21789,N_21131);
or U22975 (N_22975,N_21805,N_21885);
and U22976 (N_22976,N_20510,N_21005);
or U22977 (N_22977,N_20646,N_21997);
nand U22978 (N_22978,N_20565,N_21477);
nand U22979 (N_22979,N_20015,N_20309);
nand U22980 (N_22980,N_20315,N_20781);
and U22981 (N_22981,N_20760,N_20254);
nor U22982 (N_22982,N_20643,N_21712);
and U22983 (N_22983,N_21959,N_20290);
or U22984 (N_22984,N_20253,N_21255);
nor U22985 (N_22985,N_21452,N_20367);
xnor U22986 (N_22986,N_20147,N_20641);
and U22987 (N_22987,N_21243,N_20750);
or U22988 (N_22988,N_20925,N_20075);
and U22989 (N_22989,N_21139,N_21796);
and U22990 (N_22990,N_21551,N_21175);
nand U22991 (N_22991,N_20083,N_20263);
nor U22992 (N_22992,N_20658,N_20851);
and U22993 (N_22993,N_20828,N_21402);
nand U22994 (N_22994,N_21548,N_20808);
and U22995 (N_22995,N_21711,N_20931);
and U22996 (N_22996,N_21366,N_21311);
or U22997 (N_22997,N_21685,N_21852);
xnor U22998 (N_22998,N_21765,N_21106);
and U22999 (N_22999,N_20521,N_20530);
nor U23000 (N_23000,N_20629,N_21523);
nand U23001 (N_23001,N_20330,N_20418);
nor U23002 (N_23002,N_20350,N_20319);
or U23003 (N_23003,N_21234,N_21299);
xnor U23004 (N_23004,N_21736,N_20807);
nand U23005 (N_23005,N_21022,N_20717);
or U23006 (N_23006,N_20627,N_20069);
or U23007 (N_23007,N_20933,N_21354);
nand U23008 (N_23008,N_21471,N_21547);
and U23009 (N_23009,N_21444,N_21057);
and U23010 (N_23010,N_20039,N_20958);
xnor U23011 (N_23011,N_21706,N_21527);
or U23012 (N_23012,N_21792,N_21396);
and U23013 (N_23013,N_20021,N_21921);
nand U23014 (N_23014,N_20646,N_21611);
nand U23015 (N_23015,N_20684,N_20229);
xor U23016 (N_23016,N_20591,N_20306);
nor U23017 (N_23017,N_20212,N_21413);
and U23018 (N_23018,N_21090,N_20122);
xnor U23019 (N_23019,N_20715,N_21955);
nor U23020 (N_23020,N_21632,N_20682);
xor U23021 (N_23021,N_21204,N_21758);
nor U23022 (N_23022,N_21742,N_21718);
or U23023 (N_23023,N_21637,N_21493);
nand U23024 (N_23024,N_21742,N_21610);
xnor U23025 (N_23025,N_20403,N_21904);
or U23026 (N_23026,N_21994,N_21801);
xnor U23027 (N_23027,N_20204,N_20092);
nand U23028 (N_23028,N_20321,N_20512);
nor U23029 (N_23029,N_20467,N_20728);
nor U23030 (N_23030,N_20751,N_20914);
nand U23031 (N_23031,N_20979,N_20052);
nand U23032 (N_23032,N_20859,N_20123);
xor U23033 (N_23033,N_20727,N_20699);
nor U23034 (N_23034,N_20792,N_21390);
nor U23035 (N_23035,N_21291,N_21949);
nor U23036 (N_23036,N_21003,N_20918);
or U23037 (N_23037,N_20954,N_20147);
and U23038 (N_23038,N_21310,N_20537);
and U23039 (N_23039,N_20870,N_21470);
or U23040 (N_23040,N_21017,N_20638);
xnor U23041 (N_23041,N_20813,N_20827);
nor U23042 (N_23042,N_21567,N_20264);
or U23043 (N_23043,N_20987,N_21428);
and U23044 (N_23044,N_20793,N_20744);
xor U23045 (N_23045,N_20773,N_21985);
and U23046 (N_23046,N_21248,N_20623);
or U23047 (N_23047,N_21342,N_21750);
nand U23048 (N_23048,N_21091,N_20286);
or U23049 (N_23049,N_20662,N_21395);
nand U23050 (N_23050,N_20494,N_20056);
nor U23051 (N_23051,N_20143,N_20551);
nor U23052 (N_23052,N_20403,N_20394);
and U23053 (N_23053,N_21851,N_20164);
or U23054 (N_23054,N_21871,N_21732);
nor U23055 (N_23055,N_21202,N_21170);
nor U23056 (N_23056,N_21579,N_21333);
xor U23057 (N_23057,N_20816,N_20390);
nand U23058 (N_23058,N_20513,N_20656);
nand U23059 (N_23059,N_20966,N_21964);
xor U23060 (N_23060,N_21390,N_21897);
nor U23061 (N_23061,N_21026,N_20747);
xor U23062 (N_23062,N_21536,N_20444);
and U23063 (N_23063,N_21327,N_20953);
nor U23064 (N_23064,N_20208,N_21178);
or U23065 (N_23065,N_21663,N_20392);
nand U23066 (N_23066,N_21737,N_20356);
xor U23067 (N_23067,N_21698,N_20560);
xor U23068 (N_23068,N_20557,N_20020);
xnor U23069 (N_23069,N_20475,N_20376);
nand U23070 (N_23070,N_20825,N_20371);
and U23071 (N_23071,N_20211,N_20359);
nand U23072 (N_23072,N_21210,N_20815);
xnor U23073 (N_23073,N_20675,N_21980);
nand U23074 (N_23074,N_20463,N_21102);
nor U23075 (N_23075,N_21287,N_21732);
or U23076 (N_23076,N_21680,N_21031);
and U23077 (N_23077,N_21936,N_20879);
nor U23078 (N_23078,N_20052,N_21004);
nand U23079 (N_23079,N_21692,N_20151);
and U23080 (N_23080,N_21203,N_21803);
nand U23081 (N_23081,N_21451,N_20477);
nand U23082 (N_23082,N_21202,N_21529);
and U23083 (N_23083,N_20417,N_21620);
xnor U23084 (N_23084,N_21862,N_21815);
nand U23085 (N_23085,N_20975,N_20165);
and U23086 (N_23086,N_21398,N_20689);
xor U23087 (N_23087,N_21252,N_20684);
or U23088 (N_23088,N_20305,N_20695);
nand U23089 (N_23089,N_20048,N_21835);
and U23090 (N_23090,N_21109,N_21057);
nor U23091 (N_23091,N_21727,N_21365);
and U23092 (N_23092,N_21397,N_21106);
nor U23093 (N_23093,N_20690,N_20521);
or U23094 (N_23094,N_21079,N_20699);
nor U23095 (N_23095,N_20029,N_20781);
or U23096 (N_23096,N_21166,N_20133);
and U23097 (N_23097,N_21786,N_20709);
and U23098 (N_23098,N_20749,N_21374);
or U23099 (N_23099,N_21148,N_20207);
xor U23100 (N_23100,N_20905,N_21899);
nand U23101 (N_23101,N_21777,N_20776);
or U23102 (N_23102,N_21588,N_20213);
and U23103 (N_23103,N_21840,N_20505);
nand U23104 (N_23104,N_20185,N_20404);
nor U23105 (N_23105,N_20144,N_20947);
and U23106 (N_23106,N_21757,N_21176);
nand U23107 (N_23107,N_20949,N_20823);
or U23108 (N_23108,N_20207,N_20502);
and U23109 (N_23109,N_21981,N_20302);
nor U23110 (N_23110,N_21496,N_21798);
nand U23111 (N_23111,N_20336,N_20991);
nor U23112 (N_23112,N_21370,N_21845);
xnor U23113 (N_23113,N_20359,N_20292);
xor U23114 (N_23114,N_21080,N_21274);
nand U23115 (N_23115,N_21333,N_21158);
and U23116 (N_23116,N_20777,N_21637);
and U23117 (N_23117,N_20903,N_20512);
nand U23118 (N_23118,N_20808,N_20214);
nand U23119 (N_23119,N_20728,N_20688);
or U23120 (N_23120,N_20176,N_20855);
or U23121 (N_23121,N_21010,N_21463);
or U23122 (N_23122,N_21460,N_21706);
and U23123 (N_23123,N_21192,N_20454);
xnor U23124 (N_23124,N_21832,N_20930);
or U23125 (N_23125,N_20986,N_21641);
and U23126 (N_23126,N_20247,N_21543);
nor U23127 (N_23127,N_21908,N_20574);
nand U23128 (N_23128,N_21200,N_20897);
nand U23129 (N_23129,N_21658,N_20760);
nor U23130 (N_23130,N_20021,N_20988);
or U23131 (N_23131,N_21088,N_21539);
or U23132 (N_23132,N_20593,N_20970);
nand U23133 (N_23133,N_21772,N_21860);
and U23134 (N_23134,N_20230,N_21346);
and U23135 (N_23135,N_20057,N_20276);
nand U23136 (N_23136,N_20524,N_21344);
nand U23137 (N_23137,N_21850,N_21972);
or U23138 (N_23138,N_20113,N_21241);
xnor U23139 (N_23139,N_21831,N_20530);
and U23140 (N_23140,N_21578,N_20942);
xor U23141 (N_23141,N_21804,N_20099);
and U23142 (N_23142,N_21101,N_20607);
or U23143 (N_23143,N_21953,N_20501);
nand U23144 (N_23144,N_20650,N_21672);
or U23145 (N_23145,N_21169,N_21050);
nor U23146 (N_23146,N_21304,N_21354);
nor U23147 (N_23147,N_20573,N_21607);
and U23148 (N_23148,N_20971,N_20240);
nor U23149 (N_23149,N_21459,N_20694);
and U23150 (N_23150,N_20387,N_20982);
xor U23151 (N_23151,N_20217,N_21025);
nor U23152 (N_23152,N_21434,N_20315);
nand U23153 (N_23153,N_21040,N_20973);
nor U23154 (N_23154,N_21953,N_20821);
or U23155 (N_23155,N_21510,N_20393);
nor U23156 (N_23156,N_21267,N_20033);
nand U23157 (N_23157,N_20257,N_21567);
nor U23158 (N_23158,N_20476,N_20760);
xor U23159 (N_23159,N_21548,N_20227);
or U23160 (N_23160,N_20443,N_21391);
nor U23161 (N_23161,N_21381,N_20440);
xor U23162 (N_23162,N_21464,N_21968);
or U23163 (N_23163,N_21316,N_21200);
and U23164 (N_23164,N_20149,N_20360);
nor U23165 (N_23165,N_21935,N_21002);
or U23166 (N_23166,N_21399,N_21646);
nor U23167 (N_23167,N_20722,N_21004);
nand U23168 (N_23168,N_21882,N_20468);
nor U23169 (N_23169,N_20625,N_20815);
xnor U23170 (N_23170,N_20886,N_21131);
or U23171 (N_23171,N_20965,N_20521);
and U23172 (N_23172,N_20638,N_20438);
and U23173 (N_23173,N_21362,N_20923);
nand U23174 (N_23174,N_20612,N_20471);
and U23175 (N_23175,N_21239,N_21251);
and U23176 (N_23176,N_21377,N_20646);
xor U23177 (N_23177,N_20346,N_20250);
nand U23178 (N_23178,N_20475,N_21196);
or U23179 (N_23179,N_20014,N_21921);
and U23180 (N_23180,N_21306,N_21757);
nand U23181 (N_23181,N_20210,N_21807);
nand U23182 (N_23182,N_20863,N_21895);
or U23183 (N_23183,N_21597,N_21692);
xor U23184 (N_23184,N_21122,N_21334);
and U23185 (N_23185,N_20823,N_20391);
and U23186 (N_23186,N_20043,N_21398);
nand U23187 (N_23187,N_21878,N_20853);
and U23188 (N_23188,N_20637,N_21525);
xor U23189 (N_23189,N_20581,N_20869);
or U23190 (N_23190,N_20415,N_20129);
or U23191 (N_23191,N_21416,N_21359);
xor U23192 (N_23192,N_20465,N_21759);
or U23193 (N_23193,N_21092,N_20957);
nand U23194 (N_23194,N_20684,N_20285);
nand U23195 (N_23195,N_21552,N_20847);
or U23196 (N_23196,N_20658,N_21089);
and U23197 (N_23197,N_20268,N_21491);
nor U23198 (N_23198,N_20270,N_20264);
nand U23199 (N_23199,N_21816,N_20842);
or U23200 (N_23200,N_21645,N_21865);
xor U23201 (N_23201,N_20300,N_20039);
or U23202 (N_23202,N_21534,N_21411);
and U23203 (N_23203,N_20839,N_20770);
nor U23204 (N_23204,N_20279,N_20228);
nand U23205 (N_23205,N_21269,N_20949);
xor U23206 (N_23206,N_21161,N_20516);
or U23207 (N_23207,N_20264,N_20056);
nand U23208 (N_23208,N_20022,N_21103);
nor U23209 (N_23209,N_21628,N_21980);
xnor U23210 (N_23210,N_20560,N_20156);
nor U23211 (N_23211,N_20513,N_21433);
nor U23212 (N_23212,N_20052,N_20740);
or U23213 (N_23213,N_20078,N_21709);
nor U23214 (N_23214,N_21181,N_21271);
xor U23215 (N_23215,N_21314,N_21216);
nor U23216 (N_23216,N_20368,N_21528);
or U23217 (N_23217,N_21537,N_20050);
or U23218 (N_23218,N_20913,N_21529);
nand U23219 (N_23219,N_21111,N_21161);
nor U23220 (N_23220,N_20405,N_20220);
or U23221 (N_23221,N_21134,N_20093);
or U23222 (N_23222,N_20388,N_20923);
or U23223 (N_23223,N_20545,N_21006);
nand U23224 (N_23224,N_20804,N_21961);
nor U23225 (N_23225,N_20145,N_21855);
and U23226 (N_23226,N_20246,N_20159);
and U23227 (N_23227,N_20130,N_20438);
nand U23228 (N_23228,N_20883,N_21894);
xnor U23229 (N_23229,N_20625,N_20769);
nand U23230 (N_23230,N_20602,N_21632);
xor U23231 (N_23231,N_20850,N_21074);
or U23232 (N_23232,N_20864,N_21872);
and U23233 (N_23233,N_21326,N_21594);
and U23234 (N_23234,N_21948,N_21359);
and U23235 (N_23235,N_21560,N_21862);
xor U23236 (N_23236,N_21901,N_20081);
and U23237 (N_23237,N_21497,N_21016);
xor U23238 (N_23238,N_20687,N_20351);
and U23239 (N_23239,N_20370,N_21299);
nor U23240 (N_23240,N_20499,N_21194);
and U23241 (N_23241,N_21920,N_20348);
nor U23242 (N_23242,N_21585,N_21189);
and U23243 (N_23243,N_21006,N_20126);
nand U23244 (N_23244,N_21194,N_20041);
xor U23245 (N_23245,N_20828,N_21116);
xor U23246 (N_23246,N_20461,N_20796);
and U23247 (N_23247,N_21789,N_21031);
nor U23248 (N_23248,N_21138,N_20181);
nand U23249 (N_23249,N_21677,N_20547);
or U23250 (N_23250,N_21354,N_20201);
nand U23251 (N_23251,N_21362,N_21516);
nor U23252 (N_23252,N_20219,N_21745);
xor U23253 (N_23253,N_21640,N_20570);
nor U23254 (N_23254,N_20939,N_21969);
nand U23255 (N_23255,N_20661,N_21008);
nand U23256 (N_23256,N_21221,N_21042);
xnor U23257 (N_23257,N_20518,N_21311);
xor U23258 (N_23258,N_21435,N_20192);
nor U23259 (N_23259,N_21537,N_21640);
nand U23260 (N_23260,N_20949,N_21517);
nand U23261 (N_23261,N_20079,N_20706);
xor U23262 (N_23262,N_21350,N_21971);
nor U23263 (N_23263,N_20728,N_21750);
and U23264 (N_23264,N_20841,N_21156);
or U23265 (N_23265,N_21366,N_21481);
or U23266 (N_23266,N_20125,N_21117);
nor U23267 (N_23267,N_20742,N_20265);
or U23268 (N_23268,N_21730,N_20614);
or U23269 (N_23269,N_20059,N_21792);
xnor U23270 (N_23270,N_20471,N_20240);
nor U23271 (N_23271,N_20840,N_21293);
xnor U23272 (N_23272,N_20338,N_21082);
nand U23273 (N_23273,N_20686,N_20159);
nor U23274 (N_23274,N_20892,N_21591);
xor U23275 (N_23275,N_21760,N_21247);
nand U23276 (N_23276,N_20237,N_21683);
nand U23277 (N_23277,N_20903,N_20613);
nor U23278 (N_23278,N_20612,N_20322);
xor U23279 (N_23279,N_20832,N_20343);
nor U23280 (N_23280,N_20332,N_21957);
xor U23281 (N_23281,N_20797,N_20697);
nor U23282 (N_23282,N_21602,N_20470);
xnor U23283 (N_23283,N_21387,N_20083);
nor U23284 (N_23284,N_21177,N_21610);
nor U23285 (N_23285,N_21634,N_20456);
xnor U23286 (N_23286,N_21126,N_21866);
xnor U23287 (N_23287,N_21096,N_20418);
or U23288 (N_23288,N_20005,N_20750);
nand U23289 (N_23289,N_20609,N_21142);
or U23290 (N_23290,N_21810,N_20391);
nor U23291 (N_23291,N_21701,N_21489);
xor U23292 (N_23292,N_20862,N_21351);
nor U23293 (N_23293,N_21189,N_21725);
nand U23294 (N_23294,N_20376,N_20297);
nor U23295 (N_23295,N_20336,N_21982);
nor U23296 (N_23296,N_21625,N_21034);
nand U23297 (N_23297,N_21024,N_21599);
nand U23298 (N_23298,N_21266,N_21009);
xor U23299 (N_23299,N_20279,N_21084);
xnor U23300 (N_23300,N_21924,N_21894);
nand U23301 (N_23301,N_21037,N_21711);
xnor U23302 (N_23302,N_21732,N_20846);
xnor U23303 (N_23303,N_21435,N_21160);
nor U23304 (N_23304,N_21582,N_21225);
or U23305 (N_23305,N_21062,N_20661);
xor U23306 (N_23306,N_20621,N_21959);
or U23307 (N_23307,N_21009,N_20198);
and U23308 (N_23308,N_20191,N_20899);
nor U23309 (N_23309,N_20640,N_20430);
nand U23310 (N_23310,N_20738,N_21350);
xnor U23311 (N_23311,N_20884,N_21087);
and U23312 (N_23312,N_20333,N_21622);
and U23313 (N_23313,N_20853,N_20640);
or U23314 (N_23314,N_21464,N_21155);
xnor U23315 (N_23315,N_20063,N_21489);
and U23316 (N_23316,N_21087,N_20211);
or U23317 (N_23317,N_21731,N_21450);
xor U23318 (N_23318,N_20625,N_20118);
nand U23319 (N_23319,N_21256,N_21990);
or U23320 (N_23320,N_20321,N_21327);
and U23321 (N_23321,N_20977,N_21273);
xor U23322 (N_23322,N_21613,N_20471);
nand U23323 (N_23323,N_20204,N_21426);
and U23324 (N_23324,N_20874,N_20826);
nor U23325 (N_23325,N_21242,N_21952);
and U23326 (N_23326,N_20680,N_21417);
nor U23327 (N_23327,N_20701,N_21656);
or U23328 (N_23328,N_20965,N_21838);
nor U23329 (N_23329,N_21211,N_21804);
or U23330 (N_23330,N_20997,N_21102);
or U23331 (N_23331,N_20230,N_21238);
xnor U23332 (N_23332,N_21485,N_20648);
nor U23333 (N_23333,N_20339,N_20020);
nand U23334 (N_23334,N_20532,N_20948);
and U23335 (N_23335,N_20749,N_21181);
nand U23336 (N_23336,N_21648,N_21488);
and U23337 (N_23337,N_20772,N_20240);
nand U23338 (N_23338,N_20891,N_20069);
or U23339 (N_23339,N_20538,N_20930);
and U23340 (N_23340,N_21255,N_20431);
nor U23341 (N_23341,N_20008,N_21790);
and U23342 (N_23342,N_20267,N_21602);
xor U23343 (N_23343,N_21765,N_21563);
xnor U23344 (N_23344,N_21046,N_20815);
nor U23345 (N_23345,N_21290,N_21360);
nor U23346 (N_23346,N_20101,N_21843);
and U23347 (N_23347,N_21485,N_20828);
nor U23348 (N_23348,N_21518,N_21542);
nor U23349 (N_23349,N_20713,N_21886);
and U23350 (N_23350,N_21234,N_20624);
nor U23351 (N_23351,N_21563,N_21472);
or U23352 (N_23352,N_20393,N_20695);
or U23353 (N_23353,N_20551,N_20845);
and U23354 (N_23354,N_21125,N_20889);
nand U23355 (N_23355,N_21929,N_21042);
or U23356 (N_23356,N_20464,N_20875);
nor U23357 (N_23357,N_21742,N_20470);
and U23358 (N_23358,N_20193,N_21042);
xnor U23359 (N_23359,N_21059,N_20953);
or U23360 (N_23360,N_20775,N_21379);
or U23361 (N_23361,N_21553,N_20568);
nor U23362 (N_23362,N_20147,N_21306);
and U23363 (N_23363,N_21932,N_21228);
nor U23364 (N_23364,N_21435,N_21115);
and U23365 (N_23365,N_21933,N_21614);
or U23366 (N_23366,N_20164,N_20833);
or U23367 (N_23367,N_20884,N_21081);
and U23368 (N_23368,N_21268,N_21103);
or U23369 (N_23369,N_20867,N_21653);
nor U23370 (N_23370,N_20905,N_20954);
and U23371 (N_23371,N_21826,N_21496);
nor U23372 (N_23372,N_20622,N_20152);
nand U23373 (N_23373,N_21154,N_20689);
and U23374 (N_23374,N_20840,N_21110);
xor U23375 (N_23375,N_20662,N_21188);
or U23376 (N_23376,N_21521,N_21459);
or U23377 (N_23377,N_20249,N_21633);
nand U23378 (N_23378,N_20985,N_21933);
xor U23379 (N_23379,N_21367,N_20345);
xnor U23380 (N_23380,N_21930,N_21409);
nand U23381 (N_23381,N_21424,N_20304);
and U23382 (N_23382,N_21305,N_20776);
nand U23383 (N_23383,N_21326,N_20608);
nor U23384 (N_23384,N_21211,N_20513);
xnor U23385 (N_23385,N_21015,N_21761);
nand U23386 (N_23386,N_20776,N_21541);
nand U23387 (N_23387,N_20538,N_21568);
and U23388 (N_23388,N_20736,N_20785);
nor U23389 (N_23389,N_21594,N_20970);
and U23390 (N_23390,N_20404,N_21386);
nand U23391 (N_23391,N_21613,N_20105);
nand U23392 (N_23392,N_20468,N_21249);
and U23393 (N_23393,N_21017,N_20882);
nand U23394 (N_23394,N_20944,N_21052);
and U23395 (N_23395,N_21698,N_21028);
nor U23396 (N_23396,N_20247,N_21331);
nor U23397 (N_23397,N_20461,N_21053);
nor U23398 (N_23398,N_21110,N_20641);
nand U23399 (N_23399,N_21186,N_21128);
and U23400 (N_23400,N_21482,N_21065);
nor U23401 (N_23401,N_20508,N_20164);
xnor U23402 (N_23402,N_21338,N_21370);
or U23403 (N_23403,N_20698,N_20176);
nor U23404 (N_23404,N_21478,N_20881);
or U23405 (N_23405,N_20725,N_21789);
or U23406 (N_23406,N_21324,N_20071);
and U23407 (N_23407,N_20588,N_21591);
nor U23408 (N_23408,N_20665,N_20363);
xor U23409 (N_23409,N_21334,N_21634);
or U23410 (N_23410,N_21224,N_20892);
nor U23411 (N_23411,N_20750,N_20605);
or U23412 (N_23412,N_21177,N_21266);
xnor U23413 (N_23413,N_20767,N_21167);
nor U23414 (N_23414,N_20452,N_21919);
nor U23415 (N_23415,N_20744,N_20425);
nor U23416 (N_23416,N_21410,N_20793);
and U23417 (N_23417,N_20538,N_20642);
xnor U23418 (N_23418,N_21959,N_20481);
and U23419 (N_23419,N_20169,N_21553);
nor U23420 (N_23420,N_21632,N_20670);
or U23421 (N_23421,N_21841,N_21584);
nand U23422 (N_23422,N_20092,N_20787);
or U23423 (N_23423,N_20437,N_20549);
xnor U23424 (N_23424,N_21862,N_20594);
nor U23425 (N_23425,N_21750,N_21974);
nor U23426 (N_23426,N_21922,N_21773);
nand U23427 (N_23427,N_20210,N_21314);
or U23428 (N_23428,N_20533,N_21069);
nand U23429 (N_23429,N_21706,N_20870);
nor U23430 (N_23430,N_21613,N_20563);
nand U23431 (N_23431,N_20465,N_20679);
nand U23432 (N_23432,N_21826,N_21724);
and U23433 (N_23433,N_20327,N_20908);
xor U23434 (N_23434,N_20514,N_20466);
xnor U23435 (N_23435,N_21745,N_20725);
xnor U23436 (N_23436,N_21901,N_20555);
nand U23437 (N_23437,N_20224,N_21833);
xor U23438 (N_23438,N_21540,N_20694);
and U23439 (N_23439,N_21831,N_20219);
nand U23440 (N_23440,N_20726,N_20150);
and U23441 (N_23441,N_20917,N_21925);
nor U23442 (N_23442,N_21228,N_20132);
nand U23443 (N_23443,N_20454,N_20786);
nand U23444 (N_23444,N_21798,N_21605);
nor U23445 (N_23445,N_20627,N_20326);
and U23446 (N_23446,N_21603,N_20068);
nor U23447 (N_23447,N_21951,N_20524);
nand U23448 (N_23448,N_20866,N_21373);
nand U23449 (N_23449,N_21951,N_20662);
and U23450 (N_23450,N_21660,N_21560);
nor U23451 (N_23451,N_20645,N_21500);
and U23452 (N_23452,N_20172,N_20020);
xor U23453 (N_23453,N_21394,N_20342);
nand U23454 (N_23454,N_20421,N_21744);
nand U23455 (N_23455,N_21658,N_20834);
and U23456 (N_23456,N_21738,N_21907);
xnor U23457 (N_23457,N_21514,N_21510);
nand U23458 (N_23458,N_21159,N_21499);
and U23459 (N_23459,N_20113,N_20411);
nor U23460 (N_23460,N_20888,N_21035);
or U23461 (N_23461,N_21001,N_21747);
xor U23462 (N_23462,N_20485,N_21089);
and U23463 (N_23463,N_20329,N_21847);
and U23464 (N_23464,N_20522,N_20985);
xnor U23465 (N_23465,N_20437,N_21379);
or U23466 (N_23466,N_20408,N_20242);
nor U23467 (N_23467,N_20565,N_20658);
nor U23468 (N_23468,N_21708,N_20249);
nand U23469 (N_23469,N_21526,N_21976);
xor U23470 (N_23470,N_20917,N_20939);
nand U23471 (N_23471,N_20940,N_20460);
xor U23472 (N_23472,N_21700,N_21826);
nor U23473 (N_23473,N_21768,N_21749);
or U23474 (N_23474,N_21199,N_20006);
nand U23475 (N_23475,N_21755,N_21411);
or U23476 (N_23476,N_20687,N_21054);
or U23477 (N_23477,N_21215,N_21710);
or U23478 (N_23478,N_21469,N_20793);
or U23479 (N_23479,N_20816,N_21345);
nor U23480 (N_23480,N_20735,N_20127);
or U23481 (N_23481,N_20201,N_21438);
or U23482 (N_23482,N_20339,N_21358);
nand U23483 (N_23483,N_20449,N_21974);
or U23484 (N_23484,N_21556,N_20796);
xor U23485 (N_23485,N_21726,N_21261);
and U23486 (N_23486,N_21597,N_20097);
nand U23487 (N_23487,N_20115,N_21452);
or U23488 (N_23488,N_21414,N_21007);
and U23489 (N_23489,N_20003,N_21419);
nand U23490 (N_23490,N_20705,N_20580);
nand U23491 (N_23491,N_20085,N_21190);
and U23492 (N_23492,N_20487,N_20120);
or U23493 (N_23493,N_20597,N_20150);
or U23494 (N_23494,N_21328,N_21647);
nor U23495 (N_23495,N_21943,N_20921);
nand U23496 (N_23496,N_21097,N_21815);
xor U23497 (N_23497,N_20971,N_21868);
and U23498 (N_23498,N_21572,N_21804);
and U23499 (N_23499,N_20690,N_20630);
xnor U23500 (N_23500,N_21006,N_21263);
and U23501 (N_23501,N_20664,N_21065);
xnor U23502 (N_23502,N_21182,N_20576);
and U23503 (N_23503,N_20934,N_21353);
xnor U23504 (N_23504,N_20940,N_20095);
xor U23505 (N_23505,N_21490,N_20260);
and U23506 (N_23506,N_20528,N_21202);
and U23507 (N_23507,N_21847,N_20798);
and U23508 (N_23508,N_20096,N_20599);
and U23509 (N_23509,N_21855,N_20176);
and U23510 (N_23510,N_21657,N_21146);
nand U23511 (N_23511,N_21652,N_20335);
and U23512 (N_23512,N_21933,N_20054);
and U23513 (N_23513,N_20318,N_21707);
and U23514 (N_23514,N_21627,N_20942);
nand U23515 (N_23515,N_20788,N_21277);
nor U23516 (N_23516,N_20860,N_21769);
nand U23517 (N_23517,N_20138,N_20939);
and U23518 (N_23518,N_21316,N_21578);
nand U23519 (N_23519,N_20736,N_20776);
nor U23520 (N_23520,N_20828,N_20983);
xor U23521 (N_23521,N_21833,N_21411);
nor U23522 (N_23522,N_21785,N_20543);
xor U23523 (N_23523,N_21686,N_20299);
nor U23524 (N_23524,N_20807,N_20549);
or U23525 (N_23525,N_20256,N_21974);
xnor U23526 (N_23526,N_20414,N_20394);
or U23527 (N_23527,N_21110,N_21233);
or U23528 (N_23528,N_21244,N_21909);
or U23529 (N_23529,N_21271,N_21002);
and U23530 (N_23530,N_21754,N_20466);
and U23531 (N_23531,N_21804,N_21459);
and U23532 (N_23532,N_21280,N_21633);
or U23533 (N_23533,N_21522,N_21305);
xnor U23534 (N_23534,N_20893,N_20978);
xor U23535 (N_23535,N_21892,N_21107);
nor U23536 (N_23536,N_21863,N_21430);
nor U23537 (N_23537,N_21606,N_20865);
and U23538 (N_23538,N_20936,N_21551);
xnor U23539 (N_23539,N_21591,N_20424);
or U23540 (N_23540,N_20778,N_21859);
nor U23541 (N_23541,N_21149,N_21105);
nand U23542 (N_23542,N_21846,N_20999);
xnor U23543 (N_23543,N_20863,N_21110);
nor U23544 (N_23544,N_21633,N_20811);
nor U23545 (N_23545,N_21464,N_21488);
or U23546 (N_23546,N_21134,N_21393);
nor U23547 (N_23547,N_21466,N_20676);
nor U23548 (N_23548,N_21394,N_20918);
nor U23549 (N_23549,N_21836,N_20717);
and U23550 (N_23550,N_21148,N_20636);
nand U23551 (N_23551,N_20442,N_20523);
and U23552 (N_23552,N_20032,N_20256);
nand U23553 (N_23553,N_20429,N_20168);
or U23554 (N_23554,N_20748,N_21035);
xnor U23555 (N_23555,N_20828,N_21599);
xnor U23556 (N_23556,N_20639,N_20401);
nand U23557 (N_23557,N_21808,N_20719);
xor U23558 (N_23558,N_20683,N_20622);
nor U23559 (N_23559,N_20319,N_21869);
and U23560 (N_23560,N_20742,N_21932);
and U23561 (N_23561,N_20302,N_20012);
nand U23562 (N_23562,N_21300,N_21682);
nor U23563 (N_23563,N_20623,N_20992);
or U23564 (N_23564,N_21071,N_20410);
and U23565 (N_23565,N_20923,N_21628);
nand U23566 (N_23566,N_21310,N_20665);
and U23567 (N_23567,N_20035,N_21979);
nand U23568 (N_23568,N_20778,N_21112);
xnor U23569 (N_23569,N_20292,N_21013);
nor U23570 (N_23570,N_20879,N_21560);
nor U23571 (N_23571,N_21368,N_21583);
and U23572 (N_23572,N_20248,N_20354);
nor U23573 (N_23573,N_20348,N_20739);
xnor U23574 (N_23574,N_21747,N_21425);
and U23575 (N_23575,N_20171,N_21885);
or U23576 (N_23576,N_21870,N_20380);
and U23577 (N_23577,N_21370,N_20106);
xnor U23578 (N_23578,N_21828,N_21802);
or U23579 (N_23579,N_21771,N_21931);
or U23580 (N_23580,N_20431,N_21610);
nand U23581 (N_23581,N_21773,N_20064);
and U23582 (N_23582,N_20863,N_21789);
or U23583 (N_23583,N_20560,N_21552);
xnor U23584 (N_23584,N_21269,N_20793);
and U23585 (N_23585,N_20998,N_20374);
nand U23586 (N_23586,N_20164,N_21124);
nor U23587 (N_23587,N_21352,N_20192);
nand U23588 (N_23588,N_20924,N_20719);
xnor U23589 (N_23589,N_21041,N_21791);
nand U23590 (N_23590,N_21259,N_20903);
nand U23591 (N_23591,N_20905,N_21431);
or U23592 (N_23592,N_20966,N_21422);
or U23593 (N_23593,N_20219,N_20571);
xnor U23594 (N_23594,N_21351,N_21626);
or U23595 (N_23595,N_20758,N_20420);
xnor U23596 (N_23596,N_21372,N_20646);
xor U23597 (N_23597,N_21596,N_21704);
or U23598 (N_23598,N_21813,N_20907);
nand U23599 (N_23599,N_20106,N_21680);
and U23600 (N_23600,N_20468,N_21865);
nor U23601 (N_23601,N_21473,N_20505);
or U23602 (N_23602,N_20638,N_20615);
nor U23603 (N_23603,N_20041,N_20476);
nor U23604 (N_23604,N_20270,N_20726);
nor U23605 (N_23605,N_20759,N_20084);
and U23606 (N_23606,N_21435,N_20749);
or U23607 (N_23607,N_20145,N_20885);
nand U23608 (N_23608,N_21530,N_21620);
nor U23609 (N_23609,N_20009,N_21317);
nand U23610 (N_23610,N_21167,N_21794);
nand U23611 (N_23611,N_21452,N_20442);
nor U23612 (N_23612,N_21978,N_20163);
or U23613 (N_23613,N_21475,N_21517);
nor U23614 (N_23614,N_21367,N_20952);
or U23615 (N_23615,N_20588,N_20671);
and U23616 (N_23616,N_20279,N_20077);
nor U23617 (N_23617,N_21177,N_20949);
nand U23618 (N_23618,N_21386,N_20436);
xor U23619 (N_23619,N_21837,N_21596);
nand U23620 (N_23620,N_20869,N_20419);
nor U23621 (N_23621,N_20703,N_21778);
nand U23622 (N_23622,N_21136,N_21313);
or U23623 (N_23623,N_21742,N_21015);
nand U23624 (N_23624,N_20477,N_20284);
and U23625 (N_23625,N_21981,N_20060);
or U23626 (N_23626,N_21131,N_20002);
and U23627 (N_23627,N_20940,N_21531);
or U23628 (N_23628,N_20545,N_20587);
nand U23629 (N_23629,N_20920,N_21817);
nor U23630 (N_23630,N_21667,N_21002);
xor U23631 (N_23631,N_21374,N_21373);
nor U23632 (N_23632,N_21682,N_20283);
nand U23633 (N_23633,N_21594,N_21147);
nand U23634 (N_23634,N_21985,N_21967);
or U23635 (N_23635,N_21540,N_20669);
nand U23636 (N_23636,N_21984,N_21106);
and U23637 (N_23637,N_20062,N_20870);
nand U23638 (N_23638,N_21160,N_21607);
nor U23639 (N_23639,N_21384,N_20719);
nand U23640 (N_23640,N_20932,N_21529);
xnor U23641 (N_23641,N_21150,N_21056);
and U23642 (N_23642,N_20347,N_21674);
nor U23643 (N_23643,N_20339,N_21179);
and U23644 (N_23644,N_21406,N_21158);
nor U23645 (N_23645,N_20931,N_21609);
nand U23646 (N_23646,N_20485,N_20743);
nand U23647 (N_23647,N_21250,N_20615);
or U23648 (N_23648,N_20893,N_21388);
nor U23649 (N_23649,N_21349,N_20371);
nand U23650 (N_23650,N_21903,N_21828);
nand U23651 (N_23651,N_20082,N_21337);
nor U23652 (N_23652,N_21224,N_20675);
nand U23653 (N_23653,N_21057,N_21536);
nor U23654 (N_23654,N_21188,N_20451);
and U23655 (N_23655,N_20305,N_21174);
nand U23656 (N_23656,N_21392,N_21195);
and U23657 (N_23657,N_20600,N_21425);
nand U23658 (N_23658,N_21952,N_21409);
and U23659 (N_23659,N_20858,N_21454);
or U23660 (N_23660,N_20388,N_21913);
xor U23661 (N_23661,N_20067,N_21443);
nand U23662 (N_23662,N_21669,N_21564);
and U23663 (N_23663,N_21546,N_20949);
and U23664 (N_23664,N_20541,N_20004);
nor U23665 (N_23665,N_20182,N_20721);
xor U23666 (N_23666,N_20359,N_21911);
and U23667 (N_23667,N_20265,N_20981);
and U23668 (N_23668,N_21306,N_21914);
nor U23669 (N_23669,N_20638,N_21278);
nor U23670 (N_23670,N_20422,N_20125);
and U23671 (N_23671,N_20998,N_20973);
nand U23672 (N_23672,N_21131,N_21239);
or U23673 (N_23673,N_20436,N_21701);
nor U23674 (N_23674,N_21304,N_21843);
and U23675 (N_23675,N_20807,N_20778);
and U23676 (N_23676,N_20874,N_20045);
xor U23677 (N_23677,N_20207,N_21333);
nor U23678 (N_23678,N_20543,N_21198);
nand U23679 (N_23679,N_21094,N_21917);
nand U23680 (N_23680,N_20977,N_20859);
nor U23681 (N_23681,N_20310,N_20081);
and U23682 (N_23682,N_20978,N_21221);
nor U23683 (N_23683,N_20410,N_21948);
or U23684 (N_23684,N_21610,N_20997);
xor U23685 (N_23685,N_21049,N_20843);
xor U23686 (N_23686,N_20082,N_20606);
and U23687 (N_23687,N_21349,N_20039);
nand U23688 (N_23688,N_21828,N_20449);
nor U23689 (N_23689,N_21241,N_21225);
nand U23690 (N_23690,N_21012,N_21028);
xor U23691 (N_23691,N_21986,N_20391);
and U23692 (N_23692,N_20374,N_21212);
and U23693 (N_23693,N_20761,N_21080);
or U23694 (N_23694,N_20584,N_21625);
or U23695 (N_23695,N_20990,N_20340);
and U23696 (N_23696,N_20194,N_21875);
xnor U23697 (N_23697,N_20989,N_21091);
nand U23698 (N_23698,N_21664,N_20689);
or U23699 (N_23699,N_20061,N_20886);
or U23700 (N_23700,N_21549,N_20406);
and U23701 (N_23701,N_21152,N_20708);
xor U23702 (N_23702,N_21735,N_20160);
nand U23703 (N_23703,N_21314,N_21907);
nand U23704 (N_23704,N_21707,N_21004);
and U23705 (N_23705,N_20862,N_21849);
xor U23706 (N_23706,N_20213,N_21088);
nor U23707 (N_23707,N_20654,N_21530);
xnor U23708 (N_23708,N_20439,N_21315);
and U23709 (N_23709,N_20583,N_20698);
nand U23710 (N_23710,N_21706,N_20390);
xor U23711 (N_23711,N_20769,N_20639);
and U23712 (N_23712,N_20586,N_20237);
nand U23713 (N_23713,N_20808,N_21565);
and U23714 (N_23714,N_21186,N_20706);
xor U23715 (N_23715,N_20965,N_20696);
xor U23716 (N_23716,N_20726,N_21426);
nand U23717 (N_23717,N_20953,N_21145);
xor U23718 (N_23718,N_21860,N_20900);
or U23719 (N_23719,N_20989,N_20056);
or U23720 (N_23720,N_20934,N_21264);
nor U23721 (N_23721,N_21089,N_20229);
nand U23722 (N_23722,N_20283,N_20021);
nand U23723 (N_23723,N_21235,N_21709);
and U23724 (N_23724,N_20437,N_21776);
xnor U23725 (N_23725,N_20348,N_21617);
and U23726 (N_23726,N_20400,N_20409);
xor U23727 (N_23727,N_20753,N_21145);
or U23728 (N_23728,N_20322,N_21354);
and U23729 (N_23729,N_20987,N_21481);
or U23730 (N_23730,N_21264,N_20129);
or U23731 (N_23731,N_21381,N_20506);
or U23732 (N_23732,N_20565,N_20894);
and U23733 (N_23733,N_20693,N_20694);
xnor U23734 (N_23734,N_21764,N_21347);
nor U23735 (N_23735,N_20276,N_20595);
nor U23736 (N_23736,N_21768,N_21902);
and U23737 (N_23737,N_20316,N_21344);
or U23738 (N_23738,N_20483,N_21042);
or U23739 (N_23739,N_20144,N_21998);
xor U23740 (N_23740,N_20371,N_21559);
nand U23741 (N_23741,N_20762,N_21739);
and U23742 (N_23742,N_21046,N_20048);
xnor U23743 (N_23743,N_21120,N_21152);
and U23744 (N_23744,N_20872,N_20710);
and U23745 (N_23745,N_20409,N_21353);
or U23746 (N_23746,N_21222,N_21494);
and U23747 (N_23747,N_20233,N_20438);
nor U23748 (N_23748,N_20099,N_20062);
xnor U23749 (N_23749,N_21841,N_20133);
and U23750 (N_23750,N_21216,N_20811);
xor U23751 (N_23751,N_20587,N_21068);
nor U23752 (N_23752,N_20991,N_21183);
nor U23753 (N_23753,N_20514,N_21481);
nand U23754 (N_23754,N_20138,N_21554);
xnor U23755 (N_23755,N_20343,N_20778);
nor U23756 (N_23756,N_21353,N_21531);
and U23757 (N_23757,N_21049,N_20658);
nor U23758 (N_23758,N_20156,N_21738);
and U23759 (N_23759,N_20648,N_21326);
and U23760 (N_23760,N_20216,N_20592);
nand U23761 (N_23761,N_20877,N_21813);
nand U23762 (N_23762,N_21840,N_21938);
or U23763 (N_23763,N_21186,N_20361);
and U23764 (N_23764,N_21590,N_20448);
and U23765 (N_23765,N_21312,N_20051);
xor U23766 (N_23766,N_21774,N_20089);
xor U23767 (N_23767,N_21292,N_20056);
nor U23768 (N_23768,N_21916,N_21841);
nor U23769 (N_23769,N_21689,N_21204);
or U23770 (N_23770,N_20297,N_21458);
and U23771 (N_23771,N_20960,N_20275);
xnor U23772 (N_23772,N_21385,N_20131);
nand U23773 (N_23773,N_21534,N_21986);
or U23774 (N_23774,N_20419,N_20609);
nand U23775 (N_23775,N_21610,N_21974);
and U23776 (N_23776,N_21449,N_20196);
nand U23777 (N_23777,N_21017,N_20778);
nand U23778 (N_23778,N_21936,N_21397);
nand U23779 (N_23779,N_21141,N_21599);
or U23780 (N_23780,N_20258,N_21865);
nor U23781 (N_23781,N_20929,N_21205);
nand U23782 (N_23782,N_21161,N_20153);
and U23783 (N_23783,N_20294,N_21797);
or U23784 (N_23784,N_20017,N_20751);
xor U23785 (N_23785,N_21224,N_20756);
nor U23786 (N_23786,N_20974,N_21615);
nand U23787 (N_23787,N_21902,N_21640);
nand U23788 (N_23788,N_20403,N_20318);
xor U23789 (N_23789,N_20567,N_20787);
and U23790 (N_23790,N_21642,N_21168);
nand U23791 (N_23791,N_21112,N_20590);
and U23792 (N_23792,N_20923,N_20753);
nand U23793 (N_23793,N_21221,N_20719);
and U23794 (N_23794,N_21067,N_20724);
and U23795 (N_23795,N_20258,N_21052);
or U23796 (N_23796,N_21750,N_21393);
xor U23797 (N_23797,N_20848,N_20032);
nor U23798 (N_23798,N_20193,N_21312);
nand U23799 (N_23799,N_21530,N_20543);
or U23800 (N_23800,N_20595,N_20949);
nor U23801 (N_23801,N_20502,N_20462);
nor U23802 (N_23802,N_20081,N_21198);
or U23803 (N_23803,N_20109,N_20896);
and U23804 (N_23804,N_21055,N_20248);
or U23805 (N_23805,N_20902,N_20112);
nand U23806 (N_23806,N_20131,N_21752);
or U23807 (N_23807,N_20667,N_21590);
nand U23808 (N_23808,N_20592,N_21567);
and U23809 (N_23809,N_21947,N_20302);
or U23810 (N_23810,N_20415,N_21382);
nor U23811 (N_23811,N_20326,N_20642);
nor U23812 (N_23812,N_20230,N_20705);
xor U23813 (N_23813,N_21891,N_21080);
xor U23814 (N_23814,N_20029,N_20256);
nand U23815 (N_23815,N_20527,N_21920);
or U23816 (N_23816,N_20212,N_20882);
and U23817 (N_23817,N_21306,N_21661);
or U23818 (N_23818,N_20957,N_21083);
and U23819 (N_23819,N_21460,N_21604);
nor U23820 (N_23820,N_20014,N_21776);
nor U23821 (N_23821,N_20704,N_20888);
nand U23822 (N_23822,N_20654,N_20584);
xor U23823 (N_23823,N_20023,N_20965);
or U23824 (N_23824,N_21710,N_20146);
nor U23825 (N_23825,N_21328,N_20491);
nor U23826 (N_23826,N_20170,N_20949);
xnor U23827 (N_23827,N_20332,N_20267);
and U23828 (N_23828,N_20571,N_21714);
or U23829 (N_23829,N_20981,N_21029);
or U23830 (N_23830,N_21919,N_21569);
xor U23831 (N_23831,N_20554,N_20512);
and U23832 (N_23832,N_20016,N_20136);
and U23833 (N_23833,N_21386,N_21151);
xnor U23834 (N_23834,N_20665,N_21468);
and U23835 (N_23835,N_21107,N_20324);
xnor U23836 (N_23836,N_21883,N_20572);
and U23837 (N_23837,N_21320,N_21171);
nand U23838 (N_23838,N_21840,N_20880);
xnor U23839 (N_23839,N_20925,N_20574);
and U23840 (N_23840,N_20717,N_20607);
nand U23841 (N_23841,N_21890,N_20657);
nor U23842 (N_23842,N_20175,N_20942);
xnor U23843 (N_23843,N_21548,N_21946);
and U23844 (N_23844,N_20374,N_21801);
or U23845 (N_23845,N_21024,N_21853);
and U23846 (N_23846,N_20244,N_21417);
and U23847 (N_23847,N_20967,N_21109);
xor U23848 (N_23848,N_20867,N_21185);
nand U23849 (N_23849,N_20262,N_21789);
nand U23850 (N_23850,N_21614,N_21388);
and U23851 (N_23851,N_20849,N_20050);
nor U23852 (N_23852,N_20844,N_20816);
or U23853 (N_23853,N_21157,N_20310);
xnor U23854 (N_23854,N_21663,N_20063);
xor U23855 (N_23855,N_20495,N_21700);
nand U23856 (N_23856,N_20436,N_21546);
and U23857 (N_23857,N_20129,N_21288);
nor U23858 (N_23858,N_21158,N_20780);
and U23859 (N_23859,N_21596,N_21350);
or U23860 (N_23860,N_20316,N_21484);
and U23861 (N_23861,N_21084,N_21987);
nor U23862 (N_23862,N_20992,N_20940);
nand U23863 (N_23863,N_20632,N_21914);
nor U23864 (N_23864,N_20190,N_21843);
nand U23865 (N_23865,N_21809,N_21810);
xnor U23866 (N_23866,N_20890,N_20084);
or U23867 (N_23867,N_21856,N_21719);
and U23868 (N_23868,N_21563,N_21236);
or U23869 (N_23869,N_21348,N_21923);
and U23870 (N_23870,N_21201,N_21940);
and U23871 (N_23871,N_20145,N_21960);
or U23872 (N_23872,N_21681,N_20221);
or U23873 (N_23873,N_20548,N_21176);
or U23874 (N_23874,N_21681,N_21193);
and U23875 (N_23875,N_20126,N_20320);
nor U23876 (N_23876,N_20181,N_20001);
nor U23877 (N_23877,N_21419,N_21035);
nor U23878 (N_23878,N_21825,N_20404);
or U23879 (N_23879,N_21416,N_21873);
nand U23880 (N_23880,N_20167,N_20510);
xor U23881 (N_23881,N_21310,N_20598);
or U23882 (N_23882,N_21875,N_20786);
nor U23883 (N_23883,N_21137,N_21901);
or U23884 (N_23884,N_21036,N_20542);
and U23885 (N_23885,N_21755,N_20281);
nand U23886 (N_23886,N_21282,N_21807);
or U23887 (N_23887,N_20429,N_21195);
nor U23888 (N_23888,N_21506,N_21546);
and U23889 (N_23889,N_20882,N_20256);
nand U23890 (N_23890,N_21741,N_20140);
nor U23891 (N_23891,N_21046,N_21714);
nand U23892 (N_23892,N_20101,N_20936);
nand U23893 (N_23893,N_21741,N_20946);
nand U23894 (N_23894,N_21175,N_20966);
nand U23895 (N_23895,N_21566,N_21920);
nand U23896 (N_23896,N_21444,N_21172);
nand U23897 (N_23897,N_21466,N_20009);
nand U23898 (N_23898,N_21284,N_20484);
nor U23899 (N_23899,N_21092,N_20035);
and U23900 (N_23900,N_21250,N_21679);
nand U23901 (N_23901,N_20318,N_20799);
nand U23902 (N_23902,N_20591,N_21956);
nand U23903 (N_23903,N_21005,N_20313);
nor U23904 (N_23904,N_20162,N_21877);
xnor U23905 (N_23905,N_21007,N_21716);
and U23906 (N_23906,N_20000,N_20474);
nor U23907 (N_23907,N_20961,N_21897);
nand U23908 (N_23908,N_20891,N_20643);
xor U23909 (N_23909,N_21999,N_20497);
xnor U23910 (N_23910,N_21543,N_20942);
nor U23911 (N_23911,N_20839,N_21805);
nand U23912 (N_23912,N_21539,N_20474);
and U23913 (N_23913,N_21656,N_21607);
nand U23914 (N_23914,N_21079,N_21101);
nand U23915 (N_23915,N_21144,N_21466);
nand U23916 (N_23916,N_21638,N_20055);
or U23917 (N_23917,N_20596,N_20094);
nand U23918 (N_23918,N_21409,N_20598);
or U23919 (N_23919,N_20681,N_21651);
and U23920 (N_23920,N_21807,N_21456);
xnor U23921 (N_23921,N_20410,N_21540);
xor U23922 (N_23922,N_20732,N_21291);
and U23923 (N_23923,N_21054,N_20320);
and U23924 (N_23924,N_20556,N_20774);
or U23925 (N_23925,N_21179,N_20113);
xor U23926 (N_23926,N_20762,N_20352);
or U23927 (N_23927,N_21177,N_20574);
xor U23928 (N_23928,N_20240,N_21238);
xor U23929 (N_23929,N_20447,N_20585);
and U23930 (N_23930,N_20793,N_20206);
nor U23931 (N_23931,N_21989,N_21024);
nor U23932 (N_23932,N_20582,N_21129);
nand U23933 (N_23933,N_20696,N_20529);
and U23934 (N_23934,N_21144,N_20377);
and U23935 (N_23935,N_20029,N_21106);
and U23936 (N_23936,N_20319,N_20540);
or U23937 (N_23937,N_20825,N_21018);
nor U23938 (N_23938,N_21838,N_20393);
xor U23939 (N_23939,N_21352,N_21051);
or U23940 (N_23940,N_20564,N_20604);
and U23941 (N_23941,N_21675,N_21766);
or U23942 (N_23942,N_20834,N_21734);
xnor U23943 (N_23943,N_21900,N_21330);
and U23944 (N_23944,N_21957,N_21505);
xnor U23945 (N_23945,N_20456,N_21361);
nand U23946 (N_23946,N_20376,N_20280);
and U23947 (N_23947,N_21471,N_21299);
xor U23948 (N_23948,N_21344,N_20233);
nand U23949 (N_23949,N_21398,N_20191);
nor U23950 (N_23950,N_20618,N_20263);
nor U23951 (N_23951,N_20814,N_21979);
nor U23952 (N_23952,N_21578,N_20413);
xnor U23953 (N_23953,N_20927,N_20603);
and U23954 (N_23954,N_20537,N_20652);
and U23955 (N_23955,N_21404,N_21707);
nand U23956 (N_23956,N_20931,N_20226);
nor U23957 (N_23957,N_20910,N_21046);
nor U23958 (N_23958,N_21304,N_21603);
xnor U23959 (N_23959,N_20232,N_20882);
nand U23960 (N_23960,N_21095,N_21273);
nor U23961 (N_23961,N_21610,N_20852);
or U23962 (N_23962,N_21785,N_21866);
nor U23963 (N_23963,N_20586,N_20771);
xnor U23964 (N_23964,N_21169,N_21683);
or U23965 (N_23965,N_20094,N_21972);
nand U23966 (N_23966,N_20986,N_21879);
and U23967 (N_23967,N_20164,N_20435);
or U23968 (N_23968,N_21465,N_21603);
nor U23969 (N_23969,N_21900,N_20013);
and U23970 (N_23970,N_20453,N_20401);
xor U23971 (N_23971,N_20510,N_20939);
or U23972 (N_23972,N_20838,N_21774);
nor U23973 (N_23973,N_20348,N_21202);
xor U23974 (N_23974,N_21093,N_20292);
xor U23975 (N_23975,N_20068,N_20741);
nor U23976 (N_23976,N_21984,N_20387);
or U23977 (N_23977,N_21158,N_20098);
nand U23978 (N_23978,N_21894,N_21839);
nor U23979 (N_23979,N_21242,N_21618);
and U23980 (N_23980,N_21082,N_21720);
xnor U23981 (N_23981,N_21359,N_21882);
or U23982 (N_23982,N_21118,N_21651);
xnor U23983 (N_23983,N_21229,N_20882);
nor U23984 (N_23984,N_20555,N_21776);
nor U23985 (N_23985,N_20082,N_20324);
or U23986 (N_23986,N_21829,N_20338);
xor U23987 (N_23987,N_21843,N_20612);
nor U23988 (N_23988,N_21878,N_20843);
nand U23989 (N_23989,N_21448,N_21466);
and U23990 (N_23990,N_20509,N_21486);
nor U23991 (N_23991,N_21225,N_20302);
xor U23992 (N_23992,N_21619,N_20156);
nand U23993 (N_23993,N_20725,N_20738);
xnor U23994 (N_23994,N_20037,N_21753);
nor U23995 (N_23995,N_20065,N_21267);
nor U23996 (N_23996,N_21131,N_20074);
nand U23997 (N_23997,N_21509,N_21268);
nor U23998 (N_23998,N_20071,N_21321);
or U23999 (N_23999,N_21273,N_21422);
nor U24000 (N_24000,N_23030,N_22221);
or U24001 (N_24001,N_23168,N_22204);
or U24002 (N_24002,N_23028,N_22630);
and U24003 (N_24003,N_22326,N_22044);
or U24004 (N_24004,N_23719,N_22773);
and U24005 (N_24005,N_23761,N_22647);
nand U24006 (N_24006,N_23391,N_23058);
or U24007 (N_24007,N_23104,N_23446);
nor U24008 (N_24008,N_22369,N_22165);
nor U24009 (N_24009,N_23416,N_22840);
xnor U24010 (N_24010,N_22817,N_23949);
nand U24011 (N_24011,N_23925,N_22663);
xnor U24012 (N_24012,N_23882,N_23677);
xnor U24013 (N_24013,N_22091,N_23203);
xor U24014 (N_24014,N_23940,N_23723);
or U24015 (N_24015,N_22857,N_22998);
or U24016 (N_24016,N_22517,N_22714);
nand U24017 (N_24017,N_22427,N_22246);
and U24018 (N_24018,N_23773,N_22018);
nor U24019 (N_24019,N_22980,N_23824);
and U24020 (N_24020,N_23867,N_23418);
and U24021 (N_24021,N_23673,N_22548);
or U24022 (N_24022,N_22977,N_23669);
and U24023 (N_24023,N_22762,N_22585);
nand U24024 (N_24024,N_22890,N_22706);
nand U24025 (N_24025,N_22421,N_23860);
nand U24026 (N_24026,N_23414,N_22434);
nand U24027 (N_24027,N_22151,N_23924);
xnor U24028 (N_24028,N_23785,N_22832);
nor U24029 (N_24029,N_23731,N_23385);
nand U24030 (N_24030,N_23345,N_22925);
nand U24031 (N_24031,N_22511,N_22786);
nand U24032 (N_24032,N_23965,N_23498);
or U24033 (N_24033,N_23795,N_23307);
nand U24034 (N_24034,N_22041,N_23433);
nand U24035 (N_24035,N_22156,N_23331);
or U24036 (N_24036,N_22361,N_22464);
and U24037 (N_24037,N_22894,N_22090);
and U24038 (N_24038,N_23623,N_23614);
or U24039 (N_24039,N_23244,N_22742);
nor U24040 (N_24040,N_22653,N_23943);
and U24041 (N_24041,N_22073,N_22214);
and U24042 (N_24042,N_23080,N_22051);
xnor U24043 (N_24043,N_22268,N_23332);
and U24044 (N_24044,N_23458,N_23655);
nor U24045 (N_24045,N_23410,N_22937);
and U24046 (N_24046,N_22420,N_23143);
and U24047 (N_24047,N_22978,N_23271);
nor U24048 (N_24048,N_23703,N_22360);
or U24049 (N_24049,N_23077,N_23076);
or U24050 (N_24050,N_22061,N_22198);
or U24051 (N_24051,N_22191,N_22848);
nand U24052 (N_24052,N_22498,N_22929);
or U24053 (N_24053,N_22851,N_22605);
nand U24054 (N_24054,N_23341,N_22478);
xnor U24055 (N_24055,N_22907,N_23682);
or U24056 (N_24056,N_23147,N_23989);
xor U24057 (N_24057,N_23564,N_22744);
nor U24058 (N_24058,N_23969,N_22648);
and U24059 (N_24059,N_23031,N_22607);
nor U24060 (N_24060,N_23704,N_23960);
nand U24061 (N_24061,N_23840,N_23891);
nand U24062 (N_24062,N_23629,N_23473);
nand U24063 (N_24063,N_22599,N_23641);
nand U24064 (N_24064,N_22696,N_23634);
nand U24065 (N_24065,N_22778,N_23643);
or U24066 (N_24066,N_23217,N_22956);
or U24067 (N_24067,N_23119,N_23872);
nor U24068 (N_24068,N_22170,N_23199);
xor U24069 (N_24069,N_23585,N_22513);
and U24070 (N_24070,N_22408,N_22260);
xnor U24071 (N_24071,N_23277,N_23432);
xnor U24072 (N_24072,N_22602,N_23776);
and U24073 (N_24073,N_23409,N_22486);
xnor U24074 (N_24074,N_23532,N_23664);
nor U24075 (N_24075,N_22495,N_22070);
nor U24076 (N_24076,N_22912,N_22885);
or U24077 (N_24077,N_23695,N_22231);
nand U24078 (N_24078,N_23048,N_22333);
xnor U24079 (N_24079,N_23845,N_23308);
nor U24080 (N_24080,N_22891,N_23211);
nand U24081 (N_24081,N_22945,N_22641);
nor U24082 (N_24082,N_22645,N_22068);
and U24083 (N_24083,N_22604,N_23090);
xnor U24084 (N_24084,N_22021,N_23861);
nor U24085 (N_24085,N_23791,N_22487);
nand U24086 (N_24086,N_23648,N_23092);
nor U24087 (N_24087,N_23068,N_22757);
or U24088 (N_24088,N_23977,N_22723);
xnor U24089 (N_24089,N_22780,N_23393);
or U24090 (N_24090,N_23871,N_23646);
xor U24091 (N_24091,N_22088,N_22356);
nand U24092 (N_24092,N_23610,N_22280);
nand U24093 (N_24093,N_22892,N_22127);
nor U24094 (N_24094,N_23691,N_22700);
nor U24095 (N_24095,N_23661,N_23036);
or U24096 (N_24096,N_22066,N_22277);
nor U24097 (N_24097,N_22425,N_22102);
nor U24098 (N_24098,N_22065,N_23053);
and U24099 (N_24099,N_22923,N_23841);
or U24100 (N_24100,N_22330,N_22534);
and U24101 (N_24101,N_23388,N_23477);
nand U24102 (N_24102,N_22566,N_23093);
nor U24103 (N_24103,N_22272,N_23656);
or U24104 (N_24104,N_23169,N_22947);
nor U24105 (N_24105,N_23676,N_22884);
nand U24106 (N_24106,N_22235,N_22867);
and U24107 (N_24107,N_23040,N_22397);
or U24108 (N_24108,N_23497,N_23707);
or U24109 (N_24109,N_23503,N_22676);
xnor U24110 (N_24110,N_23352,N_23120);
nand U24111 (N_24111,N_22019,N_23054);
nor U24112 (N_24112,N_22684,N_23946);
nor U24113 (N_24113,N_23400,N_23278);
and U24114 (N_24114,N_23316,N_22036);
nand U24115 (N_24115,N_23511,N_22568);
or U24116 (N_24116,N_22573,N_23770);
xnor U24117 (N_24117,N_22753,N_23567);
or U24118 (N_24118,N_22347,N_22507);
and U24119 (N_24119,N_23866,N_22512);
xnor U24120 (N_24120,N_23750,N_23320);
or U24121 (N_24121,N_23530,N_22880);
xor U24122 (N_24122,N_22270,N_22193);
or U24123 (N_24123,N_23378,N_22172);
nor U24124 (N_24124,N_23253,N_23263);
nor U24125 (N_24125,N_23550,N_23494);
or U24126 (N_24126,N_23539,N_22841);
and U24127 (N_24127,N_23995,N_23584);
xnor U24128 (N_24128,N_23173,N_22805);
or U24129 (N_24129,N_22355,N_22426);
nand U24130 (N_24130,N_22001,N_22962);
or U24131 (N_24131,N_23678,N_23789);
nor U24132 (N_24132,N_22323,N_22643);
or U24133 (N_24133,N_23113,N_23578);
nand U24134 (N_24134,N_23484,N_22847);
nor U24135 (N_24135,N_22827,N_22362);
nand U24136 (N_24136,N_22422,N_23232);
or U24137 (N_24137,N_23681,N_22358);
xnor U24138 (N_24138,N_22940,N_23210);
or U24139 (N_24139,N_22692,N_23602);
or U24140 (N_24140,N_23024,N_23601);
nor U24141 (N_24141,N_23008,N_23847);
or U24142 (N_24142,N_22881,N_22610);
nor U24143 (N_24143,N_22447,N_23073);
nor U24144 (N_24144,N_23548,N_22159);
or U24145 (N_24145,N_23241,N_23248);
nor U24146 (N_24146,N_22441,N_23094);
or U24147 (N_24147,N_23043,N_22410);
or U24148 (N_24148,N_23800,N_23716);
nor U24149 (N_24149,N_22710,N_22190);
nand U24150 (N_24150,N_23524,N_22242);
nor U24151 (N_24151,N_22083,N_23125);
nor U24152 (N_24152,N_23496,N_22154);
xnor U24153 (N_24153,N_22886,N_23038);
or U24154 (N_24154,N_23366,N_22289);
or U24155 (N_24155,N_23144,N_23504);
nand U24156 (N_24156,N_23534,N_23383);
xnor U24157 (N_24157,N_22882,N_22140);
nand U24158 (N_24158,N_23899,N_22842);
xnor U24159 (N_24159,N_23665,N_23829);
or U24160 (N_24160,N_22921,N_22717);
nand U24161 (N_24161,N_22626,N_22711);
xnor U24162 (N_24162,N_23177,N_22934);
xnor U24163 (N_24163,N_23442,N_23025);
nor U24164 (N_24164,N_22915,N_23023);
or U24165 (N_24165,N_23423,N_22265);
xor U24166 (N_24166,N_22699,N_23460);
nor U24167 (N_24167,N_23455,N_23175);
and U24168 (N_24168,N_23842,N_23285);
nor U24169 (N_24169,N_23486,N_23126);
xor U24170 (N_24170,N_23813,N_22698);
and U24171 (N_24171,N_23212,N_22839);
and U24172 (N_24172,N_22679,N_23659);
xnor U24173 (N_24173,N_23583,N_22314);
nor U24174 (N_24174,N_23022,N_23815);
nand U24175 (N_24175,N_22955,N_22729);
nand U24176 (N_24176,N_23349,N_23062);
nand U24177 (N_24177,N_22831,N_23150);
xor U24178 (N_24178,N_23868,N_23215);
and U24179 (N_24179,N_23228,N_22116);
xor U24180 (N_24180,N_22402,N_22536);
or U24181 (N_24181,N_22485,N_22126);
nand U24182 (N_24182,N_23873,N_22524);
nor U24183 (N_24183,N_22301,N_22737);
and U24184 (N_24184,N_22476,N_22549);
or U24185 (N_24185,N_23926,N_22735);
or U24186 (N_24186,N_23148,N_23754);
nor U24187 (N_24187,N_23330,N_22878);
nand U24188 (N_24188,N_23559,N_23931);
xor U24189 (N_24189,N_23766,N_22303);
and U24190 (N_24190,N_23359,N_22327);
nand U24191 (N_24191,N_22031,N_23923);
and U24192 (N_24192,N_23741,N_22097);
xnor U24193 (N_24193,N_22129,N_23507);
xnor U24194 (N_24194,N_22572,N_22959);
xor U24195 (N_24195,N_23354,N_23338);
nor U24196 (N_24196,N_23927,N_22467);
nand U24197 (N_24197,N_23980,N_23667);
xor U24198 (N_24198,N_23415,N_22379);
and U24199 (N_24199,N_22725,N_22822);
and U24200 (N_24200,N_23749,N_22057);
nand U24201 (N_24201,N_23012,N_23535);
nor U24202 (N_24202,N_22344,N_23051);
nand U24203 (N_24203,N_22466,N_22423);
xnor U24204 (N_24204,N_22244,N_23767);
xnor U24205 (N_24205,N_22695,N_23123);
nand U24206 (N_24206,N_22730,N_22689);
or U24207 (N_24207,N_22559,N_23017);
or U24208 (N_24208,N_22285,N_23326);
and U24209 (N_24209,N_23945,N_22519);
and U24210 (N_24210,N_23586,N_22975);
and U24211 (N_24211,N_23774,N_23260);
xnor U24212 (N_24212,N_22670,N_22877);
xor U24213 (N_24213,N_23440,N_22888);
or U24214 (N_24214,N_23961,N_23171);
nand U24215 (N_24215,N_22400,N_22815);
or U24216 (N_24216,N_22042,N_23258);
and U24217 (N_24217,N_22320,N_23334);
and U24218 (N_24218,N_22110,N_22691);
and U24219 (N_24219,N_22781,N_22401);
and U24220 (N_24220,N_22681,N_22286);
xnor U24221 (N_24221,N_22720,N_22500);
nor U24222 (N_24222,N_22058,N_22721);
nand U24223 (N_24223,N_22652,N_22248);
xor U24224 (N_24224,N_23371,N_22835);
or U24225 (N_24225,N_23450,N_22859);
and U24226 (N_24226,N_23527,N_22206);
and U24227 (N_24227,N_22098,N_22953);
nor U24228 (N_24228,N_23981,N_23856);
xor U24229 (N_24229,N_23097,N_23552);
nor U24230 (N_24230,N_23417,N_22112);
nor U24231 (N_24231,N_23389,N_23172);
nand U24232 (N_24232,N_23708,N_22943);
xor U24233 (N_24233,N_22203,N_23060);
nand U24234 (N_24234,N_22176,N_23930);
xor U24235 (N_24235,N_23010,N_22919);
and U24236 (N_24236,N_22726,N_22171);
or U24237 (N_24237,N_23321,N_23255);
nand U24238 (N_24238,N_23102,N_23745);
and U24239 (N_24239,N_23597,N_22571);
and U24240 (N_24240,N_22146,N_23674);
and U24241 (N_24241,N_22480,N_23457);
nor U24242 (N_24242,N_23002,N_23663);
and U24243 (N_24243,N_23499,N_22124);
nand U24244 (N_24244,N_23361,N_22869);
xor U24245 (N_24245,N_23465,N_23701);
nor U24246 (N_24246,N_23122,N_23908);
or U24247 (N_24247,N_23650,N_23974);
and U24248 (N_24248,N_23651,N_23500);
or U24249 (N_24249,N_23760,N_23765);
or U24250 (N_24250,N_22690,N_22678);
and U24251 (N_24251,N_23950,N_23686);
nand U24252 (N_24252,N_22037,N_22905);
nor U24253 (N_24253,N_22521,N_23236);
nor U24254 (N_24254,N_22939,N_23342);
xor U24255 (N_24255,N_22284,N_22821);
xnor U24256 (N_24256,N_22768,N_22409);
or U24257 (N_24257,N_23549,N_23600);
nand U24258 (N_24258,N_22387,N_23830);
nand U24259 (N_24259,N_23219,N_22814);
nand U24260 (N_24260,N_23518,N_23447);
or U24261 (N_24261,N_22025,N_22252);
nor U24262 (N_24262,N_23603,N_22618);
nor U24263 (N_24263,N_23702,N_23374);
nor U24264 (N_24264,N_22642,N_22331);
or U24265 (N_24265,N_23859,N_22812);
and U24266 (N_24266,N_22688,N_22461);
nor U24267 (N_24267,N_23807,N_22846);
and U24268 (N_24268,N_23521,N_23713);
xnor U24269 (N_24269,N_22577,N_22639);
or U24270 (N_24270,N_23660,N_22899);
or U24271 (N_24271,N_23902,N_22381);
xnor U24272 (N_24272,N_22094,N_23968);
and U24273 (N_24273,N_22290,N_23613);
nor U24274 (N_24274,N_22095,N_22810);
nor U24275 (N_24275,N_22796,N_22697);
and U24276 (N_24276,N_22357,N_23174);
xnor U24277 (N_24277,N_23343,N_23289);
nand U24278 (N_24278,N_23114,N_23495);
and U24279 (N_24279,N_22555,N_23957);
nor U24280 (N_24280,N_22342,N_23846);
xnor U24281 (N_24281,N_22311,N_22174);
nand U24282 (N_24282,N_22654,N_22067);
or U24283 (N_24283,N_23734,N_23061);
and U24284 (N_24284,N_23194,N_22764);
nor U24285 (N_24285,N_23652,N_23089);
nand U24286 (N_24286,N_23441,N_22579);
or U24287 (N_24287,N_22393,N_23594);
and U24288 (N_24288,N_23149,N_23922);
and U24289 (N_24289,N_23710,N_23287);
nand U24290 (N_24290,N_23408,N_23117);
xor U24291 (N_24291,N_22125,N_22103);
nand U24292 (N_24292,N_23933,N_23261);
nand U24293 (N_24293,N_22704,N_22924);
nand U24294 (N_24294,N_23555,N_22554);
and U24295 (N_24295,N_23112,N_23376);
xor U24296 (N_24296,N_23300,N_22801);
and U24297 (N_24297,N_23124,N_23347);
nor U24298 (N_24298,N_22218,N_23565);
or U24299 (N_24299,N_23170,N_22510);
xnor U24300 (N_24300,N_23640,N_23833);
nand U24301 (N_24301,N_23537,N_22034);
xnor U24302 (N_24302,N_22489,N_23176);
or U24303 (N_24303,N_23242,N_22685);
nand U24304 (N_24304,N_23733,N_22373);
or U24305 (N_24305,N_22366,N_23201);
nor U24306 (N_24306,N_23853,N_23921);
xnor U24307 (N_24307,N_23154,N_22300);
nor U24308 (N_24308,N_23070,N_22234);
and U24309 (N_24309,N_23454,N_23317);
and U24310 (N_24310,N_22603,N_22414);
nand U24311 (N_24311,N_23786,N_22199);
nor U24312 (N_24312,N_22296,N_22050);
and U24313 (N_24313,N_22747,N_23592);
nor U24314 (N_24314,N_23195,N_23875);
or U24315 (N_24315,N_23540,N_23998);
and U24316 (N_24316,N_22315,N_23720);
or U24317 (N_24317,N_23898,N_22520);
or U24318 (N_24318,N_22281,N_22115);
and U24319 (N_24319,N_23283,N_23456);
xor U24320 (N_24320,N_22637,N_23913);
and U24321 (N_24321,N_23528,N_22027);
or U24322 (N_24322,N_22732,N_23879);
nor U24323 (N_24323,N_22694,N_22537);
and U24324 (N_24324,N_23480,N_22665);
nor U24325 (N_24325,N_23306,N_22106);
nor U24326 (N_24326,N_22659,N_23762);
nand U24327 (N_24327,N_22189,N_23240);
and U24328 (N_24328,N_23746,N_23787);
nor U24329 (N_24329,N_22990,N_22826);
or U24330 (N_24330,N_22403,N_22318);
xor U24331 (N_24331,N_22553,N_23384);
nor U24332 (N_24332,N_22633,N_23368);
and U24333 (N_24333,N_23290,N_23291);
xnor U24334 (N_24334,N_23186,N_23997);
nand U24335 (N_24335,N_23139,N_23910);
nor U24336 (N_24336,N_22656,N_22005);
nor U24337 (N_24337,N_23430,N_22541);
nor U24338 (N_24338,N_23482,N_23204);
xnor U24339 (N_24339,N_22702,N_22371);
nand U24340 (N_24340,N_22121,N_23852);
nor U24341 (N_24341,N_23403,N_23336);
nor U24342 (N_24342,N_23501,N_23346);
or U24343 (N_24343,N_23658,N_23693);
nor U24344 (N_24344,N_22264,N_23009);
and U24345 (N_24345,N_22349,N_22979);
and U24346 (N_24346,N_23814,N_23560);
and U24347 (N_24347,N_22359,N_22712);
xor U24348 (N_24348,N_22635,N_22576);
xor U24349 (N_24349,N_23911,N_22531);
nand U24350 (N_24350,N_22895,N_22650);
or U24351 (N_24351,N_23404,N_23579);
or U24352 (N_24352,N_23647,N_22946);
nor U24353 (N_24353,N_22328,N_23066);
xnor U24354 (N_24354,N_23914,N_23188);
xnor U24355 (N_24355,N_23865,N_23425);
xnor U24356 (N_24356,N_22767,N_23675);
or U24357 (N_24357,N_22207,N_23302);
nor U24358 (N_24358,N_23226,N_23018);
and U24359 (N_24359,N_23576,N_22453);
or U24360 (N_24360,N_22514,N_23580);
or U24361 (N_24361,N_23901,N_22039);
xnor U24362 (N_24362,N_23363,N_23880);
xor U24363 (N_24363,N_22936,N_23282);
xor U24364 (N_24364,N_22388,N_22854);
or U24365 (N_24365,N_22343,N_22307);
nand U24366 (N_24366,N_22621,N_22855);
nand U24367 (N_24367,N_22166,N_22139);
nor U24368 (N_24368,N_23355,N_22623);
or U24369 (N_24369,N_23137,N_23607);
nand U24370 (N_24370,N_23305,N_22384);
or U24371 (N_24371,N_22734,N_23075);
or U24372 (N_24372,N_23615,N_23959);
or U24373 (N_24373,N_22535,N_22321);
xnor U24374 (N_24374,N_23420,N_22078);
or U24375 (N_24375,N_23625,N_22561);
or U24376 (N_24376,N_22370,N_23488);
nand U24377 (N_24377,N_23869,N_22263);
and U24378 (N_24378,N_23015,N_22988);
or U24379 (N_24379,N_22266,N_23966);
nand U24380 (N_24380,N_22111,N_23319);
or U24381 (N_24381,N_23805,N_22064);
nand U24382 (N_24382,N_22597,N_22294);
or U24383 (N_24383,N_23325,N_23111);
nand U24384 (N_24384,N_22392,N_22523);
xnor U24385 (N_24385,N_22475,N_23755);
xnor U24386 (N_24386,N_22123,N_22844);
xor U24387 (N_24387,N_22047,N_23728);
xnor U24388 (N_24388,N_23471,N_22611);
nor U24389 (N_24389,N_22829,N_22999);
or U24390 (N_24390,N_23545,N_22122);
and U24391 (N_24391,N_22014,N_23134);
nor U24392 (N_24392,N_23929,N_22933);
and U24393 (N_24393,N_23461,N_22227);
xor U24394 (N_24394,N_23777,N_23042);
nor U24395 (N_24395,N_23803,N_22589);
or U24396 (N_24396,N_23724,N_23078);
xnor U24397 (N_24397,N_23680,N_22614);
or U24398 (N_24398,N_22966,N_23905);
nor U24399 (N_24399,N_22440,N_23907);
or U24400 (N_24400,N_23470,N_23313);
xor U24401 (N_24401,N_22063,N_22911);
and U24402 (N_24402,N_23027,N_23165);
xnor U24403 (N_24403,N_22861,N_23904);
or U24404 (N_24404,N_22000,N_23864);
nand U24405 (N_24405,N_22229,N_23353);
and U24406 (N_24406,N_23294,N_22967);
nor U24407 (N_24407,N_23897,N_22790);
or U24408 (N_24408,N_23303,N_22375);
nor U24409 (N_24409,N_22926,N_23451);
xor U24410 (N_24410,N_22177,N_22913);
nor U24411 (N_24411,N_23127,N_22987);
and U24412 (N_24412,N_22662,N_23581);
nand U24413 (N_24413,N_23620,N_22395);
nor U24414 (N_24414,N_23611,N_22219);
nand U24415 (N_24415,N_22743,N_22228);
or U24416 (N_24416,N_23915,N_22687);
xor U24417 (N_24417,N_23717,N_22144);
xor U24418 (N_24418,N_23963,N_22874);
nand U24419 (N_24419,N_22631,N_22169);
or U24420 (N_24420,N_23227,N_23820);
and U24421 (N_24421,N_23573,N_23772);
and U24422 (N_24422,N_22758,N_23958);
or U24423 (N_24423,N_23844,N_22843);
xnor U24424 (N_24424,N_22096,N_22319);
nor U24425 (N_24425,N_23874,N_23155);
or U24426 (N_24426,N_22108,N_23608);
nand U24427 (N_24427,N_22615,N_23178);
or U24428 (N_24428,N_23737,N_22713);
nand U24429 (N_24429,N_23407,N_22215);
or U24430 (N_24430,N_22863,N_22033);
xnor U24431 (N_24431,N_23775,N_22223);
nor U24432 (N_24432,N_23026,N_23485);
xnor U24433 (N_24433,N_23599,N_23947);
xnor U24434 (N_24434,N_23034,N_22469);
or U24435 (N_24435,N_22794,N_23462);
or U24436 (N_24436,N_23167,N_22763);
or U24437 (N_24437,N_23509,N_23542);
or U24438 (N_24438,N_22406,N_22150);
or U24439 (N_24439,N_23574,N_23158);
nor U24440 (N_24440,N_23132,N_22114);
and U24441 (N_24441,N_22372,N_22870);
or U24442 (N_24442,N_22309,N_22750);
xor U24443 (N_24443,N_23340,N_22897);
nand U24444 (N_24444,N_23683,N_23952);
and U24445 (N_24445,N_22118,N_23293);
or U24446 (N_24446,N_23357,N_23358);
nand U24447 (N_24447,N_22993,N_22580);
or U24448 (N_24448,N_22340,N_23225);
or U24449 (N_24449,N_22952,N_22465);
nor U24450 (N_24450,N_22105,N_23084);
and U24451 (N_24451,N_23515,N_23801);
xnor U24452 (N_24452,N_22590,N_23479);
nand U24453 (N_24453,N_23711,N_22405);
nand U24454 (N_24454,N_22596,N_22569);
and U24455 (N_24455,N_23821,N_22961);
and U24456 (N_24456,N_23160,N_22162);
nand U24457 (N_24457,N_23510,N_23223);
or U24458 (N_24458,N_22501,N_22293);
xnor U24459 (N_24459,N_22992,N_22181);
nand U24460 (N_24460,N_23523,N_22378);
nor U24461 (N_24461,N_22601,N_22238);
and U24462 (N_24462,N_22527,N_22302);
xnor U24463 (N_24463,N_23329,N_22530);
nor U24464 (N_24464,N_23920,N_23207);
or U24465 (N_24465,N_22186,N_22745);
nor U24466 (N_24466,N_22738,N_22481);
nor U24467 (N_24467,N_23396,N_22138);
and U24468 (N_24468,N_22491,N_23627);
nand U24469 (N_24469,N_23292,N_23516);
and U24470 (N_24470,N_22398,N_22077);
nand U24471 (N_24471,N_23793,N_23327);
xor U24472 (N_24472,N_23973,N_22304);
nand U24473 (N_24473,N_23337,N_22438);
or U24474 (N_24474,N_23883,N_23214);
xnor U24475 (N_24475,N_23431,N_23605);
or U24476 (N_24476,N_22224,N_23279);
xor U24477 (N_24477,N_22889,N_22499);
xnor U24478 (N_24478,N_22594,N_22184);
nor U24479 (N_24479,N_22724,N_22660);
nor U24480 (N_24480,N_23729,N_23364);
nor U24481 (N_24481,N_22256,N_22205);
or U24482 (N_24482,N_23780,N_22101);
or U24483 (N_24483,N_23045,N_23505);
or U24484 (N_24484,N_23179,N_23370);
and U24485 (N_24485,N_23397,N_22325);
or U24486 (N_24486,N_23422,N_23096);
nor U24487 (N_24487,N_23115,N_23763);
nor U24488 (N_24488,N_22625,N_23453);
nor U24489 (N_24489,N_23333,N_22173);
or U24490 (N_24490,N_23863,N_22072);
nand U24491 (N_24491,N_22463,N_22871);
nor U24492 (N_24492,N_22741,N_23351);
nand U24493 (N_24493,N_22651,N_22994);
nand U24494 (N_24494,N_23100,N_22188);
or U24495 (N_24495,N_23967,N_23056);
nor U24496 (N_24496,N_23474,N_23999);
nor U24497 (N_24497,N_23138,N_22551);
xnor U24498 (N_24498,N_23624,N_22666);
nand U24499 (N_24499,N_23582,N_23163);
nor U24500 (N_24500,N_23764,N_23526);
nor U24501 (N_24501,N_23944,N_23413);
and U24502 (N_24502,N_22305,N_23032);
xnor U24503 (N_24503,N_22306,N_23621);
xor U24504 (N_24504,N_23348,N_22986);
nand U24505 (N_24505,N_23490,N_23213);
nand U24506 (N_24506,N_23088,N_22503);
or U24507 (N_24507,N_23133,N_23019);
nor U24508 (N_24508,N_23218,N_23424);
nor U24509 (N_24509,N_22969,N_23637);
or U24510 (N_24510,N_23047,N_23954);
nor U24511 (N_24511,N_22099,N_22686);
or U24512 (N_24512,N_22671,N_23399);
nand U24513 (N_24513,N_23398,N_22161);
or U24514 (N_24514,N_22069,N_22135);
and U24515 (N_24515,N_22008,N_23788);
nand U24516 (N_24516,N_22149,N_22896);
xnor U24517 (N_24517,N_22380,N_23569);
nand U24518 (N_24518,N_22930,N_23311);
nand U24519 (N_24519,N_22335,N_22505);
xor U24520 (N_24520,N_22386,N_23895);
and U24521 (N_24521,N_22194,N_23448);
xor U24522 (N_24522,N_22920,N_23046);
nand U24523 (N_24523,N_22460,N_23744);
or U24524 (N_24524,N_22071,N_23543);
nand U24525 (N_24525,N_22705,N_22799);
nand U24526 (N_24526,N_23726,N_22100);
nand U24527 (N_24527,N_22632,N_22233);
nand U24528 (N_24528,N_22365,N_23064);
and U24529 (N_24529,N_23251,N_23041);
nor U24530 (N_24530,N_22444,N_22903);
or U24531 (N_24531,N_23832,N_22901);
or U24532 (N_24532,N_22490,N_22984);
or U24533 (N_24533,N_22258,N_22298);
and U24534 (N_24534,N_22765,N_22795);
or U24535 (N_24535,N_23237,N_23221);
nor U24536 (N_24536,N_23941,N_22415);
nand U24537 (N_24537,N_23235,N_22760);
and U24538 (N_24538,N_22383,N_22991);
nand U24539 (N_24539,N_22182,N_23426);
nand U24540 (N_24540,N_22137,N_22389);
and U24541 (N_24541,N_22329,N_23381);
or U24542 (N_24542,N_22550,N_22374);
or U24543 (N_24543,N_22479,N_22497);
and U24544 (N_24544,N_23362,N_23464);
nand U24545 (N_24545,N_22002,N_22985);
nor U24546 (N_24546,N_22179,N_23268);
nand U24547 (N_24547,N_23684,N_22287);
xnor U24548 (N_24548,N_23992,N_23557);
nor U24549 (N_24549,N_23281,N_23246);
xor U24550 (N_24550,N_22838,N_23491);
nor U24551 (N_24551,N_22606,N_23003);
xor U24552 (N_24552,N_22789,N_23252);
xor U24553 (N_24553,N_22085,N_23136);
and U24554 (N_24554,N_23689,N_23739);
and U24555 (N_24555,N_22797,N_22837);
and U24556 (N_24556,N_23638,N_23135);
or U24557 (N_24557,N_22655,N_22351);
and U24558 (N_24558,N_23492,N_23753);
and U24559 (N_24559,N_23369,N_22417);
xor U24560 (N_24560,N_22046,N_23059);
and U24561 (N_24561,N_23044,N_22565);
and U24562 (N_24562,N_22017,N_22316);
nand U24563 (N_24563,N_23759,N_22168);
nor U24564 (N_24564,N_22022,N_22411);
nor U24565 (N_24565,N_23982,N_22007);
nand U24566 (N_24566,N_23668,N_23109);
or U24567 (N_24567,N_23593,N_22995);
xnor U24568 (N_24568,N_23976,N_23493);
xnor U24569 (N_24569,N_23013,N_23609);
nand U24570 (N_24570,N_22212,N_22616);
xnor U24571 (N_24571,N_23808,N_22225);
and U24572 (N_24572,N_22748,N_23315);
and U24573 (N_24573,N_23402,N_22516);
xnor U24574 (N_24574,N_23942,N_23004);
xor U24575 (N_24575,N_22086,N_22556);
nand U24576 (N_24576,N_23419,N_23747);
or U24577 (N_24577,N_23151,N_23666);
and U24578 (N_24578,N_22617,N_22131);
or U24579 (N_24579,N_22310,N_23630);
and U24580 (N_24580,N_22043,N_22820);
nor U24581 (N_24581,N_23196,N_23264);
xnor U24582 (N_24582,N_23705,N_23231);
nor U24583 (N_24583,N_22640,N_22167);
nor U24584 (N_24584,N_22437,N_23598);
nor U24585 (N_24585,N_23091,N_22250);
xnor U24586 (N_24586,N_23819,N_22964);
nand U24587 (N_24587,N_23222,N_23508);
nor U24588 (N_24588,N_22055,N_23809);
nand U24589 (N_24589,N_22627,N_23671);
nor U24590 (N_24590,N_22887,N_22251);
xor U24591 (N_24591,N_22542,N_23622);
and U24592 (N_24592,N_22211,N_23831);
xor U24593 (N_24593,N_23890,N_22377);
nor U24594 (N_24594,N_23262,N_22484);
xnor U24595 (N_24595,N_22672,N_22436);
or U24596 (N_24596,N_23103,N_22142);
nand U24597 (N_24597,N_22496,N_23878);
xnor U24598 (N_24598,N_23506,N_22079);
or U24599 (N_24599,N_22332,N_23993);
xor U24600 (N_24600,N_22574,N_22954);
xnor U24601 (N_24601,N_22728,N_23514);
or U24602 (N_24602,N_22431,N_22201);
and U24603 (N_24603,N_22949,N_23595);
and U24604 (N_24604,N_23743,N_23577);
nor U24605 (N_24605,N_23467,N_22093);
or U24606 (N_24606,N_23274,N_23888);
xor U24607 (N_24607,N_23021,N_23690);
nand U24608 (N_24608,N_22222,N_22803);
or U24609 (N_24609,N_22667,N_22241);
and U24610 (N_24610,N_22253,N_23828);
nor U24611 (N_24611,N_22493,N_22922);
xor U24612 (N_24612,N_22893,N_22011);
xor U24613 (N_24613,N_23826,N_23067);
xnor U24614 (N_24614,N_22341,N_22062);
xor U24615 (N_24615,N_23487,N_23928);
nor U24616 (N_24616,N_23522,N_23688);
and U24617 (N_24617,N_23129,N_23802);
or U24618 (N_24618,N_23591,N_22087);
xor U24619 (N_24619,N_23063,N_23551);
nand U24620 (N_24620,N_22213,N_23919);
and U24621 (N_24621,N_23257,N_23270);
nand U24622 (N_24622,N_22749,N_22824);
nor U24623 (N_24623,N_23893,N_22876);
xnor U24624 (N_24624,N_22217,N_22472);
and U24625 (N_24625,N_22825,N_23020);
nand U24626 (N_24626,N_22020,N_23118);
and U24627 (N_24627,N_22664,N_22210);
and U24628 (N_24628,N_23344,N_22708);
or U24629 (N_24629,N_23014,N_22581);
or U24630 (N_24630,N_23273,N_23057);
xnor U24631 (N_24631,N_22963,N_23373);
nand U24632 (N_24632,N_22473,N_22339);
xnor U24633 (N_24633,N_23220,N_23110);
and U24634 (N_24634,N_23538,N_22981);
and U24635 (N_24635,N_23085,N_22451);
and U24636 (N_24636,N_23851,N_23142);
xor U24637 (N_24637,N_22701,N_22739);
xnor U24638 (N_24638,N_22783,N_23481);
xnor U24639 (N_24639,N_23247,N_22983);
xnor U24640 (N_24640,N_23964,N_23463);
nor U24641 (N_24641,N_23706,N_22492);
and U24642 (N_24642,N_22030,N_22482);
xnor U24643 (N_24643,N_23699,N_23502);
nand U24644 (N_24644,N_22113,N_22872);
nor U24645 (N_24645,N_23635,N_23990);
or U24646 (N_24646,N_23339,N_23099);
xor U24647 (N_24647,N_22240,N_23185);
xnor U24648 (N_24648,N_23740,N_23131);
nor U24649 (N_24649,N_23672,N_22883);
nor U24650 (N_24650,N_23164,N_23324);
or U24651 (N_24651,N_23360,N_22026);
or U24652 (N_24652,N_22779,N_22928);
nand U24653 (N_24653,N_23616,N_22104);
and U24654 (N_24654,N_23065,N_23533);
and U24655 (N_24655,N_22367,N_23779);
nand U24656 (N_24656,N_23698,N_23401);
nand U24657 (N_24657,N_23876,N_22629);
nor U24658 (N_24658,N_22751,N_23996);
or U24659 (N_24659,N_23428,N_22348);
xor U24660 (N_24660,N_23238,N_23145);
nor U24661 (N_24661,N_22628,N_23735);
or U24662 (N_24662,N_22148,N_22529);
xnor U24663 (N_24663,N_23011,N_22680);
xnor U24664 (N_24664,N_23209,N_23645);
or U24665 (N_24665,N_23906,N_22040);
or U24666 (N_24666,N_22130,N_22028);
nand U24667 (N_24667,N_22776,N_22772);
and U24668 (N_24668,N_22132,N_23536);
nor U24669 (N_24669,N_23128,N_23180);
xor U24670 (N_24670,N_23037,N_22902);
and U24671 (N_24671,N_22752,N_23280);
or U24672 (N_24672,N_23934,N_23590);
or U24673 (N_24673,N_22382,N_22187);
nor U24674 (N_24674,N_22800,N_23757);
xnor U24675 (N_24675,N_23229,N_23654);
nor U24676 (N_24676,N_22570,N_22141);
or U24677 (N_24677,N_22914,N_22038);
nand U24678 (N_24678,N_23685,N_22592);
and U24679 (N_24679,N_23190,N_23478);
or U24680 (N_24680,N_22353,N_23367);
nor U24681 (N_24681,N_23243,N_23714);
nor U24682 (N_24682,N_23434,N_23835);
or U24683 (N_24683,N_22424,N_22435);
and U24684 (N_24684,N_22931,N_22430);
or U24685 (N_24685,N_23756,N_22539);
nand U24686 (N_24686,N_23626,N_23909);
nand U24687 (N_24687,N_23443,N_23848);
or U24688 (N_24688,N_22722,N_23520);
nor U24689 (N_24689,N_22185,N_22575);
or U24690 (N_24690,N_22013,N_23596);
or U24691 (N_24691,N_22624,N_22583);
nand U24692 (N_24692,N_22143,N_23700);
and U24693 (N_24693,N_22254,N_22898);
nand U24694 (N_24694,N_22276,N_22504);
nand U24695 (N_24695,N_22428,N_23799);
or U24696 (N_24696,N_23792,N_23105);
or U24697 (N_24697,N_23230,N_23106);
nor U24698 (N_24698,N_22334,N_22661);
or U24699 (N_24699,N_22418,N_22336);
nand U24700 (N_24700,N_23392,N_23249);
nand U24701 (N_24701,N_23953,N_22774);
or U24702 (N_24702,N_22120,N_22192);
or U24703 (N_24703,N_23216,N_22230);
nor U24704 (N_24704,N_22813,N_23452);
xnor U24705 (N_24705,N_22232,N_23130);
nand U24706 (N_24706,N_22259,N_23483);
nand U24707 (N_24707,N_22035,N_22200);
and U24708 (N_24708,N_23156,N_23429);
or U24709 (N_24709,N_22715,N_23162);
or U24710 (N_24710,N_22968,N_23439);
nand U24711 (N_24711,N_22474,N_22455);
nand U24712 (N_24712,N_22271,N_23712);
or U24713 (N_24713,N_23233,N_23049);
nand U24714 (N_24714,N_23633,N_23386);
nand U24715 (N_24715,N_22769,N_23751);
nand U24716 (N_24716,N_22004,N_23742);
nand U24717 (N_24717,N_22468,N_23644);
nand U24718 (N_24718,N_22449,N_22350);
nand U24719 (N_24719,N_22598,N_22657);
nor U24720 (N_24720,N_22649,N_22613);
or U24721 (N_24721,N_23298,N_22178);
and U24722 (N_24722,N_22419,N_23721);
xor U24723 (N_24723,N_23192,N_23696);
or U24724 (N_24724,N_22295,N_23887);
xor U24725 (N_24725,N_23855,N_23006);
nand U24726 (N_24726,N_22868,N_22288);
or U24727 (N_24727,N_22546,N_22816);
nor U24728 (N_24728,N_22771,N_22682);
nand U24729 (N_24729,N_22024,N_23295);
nor U24730 (N_24730,N_23529,N_23715);
nor U24731 (N_24731,N_23087,N_22636);
xnor U24732 (N_24732,N_22445,N_22558);
xnor U24733 (N_24733,N_22404,N_22255);
nor U24734 (N_24734,N_22442,N_23806);
nor U24735 (N_24735,N_23758,N_22588);
nor U24736 (N_24736,N_22864,N_23166);
and U24737 (N_24737,N_22376,N_22528);
nor U24738 (N_24738,N_23854,N_22756);
nor U24739 (N_24739,N_23072,N_23007);
or U24740 (N_24740,N_22782,N_22544);
and U24741 (N_24741,N_23157,N_22675);
nand U24742 (N_24742,N_23804,N_23382);
and U24743 (N_24743,N_23071,N_23513);
and U24744 (N_24744,N_23975,N_22153);
nor U24745 (N_24745,N_23208,N_22718);
or U24746 (N_24746,N_22916,N_23679);
nand U24747 (N_24747,N_23193,N_22175);
and U24748 (N_24748,N_23781,N_23748);
nor U24749 (N_24749,N_23519,N_22746);
or U24750 (N_24750,N_23894,N_22941);
and U24751 (N_24751,N_23512,N_23301);
and U24752 (N_24752,N_22875,N_23571);
nand U24753 (N_24753,N_23991,N_23849);
nor U24754 (N_24754,N_22457,N_22777);
or U24755 (N_24755,N_23069,N_22278);
nor U24756 (N_24756,N_22518,N_23489);
nor U24757 (N_24757,N_23121,N_23732);
xor U24758 (N_24758,N_22128,N_23972);
xnor U24759 (N_24759,N_23250,N_22608);
or U24760 (N_24760,N_22364,N_23870);
and U24761 (N_24761,N_23254,N_23083);
xnor U24762 (N_24762,N_22828,N_22257);
or U24763 (N_24763,N_23421,N_23286);
xnor U24764 (N_24764,N_22971,N_22502);
nand U24765 (N_24765,N_23588,N_23323);
and U24766 (N_24766,N_23769,N_23224);
xor U24767 (N_24767,N_22016,N_23438);
nand U24768 (N_24768,N_23984,N_23935);
nand U24769 (N_24769,N_22006,N_23951);
and U24770 (N_24770,N_23296,N_22092);
and U24771 (N_24771,N_22522,N_23297);
or U24772 (N_24772,N_22802,N_22818);
or U24773 (N_24773,N_22483,N_22136);
nor U24774 (N_24774,N_23568,N_23335);
or U24775 (N_24775,N_23939,N_22299);
and U24776 (N_24776,N_22560,N_23771);
and U24777 (N_24777,N_23618,N_22567);
nand U24778 (N_24778,N_23752,N_22646);
nand U24779 (N_24779,N_23039,N_22412);
or U24780 (N_24780,N_23725,N_23825);
nor U24781 (N_24781,N_23184,N_22312);
or U24782 (N_24782,N_23606,N_23778);
nand U24783 (N_24783,N_23727,N_23670);
and U24784 (N_24784,N_22784,N_22282);
xnor U24785 (N_24785,N_22237,N_23558);
or U24786 (N_24786,N_22584,N_22338);
nor U24787 (N_24787,N_23784,N_23839);
nor U24788 (N_24788,N_22830,N_22107);
nand U24789 (N_24789,N_23198,N_22736);
nor U24790 (N_24790,N_22508,N_22413);
and U24791 (N_24791,N_22798,N_23310);
nand U24792 (N_24792,N_22279,N_23052);
nand U24793 (N_24793,N_23033,N_22865);
xnor U24794 (N_24794,N_23970,N_23152);
nand U24795 (N_24795,N_22352,N_22477);
and U24796 (N_24796,N_22236,N_23572);
xor U24797 (N_24797,N_22709,N_23730);
nand U24798 (N_24798,N_23200,N_22308);
nand U24799 (N_24799,N_22819,N_23900);
nand U24800 (N_24800,N_23146,N_23153);
xor U24801 (N_24801,N_23531,N_23544);
nor U24802 (N_24802,N_22267,N_22853);
nor U24803 (N_24803,N_22850,N_23632);
xnor U24804 (N_24804,N_23275,N_23379);
nand U24805 (N_24805,N_22470,N_23468);
or U24806 (N_24806,N_22459,N_23546);
nand U24807 (N_24807,N_23736,N_23266);
xnor U24808 (N_24808,N_23709,N_22674);
nor U24809 (N_24809,N_22563,N_23639);
or U24810 (N_24810,N_23444,N_23843);
or U24811 (N_24811,N_23979,N_22164);
and U24812 (N_24812,N_22860,N_23978);
nor U24813 (N_24813,N_22337,N_23050);
or U24814 (N_24814,N_22644,N_23086);
xor U24815 (N_24815,N_23994,N_22297);
nor U24816 (N_24816,N_22049,N_23768);
xnor U24817 (N_24817,N_22906,N_22856);
or U24818 (N_24818,N_23916,N_22806);
or U24819 (N_24819,N_23653,N_22448);
or U24820 (N_24820,N_22543,N_23794);
nor U24821 (N_24821,N_23299,N_23029);
xor U24822 (N_24822,N_23016,N_23575);
nand U24823 (N_24823,N_22391,N_23267);
xor U24824 (N_24824,N_23140,N_23587);
xor U24825 (N_24825,N_23390,N_22910);
xor U24826 (N_24826,N_23896,N_22075);
or U24827 (N_24827,N_23436,N_22593);
nand U24828 (N_24828,N_22015,N_22900);
nor U24829 (N_24829,N_23541,N_23276);
nand U24830 (N_24830,N_22084,N_22620);
nor U24831 (N_24831,N_23827,N_23406);
and U24832 (N_24832,N_22494,N_22345);
or U24833 (N_24833,N_23917,N_22833);
and U24834 (N_24834,N_22454,N_23547);
and U24835 (N_24835,N_22134,N_22770);
or U24836 (N_24836,N_23850,N_22117);
nor U24837 (N_24837,N_22385,N_23427);
nand U24838 (N_24838,N_22740,N_22638);
or U24839 (N_24839,N_22243,N_23182);
nand U24840 (N_24840,N_22591,N_23375);
and U24841 (N_24841,N_23798,N_22109);
or U24842 (N_24842,N_22089,N_22788);
xor U24843 (N_24843,N_22733,N_22619);
or U24844 (N_24844,N_22958,N_22564);
and U24845 (N_24845,N_22291,N_23834);
or U24846 (N_24846,N_23936,N_23885);
nand U24847 (N_24847,N_22811,N_23811);
or U24848 (N_24848,N_23697,N_22997);
nor U24849 (N_24849,N_23191,N_22586);
nand U24850 (N_24850,N_22450,N_22390);
or U24851 (N_24851,N_23161,N_23822);
and U24852 (N_24852,N_22849,N_23141);
and U24853 (N_24853,N_23245,N_23589);
xnor U24854 (N_24854,N_22456,N_23055);
xor U24855 (N_24855,N_22269,N_22525);
or U24856 (N_24856,N_22509,N_23812);
xnor U24857 (N_24857,N_22918,N_22048);
nand U24858 (N_24858,N_22808,N_23074);
nand U24859 (N_24859,N_22488,N_22152);
and U24860 (N_24860,N_23553,N_22158);
or U24861 (N_24861,N_22582,N_22119);
and U24862 (N_24862,N_23189,N_22707);
or U24863 (N_24863,N_23466,N_22834);
and U24864 (N_24864,N_22407,N_23318);
or U24865 (N_24865,N_23817,N_22787);
xnor U24866 (N_24866,N_23862,N_23202);
and U24867 (N_24867,N_22245,N_22622);
and U24868 (N_24868,N_22540,N_22195);
nor U24869 (N_24869,N_22216,N_23356);
or U24870 (N_24870,N_22145,N_23782);
nand U24871 (N_24871,N_23256,N_22562);
and U24872 (N_24872,N_23000,N_23797);
or U24873 (N_24873,N_22273,N_22274);
or U24874 (N_24874,N_22354,N_22059);
nand U24875 (N_24875,N_23642,N_22368);
or U24876 (N_24876,N_22197,N_23082);
nor U24877 (N_24877,N_22935,N_23394);
nand U24878 (N_24878,N_23001,N_23988);
nand U24879 (N_24879,N_22970,N_22160);
or U24880 (N_24880,N_23265,N_22658);
and U24881 (N_24881,N_22080,N_23657);
and U24882 (N_24882,N_23108,N_22785);
nor U24883 (N_24883,N_22845,N_23881);
xnor U24884 (N_24884,N_22202,N_22076);
or U24885 (N_24885,N_22247,N_22673);
and U24886 (N_24886,N_22533,N_22292);
nor U24887 (N_24887,N_23932,N_23956);
and U24888 (N_24888,N_22960,N_23837);
nand U24889 (N_24889,N_23566,N_23918);
and U24890 (N_24890,N_23857,N_23259);
nand U24891 (N_24891,N_23476,N_22754);
and U24892 (N_24892,N_23617,N_23405);
nand U24893 (N_24893,N_23838,N_23035);
and U24894 (N_24894,N_23570,N_22974);
or U24895 (N_24895,N_22792,N_23955);
or U24896 (N_24896,N_22873,N_22879);
and U24897 (N_24897,N_23372,N_22683);
and U24898 (N_24898,N_23823,N_22761);
nor U24899 (N_24899,N_22009,N_22399);
nor U24900 (N_24900,N_22950,N_22545);
nand U24901 (N_24901,N_23561,N_23449);
nand U24902 (N_24902,N_23604,N_23662);
nor U24903 (N_24903,N_23269,N_23718);
nand U24904 (N_24904,N_23687,N_22538);
nand U24905 (N_24905,N_22957,N_23790);
nor U24906 (N_24906,N_22862,N_23612);
nand U24907 (N_24907,N_22965,N_22032);
nor U24908 (N_24908,N_22183,N_22731);
xnor U24909 (N_24909,N_23836,N_23187);
nor U24910 (N_24910,N_22634,N_22609);
xor U24911 (N_24911,N_23206,N_22587);
xnor U24912 (N_24912,N_22938,N_23631);
xor U24913 (N_24913,N_23858,N_23272);
or U24914 (N_24914,N_22208,N_22972);
and U24915 (N_24915,N_23116,N_23328);
xor U24916 (N_24916,N_22858,N_22082);
or U24917 (N_24917,N_22791,N_22532);
or U24918 (N_24918,N_22439,N_22996);
nor U24919 (N_24919,N_23314,N_23445);
and U24920 (N_24920,N_22239,N_22852);
nand U24921 (N_24921,N_23098,N_22196);
xor U24922 (N_24922,N_23181,N_22755);
or U24923 (N_24923,N_23903,N_22003);
and U24924 (N_24924,N_22578,N_23380);
or U24925 (N_24925,N_22973,N_23469);
or U24926 (N_24926,N_23107,N_22180);
or U24927 (N_24927,N_23783,N_22053);
or U24928 (N_24928,N_22324,N_23938);
xnor U24929 (N_24929,N_22052,N_23738);
or U24930 (N_24930,N_22677,N_23554);
or U24931 (N_24931,N_22989,N_23563);
nor U24932 (N_24932,N_23183,N_22322);
nor U24933 (N_24933,N_23816,N_23079);
and U24934 (N_24934,N_23350,N_22313);
nand U24935 (N_24935,N_22471,N_23556);
nor U24936 (N_24936,N_22056,N_23205);
nor U24937 (N_24937,N_22793,N_23525);
nand U24938 (N_24938,N_23101,N_22443);
or U24939 (N_24939,N_22010,N_22600);
and U24940 (N_24940,N_22029,N_22283);
nor U24941 (N_24941,N_22932,N_22363);
nor U24942 (N_24942,N_22904,N_22766);
nand U24943 (N_24943,N_23159,N_23081);
and U24944 (N_24944,N_22054,N_22458);
nor U24945 (N_24945,N_22506,N_23619);
nor U24946 (N_24946,N_22163,N_22157);
or U24947 (N_24947,N_22669,N_22433);
nor U24948 (N_24948,N_23692,N_22394);
xor U24949 (N_24949,N_23304,N_22547);
xnor U24950 (N_24950,N_22317,N_22703);
nor U24951 (N_24951,N_23411,N_22209);
nor U24952 (N_24952,N_22951,N_22693);
nor U24953 (N_24953,N_22612,N_23517);
and U24954 (N_24954,N_23983,N_23412);
or U24955 (N_24955,N_22220,N_22775);
nand U24956 (N_24956,N_23435,N_23877);
xnor U24957 (N_24957,N_22226,N_22515);
nand U24958 (N_24958,N_23810,N_23475);
or U24959 (N_24959,N_22012,N_22275);
or U24960 (N_24960,N_22249,N_23197);
and U24961 (N_24961,N_22396,N_22045);
and U24962 (N_24962,N_23459,N_23472);
or U24963 (N_24963,N_22462,N_22866);
or U24964 (N_24964,N_22719,N_22976);
nand U24965 (N_24965,N_22595,N_22262);
or U24966 (N_24966,N_23365,N_22823);
nand U24967 (N_24967,N_22909,N_22727);
or U24968 (N_24968,N_23694,N_22432);
nor U24969 (N_24969,N_22346,N_22917);
or U24970 (N_24970,N_22429,N_22074);
or U24971 (N_24971,N_22023,N_23095);
and U24972 (N_24972,N_22081,N_23892);
nor U24973 (N_24973,N_22759,N_22668);
xnor U24974 (N_24974,N_23284,N_23722);
and U24975 (N_24975,N_22526,N_23288);
and U24976 (N_24976,N_22552,N_23437);
or U24977 (N_24977,N_23962,N_23948);
or U24978 (N_24978,N_22716,N_22944);
nand U24979 (N_24979,N_22452,N_23818);
nand U24980 (N_24980,N_23986,N_22942);
xor U24981 (N_24981,N_22908,N_22155);
nand U24982 (N_24982,N_22416,N_22060);
or U24983 (N_24983,N_23312,N_22147);
nand U24984 (N_24984,N_23971,N_23987);
nand U24985 (N_24985,N_22133,N_23636);
and U24986 (N_24986,N_23239,N_23985);
and U24987 (N_24987,N_22557,N_22948);
nor U24988 (N_24988,N_23377,N_23912);
nand U24989 (N_24989,N_23562,N_22836);
nor U24990 (N_24990,N_22261,N_23937);
nand U24991 (N_24991,N_23005,N_23395);
nor U24992 (N_24992,N_23322,N_23884);
nand U24993 (N_24993,N_23628,N_22927);
or U24994 (N_24994,N_23796,N_23309);
nor U24995 (N_24995,N_23886,N_23889);
and U24996 (N_24996,N_22807,N_22446);
nand U24997 (N_24997,N_23387,N_22804);
nand U24998 (N_24998,N_22809,N_23234);
or U24999 (N_24999,N_23649,N_22982);
or U25000 (N_25000,N_22569,N_23188);
or U25001 (N_25001,N_22619,N_23442);
and U25002 (N_25002,N_22563,N_22364);
and U25003 (N_25003,N_23458,N_23072);
or U25004 (N_25004,N_23430,N_22578);
nor U25005 (N_25005,N_22969,N_23979);
xnor U25006 (N_25006,N_22219,N_22702);
xor U25007 (N_25007,N_22977,N_23633);
xor U25008 (N_25008,N_22462,N_23568);
xor U25009 (N_25009,N_22326,N_23378);
or U25010 (N_25010,N_22510,N_23151);
nand U25011 (N_25011,N_22659,N_23108);
nand U25012 (N_25012,N_23810,N_23383);
nor U25013 (N_25013,N_22828,N_22181);
xnor U25014 (N_25014,N_23759,N_22636);
or U25015 (N_25015,N_23788,N_23503);
xor U25016 (N_25016,N_22064,N_23399);
or U25017 (N_25017,N_22010,N_22260);
nor U25018 (N_25018,N_23449,N_22969);
and U25019 (N_25019,N_22491,N_23058);
or U25020 (N_25020,N_23176,N_22084);
nand U25021 (N_25021,N_22367,N_23523);
or U25022 (N_25022,N_23135,N_22931);
nand U25023 (N_25023,N_23627,N_23100);
xnor U25024 (N_25024,N_22216,N_22081);
nor U25025 (N_25025,N_23051,N_23038);
or U25026 (N_25026,N_23548,N_22452);
xor U25027 (N_25027,N_23919,N_23540);
nand U25028 (N_25028,N_22976,N_22691);
and U25029 (N_25029,N_23726,N_22437);
and U25030 (N_25030,N_23860,N_23710);
nand U25031 (N_25031,N_23556,N_22978);
xor U25032 (N_25032,N_23106,N_22421);
or U25033 (N_25033,N_22443,N_22873);
or U25034 (N_25034,N_23015,N_22448);
nor U25035 (N_25035,N_23187,N_22888);
nand U25036 (N_25036,N_22126,N_23552);
and U25037 (N_25037,N_22220,N_23933);
and U25038 (N_25038,N_22807,N_23929);
and U25039 (N_25039,N_22454,N_22766);
and U25040 (N_25040,N_23154,N_22440);
nand U25041 (N_25041,N_23783,N_23572);
nand U25042 (N_25042,N_22550,N_22632);
or U25043 (N_25043,N_22002,N_22187);
or U25044 (N_25044,N_22698,N_22725);
and U25045 (N_25045,N_22376,N_22518);
and U25046 (N_25046,N_22083,N_23827);
nand U25047 (N_25047,N_23460,N_23602);
or U25048 (N_25048,N_23878,N_23306);
and U25049 (N_25049,N_22774,N_22541);
and U25050 (N_25050,N_23795,N_22874);
and U25051 (N_25051,N_23303,N_22521);
nor U25052 (N_25052,N_22709,N_22869);
and U25053 (N_25053,N_22073,N_22585);
nand U25054 (N_25054,N_23373,N_22423);
and U25055 (N_25055,N_22842,N_23764);
nand U25056 (N_25056,N_23893,N_22540);
xnor U25057 (N_25057,N_23973,N_22261);
and U25058 (N_25058,N_23399,N_22152);
nand U25059 (N_25059,N_23707,N_22985);
nand U25060 (N_25060,N_22391,N_22439);
xnor U25061 (N_25061,N_22391,N_23624);
and U25062 (N_25062,N_23797,N_22400);
nor U25063 (N_25063,N_22958,N_22070);
xnor U25064 (N_25064,N_22412,N_23235);
and U25065 (N_25065,N_22663,N_22456);
nand U25066 (N_25066,N_22005,N_22989);
xnor U25067 (N_25067,N_23925,N_23117);
and U25068 (N_25068,N_23221,N_23028);
xnor U25069 (N_25069,N_23411,N_22570);
xnor U25070 (N_25070,N_22437,N_23212);
nor U25071 (N_25071,N_23654,N_23472);
nor U25072 (N_25072,N_23481,N_23989);
and U25073 (N_25073,N_22785,N_22371);
or U25074 (N_25074,N_23377,N_22406);
or U25075 (N_25075,N_22747,N_22485);
and U25076 (N_25076,N_22331,N_22054);
nor U25077 (N_25077,N_22479,N_22146);
nand U25078 (N_25078,N_22979,N_22478);
or U25079 (N_25079,N_23516,N_22774);
and U25080 (N_25080,N_22167,N_22399);
nor U25081 (N_25081,N_23666,N_22184);
or U25082 (N_25082,N_23232,N_22578);
nand U25083 (N_25083,N_22901,N_22843);
nor U25084 (N_25084,N_22425,N_22449);
xnor U25085 (N_25085,N_22371,N_22381);
and U25086 (N_25086,N_23567,N_23137);
xnor U25087 (N_25087,N_22341,N_22780);
and U25088 (N_25088,N_22233,N_22296);
or U25089 (N_25089,N_22159,N_23657);
xor U25090 (N_25090,N_23021,N_22361);
and U25091 (N_25091,N_23396,N_22084);
nand U25092 (N_25092,N_22031,N_22385);
nor U25093 (N_25093,N_23914,N_22420);
nor U25094 (N_25094,N_22161,N_22624);
xor U25095 (N_25095,N_22776,N_23593);
nor U25096 (N_25096,N_23130,N_23016);
or U25097 (N_25097,N_23390,N_23864);
nor U25098 (N_25098,N_23042,N_23195);
nand U25099 (N_25099,N_22257,N_23794);
nand U25100 (N_25100,N_22008,N_23404);
xnor U25101 (N_25101,N_23350,N_23223);
or U25102 (N_25102,N_22738,N_23639);
and U25103 (N_25103,N_23179,N_23861);
nor U25104 (N_25104,N_23266,N_23233);
or U25105 (N_25105,N_23138,N_23773);
or U25106 (N_25106,N_22832,N_23790);
and U25107 (N_25107,N_23399,N_22361);
and U25108 (N_25108,N_22214,N_23413);
nand U25109 (N_25109,N_23919,N_22185);
or U25110 (N_25110,N_23598,N_23004);
and U25111 (N_25111,N_23524,N_22879);
or U25112 (N_25112,N_23262,N_22947);
xor U25113 (N_25113,N_22501,N_23532);
nor U25114 (N_25114,N_23161,N_23019);
and U25115 (N_25115,N_22928,N_22368);
nand U25116 (N_25116,N_23771,N_23580);
nor U25117 (N_25117,N_23766,N_22568);
xnor U25118 (N_25118,N_23489,N_23487);
nor U25119 (N_25119,N_22430,N_22955);
and U25120 (N_25120,N_23930,N_22883);
nor U25121 (N_25121,N_23432,N_23597);
xor U25122 (N_25122,N_23791,N_22800);
nand U25123 (N_25123,N_22306,N_22999);
nor U25124 (N_25124,N_23670,N_23019);
nand U25125 (N_25125,N_22513,N_22557);
and U25126 (N_25126,N_23637,N_23600);
and U25127 (N_25127,N_23306,N_23047);
nor U25128 (N_25128,N_23630,N_23635);
nor U25129 (N_25129,N_23721,N_22086);
xor U25130 (N_25130,N_23943,N_22587);
nor U25131 (N_25131,N_22098,N_22106);
xor U25132 (N_25132,N_22993,N_22502);
or U25133 (N_25133,N_23509,N_22059);
and U25134 (N_25134,N_22126,N_22384);
or U25135 (N_25135,N_23131,N_22317);
xor U25136 (N_25136,N_23083,N_23779);
xor U25137 (N_25137,N_23866,N_23282);
nand U25138 (N_25138,N_22231,N_22841);
nor U25139 (N_25139,N_22241,N_22357);
nand U25140 (N_25140,N_22568,N_22139);
and U25141 (N_25141,N_22892,N_23783);
or U25142 (N_25142,N_22024,N_23012);
and U25143 (N_25143,N_22594,N_23464);
nand U25144 (N_25144,N_22707,N_22142);
or U25145 (N_25145,N_23667,N_22444);
nand U25146 (N_25146,N_22504,N_23983);
and U25147 (N_25147,N_23314,N_22469);
xnor U25148 (N_25148,N_22653,N_22983);
nor U25149 (N_25149,N_23170,N_22734);
nand U25150 (N_25150,N_22221,N_22187);
nor U25151 (N_25151,N_23515,N_22172);
xnor U25152 (N_25152,N_23291,N_23585);
nand U25153 (N_25153,N_22521,N_22086);
nand U25154 (N_25154,N_22864,N_22452);
or U25155 (N_25155,N_23897,N_22282);
or U25156 (N_25156,N_22207,N_23707);
or U25157 (N_25157,N_23028,N_22226);
nor U25158 (N_25158,N_23558,N_23094);
and U25159 (N_25159,N_22427,N_22248);
or U25160 (N_25160,N_23255,N_23921);
nand U25161 (N_25161,N_23054,N_22723);
and U25162 (N_25162,N_22259,N_22514);
and U25163 (N_25163,N_22590,N_22714);
nor U25164 (N_25164,N_22043,N_23622);
nor U25165 (N_25165,N_23307,N_23208);
nor U25166 (N_25166,N_22269,N_22286);
xnor U25167 (N_25167,N_23511,N_23211);
and U25168 (N_25168,N_22092,N_22490);
nor U25169 (N_25169,N_22944,N_23084);
nor U25170 (N_25170,N_23961,N_22120);
or U25171 (N_25171,N_23509,N_22843);
xor U25172 (N_25172,N_22338,N_22796);
and U25173 (N_25173,N_22124,N_22662);
and U25174 (N_25174,N_22668,N_22930);
nand U25175 (N_25175,N_23507,N_23449);
nor U25176 (N_25176,N_23443,N_22940);
and U25177 (N_25177,N_22215,N_23417);
nor U25178 (N_25178,N_22919,N_23754);
nand U25179 (N_25179,N_22224,N_23021);
nor U25180 (N_25180,N_22603,N_23119);
xnor U25181 (N_25181,N_23784,N_23177);
or U25182 (N_25182,N_23089,N_22322);
nand U25183 (N_25183,N_22664,N_23793);
nor U25184 (N_25184,N_22216,N_22457);
or U25185 (N_25185,N_23323,N_22599);
and U25186 (N_25186,N_23695,N_22783);
and U25187 (N_25187,N_23842,N_23160);
and U25188 (N_25188,N_22371,N_23072);
or U25189 (N_25189,N_22269,N_23126);
nand U25190 (N_25190,N_23947,N_23364);
or U25191 (N_25191,N_23417,N_23497);
nor U25192 (N_25192,N_23863,N_23685);
nor U25193 (N_25193,N_23568,N_23542);
xnor U25194 (N_25194,N_22178,N_23224);
xor U25195 (N_25195,N_22528,N_22524);
nor U25196 (N_25196,N_23366,N_23699);
nand U25197 (N_25197,N_22643,N_23662);
nor U25198 (N_25198,N_23204,N_22337);
xnor U25199 (N_25199,N_23588,N_22083);
or U25200 (N_25200,N_22201,N_23980);
or U25201 (N_25201,N_23924,N_22231);
or U25202 (N_25202,N_22774,N_23808);
nor U25203 (N_25203,N_22948,N_23192);
nand U25204 (N_25204,N_22718,N_22356);
nor U25205 (N_25205,N_22036,N_22349);
and U25206 (N_25206,N_23555,N_23854);
or U25207 (N_25207,N_23259,N_22673);
or U25208 (N_25208,N_22251,N_23798);
nor U25209 (N_25209,N_22677,N_22345);
nor U25210 (N_25210,N_23053,N_22331);
or U25211 (N_25211,N_23912,N_23771);
nor U25212 (N_25212,N_22068,N_22950);
and U25213 (N_25213,N_23725,N_23523);
or U25214 (N_25214,N_23541,N_22526);
xnor U25215 (N_25215,N_22569,N_22147);
nand U25216 (N_25216,N_22538,N_22262);
or U25217 (N_25217,N_23317,N_23341);
nor U25218 (N_25218,N_23609,N_23896);
and U25219 (N_25219,N_23467,N_23199);
and U25220 (N_25220,N_22060,N_22395);
xor U25221 (N_25221,N_23573,N_22367);
nand U25222 (N_25222,N_22876,N_22195);
nand U25223 (N_25223,N_22850,N_23952);
xor U25224 (N_25224,N_23636,N_22049);
or U25225 (N_25225,N_23814,N_22652);
and U25226 (N_25226,N_22218,N_23897);
or U25227 (N_25227,N_22424,N_22308);
and U25228 (N_25228,N_22106,N_22217);
nor U25229 (N_25229,N_22224,N_23921);
nor U25230 (N_25230,N_22604,N_23793);
nand U25231 (N_25231,N_23687,N_22801);
and U25232 (N_25232,N_22514,N_23308);
or U25233 (N_25233,N_23368,N_22991);
and U25234 (N_25234,N_23745,N_22447);
or U25235 (N_25235,N_22680,N_23630);
and U25236 (N_25236,N_22050,N_22604);
nand U25237 (N_25237,N_22685,N_22848);
xor U25238 (N_25238,N_23435,N_22434);
or U25239 (N_25239,N_23101,N_23874);
nand U25240 (N_25240,N_22538,N_23941);
nand U25241 (N_25241,N_22678,N_23042);
and U25242 (N_25242,N_23219,N_22437);
nand U25243 (N_25243,N_22784,N_22909);
nor U25244 (N_25244,N_22310,N_22748);
nor U25245 (N_25245,N_22416,N_23625);
or U25246 (N_25246,N_23097,N_23079);
nor U25247 (N_25247,N_23844,N_22630);
nor U25248 (N_25248,N_22166,N_22494);
or U25249 (N_25249,N_22924,N_23029);
xor U25250 (N_25250,N_23085,N_22670);
or U25251 (N_25251,N_23666,N_22483);
nand U25252 (N_25252,N_23458,N_23982);
nor U25253 (N_25253,N_22925,N_23198);
nor U25254 (N_25254,N_22326,N_23498);
and U25255 (N_25255,N_23438,N_22186);
xor U25256 (N_25256,N_23558,N_22067);
and U25257 (N_25257,N_23427,N_23073);
or U25258 (N_25258,N_22207,N_22321);
or U25259 (N_25259,N_23033,N_23596);
and U25260 (N_25260,N_23356,N_23244);
and U25261 (N_25261,N_23882,N_23767);
or U25262 (N_25262,N_22508,N_22011);
or U25263 (N_25263,N_23131,N_23393);
or U25264 (N_25264,N_23393,N_23146);
nand U25265 (N_25265,N_22951,N_23895);
and U25266 (N_25266,N_22058,N_23130);
xnor U25267 (N_25267,N_23563,N_23472);
and U25268 (N_25268,N_23005,N_22538);
or U25269 (N_25269,N_23489,N_22189);
or U25270 (N_25270,N_23870,N_23020);
and U25271 (N_25271,N_23131,N_23648);
nand U25272 (N_25272,N_22024,N_22814);
nor U25273 (N_25273,N_22045,N_23951);
or U25274 (N_25274,N_23464,N_23546);
xnor U25275 (N_25275,N_23958,N_22526);
xor U25276 (N_25276,N_23980,N_23083);
or U25277 (N_25277,N_23051,N_22090);
and U25278 (N_25278,N_22460,N_22947);
or U25279 (N_25279,N_23931,N_23608);
nor U25280 (N_25280,N_23465,N_22518);
xor U25281 (N_25281,N_22421,N_22510);
nand U25282 (N_25282,N_23747,N_22361);
or U25283 (N_25283,N_23960,N_22683);
or U25284 (N_25284,N_22102,N_23212);
nand U25285 (N_25285,N_22098,N_22601);
nor U25286 (N_25286,N_22473,N_23870);
xnor U25287 (N_25287,N_23310,N_22586);
xor U25288 (N_25288,N_23143,N_22710);
nor U25289 (N_25289,N_23206,N_22971);
nor U25290 (N_25290,N_23406,N_22521);
xor U25291 (N_25291,N_22996,N_23785);
and U25292 (N_25292,N_22452,N_23564);
xnor U25293 (N_25293,N_23005,N_22604);
nand U25294 (N_25294,N_22365,N_23681);
and U25295 (N_25295,N_23204,N_23103);
and U25296 (N_25296,N_23702,N_23544);
or U25297 (N_25297,N_23831,N_22353);
and U25298 (N_25298,N_22666,N_22096);
and U25299 (N_25299,N_23310,N_22615);
xor U25300 (N_25300,N_23682,N_22766);
or U25301 (N_25301,N_23935,N_23464);
and U25302 (N_25302,N_22960,N_23855);
nand U25303 (N_25303,N_22477,N_22333);
and U25304 (N_25304,N_22719,N_23301);
nor U25305 (N_25305,N_23882,N_23129);
and U25306 (N_25306,N_23551,N_23897);
or U25307 (N_25307,N_22482,N_22666);
or U25308 (N_25308,N_22387,N_23640);
xor U25309 (N_25309,N_23095,N_22414);
nand U25310 (N_25310,N_23552,N_23485);
or U25311 (N_25311,N_23177,N_23473);
nor U25312 (N_25312,N_23191,N_22308);
nand U25313 (N_25313,N_22857,N_22709);
nand U25314 (N_25314,N_22266,N_23404);
or U25315 (N_25315,N_22868,N_22075);
or U25316 (N_25316,N_22696,N_22808);
xor U25317 (N_25317,N_22857,N_23455);
or U25318 (N_25318,N_23635,N_23431);
nor U25319 (N_25319,N_22654,N_22211);
nand U25320 (N_25320,N_23415,N_23384);
or U25321 (N_25321,N_22850,N_23670);
xor U25322 (N_25322,N_23191,N_23802);
nand U25323 (N_25323,N_23842,N_23022);
nand U25324 (N_25324,N_23165,N_23077);
and U25325 (N_25325,N_22622,N_22197);
xnor U25326 (N_25326,N_22986,N_23942);
and U25327 (N_25327,N_22758,N_23478);
nor U25328 (N_25328,N_22630,N_23280);
nor U25329 (N_25329,N_22092,N_22956);
and U25330 (N_25330,N_23410,N_22760);
and U25331 (N_25331,N_23081,N_22544);
xor U25332 (N_25332,N_23214,N_22782);
nor U25333 (N_25333,N_23235,N_22500);
nor U25334 (N_25334,N_23502,N_23473);
xnor U25335 (N_25335,N_23644,N_23120);
nand U25336 (N_25336,N_22174,N_22519);
nor U25337 (N_25337,N_23144,N_22381);
xor U25338 (N_25338,N_22544,N_22009);
xor U25339 (N_25339,N_22474,N_22931);
or U25340 (N_25340,N_22952,N_22334);
and U25341 (N_25341,N_23248,N_22672);
nor U25342 (N_25342,N_23626,N_23441);
and U25343 (N_25343,N_22811,N_22265);
and U25344 (N_25344,N_23413,N_22797);
or U25345 (N_25345,N_23056,N_23830);
and U25346 (N_25346,N_23830,N_22737);
nor U25347 (N_25347,N_22599,N_22629);
nor U25348 (N_25348,N_23151,N_23881);
xnor U25349 (N_25349,N_22320,N_23026);
nor U25350 (N_25350,N_22827,N_23923);
or U25351 (N_25351,N_23221,N_23915);
nand U25352 (N_25352,N_23335,N_23947);
nor U25353 (N_25353,N_23130,N_22436);
or U25354 (N_25354,N_23172,N_22761);
and U25355 (N_25355,N_22362,N_23798);
nor U25356 (N_25356,N_22336,N_22901);
or U25357 (N_25357,N_23446,N_23360);
and U25358 (N_25358,N_22435,N_22365);
xor U25359 (N_25359,N_22572,N_22617);
xnor U25360 (N_25360,N_22756,N_23406);
or U25361 (N_25361,N_22022,N_23266);
xor U25362 (N_25362,N_23269,N_23761);
and U25363 (N_25363,N_22792,N_22564);
or U25364 (N_25364,N_23540,N_23249);
xnor U25365 (N_25365,N_23075,N_23619);
or U25366 (N_25366,N_23318,N_23396);
nor U25367 (N_25367,N_23118,N_23534);
or U25368 (N_25368,N_23206,N_23904);
nand U25369 (N_25369,N_23941,N_22752);
xnor U25370 (N_25370,N_23964,N_22639);
nor U25371 (N_25371,N_23715,N_23048);
and U25372 (N_25372,N_22957,N_22523);
nor U25373 (N_25373,N_22350,N_22338);
and U25374 (N_25374,N_22235,N_23416);
nand U25375 (N_25375,N_22776,N_22689);
and U25376 (N_25376,N_23330,N_23282);
and U25377 (N_25377,N_23435,N_23532);
and U25378 (N_25378,N_23054,N_23260);
nand U25379 (N_25379,N_22512,N_22569);
and U25380 (N_25380,N_22812,N_22172);
xnor U25381 (N_25381,N_22486,N_23999);
xnor U25382 (N_25382,N_23570,N_22812);
xor U25383 (N_25383,N_23342,N_23010);
nor U25384 (N_25384,N_23226,N_23753);
and U25385 (N_25385,N_23625,N_22283);
xor U25386 (N_25386,N_23058,N_22145);
nand U25387 (N_25387,N_22917,N_23010);
and U25388 (N_25388,N_22127,N_22255);
nor U25389 (N_25389,N_22605,N_23099);
and U25390 (N_25390,N_23095,N_23707);
nor U25391 (N_25391,N_23683,N_23908);
xor U25392 (N_25392,N_22490,N_22355);
nor U25393 (N_25393,N_22455,N_22728);
and U25394 (N_25394,N_23458,N_23960);
and U25395 (N_25395,N_22921,N_23547);
xor U25396 (N_25396,N_23760,N_23614);
xor U25397 (N_25397,N_22280,N_22721);
and U25398 (N_25398,N_22280,N_23251);
nand U25399 (N_25399,N_23461,N_22355);
nor U25400 (N_25400,N_23846,N_23747);
nor U25401 (N_25401,N_22165,N_23888);
nor U25402 (N_25402,N_23436,N_22009);
and U25403 (N_25403,N_23584,N_23564);
nand U25404 (N_25404,N_23466,N_23817);
nand U25405 (N_25405,N_22873,N_22570);
xor U25406 (N_25406,N_22717,N_23988);
nand U25407 (N_25407,N_22024,N_23240);
nand U25408 (N_25408,N_22276,N_23484);
and U25409 (N_25409,N_22703,N_23319);
xnor U25410 (N_25410,N_23482,N_22287);
or U25411 (N_25411,N_23808,N_22867);
nor U25412 (N_25412,N_23747,N_23581);
or U25413 (N_25413,N_23938,N_22718);
nand U25414 (N_25414,N_22700,N_23046);
nand U25415 (N_25415,N_23235,N_22619);
and U25416 (N_25416,N_22967,N_22170);
or U25417 (N_25417,N_23189,N_22567);
nor U25418 (N_25418,N_22942,N_22695);
or U25419 (N_25419,N_23676,N_23875);
or U25420 (N_25420,N_23482,N_23976);
or U25421 (N_25421,N_23180,N_23030);
nand U25422 (N_25422,N_23531,N_22743);
xor U25423 (N_25423,N_23436,N_23611);
or U25424 (N_25424,N_23241,N_22625);
and U25425 (N_25425,N_22992,N_23979);
nor U25426 (N_25426,N_23172,N_22372);
nand U25427 (N_25427,N_23127,N_22214);
or U25428 (N_25428,N_23855,N_23126);
nor U25429 (N_25429,N_23160,N_23739);
nand U25430 (N_25430,N_23856,N_23605);
or U25431 (N_25431,N_23421,N_22563);
or U25432 (N_25432,N_23458,N_23984);
or U25433 (N_25433,N_22133,N_22923);
nor U25434 (N_25434,N_22031,N_23839);
or U25435 (N_25435,N_23386,N_23651);
nand U25436 (N_25436,N_23680,N_22258);
xnor U25437 (N_25437,N_22160,N_22884);
and U25438 (N_25438,N_22185,N_23788);
and U25439 (N_25439,N_23312,N_22987);
nor U25440 (N_25440,N_22631,N_22443);
nor U25441 (N_25441,N_22107,N_23318);
nor U25442 (N_25442,N_22013,N_22490);
xnor U25443 (N_25443,N_22982,N_22273);
nand U25444 (N_25444,N_23718,N_23511);
xor U25445 (N_25445,N_23608,N_22038);
nor U25446 (N_25446,N_23726,N_23300);
or U25447 (N_25447,N_22581,N_23888);
and U25448 (N_25448,N_22049,N_22754);
nand U25449 (N_25449,N_23261,N_23367);
or U25450 (N_25450,N_23880,N_22654);
xnor U25451 (N_25451,N_23881,N_22783);
and U25452 (N_25452,N_23424,N_22125);
and U25453 (N_25453,N_23035,N_22566);
xor U25454 (N_25454,N_23248,N_22807);
and U25455 (N_25455,N_23812,N_23650);
or U25456 (N_25456,N_23981,N_23615);
nor U25457 (N_25457,N_22861,N_23475);
nor U25458 (N_25458,N_23344,N_23002);
nand U25459 (N_25459,N_22077,N_23355);
xor U25460 (N_25460,N_22824,N_23475);
or U25461 (N_25461,N_22604,N_23598);
or U25462 (N_25462,N_22847,N_22011);
and U25463 (N_25463,N_22841,N_22490);
and U25464 (N_25464,N_23659,N_23154);
nand U25465 (N_25465,N_22461,N_23782);
and U25466 (N_25466,N_22389,N_22930);
or U25467 (N_25467,N_22781,N_23647);
xnor U25468 (N_25468,N_22919,N_22519);
nor U25469 (N_25469,N_22154,N_23373);
and U25470 (N_25470,N_22007,N_22039);
nor U25471 (N_25471,N_22979,N_23211);
or U25472 (N_25472,N_22451,N_22886);
nand U25473 (N_25473,N_23034,N_22435);
nor U25474 (N_25474,N_22278,N_23665);
nand U25475 (N_25475,N_22012,N_22286);
or U25476 (N_25476,N_22189,N_22550);
or U25477 (N_25477,N_23171,N_23394);
xor U25478 (N_25478,N_23774,N_23414);
nand U25479 (N_25479,N_22566,N_22620);
or U25480 (N_25480,N_23879,N_22613);
or U25481 (N_25481,N_23030,N_22574);
xor U25482 (N_25482,N_22339,N_23694);
nand U25483 (N_25483,N_23035,N_23244);
or U25484 (N_25484,N_23884,N_22569);
nand U25485 (N_25485,N_23936,N_22818);
nand U25486 (N_25486,N_23989,N_23071);
nand U25487 (N_25487,N_22303,N_23319);
nor U25488 (N_25488,N_22311,N_23893);
and U25489 (N_25489,N_23734,N_23250);
nor U25490 (N_25490,N_22274,N_22650);
or U25491 (N_25491,N_23826,N_22880);
nor U25492 (N_25492,N_23419,N_22686);
nor U25493 (N_25493,N_22213,N_23901);
or U25494 (N_25494,N_23545,N_22123);
nor U25495 (N_25495,N_22464,N_22608);
or U25496 (N_25496,N_23719,N_22218);
nand U25497 (N_25497,N_23038,N_22863);
xnor U25498 (N_25498,N_22264,N_22395);
nand U25499 (N_25499,N_23765,N_23324);
or U25500 (N_25500,N_22908,N_22304);
nand U25501 (N_25501,N_23287,N_23206);
nor U25502 (N_25502,N_22475,N_22011);
and U25503 (N_25503,N_22128,N_23211);
xnor U25504 (N_25504,N_23549,N_22676);
nor U25505 (N_25505,N_22411,N_23143);
xnor U25506 (N_25506,N_23305,N_23072);
xnor U25507 (N_25507,N_23027,N_23331);
xor U25508 (N_25508,N_22505,N_22286);
or U25509 (N_25509,N_23283,N_22996);
nor U25510 (N_25510,N_23015,N_22661);
or U25511 (N_25511,N_23809,N_22901);
or U25512 (N_25512,N_22717,N_22361);
xnor U25513 (N_25513,N_23339,N_23450);
xnor U25514 (N_25514,N_23877,N_22402);
xor U25515 (N_25515,N_23595,N_23771);
or U25516 (N_25516,N_22722,N_23425);
and U25517 (N_25517,N_23301,N_22352);
nand U25518 (N_25518,N_23427,N_22277);
nand U25519 (N_25519,N_23980,N_22098);
and U25520 (N_25520,N_23861,N_22186);
xnor U25521 (N_25521,N_23697,N_23726);
nand U25522 (N_25522,N_23496,N_23176);
or U25523 (N_25523,N_22410,N_23536);
xor U25524 (N_25524,N_22333,N_23206);
and U25525 (N_25525,N_22253,N_23494);
nand U25526 (N_25526,N_22498,N_22707);
xnor U25527 (N_25527,N_22375,N_23232);
xor U25528 (N_25528,N_23448,N_22786);
xor U25529 (N_25529,N_23575,N_22169);
nand U25530 (N_25530,N_22623,N_23571);
or U25531 (N_25531,N_22716,N_22764);
and U25532 (N_25532,N_23714,N_23177);
xor U25533 (N_25533,N_23630,N_23947);
or U25534 (N_25534,N_23625,N_23532);
nor U25535 (N_25535,N_23876,N_23712);
nand U25536 (N_25536,N_23178,N_22642);
nand U25537 (N_25537,N_23723,N_23895);
and U25538 (N_25538,N_23517,N_23349);
nor U25539 (N_25539,N_23185,N_22008);
and U25540 (N_25540,N_22618,N_22306);
nor U25541 (N_25541,N_23799,N_22743);
and U25542 (N_25542,N_23569,N_23456);
xnor U25543 (N_25543,N_23185,N_23459);
and U25544 (N_25544,N_23737,N_22895);
nand U25545 (N_25545,N_22585,N_23990);
xor U25546 (N_25546,N_23885,N_23874);
nor U25547 (N_25547,N_23401,N_23160);
and U25548 (N_25548,N_23969,N_22919);
nand U25549 (N_25549,N_22133,N_22233);
and U25550 (N_25550,N_23705,N_22695);
nand U25551 (N_25551,N_22560,N_23894);
nor U25552 (N_25552,N_22094,N_23722);
xor U25553 (N_25553,N_23601,N_23646);
nor U25554 (N_25554,N_23690,N_22467);
nor U25555 (N_25555,N_22922,N_22145);
or U25556 (N_25556,N_22670,N_23039);
xnor U25557 (N_25557,N_22113,N_22166);
and U25558 (N_25558,N_23994,N_22016);
or U25559 (N_25559,N_22164,N_23386);
xor U25560 (N_25560,N_22548,N_23073);
nand U25561 (N_25561,N_22193,N_23564);
xnor U25562 (N_25562,N_22339,N_22821);
nor U25563 (N_25563,N_23756,N_23017);
or U25564 (N_25564,N_23488,N_23979);
nand U25565 (N_25565,N_22290,N_22780);
nor U25566 (N_25566,N_23578,N_22743);
xnor U25567 (N_25567,N_22923,N_22952);
xnor U25568 (N_25568,N_22462,N_22102);
nand U25569 (N_25569,N_23822,N_23538);
nand U25570 (N_25570,N_23114,N_23339);
xor U25571 (N_25571,N_22521,N_23163);
nand U25572 (N_25572,N_23031,N_23909);
nand U25573 (N_25573,N_22203,N_23960);
xnor U25574 (N_25574,N_22744,N_22419);
and U25575 (N_25575,N_22188,N_22000);
or U25576 (N_25576,N_23546,N_23879);
and U25577 (N_25577,N_23980,N_22212);
and U25578 (N_25578,N_22362,N_23040);
nor U25579 (N_25579,N_22444,N_23063);
or U25580 (N_25580,N_23694,N_22919);
nor U25581 (N_25581,N_23416,N_23215);
nor U25582 (N_25582,N_23881,N_22612);
xor U25583 (N_25583,N_22007,N_22752);
nand U25584 (N_25584,N_23257,N_22614);
nor U25585 (N_25585,N_22110,N_23302);
nor U25586 (N_25586,N_22385,N_22894);
xor U25587 (N_25587,N_22094,N_22601);
nor U25588 (N_25588,N_22228,N_22082);
xor U25589 (N_25589,N_22909,N_23636);
nor U25590 (N_25590,N_22649,N_23666);
xnor U25591 (N_25591,N_23431,N_23677);
xor U25592 (N_25592,N_22663,N_22189);
xnor U25593 (N_25593,N_22560,N_23980);
xor U25594 (N_25594,N_22078,N_22678);
xor U25595 (N_25595,N_22450,N_23045);
and U25596 (N_25596,N_22554,N_23169);
nand U25597 (N_25597,N_22547,N_23253);
or U25598 (N_25598,N_22119,N_22998);
nand U25599 (N_25599,N_22115,N_22691);
and U25600 (N_25600,N_23207,N_23998);
nor U25601 (N_25601,N_22470,N_22213);
nor U25602 (N_25602,N_22164,N_22574);
or U25603 (N_25603,N_23756,N_22093);
or U25604 (N_25604,N_23273,N_23766);
nand U25605 (N_25605,N_22344,N_22235);
nor U25606 (N_25606,N_23879,N_22104);
nor U25607 (N_25607,N_22857,N_23388);
nor U25608 (N_25608,N_23694,N_23937);
nand U25609 (N_25609,N_22362,N_23109);
and U25610 (N_25610,N_23369,N_23965);
xor U25611 (N_25611,N_23304,N_23118);
xor U25612 (N_25612,N_23896,N_22761);
nor U25613 (N_25613,N_22203,N_22567);
nor U25614 (N_25614,N_22567,N_22979);
nand U25615 (N_25615,N_23250,N_23652);
or U25616 (N_25616,N_22850,N_23398);
or U25617 (N_25617,N_22455,N_23571);
nand U25618 (N_25618,N_23077,N_23836);
and U25619 (N_25619,N_22963,N_22854);
xnor U25620 (N_25620,N_23783,N_22737);
and U25621 (N_25621,N_22964,N_22696);
or U25622 (N_25622,N_22406,N_23873);
nand U25623 (N_25623,N_22431,N_23515);
nor U25624 (N_25624,N_22064,N_22132);
nand U25625 (N_25625,N_23817,N_22645);
nand U25626 (N_25626,N_22685,N_23281);
nor U25627 (N_25627,N_23113,N_22501);
and U25628 (N_25628,N_22274,N_22852);
nand U25629 (N_25629,N_23148,N_22651);
xor U25630 (N_25630,N_23897,N_23634);
xor U25631 (N_25631,N_23932,N_23063);
and U25632 (N_25632,N_23045,N_22546);
nand U25633 (N_25633,N_23530,N_23633);
nor U25634 (N_25634,N_22616,N_22647);
nor U25635 (N_25635,N_23546,N_22237);
nor U25636 (N_25636,N_22870,N_22338);
xor U25637 (N_25637,N_22764,N_23955);
xor U25638 (N_25638,N_22130,N_22255);
or U25639 (N_25639,N_23567,N_23447);
xnor U25640 (N_25640,N_22110,N_22034);
and U25641 (N_25641,N_23159,N_23133);
and U25642 (N_25642,N_22259,N_22742);
nor U25643 (N_25643,N_22464,N_22512);
or U25644 (N_25644,N_22725,N_22911);
or U25645 (N_25645,N_23935,N_22532);
nor U25646 (N_25646,N_23643,N_22378);
or U25647 (N_25647,N_23479,N_23579);
or U25648 (N_25648,N_23862,N_23688);
or U25649 (N_25649,N_22457,N_23647);
or U25650 (N_25650,N_23040,N_22882);
nand U25651 (N_25651,N_23044,N_22005);
and U25652 (N_25652,N_22330,N_22339);
or U25653 (N_25653,N_22291,N_23861);
and U25654 (N_25654,N_22195,N_22558);
nand U25655 (N_25655,N_23062,N_22967);
or U25656 (N_25656,N_23555,N_23453);
and U25657 (N_25657,N_23709,N_22222);
xor U25658 (N_25658,N_22053,N_22259);
or U25659 (N_25659,N_22445,N_23790);
xnor U25660 (N_25660,N_23147,N_22756);
and U25661 (N_25661,N_23411,N_22327);
or U25662 (N_25662,N_23277,N_22120);
nor U25663 (N_25663,N_23352,N_23686);
or U25664 (N_25664,N_22647,N_23242);
and U25665 (N_25665,N_23537,N_22179);
or U25666 (N_25666,N_23035,N_22952);
xor U25667 (N_25667,N_22775,N_23816);
nor U25668 (N_25668,N_22422,N_23586);
or U25669 (N_25669,N_22157,N_23667);
or U25670 (N_25670,N_22122,N_22804);
xnor U25671 (N_25671,N_23368,N_22709);
nor U25672 (N_25672,N_23551,N_22144);
nand U25673 (N_25673,N_22843,N_23699);
nand U25674 (N_25674,N_23971,N_22983);
and U25675 (N_25675,N_22645,N_22297);
nand U25676 (N_25676,N_22000,N_23856);
nor U25677 (N_25677,N_22808,N_23493);
and U25678 (N_25678,N_22237,N_23770);
nor U25679 (N_25679,N_23706,N_23276);
xnor U25680 (N_25680,N_22665,N_22846);
nor U25681 (N_25681,N_23939,N_23705);
xor U25682 (N_25682,N_22799,N_22287);
and U25683 (N_25683,N_22280,N_22636);
and U25684 (N_25684,N_23295,N_22925);
nor U25685 (N_25685,N_22004,N_23890);
nand U25686 (N_25686,N_23636,N_23706);
or U25687 (N_25687,N_22246,N_23499);
and U25688 (N_25688,N_22371,N_23817);
or U25689 (N_25689,N_23604,N_23992);
nor U25690 (N_25690,N_22127,N_23543);
nand U25691 (N_25691,N_22729,N_23228);
or U25692 (N_25692,N_22461,N_22436);
or U25693 (N_25693,N_22420,N_22088);
nor U25694 (N_25694,N_22149,N_23555);
nand U25695 (N_25695,N_23658,N_22490);
or U25696 (N_25696,N_22466,N_22607);
xor U25697 (N_25697,N_23071,N_22404);
nor U25698 (N_25698,N_23371,N_22630);
nor U25699 (N_25699,N_22846,N_23604);
or U25700 (N_25700,N_23011,N_23093);
nand U25701 (N_25701,N_22247,N_23442);
or U25702 (N_25702,N_23057,N_22820);
nor U25703 (N_25703,N_22584,N_22488);
and U25704 (N_25704,N_23823,N_22419);
and U25705 (N_25705,N_22870,N_23288);
nor U25706 (N_25706,N_23517,N_23252);
nor U25707 (N_25707,N_22181,N_23846);
or U25708 (N_25708,N_23390,N_22533);
or U25709 (N_25709,N_23524,N_22461);
nand U25710 (N_25710,N_23795,N_22126);
nand U25711 (N_25711,N_22181,N_23354);
nor U25712 (N_25712,N_23358,N_23272);
nand U25713 (N_25713,N_23464,N_23314);
and U25714 (N_25714,N_22547,N_22077);
and U25715 (N_25715,N_22661,N_22938);
nand U25716 (N_25716,N_23412,N_22008);
or U25717 (N_25717,N_22396,N_23512);
xor U25718 (N_25718,N_22509,N_23509);
xnor U25719 (N_25719,N_22716,N_23546);
or U25720 (N_25720,N_22141,N_23394);
nand U25721 (N_25721,N_22298,N_22575);
and U25722 (N_25722,N_23409,N_22431);
and U25723 (N_25723,N_23692,N_23815);
and U25724 (N_25724,N_22306,N_23277);
and U25725 (N_25725,N_23806,N_22745);
and U25726 (N_25726,N_23060,N_23824);
or U25727 (N_25727,N_22192,N_23530);
xor U25728 (N_25728,N_22581,N_23869);
nand U25729 (N_25729,N_22058,N_23303);
nor U25730 (N_25730,N_22591,N_22253);
and U25731 (N_25731,N_23794,N_23821);
xnor U25732 (N_25732,N_22036,N_23584);
nor U25733 (N_25733,N_23892,N_23004);
nand U25734 (N_25734,N_23958,N_23755);
or U25735 (N_25735,N_22873,N_22530);
or U25736 (N_25736,N_22850,N_22864);
nand U25737 (N_25737,N_23773,N_23339);
nor U25738 (N_25738,N_23119,N_22475);
nor U25739 (N_25739,N_22121,N_22765);
nor U25740 (N_25740,N_23134,N_23847);
nand U25741 (N_25741,N_23263,N_23536);
nor U25742 (N_25742,N_22770,N_22419);
nand U25743 (N_25743,N_22346,N_22640);
nor U25744 (N_25744,N_22554,N_22193);
and U25745 (N_25745,N_22215,N_22813);
or U25746 (N_25746,N_23036,N_23571);
nand U25747 (N_25747,N_22799,N_22419);
nand U25748 (N_25748,N_23867,N_22242);
and U25749 (N_25749,N_22378,N_23535);
or U25750 (N_25750,N_23146,N_22081);
xnor U25751 (N_25751,N_23740,N_22294);
or U25752 (N_25752,N_22970,N_23839);
or U25753 (N_25753,N_23954,N_22340);
xnor U25754 (N_25754,N_22744,N_23118);
nor U25755 (N_25755,N_23287,N_22466);
xor U25756 (N_25756,N_23843,N_23346);
or U25757 (N_25757,N_22744,N_23067);
or U25758 (N_25758,N_23878,N_23055);
nand U25759 (N_25759,N_23053,N_23515);
or U25760 (N_25760,N_23245,N_22794);
xnor U25761 (N_25761,N_23991,N_22884);
nand U25762 (N_25762,N_22465,N_22333);
and U25763 (N_25763,N_23404,N_22851);
and U25764 (N_25764,N_22888,N_22659);
or U25765 (N_25765,N_22328,N_22669);
nand U25766 (N_25766,N_22375,N_23056);
or U25767 (N_25767,N_23917,N_22925);
or U25768 (N_25768,N_22037,N_22103);
nor U25769 (N_25769,N_23825,N_22140);
or U25770 (N_25770,N_22264,N_23146);
or U25771 (N_25771,N_22465,N_23673);
and U25772 (N_25772,N_23107,N_22156);
or U25773 (N_25773,N_22175,N_23018);
nand U25774 (N_25774,N_22217,N_23949);
xor U25775 (N_25775,N_23131,N_22377);
nor U25776 (N_25776,N_22022,N_23032);
or U25777 (N_25777,N_23312,N_22275);
or U25778 (N_25778,N_23504,N_23141);
nand U25779 (N_25779,N_22367,N_23335);
xnor U25780 (N_25780,N_22523,N_23987);
and U25781 (N_25781,N_22635,N_22207);
nand U25782 (N_25782,N_23745,N_23480);
nor U25783 (N_25783,N_23751,N_23296);
and U25784 (N_25784,N_22050,N_22176);
and U25785 (N_25785,N_23654,N_22326);
nand U25786 (N_25786,N_22270,N_22214);
or U25787 (N_25787,N_23965,N_23020);
or U25788 (N_25788,N_23146,N_22045);
or U25789 (N_25789,N_23175,N_23597);
and U25790 (N_25790,N_23822,N_22506);
xor U25791 (N_25791,N_23226,N_22901);
nor U25792 (N_25792,N_22645,N_23220);
or U25793 (N_25793,N_22426,N_22976);
xnor U25794 (N_25794,N_23599,N_22360);
nor U25795 (N_25795,N_23899,N_23165);
nand U25796 (N_25796,N_22436,N_23957);
nor U25797 (N_25797,N_23437,N_22251);
and U25798 (N_25798,N_23706,N_23642);
nor U25799 (N_25799,N_22766,N_23559);
nand U25800 (N_25800,N_22546,N_23232);
nand U25801 (N_25801,N_23319,N_23878);
xor U25802 (N_25802,N_22355,N_23852);
xor U25803 (N_25803,N_22510,N_23284);
nand U25804 (N_25804,N_23262,N_23492);
or U25805 (N_25805,N_23204,N_23972);
or U25806 (N_25806,N_22911,N_23362);
or U25807 (N_25807,N_22887,N_22197);
nor U25808 (N_25808,N_23713,N_23606);
or U25809 (N_25809,N_23820,N_22097);
and U25810 (N_25810,N_22027,N_22880);
nand U25811 (N_25811,N_23147,N_22485);
nand U25812 (N_25812,N_23613,N_22147);
and U25813 (N_25813,N_23613,N_23577);
xor U25814 (N_25814,N_22868,N_22465);
nor U25815 (N_25815,N_22194,N_22102);
and U25816 (N_25816,N_23000,N_22967);
xor U25817 (N_25817,N_22916,N_23150);
and U25818 (N_25818,N_23499,N_22529);
xnor U25819 (N_25819,N_23569,N_23007);
or U25820 (N_25820,N_22371,N_22576);
nand U25821 (N_25821,N_23694,N_23733);
or U25822 (N_25822,N_23790,N_23191);
and U25823 (N_25823,N_22909,N_22560);
nand U25824 (N_25824,N_22835,N_23491);
nor U25825 (N_25825,N_22141,N_23497);
xnor U25826 (N_25826,N_22762,N_23825);
and U25827 (N_25827,N_22691,N_23651);
or U25828 (N_25828,N_23406,N_23708);
or U25829 (N_25829,N_23801,N_23115);
nand U25830 (N_25830,N_22995,N_23441);
nand U25831 (N_25831,N_23207,N_23950);
or U25832 (N_25832,N_23093,N_23335);
nor U25833 (N_25833,N_23219,N_23960);
and U25834 (N_25834,N_22308,N_22195);
nor U25835 (N_25835,N_23781,N_22510);
nor U25836 (N_25836,N_22921,N_22754);
nor U25837 (N_25837,N_23001,N_22160);
and U25838 (N_25838,N_22839,N_22707);
and U25839 (N_25839,N_22563,N_22227);
and U25840 (N_25840,N_22607,N_23747);
or U25841 (N_25841,N_22756,N_23074);
or U25842 (N_25842,N_23474,N_22003);
nand U25843 (N_25843,N_22019,N_22600);
xnor U25844 (N_25844,N_22915,N_22976);
or U25845 (N_25845,N_22870,N_22425);
xnor U25846 (N_25846,N_23332,N_23822);
or U25847 (N_25847,N_23506,N_23524);
nor U25848 (N_25848,N_23866,N_22241);
nor U25849 (N_25849,N_23314,N_23600);
or U25850 (N_25850,N_23529,N_22128);
xnor U25851 (N_25851,N_22295,N_23736);
or U25852 (N_25852,N_23616,N_22765);
or U25853 (N_25853,N_23162,N_23760);
nand U25854 (N_25854,N_22653,N_22353);
or U25855 (N_25855,N_22522,N_22468);
nand U25856 (N_25856,N_23450,N_23015);
nor U25857 (N_25857,N_22684,N_22820);
and U25858 (N_25858,N_22267,N_22605);
nand U25859 (N_25859,N_22731,N_23139);
nand U25860 (N_25860,N_23898,N_22671);
xor U25861 (N_25861,N_23158,N_22753);
nor U25862 (N_25862,N_23509,N_22767);
nand U25863 (N_25863,N_23546,N_23905);
nor U25864 (N_25864,N_23675,N_23775);
xnor U25865 (N_25865,N_22631,N_22587);
xor U25866 (N_25866,N_23177,N_22478);
xor U25867 (N_25867,N_22112,N_23844);
nand U25868 (N_25868,N_23737,N_22701);
nor U25869 (N_25869,N_22307,N_23645);
and U25870 (N_25870,N_22485,N_22008);
nand U25871 (N_25871,N_22656,N_23776);
and U25872 (N_25872,N_23805,N_22272);
and U25873 (N_25873,N_22491,N_22446);
and U25874 (N_25874,N_23142,N_23829);
nor U25875 (N_25875,N_23607,N_23370);
xor U25876 (N_25876,N_23251,N_22878);
xnor U25877 (N_25877,N_22090,N_22446);
and U25878 (N_25878,N_23300,N_22321);
and U25879 (N_25879,N_23343,N_23057);
nand U25880 (N_25880,N_23561,N_22166);
xor U25881 (N_25881,N_23069,N_23189);
nand U25882 (N_25882,N_22066,N_23251);
nor U25883 (N_25883,N_22715,N_22087);
or U25884 (N_25884,N_23595,N_22363);
or U25885 (N_25885,N_23397,N_22396);
xnor U25886 (N_25886,N_23871,N_22907);
nand U25887 (N_25887,N_23639,N_23903);
nor U25888 (N_25888,N_22527,N_23412);
xor U25889 (N_25889,N_23969,N_22570);
xnor U25890 (N_25890,N_22924,N_23365);
and U25891 (N_25891,N_22992,N_22267);
or U25892 (N_25892,N_23539,N_23999);
nand U25893 (N_25893,N_23976,N_23408);
xnor U25894 (N_25894,N_23556,N_23331);
and U25895 (N_25895,N_22518,N_23439);
or U25896 (N_25896,N_22270,N_23816);
xor U25897 (N_25897,N_23387,N_23264);
and U25898 (N_25898,N_22909,N_22492);
or U25899 (N_25899,N_22717,N_22093);
xnor U25900 (N_25900,N_23626,N_22351);
nor U25901 (N_25901,N_23614,N_23813);
nand U25902 (N_25902,N_22765,N_22530);
and U25903 (N_25903,N_23207,N_22862);
xor U25904 (N_25904,N_23630,N_23958);
and U25905 (N_25905,N_22221,N_22682);
or U25906 (N_25906,N_23896,N_23497);
and U25907 (N_25907,N_22727,N_22697);
nor U25908 (N_25908,N_23043,N_23489);
or U25909 (N_25909,N_22370,N_22006);
and U25910 (N_25910,N_23042,N_23824);
nor U25911 (N_25911,N_23674,N_23479);
and U25912 (N_25912,N_22845,N_22904);
nand U25913 (N_25913,N_22395,N_23427);
nand U25914 (N_25914,N_23918,N_22098);
xnor U25915 (N_25915,N_22063,N_23779);
and U25916 (N_25916,N_22126,N_23501);
xnor U25917 (N_25917,N_23725,N_23148);
nor U25918 (N_25918,N_22902,N_23050);
or U25919 (N_25919,N_23354,N_23635);
and U25920 (N_25920,N_23935,N_23755);
nand U25921 (N_25921,N_23693,N_23293);
and U25922 (N_25922,N_23768,N_22231);
xor U25923 (N_25923,N_22433,N_22293);
nand U25924 (N_25924,N_23163,N_22138);
nand U25925 (N_25925,N_23084,N_22360);
or U25926 (N_25926,N_22493,N_23946);
or U25927 (N_25927,N_23072,N_22249);
or U25928 (N_25928,N_23645,N_23386);
and U25929 (N_25929,N_23386,N_22851);
nor U25930 (N_25930,N_22342,N_22858);
and U25931 (N_25931,N_23961,N_22905);
nor U25932 (N_25932,N_22805,N_22621);
nand U25933 (N_25933,N_23260,N_22661);
nor U25934 (N_25934,N_23947,N_22199);
or U25935 (N_25935,N_23959,N_22285);
xor U25936 (N_25936,N_23582,N_23201);
or U25937 (N_25937,N_22822,N_22559);
and U25938 (N_25938,N_23524,N_23744);
xor U25939 (N_25939,N_22144,N_22802);
and U25940 (N_25940,N_23505,N_22857);
and U25941 (N_25941,N_23600,N_23811);
and U25942 (N_25942,N_22953,N_23668);
and U25943 (N_25943,N_22508,N_23934);
nor U25944 (N_25944,N_23348,N_22749);
and U25945 (N_25945,N_22580,N_23358);
and U25946 (N_25946,N_23351,N_23844);
xnor U25947 (N_25947,N_23084,N_22544);
nand U25948 (N_25948,N_22067,N_23951);
or U25949 (N_25949,N_23867,N_23803);
or U25950 (N_25950,N_23151,N_22548);
and U25951 (N_25951,N_23473,N_22552);
nand U25952 (N_25952,N_23782,N_22637);
nor U25953 (N_25953,N_23855,N_23069);
and U25954 (N_25954,N_23950,N_23906);
xor U25955 (N_25955,N_23151,N_23484);
nand U25956 (N_25956,N_22054,N_23390);
or U25957 (N_25957,N_22034,N_23241);
or U25958 (N_25958,N_22860,N_23598);
xnor U25959 (N_25959,N_23921,N_22254);
nand U25960 (N_25960,N_23378,N_22450);
or U25961 (N_25961,N_22672,N_23951);
xor U25962 (N_25962,N_23312,N_23810);
xnor U25963 (N_25963,N_23396,N_23970);
nand U25964 (N_25964,N_22200,N_23432);
and U25965 (N_25965,N_23115,N_22224);
or U25966 (N_25966,N_23911,N_23996);
nor U25967 (N_25967,N_22836,N_22613);
nand U25968 (N_25968,N_23904,N_23176);
nand U25969 (N_25969,N_22399,N_23780);
xnor U25970 (N_25970,N_23533,N_22704);
nor U25971 (N_25971,N_23824,N_22181);
nor U25972 (N_25972,N_23142,N_23425);
xnor U25973 (N_25973,N_22153,N_23810);
nor U25974 (N_25974,N_23278,N_22312);
nand U25975 (N_25975,N_23151,N_22606);
or U25976 (N_25976,N_22697,N_23169);
nand U25977 (N_25977,N_22513,N_22597);
nor U25978 (N_25978,N_22493,N_23464);
and U25979 (N_25979,N_23838,N_22921);
and U25980 (N_25980,N_23702,N_23126);
or U25981 (N_25981,N_23119,N_23358);
nand U25982 (N_25982,N_23270,N_23244);
nor U25983 (N_25983,N_23410,N_23751);
and U25984 (N_25984,N_23397,N_23186);
and U25985 (N_25985,N_23146,N_23287);
or U25986 (N_25986,N_22213,N_23004);
and U25987 (N_25987,N_22682,N_23285);
or U25988 (N_25988,N_22579,N_23687);
or U25989 (N_25989,N_22704,N_23447);
nand U25990 (N_25990,N_23618,N_22280);
nor U25991 (N_25991,N_22556,N_22510);
nand U25992 (N_25992,N_22176,N_22329);
and U25993 (N_25993,N_22460,N_23391);
and U25994 (N_25994,N_23075,N_23116);
nor U25995 (N_25995,N_22503,N_22335);
nand U25996 (N_25996,N_22660,N_22805);
xor U25997 (N_25997,N_22905,N_23936);
xnor U25998 (N_25998,N_22063,N_23055);
or U25999 (N_25999,N_22801,N_22486);
nand U26000 (N_26000,N_25622,N_25367);
nor U26001 (N_26001,N_24141,N_24840);
or U26002 (N_26002,N_25901,N_24559);
and U26003 (N_26003,N_25012,N_24556);
and U26004 (N_26004,N_25785,N_25372);
xnor U26005 (N_26005,N_24468,N_25655);
xnor U26006 (N_26006,N_24717,N_25362);
nand U26007 (N_26007,N_25846,N_25506);
xor U26008 (N_26008,N_24378,N_24104);
and U26009 (N_26009,N_24790,N_24457);
or U26010 (N_26010,N_25561,N_24059);
nor U26011 (N_26011,N_24796,N_25382);
xor U26012 (N_26012,N_25388,N_25228);
xnor U26013 (N_26013,N_24883,N_24052);
xor U26014 (N_26014,N_24508,N_25557);
xor U26015 (N_26015,N_25448,N_24325);
and U26016 (N_26016,N_24653,N_25498);
nor U26017 (N_26017,N_25163,N_24342);
and U26018 (N_26018,N_24408,N_24925);
xor U26019 (N_26019,N_25040,N_24304);
and U26020 (N_26020,N_25606,N_24595);
nor U26021 (N_26021,N_24841,N_24326);
or U26022 (N_26022,N_25106,N_24934);
or U26023 (N_26023,N_24194,N_25529);
and U26024 (N_26024,N_24176,N_25019);
nor U26025 (N_26025,N_25425,N_24709);
nand U26026 (N_26026,N_24875,N_24732);
nor U26027 (N_26027,N_24007,N_24598);
and U26028 (N_26028,N_25167,N_24880);
or U26029 (N_26029,N_24546,N_24578);
nor U26030 (N_26030,N_24624,N_25126);
or U26031 (N_26031,N_24359,N_24881);
xor U26032 (N_26032,N_24368,N_24096);
and U26033 (N_26033,N_24407,N_25240);
xnor U26034 (N_26034,N_24332,N_25594);
or U26035 (N_26035,N_25679,N_24908);
and U26036 (N_26036,N_24258,N_24714);
and U26037 (N_26037,N_25883,N_24197);
xnor U26038 (N_26038,N_24943,N_25495);
and U26039 (N_26039,N_25299,N_25755);
xor U26040 (N_26040,N_25139,N_24480);
and U26041 (N_26041,N_25663,N_24754);
nor U26042 (N_26042,N_25194,N_24386);
xnor U26043 (N_26043,N_25733,N_24092);
nand U26044 (N_26044,N_24370,N_24552);
nand U26045 (N_26045,N_25624,N_24612);
nor U26046 (N_26046,N_25693,N_25036);
nor U26047 (N_26047,N_24038,N_25055);
or U26048 (N_26048,N_25922,N_25789);
or U26049 (N_26049,N_25061,N_25598);
xor U26050 (N_26050,N_25107,N_24154);
and U26051 (N_26051,N_24244,N_25482);
or U26052 (N_26052,N_24954,N_24126);
nand U26053 (N_26053,N_24023,N_24681);
and U26054 (N_26054,N_25689,N_24355);
and U26055 (N_26055,N_25898,N_25586);
nor U26056 (N_26056,N_24662,N_24063);
xor U26057 (N_26057,N_25944,N_24238);
or U26058 (N_26058,N_25802,N_24808);
and U26059 (N_26059,N_24047,N_25373);
or U26060 (N_26060,N_25199,N_24986);
or U26061 (N_26061,N_25302,N_24240);
nor U26062 (N_26062,N_25083,N_24324);
or U26063 (N_26063,N_25026,N_24173);
or U26064 (N_26064,N_24418,N_25722);
nor U26065 (N_26065,N_25174,N_25831);
or U26066 (N_26066,N_25243,N_25977);
or U26067 (N_26067,N_24167,N_25236);
nand U26068 (N_26068,N_25763,N_24311);
and U26069 (N_26069,N_25752,N_24530);
nor U26070 (N_26070,N_24466,N_24435);
or U26071 (N_26071,N_25232,N_25468);
or U26072 (N_26072,N_25874,N_24810);
or U26073 (N_26073,N_24540,N_24235);
nand U26074 (N_26074,N_24011,N_25278);
and U26075 (N_26075,N_25133,N_24737);
xor U26076 (N_26076,N_24242,N_25027);
nor U26077 (N_26077,N_24688,N_25966);
nand U26078 (N_26078,N_25079,N_24006);
and U26079 (N_26079,N_25738,N_24032);
xnor U26080 (N_26080,N_24166,N_25974);
nand U26081 (N_26081,N_24294,N_24895);
nor U26082 (N_26082,N_25513,N_25590);
or U26083 (N_26083,N_24222,N_24781);
or U26084 (N_26084,N_24297,N_25021);
xnor U26085 (N_26085,N_25345,N_25400);
or U26086 (N_26086,N_25016,N_24536);
xnor U26087 (N_26087,N_24769,N_25955);
nand U26088 (N_26088,N_24017,N_24267);
nand U26089 (N_26089,N_25409,N_25288);
xor U26090 (N_26090,N_24905,N_25798);
or U26091 (N_26091,N_25125,N_24163);
nor U26092 (N_26092,N_24093,N_24272);
nand U26093 (N_26093,N_25249,N_24973);
nand U26094 (N_26094,N_24392,N_24147);
and U26095 (N_26095,N_25701,N_24060);
nand U26096 (N_26096,N_24089,N_25554);
nand U26097 (N_26097,N_25092,N_25844);
nor U26098 (N_26098,N_25749,N_24557);
xnor U26099 (N_26099,N_24462,N_25993);
and U26100 (N_26100,N_25503,N_24286);
nand U26101 (N_26101,N_25587,N_24682);
xor U26102 (N_26102,N_24277,N_25671);
or U26103 (N_26103,N_24562,N_25029);
xor U26104 (N_26104,N_25958,N_24886);
and U26105 (N_26105,N_24597,N_25965);
xor U26106 (N_26106,N_25782,N_25295);
nor U26107 (N_26107,N_25322,N_25810);
nand U26108 (N_26108,N_25218,N_24478);
xor U26109 (N_26109,N_25850,N_25268);
nor U26110 (N_26110,N_24005,N_25775);
xnor U26111 (N_26111,N_25245,N_24170);
and U26112 (N_26112,N_25632,N_24581);
xnor U26113 (N_26113,N_25510,N_24892);
nor U26114 (N_26114,N_24069,N_25523);
and U26115 (N_26115,N_25215,N_24471);
or U26116 (N_26116,N_24700,N_25207);
xnor U26117 (N_26117,N_24202,N_24078);
nor U26118 (N_26118,N_24554,N_25313);
nor U26119 (N_26119,N_24763,N_25686);
or U26120 (N_26120,N_25178,N_25328);
nor U26121 (N_26121,N_25481,N_25073);
nand U26122 (N_26122,N_24499,N_25975);
or U26123 (N_26123,N_24136,N_25407);
xor U26124 (N_26124,N_25766,N_24169);
and U26125 (N_26125,N_25282,N_25332);
nand U26126 (N_26126,N_25496,N_24778);
xor U26127 (N_26127,N_25440,N_25337);
and U26128 (N_26128,N_25238,N_25334);
nor U26129 (N_26129,N_25880,N_25473);
xnor U26130 (N_26130,N_24659,N_24230);
nand U26131 (N_26131,N_25104,N_25378);
or U26132 (N_26132,N_25540,N_24551);
xor U26133 (N_26133,N_24834,N_25556);
and U26134 (N_26134,N_25475,N_24181);
or U26135 (N_26135,N_25274,N_25369);
and U26136 (N_26136,N_24034,N_24627);
or U26137 (N_26137,N_24817,N_24933);
or U26138 (N_26138,N_25786,N_24292);
or U26139 (N_26139,N_24850,N_24381);
nand U26140 (N_26140,N_24931,N_25262);
nand U26141 (N_26141,N_25401,N_25978);
or U26142 (N_26142,N_25152,N_25264);
nand U26143 (N_26143,N_24560,N_25197);
nand U26144 (N_26144,N_25287,N_25768);
and U26145 (N_26145,N_25939,N_24869);
xor U26146 (N_26146,N_24485,N_25921);
nand U26147 (N_26147,N_24847,N_24839);
xor U26148 (N_26148,N_25374,N_24882);
nand U26149 (N_26149,N_24582,N_24003);
or U26150 (N_26150,N_24511,N_25331);
and U26151 (N_26151,N_24199,N_25805);
nor U26152 (N_26152,N_25416,N_24358);
nand U26153 (N_26153,N_25971,N_24549);
nand U26154 (N_26154,N_25934,N_25698);
xnor U26155 (N_26155,N_24906,N_24309);
xor U26156 (N_26156,N_25682,N_24842);
or U26157 (N_26157,N_25354,N_25000);
xnor U26158 (N_26158,N_24362,N_24844);
xnor U26159 (N_26159,N_24125,N_24164);
nor U26160 (N_26160,N_25269,N_25572);
nor U26161 (N_26161,N_25998,N_25352);
nand U26162 (N_26162,N_24716,N_24264);
nand U26163 (N_26163,N_25414,N_25730);
xor U26164 (N_26164,N_25518,N_24045);
nand U26165 (N_26165,N_24432,N_24901);
or U26166 (N_26166,N_25060,N_25509);
xor U26167 (N_26167,N_25108,N_24155);
nand U26168 (N_26168,N_25246,N_24062);
xor U26169 (N_26169,N_24116,N_24467);
and U26170 (N_26170,N_24723,N_24000);
xnor U26171 (N_26171,N_25987,N_24864);
and U26172 (N_26172,N_25899,N_24777);
nor U26173 (N_26173,N_25402,N_24140);
and U26174 (N_26174,N_24733,N_24825);
xnor U26175 (N_26175,N_24833,N_24831);
nand U26176 (N_26176,N_24520,N_24448);
nand U26177 (N_26177,N_24268,N_24870);
nor U26178 (N_26178,N_24541,N_24036);
nor U26179 (N_26179,N_24106,N_24745);
nor U26180 (N_26180,N_24192,N_24305);
xor U26181 (N_26181,N_24132,N_25216);
or U26182 (N_26182,N_24439,N_25330);
and U26183 (N_26183,N_25521,N_24879);
and U26184 (N_26184,N_25289,N_25643);
xnor U26185 (N_26185,N_25032,N_25592);
xor U26186 (N_26186,N_24018,N_25001);
nor U26187 (N_26187,N_25989,N_24385);
nand U26188 (N_26188,N_24718,N_25186);
xnor U26189 (N_26189,N_25210,N_25852);
xnor U26190 (N_26190,N_25385,N_24066);
nand U26191 (N_26191,N_25563,N_25739);
or U26192 (N_26192,N_25536,N_25371);
or U26193 (N_26193,N_25484,N_25648);
nor U26194 (N_26194,N_24608,N_24698);
nor U26195 (N_26195,N_24535,N_24832);
nand U26196 (N_26196,N_25076,N_24758);
or U26197 (N_26197,N_24261,N_25415);
or U26198 (N_26198,N_25122,N_24633);
or U26199 (N_26199,N_25910,N_24487);
nand U26200 (N_26200,N_24942,N_24110);
xnor U26201 (N_26201,N_24214,N_25062);
or U26202 (N_26202,N_25166,N_24975);
nor U26203 (N_26203,N_24306,N_24295);
nand U26204 (N_26204,N_25926,N_24959);
nor U26205 (N_26205,N_24053,N_25875);
nand U26206 (N_26206,N_25773,N_24755);
or U26207 (N_26207,N_25028,N_25273);
and U26208 (N_26208,N_24970,N_24372);
and U26209 (N_26209,N_25658,N_25239);
nand U26210 (N_26210,N_24437,N_24412);
and U26211 (N_26211,N_24013,N_24186);
nor U26212 (N_26212,N_25584,N_24803);
and U26213 (N_26213,N_25830,N_25960);
and U26214 (N_26214,N_25145,N_25767);
or U26215 (N_26215,N_25726,N_25353);
or U26216 (N_26216,N_24419,N_24730);
nand U26217 (N_26217,N_25010,N_25422);
nand U26218 (N_26218,N_24746,N_24087);
xnor U26219 (N_26219,N_25680,N_25790);
or U26220 (N_26220,N_25255,N_25728);
nor U26221 (N_26221,N_25427,N_25602);
and U26222 (N_26222,N_24494,N_25717);
and U26223 (N_26223,N_24914,N_25368);
and U26224 (N_26224,N_24231,N_24009);
nand U26225 (N_26225,N_24791,N_24016);
nand U26226 (N_26226,N_25408,N_24657);
nor U26227 (N_26227,N_24955,N_24739);
nor U26228 (N_26228,N_24293,N_24981);
or U26229 (N_26229,N_25150,N_24204);
or U26230 (N_26230,N_24191,N_24585);
nand U26231 (N_26231,N_24428,N_25450);
nand U26232 (N_26232,N_25996,N_24450);
nand U26233 (N_26233,N_24134,N_25031);
nand U26234 (N_26234,N_25222,N_25777);
xnor U26235 (N_26235,N_25277,N_25668);
nor U26236 (N_26236,N_25033,N_24524);
or U26237 (N_26237,N_24650,N_24940);
or U26238 (N_26238,N_25653,N_25872);
and U26239 (N_26239,N_25393,N_25864);
xnor U26240 (N_26240,N_25142,N_25307);
or U26241 (N_26241,N_24610,N_25300);
or U26242 (N_26242,N_24097,N_25636);
nor U26243 (N_26243,N_25237,N_24082);
nor U26244 (N_26244,N_24918,N_24399);
xor U26245 (N_26245,N_25477,N_25603);
xor U26246 (N_26246,N_24949,N_25363);
xnor U26247 (N_26247,N_24960,N_24697);
nor U26248 (N_26248,N_24517,N_25044);
or U26249 (N_26249,N_25100,N_25570);
nand U26250 (N_26250,N_24902,N_25615);
and U26251 (N_26251,N_25946,N_25418);
nand U26252 (N_26252,N_25014,N_25641);
xor U26253 (N_26253,N_24491,N_24426);
and U26254 (N_26254,N_24587,N_24247);
and U26255 (N_26255,N_24002,N_25847);
nor U26256 (N_26256,N_24794,N_25213);
xor U26257 (N_26257,N_24656,N_25630);
xnor U26258 (N_26258,N_25054,N_25169);
nand U26259 (N_26259,N_25203,N_25911);
or U26260 (N_26260,N_24396,N_25897);
or U26261 (N_26261,N_24857,N_24804);
or U26262 (N_26262,N_24458,N_25067);
xnor U26263 (N_26263,N_25135,N_24276);
nor U26264 (N_26264,N_25346,N_24775);
xnor U26265 (N_26265,N_25357,N_25608);
nand U26266 (N_26266,N_25294,N_25168);
xor U26267 (N_26267,N_24686,N_24665);
nor U26268 (N_26268,N_25544,N_25140);
xnor U26269 (N_26269,N_25283,N_24065);
nand U26270 (N_26270,N_24724,N_25404);
xnor U26271 (N_26271,N_25355,N_25182);
nand U26272 (N_26272,N_25486,N_25549);
xnor U26273 (N_26273,N_24427,N_25480);
xor U26274 (N_26274,N_25659,N_24913);
and U26275 (N_26275,N_25924,N_24376);
xnor U26276 (N_26276,N_24489,N_25799);
nand U26277 (N_26277,N_24084,N_25008);
nand U26278 (N_26278,N_25751,N_24707);
and U26279 (N_26279,N_25543,N_25131);
or U26280 (N_26280,N_24798,N_25015);
and U26281 (N_26281,N_25928,N_24492);
xor U26282 (N_26282,N_25715,N_25758);
nand U26283 (N_26283,N_24932,N_25979);
nor U26284 (N_26284,N_25644,N_25596);
or U26285 (N_26285,N_25565,N_24938);
nor U26286 (N_26286,N_24976,N_25320);
xor U26287 (N_26287,N_24014,N_25128);
xor U26288 (N_26288,N_24507,N_25149);
nor U26289 (N_26289,N_25241,N_25419);
and U26290 (N_26290,N_24460,N_25259);
nand U26291 (N_26291,N_24980,N_24979);
xnor U26292 (N_26292,N_24805,N_24671);
xor U26293 (N_26293,N_25716,N_24690);
or U26294 (N_26294,N_24843,N_24958);
or U26295 (N_26295,N_24056,N_24080);
nand U26296 (N_26296,N_25059,N_25386);
or U26297 (N_26297,N_25957,N_24122);
nor U26298 (N_26298,N_25562,N_24811);
nor U26299 (N_26299,N_25547,N_24547);
or U26300 (N_26300,N_24788,N_25508);
and U26301 (N_26301,N_25146,N_25248);
and U26302 (N_26302,N_25711,N_24022);
or U26303 (N_26303,N_24074,N_24505);
or U26304 (N_26304,N_25629,N_25639);
xor U26305 (N_26305,N_24413,N_24635);
nand U26306 (N_26306,N_25022,N_25360);
xor U26307 (N_26307,N_24675,N_24626);
or U26308 (N_26308,N_25493,N_24433);
and U26309 (N_26309,N_25905,N_24897);
xnor U26310 (N_26310,N_24298,N_25976);
or U26311 (N_26311,N_25896,N_24229);
xor U26312 (N_26312,N_25390,N_24838);
and U26313 (N_26313,N_25856,N_24691);
xor U26314 (N_26314,N_25023,N_25765);
nor U26315 (N_26315,N_24701,N_25500);
nor U26316 (N_26316,N_25340,N_25754);
xnor U26317 (N_26317,N_25172,N_24565);
or U26318 (N_26318,N_25938,N_25980);
nor U26319 (N_26319,N_25963,N_24592);
or U26320 (N_26320,N_24638,N_25610);
nand U26321 (N_26321,N_24713,N_25075);
and U26322 (N_26322,N_25490,N_24274);
or U26323 (N_26323,N_24421,N_25187);
or U26324 (N_26324,N_25969,N_25311);
and U26325 (N_26325,N_25970,N_24951);
nor U26326 (N_26326,N_24211,N_24963);
xor U26327 (N_26327,N_25826,N_24534);
xor U26328 (N_26328,N_25165,N_24177);
and U26329 (N_26329,N_25815,N_25375);
or U26330 (N_26330,N_24072,N_24137);
nor U26331 (N_26331,N_24406,N_24878);
and U26332 (N_26332,N_25553,N_24148);
xnor U26333 (N_26333,N_25058,N_24890);
nor U26334 (N_26334,N_25449,N_25464);
xor U26335 (N_26335,N_24631,N_24178);
or U26336 (N_26336,N_25838,N_25209);
or U26337 (N_26337,N_25784,N_25515);
nand U26338 (N_26338,N_25051,N_25545);
and U26339 (N_26339,N_24785,N_24307);
and U26340 (N_26340,N_25964,N_25792);
or U26341 (N_26341,N_24899,N_25942);
nand U26342 (N_26342,N_24498,N_25379);
nand U26343 (N_26343,N_24795,N_24422);
xor U26344 (N_26344,N_25551,N_25217);
xnor U26345 (N_26345,N_25229,N_24188);
nand U26346 (N_26346,N_24389,N_25256);
or U26347 (N_26347,N_25310,N_24030);
and U26348 (N_26348,N_24699,N_25293);
nand U26349 (N_26349,N_25667,N_24715);
and U26350 (N_26350,N_25077,N_24826);
nor U26351 (N_26351,N_24175,N_24083);
xor U26352 (N_26352,N_24760,N_25552);
or U26353 (N_26353,N_24361,N_25907);
and U26354 (N_26354,N_24900,N_25635);
nand U26355 (N_26355,N_24752,N_25043);
xnor U26356 (N_26356,N_25941,N_25861);
xnor U26357 (N_26357,N_25589,N_24430);
or U26358 (N_26358,N_25651,N_24319);
or U26359 (N_26359,N_25338,N_25597);
xnor U26360 (N_26360,N_24996,N_24377);
or U26361 (N_26361,N_24569,N_24680);
and U26362 (N_26362,N_24600,N_24004);
and U26363 (N_26363,N_25528,N_24367);
nand U26364 (N_26364,N_25524,N_25951);
nor U26365 (N_26365,N_25640,N_24866);
and U26366 (N_26366,N_25889,N_25753);
or U26367 (N_26367,N_25292,N_24772);
nand U26368 (N_26368,N_25647,N_24607);
and U26369 (N_26369,N_25699,N_24010);
and U26370 (N_26370,N_25984,N_24320);
nand U26371 (N_26371,N_24454,N_25746);
and U26372 (N_26372,N_24269,N_24046);
xnor U26373 (N_26373,N_24246,N_24613);
xnor U26374 (N_26374,N_25392,N_24997);
nand U26375 (N_26375,N_24363,N_25607);
and U26376 (N_26376,N_25638,N_25162);
nor U26377 (N_26377,N_25297,N_25961);
nor U26378 (N_26378,N_24260,N_25115);
or U26379 (N_26379,N_24497,N_24510);
xor U26380 (N_26380,N_24995,N_25931);
and U26381 (N_26381,N_24216,N_25406);
and U26382 (N_26382,N_25727,N_25492);
or U26383 (N_26383,N_24139,N_25483);
and U26384 (N_26384,N_24232,N_25933);
nand U26385 (N_26385,N_24917,N_24220);
xnor U26386 (N_26386,N_24217,N_25575);
nand U26387 (N_26387,N_25835,N_24887);
xor U26388 (N_26388,N_25394,N_25116);
and U26389 (N_26389,N_25892,N_24473);
xor U26390 (N_26390,N_25441,N_24584);
xor U26391 (N_26391,N_25954,N_24088);
and U26392 (N_26392,N_25319,N_25814);
nand U26393 (N_26393,N_24212,N_24543);
xor U26394 (N_26394,N_25411,N_25772);
nand U26395 (N_26395,N_25837,N_25403);
or U26396 (N_26396,N_25621,N_24764);
xnor U26397 (N_26397,N_25451,N_25863);
nor U26398 (N_26398,N_25020,N_24356);
nor U26399 (N_26399,N_24513,N_25323);
nor U26400 (N_26400,N_25176,N_24770);
xnor U26401 (N_26401,N_24904,N_24742);
xor U26402 (N_26402,N_24652,N_24663);
nor U26403 (N_26403,N_24567,N_24153);
xor U26404 (N_26404,N_25309,N_24391);
nand U26405 (N_26405,N_24079,N_24636);
or U26406 (N_26406,N_25432,N_24371);
and U26407 (N_26407,N_24446,N_25456);
nor U26408 (N_26408,N_24865,N_25770);
or U26409 (N_26409,N_24693,N_25779);
nor U26410 (N_26410,N_25819,N_24133);
and U26411 (N_26411,N_25823,N_24364);
or U26412 (N_26412,N_25927,N_24678);
and U26413 (N_26413,N_25462,N_25325);
xnor U26414 (N_26414,N_25737,N_25223);
or U26415 (N_26415,N_24150,N_24621);
nand U26416 (N_26416,N_24819,N_24874);
or U26417 (N_26417,N_25709,N_24666);
nor U26418 (N_26418,N_24784,N_25291);
nand U26419 (N_26419,N_24187,N_25821);
xor U26420 (N_26420,N_24655,N_24720);
xor U26421 (N_26421,N_25646,N_25081);
nor U26422 (N_26422,N_24035,N_25327);
nand U26423 (N_26423,N_24509,N_25817);
nor U26424 (N_26424,N_25522,N_24317);
xnor U26425 (N_26425,N_25003,N_24486);
xnor U26426 (N_26426,N_24369,N_24296);
xor U26427 (N_26427,N_24189,N_25049);
or U26428 (N_26428,N_25806,N_24206);
nor U26429 (N_26429,N_24158,N_24401);
or U26430 (N_26430,N_25206,N_24330);
nor U26431 (N_26431,N_24257,N_24395);
and U26432 (N_26432,N_24768,N_25445);
and U26433 (N_26433,N_24112,N_24165);
and U26434 (N_26434,N_25041,N_24818);
nor U26435 (N_26435,N_24783,N_24251);
xor U26436 (N_26436,N_25258,N_25499);
and U26437 (N_26437,N_25913,N_25383);
or U26438 (N_26438,N_25748,N_25617);
nand U26439 (N_26439,N_25064,N_25326);
xnor U26440 (N_26440,N_25613,N_24321);
and U26441 (N_26441,N_24920,N_24452);
and U26442 (N_26442,N_25343,N_25380);
nand U26443 (N_26443,N_25953,N_25950);
and U26444 (N_26444,N_24533,N_25488);
nand U26445 (N_26445,N_24226,N_24210);
or U26446 (N_26446,N_24314,N_24806);
or U26447 (N_26447,N_24512,N_24807);
xnor U26448 (N_26448,N_24442,N_25395);
or U26449 (N_26449,N_24252,N_25398);
nor U26450 (N_26450,N_25242,N_25042);
nand U26451 (N_26451,N_24606,N_24503);
xor U26452 (N_26452,N_25858,N_25376);
and U26453 (N_26453,N_25886,N_24278);
xnor U26454 (N_26454,N_25705,N_24704);
or U26455 (N_26455,N_24644,N_24623);
or U26456 (N_26456,N_24926,N_25878);
nand U26457 (N_26457,N_25202,N_25566);
or U26458 (N_26458,N_25829,N_25860);
nor U26459 (N_26459,N_24989,N_25038);
or U26460 (N_26460,N_24459,N_25902);
and U26461 (N_26461,N_25633,N_25112);
or U26462 (N_26462,N_24207,N_24984);
nand U26463 (N_26463,N_24521,N_25849);
nor U26464 (N_26464,N_25691,N_24402);
or U26465 (N_26465,N_25904,N_24922);
xor U26466 (N_26466,N_25891,N_24425);
or U26467 (N_26467,N_25072,N_25795);
nand U26468 (N_26468,N_24143,N_25917);
or U26469 (N_26469,N_24771,N_25595);
nor U26470 (N_26470,N_24779,N_25855);
xnor U26471 (N_26471,N_25429,N_25571);
and U26472 (N_26472,N_25600,N_25903);
nor U26473 (N_26473,N_24256,N_25949);
nor U26474 (N_26474,N_25339,N_25712);
xor U26475 (N_26475,N_24345,N_25442);
and U26476 (N_26476,N_25577,N_24113);
nand U26477 (N_26477,N_25143,N_24930);
nor U26478 (N_26478,N_24893,N_25656);
nor U26479 (N_26479,N_24916,N_25505);
xor U26480 (N_26480,N_25614,N_24537);
xnor U26481 (N_26481,N_24673,N_25947);
nand U26482 (N_26482,N_25757,N_25487);
nor U26483 (N_26483,N_25736,N_24328);
and U26484 (N_26484,N_25895,N_25284);
or U26485 (N_26485,N_25714,N_25454);
xor U26486 (N_26486,N_24077,N_24145);
and U26487 (N_26487,N_24338,N_25281);
xor U26488 (N_26488,N_25191,N_25006);
and U26489 (N_26489,N_24625,N_25873);
xor U26490 (N_26490,N_24195,N_24928);
nor U26491 (N_26491,N_24390,N_24453);
nand U26492 (N_26492,N_24168,N_24646);
nand U26493 (N_26493,N_24862,N_24484);
xnor U26494 (N_26494,N_24308,N_24964);
xnor U26495 (N_26495,N_24957,N_24651);
or U26496 (N_26496,N_24179,N_25723);
nor U26497 (N_26497,N_24941,N_24741);
nor U26498 (N_26498,N_25173,N_25205);
nand U26499 (N_26499,N_25700,N_25560);
and U26500 (N_26500,N_24042,N_25208);
nand U26501 (N_26501,N_25431,N_25308);
and U26502 (N_26502,N_24209,N_25672);
nor U26503 (N_26503,N_24873,N_24670);
and U26504 (N_26504,N_24953,N_25219);
or U26505 (N_26505,N_24375,N_24360);
or U26506 (N_26506,N_24993,N_24266);
or U26507 (N_26507,N_25457,N_25783);
or U26508 (N_26508,N_24828,N_25110);
and U26509 (N_26509,N_24579,N_25485);
nor U26510 (N_26510,N_24275,N_24303);
xnor U26511 (N_26511,N_24645,N_25421);
and U26512 (N_26512,N_25193,N_25096);
nand U26513 (N_26513,N_24493,N_24012);
nand U26514 (N_26514,N_24568,N_24849);
nor U26515 (N_26515,N_25198,N_25265);
nand U26516 (N_26516,N_25695,N_25718);
nor U26517 (N_26517,N_25099,N_24851);
nand U26518 (N_26518,N_25234,N_24519);
and U26519 (N_26519,N_25520,N_25270);
or U26520 (N_26520,N_25780,N_25568);
nor U26521 (N_26521,N_25546,N_24228);
and U26522 (N_26522,N_24602,N_25344);
and U26523 (N_26523,N_25781,N_25065);
xnor U26524 (N_26524,N_24431,N_24664);
nor U26525 (N_26525,N_24872,N_25195);
nor U26526 (N_26526,N_25113,N_25759);
or U26527 (N_26527,N_24479,N_24766);
and U26528 (N_26528,N_25654,N_24273);
xnor U26529 (N_26529,N_24159,N_24868);
and U26530 (N_26530,N_25359,N_25588);
and U26531 (N_26531,N_25517,N_24820);
nor U26532 (N_26532,N_24637,N_24039);
or U26533 (N_26533,N_25230,N_25894);
and U26534 (N_26534,N_24383,N_25697);
and U26535 (N_26535,N_24365,N_25366);
or U26536 (N_26536,N_24835,N_25155);
nor U26537 (N_26537,N_24793,N_24661);
xnor U26538 (N_26538,N_24405,N_25093);
nand U26539 (N_26539,N_25053,N_24138);
nor U26540 (N_26540,N_25356,N_25439);
and U26541 (N_26541,N_25111,N_24020);
or U26542 (N_26542,N_24910,N_25141);
or U26543 (N_26543,N_24837,N_25720);
and U26544 (N_26544,N_24135,N_25533);
xnor U26545 (N_26545,N_24118,N_24982);
and U26546 (N_26546,N_24738,N_24531);
nand U26547 (N_26547,N_24692,N_25009);
or U26548 (N_26548,N_25599,N_24853);
or U26549 (N_26549,N_24394,N_25102);
xor U26550 (N_26550,N_24966,N_25007);
xnor U26551 (N_26551,N_24105,N_24921);
or U26552 (N_26552,N_25455,N_24331);
and U26553 (N_26553,N_24765,N_24313);
xnor U26554 (N_26554,N_25986,N_25685);
nand U26555 (N_26555,N_25436,N_25084);
nor U26556 (N_26556,N_25760,N_25593);
and U26557 (N_26557,N_24722,N_24436);
xnor U26558 (N_26558,N_25034,N_25804);
or U26559 (N_26559,N_25868,N_24776);
and U26560 (N_26560,N_24403,N_24617);
or U26561 (N_26561,N_25925,N_24750);
and U26562 (N_26562,N_25842,N_24860);
or U26563 (N_26563,N_24640,N_24992);
and U26564 (N_26564,N_25999,N_24124);
xor U26565 (N_26565,N_24101,N_25800);
nand U26566 (N_26566,N_24117,N_25843);
xor U26567 (N_26567,N_25550,N_24696);
or U26568 (N_26568,N_25558,N_24762);
nor U26569 (N_26569,N_24388,N_25349);
or U26570 (N_26570,N_24915,N_25579);
or U26571 (N_26571,N_25063,N_24824);
nand U26572 (N_26572,N_25879,N_25652);
xnor U26573 (N_26573,N_24877,N_25918);
and U26574 (N_26574,N_25756,N_24049);
xnor U26575 (N_26575,N_24854,N_25512);
or U26576 (N_26576,N_25024,N_25690);
nand U26577 (N_26577,N_24911,N_25650);
and U26578 (N_26578,N_25035,N_25526);
or U26579 (N_26579,N_25134,N_24756);
or U26580 (N_26580,N_24352,N_25809);
nor U26581 (N_26581,N_25438,N_25890);
and U26582 (N_26582,N_25426,N_25272);
xor U26583 (N_26583,N_25389,N_24288);
or U26584 (N_26584,N_24262,N_25312);
or U26585 (N_26585,N_24474,N_24603);
and U26586 (N_26586,N_24284,N_25479);
and U26587 (N_26587,N_25491,N_24225);
nand U26588 (N_26588,N_24310,N_25665);
and U26589 (N_26589,N_24289,N_25410);
nor U26590 (N_26590,N_24496,N_25444);
or U26591 (N_26591,N_24797,N_24366);
xnor U26592 (N_26592,N_24316,N_24705);
xnor U26593 (N_26593,N_24068,N_24414);
or U26594 (N_26594,N_24130,N_25185);
xor U26595 (N_26595,N_24945,N_25494);
or U26596 (N_26596,N_24669,N_24028);
nand U26597 (N_26597,N_24064,N_24978);
or U26598 (N_26598,N_25916,N_25527);
nand U26599 (N_26599,N_25888,N_25179);
nor U26600 (N_26600,N_24729,N_25764);
nor U26601 (N_26601,N_24146,N_25183);
and U26602 (N_26602,N_24411,N_25721);
xor U26603 (N_26603,N_25318,N_25734);
xnor U26604 (N_26604,N_25220,N_25078);
and U26605 (N_26605,N_24944,N_25580);
nor U26606 (N_26606,N_24107,N_25201);
or U26607 (N_26607,N_24703,N_25157);
or U26608 (N_26608,N_25834,N_25005);
or U26609 (N_26609,N_24563,N_25350);
nand U26610 (N_26610,N_24050,N_24236);
and U26611 (N_26611,N_25625,N_24200);
and U26612 (N_26612,N_25661,N_24863);
or U26613 (N_26613,N_24008,N_24115);
or U26614 (N_26614,N_24354,N_25707);
or U26615 (N_26615,N_25303,N_24348);
or U26616 (N_26616,N_25567,N_25719);
nor U26617 (N_26617,N_25154,N_25688);
nand U26618 (N_26618,N_25250,N_25818);
or U26619 (N_26619,N_25853,N_24387);
and U26620 (N_26620,N_25342,N_25447);
and U26621 (N_26621,N_24103,N_24575);
or U26622 (N_26622,N_24786,N_24526);
nor U26623 (N_26623,N_24263,N_24987);
nand U26624 (N_26624,N_24894,N_25666);
nor U26625 (N_26625,N_24570,N_25097);
xnor U26626 (N_26626,N_25086,N_25271);
or U26627 (N_26627,N_25627,N_25387);
nand U26628 (N_26628,N_25459,N_24301);
nand U26629 (N_26629,N_24271,N_24205);
and U26630 (N_26630,N_24912,N_25988);
or U26631 (N_26631,N_24329,N_24031);
or U26632 (N_26632,N_24037,N_25467);
or U26633 (N_26633,N_24208,N_24708);
or U26634 (N_26634,N_25474,N_25745);
nor U26635 (N_26635,N_25333,N_24451);
xnor U26636 (N_26636,N_25329,N_25869);
or U26637 (N_26637,N_24239,N_25618);
nor U26638 (N_26638,N_24735,N_24641);
nor U26639 (N_26639,N_24174,N_25612);
nand U26640 (N_26640,N_24907,N_24111);
and U26641 (N_26641,N_25321,N_24241);
xor U26642 (N_26642,N_25813,N_25391);
xnor U26643 (N_26643,N_24812,N_25839);
nor U26644 (N_26644,N_24586,N_25871);
nand U26645 (N_26645,N_25489,N_25801);
nand U26646 (N_26646,N_24572,N_25836);
xor U26647 (N_26647,N_24799,N_25351);
or U26648 (N_26648,N_24999,N_24054);
or U26649 (N_26649,N_25181,N_25233);
or U26650 (N_26650,N_25018,N_24234);
nand U26651 (N_26651,N_24827,N_24761);
nor U26652 (N_26652,N_25068,N_25088);
or U26653 (N_26653,N_25724,N_25037);
and U26654 (N_26654,N_25011,N_25530);
nand U26655 (N_26655,N_25787,N_25982);
xnor U26656 (N_26656,N_25405,N_24152);
and U26657 (N_26657,N_25260,N_24470);
or U26658 (N_26658,N_25094,N_25423);
or U26659 (N_26659,N_25609,N_24649);
and U26660 (N_26660,N_24867,N_25909);
or U26661 (N_26661,N_24198,N_25472);
or U26662 (N_26662,N_24336,N_25583);
nor U26663 (N_26663,N_24203,N_24971);
or U26664 (N_26664,N_25692,N_25514);
xnor U26665 (N_26665,N_24947,N_25252);
nor U26666 (N_26666,N_25257,N_25361);
and U26667 (N_26667,N_25119,N_24075);
nor U26668 (N_26668,N_24668,N_24564);
nor U26669 (N_26669,N_25591,N_24990);
xor U26670 (N_26670,N_25247,N_25981);
nor U26671 (N_26671,N_24033,N_25601);
and U26672 (N_26672,N_24343,N_24090);
nor U26673 (N_26673,N_24972,N_24506);
and U26674 (N_26674,N_25315,N_25776);
or U26675 (N_26675,N_25816,N_24527);
or U26676 (N_26676,N_25914,N_24337);
nor U26677 (N_26677,N_24393,N_25130);
and U26678 (N_26678,N_25915,N_25825);
and U26679 (N_26679,N_25581,N_25254);
and U26680 (N_26680,N_25696,N_25778);
xnor U26681 (N_26681,N_25893,N_24561);
xor U26682 (N_26682,N_25266,N_25069);
or U26683 (N_26683,N_25151,N_24550);
nor U26684 (N_26684,N_25170,N_25267);
and U26685 (N_26685,N_25532,N_25261);
or U26686 (N_26686,N_24710,N_25147);
nor U26687 (N_26687,N_25620,N_25740);
nor U26688 (N_26688,N_25413,N_25525);
nor U26689 (N_26689,N_24687,N_24250);
xor U26690 (N_26690,N_24576,N_25251);
nor U26691 (N_26691,N_24119,N_25453);
and U26692 (N_26692,N_24099,N_24856);
xnor U26693 (N_26693,N_25743,N_25985);
nor U26694 (N_26694,N_24322,N_25945);
nand U26695 (N_26695,N_24889,N_24410);
xnor U26696 (N_26696,N_25095,N_24120);
and U26697 (N_26697,N_25936,N_25091);
nor U26698 (N_26698,N_25729,N_24936);
and U26699 (N_26699,N_24759,N_24939);
and U26700 (N_26700,N_25747,N_24919);
nand U26701 (N_26701,N_24183,N_24265);
nor U26702 (N_26702,N_25735,N_25678);
and U26703 (N_26703,N_24757,N_24753);
or U26704 (N_26704,N_25862,N_24254);
or U26705 (N_26705,N_25997,N_24544);
or U26706 (N_26706,N_24071,N_25706);
and U26707 (N_26707,N_24438,N_24525);
xnor U26708 (N_26708,N_25158,N_24548);
nor U26709 (N_26709,N_24601,N_24490);
or U26710 (N_26710,N_24456,N_24040);
and U26711 (N_26711,N_24719,N_24350);
xnor U26712 (N_26712,N_24726,N_24464);
xnor U26713 (N_26713,N_25791,N_24475);
nor U26714 (N_26714,N_24590,N_25676);
or U26715 (N_26715,N_24836,N_25948);
nor U26716 (N_26716,N_25046,N_24846);
xor U26717 (N_26717,N_25039,N_25397);
nor U26718 (N_26718,N_24983,N_24529);
nor U26719 (N_26719,N_24058,N_24353);
nor U26720 (N_26720,N_25866,N_24792);
or U26721 (N_26721,N_25460,N_24632);
and U26722 (N_26722,N_24823,N_25304);
xnor U26723 (N_26723,N_24620,N_24379);
nand U26724 (N_26724,N_24962,N_24859);
nand U26725 (N_26725,N_25929,N_24566);
and U26726 (N_26726,N_25160,N_25807);
nand U26727 (N_26727,N_24424,N_24956);
or U26728 (N_26728,N_25865,N_25066);
or U26729 (N_26729,N_25732,N_25013);
or U26730 (N_26730,N_25516,N_25435);
and U26731 (N_26731,N_25365,N_24495);
or U26732 (N_26732,N_24504,N_24346);
nor U26733 (N_26733,N_24291,N_25501);
nand U26734 (N_26734,N_25796,N_24946);
nand U26735 (N_26735,N_24583,N_24515);
nand U26736 (N_26736,N_24312,N_24333);
nand U26737 (N_26737,N_24327,N_24634);
nor U26738 (N_26738,N_25870,N_25396);
xnor U26739 (N_26739,N_24340,N_24001);
or U26740 (N_26740,N_24514,N_24357);
or U26741 (N_26741,N_25180,N_24149);
xnor U26742 (N_26742,N_24594,N_25502);
nor U26743 (N_26743,N_25148,N_25708);
xor U26744 (N_26744,N_25832,N_24123);
nand U26745 (N_26745,N_24577,N_25279);
or U26746 (N_26746,N_24830,N_24019);
or U26747 (N_26747,N_25660,N_24740);
nor U26748 (N_26748,N_25306,N_25117);
and U26749 (N_26749,N_24518,N_24736);
nor U26750 (N_26750,N_24374,N_24848);
or U26751 (N_26751,N_25070,N_24516);
nand U26752 (N_26752,N_24142,N_25507);
nand U26753 (N_26753,N_24948,N_25121);
xor U26754 (N_26754,N_24185,N_25463);
and U26755 (N_26755,N_24988,N_24542);
and U26756 (N_26756,N_24800,N_24481);
or U26757 (N_26757,N_25662,N_24580);
and U26758 (N_26758,N_25275,N_25437);
nand U26759 (N_26759,N_24896,N_25808);
nor U26760 (N_26760,N_25192,N_24127);
xor U26761 (N_26761,N_25694,N_25047);
nor U26762 (N_26762,N_24829,N_24334);
nor U26763 (N_26763,N_24397,N_25317);
nor U26764 (N_26764,N_24015,N_24044);
and U26765 (N_26765,N_24447,N_24773);
and U26766 (N_26766,N_25285,N_24461);
nor U26767 (N_26767,N_24706,N_25919);
nor U26768 (N_26768,N_25458,N_24341);
or U26769 (N_26769,N_24909,N_25244);
nor U26770 (N_26770,N_24642,N_25623);
xnor U26771 (N_26771,N_24961,N_25159);
nand U26772 (N_26772,N_25702,N_24455);
or U26773 (N_26773,N_24774,N_24041);
nand U26774 (N_26774,N_24404,N_24184);
and U26775 (N_26775,N_25574,N_24615);
and U26776 (N_26776,N_25848,N_24221);
xor U26777 (N_26777,N_25212,N_25683);
and U26778 (N_26778,N_25642,N_24815);
and U26779 (N_26779,N_25761,N_24609);
and U26780 (N_26780,N_25253,N_24888);
nand U26781 (N_26781,N_24639,N_25090);
or U26782 (N_26782,N_25030,N_25674);
and U26783 (N_26783,N_25876,N_25833);
nand U26784 (N_26784,N_25822,N_24076);
xor U26785 (N_26785,N_24067,N_25476);
xnor U26786 (N_26786,N_24476,N_24952);
and U26787 (N_26787,N_25710,N_25884);
or U26788 (N_26788,N_24891,N_24596);
or U26789 (N_26789,N_25750,N_24081);
nor U26790 (N_26790,N_24151,N_24156);
nand U26791 (N_26791,N_24415,N_25990);
or U26792 (N_26792,N_24985,N_24553);
or U26793 (N_26793,N_25713,N_25200);
or U26794 (N_26794,N_24201,N_24898);
xnor U26795 (N_26795,N_24574,N_25071);
nor U26796 (N_26796,N_24802,N_25742);
nor U26797 (N_26797,N_25995,N_25335);
nor U26798 (N_26798,N_25424,N_24677);
nand U26799 (N_26799,N_24622,N_24249);
nand U26800 (N_26800,N_24095,N_25703);
or U26801 (N_26801,N_24611,N_25673);
nor U26802 (N_26802,N_25114,N_24172);
nor U26803 (N_26803,N_25082,N_24528);
xnor U26804 (N_26804,N_25231,N_24287);
xor U26805 (N_26805,N_24441,N_24055);
and U26806 (N_26806,N_24299,N_24283);
xor U26807 (N_26807,N_25930,N_24676);
nor U26808 (N_26808,N_25604,N_25539);
and U26809 (N_26809,N_24373,N_24689);
xnor U26810 (N_26810,N_24991,N_24545);
xor U26811 (N_26811,N_25923,N_25619);
and U26812 (N_26812,N_24950,N_25433);
and U26813 (N_26813,N_24751,N_25542);
and U26814 (N_26814,N_25057,N_25290);
xor U26815 (N_26815,N_24695,N_25188);
xor U26816 (N_26816,N_24400,N_24809);
nand U26817 (N_26817,N_25314,N_24994);
xnor U26818 (N_26818,N_25461,N_25002);
nand U26819 (N_26819,N_25123,N_25124);
and U26820 (N_26820,N_25920,N_24969);
nand U26821 (N_26821,N_24694,N_25129);
nor U26822 (N_26822,N_25578,N_25364);
nor U26823 (N_26823,N_25555,N_24086);
nor U26824 (N_26824,N_24021,N_25967);
xor U26825 (N_26825,N_24672,N_24285);
xnor U26826 (N_26826,N_24998,N_24243);
xor U26827 (N_26827,N_25983,N_25420);
xor U26828 (N_26828,N_24323,N_24128);
nor U26829 (N_26829,N_25089,N_25744);
nand U26830 (N_26830,N_24683,N_24102);
nand U26831 (N_26831,N_25797,N_25175);
nor U26832 (N_26832,N_24604,N_25704);
or U26833 (N_26833,N_25637,N_25511);
and U26834 (N_26834,N_24218,N_25769);
xnor U26835 (N_26835,N_24213,N_25384);
or U26836 (N_26836,N_24725,N_25452);
or U26837 (N_26837,N_25109,N_24224);
and U26838 (N_26838,N_24114,N_25305);
or U26839 (N_26839,N_25296,N_24571);
nand U26840 (N_26840,N_25469,N_25017);
xor U26841 (N_26841,N_24121,N_24477);
or U26842 (N_26842,N_24488,N_25573);
nor U26843 (N_26843,N_25446,N_24923);
nor U26844 (N_26844,N_25417,N_25381);
or U26845 (N_26845,N_24727,N_24416);
nand U26846 (N_26846,N_24423,N_24248);
or U26847 (N_26847,N_24108,N_24501);
xnor U26848 (N_26848,N_25881,N_25731);
nor U26849 (N_26849,N_25675,N_24618);
and U26850 (N_26850,N_24029,N_25196);
or U26851 (N_26851,N_25085,N_24532);
nor U26852 (N_26852,N_24734,N_25774);
xnor U26853 (N_26853,N_25136,N_25358);
nand U26854 (N_26854,N_24300,N_24193);
nand U26855 (N_26855,N_24190,N_24845);
xnor U26856 (N_26856,N_24630,N_24351);
nor U26857 (N_26857,N_25120,N_25631);
xnor U26858 (N_26858,N_25628,N_25794);
nor U26859 (N_26859,N_24871,N_25687);
or U26860 (N_26860,N_25908,N_25885);
and U26861 (N_26861,N_24472,N_25370);
nand U26862 (N_26862,N_25298,N_24591);
nor U26863 (N_26863,N_24469,N_25669);
nand U26864 (N_26864,N_25050,N_24098);
nor U26865 (N_26865,N_25137,N_24073);
or U26866 (N_26866,N_24085,N_25138);
and U26867 (N_26867,N_24667,N_24502);
or U26868 (N_26868,N_24043,N_25466);
xnor U26869 (N_26869,N_24051,N_25412);
nor U26870 (N_26870,N_24180,N_25153);
nand U26871 (N_26871,N_24658,N_25190);
nor U26872 (N_26872,N_24555,N_24884);
nand U26873 (N_26873,N_24259,N_25098);
xnor U26874 (N_26874,N_25585,N_25048);
xnor U26875 (N_26875,N_24628,N_24109);
or U26876 (N_26876,N_24968,N_25616);
nor U26877 (N_26877,N_24445,N_25991);
and U26878 (N_26878,N_24821,N_24679);
xnor U26879 (N_26879,N_24290,N_24380);
nor U26880 (N_26880,N_25103,N_24245);
nor U26881 (N_26881,N_24974,N_24789);
and U26882 (N_26882,N_24977,N_25430);
or U26883 (N_26883,N_24801,N_25127);
nor U26884 (N_26884,N_25882,N_25677);
nand U26885 (N_26885,N_25214,N_24347);
nand U26886 (N_26886,N_25324,N_24712);
xor U26887 (N_26887,N_24100,N_24589);
and U26888 (N_26888,N_24643,N_25956);
nor U26889 (N_26889,N_24279,N_25118);
nand U26890 (N_26890,N_25824,N_24614);
nor U26891 (N_26891,N_24539,N_25828);
xnor U26892 (N_26892,N_24558,N_24409);
nor U26893 (N_26893,N_24500,N_25156);
xnor U26894 (N_26894,N_25211,N_24685);
nor U26895 (N_26895,N_24443,N_24349);
or U26896 (N_26896,N_25812,N_25935);
nor U26897 (N_26897,N_25582,N_25670);
xor U26898 (N_26898,N_25912,N_24160);
and U26899 (N_26899,N_24523,N_24858);
or U26900 (N_26900,N_25286,N_25348);
nand U26901 (N_26901,N_25906,N_24814);
xnor U26902 (N_26902,N_24219,N_24965);
or U26903 (N_26903,N_25943,N_25684);
nand U26904 (N_26904,N_25164,N_24057);
or U26905 (N_26905,N_25471,N_25235);
and U26906 (N_26906,N_24967,N_25962);
or U26907 (N_26907,N_25626,N_25857);
or U26908 (N_26908,N_25771,N_24048);
nor U26909 (N_26909,N_24813,N_25074);
or U26910 (N_26910,N_25605,N_25465);
or U26911 (N_26911,N_25940,N_24384);
and U26912 (N_26912,N_25184,N_25161);
and U26913 (N_26913,N_24885,N_25171);
xnor U26914 (N_26914,N_25434,N_25657);
or U26915 (N_26915,N_24171,N_24852);
nand U26916 (N_26916,N_24482,N_25887);
nand U26917 (N_26917,N_24929,N_25576);
or U26918 (N_26918,N_25788,N_25994);
and U26919 (N_26919,N_25336,N_25531);
nand U26920 (N_26920,N_25952,N_24434);
nand U26921 (N_26921,N_25470,N_24702);
xnor U26922 (N_26922,N_24024,N_25534);
nand U26923 (N_26923,N_25937,N_25548);
or U26924 (N_26924,N_25564,N_25900);
and U26925 (N_26925,N_25811,N_24855);
or U26926 (N_26926,N_24684,N_24417);
nand U26927 (N_26927,N_25845,N_24660);
xor U26928 (N_26928,N_24025,N_24339);
and U26929 (N_26929,N_25725,N_24463);
nor U26930 (N_26930,N_25227,N_24747);
or U26931 (N_26931,N_24782,N_25741);
xnor U26932 (N_26932,N_24780,N_24647);
and U26933 (N_26933,N_25504,N_25399);
nand U26934 (N_26934,N_24593,N_24280);
or U26935 (N_26935,N_24335,N_24027);
or U26936 (N_26936,N_25867,N_25497);
nand U26937 (N_26937,N_24161,N_24629);
xor U26938 (N_26938,N_25840,N_25377);
nand U26939 (N_26939,N_24599,N_24927);
or U26940 (N_26940,N_24182,N_25226);
or U26941 (N_26941,N_25973,N_24237);
nor U26942 (N_26942,N_24215,N_24196);
or U26943 (N_26943,N_24282,N_24129);
nor U26944 (N_26944,N_24440,N_25224);
or U26945 (N_26945,N_25649,N_24744);
or U26946 (N_26946,N_25841,N_24822);
nand U26947 (N_26947,N_24654,N_24924);
or U26948 (N_26948,N_25301,N_24302);
nor U26949 (N_26949,N_24344,N_24465);
nor U26950 (N_26950,N_24731,N_25087);
nor U26951 (N_26951,N_25519,N_24674);
or U26952 (N_26952,N_24318,N_25681);
and U26953 (N_26953,N_25478,N_25851);
or U26954 (N_26954,N_24711,N_25854);
nor U26955 (N_26955,N_25105,N_24382);
nor U26956 (N_26956,N_24876,N_25177);
or U26957 (N_26957,N_24444,N_24935);
or U26958 (N_26958,N_25045,N_24861);
nor U26959 (N_26959,N_25538,N_25559);
nand U26960 (N_26960,N_25316,N_25341);
xor U26961 (N_26961,N_24538,N_24816);
nor U26962 (N_26962,N_25056,N_25859);
nand U26963 (N_26963,N_25052,N_25004);
xor U26964 (N_26964,N_24070,N_25762);
or U26965 (N_26965,N_25080,N_24748);
nor U26966 (N_26966,N_25634,N_25221);
xor U26967 (N_26967,N_25443,N_25204);
nand U26968 (N_26968,N_24026,N_24157);
or U26969 (N_26969,N_24315,N_24131);
nand U26970 (N_26970,N_24255,N_25276);
nand U26971 (N_26971,N_24144,N_24483);
nand U26972 (N_26972,N_25569,N_25820);
xnor U26973 (N_26973,N_24605,N_24787);
or U26974 (N_26974,N_24937,N_25932);
xor U26975 (N_26975,N_24616,N_24767);
or U26976 (N_26976,N_24398,N_24061);
nand U26977 (N_26977,N_25803,N_24619);
or U26978 (N_26978,N_24743,N_25972);
xnor U26979 (N_26979,N_24281,N_24588);
or U26980 (N_26980,N_24728,N_24522);
nand U26981 (N_26981,N_24429,N_25827);
or U26982 (N_26982,N_25144,N_24573);
xnor U26983 (N_26983,N_24223,N_25101);
or U26984 (N_26984,N_24721,N_25992);
or U26985 (N_26985,N_24233,N_24253);
xnor U26986 (N_26986,N_24449,N_24420);
nor U26987 (N_26987,N_25968,N_24903);
nor U26988 (N_26988,N_25189,N_25535);
or U26989 (N_26989,N_25537,N_25664);
or U26990 (N_26990,N_25877,N_25347);
xor U26991 (N_26991,N_25611,N_25025);
xor U26992 (N_26992,N_24227,N_25132);
xnor U26993 (N_26993,N_24648,N_24091);
and U26994 (N_26994,N_24270,N_25263);
nand U26995 (N_26995,N_24094,N_25225);
xnor U26996 (N_26996,N_25280,N_24162);
nand U26997 (N_26997,N_25645,N_25959);
nor U26998 (N_26998,N_24749,N_25541);
and U26999 (N_26999,N_25793,N_25428);
and U27000 (N_27000,N_24518,N_24238);
and U27001 (N_27001,N_24436,N_24883);
and U27002 (N_27002,N_24469,N_24668);
xnor U27003 (N_27003,N_25100,N_24658);
xnor U27004 (N_27004,N_24768,N_25387);
nand U27005 (N_27005,N_24830,N_24124);
or U27006 (N_27006,N_24027,N_24561);
or U27007 (N_27007,N_24415,N_25694);
nand U27008 (N_27008,N_25119,N_24725);
and U27009 (N_27009,N_24155,N_24751);
and U27010 (N_27010,N_25698,N_24942);
and U27011 (N_27011,N_24208,N_25183);
xor U27012 (N_27012,N_24214,N_24698);
or U27013 (N_27013,N_24622,N_24057);
or U27014 (N_27014,N_24788,N_24980);
or U27015 (N_27015,N_24397,N_24251);
and U27016 (N_27016,N_24521,N_25981);
xnor U27017 (N_27017,N_24565,N_24573);
or U27018 (N_27018,N_25999,N_24391);
xor U27019 (N_27019,N_24598,N_25741);
or U27020 (N_27020,N_25281,N_25663);
xnor U27021 (N_27021,N_24734,N_24729);
or U27022 (N_27022,N_25622,N_25543);
xor U27023 (N_27023,N_24876,N_24847);
nor U27024 (N_27024,N_25030,N_24320);
or U27025 (N_27025,N_25423,N_25257);
or U27026 (N_27026,N_24546,N_25680);
xor U27027 (N_27027,N_24631,N_24874);
or U27028 (N_27028,N_25875,N_24569);
or U27029 (N_27029,N_24946,N_24965);
nor U27030 (N_27030,N_25412,N_24757);
nor U27031 (N_27031,N_25526,N_25905);
or U27032 (N_27032,N_24501,N_24150);
xor U27033 (N_27033,N_25988,N_24489);
and U27034 (N_27034,N_25871,N_24622);
nor U27035 (N_27035,N_25280,N_25775);
nand U27036 (N_27036,N_24632,N_25588);
nand U27037 (N_27037,N_25002,N_24161);
or U27038 (N_27038,N_25581,N_24325);
nor U27039 (N_27039,N_25212,N_25425);
nor U27040 (N_27040,N_25321,N_25464);
xor U27041 (N_27041,N_25906,N_24061);
xnor U27042 (N_27042,N_25398,N_24354);
xnor U27043 (N_27043,N_24106,N_25405);
xor U27044 (N_27044,N_25974,N_25170);
or U27045 (N_27045,N_24850,N_24158);
xor U27046 (N_27046,N_24187,N_25157);
nand U27047 (N_27047,N_24005,N_25525);
and U27048 (N_27048,N_25592,N_25415);
or U27049 (N_27049,N_25047,N_25886);
nor U27050 (N_27050,N_24819,N_25762);
or U27051 (N_27051,N_25906,N_25625);
and U27052 (N_27052,N_25032,N_24250);
or U27053 (N_27053,N_24037,N_24151);
xor U27054 (N_27054,N_25862,N_25155);
and U27055 (N_27055,N_24982,N_25692);
nand U27056 (N_27056,N_24553,N_25831);
and U27057 (N_27057,N_24812,N_24081);
or U27058 (N_27058,N_25594,N_24567);
and U27059 (N_27059,N_25124,N_24183);
xor U27060 (N_27060,N_25083,N_24545);
and U27061 (N_27061,N_25020,N_25313);
xnor U27062 (N_27062,N_25714,N_24775);
nor U27063 (N_27063,N_25388,N_25248);
and U27064 (N_27064,N_25850,N_25097);
xor U27065 (N_27065,N_24755,N_25114);
and U27066 (N_27066,N_24624,N_25089);
or U27067 (N_27067,N_25350,N_24304);
nor U27068 (N_27068,N_24918,N_25465);
xor U27069 (N_27069,N_24443,N_25769);
xor U27070 (N_27070,N_25943,N_25733);
nand U27071 (N_27071,N_24080,N_25727);
xnor U27072 (N_27072,N_24295,N_24374);
xnor U27073 (N_27073,N_25395,N_24894);
and U27074 (N_27074,N_24312,N_25819);
nor U27075 (N_27075,N_25851,N_24775);
or U27076 (N_27076,N_25331,N_25243);
xnor U27077 (N_27077,N_25345,N_24534);
and U27078 (N_27078,N_24965,N_25569);
and U27079 (N_27079,N_25374,N_25107);
nor U27080 (N_27080,N_25187,N_24959);
or U27081 (N_27081,N_25550,N_25049);
nor U27082 (N_27082,N_25807,N_25352);
or U27083 (N_27083,N_24916,N_24664);
or U27084 (N_27084,N_25034,N_25508);
nor U27085 (N_27085,N_24451,N_24963);
nand U27086 (N_27086,N_25743,N_25039);
nor U27087 (N_27087,N_25603,N_24015);
xor U27088 (N_27088,N_24514,N_24013);
and U27089 (N_27089,N_24875,N_24455);
or U27090 (N_27090,N_24297,N_25800);
nand U27091 (N_27091,N_25991,N_24394);
xor U27092 (N_27092,N_25233,N_25505);
or U27093 (N_27093,N_25253,N_25381);
or U27094 (N_27094,N_24089,N_25329);
nand U27095 (N_27095,N_24728,N_25207);
xor U27096 (N_27096,N_24802,N_25722);
nand U27097 (N_27097,N_25017,N_25398);
and U27098 (N_27098,N_25455,N_24733);
or U27099 (N_27099,N_24471,N_25072);
and U27100 (N_27100,N_24585,N_25212);
or U27101 (N_27101,N_25458,N_24360);
or U27102 (N_27102,N_24454,N_25895);
or U27103 (N_27103,N_24126,N_25675);
nand U27104 (N_27104,N_24352,N_25134);
nor U27105 (N_27105,N_25967,N_24627);
nor U27106 (N_27106,N_24230,N_25476);
xor U27107 (N_27107,N_25316,N_24649);
nor U27108 (N_27108,N_25157,N_25487);
or U27109 (N_27109,N_24471,N_25634);
xnor U27110 (N_27110,N_24336,N_24343);
nand U27111 (N_27111,N_24991,N_25238);
or U27112 (N_27112,N_25572,N_25466);
nand U27113 (N_27113,N_25443,N_24088);
and U27114 (N_27114,N_25330,N_25101);
nor U27115 (N_27115,N_25014,N_25266);
xnor U27116 (N_27116,N_24180,N_24432);
or U27117 (N_27117,N_25053,N_25800);
nand U27118 (N_27118,N_25820,N_25665);
or U27119 (N_27119,N_25141,N_24154);
nand U27120 (N_27120,N_24973,N_24281);
nor U27121 (N_27121,N_25524,N_25019);
or U27122 (N_27122,N_24249,N_25704);
xnor U27123 (N_27123,N_25247,N_25119);
xor U27124 (N_27124,N_24689,N_25280);
nor U27125 (N_27125,N_24534,N_25721);
and U27126 (N_27126,N_24175,N_24990);
nor U27127 (N_27127,N_24196,N_24507);
and U27128 (N_27128,N_24021,N_24374);
nor U27129 (N_27129,N_24834,N_25215);
nor U27130 (N_27130,N_25901,N_24556);
and U27131 (N_27131,N_24967,N_24455);
and U27132 (N_27132,N_24660,N_25143);
and U27133 (N_27133,N_25977,N_24136);
and U27134 (N_27134,N_24551,N_24154);
and U27135 (N_27135,N_24864,N_25877);
and U27136 (N_27136,N_24659,N_24880);
xor U27137 (N_27137,N_25085,N_24304);
nor U27138 (N_27138,N_24893,N_25334);
or U27139 (N_27139,N_24675,N_25343);
and U27140 (N_27140,N_24354,N_24855);
xnor U27141 (N_27141,N_25697,N_25213);
and U27142 (N_27142,N_24269,N_24391);
nand U27143 (N_27143,N_25347,N_25480);
nor U27144 (N_27144,N_25031,N_24950);
nor U27145 (N_27145,N_24848,N_25629);
and U27146 (N_27146,N_25685,N_25407);
xor U27147 (N_27147,N_25839,N_24626);
nand U27148 (N_27148,N_24538,N_25274);
or U27149 (N_27149,N_25461,N_24681);
xnor U27150 (N_27150,N_24166,N_25794);
and U27151 (N_27151,N_25273,N_25137);
nand U27152 (N_27152,N_24510,N_24390);
xnor U27153 (N_27153,N_25667,N_24107);
and U27154 (N_27154,N_25822,N_24740);
nand U27155 (N_27155,N_25764,N_25177);
nor U27156 (N_27156,N_24654,N_24512);
or U27157 (N_27157,N_24213,N_25422);
xnor U27158 (N_27158,N_25900,N_24577);
nor U27159 (N_27159,N_24759,N_24794);
and U27160 (N_27160,N_25502,N_25523);
nand U27161 (N_27161,N_24237,N_24722);
nor U27162 (N_27162,N_25819,N_25405);
or U27163 (N_27163,N_24286,N_24841);
or U27164 (N_27164,N_25635,N_24772);
xor U27165 (N_27165,N_25987,N_25844);
nand U27166 (N_27166,N_25438,N_25073);
and U27167 (N_27167,N_25653,N_25638);
xor U27168 (N_27168,N_24528,N_24302);
xnor U27169 (N_27169,N_25737,N_24375);
xor U27170 (N_27170,N_25516,N_24343);
nor U27171 (N_27171,N_24893,N_24304);
or U27172 (N_27172,N_25638,N_24184);
and U27173 (N_27173,N_24360,N_25638);
xnor U27174 (N_27174,N_24258,N_25363);
nor U27175 (N_27175,N_24113,N_24122);
or U27176 (N_27176,N_25440,N_25569);
and U27177 (N_27177,N_25123,N_25869);
or U27178 (N_27178,N_25310,N_25223);
or U27179 (N_27179,N_24899,N_24431);
or U27180 (N_27180,N_25851,N_25668);
xor U27181 (N_27181,N_25164,N_24593);
nor U27182 (N_27182,N_24520,N_25968);
xor U27183 (N_27183,N_24328,N_25930);
and U27184 (N_27184,N_25317,N_25982);
or U27185 (N_27185,N_24021,N_24859);
or U27186 (N_27186,N_24891,N_25686);
nor U27187 (N_27187,N_25149,N_25270);
nor U27188 (N_27188,N_25981,N_25970);
or U27189 (N_27189,N_25091,N_25202);
and U27190 (N_27190,N_25429,N_24867);
and U27191 (N_27191,N_24517,N_25624);
or U27192 (N_27192,N_25915,N_24240);
or U27193 (N_27193,N_24658,N_25895);
nand U27194 (N_27194,N_24142,N_24339);
and U27195 (N_27195,N_24876,N_25700);
or U27196 (N_27196,N_24620,N_25157);
and U27197 (N_27197,N_24939,N_25557);
nor U27198 (N_27198,N_25625,N_25040);
nand U27199 (N_27199,N_24570,N_24759);
nor U27200 (N_27200,N_25983,N_24363);
nor U27201 (N_27201,N_25705,N_25787);
and U27202 (N_27202,N_25570,N_24362);
or U27203 (N_27203,N_25005,N_25353);
xor U27204 (N_27204,N_24216,N_25014);
or U27205 (N_27205,N_24003,N_25762);
nand U27206 (N_27206,N_24888,N_24360);
nand U27207 (N_27207,N_24363,N_24318);
or U27208 (N_27208,N_25052,N_25633);
nor U27209 (N_27209,N_24140,N_24021);
nor U27210 (N_27210,N_24356,N_25497);
or U27211 (N_27211,N_25914,N_25318);
xor U27212 (N_27212,N_24587,N_25981);
nor U27213 (N_27213,N_24669,N_24457);
nand U27214 (N_27214,N_24820,N_24135);
nand U27215 (N_27215,N_25403,N_25467);
or U27216 (N_27216,N_24550,N_24113);
or U27217 (N_27217,N_24036,N_24516);
nand U27218 (N_27218,N_25306,N_25180);
xor U27219 (N_27219,N_25568,N_24350);
nor U27220 (N_27220,N_24227,N_25422);
and U27221 (N_27221,N_25599,N_24528);
nand U27222 (N_27222,N_25642,N_25024);
xnor U27223 (N_27223,N_24935,N_25569);
or U27224 (N_27224,N_25868,N_24321);
and U27225 (N_27225,N_25022,N_25463);
xnor U27226 (N_27226,N_25252,N_25119);
and U27227 (N_27227,N_24357,N_24384);
or U27228 (N_27228,N_25472,N_24558);
nor U27229 (N_27229,N_25692,N_25347);
nand U27230 (N_27230,N_25287,N_25590);
nor U27231 (N_27231,N_24391,N_24041);
nor U27232 (N_27232,N_25748,N_25129);
xnor U27233 (N_27233,N_24644,N_24474);
and U27234 (N_27234,N_25876,N_24563);
and U27235 (N_27235,N_25104,N_25099);
xor U27236 (N_27236,N_24195,N_25720);
nor U27237 (N_27237,N_25177,N_25660);
nor U27238 (N_27238,N_25165,N_25196);
and U27239 (N_27239,N_25296,N_24470);
or U27240 (N_27240,N_24502,N_24361);
or U27241 (N_27241,N_25692,N_25666);
xnor U27242 (N_27242,N_25956,N_25724);
nor U27243 (N_27243,N_24162,N_25586);
and U27244 (N_27244,N_25499,N_25767);
nor U27245 (N_27245,N_25979,N_24699);
xnor U27246 (N_27246,N_24650,N_25582);
and U27247 (N_27247,N_24217,N_24158);
or U27248 (N_27248,N_24713,N_24024);
nor U27249 (N_27249,N_24451,N_25667);
or U27250 (N_27250,N_24621,N_25929);
nor U27251 (N_27251,N_25428,N_24561);
nor U27252 (N_27252,N_25459,N_25220);
and U27253 (N_27253,N_25315,N_25188);
nand U27254 (N_27254,N_24386,N_25375);
or U27255 (N_27255,N_25686,N_24790);
nor U27256 (N_27256,N_25747,N_25142);
nor U27257 (N_27257,N_25951,N_24883);
and U27258 (N_27258,N_25994,N_24891);
and U27259 (N_27259,N_24086,N_24595);
or U27260 (N_27260,N_24416,N_24991);
xor U27261 (N_27261,N_25800,N_25188);
xnor U27262 (N_27262,N_25854,N_25284);
and U27263 (N_27263,N_24478,N_24090);
xnor U27264 (N_27264,N_24561,N_25265);
or U27265 (N_27265,N_25433,N_25209);
nand U27266 (N_27266,N_24007,N_24138);
or U27267 (N_27267,N_25949,N_25212);
nand U27268 (N_27268,N_24321,N_25764);
or U27269 (N_27269,N_25926,N_25948);
nor U27270 (N_27270,N_24119,N_24529);
and U27271 (N_27271,N_25204,N_25554);
nand U27272 (N_27272,N_24262,N_24110);
nor U27273 (N_27273,N_24526,N_24135);
or U27274 (N_27274,N_25647,N_24545);
nand U27275 (N_27275,N_25258,N_24646);
or U27276 (N_27276,N_24179,N_24993);
nand U27277 (N_27277,N_25723,N_25808);
and U27278 (N_27278,N_25520,N_24940);
nand U27279 (N_27279,N_24579,N_24873);
nor U27280 (N_27280,N_24012,N_25365);
xor U27281 (N_27281,N_25571,N_24395);
xor U27282 (N_27282,N_25673,N_25215);
xnor U27283 (N_27283,N_24493,N_25077);
nand U27284 (N_27284,N_24142,N_24227);
nand U27285 (N_27285,N_24411,N_24008);
xnor U27286 (N_27286,N_24857,N_24730);
or U27287 (N_27287,N_24641,N_24354);
or U27288 (N_27288,N_25321,N_24570);
nand U27289 (N_27289,N_24587,N_25455);
xnor U27290 (N_27290,N_24384,N_24326);
nand U27291 (N_27291,N_25334,N_25543);
nor U27292 (N_27292,N_25985,N_25225);
nor U27293 (N_27293,N_25291,N_24403);
xnor U27294 (N_27294,N_24479,N_24881);
xor U27295 (N_27295,N_24081,N_25542);
xor U27296 (N_27296,N_25709,N_24107);
nand U27297 (N_27297,N_25712,N_25277);
and U27298 (N_27298,N_25906,N_24629);
xnor U27299 (N_27299,N_24232,N_24123);
or U27300 (N_27300,N_24922,N_25188);
nand U27301 (N_27301,N_24177,N_24481);
and U27302 (N_27302,N_25027,N_25333);
or U27303 (N_27303,N_24394,N_25202);
or U27304 (N_27304,N_25976,N_25585);
xnor U27305 (N_27305,N_25943,N_24237);
or U27306 (N_27306,N_25691,N_25184);
xnor U27307 (N_27307,N_25475,N_24681);
nor U27308 (N_27308,N_25670,N_25855);
xor U27309 (N_27309,N_24495,N_25339);
or U27310 (N_27310,N_25365,N_24085);
or U27311 (N_27311,N_25261,N_24824);
nor U27312 (N_27312,N_24986,N_24565);
nand U27313 (N_27313,N_25339,N_25763);
and U27314 (N_27314,N_25932,N_24290);
or U27315 (N_27315,N_25372,N_24581);
or U27316 (N_27316,N_24013,N_24268);
nor U27317 (N_27317,N_24643,N_25128);
or U27318 (N_27318,N_25787,N_24191);
nor U27319 (N_27319,N_24383,N_24551);
nor U27320 (N_27320,N_24148,N_25485);
or U27321 (N_27321,N_24992,N_24331);
xor U27322 (N_27322,N_24377,N_25033);
and U27323 (N_27323,N_25611,N_25004);
and U27324 (N_27324,N_25901,N_25321);
nor U27325 (N_27325,N_25470,N_25278);
nand U27326 (N_27326,N_25986,N_25394);
or U27327 (N_27327,N_24861,N_25839);
nor U27328 (N_27328,N_25607,N_25636);
nor U27329 (N_27329,N_24559,N_24801);
and U27330 (N_27330,N_25001,N_24566);
nor U27331 (N_27331,N_24088,N_24618);
xor U27332 (N_27332,N_24672,N_24914);
nand U27333 (N_27333,N_25731,N_25649);
or U27334 (N_27334,N_25823,N_25894);
nand U27335 (N_27335,N_24936,N_25231);
and U27336 (N_27336,N_25470,N_25999);
nand U27337 (N_27337,N_25075,N_24360);
or U27338 (N_27338,N_25693,N_25458);
or U27339 (N_27339,N_25618,N_25508);
and U27340 (N_27340,N_24663,N_25904);
or U27341 (N_27341,N_25959,N_25437);
nor U27342 (N_27342,N_25988,N_24254);
or U27343 (N_27343,N_24392,N_25981);
or U27344 (N_27344,N_25613,N_25764);
nand U27345 (N_27345,N_25418,N_24081);
or U27346 (N_27346,N_25055,N_24544);
xor U27347 (N_27347,N_25548,N_24274);
and U27348 (N_27348,N_24547,N_25680);
and U27349 (N_27349,N_24847,N_25468);
nand U27350 (N_27350,N_25244,N_25249);
xnor U27351 (N_27351,N_25483,N_25706);
nand U27352 (N_27352,N_25943,N_25179);
and U27353 (N_27353,N_24941,N_24143);
or U27354 (N_27354,N_24739,N_25401);
nor U27355 (N_27355,N_24395,N_24559);
nand U27356 (N_27356,N_24790,N_25607);
xor U27357 (N_27357,N_25919,N_25894);
or U27358 (N_27358,N_25897,N_25297);
or U27359 (N_27359,N_25489,N_25680);
xor U27360 (N_27360,N_25562,N_24493);
xor U27361 (N_27361,N_25779,N_24648);
nand U27362 (N_27362,N_25677,N_25543);
nor U27363 (N_27363,N_25895,N_25289);
nor U27364 (N_27364,N_24607,N_25668);
nor U27365 (N_27365,N_25806,N_24929);
or U27366 (N_27366,N_25599,N_24038);
xor U27367 (N_27367,N_25500,N_24041);
xnor U27368 (N_27368,N_25108,N_24564);
xnor U27369 (N_27369,N_24277,N_25892);
nor U27370 (N_27370,N_25512,N_24293);
xor U27371 (N_27371,N_25092,N_24148);
and U27372 (N_27372,N_24780,N_25837);
xnor U27373 (N_27373,N_24817,N_24830);
nand U27374 (N_27374,N_25075,N_25254);
xnor U27375 (N_27375,N_25414,N_25995);
and U27376 (N_27376,N_24935,N_25304);
nor U27377 (N_27377,N_24637,N_24166);
nand U27378 (N_27378,N_24392,N_24715);
nor U27379 (N_27379,N_25695,N_24054);
and U27380 (N_27380,N_25432,N_25527);
nand U27381 (N_27381,N_25141,N_25360);
xor U27382 (N_27382,N_24425,N_24054);
xor U27383 (N_27383,N_25426,N_24042);
and U27384 (N_27384,N_24972,N_25508);
or U27385 (N_27385,N_24159,N_25670);
and U27386 (N_27386,N_25397,N_25062);
and U27387 (N_27387,N_24063,N_25543);
xor U27388 (N_27388,N_24190,N_24392);
xnor U27389 (N_27389,N_24091,N_24464);
and U27390 (N_27390,N_24521,N_25445);
nand U27391 (N_27391,N_25603,N_24951);
nand U27392 (N_27392,N_24317,N_24497);
nor U27393 (N_27393,N_25624,N_25956);
xnor U27394 (N_27394,N_24411,N_25188);
nand U27395 (N_27395,N_24118,N_25929);
or U27396 (N_27396,N_24170,N_24366);
xnor U27397 (N_27397,N_25315,N_24032);
xnor U27398 (N_27398,N_24682,N_24386);
and U27399 (N_27399,N_25940,N_24211);
xnor U27400 (N_27400,N_24711,N_25085);
or U27401 (N_27401,N_24405,N_24161);
nand U27402 (N_27402,N_24501,N_25095);
nand U27403 (N_27403,N_24512,N_24827);
xnor U27404 (N_27404,N_24934,N_24117);
nor U27405 (N_27405,N_24758,N_24316);
or U27406 (N_27406,N_24035,N_25790);
and U27407 (N_27407,N_25875,N_25520);
or U27408 (N_27408,N_25143,N_25893);
or U27409 (N_27409,N_25483,N_24244);
nand U27410 (N_27410,N_25576,N_25394);
nand U27411 (N_27411,N_24972,N_25512);
and U27412 (N_27412,N_25653,N_24825);
nor U27413 (N_27413,N_24049,N_24741);
and U27414 (N_27414,N_25603,N_24120);
nor U27415 (N_27415,N_25480,N_25651);
or U27416 (N_27416,N_24347,N_24904);
nor U27417 (N_27417,N_25088,N_24197);
nor U27418 (N_27418,N_24012,N_24602);
nor U27419 (N_27419,N_24877,N_24167);
xor U27420 (N_27420,N_24842,N_24107);
xor U27421 (N_27421,N_25462,N_25707);
or U27422 (N_27422,N_24425,N_24085);
xor U27423 (N_27423,N_25103,N_25342);
nor U27424 (N_27424,N_25868,N_24437);
nor U27425 (N_27425,N_24330,N_25435);
or U27426 (N_27426,N_25495,N_24284);
or U27427 (N_27427,N_25871,N_24543);
or U27428 (N_27428,N_25547,N_24594);
and U27429 (N_27429,N_25418,N_24279);
or U27430 (N_27430,N_25137,N_25131);
xor U27431 (N_27431,N_25243,N_24635);
xnor U27432 (N_27432,N_24348,N_24983);
or U27433 (N_27433,N_24517,N_25680);
and U27434 (N_27434,N_24699,N_24036);
xnor U27435 (N_27435,N_24983,N_24143);
xnor U27436 (N_27436,N_24097,N_24717);
xnor U27437 (N_27437,N_25854,N_25774);
nand U27438 (N_27438,N_25101,N_25681);
xor U27439 (N_27439,N_25686,N_24259);
nor U27440 (N_27440,N_25841,N_25374);
nand U27441 (N_27441,N_25108,N_24916);
xnor U27442 (N_27442,N_25698,N_25481);
and U27443 (N_27443,N_24403,N_25185);
nand U27444 (N_27444,N_24005,N_25011);
xor U27445 (N_27445,N_25208,N_24592);
nand U27446 (N_27446,N_24646,N_25445);
nor U27447 (N_27447,N_25400,N_24304);
and U27448 (N_27448,N_24794,N_25657);
xor U27449 (N_27449,N_24938,N_24172);
xor U27450 (N_27450,N_24043,N_25405);
and U27451 (N_27451,N_25431,N_25100);
nor U27452 (N_27452,N_24517,N_24378);
or U27453 (N_27453,N_24856,N_25166);
nor U27454 (N_27454,N_24971,N_25750);
nand U27455 (N_27455,N_25845,N_25469);
nor U27456 (N_27456,N_25048,N_24884);
nor U27457 (N_27457,N_25418,N_24540);
nor U27458 (N_27458,N_25683,N_25299);
or U27459 (N_27459,N_25537,N_25721);
or U27460 (N_27460,N_24428,N_24001);
xor U27461 (N_27461,N_25514,N_25389);
nor U27462 (N_27462,N_24854,N_24122);
and U27463 (N_27463,N_25118,N_25501);
nor U27464 (N_27464,N_25380,N_24357);
or U27465 (N_27465,N_24622,N_24436);
and U27466 (N_27466,N_25641,N_24086);
nand U27467 (N_27467,N_25551,N_25133);
or U27468 (N_27468,N_24584,N_25716);
or U27469 (N_27469,N_24315,N_25178);
nor U27470 (N_27470,N_24725,N_25182);
nand U27471 (N_27471,N_24287,N_24718);
or U27472 (N_27472,N_24230,N_25661);
and U27473 (N_27473,N_25001,N_24181);
nand U27474 (N_27474,N_24878,N_24567);
nor U27475 (N_27475,N_25085,N_24164);
nand U27476 (N_27476,N_24837,N_24301);
or U27477 (N_27477,N_25591,N_25923);
or U27478 (N_27478,N_24784,N_25760);
nand U27479 (N_27479,N_24003,N_25232);
and U27480 (N_27480,N_25747,N_24541);
or U27481 (N_27481,N_24955,N_24288);
xor U27482 (N_27482,N_25943,N_24795);
or U27483 (N_27483,N_25657,N_24504);
nor U27484 (N_27484,N_25042,N_24288);
xnor U27485 (N_27485,N_24092,N_25624);
nor U27486 (N_27486,N_24992,N_24677);
xor U27487 (N_27487,N_25317,N_25539);
nor U27488 (N_27488,N_25506,N_24385);
nor U27489 (N_27489,N_25645,N_24069);
or U27490 (N_27490,N_24171,N_25003);
nand U27491 (N_27491,N_25794,N_25029);
or U27492 (N_27492,N_25377,N_24915);
and U27493 (N_27493,N_24352,N_24129);
nor U27494 (N_27494,N_24846,N_25810);
xor U27495 (N_27495,N_25756,N_25695);
and U27496 (N_27496,N_24666,N_24228);
xor U27497 (N_27497,N_24091,N_25470);
nor U27498 (N_27498,N_24871,N_25302);
and U27499 (N_27499,N_24294,N_24310);
or U27500 (N_27500,N_25024,N_24605);
xnor U27501 (N_27501,N_25399,N_24400);
and U27502 (N_27502,N_24330,N_24927);
and U27503 (N_27503,N_25976,N_25458);
xor U27504 (N_27504,N_25188,N_25127);
or U27505 (N_27505,N_25714,N_25755);
nor U27506 (N_27506,N_24285,N_24702);
or U27507 (N_27507,N_25282,N_24504);
nand U27508 (N_27508,N_24537,N_24073);
and U27509 (N_27509,N_25884,N_24837);
nand U27510 (N_27510,N_25970,N_25986);
xnor U27511 (N_27511,N_25177,N_24975);
nor U27512 (N_27512,N_25793,N_25498);
and U27513 (N_27513,N_25709,N_24148);
nor U27514 (N_27514,N_25192,N_24048);
xor U27515 (N_27515,N_24192,N_25858);
xnor U27516 (N_27516,N_25314,N_24298);
nor U27517 (N_27517,N_25610,N_25969);
nand U27518 (N_27518,N_24006,N_24198);
nor U27519 (N_27519,N_25409,N_25735);
and U27520 (N_27520,N_25566,N_25849);
nand U27521 (N_27521,N_25732,N_24319);
xnor U27522 (N_27522,N_25192,N_24707);
xor U27523 (N_27523,N_24942,N_24026);
or U27524 (N_27524,N_25520,N_25710);
xnor U27525 (N_27525,N_25933,N_25804);
xnor U27526 (N_27526,N_25396,N_24926);
xnor U27527 (N_27527,N_25936,N_25106);
and U27528 (N_27528,N_24451,N_25297);
and U27529 (N_27529,N_25597,N_25833);
and U27530 (N_27530,N_25840,N_24765);
and U27531 (N_27531,N_24305,N_25411);
nor U27532 (N_27532,N_25310,N_25521);
xnor U27533 (N_27533,N_24384,N_25389);
and U27534 (N_27534,N_25586,N_24927);
and U27535 (N_27535,N_25414,N_25826);
nor U27536 (N_27536,N_25670,N_25042);
nor U27537 (N_27537,N_24469,N_25957);
or U27538 (N_27538,N_25253,N_25580);
or U27539 (N_27539,N_25364,N_24706);
xor U27540 (N_27540,N_25817,N_24044);
nor U27541 (N_27541,N_24635,N_24464);
nand U27542 (N_27542,N_25578,N_24215);
nor U27543 (N_27543,N_25034,N_24461);
or U27544 (N_27544,N_24106,N_25714);
nor U27545 (N_27545,N_24688,N_24563);
xnor U27546 (N_27546,N_24438,N_24297);
nand U27547 (N_27547,N_24587,N_24399);
and U27548 (N_27548,N_25353,N_25636);
nand U27549 (N_27549,N_24980,N_25035);
nor U27550 (N_27550,N_24791,N_25025);
nor U27551 (N_27551,N_25175,N_25791);
and U27552 (N_27552,N_25478,N_24302);
and U27553 (N_27553,N_24601,N_24603);
nor U27554 (N_27554,N_25525,N_25887);
nand U27555 (N_27555,N_25031,N_25767);
or U27556 (N_27556,N_24925,N_25088);
or U27557 (N_27557,N_24601,N_24348);
or U27558 (N_27558,N_24872,N_25508);
or U27559 (N_27559,N_24916,N_24487);
xnor U27560 (N_27560,N_24845,N_25898);
nor U27561 (N_27561,N_25013,N_24397);
xnor U27562 (N_27562,N_24060,N_24393);
nor U27563 (N_27563,N_24297,N_24320);
nor U27564 (N_27564,N_25996,N_24296);
nand U27565 (N_27565,N_25387,N_24252);
and U27566 (N_27566,N_25884,N_24403);
nor U27567 (N_27567,N_24805,N_25378);
xnor U27568 (N_27568,N_25772,N_25583);
or U27569 (N_27569,N_25568,N_24040);
nand U27570 (N_27570,N_25498,N_24042);
nor U27571 (N_27571,N_25632,N_24674);
nand U27572 (N_27572,N_25462,N_25131);
and U27573 (N_27573,N_24539,N_24326);
nand U27574 (N_27574,N_25812,N_25608);
xnor U27575 (N_27575,N_24512,N_24131);
nand U27576 (N_27576,N_25606,N_24248);
and U27577 (N_27577,N_24919,N_25390);
nor U27578 (N_27578,N_25693,N_25903);
nand U27579 (N_27579,N_24910,N_25982);
xnor U27580 (N_27580,N_25956,N_25155);
xor U27581 (N_27581,N_24679,N_24029);
nand U27582 (N_27582,N_24128,N_25042);
and U27583 (N_27583,N_25195,N_25261);
xnor U27584 (N_27584,N_25543,N_24178);
nor U27585 (N_27585,N_24446,N_24042);
nand U27586 (N_27586,N_24012,N_25844);
and U27587 (N_27587,N_25793,N_25304);
and U27588 (N_27588,N_24091,N_24365);
or U27589 (N_27589,N_25375,N_24893);
nor U27590 (N_27590,N_24906,N_25552);
and U27591 (N_27591,N_25008,N_24867);
xnor U27592 (N_27592,N_24790,N_24549);
and U27593 (N_27593,N_25426,N_25894);
xor U27594 (N_27594,N_24023,N_24916);
nor U27595 (N_27595,N_25516,N_25911);
nor U27596 (N_27596,N_25208,N_24079);
nor U27597 (N_27597,N_24554,N_24869);
or U27598 (N_27598,N_24612,N_24983);
and U27599 (N_27599,N_25013,N_24947);
xor U27600 (N_27600,N_24925,N_24763);
xnor U27601 (N_27601,N_25929,N_25680);
xnor U27602 (N_27602,N_24077,N_25716);
nand U27603 (N_27603,N_25769,N_25255);
nand U27604 (N_27604,N_25801,N_25234);
xor U27605 (N_27605,N_25196,N_24128);
nor U27606 (N_27606,N_25403,N_24702);
xnor U27607 (N_27607,N_24215,N_25849);
nand U27608 (N_27608,N_25498,N_24001);
or U27609 (N_27609,N_25799,N_24238);
nor U27610 (N_27610,N_24810,N_25582);
nand U27611 (N_27611,N_24449,N_24049);
xnor U27612 (N_27612,N_24247,N_25619);
and U27613 (N_27613,N_24797,N_24273);
and U27614 (N_27614,N_24964,N_25103);
and U27615 (N_27615,N_25856,N_24399);
and U27616 (N_27616,N_24740,N_24746);
xor U27617 (N_27617,N_24146,N_25666);
or U27618 (N_27618,N_24143,N_25278);
nand U27619 (N_27619,N_25192,N_24596);
xnor U27620 (N_27620,N_24245,N_25235);
and U27621 (N_27621,N_24634,N_25621);
nor U27622 (N_27622,N_25816,N_24891);
and U27623 (N_27623,N_24210,N_24994);
and U27624 (N_27624,N_25009,N_25568);
xor U27625 (N_27625,N_24052,N_25716);
xnor U27626 (N_27626,N_24676,N_24065);
nand U27627 (N_27627,N_24451,N_24438);
nand U27628 (N_27628,N_24581,N_25740);
nor U27629 (N_27629,N_25689,N_25484);
or U27630 (N_27630,N_25814,N_24186);
xnor U27631 (N_27631,N_24484,N_24211);
nor U27632 (N_27632,N_24206,N_24830);
xor U27633 (N_27633,N_24975,N_25578);
nor U27634 (N_27634,N_24805,N_25102);
nor U27635 (N_27635,N_24542,N_25610);
nor U27636 (N_27636,N_25202,N_25702);
nand U27637 (N_27637,N_24054,N_24987);
nor U27638 (N_27638,N_25355,N_24276);
nor U27639 (N_27639,N_24866,N_24024);
and U27640 (N_27640,N_24191,N_24359);
and U27641 (N_27641,N_25580,N_24428);
or U27642 (N_27642,N_25685,N_24021);
and U27643 (N_27643,N_25533,N_24478);
and U27644 (N_27644,N_25060,N_25408);
and U27645 (N_27645,N_24716,N_25955);
and U27646 (N_27646,N_25269,N_25079);
nor U27647 (N_27647,N_24168,N_24118);
nand U27648 (N_27648,N_24005,N_24360);
or U27649 (N_27649,N_24089,N_25681);
or U27650 (N_27650,N_24921,N_25435);
and U27651 (N_27651,N_25300,N_25867);
or U27652 (N_27652,N_24742,N_24987);
xnor U27653 (N_27653,N_25433,N_25618);
nand U27654 (N_27654,N_25671,N_25482);
nand U27655 (N_27655,N_24097,N_24825);
or U27656 (N_27656,N_25169,N_25443);
nor U27657 (N_27657,N_24093,N_25641);
or U27658 (N_27658,N_25706,N_25223);
nand U27659 (N_27659,N_24230,N_24052);
nor U27660 (N_27660,N_25873,N_24798);
and U27661 (N_27661,N_24079,N_24235);
xnor U27662 (N_27662,N_24006,N_25857);
and U27663 (N_27663,N_25189,N_24415);
nor U27664 (N_27664,N_24864,N_25479);
nor U27665 (N_27665,N_25325,N_25814);
or U27666 (N_27666,N_25054,N_24206);
nand U27667 (N_27667,N_24722,N_24650);
xnor U27668 (N_27668,N_24834,N_24195);
nand U27669 (N_27669,N_24934,N_25431);
or U27670 (N_27670,N_25202,N_24726);
and U27671 (N_27671,N_24308,N_25042);
xnor U27672 (N_27672,N_24473,N_24786);
or U27673 (N_27673,N_25995,N_25131);
or U27674 (N_27674,N_25237,N_24479);
nor U27675 (N_27675,N_25418,N_24638);
nor U27676 (N_27676,N_24243,N_24482);
xor U27677 (N_27677,N_25874,N_24963);
xor U27678 (N_27678,N_24914,N_25037);
nand U27679 (N_27679,N_24006,N_25530);
nand U27680 (N_27680,N_25917,N_24767);
nor U27681 (N_27681,N_24953,N_25855);
and U27682 (N_27682,N_24427,N_25208);
or U27683 (N_27683,N_24238,N_25095);
or U27684 (N_27684,N_24744,N_25229);
nor U27685 (N_27685,N_25847,N_25266);
nand U27686 (N_27686,N_24003,N_25392);
and U27687 (N_27687,N_24219,N_24452);
nor U27688 (N_27688,N_25934,N_25151);
and U27689 (N_27689,N_25026,N_25741);
nand U27690 (N_27690,N_24703,N_24121);
xor U27691 (N_27691,N_24958,N_25500);
xnor U27692 (N_27692,N_25044,N_24959);
or U27693 (N_27693,N_24999,N_24393);
or U27694 (N_27694,N_24424,N_25654);
nor U27695 (N_27695,N_24330,N_25346);
and U27696 (N_27696,N_24089,N_24295);
and U27697 (N_27697,N_24513,N_24035);
nand U27698 (N_27698,N_25684,N_25533);
and U27699 (N_27699,N_24571,N_24114);
nor U27700 (N_27700,N_24714,N_24935);
nor U27701 (N_27701,N_25370,N_25170);
nand U27702 (N_27702,N_25494,N_25011);
nor U27703 (N_27703,N_24841,N_25520);
or U27704 (N_27704,N_25431,N_24615);
nand U27705 (N_27705,N_24640,N_24303);
or U27706 (N_27706,N_24512,N_25030);
and U27707 (N_27707,N_24543,N_25628);
nand U27708 (N_27708,N_24488,N_25261);
and U27709 (N_27709,N_24924,N_25476);
and U27710 (N_27710,N_24593,N_25941);
and U27711 (N_27711,N_24974,N_25460);
xor U27712 (N_27712,N_25337,N_25392);
nand U27713 (N_27713,N_25365,N_25156);
nand U27714 (N_27714,N_25731,N_24015);
nand U27715 (N_27715,N_25490,N_25963);
xnor U27716 (N_27716,N_25251,N_24966);
or U27717 (N_27717,N_25518,N_25256);
nor U27718 (N_27718,N_25942,N_25223);
xor U27719 (N_27719,N_25587,N_25975);
nand U27720 (N_27720,N_24998,N_25115);
nor U27721 (N_27721,N_25421,N_25935);
xnor U27722 (N_27722,N_24184,N_24555);
or U27723 (N_27723,N_25411,N_24986);
nand U27724 (N_27724,N_25908,N_25653);
nor U27725 (N_27725,N_24589,N_25892);
and U27726 (N_27726,N_24197,N_24622);
nand U27727 (N_27727,N_25283,N_24912);
xnor U27728 (N_27728,N_25674,N_24325);
and U27729 (N_27729,N_24637,N_25989);
or U27730 (N_27730,N_25414,N_25728);
xnor U27731 (N_27731,N_24949,N_24385);
or U27732 (N_27732,N_25859,N_24917);
and U27733 (N_27733,N_24558,N_24192);
nor U27734 (N_27734,N_24936,N_25509);
nor U27735 (N_27735,N_25545,N_25267);
or U27736 (N_27736,N_25554,N_25664);
nand U27737 (N_27737,N_25210,N_25907);
xor U27738 (N_27738,N_24357,N_24200);
or U27739 (N_27739,N_25094,N_24583);
nor U27740 (N_27740,N_25675,N_24276);
or U27741 (N_27741,N_25917,N_24332);
nor U27742 (N_27742,N_25395,N_25836);
and U27743 (N_27743,N_25819,N_24753);
xnor U27744 (N_27744,N_25542,N_25674);
xnor U27745 (N_27745,N_25754,N_25346);
or U27746 (N_27746,N_25428,N_25456);
and U27747 (N_27747,N_25122,N_25343);
xnor U27748 (N_27748,N_25602,N_24840);
and U27749 (N_27749,N_25579,N_25006);
xnor U27750 (N_27750,N_24455,N_24661);
nand U27751 (N_27751,N_24289,N_25996);
xnor U27752 (N_27752,N_25366,N_24067);
xor U27753 (N_27753,N_24848,N_25995);
nor U27754 (N_27754,N_24452,N_25980);
and U27755 (N_27755,N_24994,N_24045);
and U27756 (N_27756,N_25864,N_25496);
xnor U27757 (N_27757,N_25045,N_25385);
nor U27758 (N_27758,N_24307,N_24933);
nand U27759 (N_27759,N_24681,N_24451);
nor U27760 (N_27760,N_24267,N_24849);
and U27761 (N_27761,N_24041,N_25852);
nor U27762 (N_27762,N_24805,N_25663);
xor U27763 (N_27763,N_24640,N_25947);
and U27764 (N_27764,N_25625,N_24654);
nand U27765 (N_27765,N_25823,N_24344);
nor U27766 (N_27766,N_24544,N_25758);
xor U27767 (N_27767,N_24378,N_24552);
xor U27768 (N_27768,N_25437,N_25258);
nand U27769 (N_27769,N_25408,N_25201);
nand U27770 (N_27770,N_24940,N_25507);
or U27771 (N_27771,N_25049,N_25565);
nor U27772 (N_27772,N_25021,N_25713);
nor U27773 (N_27773,N_25142,N_24438);
nand U27774 (N_27774,N_24796,N_25067);
xor U27775 (N_27775,N_24588,N_25759);
nor U27776 (N_27776,N_25539,N_24694);
and U27777 (N_27777,N_24672,N_25027);
and U27778 (N_27778,N_24644,N_24333);
and U27779 (N_27779,N_25128,N_25129);
and U27780 (N_27780,N_25307,N_25364);
xor U27781 (N_27781,N_25721,N_25963);
nor U27782 (N_27782,N_25227,N_25266);
or U27783 (N_27783,N_24263,N_24331);
and U27784 (N_27784,N_24928,N_24206);
and U27785 (N_27785,N_24557,N_24696);
nand U27786 (N_27786,N_25860,N_25745);
nand U27787 (N_27787,N_24257,N_24438);
and U27788 (N_27788,N_24864,N_25132);
and U27789 (N_27789,N_24399,N_24381);
nor U27790 (N_27790,N_25476,N_25003);
nor U27791 (N_27791,N_24980,N_25871);
and U27792 (N_27792,N_25323,N_25585);
xnor U27793 (N_27793,N_25456,N_24047);
and U27794 (N_27794,N_25610,N_24132);
xnor U27795 (N_27795,N_25204,N_24389);
xor U27796 (N_27796,N_25622,N_25400);
xor U27797 (N_27797,N_24911,N_25880);
and U27798 (N_27798,N_25123,N_24584);
and U27799 (N_27799,N_25431,N_24704);
xnor U27800 (N_27800,N_25057,N_24558);
nand U27801 (N_27801,N_25289,N_24789);
nand U27802 (N_27802,N_24686,N_24708);
and U27803 (N_27803,N_24352,N_25593);
nand U27804 (N_27804,N_25718,N_25873);
xor U27805 (N_27805,N_24574,N_25035);
and U27806 (N_27806,N_24363,N_25821);
and U27807 (N_27807,N_24931,N_24654);
nand U27808 (N_27808,N_24383,N_24347);
nand U27809 (N_27809,N_24158,N_25579);
or U27810 (N_27810,N_25352,N_25198);
xnor U27811 (N_27811,N_24457,N_25060);
xor U27812 (N_27812,N_24341,N_25551);
xor U27813 (N_27813,N_25593,N_25363);
and U27814 (N_27814,N_24954,N_24830);
nor U27815 (N_27815,N_25192,N_25511);
nor U27816 (N_27816,N_24183,N_24408);
xor U27817 (N_27817,N_25287,N_24411);
or U27818 (N_27818,N_24470,N_24773);
or U27819 (N_27819,N_24873,N_24675);
and U27820 (N_27820,N_24080,N_25020);
nor U27821 (N_27821,N_24109,N_24324);
and U27822 (N_27822,N_24405,N_25532);
xnor U27823 (N_27823,N_24554,N_24638);
nand U27824 (N_27824,N_25536,N_24374);
xor U27825 (N_27825,N_24420,N_24184);
nor U27826 (N_27826,N_24168,N_24725);
and U27827 (N_27827,N_24331,N_25746);
xor U27828 (N_27828,N_25629,N_25825);
xnor U27829 (N_27829,N_25050,N_25319);
nand U27830 (N_27830,N_24627,N_24246);
xnor U27831 (N_27831,N_25987,N_25002);
nor U27832 (N_27832,N_24366,N_24584);
xor U27833 (N_27833,N_24146,N_24663);
nor U27834 (N_27834,N_24398,N_25815);
and U27835 (N_27835,N_24545,N_25296);
and U27836 (N_27836,N_24981,N_24319);
or U27837 (N_27837,N_25460,N_24964);
or U27838 (N_27838,N_24256,N_25896);
nor U27839 (N_27839,N_24131,N_24025);
or U27840 (N_27840,N_25188,N_24026);
and U27841 (N_27841,N_24809,N_24637);
or U27842 (N_27842,N_24981,N_24450);
and U27843 (N_27843,N_24990,N_25914);
xnor U27844 (N_27844,N_25406,N_24735);
nor U27845 (N_27845,N_25758,N_24994);
or U27846 (N_27846,N_25582,N_24567);
nor U27847 (N_27847,N_24297,N_24241);
and U27848 (N_27848,N_25465,N_25116);
nand U27849 (N_27849,N_24079,N_25351);
or U27850 (N_27850,N_25815,N_25150);
nor U27851 (N_27851,N_24277,N_25230);
xnor U27852 (N_27852,N_25131,N_24697);
or U27853 (N_27853,N_25974,N_25395);
xnor U27854 (N_27854,N_24056,N_25407);
xor U27855 (N_27855,N_24805,N_25599);
nand U27856 (N_27856,N_25232,N_24877);
or U27857 (N_27857,N_24432,N_25786);
and U27858 (N_27858,N_24479,N_24743);
xor U27859 (N_27859,N_24561,N_25743);
or U27860 (N_27860,N_25673,N_24809);
xnor U27861 (N_27861,N_24035,N_24709);
xnor U27862 (N_27862,N_25937,N_25896);
xor U27863 (N_27863,N_24853,N_24017);
xor U27864 (N_27864,N_25415,N_25558);
nor U27865 (N_27865,N_25569,N_24081);
and U27866 (N_27866,N_25411,N_24564);
xnor U27867 (N_27867,N_24455,N_24448);
and U27868 (N_27868,N_25198,N_24565);
or U27869 (N_27869,N_25460,N_24382);
nand U27870 (N_27870,N_24033,N_24958);
or U27871 (N_27871,N_25073,N_25678);
nand U27872 (N_27872,N_25316,N_25256);
and U27873 (N_27873,N_24660,N_24215);
or U27874 (N_27874,N_25454,N_24053);
nor U27875 (N_27875,N_25790,N_24101);
nand U27876 (N_27876,N_24766,N_24475);
or U27877 (N_27877,N_24229,N_25257);
nor U27878 (N_27878,N_25236,N_25884);
nand U27879 (N_27879,N_25263,N_24673);
nand U27880 (N_27880,N_25427,N_24322);
nor U27881 (N_27881,N_25079,N_25595);
nor U27882 (N_27882,N_24183,N_24558);
and U27883 (N_27883,N_24515,N_25762);
nor U27884 (N_27884,N_24163,N_25132);
xor U27885 (N_27885,N_25968,N_24560);
and U27886 (N_27886,N_25454,N_25136);
xor U27887 (N_27887,N_24413,N_25602);
and U27888 (N_27888,N_25187,N_25423);
or U27889 (N_27889,N_25243,N_24394);
nand U27890 (N_27890,N_24032,N_24876);
nor U27891 (N_27891,N_25530,N_24107);
nor U27892 (N_27892,N_24368,N_24944);
nor U27893 (N_27893,N_25193,N_25612);
xnor U27894 (N_27894,N_25849,N_24550);
and U27895 (N_27895,N_24099,N_25552);
nor U27896 (N_27896,N_25210,N_24484);
xnor U27897 (N_27897,N_24347,N_25536);
or U27898 (N_27898,N_25426,N_25206);
nand U27899 (N_27899,N_24182,N_24869);
nand U27900 (N_27900,N_24009,N_25939);
or U27901 (N_27901,N_25631,N_25011);
xor U27902 (N_27902,N_25565,N_24721);
xnor U27903 (N_27903,N_25611,N_25506);
nor U27904 (N_27904,N_24434,N_24058);
or U27905 (N_27905,N_24385,N_24416);
nand U27906 (N_27906,N_24486,N_24675);
and U27907 (N_27907,N_25212,N_24534);
and U27908 (N_27908,N_25173,N_24027);
and U27909 (N_27909,N_25283,N_24699);
and U27910 (N_27910,N_25610,N_24448);
xnor U27911 (N_27911,N_25885,N_24554);
and U27912 (N_27912,N_25560,N_24597);
xor U27913 (N_27913,N_25640,N_25897);
or U27914 (N_27914,N_24400,N_24026);
or U27915 (N_27915,N_24251,N_25499);
and U27916 (N_27916,N_25359,N_25882);
nor U27917 (N_27917,N_25883,N_24911);
nor U27918 (N_27918,N_25026,N_25620);
and U27919 (N_27919,N_24806,N_24981);
or U27920 (N_27920,N_24438,N_25224);
nor U27921 (N_27921,N_24383,N_25021);
and U27922 (N_27922,N_24485,N_24845);
xor U27923 (N_27923,N_24581,N_24275);
nand U27924 (N_27924,N_25952,N_24436);
nor U27925 (N_27925,N_25676,N_24819);
or U27926 (N_27926,N_24626,N_24622);
and U27927 (N_27927,N_24277,N_25246);
nor U27928 (N_27928,N_24844,N_24976);
or U27929 (N_27929,N_24551,N_25514);
xor U27930 (N_27930,N_25065,N_25323);
xor U27931 (N_27931,N_25492,N_25830);
or U27932 (N_27932,N_24622,N_25759);
and U27933 (N_27933,N_25806,N_24213);
nand U27934 (N_27934,N_25051,N_25858);
nor U27935 (N_27935,N_25655,N_25338);
xnor U27936 (N_27936,N_25072,N_25745);
nor U27937 (N_27937,N_24289,N_25244);
xnor U27938 (N_27938,N_24079,N_25492);
nor U27939 (N_27939,N_24537,N_25610);
and U27940 (N_27940,N_24266,N_24468);
xnor U27941 (N_27941,N_24516,N_24300);
nand U27942 (N_27942,N_24026,N_24298);
nand U27943 (N_27943,N_25574,N_25812);
nor U27944 (N_27944,N_25018,N_25289);
nor U27945 (N_27945,N_25179,N_25017);
nor U27946 (N_27946,N_25302,N_25380);
nand U27947 (N_27947,N_24841,N_24444);
xnor U27948 (N_27948,N_24923,N_24096);
and U27949 (N_27949,N_25366,N_25089);
nor U27950 (N_27950,N_25990,N_24644);
xnor U27951 (N_27951,N_24411,N_24470);
nand U27952 (N_27952,N_25614,N_24414);
nor U27953 (N_27953,N_25750,N_25077);
nand U27954 (N_27954,N_25674,N_25990);
nand U27955 (N_27955,N_24726,N_24046);
xnor U27956 (N_27956,N_24863,N_25571);
and U27957 (N_27957,N_25938,N_25758);
nor U27958 (N_27958,N_24213,N_24251);
nor U27959 (N_27959,N_24928,N_24373);
or U27960 (N_27960,N_25976,N_24061);
and U27961 (N_27961,N_24928,N_25854);
and U27962 (N_27962,N_24804,N_24135);
and U27963 (N_27963,N_24951,N_25231);
or U27964 (N_27964,N_24659,N_25603);
nor U27965 (N_27965,N_25606,N_24564);
xnor U27966 (N_27966,N_25732,N_25149);
xor U27967 (N_27967,N_24832,N_25601);
nand U27968 (N_27968,N_24786,N_24619);
nand U27969 (N_27969,N_24931,N_24543);
nand U27970 (N_27970,N_25202,N_25313);
nor U27971 (N_27971,N_24228,N_25726);
xor U27972 (N_27972,N_25565,N_25113);
or U27973 (N_27973,N_24780,N_25115);
or U27974 (N_27974,N_24542,N_24186);
or U27975 (N_27975,N_25843,N_24143);
nor U27976 (N_27976,N_25404,N_25009);
nand U27977 (N_27977,N_24282,N_25762);
xnor U27978 (N_27978,N_24095,N_25985);
or U27979 (N_27979,N_25197,N_25909);
nor U27980 (N_27980,N_24492,N_25046);
nand U27981 (N_27981,N_25253,N_24605);
xnor U27982 (N_27982,N_24176,N_24760);
xnor U27983 (N_27983,N_24707,N_25882);
or U27984 (N_27984,N_25984,N_25306);
and U27985 (N_27985,N_24045,N_24791);
nand U27986 (N_27986,N_24929,N_25640);
and U27987 (N_27987,N_24383,N_24980);
nand U27988 (N_27988,N_24876,N_25248);
nor U27989 (N_27989,N_24133,N_25188);
nor U27990 (N_27990,N_25978,N_25407);
xor U27991 (N_27991,N_24580,N_24548);
or U27992 (N_27992,N_24960,N_25508);
nand U27993 (N_27993,N_25949,N_25763);
or U27994 (N_27994,N_25501,N_24072);
and U27995 (N_27995,N_25885,N_24184);
xnor U27996 (N_27996,N_24990,N_24263);
and U27997 (N_27997,N_24242,N_24414);
nand U27998 (N_27998,N_25663,N_24260);
nand U27999 (N_27999,N_25755,N_24977);
nor U28000 (N_28000,N_26881,N_26073);
and U28001 (N_28001,N_26564,N_26316);
nand U28002 (N_28002,N_26311,N_26972);
or U28003 (N_28003,N_27488,N_27794);
xnor U28004 (N_28004,N_26514,N_26076);
nor U28005 (N_28005,N_27973,N_26150);
and U28006 (N_28006,N_27838,N_27668);
nand U28007 (N_28007,N_26672,N_27114);
xor U28008 (N_28008,N_27185,N_27879);
or U28009 (N_28009,N_26622,N_27005);
nor U28010 (N_28010,N_27239,N_27715);
and U28011 (N_28011,N_26499,N_26847);
nor U28012 (N_28012,N_26159,N_27015);
and U28013 (N_28013,N_26268,N_27186);
nand U28014 (N_28014,N_26107,N_26758);
nor U28015 (N_28015,N_27483,N_26255);
nand U28016 (N_28016,N_27354,N_27828);
or U28017 (N_28017,N_26208,N_27583);
or U28018 (N_28018,N_27642,N_26968);
or U28019 (N_28019,N_27027,N_26318);
and U28020 (N_28020,N_26433,N_26781);
xor U28021 (N_28021,N_26606,N_27290);
and U28022 (N_28022,N_27166,N_26686);
or U28023 (N_28023,N_26590,N_26331);
or U28024 (N_28024,N_26414,N_27825);
xor U28025 (N_28025,N_27970,N_26504);
nand U28026 (N_28026,N_27150,N_27842);
xnor U28027 (N_28027,N_26443,N_26647);
nor U28028 (N_28028,N_26532,N_27826);
and U28029 (N_28029,N_26179,N_27883);
or U28030 (N_28030,N_26120,N_26144);
xnor U28031 (N_28031,N_27292,N_26645);
and U28032 (N_28032,N_26767,N_27938);
and U28033 (N_28033,N_27587,N_26244);
or U28034 (N_28034,N_26229,N_27368);
xor U28035 (N_28035,N_27361,N_27038);
or U28036 (N_28036,N_26842,N_27796);
xor U28037 (N_28037,N_27533,N_27846);
xnor U28038 (N_28038,N_26792,N_26997);
or U28039 (N_28039,N_27785,N_27907);
nand U28040 (N_28040,N_27744,N_27873);
nand U28041 (N_28041,N_26247,N_26552);
nor U28042 (N_28042,N_27051,N_26367);
nor U28043 (N_28043,N_27500,N_26475);
xor U28044 (N_28044,N_26115,N_27236);
or U28045 (N_28045,N_26542,N_26990);
and U28046 (N_28046,N_27460,N_26026);
xor U28047 (N_28047,N_26184,N_26954);
nor U28048 (N_28048,N_26512,N_26498);
nand U28049 (N_28049,N_27517,N_26085);
nor U28050 (N_28050,N_26832,N_26691);
nand U28051 (N_28051,N_26624,N_26041);
and U28052 (N_28052,N_26882,N_26711);
nand U28053 (N_28053,N_26416,N_27248);
and U28054 (N_28054,N_27058,N_26299);
or U28055 (N_28055,N_26520,N_27891);
xor U28056 (N_28056,N_26503,N_26977);
nor U28057 (N_28057,N_26217,N_26518);
nor U28058 (N_28058,N_26509,N_26690);
xor U28059 (N_28059,N_27733,N_26826);
nand U28060 (N_28060,N_27641,N_26209);
and U28061 (N_28061,N_27366,N_26889);
nor U28062 (N_28062,N_26338,N_26019);
nor U28063 (N_28063,N_27095,N_27285);
nor U28064 (N_28064,N_27017,N_26205);
nor U28065 (N_28065,N_26821,N_26613);
nor U28066 (N_28066,N_27676,N_26707);
xor U28067 (N_28067,N_27060,N_27103);
or U28068 (N_28068,N_26770,N_26204);
or U28069 (N_28069,N_26133,N_26040);
nor U28070 (N_28070,N_26480,N_26407);
or U28071 (N_28071,N_26719,N_27718);
nor U28072 (N_28072,N_27824,N_26359);
xnor U28073 (N_28073,N_26105,N_26478);
xor U28074 (N_28074,N_26627,N_26259);
or U28075 (N_28075,N_27886,N_27313);
or U28076 (N_28076,N_26103,N_27735);
nand U28077 (N_28077,N_26699,N_26701);
and U28078 (N_28078,N_26904,N_27013);
nand U28079 (N_28079,N_26315,N_27072);
nor U28080 (N_28080,N_26530,N_26570);
nor U28081 (N_28081,N_27801,N_26232);
and U28082 (N_28082,N_27155,N_26868);
or U28083 (N_28083,N_27905,N_27463);
and U28084 (N_28084,N_27710,N_26174);
and U28085 (N_28085,N_26397,N_26959);
nand U28086 (N_28086,N_26546,N_26740);
nand U28087 (N_28087,N_27756,N_27924);
xnor U28088 (N_28088,N_27009,N_26181);
xnor U28089 (N_28089,N_27277,N_27346);
nor U28090 (N_28090,N_26079,N_26093);
or U28091 (N_28091,N_27048,N_26974);
and U28092 (N_28092,N_26886,N_26097);
nand U28093 (N_28093,N_27403,N_26537);
nor U28094 (N_28094,N_27479,N_27031);
nor U28095 (N_28095,N_26545,N_27142);
and U28096 (N_28096,N_27570,N_27991);
nand U28097 (N_28097,N_27267,N_26577);
and U28098 (N_28098,N_27566,N_26907);
or U28099 (N_28099,N_27437,N_27790);
nand U28100 (N_28100,N_26598,N_26892);
nand U28101 (N_28101,N_27082,N_27025);
or U28102 (N_28102,N_27326,N_26063);
and U28103 (N_28103,N_26698,N_27163);
nand U28104 (N_28104,N_27011,N_26372);
nand U28105 (N_28105,N_27680,N_27887);
or U28106 (N_28106,N_26484,N_27432);
nand U28107 (N_28107,N_27063,N_26724);
or U28108 (N_28108,N_26243,N_27309);
xnor U28109 (N_28109,N_26845,N_26938);
xnor U28110 (N_28110,N_27995,N_26389);
or U28111 (N_28111,N_26313,N_27521);
nand U28112 (N_28112,N_27493,N_27107);
or U28113 (N_28113,N_27913,N_26031);
nor U28114 (N_28114,N_27141,N_26055);
xnor U28115 (N_28115,N_27921,N_26511);
xor U28116 (N_28116,N_26114,N_27211);
or U28117 (N_28117,N_27644,N_26365);
nand U28118 (N_28118,N_26576,N_27553);
or U28119 (N_28119,N_27998,N_26398);
nand U28120 (N_28120,N_27990,N_27010);
nand U28121 (N_28121,N_26800,N_26728);
and U28122 (N_28122,N_26227,N_27923);
and U28123 (N_28123,N_26075,N_27898);
nor U28124 (N_28124,N_27499,N_27764);
xnor U28125 (N_28125,N_26487,N_26177);
xor U28126 (N_28126,N_26677,N_27979);
or U28127 (N_28127,N_26777,N_27817);
or U28128 (N_28128,N_27743,N_26981);
xor U28129 (N_28129,N_27333,N_26950);
or U28130 (N_28130,N_26601,N_26898);
nand U28131 (N_28131,N_26084,N_26952);
xnor U28132 (N_28132,N_27286,N_26797);
and U28133 (N_28133,N_27509,N_27943);
or U28134 (N_28134,N_27885,N_27757);
nand U28135 (N_28135,N_26057,N_26617);
or U28136 (N_28136,N_26269,N_26322);
and U28137 (N_28137,N_27515,N_26531);
xnor U28138 (N_28138,N_27508,N_26448);
xnor U28139 (N_28139,N_27673,N_27040);
or U28140 (N_28140,N_26835,N_27853);
nor U28141 (N_28141,N_26658,N_27420);
and U28142 (N_28142,N_27199,N_27647);
or U28143 (N_28143,N_27843,N_26616);
or U28144 (N_28144,N_26429,N_27201);
nand U28145 (N_28145,N_26388,N_27593);
nor U28146 (N_28146,N_27954,N_27863);
and U28147 (N_28147,N_26580,N_27165);
nor U28148 (N_28148,N_27541,N_27330);
or U28149 (N_28149,N_26653,N_27547);
nand U28150 (N_28150,N_27297,N_27156);
and U28151 (N_28151,N_27503,N_26368);
and U28152 (N_28152,N_27404,N_26853);
nor U28153 (N_28153,N_26408,N_26104);
or U28154 (N_28154,N_27773,N_26615);
or U28155 (N_28155,N_27836,N_27104);
or U28156 (N_28156,N_26796,N_26806);
and U28157 (N_28157,N_26683,N_27430);
and U28158 (N_28158,N_26086,N_26088);
nand U28159 (N_28159,N_27901,N_26725);
and U28160 (N_28160,N_27847,N_26347);
xor U28161 (N_28161,N_26863,N_27724);
or U28162 (N_28162,N_26936,N_26377);
or U28163 (N_28163,N_26510,N_27305);
or U28164 (N_28164,N_27426,N_27270);
nor U28165 (N_28165,N_27349,N_26267);
nand U28166 (N_28166,N_27487,N_27950);
nand U28167 (N_28167,N_27257,N_27249);
and U28168 (N_28168,N_26988,N_27168);
nand U28169 (N_28169,N_26743,N_27964);
nand U28170 (N_28170,N_26696,N_27220);
and U28171 (N_28171,N_27219,N_26052);
and U28172 (N_28172,N_27262,N_27985);
xor U28173 (N_28173,N_26010,N_26854);
and U28174 (N_28174,N_26874,N_26687);
xnor U28175 (N_28175,N_27164,N_26729);
or U28176 (N_28176,N_27844,N_27288);
nor U28177 (N_28177,N_27656,N_26506);
and U28178 (N_28178,N_27465,N_26718);
or U28179 (N_28179,N_27461,N_26921);
xor U28180 (N_28180,N_26319,N_27029);
and U28181 (N_28181,N_27253,N_26231);
xor U28182 (N_28182,N_27279,N_26391);
and U28183 (N_28183,N_26638,N_27545);
nor U28184 (N_28184,N_27133,N_27878);
nand U28185 (N_28185,N_26918,N_26782);
nand U28186 (N_28186,N_27154,N_27496);
nand U28187 (N_28187,N_26681,N_27121);
nand U28188 (N_28188,N_26922,N_27428);
nand U28189 (N_28189,N_27377,N_26859);
and U28190 (N_28190,N_27822,N_27084);
xor U28191 (N_28191,N_27578,N_27525);
and U28192 (N_28192,N_27654,N_26636);
nor U28193 (N_28193,N_27352,N_26926);
nand U28194 (N_28194,N_27289,N_27085);
or U28195 (N_28195,N_26801,N_26785);
or U28196 (N_28196,N_27633,N_27685);
or U28197 (N_28197,N_26225,N_27215);
nand U28198 (N_28198,N_27221,N_27207);
nor U28199 (N_28199,N_27433,N_26287);
nor U28200 (N_28200,N_27388,N_26422);
and U28201 (N_28201,N_26342,N_27942);
and U28202 (N_28202,N_27120,N_26310);
or U28203 (N_28203,N_27391,N_27706);
nor U28204 (N_28204,N_26713,N_27064);
nor U28205 (N_28205,N_27537,N_27869);
and U28206 (N_28206,N_26945,N_27386);
nand U28207 (N_28207,N_27939,N_26817);
or U28208 (N_28208,N_26934,N_26118);
or U28209 (N_28209,N_26519,N_26112);
xnor U28210 (N_28210,N_27233,N_27606);
nor U28211 (N_28211,N_27161,N_26575);
xor U28212 (N_28212,N_27002,N_26643);
nand U28213 (N_28213,N_27535,N_26543);
nand U28214 (N_28214,N_26553,N_26682);
or U28215 (N_28215,N_26123,N_27783);
nor U28216 (N_28216,N_27694,N_26183);
or U28217 (N_28217,N_27759,N_27745);
and U28218 (N_28218,N_26251,N_26861);
nand U28219 (N_28219,N_26738,N_27044);
and U28220 (N_28220,N_26415,N_27983);
and U28221 (N_28221,N_27781,N_27395);
or U28222 (N_28222,N_26461,N_27291);
nand U28223 (N_28223,N_27284,N_26234);
nor U28224 (N_28224,N_26048,N_27926);
xor U28225 (N_28225,N_27335,N_27365);
xnor U28226 (N_28226,N_26198,N_27434);
and U28227 (N_28227,N_26369,N_27162);
and U28228 (N_28228,N_27135,N_26130);
nand U28229 (N_28229,N_27014,N_26466);
or U28230 (N_28230,N_27083,N_27971);
and U28231 (N_28231,N_26813,N_27977);
and U28232 (N_28232,N_27527,N_26089);
and U28233 (N_28233,N_27118,N_26906);
nand U28234 (N_28234,N_27740,N_27963);
or U28235 (N_28235,N_26896,N_27266);
nor U28236 (N_28236,N_27568,N_26744);
xnor U28237 (N_28237,N_27409,N_27050);
nand U28238 (N_28238,N_26051,N_27965);
or U28239 (N_28239,N_26285,N_27835);
xnor U28240 (N_28240,N_27144,N_26281);
nand U28241 (N_28241,N_27797,N_27076);
xnor U28242 (N_28242,N_27124,N_27188);
nand U28243 (N_28243,N_27555,N_26286);
xnor U28244 (N_28244,N_26432,N_26557);
and U28245 (N_28245,N_27597,N_26927);
or U28246 (N_28246,N_26166,N_27625);
xnor U28247 (N_28247,N_27287,N_27930);
nor U28248 (N_28248,N_26064,N_27876);
and U28249 (N_28249,N_27947,N_26463);
and U28250 (N_28250,N_26467,N_27176);
xor U28251 (N_28251,N_26942,N_26941);
nor U28252 (N_28252,N_26276,N_26404);
nor U28253 (N_28253,N_26016,N_26292);
and U28254 (N_28254,N_26931,N_26883);
nor U28255 (N_28255,N_26341,N_27818);
xnor U28256 (N_28256,N_26659,N_26091);
and U28257 (N_28257,N_27619,N_27484);
xor U28258 (N_28258,N_27256,N_27974);
or U28259 (N_28259,N_27269,N_27519);
or U28260 (N_28260,N_26413,N_27959);
nor U28261 (N_28261,N_26203,N_26715);
and U28262 (N_28262,N_26434,N_26015);
or U28263 (N_28263,N_27451,N_27353);
or U28264 (N_28264,N_26387,N_26910);
and U28265 (N_28265,N_27381,N_26056);
nor U28266 (N_28266,N_26399,N_27489);
xor U28267 (N_28267,N_27731,N_26454);
and U28268 (N_28268,N_27806,N_26884);
xnor U28269 (N_28269,N_27315,N_26556);
or U28270 (N_28270,N_26032,N_27053);
nand U28271 (N_28271,N_27208,N_26538);
or U28272 (N_28272,N_26129,N_27293);
or U28273 (N_28273,N_27152,N_26824);
or U28274 (N_28274,N_27960,N_26113);
nand U28275 (N_28275,N_26914,N_27345);
or U28276 (N_28276,N_26838,N_27815);
or U28277 (N_28277,N_27933,N_27695);
and U28278 (N_28278,N_26060,N_26237);
and U28279 (N_28279,N_26260,N_26333);
nor U28280 (N_28280,N_27580,N_27160);
xnor U28281 (N_28281,N_27627,N_27448);
and U28282 (N_28282,N_26862,N_27782);
nand U28283 (N_28283,N_26396,N_26737);
nand U28284 (N_28284,N_26226,N_27275);
xnor U28285 (N_28285,N_26470,N_26435);
and U28286 (N_28286,N_27247,N_26909);
or U28287 (N_28287,N_27146,N_26787);
nand U28288 (N_28288,N_27299,N_26561);
or U28289 (N_28289,N_27231,N_27094);
xnor U28290 (N_28290,N_27449,N_26212);
nor U28291 (N_28291,N_27175,N_27089);
or U28292 (N_28292,N_27019,N_27895);
nand U28293 (N_28293,N_26768,N_26102);
nor U28294 (N_28294,N_27526,N_26742);
xor U28295 (N_28295,N_27246,N_26983);
or U28296 (N_28296,N_27210,N_27523);
and U28297 (N_28297,N_26355,N_27911);
and U28298 (N_28298,N_26464,N_27855);
nor U28299 (N_28299,N_27424,N_26799);
and U28300 (N_28300,N_27475,N_27113);
xnor U28301 (N_28301,N_26160,N_27714);
nor U28302 (N_28302,N_26024,N_27799);
xor U28303 (N_28303,N_27173,N_27446);
xor U28304 (N_28304,N_27910,N_26121);
and U28305 (N_28305,N_27961,N_26825);
xnor U28306 (N_28306,N_26158,N_27693);
and U28307 (N_28307,N_27378,N_26547);
or U28308 (N_28308,N_26006,N_26665);
and U28309 (N_28309,N_27821,N_26751);
nand U28310 (N_28310,N_26439,N_26283);
and U28311 (N_28311,N_26155,N_26588);
or U28312 (N_28312,N_26955,N_26411);
and U28313 (N_28313,N_26436,N_27618);
and U28314 (N_28314,N_26236,N_26418);
xnor U28315 (N_28315,N_27573,N_26280);
xnor U28316 (N_28316,N_27872,N_26122);
nor U28317 (N_28317,N_27194,N_26619);
or U28318 (N_28318,N_26793,N_26127);
and U28319 (N_28319,N_27639,N_26899);
or U28320 (N_28320,N_26419,N_27252);
or U28321 (N_28321,N_26948,N_27791);
nor U28322 (N_28322,N_26481,N_27137);
nand U28323 (N_28323,N_26937,N_27306);
or U28324 (N_28324,N_26395,N_26193);
and U28325 (N_28325,N_27125,N_26258);
nand U28326 (N_28326,N_26189,N_27623);
xnor U28327 (N_28327,N_26152,N_26306);
nand U28328 (N_28328,N_27558,N_26873);
nor U28329 (N_28329,N_26712,N_26566);
nand U28330 (N_28330,N_26697,N_26943);
or U28331 (N_28331,N_27551,N_27522);
and U28332 (N_28332,N_27474,N_26985);
or U28333 (N_28333,N_26987,N_27786);
xnor U28334 (N_28334,N_27962,N_27455);
and U28335 (N_28335,N_26754,N_27077);
nor U28336 (N_28336,N_26437,N_27111);
xor U28337 (N_28337,N_26430,N_27511);
and U28338 (N_28338,N_27442,N_26652);
and U28339 (N_28339,N_26449,N_27068);
nor U28340 (N_28340,N_26705,N_27890);
and U28341 (N_28341,N_27039,N_27298);
nor U28342 (N_28342,N_27422,N_26505);
nor U28343 (N_28343,N_27874,N_27704);
and U28344 (N_28344,N_26651,N_26141);
xnor U28345 (N_28345,N_26059,N_27000);
and U28346 (N_28346,N_27871,N_27250);
or U28347 (N_28347,N_27045,N_27630);
nand U28348 (N_28348,N_26632,N_26649);
and U28349 (N_28349,N_27243,N_26266);
nor U28350 (N_28350,N_27746,N_26270);
xor U28351 (N_28351,N_26479,N_27258);
and U28352 (N_28352,N_27955,N_27807);
and U28353 (N_28353,N_27900,N_26117);
and U28354 (N_28354,N_27758,N_27540);
xnor U28355 (N_28355,N_27603,N_27927);
or U28356 (N_28356,N_27697,N_27478);
xnor U28357 (N_28357,N_27074,N_27638);
nor U28358 (N_28358,N_26605,N_27012);
and U28359 (N_28359,N_26305,N_26757);
nand U28360 (N_28360,N_27646,N_26381);
xnor U28361 (N_28361,N_27621,N_26471);
nand U28362 (N_28362,N_27513,N_26384);
or U28363 (N_28363,N_26095,N_26852);
nor U28364 (N_28364,N_26579,N_26521);
nor U28365 (N_28365,N_27115,N_26176);
and U28366 (N_28366,N_26039,N_27661);
nor U28367 (N_28367,N_27481,N_26223);
and U28368 (N_28368,N_26373,N_26508);
xnor U28369 (N_28369,N_27590,N_26401);
nand U28370 (N_28370,N_27753,N_27347);
xnor U28371 (N_28371,N_26074,N_26887);
or U28372 (N_28372,N_26371,N_27594);
or U28373 (N_28373,N_26607,N_27006);
and U28374 (N_28374,N_26038,N_26101);
and U28375 (N_28375,N_27097,N_27729);
or U28376 (N_28376,N_27941,N_27149);
nor U28377 (N_28377,N_26356,N_26747);
and U28378 (N_28378,N_27588,N_27203);
and U28379 (N_28379,N_26070,N_27622);
or U28380 (N_28380,N_27254,N_26288);
or U28381 (N_28381,N_27967,N_26207);
nand U28382 (N_28382,N_26168,N_26213);
and U28383 (N_28383,N_26885,N_27459);
nand U28384 (N_28384,N_26297,N_26571);
xor U28385 (N_28385,N_26332,N_27408);
or U28386 (N_28386,N_26304,N_26171);
nor U28387 (N_28387,N_26029,N_26228);
and U28388 (N_28388,N_26908,N_26895);
or U28389 (N_28389,N_27245,N_26809);
nor U28390 (N_28390,N_27389,N_26984);
and U28391 (N_28391,N_26195,N_27159);
nor U28392 (N_28392,N_27020,N_27373);
or U28393 (N_28393,N_27591,N_27261);
and U28394 (N_28394,N_26964,N_27864);
nor U28395 (N_28395,N_26210,N_27344);
nand U28396 (N_28396,N_26784,N_26406);
and U28397 (N_28397,N_26836,N_27450);
or U28398 (N_28398,N_27831,N_27812);
nor U28399 (N_28399,N_27999,N_26457);
or U28400 (N_28400,N_26253,N_27184);
nand U28401 (N_28401,N_27841,N_26412);
nor U28402 (N_28402,N_27364,N_27684);
xnor U28403 (N_28403,N_26080,N_27914);
and U28404 (N_28404,N_26774,N_27925);
nor U28405 (N_28405,N_27984,N_26993);
nor U28406 (N_28406,N_26739,N_26284);
and U28407 (N_28407,N_27419,N_27804);
xnor U28408 (N_28408,N_26917,N_26642);
nand U28409 (N_28409,N_27949,N_27809);
nand U28410 (N_28410,N_27754,N_26199);
xnor U28411 (N_28411,N_26146,N_27795);
xor U28412 (N_28412,N_26975,N_26037);
nor U28413 (N_28413,N_27884,N_27223);
or U28414 (N_28414,N_27865,N_27752);
or U28415 (N_28415,N_27439,N_26789);
nor U28416 (N_28416,N_26794,N_26308);
xor U28417 (N_28417,N_26042,N_26726);
and U28418 (N_28418,N_26137,N_26956);
and U28419 (N_28419,N_27988,N_26851);
or U28420 (N_28420,N_27110,N_27153);
and U28421 (N_28421,N_27716,N_26393);
nor U28422 (N_28422,N_27674,N_26702);
nor U28423 (N_28423,N_26164,N_27761);
xnor U28424 (N_28424,N_27690,N_26706);
and U28425 (N_28425,N_26022,N_26915);
or U28426 (N_28426,N_26901,N_27683);
xnor U28427 (N_28427,N_27875,N_26119);
or U28428 (N_28428,N_26541,N_27492);
nor U28429 (N_28429,N_26214,N_26722);
xor U28430 (N_28430,N_27096,N_27996);
and U28431 (N_28431,N_26294,N_27819);
nand U28432 (N_28432,N_27464,N_26612);
nand U28433 (N_28433,N_26971,N_26815);
xnor U28434 (N_28434,N_26216,N_26582);
xnor U28435 (N_28435,N_27671,N_27127);
xnor U28436 (N_28436,N_27981,N_27329);
nand U28437 (N_28437,N_26458,N_26354);
nand U28438 (N_28438,N_26132,N_27310);
nor U28439 (N_28439,N_27670,N_26440);
nor U28440 (N_28440,N_27604,N_26360);
xnor U28441 (N_28441,N_27538,N_26584);
and U28442 (N_28442,N_27458,N_26822);
xnor U28443 (N_28443,N_27438,N_27830);
nor U28444 (N_28444,N_27624,N_27732);
xor U28445 (N_28445,N_27400,N_27057);
xnor U28446 (N_28446,N_26820,N_27477);
and U28447 (N_28447,N_27225,N_27780);
nor U28448 (N_28448,N_27823,N_27073);
nor U28449 (N_28449,N_26805,N_26573);
nand U28450 (N_28450,N_27813,N_26264);
xnor U28451 (N_28451,N_27132,N_27383);
or U28452 (N_28452,N_26604,N_27802);
or U28453 (N_28453,N_27609,N_26593);
nor U28454 (N_28454,N_27748,N_27341);
nor U28455 (N_28455,N_27852,N_26970);
nand U28456 (N_28456,N_26978,N_26431);
or U28457 (N_28457,N_26028,N_26456);
or U28458 (N_28458,N_26200,N_27069);
or U28459 (N_28459,N_26261,N_26474);
xor U28460 (N_28460,N_26586,N_27635);
or U28461 (N_28461,N_26877,N_26054);
nand U28462 (N_28462,N_26321,N_27982);
and U28463 (N_28463,N_26599,N_26869);
and U28464 (N_28464,N_27209,N_26900);
nor U28465 (N_28465,N_26637,N_26082);
and U28466 (N_28466,N_26932,N_26661);
nand U28467 (N_28467,N_27948,N_26327);
nand U28468 (N_28468,N_27648,N_26866);
xor U28469 (N_28469,N_26403,N_26178);
or U28470 (N_28470,N_27416,N_26361);
nor U28471 (N_28471,N_27915,N_26837);
or U28472 (N_28472,N_26215,N_27490);
and U28473 (N_28473,N_26848,N_26351);
xor U28474 (N_28474,N_27994,N_27397);
nand U28475 (N_28475,N_26106,N_27506);
nor U28476 (N_28476,N_27662,N_27276);
nor U28477 (N_28477,N_26762,N_27978);
nand U28478 (N_28478,N_26376,N_27272);
and U28479 (N_28479,N_27681,N_27091);
nand U28480 (N_28480,N_26482,N_26967);
nand U28481 (N_28481,N_27222,N_26750);
and U28482 (N_28482,N_27956,N_26047);
or U28483 (N_28483,N_26961,N_27655);
nand U28484 (N_28484,N_27263,N_27966);
and U28485 (N_28485,N_26766,N_27182);
xor U28486 (N_28486,N_27061,N_26497);
xor U28487 (N_28487,N_27334,N_27968);
or U28488 (N_28488,N_27779,N_26982);
or U28489 (N_28489,N_26477,N_27858);
xor U28490 (N_28490,N_27265,N_27187);
or U28491 (N_28491,N_26081,N_26136);
or U28492 (N_28492,N_27951,N_26709);
and U28493 (N_28493,N_27302,N_27183);
and U28494 (N_28494,N_26585,N_27867);
and U28495 (N_28495,N_27859,N_27769);
xnor U28496 (N_28496,N_27579,N_26220);
nand U28497 (N_28497,N_27390,N_26625);
or U28498 (N_28498,N_27788,N_27126);
or U28499 (N_28499,N_26494,N_27571);
or U28500 (N_28500,N_26578,N_27935);
nand U28501 (N_28501,N_26100,N_27369);
and U28502 (N_28502,N_27820,N_26222);
nor U28503 (N_28503,N_27652,N_27026);
nor U28504 (N_28504,N_27237,N_26153);
nor U28505 (N_28505,N_26083,N_27557);
nor U28506 (N_28506,N_26596,N_26558);
nand U28507 (N_28507,N_26378,N_26560);
nand U28508 (N_28508,N_26574,N_26303);
nor U28509 (N_28509,N_26279,N_27709);
and U28510 (N_28510,N_26916,N_26099);
or U28511 (N_28511,N_26864,N_26329);
nand U28512 (N_28512,N_26727,N_26634);
or U28513 (N_28513,N_27087,N_26148);
and U28514 (N_28514,N_26973,N_27912);
or U28515 (N_28515,N_26224,N_27425);
xnor U28516 (N_28516,N_27940,N_27598);
nand U28517 (N_28517,N_26410,N_26383);
xnor U28518 (N_28518,N_27725,N_27877);
or U28519 (N_28519,N_27507,N_26666);
xnor U28520 (N_28520,N_27443,N_26246);
nand U28521 (N_28521,N_26043,N_26524);
xor U28522 (N_28522,N_27079,N_27359);
nor U28523 (N_28523,N_27101,N_27686);
nand U28524 (N_28524,N_26460,N_26170);
or U28525 (N_28525,N_27691,N_27372);
xor U28526 (N_28526,N_26493,N_27770);
nor U28527 (N_28527,N_27092,N_26935);
or U28528 (N_28528,N_27882,N_26468);
or U28529 (N_28529,N_27643,N_26528);
nand U28530 (N_28530,N_26721,N_27904);
xor U28531 (N_28531,N_27055,N_27849);
xor U28532 (N_28532,N_26902,N_27497);
xor U28533 (N_28533,N_27976,N_27259);
and U28534 (N_28534,N_27705,N_26343);
nor U28535 (N_28535,N_27380,N_27808);
nor U28536 (N_28536,N_26021,N_27251);
xnor U28537 (N_28537,N_26172,N_27700);
xnor U28538 (N_28538,N_27197,N_27750);
or U28539 (N_28539,N_26290,N_27041);
or U28540 (N_28540,N_26245,N_26486);
or U28541 (N_28541,N_27800,N_26472);
nor U28542 (N_28542,N_26238,N_26544);
nand U28543 (N_28543,N_26980,N_27793);
or U28544 (N_28544,N_26600,N_27608);
and U28545 (N_28545,N_27128,N_27512);
or U28546 (N_28546,N_27181,N_26523);
or U28547 (N_28547,N_26720,N_27789);
and U28548 (N_28548,N_26688,N_27634);
xor U28549 (N_28549,N_27322,N_26221);
nand U28550 (N_28550,N_26808,N_27958);
or U28551 (N_28551,N_27320,N_26072);
xor U28552 (N_28552,N_26843,N_27417);
xnor U28553 (N_28553,N_27402,N_27321);
nor U28554 (N_28554,N_27857,N_26953);
nand U28555 (N_28555,N_26345,N_26491);
xnor U28556 (N_28556,N_26366,N_26424);
nand U28557 (N_28557,N_26986,N_27549);
and U28558 (N_28558,N_26502,N_27861);
nor U28559 (N_28559,N_27520,N_27667);
nand U28560 (N_28560,N_26989,N_26810);
nor U28561 (N_28561,N_26804,N_27445);
nor U28562 (N_28562,N_27112,N_27435);
and U28563 (N_28563,N_26663,N_27880);
nand U28564 (N_28564,N_26965,N_27595);
nor U28565 (N_28565,N_27129,N_26128);
nor U28566 (N_28566,N_26180,N_26030);
xor U28567 (N_28567,N_26033,N_27080);
or U28568 (N_28568,N_26618,N_26157);
nand U28569 (N_28569,N_27675,N_26962);
nand U28570 (N_28570,N_27131,N_27688);
nor U28571 (N_28571,N_26723,N_26009);
nand U28572 (N_28572,N_26802,N_27008);
nor U28573 (N_28573,N_26749,N_26476);
or U28574 (N_28574,N_27585,N_26589);
xor U28575 (N_28575,N_27336,N_27340);
and U28576 (N_28576,N_27660,N_26353);
xnor U28577 (N_28577,N_26812,N_27431);
nand U28578 (N_28578,N_27307,N_26951);
nand U28579 (N_28579,N_27399,N_26325);
nand U28580 (N_28580,N_26816,N_27227);
nand U28581 (N_28581,N_27157,N_27143);
xor U28582 (N_28582,N_27742,N_27531);
xnor U28583 (N_28583,N_27834,N_27018);
and U28584 (N_28584,N_27385,N_26539);
nor U28585 (N_28585,N_27379,N_27837);
nor U28586 (N_28586,N_26001,N_26455);
and U28587 (N_28587,N_26888,N_26167);
nor U28588 (N_28588,N_27109,N_26752);
and U28589 (N_28589,N_27542,N_27530);
xnor U28590 (N_28590,N_26265,N_27696);
nor U28591 (N_28591,N_27544,N_26425);
nor U28592 (N_28592,N_26775,N_26441);
nor U28593 (N_28593,N_26025,N_27242);
and U28594 (N_28594,N_26716,N_26149);
xnor U28595 (N_28595,N_26348,N_27384);
and U28596 (N_28596,N_26517,N_26004);
or U28597 (N_28597,N_26646,N_27441);
xnor U28598 (N_28598,N_27102,N_26008);
xnor U28599 (N_28599,N_27316,N_27774);
or U28600 (N_28600,N_26704,N_26611);
nand U28601 (N_28601,N_27850,N_27198);
nor U28602 (N_28602,N_27510,N_27766);
or U28603 (N_28603,N_27308,N_27398);
nand U28604 (N_28604,N_27228,N_26536);
xnor U28605 (N_28605,N_27350,N_26746);
and U28606 (N_28606,N_27296,N_26263);
nand U28607 (N_28607,N_27713,N_27230);
and U28608 (N_28608,N_27637,N_26992);
or U28609 (N_28609,N_26850,N_27462);
or U28610 (N_28610,N_27003,N_27304);
nor U28611 (N_28611,N_27751,N_27719);
nor U28612 (N_28612,N_27586,N_26654);
or U28613 (N_28613,N_27888,N_26271);
nand U28614 (N_28614,N_26324,N_26034);
nand U28615 (N_28615,N_26756,N_27392);
or U28616 (N_28616,N_26459,N_27046);
and U28617 (N_28617,N_26291,N_26390);
nand U28618 (N_28618,N_27224,N_27893);
and U28619 (N_28619,N_26830,N_26254);
nand U28620 (N_28620,N_26017,N_26680);
and U28621 (N_28621,N_27734,N_27559);
xor U28622 (N_28622,N_27845,N_27894);
nor U28623 (N_28623,N_27367,N_27324);
nor U28624 (N_28624,N_26352,N_26748);
nor U28625 (N_28625,N_26187,N_27653);
and U28626 (N_28626,N_26108,N_27410);
and U28627 (N_28627,N_27174,N_26126);
xor U28628 (N_28628,N_27840,N_26309);
or U28629 (N_28629,N_26679,N_26911);
nor U28630 (N_28630,N_27777,N_27765);
or U28631 (N_28631,N_27665,N_27332);
xor U28632 (N_28632,N_27775,N_26930);
nand U28633 (N_28633,N_27274,N_26630);
or U28634 (N_28634,N_26856,N_27932);
nand U28635 (N_28635,N_27119,N_27574);
nor U28636 (N_28636,N_27909,N_26450);
xnor U28637 (N_28637,N_26078,N_26623);
nor U28638 (N_28638,N_26296,N_27429);
and U28639 (N_28639,N_27778,N_26445);
nand U28640 (N_28640,N_27556,N_26620);
nand U28641 (N_28641,N_27772,N_27616);
nand U28642 (N_28642,N_27889,N_26731);
and U28643 (N_28643,N_26452,N_27062);
nand U28644 (N_28644,N_27599,N_27552);
xnor U28645 (N_28645,N_26897,N_27139);
nor U28646 (N_28646,N_26124,N_26420);
xnor U28647 (N_28647,N_27169,N_27099);
nand U28648 (N_28648,N_27134,N_26495);
or U28649 (N_28649,N_26496,N_26949);
nor U28650 (N_28650,N_27827,N_27457);
or U28651 (N_28651,N_27575,N_27747);
or U28652 (N_28652,N_27860,N_27677);
nand U28653 (N_28653,N_26894,N_27180);
xnor U28654 (N_28654,N_27738,N_27602);
nor U28655 (N_28655,N_26012,N_26145);
nor U28656 (N_28656,N_27407,N_27712);
nand U28657 (N_28657,N_27032,N_27666);
nand U28658 (N_28658,N_27577,N_26317);
nand U28659 (N_28659,N_26442,N_26940);
nand U28660 (N_28660,N_27106,N_27421);
nor U28661 (N_28661,N_26192,N_26131);
nor U28662 (N_28662,N_27903,N_27028);
and U28663 (N_28663,N_27561,N_27412);
and U28664 (N_28664,N_26446,N_26963);
nor U28665 (N_28665,N_26664,N_26501);
nand U28666 (N_28666,N_26239,N_26295);
nor U28667 (N_28667,N_26090,N_27004);
nand U28668 (N_28668,N_26185,N_26392);
and U28669 (N_28669,N_26656,N_26818);
xnor U28670 (N_28670,N_26507,N_27792);
nand U28671 (N_28671,N_26769,N_26061);
or U28672 (N_28672,N_26289,N_26960);
xnor U28673 (N_28673,N_27629,N_26591);
nand U28674 (N_28674,N_26219,N_27030);
nand U28675 (N_28675,N_26282,N_26125);
nand U28676 (N_28676,N_26912,N_26298);
xnor U28677 (N_28677,N_27664,N_26650);
and U28678 (N_28678,N_27572,N_27811);
xor U28679 (N_28679,N_26803,N_27581);
nor U28680 (N_28680,N_27829,N_27728);
or U28681 (N_28681,N_27548,N_27001);
nor U28682 (N_28682,N_26765,N_27485);
nor U28683 (N_28683,N_27311,N_27226);
and U28684 (N_28684,N_27043,N_26891);
and U28685 (N_28685,N_26741,N_27640);
or U28686 (N_28686,N_27564,N_26839);
xnor U28687 (N_28687,N_26018,N_27049);
and U28688 (N_28688,N_27626,N_26196);
xor U28689 (N_28689,N_27178,N_27727);
nand U28690 (N_28690,N_27214,N_26991);
nand U28691 (N_28691,N_26827,N_27596);
or U28692 (N_28692,N_27972,N_27241);
nand U28693 (N_28693,N_26350,N_27200);
or U28694 (N_28694,N_26840,N_27319);
nand U28695 (N_28695,N_26169,N_26483);
nand U28696 (N_28696,N_26094,N_26714);
xnor U28697 (N_28697,N_27692,N_27612);
and U28698 (N_28698,N_27897,N_27401);
xnor U28699 (N_28699,N_26394,N_27376);
or U28700 (N_28700,N_27916,N_27022);
or U28701 (N_28701,N_26257,N_27614);
nand U28702 (N_28702,N_27205,N_27929);
xor U28703 (N_28703,N_27536,N_26640);
xor U28704 (N_28704,N_26036,N_26563);
nor U28705 (N_28705,N_27480,N_27992);
xnor U28706 (N_28706,N_27255,N_27122);
and U28707 (N_28707,N_27179,N_26628);
xnor U28708 (N_28708,N_27342,N_26905);
nand U28709 (N_28709,N_26609,N_27739);
and U28710 (N_28710,N_26087,N_27562);
nor U28711 (N_28711,N_27944,N_27768);
nor U28712 (N_28712,N_27317,N_27413);
nand U28713 (N_28713,N_26773,N_27189);
nand U28714 (N_28714,N_27620,N_27928);
nor U28715 (N_28715,N_27482,N_27658);
nor U28716 (N_28716,N_27108,N_27803);
or U28717 (N_28717,N_27172,N_26007);
nor U28718 (N_28718,N_26421,N_27196);
xnor U28719 (N_28719,N_26500,N_27814);
nor U28720 (N_28720,N_26581,N_27075);
and U28721 (N_28721,N_27870,N_27453);
xnor U28722 (N_28722,N_27375,N_27356);
nand U28723 (N_28723,N_26635,N_27516);
xor U28724 (N_28724,N_26275,N_26382);
and U28725 (N_28725,N_27632,N_26667);
or U28726 (N_28726,N_26783,N_26614);
xor U28727 (N_28727,N_26516,N_27355);
and U28728 (N_28728,N_27193,N_26924);
xor U28729 (N_28729,N_26554,N_27945);
or U28730 (N_28730,N_26027,N_26944);
nand U28731 (N_28731,N_26846,N_27504);
nor U28732 (N_28732,N_27295,N_26143);
and U28733 (N_28733,N_26011,N_26999);
nor U28734 (N_28734,N_27839,N_26423);
nand U28735 (N_28735,N_27454,N_26307);
nand U28736 (N_28736,N_27282,N_26535);
xnor U28737 (N_28737,N_27052,N_27919);
or U28738 (N_28738,N_27059,N_27232);
and U28739 (N_28739,N_26252,N_26831);
nand U28740 (N_28740,N_27701,N_26320);
nand U28741 (N_28741,N_26717,N_27539);
or U28742 (N_28742,N_27088,N_27931);
or U28743 (N_28743,N_27805,N_27560);
or U28744 (N_28744,N_26409,N_27204);
xnor U28745 (N_28745,N_27737,N_26675);
or U28746 (N_28746,N_26256,N_27524);
xnor U28747 (N_28747,N_26551,N_26893);
and U28748 (N_28748,N_27007,N_26138);
nor U28749 (N_28749,N_26876,N_27862);
xnor U28750 (N_28750,N_27702,N_26595);
xnor U28751 (N_28751,N_27090,N_27615);
nor U28752 (N_28752,N_26684,N_27171);
and U28753 (N_28753,N_26274,N_26795);
and U28754 (N_28754,N_26786,N_27358);
and U28755 (N_28755,N_27787,N_27281);
nor U28756 (N_28756,N_27679,N_27280);
or U28757 (N_28757,N_26337,N_26035);
nor U28758 (N_28758,N_26230,N_26241);
and U28759 (N_28759,N_26053,N_26323);
nand U28760 (N_28760,N_27902,N_26175);
and U28761 (N_28761,N_26165,N_26314);
or U28762 (N_28762,N_27953,N_26326);
or U28763 (N_28763,N_27405,N_26597);
xnor U28764 (N_28764,N_26206,N_26374);
xnor U28765 (N_28765,N_26194,N_27592);
xnor U28766 (N_28766,N_26525,N_26870);
or U28767 (N_28767,N_26957,N_26162);
nor U28768 (N_28768,N_26301,N_27213);
and U28769 (N_28769,N_27491,N_27440);
nand U28770 (N_28770,N_26426,N_27195);
nand U28771 (N_28771,N_26380,N_27116);
xnor U28772 (N_28772,N_26386,N_26142);
xor U28773 (N_28773,N_26522,N_27283);
nor U28774 (N_28774,N_26685,N_26689);
or U28775 (N_28775,N_26678,N_27447);
nand U28776 (N_28776,N_27711,N_27856);
nor U28777 (N_28777,N_26644,N_26760);
xnor U28778 (N_28778,N_26096,N_27117);
and U28779 (N_28779,N_27406,N_27605);
and U28780 (N_28780,N_27698,N_26020);
xor U28781 (N_28781,N_26671,N_27494);
and U28782 (N_28782,N_26417,N_27473);
nand U28783 (N_28783,N_27234,N_27730);
nand U28784 (N_28784,N_27600,N_26867);
nor U28785 (N_28785,N_27892,N_26109);
and U28786 (N_28786,N_26928,N_26092);
nand U28787 (N_28787,N_27720,N_26135);
and U28788 (N_28788,N_27047,N_26933);
xnor U28789 (N_28789,N_27946,N_26233);
nand U28790 (N_28790,N_26855,N_27343);
or U28791 (N_28791,N_27498,N_27466);
and U28792 (N_28792,N_26375,N_26334);
nor U28793 (N_28793,N_26734,N_26732);
and U28794 (N_28794,N_26339,N_26488);
nor U28795 (N_28795,N_26776,N_26791);
xnor U28796 (N_28796,N_26402,N_27145);
xor U28797 (N_28797,N_27989,N_27123);
xor U28798 (N_28798,N_26829,N_26400);
xor U28799 (N_28799,N_27707,N_27776);
or U28800 (N_28800,N_27218,N_27689);
and U28801 (N_28801,N_27357,N_26273);
and U28802 (N_28802,N_27423,N_26529);
nor U28803 (N_28803,N_27617,N_26562);
nor U28804 (N_28804,N_26878,N_26163);
or U28805 (N_28805,N_27314,N_26023);
or U28806 (N_28806,N_27130,N_27582);
nor U28807 (N_28807,N_27238,N_26703);
nand U28808 (N_28808,N_27649,N_27908);
and U28809 (N_28809,N_26111,N_27957);
xor U28810 (N_28810,N_26833,N_27937);
or U28811 (N_28811,N_26186,N_26587);
xor U28812 (N_28812,N_27138,N_27312);
and U28813 (N_28813,N_26755,N_27470);
nand U28814 (N_28814,N_26293,N_26871);
or U28815 (N_28815,N_27987,N_26191);
or U28816 (N_28816,N_26875,N_27081);
nor U28817 (N_28817,N_27023,N_26447);
nor U28818 (N_28818,N_26330,N_26633);
xnor U28819 (N_28819,N_26065,N_27980);
nand U28820 (N_28820,N_27086,N_26218);
and U28821 (N_28821,N_27016,N_26939);
or U28822 (N_28822,N_27100,N_27190);
and U28823 (N_28823,N_27784,N_26358);
and U28824 (N_28824,N_27471,N_26540);
nand U28825 (N_28825,N_26050,N_26811);
nand U28826 (N_28826,N_27033,N_26364);
nor U28827 (N_28827,N_26857,N_27567);
nand U28828 (N_28828,N_26610,N_27148);
nand U28829 (N_28829,N_27659,N_26473);
nand U28830 (N_28830,N_27717,N_26565);
xor U28831 (N_28831,N_27147,N_27505);
nand U28832 (N_28832,N_27093,N_26147);
xor U28833 (N_28833,N_26197,N_27607);
nand U28834 (N_28834,N_27244,N_26919);
xnor U28835 (N_28835,N_26077,N_27584);
xor U28836 (N_28836,N_26583,N_27362);
or U28837 (N_28837,N_27611,N_27387);
xnor U28838 (N_28838,N_27212,N_26312);
or U28839 (N_28839,N_26357,N_27037);
xor U28840 (N_28840,N_26708,N_27427);
nor U28841 (N_28841,N_26844,N_26344);
nor U28842 (N_28842,N_27669,N_26603);
or U28843 (N_28843,N_26555,N_27920);
xor U28844 (N_28844,N_27703,N_27370);
xor U28845 (N_28845,N_26515,N_26014);
or U28846 (N_28846,N_26764,N_27452);
and U28847 (N_28847,N_27749,N_26002);
and U28848 (N_28848,N_26139,N_27034);
nand U28849 (N_28849,N_26559,N_26629);
or U28850 (N_28850,N_26676,N_26005);
and U28851 (N_28851,N_27922,N_27042);
nand U28852 (N_28852,N_27723,N_26134);
nor U28853 (N_28853,N_26526,N_26242);
or U28854 (N_28854,N_27415,N_26592);
xor U28855 (N_28855,N_26979,N_27216);
or U28856 (N_28856,N_27650,N_27268);
nor U28857 (N_28857,N_27070,N_26302);
and U28858 (N_28858,N_26913,N_27273);
nor U28859 (N_28859,N_27722,N_27569);
xnor U28860 (N_28860,N_27469,N_26182);
or U28861 (N_28861,N_26778,N_26572);
nand U28862 (N_28862,N_26003,N_26920);
xnor U28863 (N_28863,N_26780,N_26300);
nand U28864 (N_28864,N_26379,N_26772);
nand U28865 (N_28865,N_26660,N_27767);
and U28866 (N_28866,N_27672,N_27848);
and U28867 (N_28867,N_27339,N_27294);
and U28868 (N_28868,N_27798,N_27105);
and U28869 (N_28869,N_26569,N_26657);
xnor U28870 (N_28870,N_26340,N_26759);
nor U28871 (N_28871,N_27936,N_27514);
nor U28872 (N_28872,N_27264,N_26490);
nor U28873 (N_28873,N_26872,N_27056);
and U28874 (N_28874,N_27771,N_26639);
and U28875 (N_28875,N_26262,N_27613);
nor U28876 (N_28876,N_27065,N_26890);
xnor U28877 (N_28877,N_27881,N_26250);
nand U28878 (N_28878,N_26000,N_27024);
and U28879 (N_28879,N_27952,N_27997);
nand U28880 (N_28880,N_27229,N_27348);
and U28881 (N_28881,N_26453,N_26527);
or U28882 (N_28882,N_26925,N_26444);
or U28883 (N_28883,N_26045,N_27468);
and U28884 (N_28884,N_27576,N_27444);
or U28885 (N_28885,N_27418,N_27374);
xnor U28886 (N_28886,N_26058,N_26966);
nor U28887 (N_28887,N_27067,N_27682);
nand U28888 (N_28888,N_26489,N_27678);
and U28889 (N_28889,N_26694,N_26788);
and U28890 (N_28890,N_27763,N_26710);
nor U28891 (N_28891,N_26451,N_27486);
nand U28892 (N_28892,N_27303,N_27906);
and U28893 (N_28893,N_27833,N_27021);
and U28894 (N_28894,N_26669,N_27035);
or U28895 (N_28895,N_27896,N_27501);
xor U28896 (N_28896,N_27140,N_26248);
xnor U28897 (N_28897,N_27687,N_27699);
xnor U28898 (N_28898,N_27338,N_26549);
and U28899 (N_28899,N_26211,N_26763);
xor U28900 (N_28900,N_26994,N_27518);
nand U28901 (N_28901,N_26568,N_26485);
and U28902 (N_28902,N_27851,N_27136);
nor U28903 (N_28903,N_26736,N_27240);
and U28904 (N_28904,N_26674,N_27170);
or U28905 (N_28905,N_27066,N_26745);
or U28906 (N_28906,N_26249,N_27328);
nor U28907 (N_28907,N_26668,N_27318);
xor U28908 (N_28908,N_26154,N_26462);
nor U28909 (N_28909,N_26385,N_27636);
nand U28910 (N_28910,N_26098,N_27934);
nand U28911 (N_28911,N_26969,N_26068);
or U28912 (N_28912,N_26621,N_26879);
nand U28913 (N_28913,N_27631,N_26110);
and U28914 (N_28914,N_26626,N_26662);
and U28915 (N_28915,N_26608,N_26673);
and U28916 (N_28916,N_26049,N_27993);
nor U28917 (N_28917,N_26753,N_26190);
or U28918 (N_28918,N_26735,N_27554);
nor U28919 (N_28919,N_27098,N_26860);
nor U28920 (N_28920,N_27327,N_27260);
nor U28921 (N_28921,N_26849,N_27495);
and U28922 (N_28922,N_26140,N_26761);
xnor U28923 (N_28923,N_27975,N_27278);
nand U28924 (N_28924,N_26602,N_26044);
or U28925 (N_28925,N_26534,N_26156);
or U28926 (N_28926,N_27071,N_26858);
xnor U28927 (N_28927,N_26798,N_27396);
or U28928 (N_28928,N_26235,N_27467);
nor U28929 (N_28929,N_26807,N_27868);
and U28930 (N_28930,N_26062,N_27456);
nand U28931 (N_28931,N_26067,N_26693);
xor U28932 (N_28932,N_26819,N_26779);
or U28933 (N_28933,N_26976,N_27325);
xor U28934 (N_28934,N_26201,N_27167);
nand U28935 (N_28935,N_27866,N_27543);
and U28936 (N_28936,N_26733,N_27360);
nor U28937 (N_28937,N_26492,N_27271);
nor U28938 (N_28938,N_27217,N_27054);
or U28939 (N_28939,N_26240,N_27158);
xnor U28940 (N_28940,N_27899,N_27563);
and U28941 (N_28941,N_26998,N_27741);
nor U28942 (N_28942,N_26346,N_26151);
nand U28943 (N_28943,N_26469,N_27917);
and U28944 (N_28944,N_26173,N_26834);
xor U28945 (N_28945,N_26533,N_26071);
nand U28946 (N_28946,N_26923,N_27721);
nor U28947 (N_28947,N_26513,N_27323);
and U28948 (N_28948,N_26695,N_27532);
or U28949 (N_28949,N_26161,N_27476);
or U28950 (N_28950,N_26272,N_26631);
or U28951 (N_28951,N_26349,N_27472);
xnor U28952 (N_28952,N_26405,N_26328);
nand U28953 (N_28953,N_26594,N_26066);
xor U28954 (N_28954,N_26946,N_26670);
and U28955 (N_28955,N_27036,N_26995);
nor U28956 (N_28956,N_27534,N_26465);
or U28957 (N_28957,N_26335,N_27601);
nand U28958 (N_28958,N_26929,N_27657);
and U28959 (N_28959,N_27760,N_26692);
nor U28960 (N_28960,N_26427,N_27550);
nor U28961 (N_28961,N_27078,N_27546);
nand U28962 (N_28962,N_26277,N_26730);
or U28963 (N_28963,N_27371,N_26865);
and U28964 (N_28964,N_26069,N_26641);
xnor U28965 (N_28965,N_27436,N_27708);
or U28966 (N_28966,N_26880,N_26363);
or U28967 (N_28967,N_26958,N_27755);
nor U28968 (N_28968,N_26648,N_26548);
and U28969 (N_28969,N_26013,N_26996);
nand U28970 (N_28970,N_26814,N_27351);
nor U28971 (N_28971,N_27918,N_26567);
nand U28972 (N_28972,N_27202,N_27816);
or U28973 (N_28973,N_26370,N_26438);
nand U28974 (N_28974,N_26046,N_27810);
and U28975 (N_28975,N_26336,N_27589);
nand U28976 (N_28976,N_27206,N_27663);
and U28977 (N_28977,N_27382,N_26947);
xor U28978 (N_28978,N_26278,N_26828);
nor U28979 (N_28979,N_26428,N_27832);
xor U28980 (N_28980,N_27502,N_27151);
nand U28981 (N_28981,N_26550,N_27969);
xnor U28982 (N_28982,N_26841,N_27363);
nand U28983 (N_28983,N_26771,N_27736);
or U28984 (N_28984,N_27337,N_27191);
nor U28985 (N_28985,N_27414,N_27854);
or U28986 (N_28986,N_27528,N_26202);
or U28987 (N_28987,N_26823,N_26655);
xnor U28988 (N_28988,N_27331,N_26903);
and U28989 (N_28989,N_27192,N_26116);
and U28990 (N_28990,N_27300,N_27645);
nand U28991 (N_28991,N_27393,N_27651);
nand U28992 (N_28992,N_27628,N_26700);
nor U28993 (N_28993,N_27394,N_26790);
xnor U28994 (N_28994,N_27610,N_27177);
xnor U28995 (N_28995,N_27411,N_27565);
and U28996 (N_28996,N_27726,N_27986);
or U28997 (N_28997,N_27529,N_27301);
nand U28998 (N_28998,N_26188,N_27235);
nand U28999 (N_28999,N_27762,N_26362);
and U29000 (N_29000,N_27346,N_27468);
and U29001 (N_29001,N_27813,N_26416);
xnor U29002 (N_29002,N_27743,N_27504);
xor U29003 (N_29003,N_26921,N_26400);
nand U29004 (N_29004,N_26399,N_27386);
xor U29005 (N_29005,N_27749,N_27213);
nand U29006 (N_29006,N_26459,N_26887);
xnor U29007 (N_29007,N_26105,N_26027);
nor U29008 (N_29008,N_26560,N_26988);
xnor U29009 (N_29009,N_26268,N_26675);
nor U29010 (N_29010,N_27032,N_27940);
nor U29011 (N_29011,N_26044,N_26755);
or U29012 (N_29012,N_27640,N_27779);
or U29013 (N_29013,N_27535,N_27001);
and U29014 (N_29014,N_26562,N_26248);
nand U29015 (N_29015,N_27742,N_27086);
xor U29016 (N_29016,N_26352,N_27281);
nor U29017 (N_29017,N_26151,N_26574);
and U29018 (N_29018,N_26548,N_26768);
nand U29019 (N_29019,N_26818,N_27554);
xnor U29020 (N_29020,N_26661,N_27818);
and U29021 (N_29021,N_26804,N_26964);
or U29022 (N_29022,N_27857,N_26316);
or U29023 (N_29023,N_27115,N_27191);
xnor U29024 (N_29024,N_27555,N_26906);
xnor U29025 (N_29025,N_27324,N_27026);
and U29026 (N_29026,N_26028,N_27585);
or U29027 (N_29027,N_27465,N_26324);
or U29028 (N_29028,N_27315,N_27964);
and U29029 (N_29029,N_26009,N_26025);
nand U29030 (N_29030,N_26792,N_27093);
and U29031 (N_29031,N_26309,N_26005);
or U29032 (N_29032,N_26508,N_27908);
nor U29033 (N_29033,N_26747,N_26477);
xnor U29034 (N_29034,N_26277,N_26254);
and U29035 (N_29035,N_27744,N_27129);
nand U29036 (N_29036,N_26641,N_27812);
nor U29037 (N_29037,N_26098,N_26192);
and U29038 (N_29038,N_26426,N_26811);
and U29039 (N_29039,N_26911,N_27254);
nor U29040 (N_29040,N_27426,N_27858);
xnor U29041 (N_29041,N_26393,N_26190);
nand U29042 (N_29042,N_26488,N_27679);
xnor U29043 (N_29043,N_26816,N_27527);
or U29044 (N_29044,N_26710,N_26377);
and U29045 (N_29045,N_26601,N_26404);
and U29046 (N_29046,N_27459,N_27055);
xnor U29047 (N_29047,N_26570,N_27557);
xnor U29048 (N_29048,N_26141,N_27384);
nand U29049 (N_29049,N_26177,N_26048);
and U29050 (N_29050,N_27044,N_26086);
or U29051 (N_29051,N_26989,N_27091);
xnor U29052 (N_29052,N_27295,N_26806);
or U29053 (N_29053,N_26872,N_27905);
nand U29054 (N_29054,N_26899,N_27587);
or U29055 (N_29055,N_26347,N_26781);
nor U29056 (N_29056,N_26782,N_27866);
and U29057 (N_29057,N_26043,N_27503);
xnor U29058 (N_29058,N_26030,N_26398);
nand U29059 (N_29059,N_26087,N_27515);
nor U29060 (N_29060,N_26234,N_26686);
and U29061 (N_29061,N_27770,N_27494);
and U29062 (N_29062,N_26376,N_27291);
nand U29063 (N_29063,N_26830,N_26313);
nand U29064 (N_29064,N_26343,N_27903);
nand U29065 (N_29065,N_26689,N_26302);
nand U29066 (N_29066,N_27826,N_27612);
and U29067 (N_29067,N_27209,N_27350);
or U29068 (N_29068,N_26864,N_27590);
and U29069 (N_29069,N_27123,N_26089);
xnor U29070 (N_29070,N_27004,N_27491);
or U29071 (N_29071,N_27040,N_26787);
xnor U29072 (N_29072,N_26549,N_26739);
xnor U29073 (N_29073,N_27014,N_27899);
nand U29074 (N_29074,N_26623,N_27464);
or U29075 (N_29075,N_27303,N_27173);
xnor U29076 (N_29076,N_27978,N_27312);
xnor U29077 (N_29077,N_26023,N_27532);
and U29078 (N_29078,N_27637,N_26744);
and U29079 (N_29079,N_27196,N_26406);
nand U29080 (N_29080,N_27240,N_26851);
nand U29081 (N_29081,N_27867,N_26209);
or U29082 (N_29082,N_26752,N_26470);
and U29083 (N_29083,N_26174,N_26309);
or U29084 (N_29084,N_26663,N_27340);
and U29085 (N_29085,N_26364,N_26921);
or U29086 (N_29086,N_27287,N_26870);
xnor U29087 (N_29087,N_26289,N_26435);
xnor U29088 (N_29088,N_27256,N_26076);
or U29089 (N_29089,N_27877,N_26183);
xnor U29090 (N_29090,N_26228,N_26964);
or U29091 (N_29091,N_27241,N_27654);
xor U29092 (N_29092,N_27526,N_27668);
xor U29093 (N_29093,N_27404,N_27771);
xnor U29094 (N_29094,N_27351,N_26257);
nor U29095 (N_29095,N_26324,N_27545);
or U29096 (N_29096,N_27775,N_27699);
nor U29097 (N_29097,N_27251,N_26272);
or U29098 (N_29098,N_27990,N_26460);
or U29099 (N_29099,N_27886,N_27785);
or U29100 (N_29100,N_27605,N_27915);
xnor U29101 (N_29101,N_27946,N_27443);
or U29102 (N_29102,N_27780,N_27975);
nand U29103 (N_29103,N_27699,N_26972);
nand U29104 (N_29104,N_27309,N_27647);
and U29105 (N_29105,N_26773,N_26481);
and U29106 (N_29106,N_26279,N_26319);
xnor U29107 (N_29107,N_27800,N_27435);
or U29108 (N_29108,N_26764,N_27331);
and U29109 (N_29109,N_26518,N_26464);
or U29110 (N_29110,N_26364,N_27142);
nand U29111 (N_29111,N_26301,N_26982);
xor U29112 (N_29112,N_26312,N_27248);
xor U29113 (N_29113,N_27199,N_27707);
xor U29114 (N_29114,N_26783,N_27186);
xnor U29115 (N_29115,N_26994,N_27483);
nand U29116 (N_29116,N_26517,N_26150);
xor U29117 (N_29117,N_26637,N_27413);
xnor U29118 (N_29118,N_27307,N_27619);
nand U29119 (N_29119,N_26263,N_27101);
or U29120 (N_29120,N_27578,N_27180);
and U29121 (N_29121,N_26410,N_26772);
nor U29122 (N_29122,N_26849,N_27778);
nand U29123 (N_29123,N_27974,N_27573);
nand U29124 (N_29124,N_27107,N_26583);
nor U29125 (N_29125,N_26050,N_27026);
xnor U29126 (N_29126,N_26332,N_26733);
and U29127 (N_29127,N_27188,N_26014);
and U29128 (N_29128,N_27945,N_26286);
nor U29129 (N_29129,N_27813,N_27420);
and U29130 (N_29130,N_26995,N_26064);
or U29131 (N_29131,N_26647,N_26530);
xnor U29132 (N_29132,N_27713,N_27007);
nand U29133 (N_29133,N_26580,N_27817);
and U29134 (N_29134,N_27026,N_26799);
nand U29135 (N_29135,N_27309,N_26493);
or U29136 (N_29136,N_27632,N_27612);
nor U29137 (N_29137,N_27654,N_27814);
nand U29138 (N_29138,N_26794,N_27145);
nand U29139 (N_29139,N_27781,N_27069);
or U29140 (N_29140,N_27983,N_27993);
and U29141 (N_29141,N_26766,N_26293);
and U29142 (N_29142,N_27231,N_27693);
or U29143 (N_29143,N_27239,N_27191);
xor U29144 (N_29144,N_26471,N_27659);
and U29145 (N_29145,N_27677,N_27902);
nor U29146 (N_29146,N_26935,N_27837);
and U29147 (N_29147,N_26175,N_26022);
nand U29148 (N_29148,N_26463,N_26563);
or U29149 (N_29149,N_27082,N_26743);
xor U29150 (N_29150,N_27806,N_27898);
xnor U29151 (N_29151,N_27746,N_26481);
and U29152 (N_29152,N_26714,N_26496);
nor U29153 (N_29153,N_26588,N_26764);
nor U29154 (N_29154,N_27959,N_26606);
or U29155 (N_29155,N_27811,N_26761);
xnor U29156 (N_29156,N_26136,N_26714);
xnor U29157 (N_29157,N_27703,N_26296);
and U29158 (N_29158,N_27796,N_27427);
nor U29159 (N_29159,N_26000,N_26548);
and U29160 (N_29160,N_27546,N_27873);
and U29161 (N_29161,N_26908,N_27905);
or U29162 (N_29162,N_27296,N_26701);
nor U29163 (N_29163,N_27961,N_27505);
and U29164 (N_29164,N_27243,N_26256);
xor U29165 (N_29165,N_26043,N_26784);
or U29166 (N_29166,N_26278,N_26940);
nand U29167 (N_29167,N_26905,N_26465);
or U29168 (N_29168,N_26363,N_27975);
nand U29169 (N_29169,N_26807,N_26192);
nor U29170 (N_29170,N_27351,N_26024);
xnor U29171 (N_29171,N_27575,N_27335);
nand U29172 (N_29172,N_26977,N_26647);
and U29173 (N_29173,N_26148,N_26111);
nor U29174 (N_29174,N_26758,N_26694);
or U29175 (N_29175,N_26943,N_27686);
xnor U29176 (N_29176,N_27421,N_26854);
nand U29177 (N_29177,N_26451,N_27803);
xor U29178 (N_29178,N_26063,N_27735);
or U29179 (N_29179,N_27878,N_27359);
xor U29180 (N_29180,N_26225,N_27587);
and U29181 (N_29181,N_26406,N_26421);
or U29182 (N_29182,N_27441,N_26028);
or U29183 (N_29183,N_26712,N_26221);
nand U29184 (N_29184,N_27757,N_26254);
and U29185 (N_29185,N_26993,N_26696);
nor U29186 (N_29186,N_27219,N_27163);
and U29187 (N_29187,N_26052,N_27810);
xnor U29188 (N_29188,N_27406,N_27728);
xnor U29189 (N_29189,N_27128,N_26231);
nor U29190 (N_29190,N_27734,N_26778);
or U29191 (N_29191,N_27661,N_26169);
nor U29192 (N_29192,N_27411,N_27156);
and U29193 (N_29193,N_27774,N_26668);
and U29194 (N_29194,N_26986,N_26877);
or U29195 (N_29195,N_26846,N_27515);
or U29196 (N_29196,N_27798,N_27645);
or U29197 (N_29197,N_26760,N_26145);
nand U29198 (N_29198,N_26894,N_27211);
or U29199 (N_29199,N_26243,N_27334);
xnor U29200 (N_29200,N_26301,N_27029);
nor U29201 (N_29201,N_27977,N_27488);
xor U29202 (N_29202,N_27419,N_26678);
and U29203 (N_29203,N_27578,N_26751);
and U29204 (N_29204,N_26373,N_27867);
nand U29205 (N_29205,N_27443,N_27048);
and U29206 (N_29206,N_26831,N_27623);
xor U29207 (N_29207,N_26946,N_26057);
nand U29208 (N_29208,N_26637,N_27845);
or U29209 (N_29209,N_27087,N_26796);
and U29210 (N_29210,N_27607,N_26216);
nor U29211 (N_29211,N_26029,N_26456);
and U29212 (N_29212,N_27193,N_26956);
and U29213 (N_29213,N_26877,N_27281);
nor U29214 (N_29214,N_26946,N_26028);
nand U29215 (N_29215,N_27167,N_26728);
or U29216 (N_29216,N_27013,N_26916);
nor U29217 (N_29217,N_26817,N_27826);
and U29218 (N_29218,N_26604,N_26695);
or U29219 (N_29219,N_27746,N_27483);
xnor U29220 (N_29220,N_27710,N_27769);
nand U29221 (N_29221,N_27048,N_26780);
xnor U29222 (N_29222,N_26702,N_26287);
and U29223 (N_29223,N_27885,N_26515);
and U29224 (N_29224,N_27245,N_26923);
nand U29225 (N_29225,N_27043,N_26633);
or U29226 (N_29226,N_27665,N_27884);
nor U29227 (N_29227,N_27561,N_27096);
and U29228 (N_29228,N_27170,N_27213);
nand U29229 (N_29229,N_26065,N_27466);
or U29230 (N_29230,N_26804,N_26220);
and U29231 (N_29231,N_27551,N_26161);
nor U29232 (N_29232,N_27744,N_26181);
or U29233 (N_29233,N_26412,N_26292);
nand U29234 (N_29234,N_26514,N_26198);
or U29235 (N_29235,N_26061,N_26695);
nand U29236 (N_29236,N_27622,N_27089);
or U29237 (N_29237,N_26181,N_27271);
and U29238 (N_29238,N_26016,N_27663);
and U29239 (N_29239,N_27994,N_27804);
and U29240 (N_29240,N_26470,N_27144);
nor U29241 (N_29241,N_27663,N_27273);
and U29242 (N_29242,N_27585,N_26917);
xnor U29243 (N_29243,N_27186,N_26065);
nand U29244 (N_29244,N_27603,N_26977);
nor U29245 (N_29245,N_27914,N_26906);
or U29246 (N_29246,N_26924,N_26027);
nor U29247 (N_29247,N_26211,N_26184);
and U29248 (N_29248,N_26950,N_27465);
or U29249 (N_29249,N_26873,N_27740);
nand U29250 (N_29250,N_26662,N_27639);
and U29251 (N_29251,N_26724,N_26919);
or U29252 (N_29252,N_27024,N_26610);
or U29253 (N_29253,N_27531,N_27982);
nand U29254 (N_29254,N_26440,N_27233);
xor U29255 (N_29255,N_26569,N_27937);
xnor U29256 (N_29256,N_27225,N_26771);
xnor U29257 (N_29257,N_26819,N_27807);
nand U29258 (N_29258,N_27257,N_26837);
or U29259 (N_29259,N_27214,N_26417);
nor U29260 (N_29260,N_27682,N_27572);
or U29261 (N_29261,N_26253,N_27720);
xnor U29262 (N_29262,N_27149,N_27743);
and U29263 (N_29263,N_26651,N_26840);
nand U29264 (N_29264,N_27079,N_26437);
or U29265 (N_29265,N_27104,N_27685);
nand U29266 (N_29266,N_26711,N_26405);
nor U29267 (N_29267,N_27649,N_27344);
nand U29268 (N_29268,N_27911,N_26150);
nor U29269 (N_29269,N_27292,N_27113);
and U29270 (N_29270,N_27549,N_26719);
and U29271 (N_29271,N_26629,N_27843);
and U29272 (N_29272,N_26168,N_26813);
xor U29273 (N_29273,N_27183,N_27222);
or U29274 (N_29274,N_26543,N_27160);
nand U29275 (N_29275,N_27345,N_26583);
nor U29276 (N_29276,N_26068,N_27193);
nor U29277 (N_29277,N_26629,N_26475);
or U29278 (N_29278,N_27731,N_27365);
and U29279 (N_29279,N_26815,N_27978);
and U29280 (N_29280,N_27673,N_27711);
xor U29281 (N_29281,N_27728,N_27488);
nor U29282 (N_29282,N_26537,N_27477);
or U29283 (N_29283,N_27057,N_27033);
nand U29284 (N_29284,N_26368,N_26652);
nand U29285 (N_29285,N_27441,N_26110);
xor U29286 (N_29286,N_27270,N_27602);
and U29287 (N_29287,N_26151,N_27489);
xnor U29288 (N_29288,N_26416,N_26537);
and U29289 (N_29289,N_26341,N_26395);
and U29290 (N_29290,N_26757,N_27223);
xor U29291 (N_29291,N_27142,N_27177);
xor U29292 (N_29292,N_26715,N_27760);
and U29293 (N_29293,N_26430,N_27440);
nand U29294 (N_29294,N_26170,N_27172);
and U29295 (N_29295,N_27638,N_26856);
nand U29296 (N_29296,N_27461,N_27068);
nor U29297 (N_29297,N_27451,N_26013);
or U29298 (N_29298,N_27881,N_27270);
and U29299 (N_29299,N_26492,N_26173);
or U29300 (N_29300,N_26539,N_27088);
xor U29301 (N_29301,N_26751,N_26305);
nand U29302 (N_29302,N_26153,N_26962);
and U29303 (N_29303,N_26341,N_27542);
nor U29304 (N_29304,N_27184,N_27957);
and U29305 (N_29305,N_27657,N_26995);
and U29306 (N_29306,N_26141,N_26510);
nor U29307 (N_29307,N_26544,N_26306);
and U29308 (N_29308,N_26785,N_26730);
nand U29309 (N_29309,N_26875,N_26551);
nor U29310 (N_29310,N_27236,N_26900);
xor U29311 (N_29311,N_26940,N_27248);
xor U29312 (N_29312,N_26010,N_26019);
and U29313 (N_29313,N_27948,N_27875);
nor U29314 (N_29314,N_27445,N_26762);
nand U29315 (N_29315,N_27685,N_27366);
xor U29316 (N_29316,N_26429,N_26313);
xor U29317 (N_29317,N_26061,N_26973);
and U29318 (N_29318,N_27329,N_27040);
nand U29319 (N_29319,N_27438,N_26060);
xnor U29320 (N_29320,N_26216,N_26621);
xor U29321 (N_29321,N_27764,N_27040);
nor U29322 (N_29322,N_27470,N_27630);
nand U29323 (N_29323,N_26262,N_26991);
and U29324 (N_29324,N_27089,N_27723);
nand U29325 (N_29325,N_26899,N_27148);
xor U29326 (N_29326,N_27279,N_26966);
and U29327 (N_29327,N_26692,N_27608);
xnor U29328 (N_29328,N_26125,N_26585);
nand U29329 (N_29329,N_26697,N_27315);
xor U29330 (N_29330,N_26699,N_27913);
xor U29331 (N_29331,N_26914,N_26222);
or U29332 (N_29332,N_26414,N_27041);
nor U29333 (N_29333,N_26709,N_26522);
and U29334 (N_29334,N_27439,N_26728);
nand U29335 (N_29335,N_27121,N_26499);
and U29336 (N_29336,N_26049,N_26978);
nand U29337 (N_29337,N_27365,N_27667);
nand U29338 (N_29338,N_26651,N_26437);
nor U29339 (N_29339,N_27134,N_27928);
xnor U29340 (N_29340,N_27955,N_26830);
xnor U29341 (N_29341,N_27062,N_27367);
xnor U29342 (N_29342,N_27890,N_27542);
nand U29343 (N_29343,N_26058,N_27765);
xor U29344 (N_29344,N_27400,N_26599);
nor U29345 (N_29345,N_26384,N_27791);
xnor U29346 (N_29346,N_27177,N_26583);
and U29347 (N_29347,N_26380,N_27531);
nand U29348 (N_29348,N_27963,N_27332);
xor U29349 (N_29349,N_27394,N_27837);
or U29350 (N_29350,N_26975,N_27564);
xor U29351 (N_29351,N_26584,N_26957);
and U29352 (N_29352,N_26267,N_27732);
xor U29353 (N_29353,N_26099,N_26255);
nor U29354 (N_29354,N_27869,N_27609);
nand U29355 (N_29355,N_26317,N_27846);
and U29356 (N_29356,N_27193,N_27519);
nor U29357 (N_29357,N_26859,N_26909);
nor U29358 (N_29358,N_27776,N_27526);
or U29359 (N_29359,N_27978,N_27916);
xnor U29360 (N_29360,N_26465,N_26287);
nor U29361 (N_29361,N_27162,N_27677);
nor U29362 (N_29362,N_26513,N_27125);
xor U29363 (N_29363,N_27572,N_26092);
nand U29364 (N_29364,N_26282,N_27733);
nand U29365 (N_29365,N_26089,N_26021);
nor U29366 (N_29366,N_27602,N_26567);
and U29367 (N_29367,N_26420,N_27207);
nor U29368 (N_29368,N_27231,N_27887);
nand U29369 (N_29369,N_27994,N_26141);
nor U29370 (N_29370,N_26111,N_27750);
xnor U29371 (N_29371,N_27052,N_26530);
nand U29372 (N_29372,N_27470,N_27098);
and U29373 (N_29373,N_26838,N_27207);
xor U29374 (N_29374,N_27476,N_27443);
nor U29375 (N_29375,N_26613,N_27102);
xor U29376 (N_29376,N_27730,N_26223);
and U29377 (N_29377,N_27621,N_26971);
and U29378 (N_29378,N_27058,N_27820);
nor U29379 (N_29379,N_26574,N_27789);
and U29380 (N_29380,N_27020,N_27631);
nor U29381 (N_29381,N_26168,N_27083);
and U29382 (N_29382,N_27568,N_26474);
or U29383 (N_29383,N_27470,N_27109);
or U29384 (N_29384,N_26886,N_27278);
xor U29385 (N_29385,N_26208,N_27941);
and U29386 (N_29386,N_26020,N_26993);
xor U29387 (N_29387,N_27439,N_27969);
xor U29388 (N_29388,N_26068,N_26924);
and U29389 (N_29389,N_27405,N_27351);
nand U29390 (N_29390,N_26821,N_27069);
and U29391 (N_29391,N_26564,N_26277);
nand U29392 (N_29392,N_27348,N_26707);
xnor U29393 (N_29393,N_27398,N_26321);
nand U29394 (N_29394,N_26633,N_27846);
xor U29395 (N_29395,N_26445,N_27968);
and U29396 (N_29396,N_26848,N_27423);
xnor U29397 (N_29397,N_27090,N_26248);
nand U29398 (N_29398,N_26184,N_27192);
and U29399 (N_29399,N_27016,N_27887);
or U29400 (N_29400,N_26168,N_26628);
nor U29401 (N_29401,N_26970,N_27912);
xor U29402 (N_29402,N_27382,N_27653);
xor U29403 (N_29403,N_26399,N_26945);
xnor U29404 (N_29404,N_27985,N_27256);
nand U29405 (N_29405,N_26252,N_27701);
nand U29406 (N_29406,N_27291,N_26839);
and U29407 (N_29407,N_26676,N_26279);
or U29408 (N_29408,N_26702,N_27885);
xor U29409 (N_29409,N_27579,N_27793);
and U29410 (N_29410,N_26879,N_27032);
nand U29411 (N_29411,N_26150,N_26426);
nand U29412 (N_29412,N_26512,N_26998);
and U29413 (N_29413,N_27743,N_26611);
and U29414 (N_29414,N_27353,N_26124);
and U29415 (N_29415,N_26669,N_26962);
and U29416 (N_29416,N_27856,N_26057);
and U29417 (N_29417,N_26108,N_27583);
xor U29418 (N_29418,N_26150,N_26295);
and U29419 (N_29419,N_26546,N_27202);
xor U29420 (N_29420,N_26641,N_27023);
xnor U29421 (N_29421,N_27580,N_26516);
nand U29422 (N_29422,N_26695,N_26911);
nand U29423 (N_29423,N_27957,N_27515);
and U29424 (N_29424,N_27162,N_26178);
or U29425 (N_29425,N_26599,N_27682);
nand U29426 (N_29426,N_27231,N_27489);
and U29427 (N_29427,N_27145,N_27346);
nor U29428 (N_29428,N_26010,N_26314);
xnor U29429 (N_29429,N_26130,N_27128);
and U29430 (N_29430,N_26948,N_26150);
xnor U29431 (N_29431,N_27832,N_26048);
or U29432 (N_29432,N_26423,N_26642);
or U29433 (N_29433,N_26924,N_26201);
and U29434 (N_29434,N_27255,N_26294);
and U29435 (N_29435,N_26830,N_26984);
or U29436 (N_29436,N_26955,N_26765);
xor U29437 (N_29437,N_26058,N_26442);
xor U29438 (N_29438,N_26391,N_27680);
xnor U29439 (N_29439,N_26460,N_27149);
and U29440 (N_29440,N_27724,N_26428);
or U29441 (N_29441,N_26756,N_26324);
nor U29442 (N_29442,N_27169,N_26292);
nor U29443 (N_29443,N_27517,N_27709);
or U29444 (N_29444,N_27140,N_27002);
or U29445 (N_29445,N_26077,N_27288);
xor U29446 (N_29446,N_27968,N_27083);
and U29447 (N_29447,N_27559,N_27681);
xor U29448 (N_29448,N_27943,N_27500);
nand U29449 (N_29449,N_27399,N_26536);
or U29450 (N_29450,N_26387,N_26848);
or U29451 (N_29451,N_26904,N_26821);
xor U29452 (N_29452,N_26391,N_26367);
and U29453 (N_29453,N_27747,N_26532);
nand U29454 (N_29454,N_26640,N_27245);
nand U29455 (N_29455,N_27735,N_26738);
and U29456 (N_29456,N_27207,N_26293);
nand U29457 (N_29457,N_27509,N_26418);
nand U29458 (N_29458,N_27351,N_26264);
nand U29459 (N_29459,N_27878,N_27754);
nor U29460 (N_29460,N_27865,N_26154);
xor U29461 (N_29461,N_26600,N_26001);
nor U29462 (N_29462,N_26448,N_27911);
nand U29463 (N_29463,N_27420,N_27917);
or U29464 (N_29464,N_26551,N_26591);
nand U29465 (N_29465,N_26845,N_27581);
nor U29466 (N_29466,N_27139,N_26116);
and U29467 (N_29467,N_26013,N_27008);
and U29468 (N_29468,N_26945,N_26136);
nor U29469 (N_29469,N_26397,N_27149);
and U29470 (N_29470,N_26273,N_26377);
and U29471 (N_29471,N_26560,N_26031);
xnor U29472 (N_29472,N_27120,N_26570);
nand U29473 (N_29473,N_26652,N_27499);
or U29474 (N_29474,N_27924,N_27136);
nand U29475 (N_29475,N_27529,N_27754);
nand U29476 (N_29476,N_26147,N_26046);
nor U29477 (N_29477,N_27809,N_27842);
or U29478 (N_29478,N_27109,N_27995);
nor U29479 (N_29479,N_27609,N_26870);
nand U29480 (N_29480,N_26363,N_26122);
or U29481 (N_29481,N_27674,N_27057);
and U29482 (N_29482,N_26805,N_26157);
nand U29483 (N_29483,N_27925,N_27443);
nand U29484 (N_29484,N_26396,N_26690);
nor U29485 (N_29485,N_26626,N_26644);
xnor U29486 (N_29486,N_27202,N_27582);
xor U29487 (N_29487,N_26014,N_27184);
and U29488 (N_29488,N_27769,N_26828);
xor U29489 (N_29489,N_26719,N_26478);
nand U29490 (N_29490,N_27000,N_27781);
and U29491 (N_29491,N_27866,N_27209);
xor U29492 (N_29492,N_27467,N_26760);
xnor U29493 (N_29493,N_26174,N_26389);
nor U29494 (N_29494,N_27471,N_27550);
and U29495 (N_29495,N_27688,N_27663);
and U29496 (N_29496,N_27549,N_27681);
xnor U29497 (N_29497,N_27643,N_26180);
and U29498 (N_29498,N_27585,N_27526);
nor U29499 (N_29499,N_26752,N_26393);
or U29500 (N_29500,N_27510,N_26033);
or U29501 (N_29501,N_27432,N_27288);
xor U29502 (N_29502,N_27181,N_27154);
nor U29503 (N_29503,N_27074,N_26334);
nand U29504 (N_29504,N_26596,N_27071);
nand U29505 (N_29505,N_26236,N_27522);
or U29506 (N_29506,N_27761,N_27375);
nand U29507 (N_29507,N_26819,N_27747);
or U29508 (N_29508,N_27924,N_26384);
and U29509 (N_29509,N_27893,N_27629);
and U29510 (N_29510,N_27796,N_26086);
and U29511 (N_29511,N_26549,N_26957);
and U29512 (N_29512,N_26372,N_27861);
nand U29513 (N_29513,N_27553,N_27239);
and U29514 (N_29514,N_27684,N_27814);
and U29515 (N_29515,N_26542,N_26271);
or U29516 (N_29516,N_27656,N_27367);
xor U29517 (N_29517,N_26665,N_27808);
nand U29518 (N_29518,N_26210,N_27470);
or U29519 (N_29519,N_27637,N_26026);
nor U29520 (N_29520,N_26228,N_26636);
nor U29521 (N_29521,N_26221,N_26126);
nor U29522 (N_29522,N_27814,N_26252);
or U29523 (N_29523,N_26452,N_27812);
or U29524 (N_29524,N_27832,N_27363);
xor U29525 (N_29525,N_27437,N_27478);
xor U29526 (N_29526,N_26059,N_26142);
xor U29527 (N_29527,N_27000,N_26774);
or U29528 (N_29528,N_27698,N_27043);
and U29529 (N_29529,N_27986,N_27803);
or U29530 (N_29530,N_27595,N_27243);
xor U29531 (N_29531,N_26611,N_27330);
nor U29532 (N_29532,N_27575,N_26584);
or U29533 (N_29533,N_26675,N_27232);
or U29534 (N_29534,N_27780,N_26097);
nand U29535 (N_29535,N_27615,N_27045);
nor U29536 (N_29536,N_27252,N_27581);
nor U29537 (N_29537,N_27986,N_27387);
or U29538 (N_29538,N_27898,N_26431);
nand U29539 (N_29539,N_27377,N_26756);
or U29540 (N_29540,N_26161,N_27393);
nor U29541 (N_29541,N_27063,N_27818);
nor U29542 (N_29542,N_26775,N_27239);
and U29543 (N_29543,N_26420,N_26648);
and U29544 (N_29544,N_26964,N_27152);
nand U29545 (N_29545,N_26948,N_26740);
nor U29546 (N_29546,N_26812,N_27637);
or U29547 (N_29547,N_27929,N_27580);
nor U29548 (N_29548,N_27322,N_26679);
or U29549 (N_29549,N_26168,N_27295);
nor U29550 (N_29550,N_26264,N_27203);
or U29551 (N_29551,N_26084,N_26301);
xor U29552 (N_29552,N_27923,N_26888);
nor U29553 (N_29553,N_27368,N_26911);
nor U29554 (N_29554,N_26794,N_27457);
or U29555 (N_29555,N_27071,N_27281);
or U29556 (N_29556,N_27997,N_27766);
nor U29557 (N_29557,N_26397,N_27005);
nor U29558 (N_29558,N_27177,N_26670);
and U29559 (N_29559,N_26277,N_26869);
nor U29560 (N_29560,N_26603,N_26974);
xor U29561 (N_29561,N_27871,N_27340);
and U29562 (N_29562,N_27563,N_26870);
nor U29563 (N_29563,N_26504,N_27208);
xnor U29564 (N_29564,N_26851,N_27632);
or U29565 (N_29565,N_27189,N_26926);
nor U29566 (N_29566,N_27869,N_26421);
nand U29567 (N_29567,N_26625,N_26653);
or U29568 (N_29568,N_27642,N_26122);
and U29569 (N_29569,N_26375,N_26712);
and U29570 (N_29570,N_26516,N_27929);
xor U29571 (N_29571,N_27856,N_26076);
xor U29572 (N_29572,N_26281,N_26705);
or U29573 (N_29573,N_26506,N_26598);
and U29574 (N_29574,N_26434,N_26827);
xor U29575 (N_29575,N_26602,N_27337);
xor U29576 (N_29576,N_26355,N_26053);
or U29577 (N_29577,N_26214,N_27733);
nand U29578 (N_29578,N_27345,N_27492);
xor U29579 (N_29579,N_27921,N_27060);
nand U29580 (N_29580,N_27922,N_26862);
or U29581 (N_29581,N_26470,N_26678);
or U29582 (N_29582,N_26035,N_27541);
nor U29583 (N_29583,N_26553,N_27687);
nor U29584 (N_29584,N_27041,N_27375);
or U29585 (N_29585,N_27540,N_26749);
nor U29586 (N_29586,N_26915,N_27061);
nor U29587 (N_29587,N_26159,N_26712);
xor U29588 (N_29588,N_26372,N_26441);
nor U29589 (N_29589,N_26930,N_26524);
or U29590 (N_29590,N_26860,N_27245);
or U29591 (N_29591,N_27547,N_27292);
or U29592 (N_29592,N_27716,N_27790);
nand U29593 (N_29593,N_26731,N_27375);
nor U29594 (N_29594,N_26876,N_26838);
xor U29595 (N_29595,N_26593,N_26017);
and U29596 (N_29596,N_26366,N_26471);
xor U29597 (N_29597,N_27029,N_26308);
and U29598 (N_29598,N_27475,N_26573);
nand U29599 (N_29599,N_27272,N_26552);
or U29600 (N_29600,N_27762,N_27040);
xnor U29601 (N_29601,N_26845,N_27558);
nand U29602 (N_29602,N_26460,N_26707);
and U29603 (N_29603,N_27822,N_27819);
xor U29604 (N_29604,N_27763,N_27449);
nor U29605 (N_29605,N_26232,N_26053);
and U29606 (N_29606,N_26820,N_27285);
or U29607 (N_29607,N_27125,N_26302);
or U29608 (N_29608,N_26957,N_27651);
nand U29609 (N_29609,N_26349,N_26379);
nand U29610 (N_29610,N_26881,N_27315);
or U29611 (N_29611,N_26333,N_26203);
xor U29612 (N_29612,N_27508,N_27285);
xnor U29613 (N_29613,N_26510,N_27273);
nand U29614 (N_29614,N_26136,N_27554);
xor U29615 (N_29615,N_26757,N_26540);
xnor U29616 (N_29616,N_27904,N_26700);
or U29617 (N_29617,N_26881,N_26705);
or U29618 (N_29618,N_26167,N_27954);
xnor U29619 (N_29619,N_26126,N_27975);
xor U29620 (N_29620,N_27243,N_26530);
and U29621 (N_29621,N_27536,N_27560);
and U29622 (N_29622,N_26337,N_26578);
xor U29623 (N_29623,N_27348,N_27180);
xnor U29624 (N_29624,N_26327,N_26822);
nand U29625 (N_29625,N_27226,N_27649);
nand U29626 (N_29626,N_26075,N_26940);
nand U29627 (N_29627,N_26495,N_26086);
nand U29628 (N_29628,N_27816,N_26670);
or U29629 (N_29629,N_26939,N_26832);
nor U29630 (N_29630,N_27387,N_27910);
or U29631 (N_29631,N_27252,N_27186);
nor U29632 (N_29632,N_27362,N_27208);
nand U29633 (N_29633,N_26109,N_26177);
xnor U29634 (N_29634,N_26087,N_26062);
or U29635 (N_29635,N_27580,N_26518);
or U29636 (N_29636,N_27361,N_26902);
nand U29637 (N_29637,N_27005,N_26249);
and U29638 (N_29638,N_26987,N_27826);
nor U29639 (N_29639,N_27090,N_27567);
and U29640 (N_29640,N_27954,N_27723);
nor U29641 (N_29641,N_27480,N_26092);
nor U29642 (N_29642,N_27445,N_27474);
xnor U29643 (N_29643,N_26545,N_27120);
nor U29644 (N_29644,N_27783,N_27315);
nor U29645 (N_29645,N_27102,N_27760);
or U29646 (N_29646,N_27697,N_27632);
nand U29647 (N_29647,N_26632,N_27720);
nand U29648 (N_29648,N_26827,N_27763);
xnor U29649 (N_29649,N_26858,N_27283);
nor U29650 (N_29650,N_27473,N_27862);
and U29651 (N_29651,N_27567,N_27132);
nand U29652 (N_29652,N_26061,N_27826);
and U29653 (N_29653,N_26884,N_26069);
nand U29654 (N_29654,N_27047,N_27743);
and U29655 (N_29655,N_27267,N_27793);
and U29656 (N_29656,N_27533,N_27467);
nand U29657 (N_29657,N_26995,N_27797);
nor U29658 (N_29658,N_27993,N_27086);
nor U29659 (N_29659,N_26941,N_26021);
nand U29660 (N_29660,N_26023,N_26918);
or U29661 (N_29661,N_26093,N_26432);
xor U29662 (N_29662,N_26512,N_26500);
nand U29663 (N_29663,N_26264,N_26686);
or U29664 (N_29664,N_26379,N_27233);
or U29665 (N_29665,N_27119,N_27866);
nand U29666 (N_29666,N_26582,N_26829);
nand U29667 (N_29667,N_27108,N_26510);
or U29668 (N_29668,N_26887,N_26505);
nor U29669 (N_29669,N_26989,N_27633);
and U29670 (N_29670,N_27597,N_26155);
xnor U29671 (N_29671,N_26480,N_26365);
nand U29672 (N_29672,N_27674,N_26811);
nor U29673 (N_29673,N_26004,N_26312);
nand U29674 (N_29674,N_27198,N_26509);
nor U29675 (N_29675,N_27203,N_27096);
and U29676 (N_29676,N_27624,N_27958);
nor U29677 (N_29677,N_27532,N_27554);
nor U29678 (N_29678,N_27176,N_27981);
and U29679 (N_29679,N_27545,N_27169);
xnor U29680 (N_29680,N_26650,N_27498);
and U29681 (N_29681,N_27352,N_26519);
or U29682 (N_29682,N_26368,N_26842);
nand U29683 (N_29683,N_27721,N_27604);
xor U29684 (N_29684,N_26706,N_27500);
xor U29685 (N_29685,N_26344,N_27445);
nor U29686 (N_29686,N_27895,N_27839);
or U29687 (N_29687,N_27763,N_27116);
or U29688 (N_29688,N_26062,N_26976);
nand U29689 (N_29689,N_26390,N_27628);
and U29690 (N_29690,N_27432,N_26989);
or U29691 (N_29691,N_27856,N_27817);
nor U29692 (N_29692,N_27982,N_27548);
xnor U29693 (N_29693,N_27791,N_27197);
and U29694 (N_29694,N_27071,N_27064);
xnor U29695 (N_29695,N_26460,N_27068);
nor U29696 (N_29696,N_27628,N_26190);
nand U29697 (N_29697,N_27183,N_26321);
and U29698 (N_29698,N_27958,N_26942);
and U29699 (N_29699,N_27024,N_26395);
nand U29700 (N_29700,N_26240,N_27415);
or U29701 (N_29701,N_26086,N_27670);
or U29702 (N_29702,N_27425,N_27064);
nor U29703 (N_29703,N_27325,N_26136);
nor U29704 (N_29704,N_27012,N_26303);
or U29705 (N_29705,N_27117,N_27923);
nor U29706 (N_29706,N_26594,N_27125);
or U29707 (N_29707,N_27349,N_26032);
or U29708 (N_29708,N_26606,N_26499);
nor U29709 (N_29709,N_27506,N_27457);
and U29710 (N_29710,N_26780,N_26490);
xor U29711 (N_29711,N_27380,N_26890);
and U29712 (N_29712,N_27886,N_26060);
or U29713 (N_29713,N_27307,N_27709);
xnor U29714 (N_29714,N_26081,N_26502);
nor U29715 (N_29715,N_27121,N_27554);
nand U29716 (N_29716,N_27813,N_27054);
and U29717 (N_29717,N_27565,N_27621);
xnor U29718 (N_29718,N_27971,N_27475);
xor U29719 (N_29719,N_27523,N_26906);
xor U29720 (N_29720,N_26161,N_26277);
nand U29721 (N_29721,N_27020,N_27457);
nor U29722 (N_29722,N_26813,N_26068);
or U29723 (N_29723,N_26605,N_27123);
or U29724 (N_29724,N_26984,N_26539);
nor U29725 (N_29725,N_27048,N_27709);
nor U29726 (N_29726,N_26634,N_26260);
nor U29727 (N_29727,N_26063,N_26342);
xnor U29728 (N_29728,N_26911,N_26968);
nand U29729 (N_29729,N_26624,N_27372);
nor U29730 (N_29730,N_26084,N_26281);
xnor U29731 (N_29731,N_26913,N_26242);
nand U29732 (N_29732,N_26425,N_26495);
nand U29733 (N_29733,N_26804,N_27949);
or U29734 (N_29734,N_27422,N_26087);
and U29735 (N_29735,N_27630,N_27189);
nand U29736 (N_29736,N_26335,N_27886);
nor U29737 (N_29737,N_26449,N_26692);
xor U29738 (N_29738,N_26675,N_27987);
and U29739 (N_29739,N_27792,N_27320);
and U29740 (N_29740,N_26031,N_27807);
or U29741 (N_29741,N_27554,N_27119);
xor U29742 (N_29742,N_26702,N_26021);
nor U29743 (N_29743,N_26851,N_26648);
and U29744 (N_29744,N_27320,N_26451);
xnor U29745 (N_29745,N_27869,N_27267);
or U29746 (N_29746,N_27431,N_27609);
and U29747 (N_29747,N_27656,N_26411);
or U29748 (N_29748,N_26248,N_27356);
nor U29749 (N_29749,N_26452,N_27336);
nor U29750 (N_29750,N_26596,N_26628);
nand U29751 (N_29751,N_26124,N_27278);
or U29752 (N_29752,N_27988,N_27775);
and U29753 (N_29753,N_27472,N_27669);
nor U29754 (N_29754,N_26174,N_27394);
xor U29755 (N_29755,N_26817,N_27645);
or U29756 (N_29756,N_26676,N_26261);
xor U29757 (N_29757,N_27755,N_26372);
and U29758 (N_29758,N_26251,N_26972);
nand U29759 (N_29759,N_26529,N_26948);
or U29760 (N_29760,N_26032,N_26777);
xor U29761 (N_29761,N_26998,N_26927);
or U29762 (N_29762,N_26444,N_26555);
or U29763 (N_29763,N_26776,N_27561);
nor U29764 (N_29764,N_26817,N_26172);
and U29765 (N_29765,N_27291,N_27081);
nor U29766 (N_29766,N_27434,N_26149);
or U29767 (N_29767,N_27626,N_26817);
nor U29768 (N_29768,N_27899,N_27129);
xnor U29769 (N_29769,N_26879,N_26303);
nand U29770 (N_29770,N_26587,N_26166);
and U29771 (N_29771,N_26053,N_27068);
or U29772 (N_29772,N_27405,N_26444);
nand U29773 (N_29773,N_26502,N_27580);
xor U29774 (N_29774,N_27583,N_26225);
nor U29775 (N_29775,N_27523,N_27814);
nor U29776 (N_29776,N_26365,N_26360);
or U29777 (N_29777,N_27994,N_26958);
or U29778 (N_29778,N_27189,N_26431);
and U29779 (N_29779,N_27420,N_27749);
xor U29780 (N_29780,N_27609,N_26136);
or U29781 (N_29781,N_26872,N_26667);
and U29782 (N_29782,N_27495,N_27066);
nand U29783 (N_29783,N_27391,N_26315);
nor U29784 (N_29784,N_26375,N_27839);
nor U29785 (N_29785,N_27605,N_26524);
nor U29786 (N_29786,N_26074,N_27935);
nand U29787 (N_29787,N_26094,N_26176);
nor U29788 (N_29788,N_27218,N_26803);
nand U29789 (N_29789,N_27410,N_26961);
nand U29790 (N_29790,N_26590,N_27133);
nor U29791 (N_29791,N_27480,N_27672);
xnor U29792 (N_29792,N_27840,N_26754);
and U29793 (N_29793,N_27238,N_26359);
xor U29794 (N_29794,N_27727,N_26910);
and U29795 (N_29795,N_27093,N_26029);
xor U29796 (N_29796,N_26166,N_26726);
nor U29797 (N_29797,N_26296,N_27206);
nand U29798 (N_29798,N_26002,N_27373);
xor U29799 (N_29799,N_27871,N_27766);
nor U29800 (N_29800,N_27233,N_26899);
or U29801 (N_29801,N_26394,N_27678);
nor U29802 (N_29802,N_26888,N_26807);
and U29803 (N_29803,N_27528,N_26452);
or U29804 (N_29804,N_27743,N_27277);
xor U29805 (N_29805,N_26763,N_27457);
nor U29806 (N_29806,N_27924,N_27104);
or U29807 (N_29807,N_27940,N_26336);
or U29808 (N_29808,N_27328,N_27459);
xor U29809 (N_29809,N_27485,N_26500);
xor U29810 (N_29810,N_26383,N_27612);
nor U29811 (N_29811,N_26705,N_26834);
xnor U29812 (N_29812,N_27223,N_27739);
and U29813 (N_29813,N_27326,N_27527);
or U29814 (N_29814,N_27184,N_26454);
nor U29815 (N_29815,N_26157,N_27038);
and U29816 (N_29816,N_27662,N_27826);
nand U29817 (N_29817,N_26493,N_27653);
nor U29818 (N_29818,N_27936,N_26089);
nor U29819 (N_29819,N_26420,N_26294);
nor U29820 (N_29820,N_26906,N_27752);
and U29821 (N_29821,N_26596,N_26521);
nor U29822 (N_29822,N_26450,N_26064);
xor U29823 (N_29823,N_27093,N_27383);
or U29824 (N_29824,N_26732,N_27563);
nor U29825 (N_29825,N_26563,N_26899);
xor U29826 (N_29826,N_26738,N_26610);
or U29827 (N_29827,N_26163,N_27459);
nor U29828 (N_29828,N_27897,N_26620);
and U29829 (N_29829,N_26745,N_26667);
and U29830 (N_29830,N_27143,N_27492);
or U29831 (N_29831,N_26343,N_26035);
nor U29832 (N_29832,N_27209,N_26402);
nand U29833 (N_29833,N_26795,N_27423);
xor U29834 (N_29834,N_26073,N_26811);
xnor U29835 (N_29835,N_27072,N_27762);
nor U29836 (N_29836,N_26849,N_27584);
nor U29837 (N_29837,N_27280,N_27552);
and U29838 (N_29838,N_26345,N_27917);
or U29839 (N_29839,N_26752,N_26130);
or U29840 (N_29840,N_27519,N_27606);
or U29841 (N_29841,N_26441,N_27851);
xnor U29842 (N_29842,N_27034,N_27047);
nand U29843 (N_29843,N_27863,N_27095);
nand U29844 (N_29844,N_27680,N_26578);
xor U29845 (N_29845,N_27595,N_27529);
and U29846 (N_29846,N_27672,N_27046);
nand U29847 (N_29847,N_27140,N_27192);
nor U29848 (N_29848,N_26004,N_26318);
or U29849 (N_29849,N_26147,N_27222);
nor U29850 (N_29850,N_27315,N_27063);
nand U29851 (N_29851,N_27828,N_26494);
or U29852 (N_29852,N_27019,N_26008);
nand U29853 (N_29853,N_26281,N_27522);
xor U29854 (N_29854,N_26399,N_27495);
nor U29855 (N_29855,N_27447,N_27880);
xor U29856 (N_29856,N_26304,N_26314);
and U29857 (N_29857,N_27272,N_26452);
and U29858 (N_29858,N_27765,N_27381);
or U29859 (N_29859,N_26884,N_26940);
nor U29860 (N_29860,N_27189,N_26839);
or U29861 (N_29861,N_26960,N_27770);
or U29862 (N_29862,N_27248,N_27290);
xor U29863 (N_29863,N_27655,N_27980);
and U29864 (N_29864,N_27660,N_26308);
and U29865 (N_29865,N_27404,N_27069);
nor U29866 (N_29866,N_27589,N_27754);
nand U29867 (N_29867,N_26720,N_27575);
or U29868 (N_29868,N_26840,N_26586);
xnor U29869 (N_29869,N_26244,N_26117);
nor U29870 (N_29870,N_26800,N_27849);
nor U29871 (N_29871,N_27868,N_26095);
and U29872 (N_29872,N_27650,N_27761);
nor U29873 (N_29873,N_26592,N_27070);
and U29874 (N_29874,N_26291,N_27159);
or U29875 (N_29875,N_27602,N_26547);
nor U29876 (N_29876,N_26073,N_26401);
nor U29877 (N_29877,N_27204,N_27393);
and U29878 (N_29878,N_27897,N_26412);
or U29879 (N_29879,N_27288,N_27261);
xor U29880 (N_29880,N_27730,N_26216);
nand U29881 (N_29881,N_27274,N_26067);
nor U29882 (N_29882,N_27336,N_26441);
nand U29883 (N_29883,N_27332,N_27300);
nor U29884 (N_29884,N_26578,N_27929);
xnor U29885 (N_29885,N_26061,N_26432);
nand U29886 (N_29886,N_27870,N_26855);
nor U29887 (N_29887,N_27561,N_26224);
nor U29888 (N_29888,N_26751,N_27905);
and U29889 (N_29889,N_27548,N_27501);
xnor U29890 (N_29890,N_27377,N_26099);
xor U29891 (N_29891,N_27170,N_27525);
or U29892 (N_29892,N_27499,N_26452);
nor U29893 (N_29893,N_27510,N_27771);
or U29894 (N_29894,N_27987,N_27789);
nand U29895 (N_29895,N_26755,N_26458);
and U29896 (N_29896,N_27675,N_27324);
and U29897 (N_29897,N_26650,N_27700);
and U29898 (N_29898,N_26611,N_27348);
or U29899 (N_29899,N_27521,N_26214);
and U29900 (N_29900,N_26490,N_26754);
nor U29901 (N_29901,N_27433,N_27494);
and U29902 (N_29902,N_26543,N_27248);
nand U29903 (N_29903,N_27030,N_27323);
xor U29904 (N_29904,N_27443,N_26833);
xnor U29905 (N_29905,N_27593,N_26262);
and U29906 (N_29906,N_26476,N_26071);
and U29907 (N_29907,N_26721,N_26589);
and U29908 (N_29908,N_27434,N_26571);
nor U29909 (N_29909,N_26310,N_27032);
nor U29910 (N_29910,N_27552,N_26100);
xor U29911 (N_29911,N_27095,N_27372);
xnor U29912 (N_29912,N_26518,N_27646);
or U29913 (N_29913,N_27314,N_26764);
xnor U29914 (N_29914,N_27597,N_26759);
or U29915 (N_29915,N_26481,N_26762);
nor U29916 (N_29916,N_26467,N_27654);
and U29917 (N_29917,N_26128,N_27789);
xor U29918 (N_29918,N_27811,N_27011);
nor U29919 (N_29919,N_26357,N_26083);
or U29920 (N_29920,N_27090,N_27946);
nor U29921 (N_29921,N_26352,N_27758);
nor U29922 (N_29922,N_27994,N_26819);
xor U29923 (N_29923,N_27003,N_26245);
or U29924 (N_29924,N_26985,N_27283);
nand U29925 (N_29925,N_26043,N_26022);
nor U29926 (N_29926,N_26444,N_27406);
nor U29927 (N_29927,N_27487,N_27272);
and U29928 (N_29928,N_27130,N_27203);
or U29929 (N_29929,N_26676,N_27678);
nand U29930 (N_29930,N_26062,N_27822);
or U29931 (N_29931,N_27797,N_27389);
or U29932 (N_29932,N_27057,N_26558);
nor U29933 (N_29933,N_26770,N_26089);
and U29934 (N_29934,N_27057,N_26561);
xor U29935 (N_29935,N_26637,N_26877);
nor U29936 (N_29936,N_26725,N_26042);
nor U29937 (N_29937,N_26331,N_26649);
and U29938 (N_29938,N_26025,N_26399);
nor U29939 (N_29939,N_27839,N_27563);
nor U29940 (N_29940,N_26143,N_27398);
nand U29941 (N_29941,N_27070,N_26467);
and U29942 (N_29942,N_26987,N_27739);
nor U29943 (N_29943,N_26839,N_26254);
xnor U29944 (N_29944,N_27732,N_27675);
and U29945 (N_29945,N_27247,N_27416);
or U29946 (N_29946,N_27017,N_27876);
and U29947 (N_29947,N_26724,N_27825);
or U29948 (N_29948,N_27488,N_26564);
xnor U29949 (N_29949,N_27909,N_26258);
and U29950 (N_29950,N_26719,N_27839);
or U29951 (N_29951,N_26918,N_26117);
nor U29952 (N_29952,N_27844,N_27681);
and U29953 (N_29953,N_27819,N_26910);
xnor U29954 (N_29954,N_26792,N_26586);
or U29955 (N_29955,N_26602,N_27039);
and U29956 (N_29956,N_26677,N_27770);
or U29957 (N_29957,N_27243,N_27540);
xor U29958 (N_29958,N_27155,N_27225);
and U29959 (N_29959,N_26786,N_27445);
xor U29960 (N_29960,N_27817,N_27171);
nand U29961 (N_29961,N_26721,N_27888);
or U29962 (N_29962,N_26602,N_26620);
nor U29963 (N_29963,N_27671,N_27574);
and U29964 (N_29964,N_27724,N_27136);
xnor U29965 (N_29965,N_27856,N_26240);
nand U29966 (N_29966,N_27746,N_27402);
xnor U29967 (N_29967,N_27046,N_27379);
nand U29968 (N_29968,N_27134,N_27198);
and U29969 (N_29969,N_27024,N_26516);
and U29970 (N_29970,N_26225,N_27120);
nand U29971 (N_29971,N_26863,N_26258);
or U29972 (N_29972,N_26832,N_27348);
nand U29973 (N_29973,N_26148,N_27089);
or U29974 (N_29974,N_27468,N_26593);
nand U29975 (N_29975,N_27731,N_26394);
nor U29976 (N_29976,N_27588,N_26127);
xor U29977 (N_29977,N_27859,N_26193);
or U29978 (N_29978,N_26611,N_26672);
xnor U29979 (N_29979,N_27107,N_27489);
nor U29980 (N_29980,N_27961,N_26401);
and U29981 (N_29981,N_26785,N_27489);
nor U29982 (N_29982,N_26670,N_26342);
or U29983 (N_29983,N_27307,N_27037);
nor U29984 (N_29984,N_26966,N_27759);
and U29985 (N_29985,N_27737,N_27419);
nor U29986 (N_29986,N_27776,N_26991);
nand U29987 (N_29987,N_26562,N_26567);
xor U29988 (N_29988,N_27722,N_27467);
nor U29989 (N_29989,N_26854,N_27901);
or U29990 (N_29990,N_26488,N_27093);
nand U29991 (N_29991,N_27365,N_26367);
nand U29992 (N_29992,N_27673,N_26320);
and U29993 (N_29993,N_27087,N_26160);
nor U29994 (N_29994,N_27261,N_27289);
xnor U29995 (N_29995,N_27108,N_26245);
or U29996 (N_29996,N_27629,N_26064);
nor U29997 (N_29997,N_26823,N_26340);
xnor U29998 (N_29998,N_26272,N_26497);
xnor U29999 (N_29999,N_26419,N_27219);
or UO_0 (O_0,N_29419,N_29674);
and UO_1 (O_1,N_29980,N_28452);
or UO_2 (O_2,N_29220,N_29261);
nand UO_3 (O_3,N_29246,N_28400);
or UO_4 (O_4,N_28633,N_28193);
or UO_5 (O_5,N_28459,N_29649);
nand UO_6 (O_6,N_28592,N_28133);
and UO_7 (O_7,N_29213,N_28440);
and UO_8 (O_8,N_29087,N_29662);
and UO_9 (O_9,N_29678,N_29596);
and UO_10 (O_10,N_29279,N_29411);
nand UO_11 (O_11,N_28090,N_28650);
nor UO_12 (O_12,N_29519,N_29946);
nand UO_13 (O_13,N_29441,N_29570);
and UO_14 (O_14,N_29354,N_28364);
xnor UO_15 (O_15,N_28281,N_28265);
xor UO_16 (O_16,N_28727,N_29810);
or UO_17 (O_17,N_28998,N_28867);
and UO_18 (O_18,N_29917,N_28016);
and UO_19 (O_19,N_29774,N_28647);
nand UO_20 (O_20,N_29539,N_28557);
xor UO_21 (O_21,N_28912,N_29637);
and UO_22 (O_22,N_29081,N_28349);
nor UO_23 (O_23,N_28218,N_28235);
or UO_24 (O_24,N_28325,N_28717);
nor UO_25 (O_25,N_29203,N_29532);
nor UO_26 (O_26,N_28162,N_29648);
nand UO_27 (O_27,N_29921,N_28961);
nand UO_28 (O_28,N_28329,N_28463);
nor UO_29 (O_29,N_28051,N_28374);
and UO_30 (O_30,N_29823,N_28763);
nand UO_31 (O_31,N_29288,N_28978);
or UO_32 (O_32,N_29859,N_28445);
xnor UO_33 (O_33,N_29128,N_28285);
and UO_34 (O_34,N_29426,N_28471);
nor UO_35 (O_35,N_29525,N_28523);
nor UO_36 (O_36,N_28357,N_28490);
xor UO_37 (O_37,N_29912,N_28426);
or UO_38 (O_38,N_29661,N_28952);
nor UO_39 (O_39,N_28262,N_28887);
xor UO_40 (O_40,N_28561,N_28497);
nand UO_41 (O_41,N_28122,N_28156);
nor UO_42 (O_42,N_28749,N_29072);
or UO_43 (O_43,N_29676,N_28052);
and UO_44 (O_44,N_28888,N_29737);
nand UO_45 (O_45,N_28754,N_29030);
or UO_46 (O_46,N_28744,N_28663);
and UO_47 (O_47,N_28014,N_29188);
or UO_48 (O_48,N_28782,N_28702);
and UO_49 (O_49,N_28322,N_28819);
or UO_50 (O_50,N_29391,N_28326);
nor UO_51 (O_51,N_29351,N_28707);
or UO_52 (O_52,N_28226,N_28672);
nor UO_53 (O_53,N_29037,N_29146);
and UO_54 (O_54,N_28829,N_29167);
or UO_55 (O_55,N_28365,N_28907);
and UO_56 (O_56,N_28033,N_28280);
nand UO_57 (O_57,N_28099,N_29704);
and UO_58 (O_58,N_29699,N_29097);
and UO_59 (O_59,N_28498,N_28905);
or UO_60 (O_60,N_28775,N_28345);
nor UO_61 (O_61,N_29984,N_29263);
or UO_62 (O_62,N_29058,N_29165);
xnor UO_63 (O_63,N_28092,N_28873);
xor UO_64 (O_64,N_29130,N_29339);
xnor UO_65 (O_65,N_29773,N_28758);
nand UO_66 (O_66,N_29355,N_29155);
nand UO_67 (O_67,N_28529,N_28288);
nor UO_68 (O_68,N_28547,N_28394);
xnor UO_69 (O_69,N_29452,N_29932);
and UO_70 (O_70,N_28435,N_28298);
nand UO_71 (O_71,N_28869,N_28958);
or UO_72 (O_72,N_29680,N_28692);
nand UO_73 (O_73,N_29707,N_29235);
xnor UO_74 (O_74,N_28768,N_28662);
nor UO_75 (O_75,N_28332,N_28060);
nor UO_76 (O_76,N_28116,N_29065);
or UO_77 (O_77,N_29159,N_29301);
or UO_78 (O_78,N_28512,N_29237);
or UO_79 (O_79,N_29991,N_28624);
xnor UO_80 (O_80,N_28865,N_29114);
or UO_81 (O_81,N_29295,N_29333);
xor UO_82 (O_82,N_28733,N_28104);
nand UO_83 (O_83,N_29177,N_28622);
nor UO_84 (O_84,N_28198,N_28344);
and UO_85 (O_85,N_28831,N_29803);
xor UO_86 (O_86,N_28446,N_29077);
nor UO_87 (O_87,N_29118,N_28355);
nor UO_88 (O_88,N_28901,N_28395);
or UO_89 (O_89,N_28974,N_29726);
nand UO_90 (O_90,N_29489,N_29546);
xor UO_91 (O_91,N_29881,N_28712);
or UO_92 (O_92,N_28227,N_28406);
and UO_93 (O_93,N_29761,N_28679);
nor UO_94 (O_94,N_28335,N_28489);
or UO_95 (O_95,N_28925,N_28111);
nor UO_96 (O_96,N_29895,N_28913);
or UO_97 (O_97,N_29698,N_29011);
or UO_98 (O_98,N_29369,N_29222);
or UO_99 (O_99,N_28738,N_28272);
nand UO_100 (O_100,N_28508,N_28922);
nand UO_101 (O_101,N_29510,N_29560);
nand UO_102 (O_102,N_29093,N_28472);
nor UO_103 (O_103,N_29013,N_29822);
and UO_104 (O_104,N_28214,N_28625);
and UO_105 (O_105,N_29292,N_29606);
nor UO_106 (O_106,N_29896,N_29384);
nand UO_107 (O_107,N_28160,N_29799);
nor UO_108 (O_108,N_28765,N_29334);
or UO_109 (O_109,N_29053,N_29112);
xnor UO_110 (O_110,N_29040,N_28276);
xor UO_111 (O_111,N_28396,N_28384);
or UO_112 (O_112,N_28821,N_29347);
or UO_113 (O_113,N_29873,N_29732);
xor UO_114 (O_114,N_28460,N_28296);
nand UO_115 (O_115,N_28771,N_29216);
or UO_116 (O_116,N_28073,N_29504);
or UO_117 (O_117,N_29583,N_29179);
and UO_118 (O_118,N_28341,N_29756);
nor UO_119 (O_119,N_29660,N_29602);
and UO_120 (O_120,N_28610,N_29863);
or UO_121 (O_121,N_29325,N_28499);
and UO_122 (O_122,N_28630,N_29587);
nand UO_123 (O_123,N_29476,N_28682);
nor UO_124 (O_124,N_28404,N_29794);
xor UO_125 (O_125,N_28811,N_29378);
or UO_126 (O_126,N_29577,N_29158);
xor UO_127 (O_127,N_29718,N_29434);
or UO_128 (O_128,N_28177,N_28436);
xnor UO_129 (O_129,N_29524,N_29124);
nand UO_130 (O_130,N_28244,N_28613);
and UO_131 (O_131,N_29722,N_29401);
and UO_132 (O_132,N_28718,N_29493);
or UO_133 (O_133,N_29436,N_29084);
nor UO_134 (O_134,N_28693,N_28209);
nor UO_135 (O_135,N_29062,N_29802);
xnor UO_136 (O_136,N_28334,N_28586);
and UO_137 (O_137,N_28796,N_29017);
and UO_138 (O_138,N_29588,N_29439);
nand UO_139 (O_139,N_29728,N_29578);
nand UO_140 (O_140,N_28963,N_28784);
or UO_141 (O_141,N_29049,N_29902);
xnor UO_142 (O_142,N_29162,N_28238);
or UO_143 (O_143,N_29184,N_28317);
or UO_144 (O_144,N_28185,N_28081);
nand UO_145 (O_145,N_29137,N_29571);
nor UO_146 (O_146,N_29372,N_29095);
and UO_147 (O_147,N_28040,N_28543);
nor UO_148 (O_148,N_29956,N_28323);
nor UO_149 (O_149,N_28591,N_28654);
nor UO_150 (O_150,N_28079,N_29536);
nor UO_151 (O_151,N_28217,N_29685);
nor UO_152 (O_152,N_28751,N_29296);
and UO_153 (O_153,N_29066,N_28059);
nand UO_154 (O_154,N_28492,N_29815);
nand UO_155 (O_155,N_28466,N_29079);
nor UO_156 (O_156,N_28239,N_28785);
nor UO_157 (O_157,N_29782,N_28739);
nor UO_158 (O_158,N_28391,N_28229);
nor UO_159 (O_159,N_28858,N_29553);
and UO_160 (O_160,N_28421,N_28130);
and UO_161 (O_161,N_29952,N_29336);
xor UO_162 (O_162,N_29168,N_28070);
nor UO_163 (O_163,N_29703,N_28856);
nor UO_164 (O_164,N_28150,N_28791);
nand UO_165 (O_165,N_29321,N_28246);
and UO_166 (O_166,N_29034,N_28947);
nor UO_167 (O_167,N_28476,N_28207);
or UO_168 (O_168,N_28169,N_28000);
and UO_169 (O_169,N_28319,N_29819);
or UO_170 (O_170,N_29437,N_29923);
nand UO_171 (O_171,N_29410,N_29242);
nand UO_172 (O_172,N_28339,N_28706);
nor UO_173 (O_173,N_28424,N_28767);
or UO_174 (O_174,N_29865,N_28792);
xor UO_175 (O_175,N_29505,N_29798);
xor UO_176 (O_176,N_28690,N_29190);
and UO_177 (O_177,N_28061,N_28756);
nor UO_178 (O_178,N_29241,N_28649);
nor UO_179 (O_179,N_29390,N_28684);
xor UO_180 (O_180,N_29608,N_29742);
or UO_181 (O_181,N_29104,N_28545);
or UO_182 (O_182,N_29556,N_29797);
xnor UO_183 (O_183,N_28255,N_28430);
and UO_184 (O_184,N_28570,N_28039);
nand UO_185 (O_185,N_29554,N_28274);
nor UO_186 (O_186,N_28627,N_29106);
nand UO_187 (O_187,N_29473,N_28259);
and UO_188 (O_188,N_28980,N_28897);
xor UO_189 (O_189,N_28954,N_29147);
nor UO_190 (O_190,N_29052,N_28921);
nand UO_191 (O_191,N_28282,N_29762);
xor UO_192 (O_192,N_29982,N_28372);
and UO_193 (O_193,N_28030,N_29134);
and UO_194 (O_194,N_29453,N_28469);
nand UO_195 (O_195,N_28202,N_28977);
nor UO_196 (O_196,N_29981,N_29857);
and UO_197 (O_197,N_29625,N_28740);
nor UO_198 (O_198,N_28386,N_28556);
nor UO_199 (O_199,N_29322,N_29974);
and UO_200 (O_200,N_28208,N_28709);
or UO_201 (O_201,N_29287,N_29717);
nand UO_202 (O_202,N_28804,N_29161);
or UO_203 (O_203,N_28063,N_29012);
nor UO_204 (O_204,N_29591,N_29818);
and UO_205 (O_205,N_29032,N_29181);
and UO_206 (O_206,N_28895,N_29752);
nor UO_207 (O_207,N_28494,N_29826);
and UO_208 (O_208,N_29089,N_29272);
or UO_209 (O_209,N_29398,N_28047);
nor UO_210 (O_210,N_28113,N_28077);
and UO_211 (O_211,N_29285,N_29963);
or UO_212 (O_212,N_29706,N_29804);
and UO_213 (O_213,N_28337,N_28535);
or UO_214 (O_214,N_29175,N_29851);
nand UO_215 (O_215,N_29422,N_28118);
nor UO_216 (O_216,N_29443,N_29145);
and UO_217 (O_217,N_28605,N_28411);
nand UO_218 (O_218,N_28936,N_29078);
or UO_219 (O_219,N_29760,N_29643);
or UO_220 (O_220,N_29266,N_28833);
and UO_221 (O_221,N_28269,N_29569);
nor UO_222 (O_222,N_29714,N_28010);
or UO_223 (O_223,N_29269,N_28546);
xnor UO_224 (O_224,N_28200,N_28753);
nand UO_225 (O_225,N_29239,N_28530);
xnor UO_226 (O_226,N_29922,N_29877);
and UO_227 (O_227,N_29136,N_29967);
nor UO_228 (O_228,N_29855,N_29644);
nand UO_229 (O_229,N_28115,N_28124);
nor UO_230 (O_230,N_29042,N_28665);
xnor UO_231 (O_231,N_29683,N_29491);
nand UO_232 (O_232,N_28760,N_28273);
nand UO_233 (O_233,N_28575,N_28898);
and UO_234 (O_234,N_28802,N_29860);
or UO_235 (O_235,N_28250,N_29265);
nor UO_236 (O_236,N_28376,N_28862);
and UO_237 (O_237,N_29694,N_29438);
nor UO_238 (O_238,N_28095,N_28772);
nor UO_239 (O_239,N_28455,N_29743);
and UO_240 (O_240,N_29357,N_28786);
and UO_241 (O_241,N_28761,N_28593);
nor UO_242 (O_242,N_29096,N_28068);
nand UO_243 (O_243,N_29615,N_29142);
and UO_244 (O_244,N_28172,N_29182);
or UO_245 (O_245,N_28505,N_28896);
and UO_246 (O_246,N_28467,N_28450);
xnor UO_247 (O_247,N_28338,N_28304);
or UO_248 (O_248,N_29132,N_29617);
nand UO_249 (O_249,N_28123,N_28278);
and UO_250 (O_250,N_29533,N_29245);
xor UO_251 (O_251,N_29467,N_28906);
and UO_252 (O_252,N_29611,N_28585);
nor UO_253 (O_253,N_29283,N_28976);
or UO_254 (O_254,N_29113,N_28544);
and UO_255 (O_255,N_29344,N_28799);
or UO_256 (O_256,N_28017,N_29827);
nand UO_257 (O_257,N_29667,N_28568);
and UO_258 (O_258,N_28598,N_28752);
nor UO_259 (O_259,N_29825,N_28602);
nand UO_260 (O_260,N_29538,N_28158);
nor UO_261 (O_261,N_29054,N_29365);
nand UO_262 (O_262,N_29101,N_28843);
or UO_263 (O_263,N_29440,N_28571);
nor UO_264 (O_264,N_29996,N_28600);
or UO_265 (O_265,N_28919,N_29568);
xor UO_266 (O_266,N_29796,N_28671);
and UO_267 (O_267,N_28559,N_28373);
nand UO_268 (O_268,N_28354,N_29497);
nand UO_269 (O_269,N_28949,N_28075);
or UO_270 (O_270,N_29367,N_29935);
or UO_271 (O_271,N_29853,N_28108);
or UO_272 (O_272,N_29721,N_29461);
xor UO_273 (O_273,N_28916,N_28840);
xor UO_274 (O_274,N_28362,N_29374);
xnor UO_275 (O_275,N_29131,N_29657);
and UO_276 (O_276,N_28661,N_29572);
xor UO_277 (O_277,N_28780,N_28161);
and UO_278 (O_278,N_28211,N_28594);
and UO_279 (O_279,N_28195,N_28962);
or UO_280 (O_280,N_29970,N_28447);
or UO_281 (O_281,N_29777,N_28578);
nor UO_282 (O_282,N_28164,N_28399);
xnor UO_283 (O_283,N_28878,N_29472);
nor UO_284 (O_284,N_28587,N_28956);
and UO_285 (O_285,N_28233,N_28563);
nand UO_286 (O_286,N_29688,N_29518);
and UO_287 (O_287,N_28581,N_29133);
nand UO_288 (O_288,N_28080,N_28057);
and UO_289 (O_289,N_29892,N_29424);
or UO_290 (O_290,N_29983,N_29460);
nor UO_291 (O_291,N_28302,N_28301);
xnor UO_292 (O_292,N_28899,N_28361);
nand UO_293 (O_293,N_29841,N_28190);
and UO_294 (O_294,N_29450,N_28909);
nand UO_295 (O_295,N_29868,N_28375);
xor UO_296 (O_296,N_28393,N_29253);
nor UO_297 (O_297,N_29197,N_28937);
nand UO_298 (O_298,N_29129,N_28363);
nand UO_299 (O_299,N_29541,N_29603);
nor UO_300 (O_300,N_28864,N_29565);
or UO_301 (O_301,N_29091,N_28049);
or UO_302 (O_302,N_28714,N_28340);
nor UO_303 (O_303,N_28170,N_29363);
or UO_304 (O_304,N_28220,N_29445);
xnor UO_305 (O_305,N_28715,N_28857);
xnor UO_306 (O_306,N_29658,N_29313);
and UO_307 (O_307,N_28850,N_29270);
and UO_308 (O_308,N_29739,N_29919);
or UO_309 (O_309,N_28903,N_29869);
xor UO_310 (O_310,N_28105,N_29421);
or UO_311 (O_311,N_29381,N_29126);
or UO_312 (O_312,N_29960,N_29817);
or UO_313 (O_313,N_28729,N_28294);
nor UO_314 (O_314,N_28417,N_29448);
or UO_315 (O_315,N_28112,N_29238);
nor UO_316 (O_316,N_28810,N_29433);
xnor UO_317 (O_317,N_29495,N_28029);
nand UO_318 (O_318,N_29361,N_29727);
or UO_319 (O_319,N_28291,N_29243);
or UO_320 (O_320,N_29928,N_28595);
and UO_321 (O_321,N_28087,N_28920);
xor UO_322 (O_322,N_29632,N_28616);
or UO_323 (O_323,N_28003,N_28611);
nor UO_324 (O_324,N_28516,N_28210);
and UO_325 (O_325,N_29858,N_28366);
or UO_326 (O_326,N_28448,N_29837);
or UO_327 (O_327,N_29080,N_29206);
and UO_328 (O_328,N_29669,N_29884);
or UO_329 (O_329,N_29370,N_29766);
xnor UO_330 (O_330,N_29936,N_29408);
xor UO_331 (O_331,N_28918,N_29063);
nor UO_332 (O_332,N_29508,N_29668);
xnor UO_333 (O_333,N_29048,N_28808);
or UO_334 (O_334,N_28945,N_29259);
nor UO_335 (O_335,N_29016,N_29891);
nand UO_336 (O_336,N_28243,N_28181);
xnor UO_337 (O_337,N_28572,N_29786);
and UO_338 (O_338,N_29523,N_28065);
xnor UO_339 (O_339,N_29447,N_29074);
xor UO_340 (O_340,N_28264,N_29305);
xor UO_341 (O_341,N_28965,N_28509);
or UO_342 (O_342,N_29228,N_28787);
nor UO_343 (O_343,N_29666,N_29675);
and UO_344 (O_344,N_28987,N_28044);
and UO_345 (O_345,N_28590,N_29913);
or UO_346 (O_346,N_28579,N_28599);
nor UO_347 (O_347,N_29600,N_29018);
or UO_348 (O_348,N_29312,N_29478);
xor UO_349 (O_349,N_28307,N_28212);
and UO_350 (O_350,N_28180,N_28501);
xor UO_351 (O_351,N_29659,N_28258);
and UO_352 (O_352,N_29620,N_29745);
or UO_353 (O_353,N_29710,N_28292);
nand UO_354 (O_354,N_29838,N_28071);
nor UO_355 (O_355,N_28995,N_29770);
and UO_356 (O_356,N_28438,N_29977);
xnor UO_357 (O_357,N_29562,N_29695);
xor UO_358 (O_358,N_28458,N_28370);
and UO_359 (O_359,N_28507,N_29399);
nand UO_360 (O_360,N_28305,N_29663);
and UO_361 (O_361,N_28187,N_29008);
and UO_362 (O_362,N_29725,N_29582);
and UO_363 (O_363,N_29613,N_29100);
or UO_364 (O_364,N_28838,N_29294);
nand UO_365 (O_365,N_29442,N_29639);
or UO_366 (O_366,N_29999,N_29552);
nor UO_367 (O_367,N_28885,N_29904);
xor UO_368 (O_368,N_28094,N_28131);
xnor UO_369 (O_369,N_29499,N_29358);
nor UO_370 (O_370,N_28656,N_28260);
and UO_371 (O_371,N_29544,N_28157);
xor UO_372 (O_372,N_29268,N_29633);
and UO_373 (O_373,N_28407,N_28367);
xor UO_374 (O_374,N_28360,N_29187);
nor UO_375 (O_375,N_28012,N_29465);
xor UO_376 (O_376,N_29102,N_29962);
nor UO_377 (O_377,N_29566,N_29466);
nor UO_378 (O_378,N_29025,N_29788);
or UO_379 (O_379,N_29907,N_28695);
or UO_380 (O_380,N_29972,N_29616);
and UO_381 (O_381,N_28025,N_29764);
or UO_382 (O_382,N_29338,N_28449);
nor UO_383 (O_383,N_29151,N_28705);
and UO_384 (O_384,N_28142,N_28168);
or UO_385 (O_385,N_29942,N_28018);
nand UO_386 (O_386,N_28560,N_28416);
nand UO_387 (O_387,N_28798,N_28027);
or UO_388 (O_388,N_28827,N_29276);
nor UO_389 (O_389,N_28554,N_28383);
nor UO_390 (O_390,N_28352,N_28062);
nor UO_391 (O_391,N_28289,N_28050);
xor UO_392 (O_392,N_29866,N_28983);
or UO_393 (O_393,N_28645,N_28390);
or UO_394 (O_394,N_28722,N_29360);
nand UO_395 (O_395,N_28688,N_29604);
nand UO_396 (O_396,N_29502,N_28097);
or UO_397 (O_397,N_29592,N_29576);
nor UO_398 (O_398,N_28950,N_29887);
nand UO_399 (O_399,N_29671,N_28648);
or UO_400 (O_400,N_28483,N_28410);
and UO_401 (O_401,N_29264,N_28434);
and UO_402 (O_402,N_29189,N_28474);
and UO_403 (O_403,N_28132,N_29807);
and UO_404 (O_404,N_29010,N_28639);
xnor UO_405 (O_405,N_29373,N_28996);
nor UO_406 (O_406,N_29985,N_28098);
and UO_407 (O_407,N_28900,N_28387);
or UO_408 (O_408,N_28007,N_28790);
nand UO_409 (O_409,N_28232,N_29925);
nand UO_410 (O_410,N_29451,N_28737);
and UO_411 (O_411,N_28088,N_28096);
xor UO_412 (O_412,N_29038,N_29004);
and UO_413 (O_413,N_28676,N_28584);
nor UO_414 (O_414,N_28675,N_29304);
nand UO_415 (O_415,N_28009,N_28267);
and UO_416 (O_416,N_29654,N_28778);
xnor UO_417 (O_417,N_29229,N_28923);
nand UO_418 (O_418,N_29345,N_28985);
nand UO_419 (O_419,N_29014,N_29406);
nand UO_420 (O_420,N_29790,N_29210);
xor UO_421 (O_421,N_29973,N_29749);
nand UO_422 (O_422,N_28066,N_28659);
nor UO_423 (O_423,N_28034,N_28640);
nand UO_424 (O_424,N_28773,N_28868);
nand UO_425 (O_425,N_29127,N_28854);
nand UO_426 (O_426,N_29995,N_28677);
xnor UO_427 (O_427,N_29073,N_29123);
and UO_428 (O_428,N_28078,N_29227);
or UO_429 (O_429,N_28670,N_29154);
and UO_430 (O_430,N_29420,N_28299);
nor UO_431 (O_431,N_29125,N_29515);
xnor UO_432 (O_432,N_28813,N_29109);
nand UO_433 (O_433,N_28491,N_28392);
nor UO_434 (O_434,N_29920,N_28726);
and UO_435 (O_435,N_28234,N_29929);
or UO_436 (O_436,N_29498,N_28836);
or UO_437 (O_437,N_29039,N_29144);
nor UO_438 (O_438,N_28927,N_28825);
nor UO_439 (O_439,N_29949,N_28762);
and UO_440 (O_440,N_28618,N_28277);
nor UO_441 (O_441,N_29629,N_28689);
or UO_442 (O_442,N_29307,N_28054);
nor UO_443 (O_443,N_28646,N_29814);
and UO_444 (O_444,N_29750,N_29319);
and UO_445 (O_445,N_29290,N_28041);
nor UO_446 (O_446,N_28940,N_28614);
nor UO_447 (O_447,N_28942,N_29009);
or UO_448 (O_448,N_29204,N_28569);
or UO_449 (O_449,N_29115,N_29696);
xor UO_450 (O_450,N_28295,N_28379);
xor UO_451 (O_451,N_29630,N_29051);
and UO_452 (O_452,N_28928,N_28194);
or UO_453 (O_453,N_29909,N_29346);
xor UO_454 (O_454,N_29208,N_28515);
and UO_455 (O_455,N_28252,N_29624);
nand UO_456 (O_456,N_29274,N_28151);
xnor UO_457 (O_457,N_28984,N_28521);
and UO_458 (O_458,N_28805,N_29483);
or UO_459 (O_459,N_29829,N_28283);
nand UO_460 (O_460,N_29734,N_29485);
and UO_461 (O_461,N_28004,N_29315);
or UO_462 (O_462,N_28271,N_29477);
or UO_463 (O_463,N_29303,N_28127);
xor UO_464 (O_464,N_29174,N_29417);
xor UO_465 (O_465,N_28794,N_28312);
nand UO_466 (O_466,N_29023,N_29171);
or UO_467 (O_467,N_28129,N_29614);
and UO_468 (O_468,N_29397,N_29156);
and UO_469 (O_469,N_29778,N_28320);
or UO_470 (O_470,N_29959,N_29914);
nand UO_471 (O_471,N_28989,N_28914);
and UO_472 (O_472,N_29889,N_29641);
nor UO_473 (O_473,N_29579,N_29083);
nand UO_474 (O_474,N_28951,N_29885);
nand UO_475 (O_475,N_28669,N_29138);
nor UO_476 (O_476,N_29061,N_29886);
xnor UO_477 (O_477,N_28889,N_28191);
xor UO_478 (O_478,N_28353,N_28713);
or UO_479 (O_479,N_28415,N_28710);
nor UO_480 (O_480,N_28520,N_28526);
or UO_481 (O_481,N_29394,N_29140);
or UO_482 (O_482,N_28832,N_29223);
xor UO_483 (O_483,N_29267,N_28245);
nor UO_484 (O_484,N_29716,N_28541);
xnor UO_485 (O_485,N_28215,N_29153);
nor UO_486 (O_486,N_29257,N_28664);
nand UO_487 (O_487,N_28818,N_29843);
or UO_488 (O_488,N_29256,N_29791);
nor UO_489 (O_489,N_28948,N_28946);
nor UO_490 (O_490,N_29000,N_29260);
and UO_491 (O_491,N_28074,N_28668);
xnor UO_492 (O_492,N_29117,N_29697);
nand UO_493 (O_493,N_29780,N_29186);
and UO_494 (O_494,N_28006,N_29723);
nand UO_495 (O_495,N_29530,N_28314);
nand UO_496 (O_496,N_29475,N_29456);
nor UO_497 (O_497,N_28330,N_29275);
or UO_498 (O_498,N_29376,N_29387);
xor UO_499 (O_499,N_29026,N_28502);
nor UO_500 (O_500,N_28359,N_28222);
or UO_501 (O_501,N_29327,N_28938);
nand UO_502 (O_502,N_28623,N_29816);
xnor UO_503 (O_503,N_28221,N_29284);
and UO_504 (O_504,N_28742,N_28552);
and UO_505 (O_505,N_28420,N_28518);
and UO_506 (O_506,N_28348,N_28894);
nor UO_507 (O_507,N_28955,N_28481);
and UO_508 (O_508,N_28972,N_29834);
or UO_509 (O_509,N_29480,N_29768);
nand UO_510 (O_510,N_28748,N_29191);
nand UO_511 (O_511,N_28957,N_28553);
nor UO_512 (O_512,N_29845,N_29832);
or UO_513 (O_513,N_29057,N_29785);
nor UO_514 (O_514,N_29705,N_28102);
or UO_515 (O_515,N_29978,N_29765);
and UO_516 (O_516,N_28153,N_29622);
nand UO_517 (O_517,N_28538,N_29652);
or UO_518 (O_518,N_29022,N_29446);
xor UO_519 (O_519,N_29522,N_28619);
nand UO_520 (O_520,N_29787,N_28634);
or UO_521 (O_521,N_29943,N_29076);
nand UO_522 (O_522,N_28893,N_29908);
nor UO_523 (O_523,N_28008,N_28536);
and UO_524 (O_524,N_29651,N_28461);
and UO_525 (O_525,N_28043,N_29840);
and UO_526 (O_526,N_28759,N_28103);
nand UO_527 (O_527,N_29874,N_29836);
nor UO_528 (O_528,N_28573,N_29883);
nand UO_529 (O_529,N_29428,N_28333);
nor UO_530 (O_530,N_28389,N_28743);
and UO_531 (O_531,N_28175,N_29690);
and UO_532 (O_532,N_28511,N_29060);
nand UO_533 (O_533,N_29413,N_28537);
nand UO_534 (O_534,N_29720,N_28929);
xnor UO_535 (O_535,N_29934,N_29800);
or UO_536 (O_536,N_29545,N_29783);
or UO_537 (O_537,N_28755,N_29610);
nand UO_538 (O_538,N_29007,N_28031);
and UO_539 (O_539,N_28596,N_28567);
nand UO_540 (O_540,N_29248,N_29314);
or UO_541 (O_541,N_28651,N_28635);
nand UO_542 (O_542,N_28636,N_28152);
nor UO_543 (O_543,N_28694,N_29306);
nor UO_544 (O_544,N_29302,N_29747);
or UO_545 (O_545,N_29691,N_29481);
or UO_546 (O_546,N_28268,N_29953);
or UO_547 (O_547,N_29687,N_28496);
xnor UO_548 (O_548,N_28328,N_28522);
xnor UO_549 (O_549,N_29811,N_28971);
and UO_550 (O_550,N_28439,N_28795);
or UO_551 (O_551,N_29335,N_28462);
xnor UO_552 (O_552,N_29219,N_28674);
nor UO_553 (O_553,N_28966,N_29484);
xor UO_554 (O_554,N_28824,N_29862);
nor UO_555 (O_555,N_28917,N_28504);
xnor UO_556 (O_556,N_28871,N_28835);
and UO_557 (O_557,N_28834,N_29482);
or UO_558 (O_558,N_28303,N_28698);
or UO_559 (O_559,N_29521,N_28464);
xnor UO_560 (O_560,N_29975,N_29820);
xnor UO_561 (O_561,N_29677,N_28524);
xor UO_562 (O_562,N_28432,N_29757);
nor UO_563 (O_563,N_29931,N_29258);
and UO_564 (O_564,N_28457,N_29163);
or UO_565 (O_565,N_28263,N_29507);
and UO_566 (O_566,N_28315,N_29071);
nand UO_567 (O_567,N_28588,N_28397);
nor UO_568 (O_568,N_28924,N_29806);
or UO_569 (O_569,N_29809,N_29645);
nor UO_570 (O_570,N_29506,N_29316);
xor UO_571 (O_571,N_29255,N_28608);
nand UO_572 (O_572,N_28242,N_29589);
or UO_573 (O_573,N_28056,N_29954);
xnor UO_574 (O_574,N_29938,N_28683);
nand UO_575 (O_575,N_29618,N_28548);
nand UO_576 (O_576,N_29563,N_29098);
and UO_577 (O_577,N_29231,N_28114);
and UO_578 (O_578,N_29700,N_29713);
nand UO_579 (O_579,N_28182,N_28414);
or UO_580 (O_580,N_28880,N_28165);
nand UO_581 (O_581,N_29251,N_29193);
nand UO_582 (O_582,N_28691,N_28484);
xor UO_583 (O_583,N_29898,N_29950);
nand UO_584 (O_584,N_28431,N_28696);
nor UO_585 (O_585,N_29462,N_28381);
xnor UO_586 (O_586,N_28028,N_29099);
or UO_587 (O_587,N_29059,N_29107);
nand UO_588 (O_588,N_28935,N_28973);
nand UO_589 (O_589,N_28011,N_29813);
xor UO_590 (O_590,N_29389,N_28697);
nand UO_591 (O_591,N_28155,N_28879);
or UO_592 (O_592,N_28866,N_29940);
or UO_593 (O_593,N_28734,N_29879);
xor UO_594 (O_594,N_29331,N_28716);
nor UO_595 (O_595,N_29211,N_29729);
nand UO_596 (O_596,N_28189,N_28915);
nand UO_597 (O_597,N_28327,N_29941);
nor UO_598 (O_598,N_29254,N_28606);
or UO_599 (O_599,N_29085,N_28701);
nand UO_600 (O_600,N_28724,N_29564);
nand UO_601 (O_601,N_29247,N_29105);
xor UO_602 (O_602,N_28667,N_29362);
xnor UO_603 (O_603,N_28644,N_28750);
and UO_604 (O_604,N_28249,N_29234);
and UO_605 (O_605,N_28279,N_28427);
xor UO_606 (O_606,N_28219,N_28216);
and UO_607 (O_607,N_28986,N_28823);
nand UO_608 (O_608,N_29015,N_29468);
nor UO_609 (O_609,N_29218,N_28800);
or UO_610 (O_610,N_29409,N_28741);
nor UO_611 (O_611,N_28855,N_29731);
nor UO_612 (O_612,N_28223,N_28628);
xor UO_613 (O_613,N_28680,N_28371);
and UO_614 (O_614,N_29875,N_29854);
or UO_615 (O_615,N_28844,N_29876);
nor UO_616 (O_616,N_28939,N_29236);
xor UO_617 (O_617,N_28137,N_29581);
nand UO_618 (O_618,N_29045,N_28479);
nand UO_619 (O_619,N_29332,N_29205);
nor UO_620 (O_620,N_28385,N_29250);
or UO_621 (O_621,N_29520,N_28540);
and UO_622 (O_622,N_28236,N_28206);
or UO_623 (O_623,N_28510,N_28781);
and UO_624 (O_624,N_29110,N_29989);
nand UO_625 (O_625,N_29490,N_29224);
nand UO_626 (O_626,N_28149,N_29763);
nor UO_627 (O_627,N_29672,N_28356);
or UO_628 (O_628,N_29621,N_28700);
or UO_629 (O_629,N_29383,N_29375);
and UO_630 (O_630,N_28468,N_28257);
nand UO_631 (O_631,N_29548,N_29528);
xor UO_632 (O_632,N_29635,N_28806);
nor UO_633 (O_633,N_29586,N_28321);
nand UO_634 (O_634,N_28001,N_29646);
xnor UO_635 (O_635,N_29537,N_28933);
nor UO_636 (O_636,N_29775,N_28107);
xor UO_637 (O_637,N_29427,N_28388);
nand UO_638 (O_638,N_29277,N_29755);
or UO_639 (O_639,N_28121,N_29689);
nand UO_640 (O_640,N_29396,N_29149);
xor UO_641 (O_641,N_28564,N_28286);
or UO_642 (O_642,N_29574,N_29043);
and UO_643 (O_643,N_28134,N_29542);
xnor UO_644 (O_644,N_29425,N_29965);
xor UO_645 (O_645,N_29636,N_29086);
and UO_646 (O_646,N_29377,N_29769);
xnor UO_647 (O_647,N_29308,N_29135);
and UO_648 (O_648,N_29415,N_29405);
nor UO_649 (O_649,N_29979,N_28256);
and UO_650 (O_650,N_28178,N_28398);
and UO_651 (O_651,N_28841,N_28485);
xnor UO_652 (O_652,N_29431,N_29214);
nand UO_653 (O_653,N_29120,N_29271);
or UO_654 (O_654,N_28069,N_29001);
nand UO_655 (O_655,N_29880,N_29557);
xor UO_656 (O_656,N_29075,N_29047);
and UO_657 (O_657,N_28024,N_28241);
nand UO_658 (O_658,N_28082,N_29998);
or UO_659 (O_659,N_28495,N_29712);
nand UO_660 (O_660,N_29653,N_29911);
xor UO_661 (O_661,N_29281,N_28807);
xnor UO_662 (O_662,N_29684,N_28128);
and UO_663 (O_663,N_28637,N_28902);
and UO_664 (O_664,N_29681,N_29730);
nand UO_665 (O_665,N_28266,N_29027);
xnor UO_666 (O_666,N_28770,N_28346);
nand UO_667 (O_667,N_29708,N_29240);
nor UO_668 (O_668,N_29561,N_28631);
nand UO_669 (O_669,N_29201,N_28429);
nor UO_670 (O_670,N_28968,N_29584);
and UO_671 (O_671,N_28580,N_29432);
nor UO_672 (O_672,N_28652,N_29386);
or UO_673 (O_673,N_29444,N_28655);
xnor UO_674 (O_674,N_28500,N_29754);
or UO_675 (O_675,N_29094,N_29531);
xnor UO_676 (O_676,N_28247,N_28859);
and UO_677 (O_677,N_28812,N_29864);
xnor UO_678 (O_678,N_29464,N_29340);
nor UO_679 (O_679,N_29634,N_29605);
xnor UO_680 (O_680,N_28230,N_29839);
nor UO_681 (O_681,N_29170,N_29846);
nor UO_682 (O_682,N_29055,N_29656);
nor UO_683 (O_683,N_29740,N_28555);
and UO_684 (O_684,N_28992,N_28072);
and UO_685 (O_685,N_29988,N_29597);
or UO_686 (O_686,N_28120,N_28171);
nand UO_687 (O_687,N_28783,N_29558);
xnor UO_688 (O_688,N_29894,N_29882);
or UO_689 (O_689,N_29119,N_29924);
xor UO_690 (O_690,N_28860,N_29280);
nand UO_691 (O_691,N_29232,N_29664);
or UO_692 (O_692,N_29400,N_29392);
xnor UO_693 (O_693,N_29955,N_28757);
or UO_694 (O_694,N_28814,N_28076);
or UO_695 (O_695,N_28849,N_29309);
and UO_696 (O_696,N_28343,N_29598);
and UO_697 (O_697,N_29751,N_28311);
and UO_698 (O_698,N_28167,N_29872);
xnor UO_699 (O_699,N_28852,N_28042);
or UO_700 (O_700,N_28465,N_28240);
or UO_701 (O_701,N_28136,N_28562);
and UO_702 (O_702,N_28183,N_29585);
nor UO_703 (O_703,N_28534,N_28711);
or UO_704 (O_704,N_28601,N_29670);
nor UO_705 (O_705,N_28119,N_29628);
and UO_706 (O_706,N_28666,N_29930);
xor UO_707 (O_707,N_29607,N_28934);
nor UO_708 (O_708,N_29753,N_28620);
nor UO_709 (O_709,N_28146,N_29792);
or UO_710 (O_710,N_29353,N_28405);
nor UO_711 (O_711,N_28045,N_29631);
nand UO_712 (O_712,N_28542,N_28532);
and UO_713 (O_713,N_29501,N_29759);
xor UO_714 (O_714,N_28037,N_29006);
or UO_715 (O_715,N_29529,N_28248);
nand UO_716 (O_716,N_28176,N_29310);
nand UO_717 (O_717,N_28603,N_29709);
or UO_718 (O_718,N_28872,N_28941);
xnor UO_719 (O_719,N_28870,N_29906);
and UO_720 (O_720,N_28621,N_28441);
xor UO_721 (O_721,N_28566,N_28192);
nand UO_722 (O_722,N_28419,N_29500);
or UO_723 (O_723,N_29323,N_28910);
or UO_724 (O_724,N_29905,N_28846);
nor UO_725 (O_725,N_28642,N_29890);
nand UO_726 (O_726,N_29805,N_28845);
and UO_727 (O_727,N_28638,N_28882);
nor UO_728 (O_728,N_29416,N_28883);
nand UO_729 (O_729,N_29986,N_29173);
xor UO_730 (O_730,N_28475,N_28533);
or UO_731 (O_731,N_29535,N_28403);
nor UO_732 (O_732,N_29601,N_29169);
and UO_733 (O_733,N_29701,N_29517);
nand UO_734 (O_734,N_28960,N_28704);
xnor UO_735 (O_735,N_28531,N_29019);
nor UO_736 (O_736,N_29459,N_28877);
xnor UO_737 (O_737,N_29987,N_28163);
and UO_738 (O_738,N_28159,N_29068);
nand UO_739 (O_739,N_29036,N_28412);
xnor UO_740 (O_740,N_29551,N_28815);
nand UO_741 (O_741,N_29692,N_29176);
xor UO_742 (O_742,N_28196,N_28731);
nand UO_743 (O_743,N_28817,N_28686);
and UO_744 (O_744,N_29711,N_28747);
nand UO_745 (O_745,N_29594,N_29273);
xor UO_746 (O_746,N_29944,N_29056);
xnor UO_747 (O_747,N_29599,N_29293);
and UO_748 (O_748,N_28488,N_28480);
and UO_749 (O_749,N_29665,N_29559);
and UO_750 (O_750,N_29002,N_28816);
nor UO_751 (O_751,N_28863,N_28609);
nor UO_752 (O_752,N_28324,N_29650);
nor UO_753 (O_753,N_28723,N_29915);
nor UO_754 (O_754,N_28036,N_28205);
nor UO_755 (O_755,N_28779,N_28261);
nand UO_756 (O_756,N_28493,N_29503);
nor UO_757 (O_757,N_29655,N_29831);
and UO_758 (O_758,N_29933,N_29593);
and UO_759 (O_759,N_29458,N_28582);
and UO_760 (O_760,N_29781,N_28470);
xnor UO_761 (O_761,N_28213,N_29359);
and UO_762 (O_762,N_29474,N_29910);
or UO_763 (O_763,N_29830,N_28607);
or UO_764 (O_764,N_29379,N_29848);
xnor UO_765 (O_765,N_29850,N_28732);
xnor UO_766 (O_766,N_28201,N_28251);
nor UO_767 (O_767,N_28612,N_28967);
xor UO_768 (O_768,N_29513,N_29198);
or UO_769 (O_769,N_29612,N_29994);
and UO_770 (O_770,N_28138,N_29738);
or UO_771 (O_771,N_28615,N_29789);
xor UO_772 (O_772,N_29199,N_29380);
or UO_773 (O_773,N_28126,N_28826);
nor UO_774 (O_774,N_29516,N_29320);
and UO_775 (O_775,N_29035,N_28617);
nand UO_776 (O_776,N_29300,N_29509);
xor UO_777 (O_777,N_28401,N_28746);
or UO_778 (O_778,N_29852,N_28145);
and UO_779 (O_779,N_28653,N_28199);
nand UO_780 (O_780,N_29627,N_28331);
xnor UO_781 (O_781,N_29455,N_29961);
or UO_782 (O_782,N_28797,N_28174);
nand UO_783 (O_783,N_29642,N_29997);
and UO_784 (O_784,N_28197,N_29329);
nor UO_785 (O_785,N_29682,N_29041);
nand UO_786 (O_786,N_29492,N_28926);
or UO_787 (O_787,N_28002,N_29916);
nand UO_788 (O_788,N_29590,N_29771);
and UO_789 (O_789,N_29356,N_28297);
or UO_790 (O_790,N_29772,N_29486);
or UO_791 (O_791,N_28306,N_28290);
nand UO_792 (O_792,N_29926,N_29337);
nand UO_793 (O_793,N_28574,N_29414);
or UO_794 (O_794,N_29454,N_29947);
nor UO_795 (O_795,N_29402,N_29990);
or UO_796 (O_796,N_29776,N_29976);
xor UO_797 (O_797,N_28026,N_29801);
or UO_798 (O_798,N_29948,N_29937);
xnor UO_799 (O_799,N_29719,N_28035);
nand UO_800 (O_800,N_28842,N_28979);
or UO_801 (O_801,N_29412,N_29070);
xnor UO_802 (O_802,N_29575,N_29647);
nand UO_803 (O_803,N_28089,N_29430);
and UO_804 (O_804,N_29900,N_29348);
xnor UO_805 (O_805,N_29139,N_28576);
and UO_806 (O_806,N_28657,N_28766);
nand UO_807 (O_807,N_28309,N_29514);
and UO_808 (O_808,N_29971,N_28685);
xnor UO_809 (O_809,N_28038,N_29945);
nor UO_810 (O_810,N_28253,N_28730);
xor UO_811 (O_811,N_29366,N_29793);
and UO_812 (O_812,N_29779,N_29090);
and UO_813 (O_813,N_29893,N_28837);
nand UO_814 (O_814,N_28876,N_29215);
nand UO_815 (O_815,N_28788,N_28736);
nand UO_816 (O_816,N_28293,N_28203);
nor UO_817 (O_817,N_29488,N_29326);
nand UO_818 (O_818,N_29939,N_28527);
xor UO_819 (O_819,N_29121,N_28184);
nor UO_820 (O_820,N_28990,N_28454);
xor UO_821 (O_821,N_28378,N_28101);
nor UO_822 (O_822,N_28019,N_28991);
or UO_823 (O_823,N_29828,N_29540);
nand UO_824 (O_824,N_28109,N_28673);
or UO_825 (O_825,N_28774,N_29262);
or UO_826 (O_826,N_29549,N_29736);
and UO_827 (O_827,N_28166,N_28368);
and UO_828 (O_828,N_29871,N_29746);
nor UO_829 (O_829,N_28275,N_28506);
nor UO_830 (O_830,N_28486,N_28970);
nor UO_831 (O_831,N_28720,N_29195);
and UO_832 (O_832,N_28437,N_29202);
nand UO_833 (O_833,N_28908,N_28482);
nand UO_834 (O_834,N_29580,N_28369);
or UO_835 (O_835,N_28931,N_28643);
nor UO_836 (O_836,N_28891,N_28944);
nor UO_837 (O_837,N_29225,N_28809);
nor UO_838 (O_838,N_28820,N_29964);
nor UO_839 (O_839,N_29543,N_29029);
and UO_840 (O_840,N_28513,N_28525);
xnor UO_841 (O_841,N_28503,N_28433);
xnor UO_842 (O_842,N_29324,N_29318);
xnor UO_843 (O_843,N_28660,N_29244);
nand UO_844 (O_844,N_29849,N_28015);
and UO_845 (O_845,N_28793,N_28377);
or UO_846 (O_846,N_29679,N_28892);
nand UO_847 (O_847,N_29108,N_28020);
xor UO_848 (O_848,N_28848,N_28048);
or UO_849 (O_849,N_28687,N_28699);
and UO_850 (O_850,N_29429,N_29194);
nor UO_851 (O_851,N_29200,N_29735);
xnor UO_852 (O_852,N_28316,N_28981);
nand UO_853 (O_853,N_29812,N_28085);
or UO_854 (O_854,N_28851,N_29527);
xnor UO_855 (O_855,N_28342,N_29371);
and UO_856 (O_856,N_28994,N_28708);
nand UO_857 (O_857,N_29297,N_29164);
and UO_858 (O_858,N_28409,N_28350);
nor UO_859 (O_859,N_28745,N_29702);
xor UO_860 (O_860,N_29547,N_29487);
and UO_861 (O_861,N_29050,N_28110);
nor UO_862 (O_862,N_29463,N_29824);
nand UO_863 (O_863,N_28147,N_28719);
nor UO_864 (O_864,N_29423,N_29192);
or UO_865 (O_865,N_28822,N_28725);
nor UO_866 (O_866,N_28100,N_29993);
nor UO_867 (O_867,N_29278,N_28144);
nor UO_868 (O_868,N_28442,N_29992);
nand UO_869 (O_869,N_28943,N_29469);
nand UO_870 (O_870,N_28086,N_28777);
nor UO_871 (O_871,N_29741,N_29861);
and UO_872 (O_872,N_28789,N_29364);
xor UO_873 (O_873,N_28083,N_28517);
nand UO_874 (O_874,N_29867,N_29368);
nand UO_875 (O_875,N_29067,N_29343);
nor UO_876 (O_876,N_28884,N_28847);
nor UO_877 (O_877,N_28764,N_29148);
or UO_878 (O_878,N_28629,N_29298);
nor UO_879 (O_879,N_29626,N_29291);
and UO_880 (O_880,N_29733,N_29157);
xor UO_881 (O_881,N_29141,N_28853);
or UO_882 (O_882,N_28886,N_28477);
and UO_883 (O_883,N_28380,N_29328);
or UO_884 (O_884,N_28583,N_29808);
xor UO_885 (O_885,N_29457,N_28382);
or UO_886 (O_886,N_29069,N_28550);
xor UO_887 (O_887,N_28408,N_28046);
xor UO_888 (O_888,N_29178,N_29418);
or UO_889 (O_889,N_28186,N_29744);
and UO_890 (O_890,N_29404,N_29103);
nor UO_891 (O_891,N_29252,N_28418);
and UO_892 (O_892,N_29842,N_29870);
nand UO_893 (O_893,N_29918,N_29330);
nand UO_894 (O_894,N_28139,N_29342);
and UO_895 (O_895,N_29555,N_29382);
or UO_896 (O_896,N_29005,N_29395);
and UO_897 (O_897,N_28890,N_28308);
xor UO_898 (O_898,N_28023,N_28964);
xor UO_899 (O_899,N_29958,N_28231);
or UO_900 (O_900,N_28728,N_28904);
xnor UO_901 (O_901,N_28318,N_28632);
and UO_902 (O_902,N_29166,N_28141);
nand UO_903 (O_903,N_29449,N_29888);
and UO_904 (O_904,N_29835,N_29388);
nor UO_905 (O_905,N_28861,N_29511);
or UO_906 (O_906,N_29470,N_28514);
nor UO_907 (O_907,N_28237,N_28188);
nand UO_908 (O_908,N_29082,N_28093);
or UO_909 (O_909,N_28735,N_29847);
or UO_910 (O_910,N_29856,N_28969);
nor UO_911 (O_911,N_29512,N_28565);
or UO_912 (O_912,N_28999,N_29044);
or UO_913 (O_913,N_29897,N_29724);
nand UO_914 (O_914,N_29249,N_29951);
nand UO_915 (O_915,N_29435,N_29064);
and UO_916 (O_916,N_28135,N_28993);
and UO_917 (O_917,N_28270,N_29289);
nor UO_918 (O_918,N_29821,N_29899);
nor UO_919 (O_919,N_28953,N_28084);
xor UO_920 (O_920,N_28519,N_29833);
and UO_921 (O_921,N_29024,N_29311);
or UO_922 (O_922,N_28839,N_29878);
nand UO_923 (O_923,N_29573,N_28423);
and UO_924 (O_924,N_28032,N_28140);
and UO_925 (O_925,N_28911,N_28284);
nor UO_926 (O_926,N_29233,N_28336);
xnor UO_927 (O_927,N_29350,N_29217);
xor UO_928 (O_928,N_28604,N_29221);
nor UO_929 (O_929,N_28005,N_28801);
nor UO_930 (O_930,N_29088,N_28982);
nand UO_931 (O_931,N_29352,N_28681);
nor UO_932 (O_932,N_29341,N_29209);
and UO_933 (O_933,N_28013,N_29111);
and UO_934 (O_934,N_29180,N_29638);
nor UO_935 (O_935,N_29033,N_28803);
and UO_936 (O_936,N_28589,N_28473);
and UO_937 (O_937,N_28358,N_29496);
nand UO_938 (O_938,N_29172,N_28875);
nor UO_939 (O_939,N_29623,N_29160);
xnor UO_940 (O_940,N_29903,N_28106);
xnor UO_941 (O_941,N_29028,N_28055);
and UO_942 (O_942,N_29393,N_29299);
and UO_943 (O_943,N_28422,N_28597);
xnor UO_944 (O_944,N_28428,N_29150);
and UO_945 (O_945,N_28117,N_29183);
or UO_946 (O_946,N_28351,N_28997);
nand UO_947 (O_947,N_29471,N_29619);
or UO_948 (O_948,N_29640,N_29020);
nor UO_949 (O_949,N_28143,N_28173);
and UO_950 (O_950,N_29385,N_28310);
and UO_951 (O_951,N_28224,N_28022);
or UO_952 (O_952,N_29407,N_29494);
nor UO_953 (O_953,N_28558,N_29550);
or UO_954 (O_954,N_29230,N_29534);
and UO_955 (O_955,N_29212,N_28988);
or UO_956 (O_956,N_28125,N_29767);
nand UO_957 (O_957,N_29758,N_28425);
xnor UO_958 (O_958,N_28451,N_29349);
nor UO_959 (O_959,N_28830,N_29479);
and UO_960 (O_960,N_28626,N_29901);
nand UO_961 (O_961,N_29021,N_29122);
nand UO_962 (O_962,N_29031,N_29196);
and UO_963 (O_963,N_28776,N_28828);
nand UO_964 (O_964,N_29143,N_28641);
and UO_965 (O_965,N_28658,N_29927);
xor UO_966 (O_966,N_28721,N_28053);
nand UO_967 (O_967,N_28154,N_28478);
and UO_968 (O_968,N_29966,N_28064);
or UO_969 (O_969,N_28551,N_29317);
nor UO_970 (O_970,N_29226,N_28549);
and UO_971 (O_971,N_28254,N_29748);
or UO_972 (O_972,N_28313,N_29693);
and UO_973 (O_973,N_29526,N_29152);
nor UO_974 (O_974,N_28347,N_28413);
xor UO_975 (O_975,N_28577,N_29003);
xnor UO_976 (O_976,N_28975,N_28148);
nor UO_977 (O_977,N_28058,N_29046);
and UO_978 (O_978,N_28930,N_28228);
nor UO_979 (O_979,N_29116,N_29957);
nand UO_980 (O_980,N_28204,N_28443);
xor UO_981 (O_981,N_29286,N_29595);
nor UO_982 (O_982,N_29282,N_28539);
or UO_983 (O_983,N_28959,N_28678);
xnor UO_984 (O_984,N_28021,N_29092);
nor UO_985 (O_985,N_28487,N_29686);
nand UO_986 (O_986,N_29567,N_28456);
or UO_987 (O_987,N_29207,N_28067);
nor UO_988 (O_988,N_28402,N_28528);
xnor UO_989 (O_989,N_29784,N_28932);
xnor UO_990 (O_990,N_28179,N_29673);
nor UO_991 (O_991,N_29403,N_28703);
xor UO_992 (O_992,N_28874,N_29968);
or UO_993 (O_993,N_29795,N_29715);
nor UO_994 (O_994,N_29969,N_28091);
and UO_995 (O_995,N_29609,N_28287);
nor UO_996 (O_996,N_28769,N_28444);
or UO_997 (O_997,N_29185,N_28225);
xor UO_998 (O_998,N_28453,N_29844);
nor UO_999 (O_999,N_28881,N_28300);
nor UO_1000 (O_1000,N_29630,N_28674);
nand UO_1001 (O_1001,N_28189,N_29548);
and UO_1002 (O_1002,N_28074,N_29722);
nor UO_1003 (O_1003,N_29516,N_29885);
xnor UO_1004 (O_1004,N_28515,N_28544);
or UO_1005 (O_1005,N_28040,N_29809);
or UO_1006 (O_1006,N_28599,N_28395);
nand UO_1007 (O_1007,N_29272,N_29684);
or UO_1008 (O_1008,N_29061,N_28626);
nor UO_1009 (O_1009,N_29040,N_29867);
and UO_1010 (O_1010,N_29603,N_29630);
xnor UO_1011 (O_1011,N_29830,N_28742);
and UO_1012 (O_1012,N_29463,N_28289);
or UO_1013 (O_1013,N_28968,N_29078);
nand UO_1014 (O_1014,N_29016,N_28354);
or UO_1015 (O_1015,N_29578,N_29136);
and UO_1016 (O_1016,N_29371,N_28170);
or UO_1017 (O_1017,N_29761,N_29450);
and UO_1018 (O_1018,N_28224,N_29565);
nand UO_1019 (O_1019,N_29102,N_28679);
nor UO_1020 (O_1020,N_28936,N_29534);
and UO_1021 (O_1021,N_28438,N_29945);
nor UO_1022 (O_1022,N_29200,N_28034);
and UO_1023 (O_1023,N_28376,N_29320);
and UO_1024 (O_1024,N_28252,N_28572);
nor UO_1025 (O_1025,N_28228,N_29267);
xor UO_1026 (O_1026,N_29233,N_28416);
nand UO_1027 (O_1027,N_29501,N_28460);
and UO_1028 (O_1028,N_29056,N_28265);
nor UO_1029 (O_1029,N_28050,N_28635);
and UO_1030 (O_1030,N_28651,N_29323);
nor UO_1031 (O_1031,N_29780,N_29820);
nand UO_1032 (O_1032,N_29226,N_28395);
nand UO_1033 (O_1033,N_29059,N_29877);
and UO_1034 (O_1034,N_28298,N_28216);
xnor UO_1035 (O_1035,N_28609,N_29466);
and UO_1036 (O_1036,N_29407,N_28441);
xor UO_1037 (O_1037,N_29348,N_29439);
nor UO_1038 (O_1038,N_29694,N_29451);
xor UO_1039 (O_1039,N_28011,N_28868);
and UO_1040 (O_1040,N_28370,N_29374);
or UO_1041 (O_1041,N_29339,N_28599);
nand UO_1042 (O_1042,N_28043,N_29748);
or UO_1043 (O_1043,N_28776,N_29549);
or UO_1044 (O_1044,N_29424,N_29231);
xnor UO_1045 (O_1045,N_28937,N_29974);
nand UO_1046 (O_1046,N_29640,N_29858);
nor UO_1047 (O_1047,N_29638,N_28179);
nor UO_1048 (O_1048,N_28568,N_28822);
nor UO_1049 (O_1049,N_29707,N_29451);
or UO_1050 (O_1050,N_28429,N_29761);
nor UO_1051 (O_1051,N_29928,N_28466);
nand UO_1052 (O_1052,N_29414,N_29542);
nand UO_1053 (O_1053,N_29188,N_28903);
nand UO_1054 (O_1054,N_29550,N_29236);
or UO_1055 (O_1055,N_28918,N_28342);
or UO_1056 (O_1056,N_29542,N_29461);
nand UO_1057 (O_1057,N_29517,N_29231);
xnor UO_1058 (O_1058,N_29536,N_28660);
and UO_1059 (O_1059,N_29833,N_29886);
nand UO_1060 (O_1060,N_28163,N_29604);
nand UO_1061 (O_1061,N_28549,N_28917);
nand UO_1062 (O_1062,N_29663,N_28097);
nor UO_1063 (O_1063,N_28296,N_28314);
or UO_1064 (O_1064,N_28791,N_29904);
nor UO_1065 (O_1065,N_28128,N_29400);
nand UO_1066 (O_1066,N_28099,N_29916);
nor UO_1067 (O_1067,N_28630,N_29927);
nor UO_1068 (O_1068,N_28182,N_28435);
nand UO_1069 (O_1069,N_29386,N_28670);
nor UO_1070 (O_1070,N_29094,N_29752);
xnor UO_1071 (O_1071,N_29006,N_28314);
or UO_1072 (O_1072,N_28841,N_28416);
and UO_1073 (O_1073,N_29438,N_29428);
xor UO_1074 (O_1074,N_28769,N_28422);
nand UO_1075 (O_1075,N_28161,N_28546);
and UO_1076 (O_1076,N_28805,N_29772);
nor UO_1077 (O_1077,N_28051,N_29272);
and UO_1078 (O_1078,N_28017,N_29363);
nor UO_1079 (O_1079,N_28774,N_28172);
or UO_1080 (O_1080,N_28000,N_28778);
or UO_1081 (O_1081,N_28542,N_29588);
nor UO_1082 (O_1082,N_28389,N_29339);
and UO_1083 (O_1083,N_29472,N_28517);
nor UO_1084 (O_1084,N_29910,N_28789);
nor UO_1085 (O_1085,N_29764,N_28869);
xnor UO_1086 (O_1086,N_28074,N_29986);
xnor UO_1087 (O_1087,N_28357,N_29805);
nand UO_1088 (O_1088,N_29166,N_28137);
nand UO_1089 (O_1089,N_29477,N_28423);
xor UO_1090 (O_1090,N_28508,N_28023);
and UO_1091 (O_1091,N_29546,N_29954);
and UO_1092 (O_1092,N_28139,N_29702);
xnor UO_1093 (O_1093,N_28491,N_28190);
nand UO_1094 (O_1094,N_28446,N_29985);
or UO_1095 (O_1095,N_29044,N_28343);
or UO_1096 (O_1096,N_28449,N_29074);
or UO_1097 (O_1097,N_29803,N_28973);
nand UO_1098 (O_1098,N_28491,N_28844);
or UO_1099 (O_1099,N_29028,N_28422);
or UO_1100 (O_1100,N_28072,N_28629);
nand UO_1101 (O_1101,N_28453,N_28839);
or UO_1102 (O_1102,N_29455,N_29476);
nor UO_1103 (O_1103,N_28959,N_29094);
and UO_1104 (O_1104,N_28016,N_28236);
nor UO_1105 (O_1105,N_28305,N_28264);
nand UO_1106 (O_1106,N_28696,N_28313);
or UO_1107 (O_1107,N_29164,N_28729);
nand UO_1108 (O_1108,N_28202,N_28998);
or UO_1109 (O_1109,N_29888,N_29664);
and UO_1110 (O_1110,N_28595,N_28042);
nand UO_1111 (O_1111,N_29014,N_28346);
xnor UO_1112 (O_1112,N_28885,N_29324);
xor UO_1113 (O_1113,N_28006,N_28027);
nor UO_1114 (O_1114,N_28791,N_29930);
nor UO_1115 (O_1115,N_29239,N_29522);
nand UO_1116 (O_1116,N_29676,N_28731);
and UO_1117 (O_1117,N_29592,N_29265);
nand UO_1118 (O_1118,N_28085,N_28080);
xnor UO_1119 (O_1119,N_29434,N_29091);
xnor UO_1120 (O_1120,N_28322,N_28603);
or UO_1121 (O_1121,N_28580,N_28895);
and UO_1122 (O_1122,N_29580,N_29233);
xnor UO_1123 (O_1123,N_29769,N_29170);
nor UO_1124 (O_1124,N_29686,N_28169);
nor UO_1125 (O_1125,N_29396,N_29558);
or UO_1126 (O_1126,N_29530,N_29490);
or UO_1127 (O_1127,N_28544,N_29131);
nor UO_1128 (O_1128,N_29259,N_28712);
nand UO_1129 (O_1129,N_29770,N_29426);
or UO_1130 (O_1130,N_29250,N_28957);
and UO_1131 (O_1131,N_29463,N_28730);
nand UO_1132 (O_1132,N_28153,N_28091);
xor UO_1133 (O_1133,N_28168,N_28760);
xor UO_1134 (O_1134,N_28201,N_28693);
or UO_1135 (O_1135,N_29343,N_28340);
nand UO_1136 (O_1136,N_29769,N_29993);
and UO_1137 (O_1137,N_29138,N_29549);
nor UO_1138 (O_1138,N_28017,N_29643);
and UO_1139 (O_1139,N_28112,N_29083);
nand UO_1140 (O_1140,N_28623,N_28897);
nor UO_1141 (O_1141,N_28838,N_29277);
xor UO_1142 (O_1142,N_28892,N_29665);
nand UO_1143 (O_1143,N_28440,N_28272);
and UO_1144 (O_1144,N_29851,N_28602);
and UO_1145 (O_1145,N_28133,N_28739);
or UO_1146 (O_1146,N_29225,N_28674);
or UO_1147 (O_1147,N_28078,N_28629);
or UO_1148 (O_1148,N_29866,N_29638);
nor UO_1149 (O_1149,N_29892,N_28920);
nand UO_1150 (O_1150,N_29221,N_28326);
or UO_1151 (O_1151,N_28637,N_29624);
nor UO_1152 (O_1152,N_29701,N_28293);
nor UO_1153 (O_1153,N_29966,N_29249);
nor UO_1154 (O_1154,N_29480,N_28427);
and UO_1155 (O_1155,N_29381,N_29715);
or UO_1156 (O_1156,N_29500,N_29153);
or UO_1157 (O_1157,N_28616,N_29067);
xor UO_1158 (O_1158,N_28303,N_29122);
and UO_1159 (O_1159,N_29215,N_28680);
nand UO_1160 (O_1160,N_28178,N_29271);
or UO_1161 (O_1161,N_29631,N_29500);
and UO_1162 (O_1162,N_29150,N_29144);
nor UO_1163 (O_1163,N_29043,N_29271);
xnor UO_1164 (O_1164,N_28969,N_29562);
xnor UO_1165 (O_1165,N_29090,N_29745);
and UO_1166 (O_1166,N_28279,N_28012);
xor UO_1167 (O_1167,N_28070,N_29736);
and UO_1168 (O_1168,N_28884,N_28699);
nand UO_1169 (O_1169,N_29493,N_28355);
nor UO_1170 (O_1170,N_29343,N_29543);
nor UO_1171 (O_1171,N_28610,N_28444);
nor UO_1172 (O_1172,N_29411,N_29191);
or UO_1173 (O_1173,N_28703,N_29831);
xor UO_1174 (O_1174,N_29984,N_29719);
nand UO_1175 (O_1175,N_28452,N_28436);
xor UO_1176 (O_1176,N_29671,N_28900);
or UO_1177 (O_1177,N_29821,N_28388);
xor UO_1178 (O_1178,N_29846,N_28789);
nor UO_1179 (O_1179,N_29540,N_29025);
or UO_1180 (O_1180,N_29336,N_28094);
nand UO_1181 (O_1181,N_28954,N_28287);
and UO_1182 (O_1182,N_29920,N_28461);
and UO_1183 (O_1183,N_29047,N_28576);
xor UO_1184 (O_1184,N_28409,N_28020);
and UO_1185 (O_1185,N_28844,N_29045);
and UO_1186 (O_1186,N_29218,N_28687);
or UO_1187 (O_1187,N_28438,N_29079);
or UO_1188 (O_1188,N_28070,N_28432);
and UO_1189 (O_1189,N_29542,N_29773);
nor UO_1190 (O_1190,N_28134,N_28346);
and UO_1191 (O_1191,N_29916,N_28948);
nand UO_1192 (O_1192,N_29825,N_28979);
nand UO_1193 (O_1193,N_28756,N_29962);
nand UO_1194 (O_1194,N_28562,N_28426);
nor UO_1195 (O_1195,N_28986,N_28241);
xor UO_1196 (O_1196,N_28020,N_29345);
xor UO_1197 (O_1197,N_28114,N_29407);
nand UO_1198 (O_1198,N_29019,N_28440);
xnor UO_1199 (O_1199,N_29315,N_28825);
nand UO_1200 (O_1200,N_29539,N_28913);
nor UO_1201 (O_1201,N_29075,N_28690);
xnor UO_1202 (O_1202,N_29108,N_28094);
and UO_1203 (O_1203,N_29830,N_28821);
or UO_1204 (O_1204,N_28211,N_28262);
or UO_1205 (O_1205,N_28312,N_28555);
and UO_1206 (O_1206,N_29982,N_29332);
xor UO_1207 (O_1207,N_29128,N_29310);
xor UO_1208 (O_1208,N_29791,N_29569);
or UO_1209 (O_1209,N_29904,N_28313);
and UO_1210 (O_1210,N_28021,N_28292);
nor UO_1211 (O_1211,N_29622,N_29074);
and UO_1212 (O_1212,N_28745,N_28538);
nand UO_1213 (O_1213,N_29722,N_29892);
and UO_1214 (O_1214,N_29525,N_28815);
nor UO_1215 (O_1215,N_28458,N_28823);
nand UO_1216 (O_1216,N_28256,N_29496);
xor UO_1217 (O_1217,N_29044,N_29959);
xnor UO_1218 (O_1218,N_28403,N_29270);
nand UO_1219 (O_1219,N_29066,N_28969);
nand UO_1220 (O_1220,N_29027,N_28386);
or UO_1221 (O_1221,N_28226,N_29919);
or UO_1222 (O_1222,N_29517,N_29927);
and UO_1223 (O_1223,N_28602,N_28765);
xor UO_1224 (O_1224,N_29047,N_29023);
nor UO_1225 (O_1225,N_28266,N_28779);
nor UO_1226 (O_1226,N_28959,N_29824);
or UO_1227 (O_1227,N_28938,N_29675);
and UO_1228 (O_1228,N_29470,N_28186);
nor UO_1229 (O_1229,N_28743,N_28461);
nor UO_1230 (O_1230,N_29271,N_28815);
nor UO_1231 (O_1231,N_29124,N_29671);
and UO_1232 (O_1232,N_29866,N_29573);
nand UO_1233 (O_1233,N_29304,N_28370);
nand UO_1234 (O_1234,N_29835,N_29880);
or UO_1235 (O_1235,N_29871,N_28248);
nand UO_1236 (O_1236,N_29525,N_29738);
and UO_1237 (O_1237,N_28605,N_28730);
or UO_1238 (O_1238,N_29866,N_28505);
xor UO_1239 (O_1239,N_29515,N_29495);
xnor UO_1240 (O_1240,N_28702,N_29217);
or UO_1241 (O_1241,N_29060,N_29598);
xnor UO_1242 (O_1242,N_29110,N_28356);
nand UO_1243 (O_1243,N_29555,N_28983);
or UO_1244 (O_1244,N_29705,N_28370);
or UO_1245 (O_1245,N_28526,N_28777);
nor UO_1246 (O_1246,N_28358,N_29195);
nand UO_1247 (O_1247,N_29976,N_29237);
xor UO_1248 (O_1248,N_28756,N_28056);
nor UO_1249 (O_1249,N_29480,N_29483);
nor UO_1250 (O_1250,N_29410,N_29185);
and UO_1251 (O_1251,N_29864,N_29287);
and UO_1252 (O_1252,N_29132,N_29848);
and UO_1253 (O_1253,N_28691,N_29157);
and UO_1254 (O_1254,N_28785,N_28456);
xor UO_1255 (O_1255,N_29723,N_29305);
nand UO_1256 (O_1256,N_29968,N_29055);
nand UO_1257 (O_1257,N_28018,N_29452);
xnor UO_1258 (O_1258,N_29386,N_28901);
and UO_1259 (O_1259,N_29890,N_29314);
nand UO_1260 (O_1260,N_28142,N_28408);
nand UO_1261 (O_1261,N_29195,N_29837);
or UO_1262 (O_1262,N_28332,N_28326);
xor UO_1263 (O_1263,N_29192,N_28865);
or UO_1264 (O_1264,N_28998,N_29632);
or UO_1265 (O_1265,N_28997,N_28134);
xnor UO_1266 (O_1266,N_29110,N_29438);
or UO_1267 (O_1267,N_28475,N_29409);
nor UO_1268 (O_1268,N_29831,N_28312);
nand UO_1269 (O_1269,N_28141,N_29404);
nor UO_1270 (O_1270,N_29516,N_29407);
nor UO_1271 (O_1271,N_28558,N_29135);
and UO_1272 (O_1272,N_28946,N_28656);
and UO_1273 (O_1273,N_28709,N_29563);
and UO_1274 (O_1274,N_28140,N_29618);
nand UO_1275 (O_1275,N_29227,N_28440);
and UO_1276 (O_1276,N_28380,N_29081);
and UO_1277 (O_1277,N_29315,N_28827);
nor UO_1278 (O_1278,N_29844,N_28602);
or UO_1279 (O_1279,N_29112,N_29523);
nor UO_1280 (O_1280,N_29356,N_29969);
and UO_1281 (O_1281,N_29009,N_29581);
nor UO_1282 (O_1282,N_28782,N_28612);
nor UO_1283 (O_1283,N_29994,N_28166);
or UO_1284 (O_1284,N_28649,N_29791);
xor UO_1285 (O_1285,N_29364,N_29577);
or UO_1286 (O_1286,N_28727,N_28653);
and UO_1287 (O_1287,N_28832,N_28283);
or UO_1288 (O_1288,N_28573,N_28815);
and UO_1289 (O_1289,N_29575,N_28068);
and UO_1290 (O_1290,N_29759,N_28523);
or UO_1291 (O_1291,N_29620,N_28754);
and UO_1292 (O_1292,N_28721,N_29994);
and UO_1293 (O_1293,N_28088,N_29231);
nor UO_1294 (O_1294,N_29851,N_29917);
xor UO_1295 (O_1295,N_29129,N_29395);
xor UO_1296 (O_1296,N_29957,N_29419);
nor UO_1297 (O_1297,N_29467,N_29530);
nor UO_1298 (O_1298,N_28342,N_28272);
xnor UO_1299 (O_1299,N_28796,N_28098);
or UO_1300 (O_1300,N_29295,N_29959);
and UO_1301 (O_1301,N_29243,N_29475);
nor UO_1302 (O_1302,N_28202,N_28877);
xor UO_1303 (O_1303,N_28778,N_29198);
or UO_1304 (O_1304,N_29203,N_28413);
nor UO_1305 (O_1305,N_28247,N_28236);
xnor UO_1306 (O_1306,N_29721,N_29321);
nand UO_1307 (O_1307,N_28876,N_28914);
or UO_1308 (O_1308,N_28245,N_28082);
and UO_1309 (O_1309,N_29109,N_28448);
and UO_1310 (O_1310,N_28562,N_29058);
xnor UO_1311 (O_1311,N_28291,N_29431);
and UO_1312 (O_1312,N_29957,N_28782);
or UO_1313 (O_1313,N_29474,N_28689);
or UO_1314 (O_1314,N_29683,N_29255);
nor UO_1315 (O_1315,N_28224,N_28310);
nor UO_1316 (O_1316,N_28172,N_28530);
and UO_1317 (O_1317,N_28036,N_29095);
nand UO_1318 (O_1318,N_29088,N_28961);
nor UO_1319 (O_1319,N_28494,N_29995);
nor UO_1320 (O_1320,N_28511,N_29357);
xor UO_1321 (O_1321,N_29741,N_28626);
or UO_1322 (O_1322,N_28992,N_29415);
and UO_1323 (O_1323,N_29645,N_28052);
and UO_1324 (O_1324,N_28548,N_29826);
nand UO_1325 (O_1325,N_28031,N_29343);
or UO_1326 (O_1326,N_28807,N_28411);
nor UO_1327 (O_1327,N_28674,N_28964);
or UO_1328 (O_1328,N_28105,N_28611);
xnor UO_1329 (O_1329,N_29585,N_29565);
and UO_1330 (O_1330,N_29079,N_28503);
xor UO_1331 (O_1331,N_29904,N_28413);
nor UO_1332 (O_1332,N_29243,N_29085);
xor UO_1333 (O_1333,N_28793,N_28199);
and UO_1334 (O_1334,N_29123,N_28933);
xnor UO_1335 (O_1335,N_29523,N_28981);
or UO_1336 (O_1336,N_28909,N_28898);
or UO_1337 (O_1337,N_28294,N_28264);
and UO_1338 (O_1338,N_29986,N_28679);
xor UO_1339 (O_1339,N_28040,N_29571);
nor UO_1340 (O_1340,N_29921,N_29781);
nor UO_1341 (O_1341,N_28248,N_29856);
and UO_1342 (O_1342,N_29540,N_29960);
nor UO_1343 (O_1343,N_28796,N_29358);
xor UO_1344 (O_1344,N_29655,N_29129);
nand UO_1345 (O_1345,N_29449,N_29783);
nor UO_1346 (O_1346,N_28377,N_29506);
and UO_1347 (O_1347,N_29692,N_28148);
or UO_1348 (O_1348,N_29270,N_29225);
xnor UO_1349 (O_1349,N_29916,N_29491);
or UO_1350 (O_1350,N_28692,N_29027);
or UO_1351 (O_1351,N_29154,N_28923);
nand UO_1352 (O_1352,N_28709,N_28119);
or UO_1353 (O_1353,N_29665,N_28943);
nand UO_1354 (O_1354,N_28061,N_29028);
or UO_1355 (O_1355,N_29593,N_28380);
nand UO_1356 (O_1356,N_28785,N_28633);
or UO_1357 (O_1357,N_29277,N_28375);
and UO_1358 (O_1358,N_29588,N_28672);
xor UO_1359 (O_1359,N_28867,N_29310);
or UO_1360 (O_1360,N_29037,N_29736);
xor UO_1361 (O_1361,N_29301,N_28302);
nor UO_1362 (O_1362,N_28381,N_29668);
nand UO_1363 (O_1363,N_28120,N_28391);
xnor UO_1364 (O_1364,N_28235,N_28310);
nand UO_1365 (O_1365,N_29511,N_28097);
or UO_1366 (O_1366,N_29195,N_28219);
or UO_1367 (O_1367,N_29098,N_28406);
or UO_1368 (O_1368,N_29699,N_29758);
nand UO_1369 (O_1369,N_29010,N_29523);
xnor UO_1370 (O_1370,N_28179,N_29040);
nor UO_1371 (O_1371,N_29857,N_29253);
nand UO_1372 (O_1372,N_28300,N_28622);
and UO_1373 (O_1373,N_28641,N_28982);
or UO_1374 (O_1374,N_29047,N_28040);
nand UO_1375 (O_1375,N_29074,N_29001);
and UO_1376 (O_1376,N_28682,N_29420);
xor UO_1377 (O_1377,N_28139,N_28751);
or UO_1378 (O_1378,N_28781,N_29266);
or UO_1379 (O_1379,N_28094,N_29894);
nand UO_1380 (O_1380,N_28195,N_28774);
xor UO_1381 (O_1381,N_29691,N_28884);
nor UO_1382 (O_1382,N_29429,N_29401);
nor UO_1383 (O_1383,N_28165,N_28009);
and UO_1384 (O_1384,N_28113,N_29482);
nand UO_1385 (O_1385,N_28819,N_28260);
or UO_1386 (O_1386,N_28803,N_28694);
and UO_1387 (O_1387,N_29916,N_28760);
and UO_1388 (O_1388,N_29525,N_28888);
or UO_1389 (O_1389,N_28999,N_28206);
or UO_1390 (O_1390,N_29483,N_29606);
xor UO_1391 (O_1391,N_29285,N_28031);
nand UO_1392 (O_1392,N_29977,N_28333);
xnor UO_1393 (O_1393,N_29015,N_29265);
xnor UO_1394 (O_1394,N_29120,N_28609);
or UO_1395 (O_1395,N_29354,N_29345);
and UO_1396 (O_1396,N_28111,N_29498);
xnor UO_1397 (O_1397,N_29803,N_29147);
nor UO_1398 (O_1398,N_29327,N_28684);
and UO_1399 (O_1399,N_28082,N_28870);
nand UO_1400 (O_1400,N_28492,N_28102);
nand UO_1401 (O_1401,N_29212,N_29520);
or UO_1402 (O_1402,N_28375,N_29138);
and UO_1403 (O_1403,N_28067,N_29349);
or UO_1404 (O_1404,N_28158,N_29683);
nor UO_1405 (O_1405,N_29059,N_28898);
nor UO_1406 (O_1406,N_29065,N_28492);
or UO_1407 (O_1407,N_28748,N_28499);
xnor UO_1408 (O_1408,N_28085,N_28409);
and UO_1409 (O_1409,N_29224,N_29747);
nand UO_1410 (O_1410,N_28322,N_29269);
xor UO_1411 (O_1411,N_28496,N_28227);
nor UO_1412 (O_1412,N_28667,N_29259);
xnor UO_1413 (O_1413,N_29156,N_29693);
xnor UO_1414 (O_1414,N_29172,N_29287);
or UO_1415 (O_1415,N_28869,N_28769);
nand UO_1416 (O_1416,N_29471,N_29498);
and UO_1417 (O_1417,N_28239,N_28246);
nor UO_1418 (O_1418,N_29379,N_29103);
nor UO_1419 (O_1419,N_29425,N_29068);
and UO_1420 (O_1420,N_28388,N_28414);
or UO_1421 (O_1421,N_29668,N_29401);
xor UO_1422 (O_1422,N_28477,N_28409);
nor UO_1423 (O_1423,N_29239,N_29126);
or UO_1424 (O_1424,N_29923,N_29085);
xor UO_1425 (O_1425,N_28726,N_28707);
nor UO_1426 (O_1426,N_28732,N_29363);
nand UO_1427 (O_1427,N_29147,N_29989);
nor UO_1428 (O_1428,N_28412,N_28913);
or UO_1429 (O_1429,N_29814,N_28144);
xor UO_1430 (O_1430,N_29523,N_29133);
xor UO_1431 (O_1431,N_28415,N_29397);
xnor UO_1432 (O_1432,N_28331,N_28225);
xor UO_1433 (O_1433,N_28993,N_29411);
xor UO_1434 (O_1434,N_29174,N_28352);
and UO_1435 (O_1435,N_28568,N_28675);
and UO_1436 (O_1436,N_28288,N_29499);
and UO_1437 (O_1437,N_29681,N_28127);
nand UO_1438 (O_1438,N_29990,N_28790);
or UO_1439 (O_1439,N_29044,N_28586);
nor UO_1440 (O_1440,N_29164,N_29419);
xnor UO_1441 (O_1441,N_29851,N_29920);
and UO_1442 (O_1442,N_28629,N_29935);
and UO_1443 (O_1443,N_28144,N_29070);
or UO_1444 (O_1444,N_28242,N_29501);
nand UO_1445 (O_1445,N_29929,N_28729);
nor UO_1446 (O_1446,N_29010,N_29422);
nand UO_1447 (O_1447,N_29531,N_28085);
nand UO_1448 (O_1448,N_28376,N_29899);
nor UO_1449 (O_1449,N_28350,N_28968);
or UO_1450 (O_1450,N_29966,N_28966);
or UO_1451 (O_1451,N_28894,N_29369);
nor UO_1452 (O_1452,N_29340,N_28171);
nand UO_1453 (O_1453,N_29734,N_29218);
nand UO_1454 (O_1454,N_29837,N_28556);
nor UO_1455 (O_1455,N_29189,N_29791);
and UO_1456 (O_1456,N_29890,N_28976);
nand UO_1457 (O_1457,N_28553,N_29814);
nor UO_1458 (O_1458,N_28382,N_29535);
or UO_1459 (O_1459,N_28996,N_29128);
and UO_1460 (O_1460,N_29511,N_28891);
nand UO_1461 (O_1461,N_28577,N_28202);
xor UO_1462 (O_1462,N_28809,N_29769);
xor UO_1463 (O_1463,N_29274,N_29578);
nand UO_1464 (O_1464,N_28264,N_29933);
nor UO_1465 (O_1465,N_29066,N_28755);
nor UO_1466 (O_1466,N_28619,N_28765);
or UO_1467 (O_1467,N_29255,N_29424);
and UO_1468 (O_1468,N_29394,N_29074);
nand UO_1469 (O_1469,N_28077,N_29419);
nor UO_1470 (O_1470,N_28499,N_28193);
nand UO_1471 (O_1471,N_29603,N_28582);
xnor UO_1472 (O_1472,N_29255,N_29904);
nand UO_1473 (O_1473,N_29798,N_28168);
and UO_1474 (O_1474,N_28134,N_29026);
nand UO_1475 (O_1475,N_29177,N_28886);
xnor UO_1476 (O_1476,N_29099,N_29004);
and UO_1477 (O_1477,N_28927,N_28195);
nor UO_1478 (O_1478,N_29954,N_28054);
nand UO_1479 (O_1479,N_29496,N_29121);
or UO_1480 (O_1480,N_29807,N_28002);
and UO_1481 (O_1481,N_29757,N_28544);
and UO_1482 (O_1482,N_28424,N_28241);
or UO_1483 (O_1483,N_28133,N_29103);
nand UO_1484 (O_1484,N_29549,N_28168);
xor UO_1485 (O_1485,N_28221,N_29900);
and UO_1486 (O_1486,N_29276,N_28842);
xor UO_1487 (O_1487,N_28655,N_28313);
nand UO_1488 (O_1488,N_28303,N_29190);
or UO_1489 (O_1489,N_29373,N_29975);
or UO_1490 (O_1490,N_28451,N_29318);
nor UO_1491 (O_1491,N_28535,N_29264);
or UO_1492 (O_1492,N_29600,N_28899);
nor UO_1493 (O_1493,N_28260,N_29677);
xor UO_1494 (O_1494,N_29125,N_28041);
nand UO_1495 (O_1495,N_28348,N_29789);
nor UO_1496 (O_1496,N_29406,N_29786);
xor UO_1497 (O_1497,N_28231,N_29738);
nand UO_1498 (O_1498,N_29471,N_29713);
or UO_1499 (O_1499,N_28714,N_28796);
or UO_1500 (O_1500,N_28174,N_29246);
nand UO_1501 (O_1501,N_29671,N_29393);
or UO_1502 (O_1502,N_29353,N_28734);
or UO_1503 (O_1503,N_28378,N_28144);
or UO_1504 (O_1504,N_29402,N_28717);
and UO_1505 (O_1505,N_28994,N_28904);
nand UO_1506 (O_1506,N_28197,N_29333);
nor UO_1507 (O_1507,N_29719,N_29214);
nand UO_1508 (O_1508,N_28705,N_28389);
and UO_1509 (O_1509,N_28360,N_28674);
nand UO_1510 (O_1510,N_28694,N_28317);
or UO_1511 (O_1511,N_29862,N_29474);
and UO_1512 (O_1512,N_28109,N_28782);
and UO_1513 (O_1513,N_29131,N_28036);
nor UO_1514 (O_1514,N_29206,N_29412);
xor UO_1515 (O_1515,N_29477,N_29552);
and UO_1516 (O_1516,N_28785,N_28030);
nor UO_1517 (O_1517,N_28162,N_29907);
nor UO_1518 (O_1518,N_29847,N_28968);
and UO_1519 (O_1519,N_29905,N_29664);
and UO_1520 (O_1520,N_29224,N_29778);
nor UO_1521 (O_1521,N_29350,N_29762);
xor UO_1522 (O_1522,N_28453,N_29779);
and UO_1523 (O_1523,N_29045,N_29510);
nand UO_1524 (O_1524,N_29766,N_29598);
nand UO_1525 (O_1525,N_28282,N_28296);
nand UO_1526 (O_1526,N_29436,N_28962);
nand UO_1527 (O_1527,N_29116,N_28970);
or UO_1528 (O_1528,N_28798,N_28872);
nor UO_1529 (O_1529,N_28090,N_29277);
xnor UO_1530 (O_1530,N_28675,N_28161);
nor UO_1531 (O_1531,N_29602,N_28352);
xor UO_1532 (O_1532,N_28701,N_28214);
and UO_1533 (O_1533,N_28265,N_28345);
nand UO_1534 (O_1534,N_29875,N_29747);
or UO_1535 (O_1535,N_29120,N_28479);
nand UO_1536 (O_1536,N_28916,N_28352);
or UO_1537 (O_1537,N_28801,N_29527);
nand UO_1538 (O_1538,N_29502,N_28365);
and UO_1539 (O_1539,N_29913,N_29835);
or UO_1540 (O_1540,N_28481,N_28129);
nand UO_1541 (O_1541,N_29328,N_28759);
nor UO_1542 (O_1542,N_29014,N_29616);
nor UO_1543 (O_1543,N_29885,N_29345);
nor UO_1544 (O_1544,N_29479,N_29273);
xnor UO_1545 (O_1545,N_28391,N_29747);
or UO_1546 (O_1546,N_28296,N_29843);
and UO_1547 (O_1547,N_28741,N_28653);
nor UO_1548 (O_1548,N_29962,N_28213);
or UO_1549 (O_1549,N_28721,N_29076);
xor UO_1550 (O_1550,N_29311,N_28750);
nand UO_1551 (O_1551,N_28291,N_28309);
and UO_1552 (O_1552,N_29768,N_28388);
and UO_1553 (O_1553,N_28069,N_28536);
xor UO_1554 (O_1554,N_28780,N_28121);
nor UO_1555 (O_1555,N_28775,N_29349);
and UO_1556 (O_1556,N_29873,N_29359);
nor UO_1557 (O_1557,N_29914,N_29255);
nand UO_1558 (O_1558,N_29784,N_29632);
nand UO_1559 (O_1559,N_29869,N_29028);
and UO_1560 (O_1560,N_28657,N_29556);
or UO_1561 (O_1561,N_29542,N_28936);
nor UO_1562 (O_1562,N_29082,N_29805);
xor UO_1563 (O_1563,N_29783,N_29807);
or UO_1564 (O_1564,N_28182,N_28472);
xnor UO_1565 (O_1565,N_29182,N_28514);
nand UO_1566 (O_1566,N_28176,N_29328);
or UO_1567 (O_1567,N_29572,N_29272);
and UO_1568 (O_1568,N_29344,N_29160);
or UO_1569 (O_1569,N_29161,N_28332);
or UO_1570 (O_1570,N_29472,N_28033);
or UO_1571 (O_1571,N_29388,N_28622);
nor UO_1572 (O_1572,N_28787,N_28372);
nor UO_1573 (O_1573,N_28806,N_29464);
nor UO_1574 (O_1574,N_28731,N_28787);
and UO_1575 (O_1575,N_29711,N_29910);
nand UO_1576 (O_1576,N_29604,N_28453);
nor UO_1577 (O_1577,N_29112,N_28930);
nand UO_1578 (O_1578,N_29907,N_29260);
nor UO_1579 (O_1579,N_29208,N_28475);
nor UO_1580 (O_1580,N_28114,N_28229);
and UO_1581 (O_1581,N_29858,N_29537);
and UO_1582 (O_1582,N_28078,N_28270);
and UO_1583 (O_1583,N_29513,N_29323);
nor UO_1584 (O_1584,N_28737,N_28119);
nor UO_1585 (O_1585,N_28112,N_28167);
or UO_1586 (O_1586,N_28329,N_29803);
or UO_1587 (O_1587,N_28190,N_28488);
xor UO_1588 (O_1588,N_28900,N_28711);
or UO_1589 (O_1589,N_28974,N_29572);
xor UO_1590 (O_1590,N_29314,N_29052);
or UO_1591 (O_1591,N_29094,N_29332);
nand UO_1592 (O_1592,N_29090,N_28108);
nand UO_1593 (O_1593,N_28195,N_29682);
nor UO_1594 (O_1594,N_29036,N_29922);
nor UO_1595 (O_1595,N_28137,N_29898);
or UO_1596 (O_1596,N_29138,N_29651);
xnor UO_1597 (O_1597,N_28694,N_29525);
nand UO_1598 (O_1598,N_28434,N_28359);
xor UO_1599 (O_1599,N_29389,N_29553);
xor UO_1600 (O_1600,N_29554,N_28401);
or UO_1601 (O_1601,N_28613,N_28583);
xnor UO_1602 (O_1602,N_28541,N_29714);
xnor UO_1603 (O_1603,N_28942,N_28604);
nor UO_1604 (O_1604,N_29184,N_29079);
nand UO_1605 (O_1605,N_29837,N_29498);
or UO_1606 (O_1606,N_29761,N_29840);
and UO_1607 (O_1607,N_28264,N_28450);
xor UO_1608 (O_1608,N_28559,N_29755);
nand UO_1609 (O_1609,N_29312,N_29779);
xor UO_1610 (O_1610,N_28566,N_28666);
and UO_1611 (O_1611,N_28394,N_28761);
nor UO_1612 (O_1612,N_29638,N_28959);
and UO_1613 (O_1613,N_28745,N_28078);
and UO_1614 (O_1614,N_29419,N_29733);
or UO_1615 (O_1615,N_29295,N_28164);
or UO_1616 (O_1616,N_28922,N_29443);
and UO_1617 (O_1617,N_28244,N_28837);
xnor UO_1618 (O_1618,N_28070,N_29668);
and UO_1619 (O_1619,N_29329,N_28223);
nor UO_1620 (O_1620,N_29930,N_28615);
nor UO_1621 (O_1621,N_29455,N_28316);
xnor UO_1622 (O_1622,N_29588,N_28514);
nor UO_1623 (O_1623,N_29048,N_28637);
or UO_1624 (O_1624,N_29392,N_28088);
and UO_1625 (O_1625,N_28822,N_29172);
xnor UO_1626 (O_1626,N_28365,N_28074);
nand UO_1627 (O_1627,N_28623,N_28451);
and UO_1628 (O_1628,N_28504,N_28063);
nor UO_1629 (O_1629,N_29496,N_29806);
or UO_1630 (O_1630,N_28924,N_29940);
or UO_1631 (O_1631,N_29040,N_28460);
nand UO_1632 (O_1632,N_29037,N_29582);
xnor UO_1633 (O_1633,N_29027,N_28265);
or UO_1634 (O_1634,N_29618,N_28812);
xnor UO_1635 (O_1635,N_29656,N_29267);
or UO_1636 (O_1636,N_29270,N_29689);
or UO_1637 (O_1637,N_28357,N_29384);
nand UO_1638 (O_1638,N_29290,N_29034);
xnor UO_1639 (O_1639,N_28613,N_29109);
nor UO_1640 (O_1640,N_29698,N_29940);
nand UO_1641 (O_1641,N_29912,N_29117);
and UO_1642 (O_1642,N_28898,N_28686);
nand UO_1643 (O_1643,N_29075,N_29586);
nor UO_1644 (O_1644,N_29873,N_28916);
xnor UO_1645 (O_1645,N_28768,N_29397);
nand UO_1646 (O_1646,N_28602,N_28997);
nor UO_1647 (O_1647,N_29875,N_28295);
and UO_1648 (O_1648,N_28832,N_28183);
nand UO_1649 (O_1649,N_29828,N_29618);
and UO_1650 (O_1650,N_29798,N_29843);
nor UO_1651 (O_1651,N_28128,N_29950);
nor UO_1652 (O_1652,N_29799,N_28591);
nor UO_1653 (O_1653,N_29863,N_28063);
nor UO_1654 (O_1654,N_28973,N_28851);
nand UO_1655 (O_1655,N_29287,N_29619);
xor UO_1656 (O_1656,N_28791,N_28570);
nand UO_1657 (O_1657,N_29266,N_28934);
xor UO_1658 (O_1658,N_28676,N_29710);
or UO_1659 (O_1659,N_28575,N_28933);
xor UO_1660 (O_1660,N_28212,N_29476);
xnor UO_1661 (O_1661,N_29364,N_28513);
and UO_1662 (O_1662,N_28646,N_28724);
nand UO_1663 (O_1663,N_29151,N_28948);
xor UO_1664 (O_1664,N_29948,N_28905);
nand UO_1665 (O_1665,N_28939,N_29062);
xor UO_1666 (O_1666,N_29146,N_29006);
nand UO_1667 (O_1667,N_28299,N_28621);
nand UO_1668 (O_1668,N_29761,N_29114);
xnor UO_1669 (O_1669,N_28363,N_28664);
nor UO_1670 (O_1670,N_28830,N_29418);
nand UO_1671 (O_1671,N_29260,N_29075);
xor UO_1672 (O_1672,N_28325,N_29089);
xor UO_1673 (O_1673,N_28339,N_29209);
and UO_1674 (O_1674,N_28519,N_29028);
or UO_1675 (O_1675,N_28565,N_29331);
nand UO_1676 (O_1676,N_28555,N_28455);
and UO_1677 (O_1677,N_28053,N_28121);
or UO_1678 (O_1678,N_28659,N_28406);
xor UO_1679 (O_1679,N_29611,N_28062);
nand UO_1680 (O_1680,N_29727,N_28501);
and UO_1681 (O_1681,N_28398,N_29044);
or UO_1682 (O_1682,N_29291,N_28384);
nor UO_1683 (O_1683,N_28074,N_28732);
nand UO_1684 (O_1684,N_29210,N_29152);
xnor UO_1685 (O_1685,N_29594,N_29491);
nor UO_1686 (O_1686,N_29383,N_29524);
nand UO_1687 (O_1687,N_29383,N_28201);
and UO_1688 (O_1688,N_28119,N_29849);
nand UO_1689 (O_1689,N_28434,N_29463);
or UO_1690 (O_1690,N_29156,N_28641);
xnor UO_1691 (O_1691,N_29941,N_29526);
nor UO_1692 (O_1692,N_28364,N_28840);
nand UO_1693 (O_1693,N_29554,N_28799);
xor UO_1694 (O_1694,N_28726,N_28427);
or UO_1695 (O_1695,N_28005,N_28600);
nor UO_1696 (O_1696,N_28523,N_29693);
or UO_1697 (O_1697,N_28785,N_29926);
xnor UO_1698 (O_1698,N_29921,N_29630);
nand UO_1699 (O_1699,N_28245,N_28167);
or UO_1700 (O_1700,N_29042,N_29239);
or UO_1701 (O_1701,N_29316,N_29452);
and UO_1702 (O_1702,N_29006,N_28901);
nand UO_1703 (O_1703,N_28154,N_28418);
or UO_1704 (O_1704,N_28067,N_28075);
or UO_1705 (O_1705,N_28461,N_29552);
or UO_1706 (O_1706,N_29940,N_29325);
nand UO_1707 (O_1707,N_28913,N_28739);
and UO_1708 (O_1708,N_28998,N_29325);
nor UO_1709 (O_1709,N_28711,N_28939);
and UO_1710 (O_1710,N_28348,N_28265);
xnor UO_1711 (O_1711,N_28916,N_29733);
or UO_1712 (O_1712,N_29051,N_29443);
nand UO_1713 (O_1713,N_29328,N_28785);
xor UO_1714 (O_1714,N_29240,N_29295);
or UO_1715 (O_1715,N_28049,N_28306);
and UO_1716 (O_1716,N_29299,N_28147);
nand UO_1717 (O_1717,N_29008,N_29704);
nor UO_1718 (O_1718,N_29081,N_29593);
xnor UO_1719 (O_1719,N_28235,N_29442);
xnor UO_1720 (O_1720,N_28470,N_29269);
xnor UO_1721 (O_1721,N_29582,N_29810);
or UO_1722 (O_1722,N_28917,N_29392);
xor UO_1723 (O_1723,N_28451,N_29917);
xnor UO_1724 (O_1724,N_28718,N_28856);
nand UO_1725 (O_1725,N_29596,N_28918);
nor UO_1726 (O_1726,N_29167,N_28661);
and UO_1727 (O_1727,N_29196,N_29345);
or UO_1728 (O_1728,N_28490,N_29487);
xnor UO_1729 (O_1729,N_28135,N_29149);
nand UO_1730 (O_1730,N_28891,N_29427);
nand UO_1731 (O_1731,N_29410,N_28188);
and UO_1732 (O_1732,N_28810,N_28527);
and UO_1733 (O_1733,N_29395,N_28254);
or UO_1734 (O_1734,N_29667,N_28111);
and UO_1735 (O_1735,N_28853,N_28773);
xnor UO_1736 (O_1736,N_29059,N_28718);
and UO_1737 (O_1737,N_28299,N_28294);
or UO_1738 (O_1738,N_29130,N_29346);
nand UO_1739 (O_1739,N_28160,N_29010);
nor UO_1740 (O_1740,N_28454,N_29463);
nor UO_1741 (O_1741,N_29721,N_28814);
xor UO_1742 (O_1742,N_29133,N_29874);
xor UO_1743 (O_1743,N_28479,N_29923);
or UO_1744 (O_1744,N_29939,N_29828);
xnor UO_1745 (O_1745,N_29464,N_28553);
nand UO_1746 (O_1746,N_28044,N_28990);
or UO_1747 (O_1747,N_29651,N_28176);
or UO_1748 (O_1748,N_28652,N_28037);
xnor UO_1749 (O_1749,N_28370,N_29070);
xor UO_1750 (O_1750,N_28298,N_29509);
and UO_1751 (O_1751,N_29032,N_29834);
and UO_1752 (O_1752,N_28277,N_29316);
or UO_1753 (O_1753,N_28730,N_29487);
xor UO_1754 (O_1754,N_28665,N_28801);
nand UO_1755 (O_1755,N_28226,N_29635);
nor UO_1756 (O_1756,N_28768,N_28386);
xor UO_1757 (O_1757,N_29902,N_28528);
and UO_1758 (O_1758,N_28539,N_28260);
nand UO_1759 (O_1759,N_29332,N_28314);
and UO_1760 (O_1760,N_29787,N_28207);
nand UO_1761 (O_1761,N_28764,N_29327);
and UO_1762 (O_1762,N_28761,N_29123);
or UO_1763 (O_1763,N_28470,N_28731);
nand UO_1764 (O_1764,N_29054,N_28994);
and UO_1765 (O_1765,N_28637,N_29595);
and UO_1766 (O_1766,N_28022,N_28051);
or UO_1767 (O_1767,N_29990,N_28978);
nor UO_1768 (O_1768,N_28283,N_29993);
nand UO_1769 (O_1769,N_29311,N_29556);
and UO_1770 (O_1770,N_28841,N_29273);
nand UO_1771 (O_1771,N_29924,N_28670);
nand UO_1772 (O_1772,N_28784,N_29382);
and UO_1773 (O_1773,N_28415,N_28365);
xnor UO_1774 (O_1774,N_29924,N_28787);
and UO_1775 (O_1775,N_28968,N_28576);
nand UO_1776 (O_1776,N_28386,N_28985);
xnor UO_1777 (O_1777,N_29545,N_29779);
nor UO_1778 (O_1778,N_28322,N_29483);
xnor UO_1779 (O_1779,N_29206,N_28220);
or UO_1780 (O_1780,N_29701,N_28498);
xnor UO_1781 (O_1781,N_28232,N_29433);
and UO_1782 (O_1782,N_29633,N_28232);
xnor UO_1783 (O_1783,N_29060,N_29243);
xor UO_1784 (O_1784,N_29398,N_29395);
xnor UO_1785 (O_1785,N_29294,N_28208);
and UO_1786 (O_1786,N_29665,N_29596);
or UO_1787 (O_1787,N_29593,N_29882);
and UO_1788 (O_1788,N_29619,N_29034);
or UO_1789 (O_1789,N_29846,N_29949);
nor UO_1790 (O_1790,N_29982,N_29652);
nor UO_1791 (O_1791,N_29200,N_29734);
and UO_1792 (O_1792,N_28288,N_29110);
and UO_1793 (O_1793,N_29646,N_29117);
and UO_1794 (O_1794,N_28756,N_28596);
or UO_1795 (O_1795,N_29709,N_29295);
xor UO_1796 (O_1796,N_29417,N_28509);
or UO_1797 (O_1797,N_28776,N_29407);
and UO_1798 (O_1798,N_29961,N_29507);
xnor UO_1799 (O_1799,N_29776,N_28089);
or UO_1800 (O_1800,N_29555,N_29203);
nand UO_1801 (O_1801,N_28081,N_28046);
xnor UO_1802 (O_1802,N_29789,N_28320);
or UO_1803 (O_1803,N_29660,N_28939);
nor UO_1804 (O_1804,N_28242,N_29942);
xnor UO_1805 (O_1805,N_29861,N_28451);
and UO_1806 (O_1806,N_29129,N_29565);
nand UO_1807 (O_1807,N_29490,N_29932);
and UO_1808 (O_1808,N_29739,N_29331);
or UO_1809 (O_1809,N_28351,N_28708);
nand UO_1810 (O_1810,N_29250,N_28072);
nand UO_1811 (O_1811,N_29844,N_28250);
xnor UO_1812 (O_1812,N_29198,N_28313);
or UO_1813 (O_1813,N_29882,N_28281);
or UO_1814 (O_1814,N_29961,N_29800);
xnor UO_1815 (O_1815,N_28039,N_28457);
xor UO_1816 (O_1816,N_28554,N_28412);
xor UO_1817 (O_1817,N_28884,N_28777);
and UO_1818 (O_1818,N_29476,N_29503);
and UO_1819 (O_1819,N_28798,N_29736);
nor UO_1820 (O_1820,N_28198,N_29625);
xnor UO_1821 (O_1821,N_29987,N_29984);
xnor UO_1822 (O_1822,N_29537,N_29294);
nand UO_1823 (O_1823,N_29453,N_29318);
nor UO_1824 (O_1824,N_28202,N_28736);
or UO_1825 (O_1825,N_28339,N_29840);
nand UO_1826 (O_1826,N_29477,N_28135);
and UO_1827 (O_1827,N_28931,N_29794);
xor UO_1828 (O_1828,N_28387,N_28821);
nor UO_1829 (O_1829,N_29050,N_28454);
and UO_1830 (O_1830,N_28431,N_29002);
and UO_1831 (O_1831,N_29858,N_28829);
or UO_1832 (O_1832,N_29978,N_28072);
and UO_1833 (O_1833,N_28253,N_29690);
and UO_1834 (O_1834,N_28603,N_28999);
and UO_1835 (O_1835,N_29200,N_29708);
nand UO_1836 (O_1836,N_28752,N_28724);
or UO_1837 (O_1837,N_28149,N_29097);
nand UO_1838 (O_1838,N_29487,N_29825);
xnor UO_1839 (O_1839,N_28961,N_28426);
xnor UO_1840 (O_1840,N_28727,N_28097);
or UO_1841 (O_1841,N_29417,N_29030);
nor UO_1842 (O_1842,N_29799,N_28579);
nand UO_1843 (O_1843,N_29676,N_28284);
and UO_1844 (O_1844,N_28937,N_28734);
nand UO_1845 (O_1845,N_29761,N_29034);
and UO_1846 (O_1846,N_29221,N_28384);
xor UO_1847 (O_1847,N_29285,N_29138);
and UO_1848 (O_1848,N_29376,N_29594);
xor UO_1849 (O_1849,N_28983,N_29017);
or UO_1850 (O_1850,N_28713,N_28720);
xnor UO_1851 (O_1851,N_29743,N_29514);
nor UO_1852 (O_1852,N_28922,N_29736);
nand UO_1853 (O_1853,N_28711,N_28829);
nor UO_1854 (O_1854,N_29727,N_28525);
and UO_1855 (O_1855,N_28666,N_28587);
or UO_1856 (O_1856,N_29795,N_29545);
or UO_1857 (O_1857,N_28064,N_28386);
or UO_1858 (O_1858,N_28993,N_28440);
or UO_1859 (O_1859,N_28066,N_29416);
nand UO_1860 (O_1860,N_29620,N_28463);
or UO_1861 (O_1861,N_28235,N_29032);
or UO_1862 (O_1862,N_28097,N_28113);
nand UO_1863 (O_1863,N_28321,N_29676);
nor UO_1864 (O_1864,N_28570,N_28847);
nand UO_1865 (O_1865,N_28360,N_29581);
nand UO_1866 (O_1866,N_28028,N_29627);
and UO_1867 (O_1867,N_28561,N_29007);
or UO_1868 (O_1868,N_29297,N_28627);
or UO_1869 (O_1869,N_29863,N_29418);
xnor UO_1870 (O_1870,N_28988,N_29202);
xor UO_1871 (O_1871,N_29174,N_28833);
xnor UO_1872 (O_1872,N_28119,N_29008);
and UO_1873 (O_1873,N_28471,N_28281);
and UO_1874 (O_1874,N_28387,N_28094);
nand UO_1875 (O_1875,N_28836,N_28789);
nor UO_1876 (O_1876,N_28033,N_28565);
and UO_1877 (O_1877,N_29405,N_28586);
and UO_1878 (O_1878,N_28891,N_29793);
or UO_1879 (O_1879,N_29162,N_29966);
and UO_1880 (O_1880,N_29652,N_28863);
nand UO_1881 (O_1881,N_28542,N_29271);
or UO_1882 (O_1882,N_28785,N_29577);
nor UO_1883 (O_1883,N_28031,N_28528);
or UO_1884 (O_1884,N_29721,N_29302);
and UO_1885 (O_1885,N_28591,N_28285);
xor UO_1886 (O_1886,N_29520,N_28574);
or UO_1887 (O_1887,N_28959,N_28566);
nand UO_1888 (O_1888,N_28795,N_28099);
nor UO_1889 (O_1889,N_28294,N_29367);
nor UO_1890 (O_1890,N_28229,N_29387);
nand UO_1891 (O_1891,N_29782,N_28158);
nor UO_1892 (O_1892,N_29978,N_29700);
nand UO_1893 (O_1893,N_28434,N_28307);
nor UO_1894 (O_1894,N_28319,N_29457);
or UO_1895 (O_1895,N_28489,N_29462);
and UO_1896 (O_1896,N_28908,N_28204);
nand UO_1897 (O_1897,N_28015,N_28034);
nor UO_1898 (O_1898,N_29564,N_28141);
nand UO_1899 (O_1899,N_28744,N_29770);
nor UO_1900 (O_1900,N_29586,N_29305);
xnor UO_1901 (O_1901,N_28197,N_28079);
nor UO_1902 (O_1902,N_29677,N_28451);
nand UO_1903 (O_1903,N_29619,N_28656);
xnor UO_1904 (O_1904,N_29827,N_29577);
or UO_1905 (O_1905,N_28970,N_28734);
xor UO_1906 (O_1906,N_28629,N_29418);
nor UO_1907 (O_1907,N_28292,N_28852);
and UO_1908 (O_1908,N_28184,N_29222);
or UO_1909 (O_1909,N_28724,N_29200);
nor UO_1910 (O_1910,N_28879,N_29004);
nor UO_1911 (O_1911,N_28270,N_29438);
xnor UO_1912 (O_1912,N_29312,N_28146);
and UO_1913 (O_1913,N_28342,N_28654);
nand UO_1914 (O_1914,N_28567,N_29054);
nor UO_1915 (O_1915,N_28007,N_28069);
nand UO_1916 (O_1916,N_28616,N_28126);
nand UO_1917 (O_1917,N_29405,N_29110);
and UO_1918 (O_1918,N_29741,N_28739);
nand UO_1919 (O_1919,N_28834,N_29686);
or UO_1920 (O_1920,N_29868,N_29273);
xor UO_1921 (O_1921,N_28371,N_29576);
nor UO_1922 (O_1922,N_29242,N_28717);
nand UO_1923 (O_1923,N_28522,N_29399);
xor UO_1924 (O_1924,N_29631,N_28860);
and UO_1925 (O_1925,N_28454,N_29969);
nor UO_1926 (O_1926,N_28315,N_28074);
nor UO_1927 (O_1927,N_29740,N_29232);
xor UO_1928 (O_1928,N_29143,N_28252);
nor UO_1929 (O_1929,N_28966,N_28934);
xnor UO_1930 (O_1930,N_28427,N_29874);
and UO_1931 (O_1931,N_28590,N_28476);
or UO_1932 (O_1932,N_29818,N_29163);
nor UO_1933 (O_1933,N_29702,N_29187);
nor UO_1934 (O_1934,N_29658,N_28899);
and UO_1935 (O_1935,N_28969,N_28512);
nor UO_1936 (O_1936,N_28922,N_28694);
nor UO_1937 (O_1937,N_28253,N_28427);
and UO_1938 (O_1938,N_29958,N_29332);
nand UO_1939 (O_1939,N_29139,N_28438);
nor UO_1940 (O_1940,N_29174,N_29815);
or UO_1941 (O_1941,N_28395,N_29741);
nand UO_1942 (O_1942,N_28295,N_28537);
xnor UO_1943 (O_1943,N_28972,N_28408);
nor UO_1944 (O_1944,N_29224,N_28473);
nor UO_1945 (O_1945,N_29525,N_29752);
and UO_1946 (O_1946,N_28709,N_28811);
nand UO_1947 (O_1947,N_28019,N_29543);
and UO_1948 (O_1948,N_28898,N_29999);
and UO_1949 (O_1949,N_29266,N_28406);
nand UO_1950 (O_1950,N_29363,N_29939);
nand UO_1951 (O_1951,N_29509,N_28402);
nand UO_1952 (O_1952,N_28454,N_29843);
nand UO_1953 (O_1953,N_29682,N_28907);
xnor UO_1954 (O_1954,N_28959,N_29145);
or UO_1955 (O_1955,N_28380,N_28137);
nand UO_1956 (O_1956,N_29986,N_29495);
and UO_1957 (O_1957,N_28701,N_28087);
xor UO_1958 (O_1958,N_28279,N_28589);
xnor UO_1959 (O_1959,N_29733,N_28586);
nand UO_1960 (O_1960,N_29973,N_28910);
or UO_1961 (O_1961,N_28903,N_28284);
xor UO_1962 (O_1962,N_28979,N_28175);
nand UO_1963 (O_1963,N_29495,N_28631);
and UO_1964 (O_1964,N_29063,N_29975);
nor UO_1965 (O_1965,N_28192,N_29527);
nand UO_1966 (O_1966,N_28509,N_28378);
or UO_1967 (O_1967,N_28701,N_29534);
xor UO_1968 (O_1968,N_28902,N_28865);
nand UO_1969 (O_1969,N_28610,N_29673);
and UO_1970 (O_1970,N_29457,N_28611);
nand UO_1971 (O_1971,N_29438,N_29913);
or UO_1972 (O_1972,N_29197,N_28425);
or UO_1973 (O_1973,N_28927,N_28295);
or UO_1974 (O_1974,N_28090,N_29758);
and UO_1975 (O_1975,N_28201,N_29147);
nor UO_1976 (O_1976,N_29210,N_28334);
xnor UO_1977 (O_1977,N_28252,N_29955);
and UO_1978 (O_1978,N_28219,N_28613);
nor UO_1979 (O_1979,N_28049,N_29119);
nor UO_1980 (O_1980,N_28054,N_28995);
or UO_1981 (O_1981,N_29939,N_28986);
xor UO_1982 (O_1982,N_28844,N_28848);
xor UO_1983 (O_1983,N_29143,N_29635);
nand UO_1984 (O_1984,N_29982,N_28040);
nor UO_1985 (O_1985,N_29314,N_28017);
and UO_1986 (O_1986,N_28946,N_29946);
nor UO_1987 (O_1987,N_29910,N_28366);
or UO_1988 (O_1988,N_28460,N_29827);
nor UO_1989 (O_1989,N_28945,N_28912);
and UO_1990 (O_1990,N_29314,N_29797);
and UO_1991 (O_1991,N_28469,N_28011);
nand UO_1992 (O_1992,N_29114,N_28953);
or UO_1993 (O_1993,N_29895,N_29198);
xnor UO_1994 (O_1994,N_29259,N_29844);
nor UO_1995 (O_1995,N_28767,N_28092);
or UO_1996 (O_1996,N_29862,N_28324);
and UO_1997 (O_1997,N_28549,N_28554);
xnor UO_1998 (O_1998,N_29948,N_29445);
and UO_1999 (O_1999,N_28394,N_28335);
and UO_2000 (O_2000,N_29423,N_29127);
nand UO_2001 (O_2001,N_28532,N_28468);
nor UO_2002 (O_2002,N_28389,N_29444);
and UO_2003 (O_2003,N_28795,N_28342);
nand UO_2004 (O_2004,N_29029,N_28853);
or UO_2005 (O_2005,N_29802,N_29864);
or UO_2006 (O_2006,N_29905,N_28521);
nor UO_2007 (O_2007,N_29017,N_29613);
xnor UO_2008 (O_2008,N_28290,N_29918);
nor UO_2009 (O_2009,N_29710,N_29518);
xor UO_2010 (O_2010,N_29914,N_28191);
or UO_2011 (O_2011,N_28335,N_29493);
and UO_2012 (O_2012,N_28134,N_29156);
nand UO_2013 (O_2013,N_29316,N_28317);
nor UO_2014 (O_2014,N_28505,N_28699);
xor UO_2015 (O_2015,N_28804,N_29696);
nand UO_2016 (O_2016,N_28137,N_28457);
and UO_2017 (O_2017,N_28203,N_28928);
nor UO_2018 (O_2018,N_29920,N_28460);
or UO_2019 (O_2019,N_29250,N_28164);
or UO_2020 (O_2020,N_29394,N_29444);
and UO_2021 (O_2021,N_28336,N_28042);
and UO_2022 (O_2022,N_28609,N_29365);
and UO_2023 (O_2023,N_29752,N_28037);
nand UO_2024 (O_2024,N_28612,N_28700);
nor UO_2025 (O_2025,N_28635,N_29831);
xnor UO_2026 (O_2026,N_28860,N_28000);
xor UO_2027 (O_2027,N_29760,N_29389);
xor UO_2028 (O_2028,N_28663,N_28269);
xnor UO_2029 (O_2029,N_28319,N_29261);
and UO_2030 (O_2030,N_29457,N_29799);
or UO_2031 (O_2031,N_28298,N_28851);
or UO_2032 (O_2032,N_29871,N_29345);
and UO_2033 (O_2033,N_29333,N_29986);
or UO_2034 (O_2034,N_29782,N_28569);
nor UO_2035 (O_2035,N_28918,N_29636);
and UO_2036 (O_2036,N_28774,N_28174);
nor UO_2037 (O_2037,N_28194,N_29462);
nand UO_2038 (O_2038,N_28932,N_29634);
or UO_2039 (O_2039,N_28458,N_28176);
nand UO_2040 (O_2040,N_28024,N_28572);
and UO_2041 (O_2041,N_28426,N_28451);
nor UO_2042 (O_2042,N_28631,N_29310);
nand UO_2043 (O_2043,N_28277,N_29327);
nor UO_2044 (O_2044,N_29065,N_28990);
or UO_2045 (O_2045,N_29478,N_29738);
nor UO_2046 (O_2046,N_28582,N_28410);
xnor UO_2047 (O_2047,N_29287,N_28623);
nor UO_2048 (O_2048,N_29411,N_29235);
and UO_2049 (O_2049,N_29461,N_28761);
or UO_2050 (O_2050,N_28606,N_28459);
or UO_2051 (O_2051,N_29064,N_29887);
xor UO_2052 (O_2052,N_29991,N_29612);
nor UO_2053 (O_2053,N_28081,N_28905);
nand UO_2054 (O_2054,N_28341,N_28888);
nor UO_2055 (O_2055,N_28138,N_29968);
or UO_2056 (O_2056,N_29792,N_29084);
and UO_2057 (O_2057,N_29217,N_29884);
nor UO_2058 (O_2058,N_29584,N_29270);
and UO_2059 (O_2059,N_28342,N_28110);
xor UO_2060 (O_2060,N_29988,N_29781);
and UO_2061 (O_2061,N_28173,N_29644);
and UO_2062 (O_2062,N_29405,N_28687);
nor UO_2063 (O_2063,N_28884,N_29957);
nand UO_2064 (O_2064,N_28502,N_29976);
nand UO_2065 (O_2065,N_28905,N_29957);
and UO_2066 (O_2066,N_29210,N_28043);
nand UO_2067 (O_2067,N_28638,N_28810);
nor UO_2068 (O_2068,N_28732,N_29600);
and UO_2069 (O_2069,N_29901,N_29161);
or UO_2070 (O_2070,N_29226,N_29231);
nor UO_2071 (O_2071,N_29460,N_28072);
and UO_2072 (O_2072,N_29655,N_28041);
xnor UO_2073 (O_2073,N_28622,N_29358);
nand UO_2074 (O_2074,N_29892,N_29131);
nand UO_2075 (O_2075,N_29172,N_28652);
nand UO_2076 (O_2076,N_29633,N_29290);
nor UO_2077 (O_2077,N_29368,N_28797);
nand UO_2078 (O_2078,N_29647,N_28745);
or UO_2079 (O_2079,N_28111,N_29232);
or UO_2080 (O_2080,N_28413,N_28586);
or UO_2081 (O_2081,N_29385,N_29302);
xnor UO_2082 (O_2082,N_28012,N_29130);
nor UO_2083 (O_2083,N_28356,N_29093);
or UO_2084 (O_2084,N_29002,N_28512);
and UO_2085 (O_2085,N_28635,N_29512);
and UO_2086 (O_2086,N_28610,N_28375);
and UO_2087 (O_2087,N_29451,N_29147);
or UO_2088 (O_2088,N_29621,N_28342);
and UO_2089 (O_2089,N_28822,N_28084);
xor UO_2090 (O_2090,N_28094,N_29291);
and UO_2091 (O_2091,N_28972,N_29788);
nor UO_2092 (O_2092,N_29352,N_29216);
nand UO_2093 (O_2093,N_29631,N_29927);
or UO_2094 (O_2094,N_28134,N_28550);
or UO_2095 (O_2095,N_28410,N_28027);
nor UO_2096 (O_2096,N_28443,N_28761);
nor UO_2097 (O_2097,N_28482,N_28063);
nand UO_2098 (O_2098,N_29126,N_28176);
nand UO_2099 (O_2099,N_28468,N_29758);
nor UO_2100 (O_2100,N_28338,N_28668);
nand UO_2101 (O_2101,N_28174,N_29154);
nand UO_2102 (O_2102,N_28171,N_29450);
xnor UO_2103 (O_2103,N_28177,N_28837);
nor UO_2104 (O_2104,N_29866,N_29042);
nand UO_2105 (O_2105,N_29453,N_29861);
and UO_2106 (O_2106,N_29897,N_28747);
nand UO_2107 (O_2107,N_28795,N_29431);
nand UO_2108 (O_2108,N_28983,N_29282);
xor UO_2109 (O_2109,N_28763,N_29205);
or UO_2110 (O_2110,N_28096,N_28053);
nor UO_2111 (O_2111,N_29033,N_29231);
xnor UO_2112 (O_2112,N_28488,N_28409);
or UO_2113 (O_2113,N_28932,N_29568);
and UO_2114 (O_2114,N_28505,N_29364);
or UO_2115 (O_2115,N_29276,N_28941);
xnor UO_2116 (O_2116,N_28768,N_29315);
nand UO_2117 (O_2117,N_29663,N_29069);
xnor UO_2118 (O_2118,N_28353,N_29615);
nand UO_2119 (O_2119,N_28516,N_29675);
xor UO_2120 (O_2120,N_28077,N_29145);
xnor UO_2121 (O_2121,N_29668,N_28242);
nand UO_2122 (O_2122,N_29920,N_28305);
or UO_2123 (O_2123,N_29473,N_29653);
and UO_2124 (O_2124,N_29839,N_29552);
and UO_2125 (O_2125,N_28887,N_28610);
and UO_2126 (O_2126,N_28880,N_28392);
or UO_2127 (O_2127,N_29702,N_28583);
nor UO_2128 (O_2128,N_29821,N_28848);
or UO_2129 (O_2129,N_28295,N_28025);
and UO_2130 (O_2130,N_28139,N_29439);
nor UO_2131 (O_2131,N_29703,N_28039);
xnor UO_2132 (O_2132,N_29838,N_28460);
nor UO_2133 (O_2133,N_28330,N_29243);
or UO_2134 (O_2134,N_28273,N_28704);
or UO_2135 (O_2135,N_29304,N_29329);
xor UO_2136 (O_2136,N_29768,N_29760);
nand UO_2137 (O_2137,N_28045,N_29501);
nand UO_2138 (O_2138,N_29280,N_29400);
and UO_2139 (O_2139,N_28931,N_29447);
nand UO_2140 (O_2140,N_28209,N_29435);
nand UO_2141 (O_2141,N_28764,N_28982);
nor UO_2142 (O_2142,N_29787,N_28074);
nand UO_2143 (O_2143,N_28470,N_29336);
and UO_2144 (O_2144,N_28566,N_28412);
nand UO_2145 (O_2145,N_29505,N_28792);
xnor UO_2146 (O_2146,N_29963,N_28081);
nand UO_2147 (O_2147,N_29605,N_29633);
nor UO_2148 (O_2148,N_29783,N_28105);
nor UO_2149 (O_2149,N_28259,N_28893);
and UO_2150 (O_2150,N_28323,N_29569);
or UO_2151 (O_2151,N_29744,N_29620);
and UO_2152 (O_2152,N_29338,N_29812);
nor UO_2153 (O_2153,N_29073,N_28477);
xor UO_2154 (O_2154,N_29673,N_28219);
xnor UO_2155 (O_2155,N_29952,N_29066);
nand UO_2156 (O_2156,N_29086,N_29458);
nand UO_2157 (O_2157,N_29391,N_28884);
nand UO_2158 (O_2158,N_29770,N_29678);
nand UO_2159 (O_2159,N_29129,N_28177);
nand UO_2160 (O_2160,N_29126,N_28012);
and UO_2161 (O_2161,N_28993,N_29178);
and UO_2162 (O_2162,N_29750,N_29945);
nand UO_2163 (O_2163,N_28138,N_29265);
and UO_2164 (O_2164,N_29454,N_29230);
and UO_2165 (O_2165,N_29192,N_29116);
or UO_2166 (O_2166,N_28402,N_28551);
nand UO_2167 (O_2167,N_29762,N_29435);
xor UO_2168 (O_2168,N_29356,N_29543);
or UO_2169 (O_2169,N_29605,N_28371);
nand UO_2170 (O_2170,N_28390,N_28613);
nor UO_2171 (O_2171,N_29168,N_29092);
nand UO_2172 (O_2172,N_28672,N_29233);
and UO_2173 (O_2173,N_28727,N_28289);
nand UO_2174 (O_2174,N_29041,N_29942);
or UO_2175 (O_2175,N_29293,N_29076);
or UO_2176 (O_2176,N_29174,N_28850);
or UO_2177 (O_2177,N_29821,N_28026);
or UO_2178 (O_2178,N_28731,N_29674);
nand UO_2179 (O_2179,N_29315,N_29229);
or UO_2180 (O_2180,N_28132,N_28795);
nand UO_2181 (O_2181,N_29534,N_28046);
xor UO_2182 (O_2182,N_28195,N_29899);
xor UO_2183 (O_2183,N_29120,N_28021);
nor UO_2184 (O_2184,N_28523,N_28568);
and UO_2185 (O_2185,N_29362,N_28567);
nor UO_2186 (O_2186,N_29865,N_29552);
and UO_2187 (O_2187,N_29751,N_29028);
nand UO_2188 (O_2188,N_28956,N_29503);
and UO_2189 (O_2189,N_28770,N_28759);
xor UO_2190 (O_2190,N_29301,N_28431);
nor UO_2191 (O_2191,N_28784,N_29531);
or UO_2192 (O_2192,N_29872,N_28589);
nand UO_2193 (O_2193,N_28354,N_29350);
nor UO_2194 (O_2194,N_28739,N_28783);
nor UO_2195 (O_2195,N_29698,N_29645);
or UO_2196 (O_2196,N_28757,N_28651);
or UO_2197 (O_2197,N_28997,N_29371);
xor UO_2198 (O_2198,N_28531,N_29587);
nand UO_2199 (O_2199,N_28859,N_28151);
nor UO_2200 (O_2200,N_28040,N_28173);
nor UO_2201 (O_2201,N_28826,N_29390);
or UO_2202 (O_2202,N_29940,N_28885);
xnor UO_2203 (O_2203,N_28598,N_29651);
and UO_2204 (O_2204,N_29824,N_29005);
xor UO_2205 (O_2205,N_28890,N_28210);
or UO_2206 (O_2206,N_28969,N_28136);
nor UO_2207 (O_2207,N_28469,N_28878);
nor UO_2208 (O_2208,N_29982,N_28651);
and UO_2209 (O_2209,N_29738,N_28197);
nor UO_2210 (O_2210,N_29060,N_28295);
or UO_2211 (O_2211,N_29533,N_29659);
xor UO_2212 (O_2212,N_29705,N_28715);
and UO_2213 (O_2213,N_29701,N_29274);
and UO_2214 (O_2214,N_28503,N_28154);
and UO_2215 (O_2215,N_29988,N_28435);
and UO_2216 (O_2216,N_28481,N_29191);
or UO_2217 (O_2217,N_29587,N_28003);
nor UO_2218 (O_2218,N_29402,N_29243);
nand UO_2219 (O_2219,N_29685,N_29681);
or UO_2220 (O_2220,N_29444,N_28947);
or UO_2221 (O_2221,N_28074,N_29454);
and UO_2222 (O_2222,N_28842,N_28558);
nand UO_2223 (O_2223,N_28076,N_28656);
nand UO_2224 (O_2224,N_29681,N_29277);
nand UO_2225 (O_2225,N_29684,N_29571);
or UO_2226 (O_2226,N_28930,N_29581);
xnor UO_2227 (O_2227,N_28890,N_28768);
and UO_2228 (O_2228,N_28296,N_29278);
and UO_2229 (O_2229,N_29676,N_28401);
xor UO_2230 (O_2230,N_28485,N_28405);
xnor UO_2231 (O_2231,N_29986,N_28543);
nand UO_2232 (O_2232,N_28028,N_28824);
nand UO_2233 (O_2233,N_29923,N_28725);
and UO_2234 (O_2234,N_29572,N_28667);
xnor UO_2235 (O_2235,N_29041,N_28276);
xnor UO_2236 (O_2236,N_28550,N_28325);
nand UO_2237 (O_2237,N_29366,N_29010);
nand UO_2238 (O_2238,N_29649,N_28479);
nand UO_2239 (O_2239,N_29637,N_28595);
or UO_2240 (O_2240,N_29704,N_29303);
nor UO_2241 (O_2241,N_28440,N_29600);
or UO_2242 (O_2242,N_29328,N_29677);
and UO_2243 (O_2243,N_28745,N_29439);
nand UO_2244 (O_2244,N_29576,N_29905);
or UO_2245 (O_2245,N_29369,N_28853);
and UO_2246 (O_2246,N_28952,N_28238);
nor UO_2247 (O_2247,N_28023,N_28133);
and UO_2248 (O_2248,N_28057,N_29523);
nand UO_2249 (O_2249,N_29199,N_29156);
xnor UO_2250 (O_2250,N_29353,N_28646);
xor UO_2251 (O_2251,N_29811,N_28522);
nor UO_2252 (O_2252,N_29146,N_29005);
nor UO_2253 (O_2253,N_29898,N_29961);
nand UO_2254 (O_2254,N_28508,N_28634);
xor UO_2255 (O_2255,N_29643,N_28403);
xnor UO_2256 (O_2256,N_28894,N_29532);
or UO_2257 (O_2257,N_29235,N_28251);
nand UO_2258 (O_2258,N_28307,N_28141);
xnor UO_2259 (O_2259,N_28677,N_29371);
nand UO_2260 (O_2260,N_28368,N_28661);
and UO_2261 (O_2261,N_28450,N_28074);
nand UO_2262 (O_2262,N_29760,N_28999);
xor UO_2263 (O_2263,N_29822,N_29655);
nor UO_2264 (O_2264,N_29542,N_28088);
or UO_2265 (O_2265,N_29114,N_29172);
nor UO_2266 (O_2266,N_29187,N_29919);
or UO_2267 (O_2267,N_28597,N_29471);
or UO_2268 (O_2268,N_29206,N_28931);
or UO_2269 (O_2269,N_28497,N_29141);
and UO_2270 (O_2270,N_28768,N_28353);
nor UO_2271 (O_2271,N_29059,N_29068);
nor UO_2272 (O_2272,N_28474,N_29312);
nand UO_2273 (O_2273,N_29221,N_29465);
or UO_2274 (O_2274,N_29826,N_29651);
and UO_2275 (O_2275,N_29139,N_28951);
or UO_2276 (O_2276,N_28128,N_29949);
and UO_2277 (O_2277,N_29835,N_28832);
xnor UO_2278 (O_2278,N_28306,N_28239);
or UO_2279 (O_2279,N_29416,N_29196);
or UO_2280 (O_2280,N_29012,N_29165);
or UO_2281 (O_2281,N_29175,N_29885);
or UO_2282 (O_2282,N_28694,N_29261);
or UO_2283 (O_2283,N_28567,N_28410);
xnor UO_2284 (O_2284,N_29098,N_29458);
nand UO_2285 (O_2285,N_28989,N_29486);
nand UO_2286 (O_2286,N_28417,N_28418);
nor UO_2287 (O_2287,N_28230,N_28225);
or UO_2288 (O_2288,N_28111,N_28236);
nor UO_2289 (O_2289,N_28280,N_29886);
xor UO_2290 (O_2290,N_28173,N_29154);
xor UO_2291 (O_2291,N_28752,N_28175);
nor UO_2292 (O_2292,N_29429,N_29901);
or UO_2293 (O_2293,N_28337,N_29036);
xor UO_2294 (O_2294,N_28150,N_28807);
nor UO_2295 (O_2295,N_28240,N_29305);
nand UO_2296 (O_2296,N_28150,N_28236);
xnor UO_2297 (O_2297,N_29283,N_29674);
nor UO_2298 (O_2298,N_28169,N_28830);
xor UO_2299 (O_2299,N_28671,N_28075);
nor UO_2300 (O_2300,N_29850,N_29086);
nand UO_2301 (O_2301,N_28169,N_28251);
or UO_2302 (O_2302,N_29862,N_28385);
nor UO_2303 (O_2303,N_28377,N_29940);
nand UO_2304 (O_2304,N_28209,N_28579);
nor UO_2305 (O_2305,N_28031,N_29139);
nor UO_2306 (O_2306,N_29640,N_29891);
nor UO_2307 (O_2307,N_28240,N_29933);
nand UO_2308 (O_2308,N_28561,N_29143);
or UO_2309 (O_2309,N_29995,N_29502);
or UO_2310 (O_2310,N_29217,N_29687);
nor UO_2311 (O_2311,N_29693,N_29957);
nand UO_2312 (O_2312,N_28056,N_28882);
or UO_2313 (O_2313,N_29220,N_28678);
or UO_2314 (O_2314,N_29342,N_29325);
and UO_2315 (O_2315,N_28507,N_29761);
xnor UO_2316 (O_2316,N_28888,N_28184);
or UO_2317 (O_2317,N_29276,N_29328);
nor UO_2318 (O_2318,N_29472,N_28339);
xor UO_2319 (O_2319,N_28451,N_29693);
nand UO_2320 (O_2320,N_29923,N_28761);
and UO_2321 (O_2321,N_29720,N_28283);
and UO_2322 (O_2322,N_29183,N_29276);
and UO_2323 (O_2323,N_28887,N_28990);
nand UO_2324 (O_2324,N_28882,N_28614);
xor UO_2325 (O_2325,N_28460,N_29293);
xor UO_2326 (O_2326,N_28806,N_28318);
and UO_2327 (O_2327,N_29977,N_28874);
nor UO_2328 (O_2328,N_29298,N_28416);
nor UO_2329 (O_2329,N_29526,N_28421);
nand UO_2330 (O_2330,N_29601,N_29856);
or UO_2331 (O_2331,N_29229,N_28388);
xnor UO_2332 (O_2332,N_29670,N_28516);
and UO_2333 (O_2333,N_28805,N_28065);
nor UO_2334 (O_2334,N_28901,N_28830);
and UO_2335 (O_2335,N_29507,N_29285);
and UO_2336 (O_2336,N_28645,N_28934);
or UO_2337 (O_2337,N_28028,N_28042);
and UO_2338 (O_2338,N_28482,N_29939);
xor UO_2339 (O_2339,N_29551,N_29276);
nand UO_2340 (O_2340,N_28303,N_29005);
nand UO_2341 (O_2341,N_29102,N_29481);
nand UO_2342 (O_2342,N_28373,N_28135);
or UO_2343 (O_2343,N_28304,N_29665);
or UO_2344 (O_2344,N_28184,N_28686);
nand UO_2345 (O_2345,N_29251,N_28203);
nand UO_2346 (O_2346,N_29157,N_29431);
nand UO_2347 (O_2347,N_29903,N_29750);
xor UO_2348 (O_2348,N_29416,N_29595);
nor UO_2349 (O_2349,N_28315,N_28833);
nand UO_2350 (O_2350,N_29762,N_29635);
nand UO_2351 (O_2351,N_28484,N_29302);
nor UO_2352 (O_2352,N_28004,N_29010);
and UO_2353 (O_2353,N_28183,N_28682);
or UO_2354 (O_2354,N_28214,N_29329);
xnor UO_2355 (O_2355,N_29812,N_29443);
nand UO_2356 (O_2356,N_28059,N_29950);
nor UO_2357 (O_2357,N_28248,N_28876);
and UO_2358 (O_2358,N_29326,N_29609);
nor UO_2359 (O_2359,N_28896,N_28988);
xor UO_2360 (O_2360,N_28664,N_29171);
nor UO_2361 (O_2361,N_28611,N_29376);
and UO_2362 (O_2362,N_28162,N_28460);
nor UO_2363 (O_2363,N_29451,N_28743);
xnor UO_2364 (O_2364,N_29431,N_28008);
or UO_2365 (O_2365,N_28463,N_28452);
xnor UO_2366 (O_2366,N_28781,N_28833);
nand UO_2367 (O_2367,N_29368,N_28267);
or UO_2368 (O_2368,N_29695,N_28167);
and UO_2369 (O_2369,N_29011,N_29192);
nand UO_2370 (O_2370,N_28328,N_29167);
nand UO_2371 (O_2371,N_29816,N_28690);
or UO_2372 (O_2372,N_29380,N_29797);
nand UO_2373 (O_2373,N_29934,N_28293);
xor UO_2374 (O_2374,N_28465,N_29067);
xnor UO_2375 (O_2375,N_28701,N_29479);
and UO_2376 (O_2376,N_29361,N_29650);
xor UO_2377 (O_2377,N_29186,N_29043);
xor UO_2378 (O_2378,N_28683,N_28845);
nand UO_2379 (O_2379,N_28537,N_28776);
or UO_2380 (O_2380,N_29055,N_29556);
nand UO_2381 (O_2381,N_29222,N_29839);
xor UO_2382 (O_2382,N_29908,N_29879);
nand UO_2383 (O_2383,N_29786,N_29827);
or UO_2384 (O_2384,N_29230,N_28893);
or UO_2385 (O_2385,N_28151,N_28873);
or UO_2386 (O_2386,N_28518,N_29505);
nand UO_2387 (O_2387,N_29617,N_29151);
xnor UO_2388 (O_2388,N_29655,N_29587);
or UO_2389 (O_2389,N_28328,N_29503);
nand UO_2390 (O_2390,N_28025,N_28036);
and UO_2391 (O_2391,N_28775,N_29283);
nor UO_2392 (O_2392,N_29011,N_29104);
xor UO_2393 (O_2393,N_28492,N_29247);
or UO_2394 (O_2394,N_29274,N_28061);
or UO_2395 (O_2395,N_29978,N_28568);
or UO_2396 (O_2396,N_28545,N_29664);
or UO_2397 (O_2397,N_29914,N_29060);
and UO_2398 (O_2398,N_28836,N_28983);
and UO_2399 (O_2399,N_29633,N_29296);
nor UO_2400 (O_2400,N_28735,N_29995);
nand UO_2401 (O_2401,N_29348,N_28405);
nand UO_2402 (O_2402,N_28164,N_29284);
nand UO_2403 (O_2403,N_28895,N_29374);
nor UO_2404 (O_2404,N_29323,N_29142);
xor UO_2405 (O_2405,N_29855,N_29528);
nor UO_2406 (O_2406,N_29295,N_28427);
and UO_2407 (O_2407,N_29353,N_28098);
or UO_2408 (O_2408,N_28687,N_29106);
nand UO_2409 (O_2409,N_29412,N_28623);
xor UO_2410 (O_2410,N_28329,N_28944);
xnor UO_2411 (O_2411,N_28747,N_29650);
nand UO_2412 (O_2412,N_29524,N_28729);
xnor UO_2413 (O_2413,N_28162,N_29369);
nor UO_2414 (O_2414,N_28138,N_29257);
nand UO_2415 (O_2415,N_28880,N_29407);
xor UO_2416 (O_2416,N_29929,N_28412);
or UO_2417 (O_2417,N_28437,N_28924);
and UO_2418 (O_2418,N_28750,N_28350);
or UO_2419 (O_2419,N_29758,N_28773);
nand UO_2420 (O_2420,N_29414,N_28255);
and UO_2421 (O_2421,N_29044,N_29969);
nor UO_2422 (O_2422,N_29980,N_28697);
nand UO_2423 (O_2423,N_28496,N_28922);
nand UO_2424 (O_2424,N_29073,N_29087);
or UO_2425 (O_2425,N_28665,N_29800);
or UO_2426 (O_2426,N_29474,N_29818);
or UO_2427 (O_2427,N_28262,N_28734);
nor UO_2428 (O_2428,N_28726,N_29828);
or UO_2429 (O_2429,N_28581,N_28218);
nor UO_2430 (O_2430,N_29783,N_29931);
or UO_2431 (O_2431,N_29203,N_29504);
nand UO_2432 (O_2432,N_29227,N_28712);
nor UO_2433 (O_2433,N_28448,N_28728);
and UO_2434 (O_2434,N_28748,N_29861);
xnor UO_2435 (O_2435,N_28170,N_28703);
and UO_2436 (O_2436,N_28909,N_29899);
and UO_2437 (O_2437,N_28880,N_29957);
xnor UO_2438 (O_2438,N_29019,N_28391);
and UO_2439 (O_2439,N_29258,N_28383);
xnor UO_2440 (O_2440,N_28172,N_29538);
nand UO_2441 (O_2441,N_29525,N_28587);
xnor UO_2442 (O_2442,N_28500,N_28525);
nand UO_2443 (O_2443,N_28123,N_28765);
or UO_2444 (O_2444,N_28055,N_28393);
nand UO_2445 (O_2445,N_28995,N_28920);
nor UO_2446 (O_2446,N_29099,N_28183);
nand UO_2447 (O_2447,N_28876,N_28096);
xor UO_2448 (O_2448,N_29042,N_29626);
nand UO_2449 (O_2449,N_28280,N_29747);
and UO_2450 (O_2450,N_29105,N_28515);
nor UO_2451 (O_2451,N_29101,N_29617);
xor UO_2452 (O_2452,N_28369,N_28814);
xor UO_2453 (O_2453,N_28923,N_28478);
xor UO_2454 (O_2454,N_28388,N_29774);
nand UO_2455 (O_2455,N_28354,N_28914);
or UO_2456 (O_2456,N_28236,N_28039);
or UO_2457 (O_2457,N_29924,N_28658);
nand UO_2458 (O_2458,N_28078,N_28960);
and UO_2459 (O_2459,N_29481,N_28504);
or UO_2460 (O_2460,N_29873,N_29777);
or UO_2461 (O_2461,N_28401,N_29383);
or UO_2462 (O_2462,N_28743,N_29158);
nor UO_2463 (O_2463,N_29463,N_29988);
nand UO_2464 (O_2464,N_29436,N_29069);
nor UO_2465 (O_2465,N_28460,N_28133);
or UO_2466 (O_2466,N_28744,N_28423);
nor UO_2467 (O_2467,N_28832,N_29754);
xor UO_2468 (O_2468,N_28200,N_29278);
xnor UO_2469 (O_2469,N_28311,N_28900);
and UO_2470 (O_2470,N_28370,N_28272);
or UO_2471 (O_2471,N_29001,N_28221);
xor UO_2472 (O_2472,N_29817,N_29612);
xnor UO_2473 (O_2473,N_29492,N_29382);
nor UO_2474 (O_2474,N_28071,N_28176);
or UO_2475 (O_2475,N_29912,N_29663);
and UO_2476 (O_2476,N_28884,N_29774);
nor UO_2477 (O_2477,N_28682,N_28732);
xor UO_2478 (O_2478,N_29491,N_28775);
or UO_2479 (O_2479,N_29019,N_28081);
nor UO_2480 (O_2480,N_28838,N_28311);
xor UO_2481 (O_2481,N_28445,N_28464);
nand UO_2482 (O_2482,N_28185,N_28379);
and UO_2483 (O_2483,N_29141,N_29506);
xor UO_2484 (O_2484,N_28934,N_29365);
and UO_2485 (O_2485,N_28790,N_29349);
and UO_2486 (O_2486,N_29080,N_28141);
xnor UO_2487 (O_2487,N_29695,N_29601);
or UO_2488 (O_2488,N_28709,N_29631);
xor UO_2489 (O_2489,N_28849,N_28118);
xnor UO_2490 (O_2490,N_28153,N_29708);
nand UO_2491 (O_2491,N_28180,N_28859);
nor UO_2492 (O_2492,N_28777,N_28421);
xnor UO_2493 (O_2493,N_28365,N_28425);
or UO_2494 (O_2494,N_28436,N_29273);
and UO_2495 (O_2495,N_29915,N_28266);
or UO_2496 (O_2496,N_29553,N_28946);
nor UO_2497 (O_2497,N_29354,N_28037);
xor UO_2498 (O_2498,N_28325,N_28563);
and UO_2499 (O_2499,N_29701,N_29943);
nor UO_2500 (O_2500,N_28337,N_29119);
nand UO_2501 (O_2501,N_28775,N_28120);
nor UO_2502 (O_2502,N_29186,N_28023);
nand UO_2503 (O_2503,N_29511,N_28772);
xor UO_2504 (O_2504,N_28306,N_28736);
nor UO_2505 (O_2505,N_29564,N_28958);
and UO_2506 (O_2506,N_28913,N_28221);
or UO_2507 (O_2507,N_29115,N_28991);
nand UO_2508 (O_2508,N_29861,N_28947);
and UO_2509 (O_2509,N_28246,N_29204);
nand UO_2510 (O_2510,N_29114,N_28882);
nand UO_2511 (O_2511,N_29041,N_28371);
nor UO_2512 (O_2512,N_29329,N_28420);
and UO_2513 (O_2513,N_28776,N_29180);
nor UO_2514 (O_2514,N_28045,N_28963);
nor UO_2515 (O_2515,N_28537,N_28837);
nor UO_2516 (O_2516,N_29264,N_28470);
xnor UO_2517 (O_2517,N_28476,N_28740);
or UO_2518 (O_2518,N_28503,N_29136);
and UO_2519 (O_2519,N_29035,N_29397);
or UO_2520 (O_2520,N_29011,N_28038);
nor UO_2521 (O_2521,N_29216,N_28903);
nor UO_2522 (O_2522,N_28456,N_28765);
or UO_2523 (O_2523,N_28272,N_29886);
xor UO_2524 (O_2524,N_29317,N_28588);
xor UO_2525 (O_2525,N_28245,N_28343);
and UO_2526 (O_2526,N_29440,N_28087);
and UO_2527 (O_2527,N_29426,N_28005);
and UO_2528 (O_2528,N_29396,N_29374);
and UO_2529 (O_2529,N_29727,N_29663);
nand UO_2530 (O_2530,N_29811,N_29833);
xnor UO_2531 (O_2531,N_28627,N_29865);
nand UO_2532 (O_2532,N_29617,N_28602);
xnor UO_2533 (O_2533,N_29371,N_28424);
nand UO_2534 (O_2534,N_28177,N_29590);
nor UO_2535 (O_2535,N_28326,N_29637);
nor UO_2536 (O_2536,N_29045,N_29695);
nand UO_2537 (O_2537,N_28255,N_28128);
and UO_2538 (O_2538,N_28331,N_29535);
nand UO_2539 (O_2539,N_28881,N_28833);
nor UO_2540 (O_2540,N_29263,N_28473);
or UO_2541 (O_2541,N_29067,N_28359);
or UO_2542 (O_2542,N_29321,N_29202);
xor UO_2543 (O_2543,N_28920,N_29750);
xnor UO_2544 (O_2544,N_28535,N_28445);
xor UO_2545 (O_2545,N_28095,N_28847);
and UO_2546 (O_2546,N_29304,N_28551);
nor UO_2547 (O_2547,N_29685,N_28755);
and UO_2548 (O_2548,N_28052,N_29641);
nor UO_2549 (O_2549,N_28159,N_28670);
xor UO_2550 (O_2550,N_29850,N_29749);
and UO_2551 (O_2551,N_28674,N_28011);
and UO_2552 (O_2552,N_29742,N_29976);
nor UO_2553 (O_2553,N_28976,N_29859);
nor UO_2554 (O_2554,N_29518,N_29976);
and UO_2555 (O_2555,N_29331,N_28836);
nand UO_2556 (O_2556,N_28021,N_29485);
or UO_2557 (O_2557,N_29571,N_29192);
nand UO_2558 (O_2558,N_29464,N_28821);
xnor UO_2559 (O_2559,N_28543,N_28824);
nor UO_2560 (O_2560,N_28605,N_29834);
xnor UO_2561 (O_2561,N_28149,N_29517);
and UO_2562 (O_2562,N_28345,N_29140);
xnor UO_2563 (O_2563,N_29568,N_28852);
xnor UO_2564 (O_2564,N_29903,N_29015);
nor UO_2565 (O_2565,N_29986,N_28515);
or UO_2566 (O_2566,N_28155,N_29236);
and UO_2567 (O_2567,N_28114,N_29393);
and UO_2568 (O_2568,N_29820,N_29362);
nand UO_2569 (O_2569,N_28667,N_29851);
xor UO_2570 (O_2570,N_29640,N_29060);
nor UO_2571 (O_2571,N_28766,N_28151);
nor UO_2572 (O_2572,N_28385,N_28344);
nor UO_2573 (O_2573,N_28512,N_28088);
nand UO_2574 (O_2574,N_28893,N_28553);
and UO_2575 (O_2575,N_29093,N_29696);
nand UO_2576 (O_2576,N_29457,N_29456);
or UO_2577 (O_2577,N_29490,N_28075);
or UO_2578 (O_2578,N_28401,N_28825);
and UO_2579 (O_2579,N_28016,N_29888);
nor UO_2580 (O_2580,N_28309,N_29542);
and UO_2581 (O_2581,N_29841,N_29193);
nand UO_2582 (O_2582,N_28858,N_28450);
or UO_2583 (O_2583,N_29859,N_29613);
xnor UO_2584 (O_2584,N_29656,N_28996);
xnor UO_2585 (O_2585,N_29874,N_28048);
xnor UO_2586 (O_2586,N_29087,N_28927);
xnor UO_2587 (O_2587,N_29258,N_28302);
and UO_2588 (O_2588,N_28384,N_28507);
nand UO_2589 (O_2589,N_28265,N_28591);
nor UO_2590 (O_2590,N_29001,N_28505);
nand UO_2591 (O_2591,N_29625,N_29312);
nor UO_2592 (O_2592,N_28056,N_28920);
and UO_2593 (O_2593,N_29978,N_29999);
and UO_2594 (O_2594,N_28219,N_28008);
xor UO_2595 (O_2595,N_29523,N_29659);
nand UO_2596 (O_2596,N_29186,N_28965);
nor UO_2597 (O_2597,N_28187,N_28288);
xor UO_2598 (O_2598,N_28964,N_29703);
nor UO_2599 (O_2599,N_29497,N_29284);
xor UO_2600 (O_2600,N_28491,N_28655);
nand UO_2601 (O_2601,N_28692,N_28251);
xor UO_2602 (O_2602,N_28170,N_28171);
nand UO_2603 (O_2603,N_29279,N_29634);
xor UO_2604 (O_2604,N_28860,N_28238);
nor UO_2605 (O_2605,N_28309,N_28358);
or UO_2606 (O_2606,N_29319,N_29518);
nor UO_2607 (O_2607,N_28009,N_29168);
or UO_2608 (O_2608,N_29602,N_28086);
nor UO_2609 (O_2609,N_28556,N_29140);
nand UO_2610 (O_2610,N_28001,N_29998);
nand UO_2611 (O_2611,N_29042,N_28871);
nor UO_2612 (O_2612,N_29425,N_29701);
xnor UO_2613 (O_2613,N_28520,N_28144);
nand UO_2614 (O_2614,N_28488,N_28907);
or UO_2615 (O_2615,N_28828,N_28602);
nor UO_2616 (O_2616,N_28728,N_29041);
nand UO_2617 (O_2617,N_28010,N_29110);
xor UO_2618 (O_2618,N_28085,N_29281);
xnor UO_2619 (O_2619,N_29134,N_29574);
nor UO_2620 (O_2620,N_28144,N_29199);
or UO_2621 (O_2621,N_29979,N_28810);
nor UO_2622 (O_2622,N_29726,N_28528);
xor UO_2623 (O_2623,N_28269,N_28912);
nor UO_2624 (O_2624,N_28556,N_28979);
xor UO_2625 (O_2625,N_29169,N_29786);
and UO_2626 (O_2626,N_29001,N_28215);
and UO_2627 (O_2627,N_29123,N_29834);
nor UO_2628 (O_2628,N_29923,N_28062);
nand UO_2629 (O_2629,N_28771,N_29362);
or UO_2630 (O_2630,N_28597,N_29063);
and UO_2631 (O_2631,N_28525,N_29094);
xnor UO_2632 (O_2632,N_29357,N_28549);
nor UO_2633 (O_2633,N_28376,N_28035);
nor UO_2634 (O_2634,N_29253,N_29283);
and UO_2635 (O_2635,N_28245,N_28029);
nand UO_2636 (O_2636,N_28340,N_29996);
nor UO_2637 (O_2637,N_28703,N_29555);
xnor UO_2638 (O_2638,N_29231,N_29910);
xor UO_2639 (O_2639,N_29389,N_28511);
and UO_2640 (O_2640,N_28339,N_29968);
xnor UO_2641 (O_2641,N_28043,N_28857);
nand UO_2642 (O_2642,N_28256,N_29119);
xor UO_2643 (O_2643,N_29417,N_29905);
or UO_2644 (O_2644,N_28069,N_29787);
or UO_2645 (O_2645,N_29450,N_28243);
or UO_2646 (O_2646,N_29016,N_28912);
nor UO_2647 (O_2647,N_28866,N_28042);
nor UO_2648 (O_2648,N_28283,N_29237);
and UO_2649 (O_2649,N_28189,N_29141);
xor UO_2650 (O_2650,N_29160,N_29616);
or UO_2651 (O_2651,N_29172,N_28363);
and UO_2652 (O_2652,N_29901,N_29052);
or UO_2653 (O_2653,N_28140,N_28838);
nand UO_2654 (O_2654,N_29330,N_29973);
xor UO_2655 (O_2655,N_28615,N_28224);
nor UO_2656 (O_2656,N_29246,N_28508);
and UO_2657 (O_2657,N_29518,N_28424);
or UO_2658 (O_2658,N_28126,N_29815);
nor UO_2659 (O_2659,N_28277,N_29872);
nand UO_2660 (O_2660,N_29642,N_29185);
or UO_2661 (O_2661,N_29503,N_29235);
xor UO_2662 (O_2662,N_29391,N_29252);
and UO_2663 (O_2663,N_28283,N_29322);
nand UO_2664 (O_2664,N_28699,N_29660);
nor UO_2665 (O_2665,N_28451,N_28932);
or UO_2666 (O_2666,N_28793,N_28099);
or UO_2667 (O_2667,N_28193,N_28621);
or UO_2668 (O_2668,N_28460,N_28727);
xnor UO_2669 (O_2669,N_28848,N_28401);
nor UO_2670 (O_2670,N_29451,N_28684);
nor UO_2671 (O_2671,N_29571,N_28968);
nor UO_2672 (O_2672,N_29342,N_28009);
or UO_2673 (O_2673,N_28295,N_29840);
nor UO_2674 (O_2674,N_29616,N_29199);
and UO_2675 (O_2675,N_28056,N_29379);
and UO_2676 (O_2676,N_28525,N_28461);
and UO_2677 (O_2677,N_29273,N_29478);
nand UO_2678 (O_2678,N_28540,N_28253);
nand UO_2679 (O_2679,N_29646,N_29455);
nor UO_2680 (O_2680,N_28287,N_29232);
or UO_2681 (O_2681,N_29616,N_28618);
xor UO_2682 (O_2682,N_28524,N_29081);
or UO_2683 (O_2683,N_29349,N_28220);
xor UO_2684 (O_2684,N_28509,N_29395);
and UO_2685 (O_2685,N_29108,N_28455);
xnor UO_2686 (O_2686,N_29821,N_28113);
nand UO_2687 (O_2687,N_29041,N_28388);
or UO_2688 (O_2688,N_29949,N_29240);
or UO_2689 (O_2689,N_29155,N_28209);
xor UO_2690 (O_2690,N_29558,N_29379);
nor UO_2691 (O_2691,N_29498,N_29205);
xor UO_2692 (O_2692,N_28497,N_29160);
nand UO_2693 (O_2693,N_28107,N_28316);
nor UO_2694 (O_2694,N_28567,N_28911);
xnor UO_2695 (O_2695,N_29043,N_28693);
xnor UO_2696 (O_2696,N_29620,N_29271);
and UO_2697 (O_2697,N_28987,N_28880);
nand UO_2698 (O_2698,N_28139,N_29412);
nand UO_2699 (O_2699,N_29980,N_28466);
nor UO_2700 (O_2700,N_29306,N_29791);
and UO_2701 (O_2701,N_28571,N_29195);
xor UO_2702 (O_2702,N_28568,N_28514);
and UO_2703 (O_2703,N_29895,N_29590);
nor UO_2704 (O_2704,N_29109,N_28483);
xnor UO_2705 (O_2705,N_28565,N_29379);
nor UO_2706 (O_2706,N_28252,N_29056);
nor UO_2707 (O_2707,N_28788,N_28886);
or UO_2708 (O_2708,N_28303,N_29055);
nand UO_2709 (O_2709,N_29145,N_29955);
xor UO_2710 (O_2710,N_28601,N_28164);
nor UO_2711 (O_2711,N_28290,N_29446);
or UO_2712 (O_2712,N_29891,N_29628);
and UO_2713 (O_2713,N_28599,N_28858);
nor UO_2714 (O_2714,N_29587,N_29250);
nor UO_2715 (O_2715,N_29780,N_28907);
xor UO_2716 (O_2716,N_29074,N_29404);
xnor UO_2717 (O_2717,N_28006,N_29465);
nand UO_2718 (O_2718,N_29370,N_28122);
or UO_2719 (O_2719,N_28631,N_28731);
and UO_2720 (O_2720,N_29529,N_28393);
nand UO_2721 (O_2721,N_29652,N_29300);
and UO_2722 (O_2722,N_28800,N_28162);
and UO_2723 (O_2723,N_28406,N_29451);
nor UO_2724 (O_2724,N_29611,N_28125);
or UO_2725 (O_2725,N_28720,N_29332);
nand UO_2726 (O_2726,N_29564,N_29321);
nand UO_2727 (O_2727,N_28762,N_29868);
xor UO_2728 (O_2728,N_29697,N_29041);
nand UO_2729 (O_2729,N_29675,N_28000);
nor UO_2730 (O_2730,N_28815,N_28026);
nand UO_2731 (O_2731,N_28329,N_28198);
or UO_2732 (O_2732,N_29569,N_28638);
and UO_2733 (O_2733,N_29088,N_28023);
and UO_2734 (O_2734,N_29563,N_29270);
or UO_2735 (O_2735,N_29718,N_28751);
and UO_2736 (O_2736,N_29323,N_28749);
or UO_2737 (O_2737,N_28110,N_29507);
xnor UO_2738 (O_2738,N_29516,N_28892);
nand UO_2739 (O_2739,N_28699,N_29786);
or UO_2740 (O_2740,N_28810,N_29500);
nor UO_2741 (O_2741,N_28456,N_29530);
xnor UO_2742 (O_2742,N_28916,N_29517);
or UO_2743 (O_2743,N_29320,N_29815);
nor UO_2744 (O_2744,N_28364,N_28407);
xor UO_2745 (O_2745,N_28603,N_28513);
xor UO_2746 (O_2746,N_28864,N_28556);
and UO_2747 (O_2747,N_28319,N_28930);
nor UO_2748 (O_2748,N_29843,N_28865);
or UO_2749 (O_2749,N_28920,N_29817);
and UO_2750 (O_2750,N_28204,N_29330);
xnor UO_2751 (O_2751,N_28954,N_29990);
nor UO_2752 (O_2752,N_28361,N_28404);
xor UO_2753 (O_2753,N_29131,N_29932);
xor UO_2754 (O_2754,N_29833,N_29212);
nor UO_2755 (O_2755,N_29135,N_28851);
nor UO_2756 (O_2756,N_28086,N_28848);
nor UO_2757 (O_2757,N_29346,N_29900);
xnor UO_2758 (O_2758,N_29115,N_29977);
or UO_2759 (O_2759,N_28286,N_28985);
and UO_2760 (O_2760,N_29473,N_28384);
or UO_2761 (O_2761,N_28637,N_29787);
and UO_2762 (O_2762,N_28625,N_28594);
and UO_2763 (O_2763,N_29981,N_29175);
nand UO_2764 (O_2764,N_28301,N_29959);
and UO_2765 (O_2765,N_28231,N_29755);
nand UO_2766 (O_2766,N_28267,N_29179);
and UO_2767 (O_2767,N_28710,N_29540);
or UO_2768 (O_2768,N_28687,N_28645);
nand UO_2769 (O_2769,N_29420,N_28780);
and UO_2770 (O_2770,N_28872,N_29603);
nor UO_2771 (O_2771,N_28359,N_28738);
xor UO_2772 (O_2772,N_28713,N_29623);
nand UO_2773 (O_2773,N_28316,N_28199);
and UO_2774 (O_2774,N_28901,N_28908);
or UO_2775 (O_2775,N_29023,N_29156);
nand UO_2776 (O_2776,N_29836,N_28342);
nand UO_2777 (O_2777,N_28007,N_29284);
nor UO_2778 (O_2778,N_29805,N_29635);
xnor UO_2779 (O_2779,N_28189,N_28853);
nor UO_2780 (O_2780,N_29285,N_28794);
or UO_2781 (O_2781,N_28483,N_28256);
xor UO_2782 (O_2782,N_29419,N_29671);
nor UO_2783 (O_2783,N_29390,N_28592);
nand UO_2784 (O_2784,N_29170,N_28102);
or UO_2785 (O_2785,N_28265,N_29390);
nand UO_2786 (O_2786,N_28721,N_29959);
nor UO_2787 (O_2787,N_28792,N_28212);
xnor UO_2788 (O_2788,N_29226,N_29095);
or UO_2789 (O_2789,N_28948,N_29679);
or UO_2790 (O_2790,N_28509,N_29835);
nor UO_2791 (O_2791,N_28857,N_28955);
xnor UO_2792 (O_2792,N_29944,N_29758);
and UO_2793 (O_2793,N_29815,N_28116);
xor UO_2794 (O_2794,N_29614,N_29646);
or UO_2795 (O_2795,N_29505,N_29909);
or UO_2796 (O_2796,N_29051,N_29216);
or UO_2797 (O_2797,N_28278,N_29945);
nor UO_2798 (O_2798,N_28914,N_28592);
nor UO_2799 (O_2799,N_28908,N_28669);
nor UO_2800 (O_2800,N_29613,N_28175);
nor UO_2801 (O_2801,N_28915,N_29601);
xnor UO_2802 (O_2802,N_28281,N_28525);
nand UO_2803 (O_2803,N_28198,N_28474);
or UO_2804 (O_2804,N_29692,N_28837);
and UO_2805 (O_2805,N_29484,N_29402);
or UO_2806 (O_2806,N_28999,N_28104);
xnor UO_2807 (O_2807,N_28759,N_29127);
or UO_2808 (O_2808,N_29646,N_29583);
xnor UO_2809 (O_2809,N_29901,N_29954);
nand UO_2810 (O_2810,N_29487,N_29852);
or UO_2811 (O_2811,N_29857,N_28387);
xor UO_2812 (O_2812,N_28211,N_29352);
nand UO_2813 (O_2813,N_29107,N_29223);
and UO_2814 (O_2814,N_28634,N_28589);
xnor UO_2815 (O_2815,N_28766,N_28936);
and UO_2816 (O_2816,N_29514,N_29859);
and UO_2817 (O_2817,N_29086,N_28513);
nor UO_2818 (O_2818,N_29721,N_28112);
and UO_2819 (O_2819,N_28432,N_28237);
xnor UO_2820 (O_2820,N_28564,N_28222);
or UO_2821 (O_2821,N_29809,N_28362);
nor UO_2822 (O_2822,N_28308,N_28035);
and UO_2823 (O_2823,N_29232,N_28865);
and UO_2824 (O_2824,N_28410,N_28820);
and UO_2825 (O_2825,N_28047,N_29734);
and UO_2826 (O_2826,N_28397,N_29063);
or UO_2827 (O_2827,N_29076,N_29016);
nand UO_2828 (O_2828,N_29995,N_28688);
xor UO_2829 (O_2829,N_28527,N_29954);
or UO_2830 (O_2830,N_28214,N_29799);
and UO_2831 (O_2831,N_29685,N_29239);
nor UO_2832 (O_2832,N_29662,N_28479);
nor UO_2833 (O_2833,N_29370,N_28888);
and UO_2834 (O_2834,N_28836,N_28529);
and UO_2835 (O_2835,N_29874,N_29932);
nor UO_2836 (O_2836,N_29481,N_29371);
and UO_2837 (O_2837,N_29220,N_28356);
xor UO_2838 (O_2838,N_28389,N_29908);
nor UO_2839 (O_2839,N_29799,N_28510);
nor UO_2840 (O_2840,N_28250,N_29764);
or UO_2841 (O_2841,N_28522,N_28019);
nand UO_2842 (O_2842,N_28422,N_28689);
nor UO_2843 (O_2843,N_28945,N_29909);
or UO_2844 (O_2844,N_28038,N_28040);
xnor UO_2845 (O_2845,N_29102,N_28053);
nor UO_2846 (O_2846,N_28676,N_29596);
nor UO_2847 (O_2847,N_28330,N_29547);
nand UO_2848 (O_2848,N_29549,N_29242);
nor UO_2849 (O_2849,N_29781,N_29208);
xor UO_2850 (O_2850,N_28039,N_28743);
xnor UO_2851 (O_2851,N_28123,N_29849);
nor UO_2852 (O_2852,N_28046,N_28796);
or UO_2853 (O_2853,N_29627,N_28941);
and UO_2854 (O_2854,N_28261,N_29420);
or UO_2855 (O_2855,N_29118,N_28208);
or UO_2856 (O_2856,N_28480,N_29377);
xnor UO_2857 (O_2857,N_28005,N_28670);
nor UO_2858 (O_2858,N_28170,N_28353);
or UO_2859 (O_2859,N_29938,N_28734);
nand UO_2860 (O_2860,N_28568,N_28919);
nand UO_2861 (O_2861,N_29091,N_28522);
or UO_2862 (O_2862,N_28591,N_29227);
nor UO_2863 (O_2863,N_29136,N_29940);
or UO_2864 (O_2864,N_29740,N_28039);
nand UO_2865 (O_2865,N_29944,N_29816);
and UO_2866 (O_2866,N_28252,N_29318);
or UO_2867 (O_2867,N_29028,N_28321);
and UO_2868 (O_2868,N_29607,N_28534);
nor UO_2869 (O_2869,N_28114,N_29083);
or UO_2870 (O_2870,N_29910,N_29703);
nor UO_2871 (O_2871,N_28742,N_28593);
or UO_2872 (O_2872,N_29301,N_28110);
nor UO_2873 (O_2873,N_29215,N_28932);
or UO_2874 (O_2874,N_29795,N_28471);
xnor UO_2875 (O_2875,N_29742,N_29982);
and UO_2876 (O_2876,N_28116,N_28924);
or UO_2877 (O_2877,N_28008,N_29115);
or UO_2878 (O_2878,N_28417,N_28325);
nor UO_2879 (O_2879,N_29616,N_29567);
or UO_2880 (O_2880,N_28411,N_28912);
nor UO_2881 (O_2881,N_29845,N_29786);
and UO_2882 (O_2882,N_29579,N_29204);
or UO_2883 (O_2883,N_29197,N_28993);
xor UO_2884 (O_2884,N_29892,N_29937);
nor UO_2885 (O_2885,N_29524,N_29022);
nor UO_2886 (O_2886,N_29971,N_29524);
nand UO_2887 (O_2887,N_28767,N_28315);
nand UO_2888 (O_2888,N_28855,N_28699);
and UO_2889 (O_2889,N_29573,N_29110);
nor UO_2890 (O_2890,N_28280,N_29471);
nand UO_2891 (O_2891,N_29988,N_28965);
and UO_2892 (O_2892,N_28333,N_28062);
nor UO_2893 (O_2893,N_29055,N_28625);
nor UO_2894 (O_2894,N_29911,N_29636);
nand UO_2895 (O_2895,N_29385,N_28088);
and UO_2896 (O_2896,N_28366,N_28408);
and UO_2897 (O_2897,N_29493,N_28546);
nor UO_2898 (O_2898,N_29255,N_28271);
nand UO_2899 (O_2899,N_28501,N_28726);
nand UO_2900 (O_2900,N_28881,N_28922);
nor UO_2901 (O_2901,N_28983,N_29975);
nand UO_2902 (O_2902,N_29804,N_29925);
or UO_2903 (O_2903,N_29692,N_29611);
nand UO_2904 (O_2904,N_28138,N_29969);
or UO_2905 (O_2905,N_28813,N_29894);
and UO_2906 (O_2906,N_28945,N_28874);
xor UO_2907 (O_2907,N_29996,N_29535);
xor UO_2908 (O_2908,N_29218,N_29322);
nor UO_2909 (O_2909,N_28032,N_28603);
nor UO_2910 (O_2910,N_28488,N_29071);
nor UO_2911 (O_2911,N_29096,N_29479);
or UO_2912 (O_2912,N_29026,N_29016);
or UO_2913 (O_2913,N_28263,N_29001);
nor UO_2914 (O_2914,N_28425,N_29121);
xor UO_2915 (O_2915,N_29196,N_29114);
and UO_2916 (O_2916,N_29108,N_28646);
nand UO_2917 (O_2917,N_29433,N_28993);
or UO_2918 (O_2918,N_28201,N_29754);
xor UO_2919 (O_2919,N_29737,N_28265);
xor UO_2920 (O_2920,N_29929,N_29294);
nor UO_2921 (O_2921,N_28585,N_29763);
xnor UO_2922 (O_2922,N_28889,N_28791);
nor UO_2923 (O_2923,N_28489,N_29355);
and UO_2924 (O_2924,N_28432,N_28152);
xnor UO_2925 (O_2925,N_28353,N_28194);
nand UO_2926 (O_2926,N_29089,N_28624);
or UO_2927 (O_2927,N_29279,N_29789);
nor UO_2928 (O_2928,N_28748,N_29791);
and UO_2929 (O_2929,N_29026,N_28458);
or UO_2930 (O_2930,N_29958,N_29011);
xnor UO_2931 (O_2931,N_29830,N_28589);
or UO_2932 (O_2932,N_28406,N_29520);
xnor UO_2933 (O_2933,N_28180,N_28313);
or UO_2934 (O_2934,N_29440,N_28771);
nor UO_2935 (O_2935,N_29810,N_28950);
or UO_2936 (O_2936,N_28050,N_29071);
and UO_2937 (O_2937,N_28488,N_29599);
or UO_2938 (O_2938,N_29627,N_29051);
nand UO_2939 (O_2939,N_28221,N_29274);
and UO_2940 (O_2940,N_28222,N_29413);
nor UO_2941 (O_2941,N_28332,N_29951);
or UO_2942 (O_2942,N_29314,N_28190);
or UO_2943 (O_2943,N_28113,N_29798);
nand UO_2944 (O_2944,N_28087,N_29093);
and UO_2945 (O_2945,N_28217,N_28491);
xor UO_2946 (O_2946,N_28649,N_29269);
nor UO_2947 (O_2947,N_29046,N_29352);
and UO_2948 (O_2948,N_29480,N_28330);
nor UO_2949 (O_2949,N_29945,N_28331);
or UO_2950 (O_2950,N_28936,N_29163);
nor UO_2951 (O_2951,N_28957,N_28791);
or UO_2952 (O_2952,N_28476,N_29312);
xor UO_2953 (O_2953,N_28995,N_29448);
xor UO_2954 (O_2954,N_29048,N_28562);
or UO_2955 (O_2955,N_28907,N_28241);
xnor UO_2956 (O_2956,N_29362,N_29773);
and UO_2957 (O_2957,N_29198,N_28418);
and UO_2958 (O_2958,N_29336,N_28927);
or UO_2959 (O_2959,N_28384,N_29034);
or UO_2960 (O_2960,N_28518,N_28197);
or UO_2961 (O_2961,N_29890,N_28005);
nor UO_2962 (O_2962,N_28113,N_29412);
nand UO_2963 (O_2963,N_29022,N_28313);
nand UO_2964 (O_2964,N_28735,N_29210);
xnor UO_2965 (O_2965,N_28303,N_29013);
xor UO_2966 (O_2966,N_28446,N_28615);
or UO_2967 (O_2967,N_28343,N_28316);
xor UO_2968 (O_2968,N_29524,N_28310);
nor UO_2969 (O_2969,N_28106,N_29562);
and UO_2970 (O_2970,N_29444,N_29737);
and UO_2971 (O_2971,N_28030,N_29645);
nand UO_2972 (O_2972,N_28783,N_29375);
xnor UO_2973 (O_2973,N_29878,N_29663);
xor UO_2974 (O_2974,N_28092,N_29831);
xnor UO_2975 (O_2975,N_29607,N_28772);
or UO_2976 (O_2976,N_28184,N_28133);
nor UO_2977 (O_2977,N_29544,N_29879);
or UO_2978 (O_2978,N_29578,N_28020);
and UO_2979 (O_2979,N_29533,N_29534);
xnor UO_2980 (O_2980,N_28508,N_29197);
or UO_2981 (O_2981,N_29842,N_29875);
and UO_2982 (O_2982,N_29909,N_29921);
or UO_2983 (O_2983,N_29487,N_28232);
nand UO_2984 (O_2984,N_29800,N_28750);
xor UO_2985 (O_2985,N_29017,N_28038);
and UO_2986 (O_2986,N_28846,N_28459);
xnor UO_2987 (O_2987,N_29236,N_28721);
xor UO_2988 (O_2988,N_29007,N_28639);
and UO_2989 (O_2989,N_28216,N_29638);
or UO_2990 (O_2990,N_29696,N_29474);
nor UO_2991 (O_2991,N_28555,N_28235);
nor UO_2992 (O_2992,N_28679,N_29798);
or UO_2993 (O_2993,N_29675,N_29084);
xor UO_2994 (O_2994,N_29988,N_29983);
and UO_2995 (O_2995,N_29828,N_29549);
and UO_2996 (O_2996,N_28415,N_29995);
nor UO_2997 (O_2997,N_29650,N_29147);
nor UO_2998 (O_2998,N_28094,N_28629);
xnor UO_2999 (O_2999,N_29775,N_28100);
and UO_3000 (O_3000,N_28193,N_29728);
and UO_3001 (O_3001,N_29648,N_28685);
xnor UO_3002 (O_3002,N_28045,N_29117);
or UO_3003 (O_3003,N_29573,N_28151);
nor UO_3004 (O_3004,N_28803,N_28433);
nor UO_3005 (O_3005,N_28453,N_28989);
or UO_3006 (O_3006,N_28484,N_28600);
nor UO_3007 (O_3007,N_29223,N_29587);
xor UO_3008 (O_3008,N_28524,N_29289);
xor UO_3009 (O_3009,N_28832,N_29514);
or UO_3010 (O_3010,N_28673,N_28743);
or UO_3011 (O_3011,N_28597,N_29459);
and UO_3012 (O_3012,N_28399,N_28582);
nand UO_3013 (O_3013,N_28783,N_29418);
and UO_3014 (O_3014,N_28261,N_29942);
xnor UO_3015 (O_3015,N_28785,N_28462);
xor UO_3016 (O_3016,N_29372,N_29816);
nor UO_3017 (O_3017,N_28876,N_28477);
nor UO_3018 (O_3018,N_28733,N_28871);
and UO_3019 (O_3019,N_28117,N_29771);
nand UO_3020 (O_3020,N_28006,N_29106);
nand UO_3021 (O_3021,N_28553,N_29303);
xor UO_3022 (O_3022,N_28237,N_28352);
xnor UO_3023 (O_3023,N_29061,N_29059);
or UO_3024 (O_3024,N_29570,N_28436);
or UO_3025 (O_3025,N_29545,N_29810);
or UO_3026 (O_3026,N_29113,N_29204);
nand UO_3027 (O_3027,N_28824,N_28382);
xnor UO_3028 (O_3028,N_29895,N_28129);
nor UO_3029 (O_3029,N_29338,N_28928);
nor UO_3030 (O_3030,N_29168,N_29191);
nand UO_3031 (O_3031,N_28063,N_29176);
or UO_3032 (O_3032,N_29064,N_29900);
nand UO_3033 (O_3033,N_28924,N_29223);
nor UO_3034 (O_3034,N_29882,N_28366);
nor UO_3035 (O_3035,N_29944,N_28964);
and UO_3036 (O_3036,N_29803,N_29402);
xnor UO_3037 (O_3037,N_29785,N_28167);
or UO_3038 (O_3038,N_28580,N_29777);
nor UO_3039 (O_3039,N_29781,N_28085);
xnor UO_3040 (O_3040,N_29677,N_28109);
nor UO_3041 (O_3041,N_28782,N_28949);
or UO_3042 (O_3042,N_28762,N_29885);
and UO_3043 (O_3043,N_28676,N_29679);
or UO_3044 (O_3044,N_28483,N_28166);
and UO_3045 (O_3045,N_29438,N_29446);
and UO_3046 (O_3046,N_29233,N_28343);
and UO_3047 (O_3047,N_29942,N_28751);
xor UO_3048 (O_3048,N_28841,N_28051);
xor UO_3049 (O_3049,N_28118,N_28279);
or UO_3050 (O_3050,N_29693,N_29883);
and UO_3051 (O_3051,N_28249,N_29479);
or UO_3052 (O_3052,N_29401,N_29713);
or UO_3053 (O_3053,N_29685,N_29103);
and UO_3054 (O_3054,N_28560,N_29378);
xor UO_3055 (O_3055,N_28239,N_28227);
or UO_3056 (O_3056,N_28224,N_29202);
xnor UO_3057 (O_3057,N_29555,N_28400);
xnor UO_3058 (O_3058,N_29486,N_28776);
and UO_3059 (O_3059,N_28306,N_28455);
nor UO_3060 (O_3060,N_29896,N_29418);
or UO_3061 (O_3061,N_29394,N_29110);
and UO_3062 (O_3062,N_29409,N_29467);
and UO_3063 (O_3063,N_28622,N_29886);
and UO_3064 (O_3064,N_29860,N_29570);
nand UO_3065 (O_3065,N_29602,N_29475);
nor UO_3066 (O_3066,N_29345,N_28805);
nand UO_3067 (O_3067,N_29907,N_29826);
xor UO_3068 (O_3068,N_28262,N_29735);
xor UO_3069 (O_3069,N_28515,N_29057);
nand UO_3070 (O_3070,N_28741,N_28906);
nand UO_3071 (O_3071,N_28493,N_28170);
or UO_3072 (O_3072,N_29681,N_28375);
and UO_3073 (O_3073,N_28740,N_28885);
and UO_3074 (O_3074,N_28448,N_28560);
xnor UO_3075 (O_3075,N_29851,N_29782);
nor UO_3076 (O_3076,N_29286,N_29535);
xor UO_3077 (O_3077,N_28738,N_29119);
nand UO_3078 (O_3078,N_29372,N_28554);
and UO_3079 (O_3079,N_28395,N_28942);
and UO_3080 (O_3080,N_28739,N_29631);
nand UO_3081 (O_3081,N_28797,N_28710);
nand UO_3082 (O_3082,N_28146,N_29837);
or UO_3083 (O_3083,N_29081,N_28154);
xnor UO_3084 (O_3084,N_28343,N_29034);
or UO_3085 (O_3085,N_28600,N_28844);
and UO_3086 (O_3086,N_28806,N_29865);
nand UO_3087 (O_3087,N_28157,N_28316);
nor UO_3088 (O_3088,N_28664,N_28106);
xor UO_3089 (O_3089,N_28266,N_29216);
or UO_3090 (O_3090,N_29834,N_29698);
and UO_3091 (O_3091,N_29174,N_29001);
and UO_3092 (O_3092,N_29805,N_28161);
xnor UO_3093 (O_3093,N_28027,N_29026);
xnor UO_3094 (O_3094,N_29768,N_28383);
xnor UO_3095 (O_3095,N_28242,N_29207);
nor UO_3096 (O_3096,N_29060,N_28443);
and UO_3097 (O_3097,N_28281,N_29959);
nor UO_3098 (O_3098,N_28874,N_29911);
and UO_3099 (O_3099,N_29197,N_29611);
nand UO_3100 (O_3100,N_28870,N_29427);
nor UO_3101 (O_3101,N_29575,N_29882);
or UO_3102 (O_3102,N_28866,N_29179);
or UO_3103 (O_3103,N_28368,N_28157);
nor UO_3104 (O_3104,N_28435,N_29052);
nand UO_3105 (O_3105,N_29173,N_29223);
nor UO_3106 (O_3106,N_29034,N_29388);
nor UO_3107 (O_3107,N_29853,N_28314);
nor UO_3108 (O_3108,N_28301,N_28823);
and UO_3109 (O_3109,N_28344,N_29383);
nor UO_3110 (O_3110,N_29382,N_28308);
nor UO_3111 (O_3111,N_29091,N_28792);
or UO_3112 (O_3112,N_29854,N_29408);
or UO_3113 (O_3113,N_28693,N_29435);
xnor UO_3114 (O_3114,N_28845,N_28596);
xnor UO_3115 (O_3115,N_28137,N_28776);
and UO_3116 (O_3116,N_28437,N_29715);
xnor UO_3117 (O_3117,N_28264,N_29171);
and UO_3118 (O_3118,N_29780,N_28798);
and UO_3119 (O_3119,N_29348,N_29251);
nand UO_3120 (O_3120,N_29396,N_29830);
nor UO_3121 (O_3121,N_28852,N_28461);
xor UO_3122 (O_3122,N_28323,N_28934);
xor UO_3123 (O_3123,N_29793,N_28324);
nor UO_3124 (O_3124,N_29659,N_28372);
nor UO_3125 (O_3125,N_28707,N_29380);
nor UO_3126 (O_3126,N_29617,N_29949);
or UO_3127 (O_3127,N_29778,N_28185);
xnor UO_3128 (O_3128,N_28970,N_29025);
nor UO_3129 (O_3129,N_28293,N_28783);
xnor UO_3130 (O_3130,N_29812,N_29043);
and UO_3131 (O_3131,N_29277,N_29260);
nor UO_3132 (O_3132,N_29855,N_29319);
and UO_3133 (O_3133,N_28360,N_29344);
nand UO_3134 (O_3134,N_29815,N_28262);
and UO_3135 (O_3135,N_28222,N_28011);
or UO_3136 (O_3136,N_28118,N_29034);
and UO_3137 (O_3137,N_28506,N_28078);
nand UO_3138 (O_3138,N_29974,N_28173);
or UO_3139 (O_3139,N_29873,N_29482);
nor UO_3140 (O_3140,N_28480,N_28942);
nor UO_3141 (O_3141,N_28755,N_28557);
and UO_3142 (O_3142,N_28613,N_29785);
nand UO_3143 (O_3143,N_28825,N_28334);
nand UO_3144 (O_3144,N_28222,N_29844);
nor UO_3145 (O_3145,N_28724,N_29097);
nor UO_3146 (O_3146,N_29585,N_28998);
xnor UO_3147 (O_3147,N_29719,N_28162);
nand UO_3148 (O_3148,N_28987,N_29179);
xnor UO_3149 (O_3149,N_28681,N_29593);
and UO_3150 (O_3150,N_29236,N_28215);
and UO_3151 (O_3151,N_28960,N_28451);
or UO_3152 (O_3152,N_28385,N_28752);
xnor UO_3153 (O_3153,N_29025,N_29145);
or UO_3154 (O_3154,N_29479,N_28733);
nor UO_3155 (O_3155,N_28324,N_28775);
nor UO_3156 (O_3156,N_28631,N_28929);
and UO_3157 (O_3157,N_29037,N_28888);
nor UO_3158 (O_3158,N_29963,N_29188);
xnor UO_3159 (O_3159,N_28886,N_28432);
xnor UO_3160 (O_3160,N_28166,N_28900);
and UO_3161 (O_3161,N_28523,N_29502);
nor UO_3162 (O_3162,N_29984,N_29927);
or UO_3163 (O_3163,N_29667,N_28427);
nor UO_3164 (O_3164,N_29658,N_28960);
nand UO_3165 (O_3165,N_29216,N_28022);
nor UO_3166 (O_3166,N_29592,N_29367);
nand UO_3167 (O_3167,N_28674,N_29461);
or UO_3168 (O_3168,N_29051,N_28366);
or UO_3169 (O_3169,N_29966,N_28669);
and UO_3170 (O_3170,N_29326,N_28695);
xor UO_3171 (O_3171,N_29892,N_29535);
or UO_3172 (O_3172,N_28624,N_29405);
xnor UO_3173 (O_3173,N_29948,N_28835);
and UO_3174 (O_3174,N_28478,N_28527);
and UO_3175 (O_3175,N_28874,N_29293);
xor UO_3176 (O_3176,N_29915,N_29434);
and UO_3177 (O_3177,N_28640,N_29207);
xnor UO_3178 (O_3178,N_28010,N_29488);
or UO_3179 (O_3179,N_28275,N_29162);
nand UO_3180 (O_3180,N_29579,N_29055);
nor UO_3181 (O_3181,N_28999,N_28003);
nand UO_3182 (O_3182,N_29843,N_29021);
xor UO_3183 (O_3183,N_29250,N_28504);
nand UO_3184 (O_3184,N_29224,N_28765);
and UO_3185 (O_3185,N_29044,N_28326);
xnor UO_3186 (O_3186,N_28353,N_29017);
xnor UO_3187 (O_3187,N_28105,N_29498);
nand UO_3188 (O_3188,N_29364,N_29224);
or UO_3189 (O_3189,N_28842,N_29659);
nor UO_3190 (O_3190,N_29529,N_28827);
xnor UO_3191 (O_3191,N_29675,N_28438);
and UO_3192 (O_3192,N_29948,N_28537);
or UO_3193 (O_3193,N_28254,N_29993);
nor UO_3194 (O_3194,N_29367,N_28902);
xor UO_3195 (O_3195,N_29478,N_28272);
nand UO_3196 (O_3196,N_28770,N_29334);
nor UO_3197 (O_3197,N_29631,N_29731);
nor UO_3198 (O_3198,N_28196,N_29287);
or UO_3199 (O_3199,N_28891,N_28583);
or UO_3200 (O_3200,N_29625,N_28534);
and UO_3201 (O_3201,N_29472,N_28505);
xor UO_3202 (O_3202,N_29493,N_28901);
nand UO_3203 (O_3203,N_28723,N_29189);
nand UO_3204 (O_3204,N_29082,N_28043);
nor UO_3205 (O_3205,N_28337,N_29080);
or UO_3206 (O_3206,N_29050,N_29180);
and UO_3207 (O_3207,N_29262,N_29959);
nand UO_3208 (O_3208,N_29870,N_28364);
or UO_3209 (O_3209,N_28774,N_28118);
xnor UO_3210 (O_3210,N_28305,N_28863);
xor UO_3211 (O_3211,N_28210,N_28277);
and UO_3212 (O_3212,N_28896,N_28337);
nand UO_3213 (O_3213,N_29498,N_28020);
or UO_3214 (O_3214,N_29860,N_28036);
nor UO_3215 (O_3215,N_28252,N_29579);
nor UO_3216 (O_3216,N_28798,N_28909);
nor UO_3217 (O_3217,N_29514,N_29413);
nand UO_3218 (O_3218,N_28834,N_28722);
and UO_3219 (O_3219,N_29436,N_29761);
nand UO_3220 (O_3220,N_28860,N_29601);
nand UO_3221 (O_3221,N_29522,N_28343);
nand UO_3222 (O_3222,N_28631,N_29045);
nor UO_3223 (O_3223,N_29559,N_28541);
or UO_3224 (O_3224,N_29366,N_29674);
or UO_3225 (O_3225,N_28461,N_28371);
nand UO_3226 (O_3226,N_29495,N_28528);
xnor UO_3227 (O_3227,N_28446,N_29123);
and UO_3228 (O_3228,N_28118,N_29772);
nand UO_3229 (O_3229,N_28508,N_28153);
nand UO_3230 (O_3230,N_29344,N_28518);
nor UO_3231 (O_3231,N_28866,N_29623);
nor UO_3232 (O_3232,N_29738,N_28469);
and UO_3233 (O_3233,N_29500,N_29315);
nand UO_3234 (O_3234,N_28976,N_28347);
xor UO_3235 (O_3235,N_28023,N_29083);
nor UO_3236 (O_3236,N_28062,N_29076);
nor UO_3237 (O_3237,N_28222,N_29628);
nand UO_3238 (O_3238,N_29209,N_29508);
nand UO_3239 (O_3239,N_29704,N_28683);
nand UO_3240 (O_3240,N_29182,N_29852);
nor UO_3241 (O_3241,N_29287,N_29326);
nand UO_3242 (O_3242,N_29164,N_28774);
xor UO_3243 (O_3243,N_28580,N_28581);
xnor UO_3244 (O_3244,N_29044,N_29580);
nand UO_3245 (O_3245,N_28689,N_29162);
or UO_3246 (O_3246,N_28768,N_28327);
nor UO_3247 (O_3247,N_29465,N_29024);
xnor UO_3248 (O_3248,N_29279,N_28950);
and UO_3249 (O_3249,N_29642,N_28320);
and UO_3250 (O_3250,N_29602,N_28869);
or UO_3251 (O_3251,N_29341,N_29182);
nand UO_3252 (O_3252,N_29791,N_29147);
or UO_3253 (O_3253,N_28363,N_29435);
and UO_3254 (O_3254,N_29419,N_29540);
and UO_3255 (O_3255,N_28258,N_28143);
and UO_3256 (O_3256,N_28158,N_28573);
nand UO_3257 (O_3257,N_28778,N_28864);
and UO_3258 (O_3258,N_29012,N_29981);
nand UO_3259 (O_3259,N_28057,N_29713);
or UO_3260 (O_3260,N_28557,N_29313);
xnor UO_3261 (O_3261,N_29447,N_29650);
nand UO_3262 (O_3262,N_29059,N_29967);
xnor UO_3263 (O_3263,N_28150,N_28918);
xor UO_3264 (O_3264,N_29503,N_29644);
and UO_3265 (O_3265,N_28785,N_28073);
xor UO_3266 (O_3266,N_28896,N_28257);
nor UO_3267 (O_3267,N_28274,N_29542);
xor UO_3268 (O_3268,N_28622,N_28955);
or UO_3269 (O_3269,N_28118,N_29324);
xnor UO_3270 (O_3270,N_28611,N_29344);
xnor UO_3271 (O_3271,N_28896,N_29251);
nor UO_3272 (O_3272,N_29378,N_28958);
or UO_3273 (O_3273,N_28643,N_29753);
and UO_3274 (O_3274,N_28987,N_29274);
or UO_3275 (O_3275,N_29449,N_28690);
nor UO_3276 (O_3276,N_29512,N_29801);
or UO_3277 (O_3277,N_29326,N_29766);
and UO_3278 (O_3278,N_28170,N_29249);
nand UO_3279 (O_3279,N_29566,N_29236);
nand UO_3280 (O_3280,N_28889,N_28211);
nand UO_3281 (O_3281,N_28264,N_29730);
and UO_3282 (O_3282,N_28421,N_29804);
nand UO_3283 (O_3283,N_29268,N_28030);
and UO_3284 (O_3284,N_29145,N_28268);
or UO_3285 (O_3285,N_29278,N_29398);
or UO_3286 (O_3286,N_29605,N_29282);
nor UO_3287 (O_3287,N_29643,N_29157);
nand UO_3288 (O_3288,N_29371,N_29474);
or UO_3289 (O_3289,N_28955,N_29795);
or UO_3290 (O_3290,N_28663,N_29609);
nand UO_3291 (O_3291,N_29212,N_28574);
xor UO_3292 (O_3292,N_29579,N_29995);
or UO_3293 (O_3293,N_29609,N_28954);
or UO_3294 (O_3294,N_28969,N_28206);
nand UO_3295 (O_3295,N_29467,N_28505);
nor UO_3296 (O_3296,N_29229,N_28938);
nor UO_3297 (O_3297,N_29565,N_29850);
nor UO_3298 (O_3298,N_29402,N_28189);
and UO_3299 (O_3299,N_29289,N_29351);
and UO_3300 (O_3300,N_28556,N_28603);
nand UO_3301 (O_3301,N_28365,N_29849);
xor UO_3302 (O_3302,N_28622,N_28870);
or UO_3303 (O_3303,N_29293,N_28569);
xor UO_3304 (O_3304,N_28406,N_29939);
nor UO_3305 (O_3305,N_29658,N_28525);
and UO_3306 (O_3306,N_29751,N_29856);
nand UO_3307 (O_3307,N_28162,N_29642);
and UO_3308 (O_3308,N_28643,N_28764);
nor UO_3309 (O_3309,N_28009,N_29141);
and UO_3310 (O_3310,N_29969,N_29270);
or UO_3311 (O_3311,N_29082,N_28263);
nand UO_3312 (O_3312,N_29522,N_28202);
xnor UO_3313 (O_3313,N_28263,N_29298);
and UO_3314 (O_3314,N_29937,N_28352);
nand UO_3315 (O_3315,N_28133,N_28263);
xnor UO_3316 (O_3316,N_29085,N_28735);
or UO_3317 (O_3317,N_28068,N_29971);
and UO_3318 (O_3318,N_28994,N_29316);
xor UO_3319 (O_3319,N_29787,N_29944);
nor UO_3320 (O_3320,N_28897,N_29352);
xor UO_3321 (O_3321,N_29595,N_29161);
xor UO_3322 (O_3322,N_29007,N_29783);
nand UO_3323 (O_3323,N_29193,N_29095);
or UO_3324 (O_3324,N_28293,N_28677);
nor UO_3325 (O_3325,N_28302,N_29218);
nand UO_3326 (O_3326,N_29452,N_28522);
nand UO_3327 (O_3327,N_29846,N_29876);
or UO_3328 (O_3328,N_29832,N_28369);
nand UO_3329 (O_3329,N_29757,N_28837);
or UO_3330 (O_3330,N_28940,N_29665);
nand UO_3331 (O_3331,N_28963,N_29167);
or UO_3332 (O_3332,N_29294,N_28129);
or UO_3333 (O_3333,N_28561,N_28311);
and UO_3334 (O_3334,N_28042,N_28275);
xnor UO_3335 (O_3335,N_29659,N_29141);
or UO_3336 (O_3336,N_28595,N_28223);
nand UO_3337 (O_3337,N_28355,N_29088);
nand UO_3338 (O_3338,N_28789,N_28197);
nor UO_3339 (O_3339,N_28718,N_29796);
or UO_3340 (O_3340,N_28810,N_28053);
nand UO_3341 (O_3341,N_28766,N_29973);
nor UO_3342 (O_3342,N_29973,N_28134);
nand UO_3343 (O_3343,N_29571,N_28362);
nor UO_3344 (O_3344,N_28822,N_29886);
nor UO_3345 (O_3345,N_29420,N_29254);
nor UO_3346 (O_3346,N_28382,N_28894);
or UO_3347 (O_3347,N_28465,N_28508);
xor UO_3348 (O_3348,N_28188,N_28146);
and UO_3349 (O_3349,N_29539,N_28392);
nand UO_3350 (O_3350,N_29772,N_29904);
nand UO_3351 (O_3351,N_28635,N_28229);
xnor UO_3352 (O_3352,N_29092,N_28191);
nor UO_3353 (O_3353,N_28337,N_28363);
xor UO_3354 (O_3354,N_29165,N_29689);
nor UO_3355 (O_3355,N_28158,N_29415);
or UO_3356 (O_3356,N_28200,N_28798);
and UO_3357 (O_3357,N_28122,N_28779);
and UO_3358 (O_3358,N_29224,N_28968);
or UO_3359 (O_3359,N_28910,N_28215);
and UO_3360 (O_3360,N_28505,N_29434);
xnor UO_3361 (O_3361,N_28997,N_28226);
or UO_3362 (O_3362,N_29310,N_29719);
xnor UO_3363 (O_3363,N_29086,N_29075);
nor UO_3364 (O_3364,N_28347,N_28189);
nor UO_3365 (O_3365,N_29851,N_28944);
nand UO_3366 (O_3366,N_28415,N_29817);
or UO_3367 (O_3367,N_28856,N_28096);
nor UO_3368 (O_3368,N_29217,N_29076);
xor UO_3369 (O_3369,N_28216,N_29756);
xnor UO_3370 (O_3370,N_29449,N_29663);
and UO_3371 (O_3371,N_29269,N_29895);
or UO_3372 (O_3372,N_29829,N_28500);
or UO_3373 (O_3373,N_28730,N_28777);
or UO_3374 (O_3374,N_29069,N_29827);
and UO_3375 (O_3375,N_29767,N_28862);
and UO_3376 (O_3376,N_28670,N_29134);
xnor UO_3377 (O_3377,N_28035,N_28022);
and UO_3378 (O_3378,N_29144,N_29024);
xnor UO_3379 (O_3379,N_29160,N_28290);
or UO_3380 (O_3380,N_28605,N_28422);
or UO_3381 (O_3381,N_29848,N_28360);
and UO_3382 (O_3382,N_28728,N_29319);
nor UO_3383 (O_3383,N_28897,N_28598);
nand UO_3384 (O_3384,N_29533,N_28124);
and UO_3385 (O_3385,N_29773,N_28993);
xor UO_3386 (O_3386,N_28238,N_29300);
and UO_3387 (O_3387,N_29230,N_28104);
and UO_3388 (O_3388,N_29234,N_28464);
nor UO_3389 (O_3389,N_28555,N_28388);
nand UO_3390 (O_3390,N_28792,N_29038);
nor UO_3391 (O_3391,N_28571,N_29764);
and UO_3392 (O_3392,N_29255,N_28269);
and UO_3393 (O_3393,N_28054,N_29462);
and UO_3394 (O_3394,N_28501,N_29638);
and UO_3395 (O_3395,N_29305,N_28221);
xnor UO_3396 (O_3396,N_28766,N_28155);
and UO_3397 (O_3397,N_29270,N_28743);
nor UO_3398 (O_3398,N_29245,N_28950);
or UO_3399 (O_3399,N_28433,N_28261);
nor UO_3400 (O_3400,N_28781,N_29868);
and UO_3401 (O_3401,N_28672,N_28112);
or UO_3402 (O_3402,N_28692,N_29147);
and UO_3403 (O_3403,N_29746,N_28943);
or UO_3404 (O_3404,N_29147,N_28357);
or UO_3405 (O_3405,N_28454,N_28725);
nor UO_3406 (O_3406,N_29382,N_28333);
nand UO_3407 (O_3407,N_28987,N_28020);
nor UO_3408 (O_3408,N_28233,N_29689);
xnor UO_3409 (O_3409,N_28859,N_29821);
xor UO_3410 (O_3410,N_28432,N_28551);
nor UO_3411 (O_3411,N_29578,N_28795);
nor UO_3412 (O_3412,N_28980,N_28927);
nor UO_3413 (O_3413,N_28430,N_28241);
and UO_3414 (O_3414,N_29055,N_29052);
and UO_3415 (O_3415,N_28433,N_28647);
xor UO_3416 (O_3416,N_29012,N_29006);
and UO_3417 (O_3417,N_28807,N_29055);
nand UO_3418 (O_3418,N_29449,N_29044);
nor UO_3419 (O_3419,N_29533,N_28994);
xnor UO_3420 (O_3420,N_29736,N_28644);
nand UO_3421 (O_3421,N_29639,N_28260);
or UO_3422 (O_3422,N_28886,N_28908);
xor UO_3423 (O_3423,N_28581,N_28024);
nand UO_3424 (O_3424,N_28505,N_29443);
nor UO_3425 (O_3425,N_28073,N_28205);
or UO_3426 (O_3426,N_29777,N_28750);
or UO_3427 (O_3427,N_28941,N_29864);
xnor UO_3428 (O_3428,N_29627,N_28599);
or UO_3429 (O_3429,N_29344,N_28389);
or UO_3430 (O_3430,N_28422,N_29024);
xnor UO_3431 (O_3431,N_29906,N_29284);
and UO_3432 (O_3432,N_29824,N_29761);
nand UO_3433 (O_3433,N_28372,N_28275);
nor UO_3434 (O_3434,N_29921,N_28679);
xor UO_3435 (O_3435,N_29807,N_28016);
nor UO_3436 (O_3436,N_29651,N_29788);
xnor UO_3437 (O_3437,N_29580,N_29878);
or UO_3438 (O_3438,N_29538,N_29916);
nand UO_3439 (O_3439,N_28266,N_28968);
nor UO_3440 (O_3440,N_28848,N_29763);
nand UO_3441 (O_3441,N_28024,N_28417);
nand UO_3442 (O_3442,N_29530,N_28462);
xor UO_3443 (O_3443,N_29495,N_28890);
xor UO_3444 (O_3444,N_29729,N_28746);
nand UO_3445 (O_3445,N_28653,N_29906);
nand UO_3446 (O_3446,N_28794,N_29601);
and UO_3447 (O_3447,N_28563,N_28338);
nand UO_3448 (O_3448,N_28085,N_29276);
nand UO_3449 (O_3449,N_29671,N_28172);
and UO_3450 (O_3450,N_28997,N_29890);
nor UO_3451 (O_3451,N_29561,N_29806);
or UO_3452 (O_3452,N_29473,N_29955);
nor UO_3453 (O_3453,N_29268,N_28461);
nor UO_3454 (O_3454,N_28962,N_28265);
or UO_3455 (O_3455,N_28500,N_28812);
and UO_3456 (O_3456,N_29678,N_28272);
nand UO_3457 (O_3457,N_29252,N_28415);
nand UO_3458 (O_3458,N_29791,N_29615);
nand UO_3459 (O_3459,N_28285,N_29222);
and UO_3460 (O_3460,N_28584,N_28413);
nand UO_3461 (O_3461,N_29199,N_29651);
nand UO_3462 (O_3462,N_28323,N_28409);
nand UO_3463 (O_3463,N_29498,N_28368);
nor UO_3464 (O_3464,N_28245,N_28580);
nor UO_3465 (O_3465,N_28840,N_28565);
and UO_3466 (O_3466,N_28161,N_28811);
nor UO_3467 (O_3467,N_29117,N_29623);
nor UO_3468 (O_3468,N_29097,N_29275);
xor UO_3469 (O_3469,N_28517,N_29232);
and UO_3470 (O_3470,N_28732,N_29806);
or UO_3471 (O_3471,N_28205,N_29829);
xor UO_3472 (O_3472,N_29022,N_29510);
and UO_3473 (O_3473,N_28093,N_28736);
nand UO_3474 (O_3474,N_29767,N_29112);
nor UO_3475 (O_3475,N_29496,N_29057);
and UO_3476 (O_3476,N_29398,N_28045);
nand UO_3477 (O_3477,N_29988,N_28341);
and UO_3478 (O_3478,N_28230,N_28811);
xor UO_3479 (O_3479,N_29090,N_28170);
and UO_3480 (O_3480,N_28836,N_29955);
or UO_3481 (O_3481,N_29006,N_29797);
nor UO_3482 (O_3482,N_28231,N_29449);
or UO_3483 (O_3483,N_28933,N_29495);
or UO_3484 (O_3484,N_28489,N_29153);
or UO_3485 (O_3485,N_29709,N_29783);
or UO_3486 (O_3486,N_28749,N_29818);
xor UO_3487 (O_3487,N_29439,N_29191);
xnor UO_3488 (O_3488,N_28782,N_28420);
nor UO_3489 (O_3489,N_29622,N_28607);
xor UO_3490 (O_3490,N_28336,N_28243);
and UO_3491 (O_3491,N_29701,N_28994);
and UO_3492 (O_3492,N_28206,N_29293);
nor UO_3493 (O_3493,N_28301,N_29054);
nor UO_3494 (O_3494,N_28309,N_28705);
and UO_3495 (O_3495,N_29879,N_28958);
nand UO_3496 (O_3496,N_29003,N_29074);
nand UO_3497 (O_3497,N_29196,N_29652);
xor UO_3498 (O_3498,N_29867,N_28775);
nand UO_3499 (O_3499,N_29771,N_28959);
endmodule