module basic_1000_10000_1500_50_levels_10xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
and U0 (N_0,In_522,In_803);
or U1 (N_1,In_554,In_760);
xor U2 (N_2,In_514,In_957);
nand U3 (N_3,In_228,In_638);
nand U4 (N_4,In_537,In_177);
nand U5 (N_5,In_26,In_156);
and U6 (N_6,In_233,In_317);
xnor U7 (N_7,In_257,In_51);
nand U8 (N_8,In_496,In_1);
xor U9 (N_9,In_405,In_446);
or U10 (N_10,In_54,In_139);
nor U11 (N_11,In_936,In_181);
and U12 (N_12,In_856,In_196);
xnor U13 (N_13,In_203,In_289);
and U14 (N_14,In_841,In_650);
nor U15 (N_15,In_999,In_597);
xnor U16 (N_16,In_74,In_690);
or U17 (N_17,In_14,In_86);
nand U18 (N_18,In_98,In_981);
and U19 (N_19,In_832,In_141);
nor U20 (N_20,In_903,In_801);
and U21 (N_21,In_774,In_933);
nor U22 (N_22,In_352,In_818);
or U23 (N_23,In_404,In_288);
nand U24 (N_24,In_114,In_807);
or U25 (N_25,In_299,In_843);
nor U26 (N_26,In_441,In_427);
nand U27 (N_27,In_385,In_886);
or U28 (N_28,In_149,In_872);
and U29 (N_29,In_195,In_244);
nand U30 (N_30,In_173,In_915);
nand U31 (N_31,In_209,In_546);
and U32 (N_32,In_587,In_65);
or U33 (N_33,In_28,In_645);
nand U34 (N_34,In_799,In_32);
or U35 (N_35,In_989,In_563);
nand U36 (N_36,In_392,In_384);
and U37 (N_37,In_855,In_148);
xor U38 (N_38,In_187,In_515);
nor U39 (N_39,In_160,In_730);
nand U40 (N_40,In_953,In_235);
xor U41 (N_41,In_585,In_155);
nor U42 (N_42,In_267,In_30);
nor U43 (N_43,In_866,In_8);
xor U44 (N_44,In_719,In_94);
or U45 (N_45,In_401,In_321);
nor U46 (N_46,In_99,In_363);
nand U47 (N_47,In_6,In_627);
or U48 (N_48,In_746,In_464);
xnor U49 (N_49,In_835,In_613);
nor U50 (N_50,In_101,In_455);
or U51 (N_51,In_10,In_304);
nand U52 (N_52,In_534,In_821);
and U53 (N_53,In_894,In_943);
or U54 (N_54,In_276,In_452);
xor U55 (N_55,In_162,In_833);
xnor U56 (N_56,In_666,In_305);
or U57 (N_57,In_408,In_225);
or U58 (N_58,In_335,In_301);
nand U59 (N_59,In_306,In_701);
and U60 (N_60,In_773,In_967);
xnor U61 (N_61,In_880,In_611);
or U62 (N_62,In_592,In_834);
nand U63 (N_63,In_751,In_247);
and U64 (N_64,In_929,In_593);
or U65 (N_65,In_105,In_179);
nand U66 (N_66,In_813,In_713);
or U67 (N_67,In_223,In_785);
and U68 (N_68,In_75,In_897);
and U69 (N_69,In_448,In_264);
xor U70 (N_70,In_964,In_81);
nand U71 (N_71,In_617,In_126);
and U72 (N_72,In_693,In_874);
nand U73 (N_73,In_870,In_313);
xnor U74 (N_74,In_202,In_914);
or U75 (N_75,In_938,In_493);
and U76 (N_76,In_70,In_579);
nor U77 (N_77,In_351,In_108);
nor U78 (N_78,In_429,In_950);
or U79 (N_79,In_35,In_836);
or U80 (N_80,In_340,In_739);
or U81 (N_81,In_940,In_643);
or U82 (N_82,In_790,In_902);
or U83 (N_83,In_227,In_918);
nand U84 (N_84,In_581,In_922);
nor U85 (N_85,In_413,In_817);
or U86 (N_86,In_814,In_402);
or U87 (N_87,In_256,In_273);
xnor U88 (N_88,In_31,In_987);
and U89 (N_89,In_876,In_649);
nand U90 (N_90,In_596,In_85);
and U91 (N_91,In_703,In_319);
nand U92 (N_92,In_697,In_170);
or U93 (N_93,In_669,In_48);
or U94 (N_94,In_147,In_823);
and U95 (N_95,In_511,In_124);
nand U96 (N_96,In_18,In_711);
xor U97 (N_97,In_186,In_398);
xor U98 (N_98,In_887,In_565);
xnor U99 (N_99,In_95,In_684);
or U100 (N_100,In_143,In_198);
xnor U101 (N_101,In_116,In_38);
or U102 (N_102,In_323,In_702);
nor U103 (N_103,In_419,In_682);
xor U104 (N_104,In_211,In_439);
nand U105 (N_105,In_300,In_412);
and U106 (N_106,In_208,In_549);
xnor U107 (N_107,In_962,In_27);
nor U108 (N_108,In_449,In_42);
xor U109 (N_109,In_142,In_120);
nand U110 (N_110,In_472,In_709);
xnor U111 (N_111,In_517,In_520);
nor U112 (N_112,In_959,In_508);
and U113 (N_113,In_978,In_296);
xnor U114 (N_114,In_111,In_923);
and U115 (N_115,In_793,In_406);
or U116 (N_116,In_62,In_325);
nand U117 (N_117,In_777,In_409);
or U118 (N_118,In_648,In_486);
xor U119 (N_119,In_188,In_373);
xnor U120 (N_120,In_491,In_260);
and U121 (N_121,In_527,In_727);
nor U122 (N_122,In_827,In_91);
or U123 (N_123,In_538,In_524);
nor U124 (N_124,In_258,In_513);
nand U125 (N_125,In_891,In_151);
and U126 (N_126,In_462,In_231);
xnor U127 (N_127,In_47,In_809);
or U128 (N_128,In_55,In_396);
nor U129 (N_129,In_123,In_646);
nor U130 (N_130,In_560,In_459);
or U131 (N_131,In_145,In_780);
xor U132 (N_132,In_368,In_926);
nand U133 (N_133,In_737,In_157);
xnor U134 (N_134,In_311,In_745);
xnor U135 (N_135,In_766,In_292);
nand U136 (N_136,In_970,In_303);
or U137 (N_137,In_348,In_444);
or U138 (N_138,In_440,In_320);
and U139 (N_139,In_61,In_488);
xor U140 (N_140,In_916,In_367);
and U141 (N_141,In_586,In_505);
nand U142 (N_142,In_394,In_115);
xnor U143 (N_143,In_826,In_206);
xnor U144 (N_144,In_269,In_332);
nor U145 (N_145,In_293,In_399);
and U146 (N_146,In_659,In_802);
xnor U147 (N_147,In_677,In_20);
nor U148 (N_148,In_360,In_204);
nand U149 (N_149,In_483,In_316);
and U150 (N_150,In_906,In_954);
nand U151 (N_151,In_469,In_457);
nor U152 (N_152,In_825,In_699);
or U153 (N_153,In_389,In_864);
and U154 (N_154,In_239,In_992);
xor U155 (N_155,In_89,In_49);
and U156 (N_156,In_342,In_536);
nor U157 (N_157,In_327,In_158);
nand U158 (N_158,In_924,In_768);
and U159 (N_159,In_948,In_951);
and U160 (N_160,In_474,In_535);
or U161 (N_161,In_822,In_21);
nor U162 (N_162,In_315,In_657);
or U163 (N_163,In_842,In_16);
xor U164 (N_164,In_84,In_96);
nor U165 (N_165,In_83,In_888);
or U166 (N_166,In_620,In_758);
or U167 (N_167,In_997,In_4);
nand U168 (N_168,In_808,In_285);
nor U169 (N_169,In_278,In_840);
or U170 (N_170,In_770,In_909);
and U171 (N_171,In_0,In_589);
and U172 (N_172,In_336,In_201);
or U173 (N_173,In_45,In_418);
xor U174 (N_174,In_512,In_221);
and U175 (N_175,In_707,In_165);
nor U176 (N_176,In_34,In_584);
xnor U177 (N_177,In_191,In_122);
nand U178 (N_178,In_465,In_744);
nor U179 (N_179,In_460,In_246);
nor U180 (N_180,In_623,In_661);
or U181 (N_181,In_601,In_397);
or U182 (N_182,In_501,In_789);
or U183 (N_183,In_507,In_991);
nor U184 (N_184,In_772,In_717);
nor U185 (N_185,In_495,In_608);
and U186 (N_186,In_686,In_622);
xor U187 (N_187,In_266,In_689);
nand U188 (N_188,In_735,In_467);
or U189 (N_189,In_154,In_607);
or U190 (N_190,In_656,In_761);
xnor U191 (N_191,In_376,In_639);
and U192 (N_192,In_787,In_757);
and U193 (N_193,In_629,In_831);
or U194 (N_194,In_605,In_574);
or U195 (N_195,In_243,In_355);
or U196 (N_196,In_456,In_844);
nor U197 (N_197,In_961,In_539);
nor U198 (N_198,In_113,In_334);
or U199 (N_199,In_271,In_810);
and U200 (N_200,In_982,In_988);
xnor U201 (N_201,In_947,In_420);
xnor U202 (N_202,In_80,In_900);
nor U203 (N_203,In_281,In_310);
nor U204 (N_204,In_566,In_850);
or U205 (N_205,In_700,In_721);
nor U206 (N_206,In_265,In_109);
xor U207 (N_207,In_354,In_272);
and U208 (N_208,In_185,N_92);
xnor U209 (N_209,N_3,N_10);
xor U210 (N_210,N_29,In_561);
or U211 (N_211,In_58,N_23);
nor U212 (N_212,In_287,N_15);
and U213 (N_213,In_286,In_482);
and U214 (N_214,In_696,N_170);
nor U215 (N_215,In_580,N_14);
nor U216 (N_216,In_338,N_24);
nand U217 (N_217,In_447,In_131);
nand U218 (N_218,N_123,In_477);
xnor U219 (N_219,In_578,In_540);
and U220 (N_220,In_740,N_155);
nand U221 (N_221,N_62,In_952);
nor U222 (N_222,In_125,N_192);
xnor U223 (N_223,N_103,In_350);
or U224 (N_224,In_956,In_895);
and U225 (N_225,In_358,In_9);
nand U226 (N_226,N_171,In_76);
xor U227 (N_227,In_36,In_224);
xnor U228 (N_228,In_865,In_706);
nand U229 (N_229,In_130,In_283);
and U230 (N_230,N_68,In_741);
and U231 (N_231,In_750,In_450);
and U232 (N_232,In_353,In_734);
nand U233 (N_233,In_972,N_95);
xor U234 (N_234,N_117,In_15);
and U235 (N_235,In_330,N_127);
nor U236 (N_236,In_712,N_80);
nor U237 (N_237,N_73,In_816);
or U238 (N_238,In_309,In_463);
and U239 (N_239,In_907,In_341);
and U240 (N_240,In_322,In_668);
or U241 (N_241,In_971,N_17);
xnor U242 (N_242,In_861,In_410);
and U243 (N_243,In_839,In_797);
or U244 (N_244,In_253,In_205);
nor U245 (N_245,In_528,In_127);
xnor U246 (N_246,In_647,In_254);
nor U247 (N_247,In_913,N_56);
nand U248 (N_248,N_5,N_72);
nor U249 (N_249,N_55,In_974);
xor U250 (N_250,In_270,N_97);
or U251 (N_251,In_983,In_800);
or U252 (N_252,In_945,In_603);
xnor U253 (N_253,N_41,In_103);
nor U254 (N_254,In_97,In_577);
xnor U255 (N_255,In_958,In_868);
or U256 (N_256,In_132,N_30);
or U257 (N_257,In_722,In_718);
and U258 (N_258,In_753,In_949);
xor U259 (N_259,In_532,In_848);
xor U260 (N_260,In_612,In_218);
nor U261 (N_261,In_892,In_297);
xor U262 (N_262,In_64,In_747);
or U263 (N_263,N_38,In_442);
xnor U264 (N_264,N_152,In_133);
and U265 (N_265,In_331,In_625);
and U266 (N_266,N_177,N_193);
and U267 (N_267,N_88,N_11);
nand U268 (N_268,In_849,In_752);
or U269 (N_269,N_142,In_487);
nand U270 (N_270,In_324,In_230);
nand U271 (N_271,In_679,In_588);
and U272 (N_272,In_771,In_912);
nor U273 (N_273,In_19,In_794);
xnor U274 (N_274,In_366,In_937);
or U275 (N_275,In_644,In_628);
nand U276 (N_276,In_518,N_105);
or U277 (N_277,In_599,N_179);
nand U278 (N_278,N_167,In_928);
and U279 (N_279,In_117,In_558);
nor U280 (N_280,N_86,In_615);
nand U281 (N_281,N_115,In_863);
and U282 (N_282,In_635,N_128);
nor U283 (N_283,N_32,In_529);
xnor U284 (N_284,In_33,N_101);
and U285 (N_285,In_87,N_27);
nand U286 (N_286,In_194,In_990);
xnor U287 (N_287,N_185,In_454);
xor U288 (N_288,In_176,In_136);
nand U289 (N_289,N_63,In_678);
nand U290 (N_290,In_234,In_653);
nor U291 (N_291,In_414,In_845);
nor U292 (N_292,In_869,In_370);
and U293 (N_293,In_248,In_343);
nand U294 (N_294,In_621,In_171);
and U295 (N_295,In_238,In_551);
or U296 (N_296,In_371,In_479);
nand U297 (N_297,N_79,N_160);
nand U298 (N_298,N_52,In_640);
nor U299 (N_299,In_798,In_37);
or U300 (N_300,In_365,In_609);
or U301 (N_301,In_180,In_901);
nand U302 (N_302,In_290,In_525);
nand U303 (N_303,In_692,In_106);
nand U304 (N_304,N_118,In_263);
or U305 (N_305,N_191,N_77);
nand U306 (N_306,In_121,N_45);
nor U307 (N_307,In_432,N_106);
nand U308 (N_308,In_393,N_124);
nor U309 (N_309,In_216,In_867);
or U310 (N_310,In_362,In_90);
xor U311 (N_311,In_860,N_132);
or U312 (N_312,N_149,In_875);
nor U313 (N_313,In_382,In_381);
and U314 (N_314,N_50,In_494);
nand U315 (N_315,In_435,N_198);
nand U316 (N_316,In_57,In_328);
nand U317 (N_317,In_553,In_134);
nor U318 (N_318,In_598,In_550);
nor U319 (N_319,In_927,In_889);
nor U320 (N_320,In_968,N_99);
nand U321 (N_321,In_688,In_2);
and U322 (N_322,In_5,In_642);
nor U323 (N_323,In_652,In_544);
xnor U324 (N_324,In_779,In_691);
or U325 (N_325,N_162,In_919);
or U326 (N_326,N_174,In_516);
or U327 (N_327,In_986,In_541);
nand U328 (N_328,In_862,N_18);
and U329 (N_329,In_667,In_161);
nand U330 (N_330,N_102,In_595);
nand U331 (N_331,In_674,In_295);
xnor U332 (N_332,N_20,N_64);
or U333 (N_333,N_25,N_35);
xnor U334 (N_334,In_167,In_425);
and U335 (N_335,In_788,N_175);
xnor U336 (N_336,N_188,In_82);
or U337 (N_337,N_48,In_219);
and U338 (N_338,In_329,In_461);
nor U339 (N_339,In_619,N_57);
or U340 (N_340,N_34,In_931);
nor U341 (N_341,N_98,In_616);
and U342 (N_342,In_391,In_673);
nand U343 (N_343,In_724,In_542);
and U344 (N_344,In_960,In_484);
nand U345 (N_345,N_139,N_137);
xnor U346 (N_346,In_634,In_379);
nor U347 (N_347,In_453,In_128);
nor U348 (N_348,N_65,In_298);
xor U349 (N_349,In_881,N_168);
nand U350 (N_350,In_102,In_655);
nand U351 (N_351,In_434,In_852);
xnor U352 (N_352,N_19,N_156);
nor U353 (N_353,In_557,In_762);
or U354 (N_354,In_359,N_8);
and U355 (N_355,In_458,N_46);
nor U356 (N_356,N_0,In_110);
and U357 (N_357,N_4,In_853);
nor U358 (N_358,N_194,In_307);
or U359 (N_359,In_275,In_476);
nor U360 (N_360,In_498,In_215);
or U361 (N_361,In_944,In_715);
xnor U362 (N_362,N_131,N_12);
and U363 (N_363,In_240,In_159);
or U364 (N_364,In_100,In_344);
nor U365 (N_365,In_291,In_680);
nor U366 (N_366,N_157,N_140);
xor U367 (N_367,In_925,In_795);
nor U368 (N_368,N_116,In_497);
and U369 (N_369,N_164,In_519);
nor U370 (N_370,In_670,In_387);
nor U371 (N_371,In_390,In_873);
xor U372 (N_372,In_998,In_898);
or U373 (N_373,In_626,In_135);
nand U374 (N_374,In_602,N_113);
xnor U375 (N_375,N_154,N_189);
nor U376 (N_376,In_312,N_58);
and U377 (N_377,In_314,In_259);
or U378 (N_378,N_83,In_641);
and U379 (N_379,In_164,In_778);
nand U380 (N_380,In_478,N_85);
nand U381 (N_381,In_52,In_658);
xor U382 (N_382,In_857,In_792);
nor U383 (N_383,In_470,N_176);
and U384 (N_384,In_610,N_40);
and U385 (N_385,In_431,In_896);
or U386 (N_386,N_74,In_78);
xnor U387 (N_387,In_731,N_104);
nor U388 (N_388,In_729,In_197);
xnor U389 (N_389,N_197,In_904);
nand U390 (N_390,In_965,In_473);
and U391 (N_391,In_72,N_2);
and U392 (N_392,In_153,In_226);
xnor U393 (N_393,N_133,N_126);
nand U394 (N_394,N_114,In_437);
or U395 (N_395,In_805,In_262);
or U396 (N_396,In_252,In_533);
nand U397 (N_397,In_137,In_490);
or U398 (N_398,In_436,In_631);
nor U399 (N_399,In_250,N_61);
nor U400 (N_400,In_973,N_130);
nand U401 (N_401,N_223,In_725);
nand U402 (N_402,In_294,In_879);
nand U403 (N_403,In_786,In_502);
nand U404 (N_404,In_166,In_764);
and U405 (N_405,In_407,N_363);
xor U406 (N_406,In_783,N_323);
or U407 (N_407,N_166,In_976);
nor U408 (N_408,In_993,In_44);
or U409 (N_409,In_893,N_276);
and U410 (N_410,In_877,In_590);
nor U411 (N_411,In_88,In_675);
and U412 (N_412,N_42,In_665);
or U413 (N_413,In_720,N_390);
xor U414 (N_414,In_468,In_884);
xor U415 (N_415,N_329,N_314);
and U416 (N_416,In_743,N_312);
and U417 (N_417,N_247,In_73);
and U418 (N_418,N_22,N_87);
xor U419 (N_419,N_237,N_373);
nand U420 (N_420,In_765,N_272);
and U421 (N_421,In_480,In_280);
nand U422 (N_422,In_146,N_364);
xnor U423 (N_423,N_275,In_383);
and U424 (N_424,In_733,N_393);
nand U425 (N_425,In_521,N_251);
and U426 (N_426,N_200,N_235);
and U427 (N_427,In_356,In_630);
nand U428 (N_428,In_624,In_29);
or U429 (N_429,In_796,In_213);
or U430 (N_430,N_357,In_985);
or U431 (N_431,In_506,In_636);
and U432 (N_432,N_75,N_16);
nand U433 (N_433,In_403,N_47);
or U434 (N_434,In_885,In_339);
xor U435 (N_435,N_362,In_582);
or U436 (N_436,In_77,N_301);
xor U437 (N_437,In_7,In_828);
xnor U438 (N_438,N_354,N_266);
xnor U439 (N_439,In_284,N_350);
xnor U440 (N_440,In_749,N_144);
or U441 (N_441,N_248,In_984);
xnor U442 (N_442,In_921,N_333);
xor U443 (N_443,N_108,In_169);
and U444 (N_444,In_614,N_136);
nor U445 (N_445,N_293,N_280);
nand U446 (N_446,N_250,N_243);
and U447 (N_447,N_383,N_7);
xnor U448 (N_448,N_297,N_330);
xor U449 (N_449,N_263,N_6);
or U450 (N_450,N_26,N_328);
and U451 (N_451,N_135,In_104);
xor U452 (N_452,N_343,In_489);
nand U453 (N_453,In_955,In_651);
nor U454 (N_454,N_360,N_145);
nand U455 (N_455,N_228,N_305);
or U456 (N_456,In_975,N_273);
nor U457 (N_457,N_110,In_979);
nand U458 (N_458,In_775,In_941);
and U459 (N_459,N_112,In_261);
nand U460 (N_460,In_564,In_129);
nand U461 (N_461,N_1,In_302);
or U462 (N_462,N_163,In_504);
and U463 (N_463,N_359,In_911);
and U464 (N_464,N_159,In_871);
nand U465 (N_465,N_107,In_934);
nand U466 (N_466,N_396,In_144);
nand U467 (N_467,In_830,In_910);
or U468 (N_468,N_219,N_349);
xor U469 (N_469,In_424,N_84);
or U470 (N_470,N_286,In_308);
nor U471 (N_471,N_324,In_274);
or U472 (N_472,N_143,In_676);
nand U473 (N_473,N_299,In_806);
and U474 (N_474,N_208,N_378);
nor U475 (N_475,N_391,In_172);
and U476 (N_476,In_175,In_43);
xnor U477 (N_477,In_333,In_672);
nor U478 (N_478,In_178,N_224);
xor U479 (N_479,In_683,N_180);
or U480 (N_480,In_25,N_211);
nor U481 (N_481,In_769,N_220);
nand U482 (N_482,N_325,N_303);
nor U483 (N_483,N_308,N_204);
nand U484 (N_484,In_68,In_59);
and U485 (N_485,In_698,N_183);
nor U486 (N_486,N_147,N_173);
xnor U487 (N_487,In_694,N_379);
nor U488 (N_488,In_13,N_181);
or U489 (N_489,N_311,N_31);
xnor U490 (N_490,In_168,In_428);
xor U491 (N_491,In_229,N_397);
xnor U492 (N_492,N_317,In_966);
nand U493 (N_493,N_399,N_212);
nor U494 (N_494,N_196,In_212);
nor U495 (N_495,In_107,In_245);
nand U496 (N_496,N_229,N_240);
xnor U497 (N_497,N_199,N_218);
nand U498 (N_498,In_776,In_687);
or U499 (N_499,N_146,In_222);
or U500 (N_500,In_236,N_277);
or U501 (N_501,In_681,In_503);
and U502 (N_502,In_374,N_331);
or U503 (N_503,In_996,N_216);
nand U504 (N_504,In_633,N_388);
and U505 (N_505,N_316,In_346);
or U506 (N_506,N_71,N_375);
nand U507 (N_507,In_695,N_366);
nor U508 (N_508,N_256,N_234);
xnor U509 (N_509,N_122,N_81);
or U510 (N_510,N_292,In_485);
and U511 (N_511,In_451,N_341);
or U512 (N_512,In_812,In_547);
nor U513 (N_513,In_251,N_239);
and U514 (N_514,In_569,In_531);
or U515 (N_515,In_364,N_288);
xnor U516 (N_516,N_213,N_54);
or U517 (N_517,N_355,In_23);
nor U518 (N_518,N_368,N_353);
or U519 (N_519,In_345,N_285);
nand U520 (N_520,In_69,N_254);
nand U521 (N_521,N_347,In_890);
nor U522 (N_522,In_152,In_811);
xor U523 (N_523,N_258,In_67);
and U524 (N_524,In_930,In_422);
or U525 (N_525,In_255,N_334);
or U526 (N_526,N_182,N_153);
nand U527 (N_527,In_604,In_56);
xnor U528 (N_528,N_96,In_193);
and U529 (N_529,N_66,In_935);
nor U530 (N_530,In_237,In_685);
xor U531 (N_531,N_129,In_475);
nor U532 (N_532,In_784,In_92);
nand U533 (N_533,N_165,N_344);
xor U534 (N_534,In_530,N_207);
and U535 (N_535,In_372,In_883);
or U536 (N_536,In_804,In_138);
and U537 (N_537,In_736,N_270);
xnor U538 (N_538,N_264,N_205);
nand U539 (N_539,N_184,In_548);
and U540 (N_540,In_763,In_782);
nand U541 (N_541,In_543,In_71);
nand U542 (N_542,N_169,N_338);
xor U543 (N_543,N_321,N_195);
or U544 (N_544,In_847,N_214);
xnor U545 (N_545,In_192,In_510);
nand U546 (N_546,N_336,N_309);
nor U547 (N_547,In_199,In_40);
xnor U548 (N_548,In_416,N_315);
or U549 (N_549,N_290,In_710);
nand U550 (N_550,In_671,N_377);
nand U551 (N_551,N_322,N_232);
or U552 (N_552,In_759,In_388);
xor U553 (N_553,In_430,N_342);
nor U554 (N_554,N_60,N_291);
or U555 (N_555,N_253,N_374);
or U556 (N_556,N_382,N_381);
and U557 (N_557,N_365,N_230);
nand U558 (N_558,In_726,In_79);
and U559 (N_559,In_552,N_39);
and U560 (N_560,In_214,N_33);
nor U561 (N_561,In_837,In_46);
nor U562 (N_562,N_318,N_269);
nor U563 (N_563,N_190,N_82);
or U564 (N_564,N_337,In_268);
or U565 (N_565,In_815,In_570);
and U566 (N_566,N_261,N_53);
and U567 (N_567,N_67,In_411);
nand U568 (N_568,In_994,In_562);
xnor U569 (N_569,In_932,N_178);
nand U570 (N_570,N_49,N_300);
xor U571 (N_571,N_231,In_326);
and U572 (N_572,N_36,N_294);
and U573 (N_573,In_663,In_499);
or U574 (N_574,N_120,In_939);
xor U575 (N_575,N_222,In_184);
nand U576 (N_576,In_22,N_367);
and U577 (N_577,N_313,In_977);
or U578 (N_578,In_163,In_748);
nand U579 (N_579,In_545,N_351);
and U580 (N_580,N_59,In_705);
nor U581 (N_581,N_186,In_438);
nand U582 (N_582,N_172,In_732);
nor U583 (N_583,N_209,N_345);
nand U584 (N_584,In_232,In_754);
xor U585 (N_585,N_380,N_262);
nand U586 (N_586,In_357,N_206);
xor U587 (N_587,N_245,N_225);
nand U588 (N_588,In_854,In_41);
nand U589 (N_589,In_708,In_714);
nand U590 (N_590,N_44,In_662);
nor U591 (N_591,In_969,N_283);
xor U592 (N_592,N_91,In_723);
nand U593 (N_593,In_660,In_3);
nor U594 (N_594,In_583,N_242);
or U595 (N_595,N_141,N_265);
xnor U596 (N_596,In_851,In_347);
and U597 (N_597,N_260,In_400);
nor U598 (N_598,In_575,In_728);
and U599 (N_599,N_310,N_51);
nand U600 (N_600,N_492,In_241);
nand U601 (N_601,N_501,N_278);
nor U602 (N_602,N_553,N_566);
and U603 (N_603,N_541,N_412);
or U604 (N_604,N_9,In_654);
nor U605 (N_605,N_557,N_304);
xnor U606 (N_606,N_430,In_11);
xor U607 (N_607,N_417,In_738);
and U608 (N_608,N_451,In_189);
and U609 (N_609,N_407,N_389);
and U610 (N_610,In_426,N_458);
xor U611 (N_611,N_298,N_221);
nand U612 (N_612,N_542,N_533);
and U613 (N_613,In_600,N_543);
xor U614 (N_614,In_572,N_518);
xnor U615 (N_615,N_503,N_570);
nand U616 (N_616,N_431,N_464);
xor U617 (N_617,N_506,N_94);
nor U618 (N_618,N_404,N_497);
and U619 (N_619,N_580,N_480);
xor U620 (N_620,In_878,N_468);
xor U621 (N_621,N_449,N_529);
xnor U622 (N_622,N_527,N_589);
xor U623 (N_623,N_517,In_39);
and U624 (N_624,N_121,In_150);
nor U625 (N_625,N_279,In_443);
nand U626 (N_626,N_462,N_400);
xnor U627 (N_627,In_492,N_282);
nand U628 (N_628,N_394,N_158);
or U629 (N_629,N_448,In_567);
nor U630 (N_630,N_487,N_93);
nand U631 (N_631,N_410,In_838);
or U632 (N_632,N_452,N_403);
or U633 (N_633,N_549,N_461);
and U634 (N_634,In_415,N_528);
nor U635 (N_635,N_13,N_327);
nor U636 (N_636,N_244,N_577);
or U637 (N_637,In_174,N_289);
xor U638 (N_638,N_561,N_320);
nor U639 (N_639,In_17,In_859);
xor U640 (N_640,In_637,In_606);
nor U641 (N_641,N_406,N_583);
and U642 (N_642,In_182,In_781);
and U643 (N_643,N_555,N_556);
xnor U644 (N_644,In_423,In_905);
and U645 (N_645,In_523,N_335);
nand U646 (N_646,N_257,N_525);
xor U647 (N_647,N_210,N_578);
and U648 (N_648,N_586,N_596);
nand U649 (N_649,N_511,N_530);
or U650 (N_650,N_274,N_597);
nor U651 (N_651,In_190,N_476);
and U652 (N_652,N_398,N_405);
nor U653 (N_653,N_238,N_339);
nand U654 (N_654,N_348,In_349);
and U655 (N_655,N_538,N_474);
or U656 (N_656,N_552,N_481);
nand U657 (N_657,In_573,In_632);
nand U658 (N_658,In_755,N_564);
xnor U659 (N_659,N_371,N_493);
nand U660 (N_660,N_361,N_457);
and U661 (N_661,N_500,N_78);
xor U662 (N_662,N_534,In_824);
nor U663 (N_663,N_587,In_395);
xor U664 (N_664,In_93,N_576);
xor U665 (N_665,N_271,In_386);
and U666 (N_666,In_716,N_425);
nor U667 (N_667,N_563,N_358);
or U668 (N_668,N_259,N_302);
nor U669 (N_669,N_537,N_70);
and U670 (N_670,N_512,N_340);
or U671 (N_671,N_284,N_427);
nand U672 (N_672,N_227,N_401);
nand U673 (N_673,N_510,N_548);
nor U674 (N_674,N_584,N_547);
nor U675 (N_675,N_513,N_411);
xnor U676 (N_676,N_252,N_489);
nand U677 (N_677,N_409,N_437);
and U678 (N_678,N_295,In_277);
nor U679 (N_679,In_282,In_571);
nand U680 (N_680,In_369,N_591);
nor U681 (N_681,N_550,In_568);
or U682 (N_682,N_496,N_241);
xnor U683 (N_683,N_233,N_572);
nor U684 (N_684,In_500,N_485);
or U685 (N_685,N_226,N_150);
nand U686 (N_686,N_148,N_486);
nor U687 (N_687,N_519,In_417);
nand U688 (N_688,N_522,N_508);
nor U689 (N_689,N_69,N_215);
and U690 (N_690,In_882,N_473);
xnor U691 (N_691,N_592,N_443);
and U692 (N_692,N_76,N_306);
or U693 (N_693,In_445,In_481);
nand U694 (N_694,N_554,N_201);
nand U695 (N_695,N_435,N_392);
xnor U696 (N_696,N_516,N_490);
nor U697 (N_697,In_820,N_429);
or U698 (N_698,N_551,N_593);
and U699 (N_699,N_287,In_200);
xor U700 (N_700,N_246,N_415);
nand U701 (N_701,N_469,N_504);
or U702 (N_702,N_439,N_372);
nand U703 (N_703,N_459,N_569);
nand U704 (N_704,In_60,N_502);
nand U705 (N_705,N_465,N_37);
nor U706 (N_706,N_356,N_539);
xnor U707 (N_707,In_829,N_416);
or U708 (N_708,N_418,In_963);
xnor U709 (N_709,In_899,N_421);
and U710 (N_710,N_571,N_21);
and U711 (N_711,N_446,N_428);
xor U712 (N_712,N_488,N_454);
xnor U713 (N_713,N_453,N_369);
and U714 (N_714,N_463,N_475);
nand U715 (N_715,N_423,In_664);
nor U716 (N_716,N_581,In_361);
or U717 (N_717,N_125,In_421);
nand U718 (N_718,In_375,In_526);
nand U719 (N_719,N_466,N_562);
and U720 (N_720,N_442,N_558);
xnor U721 (N_721,N_161,In_556);
and U722 (N_722,N_567,N_100);
nand U723 (N_723,N_507,In_12);
xor U724 (N_724,N_402,N_546);
nand U725 (N_725,In_140,N_498);
and U726 (N_726,N_267,N_484);
xnor U727 (N_727,N_440,N_509);
nor U728 (N_728,N_352,N_535);
nor U729 (N_729,N_482,N_111);
or U730 (N_730,N_151,N_574);
and U731 (N_731,In_279,N_395);
nor U732 (N_732,In_183,N_217);
and U733 (N_733,In_618,N_472);
nor U734 (N_734,In_210,N_445);
nor U735 (N_735,N_585,N_520);
and U736 (N_736,In_466,N_598);
or U737 (N_737,N_526,In_53);
or U738 (N_738,N_413,N_540);
xnor U739 (N_739,In_742,In_337);
nor U740 (N_740,N_536,N_456);
xnor U741 (N_741,N_599,N_236);
nand U742 (N_742,N_455,N_579);
nand U743 (N_743,In_24,N_434);
or U744 (N_744,In_380,N_249);
nand U745 (N_745,N_414,In_819);
nor U746 (N_746,N_531,In_249);
xor U747 (N_747,N_521,In_220);
nand U748 (N_748,In_756,In_555);
nor U749 (N_749,N_119,In_471);
or U750 (N_750,In_917,N_590);
nor U751 (N_751,N_90,N_134);
or U752 (N_752,N_203,N_255);
xor U753 (N_753,In_217,N_419);
or U754 (N_754,N_494,N_450);
nor U755 (N_755,N_296,In_50);
or U756 (N_756,In_112,In_594);
xnor U757 (N_757,N_438,In_591);
and U758 (N_758,N_524,N_575);
nor U759 (N_759,N_582,N_594);
nor U760 (N_760,In_946,N_426);
xor U761 (N_761,N_478,N_432);
and U762 (N_762,N_560,In_908);
nand U763 (N_763,N_545,In_995);
nor U764 (N_764,N_573,N_514);
nand U765 (N_765,N_281,In_942);
nand U766 (N_766,N_433,N_499);
and U767 (N_767,N_559,N_424);
xnor U768 (N_768,N_387,N_307);
xnor U769 (N_769,N_43,In_846);
xnor U770 (N_770,In_791,In_63);
and U771 (N_771,In_433,N_477);
and U772 (N_772,N_420,N_370);
xnor U773 (N_773,In_559,In_509);
or U774 (N_774,N_109,N_588);
nor U775 (N_775,N_422,N_595);
nor U776 (N_776,N_544,N_187);
nor U777 (N_777,In_980,N_467);
and U778 (N_778,In_704,N_447);
nor U779 (N_779,N_470,N_138);
nor U780 (N_780,N_532,N_28);
xnor U781 (N_781,N_346,N_202);
nor U782 (N_782,N_408,In_767);
and U783 (N_783,In_119,N_376);
or U784 (N_784,N_479,N_436);
nand U785 (N_785,N_444,N_505);
nand U786 (N_786,N_384,N_495);
and U787 (N_787,N_515,N_460);
nor U788 (N_788,In_66,N_483);
xnor U789 (N_789,N_568,N_332);
or U790 (N_790,N_471,In_118);
xor U791 (N_791,In_242,In_378);
xor U792 (N_792,N_319,In_377);
nand U793 (N_793,In_920,N_523);
and U794 (N_794,In_576,In_207);
and U795 (N_795,N_89,N_441);
nand U796 (N_796,N_565,In_858);
nand U797 (N_797,N_385,N_386);
or U798 (N_798,N_268,N_491);
nand U799 (N_799,In_318,N_326);
nand U800 (N_800,N_667,N_759);
xor U801 (N_801,N_699,N_690);
nand U802 (N_802,N_752,N_682);
nor U803 (N_803,N_732,N_642);
or U804 (N_804,N_734,N_737);
nand U805 (N_805,N_607,N_624);
xor U806 (N_806,N_795,N_742);
xor U807 (N_807,N_719,N_611);
and U808 (N_808,N_632,N_685);
xnor U809 (N_809,N_687,N_747);
nand U810 (N_810,N_622,N_681);
or U811 (N_811,N_676,N_783);
nor U812 (N_812,N_645,N_730);
or U813 (N_813,N_680,N_653);
nor U814 (N_814,N_691,N_639);
nand U815 (N_815,N_620,N_609);
or U816 (N_816,N_600,N_689);
nand U817 (N_817,N_655,N_654);
nand U818 (N_818,N_688,N_651);
or U819 (N_819,N_779,N_672);
nor U820 (N_820,N_794,N_659);
or U821 (N_821,N_608,N_677);
or U822 (N_822,N_702,N_711);
and U823 (N_823,N_623,N_604);
xor U824 (N_824,N_644,N_735);
xnor U825 (N_825,N_754,N_733);
nor U826 (N_826,N_673,N_612);
and U827 (N_827,N_780,N_731);
and U828 (N_828,N_727,N_615);
or U829 (N_829,N_774,N_728);
or U830 (N_830,N_648,N_722);
and U831 (N_831,N_698,N_618);
nand U832 (N_832,N_764,N_661);
nand U833 (N_833,N_776,N_791);
nand U834 (N_834,N_606,N_790);
and U835 (N_835,N_649,N_652);
or U836 (N_836,N_736,N_744);
nand U837 (N_837,N_769,N_671);
xnor U838 (N_838,N_700,N_758);
or U839 (N_839,N_773,N_757);
xnor U840 (N_840,N_745,N_785);
nand U841 (N_841,N_762,N_713);
nand U842 (N_842,N_631,N_772);
xnor U843 (N_843,N_637,N_692);
or U844 (N_844,N_740,N_721);
and U845 (N_845,N_704,N_646);
nor U846 (N_846,N_751,N_799);
xnor U847 (N_847,N_670,N_696);
or U848 (N_848,N_705,N_760);
xnor U849 (N_849,N_787,N_628);
and U850 (N_850,N_766,N_750);
nand U851 (N_851,N_712,N_613);
nand U852 (N_852,N_647,N_775);
xor U853 (N_853,N_788,N_703);
nor U854 (N_854,N_683,N_657);
and U855 (N_855,N_718,N_796);
nand U856 (N_856,N_658,N_694);
xnor U857 (N_857,N_669,N_708);
and U858 (N_858,N_761,N_656);
xnor U859 (N_859,N_634,N_743);
or U860 (N_860,N_725,N_605);
xnor U861 (N_861,N_602,N_638);
or U862 (N_862,N_621,N_756);
nor U863 (N_863,N_697,N_729);
nor U864 (N_864,N_636,N_633);
nor U865 (N_865,N_695,N_701);
nand U866 (N_866,N_617,N_715);
or U867 (N_867,N_753,N_716);
xor U868 (N_868,N_640,N_650);
and U869 (N_869,N_706,N_627);
and U870 (N_870,N_663,N_614);
nand U871 (N_871,N_797,N_723);
nor U872 (N_872,N_748,N_643);
nor U873 (N_873,N_789,N_684);
nor U874 (N_874,N_675,N_610);
or U875 (N_875,N_767,N_726);
nor U876 (N_876,N_770,N_777);
xnor U877 (N_877,N_601,N_741);
xor U878 (N_878,N_665,N_792);
nor U879 (N_879,N_768,N_707);
nand U880 (N_880,N_660,N_784);
and U881 (N_881,N_771,N_720);
or U882 (N_882,N_755,N_619);
or U883 (N_883,N_782,N_635);
or U884 (N_884,N_668,N_765);
nand U885 (N_885,N_662,N_746);
or U886 (N_886,N_724,N_738);
and U887 (N_887,N_603,N_625);
nand U888 (N_888,N_666,N_793);
and U889 (N_889,N_714,N_630);
nor U890 (N_890,N_709,N_798);
nor U891 (N_891,N_674,N_781);
nand U892 (N_892,N_679,N_629);
or U893 (N_893,N_641,N_763);
and U894 (N_894,N_717,N_778);
or U895 (N_895,N_616,N_678);
and U896 (N_896,N_739,N_686);
nand U897 (N_897,N_710,N_693);
nor U898 (N_898,N_626,N_749);
and U899 (N_899,N_664,N_786);
nor U900 (N_900,N_690,N_798);
xor U901 (N_901,N_612,N_782);
nand U902 (N_902,N_614,N_626);
nand U903 (N_903,N_727,N_690);
nor U904 (N_904,N_652,N_685);
or U905 (N_905,N_600,N_652);
nor U906 (N_906,N_684,N_799);
xor U907 (N_907,N_693,N_794);
nand U908 (N_908,N_600,N_764);
and U909 (N_909,N_659,N_694);
nand U910 (N_910,N_611,N_665);
nand U911 (N_911,N_643,N_644);
and U912 (N_912,N_617,N_655);
xor U913 (N_913,N_631,N_734);
nor U914 (N_914,N_645,N_638);
nand U915 (N_915,N_691,N_643);
and U916 (N_916,N_609,N_683);
or U917 (N_917,N_608,N_770);
or U918 (N_918,N_785,N_684);
xor U919 (N_919,N_747,N_658);
nor U920 (N_920,N_743,N_649);
nand U921 (N_921,N_760,N_625);
xor U922 (N_922,N_655,N_684);
and U923 (N_923,N_762,N_668);
or U924 (N_924,N_674,N_656);
nor U925 (N_925,N_744,N_749);
nor U926 (N_926,N_637,N_760);
nor U927 (N_927,N_746,N_633);
or U928 (N_928,N_785,N_662);
and U929 (N_929,N_719,N_715);
or U930 (N_930,N_658,N_724);
nand U931 (N_931,N_757,N_646);
nor U932 (N_932,N_742,N_700);
and U933 (N_933,N_739,N_748);
nand U934 (N_934,N_647,N_731);
nor U935 (N_935,N_792,N_678);
nand U936 (N_936,N_768,N_735);
nand U937 (N_937,N_759,N_698);
xor U938 (N_938,N_765,N_679);
xor U939 (N_939,N_729,N_678);
or U940 (N_940,N_745,N_774);
nand U941 (N_941,N_713,N_601);
nand U942 (N_942,N_719,N_689);
nor U943 (N_943,N_675,N_708);
nand U944 (N_944,N_775,N_670);
xor U945 (N_945,N_758,N_732);
or U946 (N_946,N_771,N_712);
xor U947 (N_947,N_742,N_686);
nor U948 (N_948,N_634,N_701);
nand U949 (N_949,N_654,N_735);
nor U950 (N_950,N_688,N_696);
nor U951 (N_951,N_615,N_637);
nor U952 (N_952,N_745,N_644);
nand U953 (N_953,N_612,N_762);
and U954 (N_954,N_642,N_767);
nand U955 (N_955,N_604,N_641);
or U956 (N_956,N_711,N_643);
nand U957 (N_957,N_723,N_762);
nand U958 (N_958,N_799,N_757);
xor U959 (N_959,N_776,N_706);
xnor U960 (N_960,N_692,N_626);
or U961 (N_961,N_771,N_616);
nor U962 (N_962,N_689,N_740);
nor U963 (N_963,N_654,N_741);
nor U964 (N_964,N_796,N_685);
nand U965 (N_965,N_612,N_798);
nor U966 (N_966,N_669,N_688);
nand U967 (N_967,N_601,N_603);
nand U968 (N_968,N_709,N_767);
nand U969 (N_969,N_666,N_712);
nor U970 (N_970,N_797,N_718);
xnor U971 (N_971,N_659,N_660);
or U972 (N_972,N_776,N_678);
nor U973 (N_973,N_687,N_629);
or U974 (N_974,N_673,N_633);
nand U975 (N_975,N_760,N_648);
nor U976 (N_976,N_699,N_745);
or U977 (N_977,N_669,N_633);
or U978 (N_978,N_668,N_619);
nand U979 (N_979,N_757,N_706);
or U980 (N_980,N_697,N_726);
nor U981 (N_981,N_677,N_783);
nand U982 (N_982,N_722,N_610);
and U983 (N_983,N_733,N_753);
nand U984 (N_984,N_669,N_714);
or U985 (N_985,N_767,N_724);
nand U986 (N_986,N_742,N_628);
or U987 (N_987,N_655,N_630);
nor U988 (N_988,N_655,N_621);
nor U989 (N_989,N_624,N_791);
xor U990 (N_990,N_752,N_732);
nand U991 (N_991,N_659,N_739);
xnor U992 (N_992,N_654,N_798);
xnor U993 (N_993,N_687,N_681);
nand U994 (N_994,N_681,N_618);
and U995 (N_995,N_754,N_656);
nor U996 (N_996,N_750,N_625);
nand U997 (N_997,N_607,N_671);
xnor U998 (N_998,N_783,N_688);
xor U999 (N_999,N_659,N_775);
nand U1000 (N_1000,N_848,N_871);
xnor U1001 (N_1001,N_812,N_890);
and U1002 (N_1002,N_979,N_868);
or U1003 (N_1003,N_875,N_949);
or U1004 (N_1004,N_866,N_847);
and U1005 (N_1005,N_938,N_973);
or U1006 (N_1006,N_860,N_894);
or U1007 (N_1007,N_915,N_869);
nor U1008 (N_1008,N_907,N_991);
nor U1009 (N_1009,N_930,N_892);
and U1010 (N_1010,N_923,N_842);
xnor U1011 (N_1011,N_966,N_925);
nand U1012 (N_1012,N_820,N_950);
xor U1013 (N_1013,N_945,N_963);
or U1014 (N_1014,N_959,N_971);
and U1015 (N_1015,N_886,N_993);
nand U1016 (N_1016,N_840,N_948);
nand U1017 (N_1017,N_934,N_805);
or U1018 (N_1018,N_839,N_821);
nand U1019 (N_1019,N_882,N_906);
nand U1020 (N_1020,N_800,N_986);
or U1021 (N_1021,N_836,N_964);
or U1022 (N_1022,N_830,N_887);
nor U1023 (N_1023,N_832,N_919);
xnor U1024 (N_1024,N_898,N_804);
xnor U1025 (N_1025,N_845,N_953);
nor U1026 (N_1026,N_811,N_889);
nand U1027 (N_1027,N_989,N_951);
nand U1028 (N_1028,N_961,N_801);
nor U1029 (N_1029,N_834,N_806);
nand U1030 (N_1030,N_992,N_859);
nand U1031 (N_1031,N_940,N_904);
nor U1032 (N_1032,N_901,N_816);
nor U1033 (N_1033,N_879,N_981);
or U1034 (N_1034,N_935,N_962);
xnor U1035 (N_1035,N_908,N_813);
and U1036 (N_1036,N_877,N_880);
nor U1037 (N_1037,N_922,N_918);
or U1038 (N_1038,N_846,N_817);
xnor U1039 (N_1039,N_823,N_911);
xnor U1040 (N_1040,N_814,N_960);
xnor U1041 (N_1041,N_888,N_807);
nor U1042 (N_1042,N_861,N_972);
nor U1043 (N_1043,N_975,N_958);
nand U1044 (N_1044,N_917,N_863);
xnor U1045 (N_1045,N_990,N_921);
nand U1046 (N_1046,N_885,N_891);
xor U1047 (N_1047,N_984,N_858);
nand U1048 (N_1048,N_974,N_946);
xnor U1049 (N_1049,N_883,N_916);
nand U1050 (N_1050,N_838,N_835);
or U1051 (N_1051,N_831,N_987);
or U1052 (N_1052,N_954,N_980);
nor U1053 (N_1053,N_909,N_867);
and U1054 (N_1054,N_941,N_955);
xnor U1055 (N_1055,N_942,N_824);
and U1056 (N_1056,N_878,N_873);
nor U1057 (N_1057,N_932,N_996);
nand U1058 (N_1058,N_976,N_927);
and U1059 (N_1059,N_998,N_822);
nor U1060 (N_1060,N_982,N_897);
and U1061 (N_1061,N_870,N_827);
or U1062 (N_1062,N_825,N_896);
xor U1063 (N_1063,N_999,N_893);
xnor U1064 (N_1064,N_850,N_970);
or U1065 (N_1065,N_829,N_881);
nand U1066 (N_1066,N_988,N_928);
or U1067 (N_1067,N_844,N_905);
nand U1068 (N_1068,N_900,N_864);
and U1069 (N_1069,N_841,N_818);
xor U1070 (N_1070,N_874,N_968);
and U1071 (N_1071,N_914,N_956);
xnor U1072 (N_1072,N_913,N_849);
nand U1073 (N_1073,N_983,N_920);
or U1074 (N_1074,N_809,N_912);
xor U1075 (N_1075,N_903,N_994);
nor U1076 (N_1076,N_895,N_828);
nor U1077 (N_1077,N_947,N_884);
and U1078 (N_1078,N_967,N_802);
and U1079 (N_1079,N_910,N_865);
nor U1080 (N_1080,N_985,N_937);
nand U1081 (N_1081,N_978,N_997);
xnor U1082 (N_1082,N_929,N_926);
and U1083 (N_1083,N_952,N_851);
nand U1084 (N_1084,N_969,N_862);
and U1085 (N_1085,N_876,N_815);
nor U1086 (N_1086,N_810,N_977);
or U1087 (N_1087,N_995,N_944);
xnor U1088 (N_1088,N_853,N_852);
xor U1089 (N_1089,N_965,N_819);
nand U1090 (N_1090,N_826,N_854);
xnor U1091 (N_1091,N_957,N_837);
nand U1092 (N_1092,N_857,N_803);
xnor U1093 (N_1093,N_833,N_808);
xnor U1094 (N_1094,N_872,N_855);
nand U1095 (N_1095,N_939,N_899);
or U1096 (N_1096,N_933,N_936);
or U1097 (N_1097,N_943,N_902);
nand U1098 (N_1098,N_856,N_843);
nor U1099 (N_1099,N_924,N_931);
xor U1100 (N_1100,N_846,N_890);
or U1101 (N_1101,N_980,N_904);
or U1102 (N_1102,N_990,N_876);
and U1103 (N_1103,N_908,N_824);
and U1104 (N_1104,N_977,N_827);
and U1105 (N_1105,N_893,N_860);
nor U1106 (N_1106,N_841,N_970);
and U1107 (N_1107,N_965,N_810);
and U1108 (N_1108,N_837,N_849);
nand U1109 (N_1109,N_845,N_904);
nor U1110 (N_1110,N_849,N_990);
or U1111 (N_1111,N_863,N_816);
or U1112 (N_1112,N_898,N_973);
or U1113 (N_1113,N_868,N_930);
or U1114 (N_1114,N_852,N_921);
nand U1115 (N_1115,N_958,N_923);
xnor U1116 (N_1116,N_960,N_817);
and U1117 (N_1117,N_942,N_905);
nor U1118 (N_1118,N_852,N_982);
nand U1119 (N_1119,N_945,N_914);
and U1120 (N_1120,N_899,N_817);
and U1121 (N_1121,N_815,N_881);
and U1122 (N_1122,N_840,N_998);
nor U1123 (N_1123,N_869,N_989);
xnor U1124 (N_1124,N_984,N_891);
and U1125 (N_1125,N_951,N_801);
nand U1126 (N_1126,N_871,N_854);
xor U1127 (N_1127,N_835,N_879);
and U1128 (N_1128,N_900,N_899);
nor U1129 (N_1129,N_893,N_971);
xor U1130 (N_1130,N_845,N_982);
nor U1131 (N_1131,N_967,N_853);
and U1132 (N_1132,N_956,N_864);
nand U1133 (N_1133,N_956,N_814);
nand U1134 (N_1134,N_829,N_805);
or U1135 (N_1135,N_847,N_867);
xor U1136 (N_1136,N_807,N_837);
xnor U1137 (N_1137,N_853,N_842);
nand U1138 (N_1138,N_950,N_964);
nor U1139 (N_1139,N_936,N_908);
or U1140 (N_1140,N_805,N_819);
nand U1141 (N_1141,N_894,N_900);
nand U1142 (N_1142,N_876,N_989);
and U1143 (N_1143,N_908,N_909);
and U1144 (N_1144,N_865,N_881);
and U1145 (N_1145,N_896,N_996);
and U1146 (N_1146,N_916,N_800);
nand U1147 (N_1147,N_955,N_881);
xnor U1148 (N_1148,N_889,N_981);
and U1149 (N_1149,N_953,N_992);
xnor U1150 (N_1150,N_800,N_835);
xor U1151 (N_1151,N_840,N_945);
xnor U1152 (N_1152,N_826,N_895);
nor U1153 (N_1153,N_987,N_884);
or U1154 (N_1154,N_875,N_819);
xor U1155 (N_1155,N_919,N_932);
nand U1156 (N_1156,N_937,N_860);
nand U1157 (N_1157,N_843,N_984);
xnor U1158 (N_1158,N_848,N_976);
or U1159 (N_1159,N_948,N_853);
xor U1160 (N_1160,N_914,N_991);
and U1161 (N_1161,N_992,N_843);
xnor U1162 (N_1162,N_914,N_977);
nand U1163 (N_1163,N_821,N_948);
or U1164 (N_1164,N_865,N_944);
and U1165 (N_1165,N_915,N_980);
or U1166 (N_1166,N_989,N_808);
nand U1167 (N_1167,N_997,N_960);
or U1168 (N_1168,N_937,N_822);
or U1169 (N_1169,N_939,N_812);
nor U1170 (N_1170,N_993,N_898);
nand U1171 (N_1171,N_897,N_896);
nand U1172 (N_1172,N_851,N_890);
nor U1173 (N_1173,N_877,N_869);
nand U1174 (N_1174,N_966,N_934);
nor U1175 (N_1175,N_828,N_968);
nor U1176 (N_1176,N_934,N_844);
nor U1177 (N_1177,N_927,N_894);
nand U1178 (N_1178,N_863,N_861);
nand U1179 (N_1179,N_832,N_957);
and U1180 (N_1180,N_875,N_835);
xnor U1181 (N_1181,N_804,N_906);
nand U1182 (N_1182,N_878,N_883);
or U1183 (N_1183,N_887,N_910);
nor U1184 (N_1184,N_870,N_869);
nor U1185 (N_1185,N_821,N_858);
nor U1186 (N_1186,N_876,N_866);
xnor U1187 (N_1187,N_870,N_929);
nor U1188 (N_1188,N_978,N_873);
and U1189 (N_1189,N_974,N_933);
xor U1190 (N_1190,N_876,N_914);
nand U1191 (N_1191,N_908,N_930);
xor U1192 (N_1192,N_811,N_802);
or U1193 (N_1193,N_862,N_878);
and U1194 (N_1194,N_908,N_884);
xor U1195 (N_1195,N_939,N_859);
nand U1196 (N_1196,N_822,N_934);
and U1197 (N_1197,N_994,N_987);
or U1198 (N_1198,N_952,N_919);
and U1199 (N_1199,N_926,N_823);
or U1200 (N_1200,N_1185,N_1105);
nand U1201 (N_1201,N_1012,N_1188);
and U1202 (N_1202,N_1135,N_1171);
nor U1203 (N_1203,N_1156,N_1179);
xnor U1204 (N_1204,N_1022,N_1057);
or U1205 (N_1205,N_1143,N_1180);
nand U1206 (N_1206,N_1147,N_1033);
and U1207 (N_1207,N_1168,N_1037);
nand U1208 (N_1208,N_1183,N_1198);
nor U1209 (N_1209,N_1187,N_1065);
or U1210 (N_1210,N_1106,N_1128);
and U1211 (N_1211,N_1148,N_1052);
nand U1212 (N_1212,N_1056,N_1005);
nor U1213 (N_1213,N_1170,N_1023);
nand U1214 (N_1214,N_1112,N_1092);
nor U1215 (N_1215,N_1080,N_1102);
nor U1216 (N_1216,N_1169,N_1027);
nor U1217 (N_1217,N_1016,N_1142);
and U1218 (N_1218,N_1197,N_1104);
and U1219 (N_1219,N_1082,N_1044);
or U1220 (N_1220,N_1091,N_1100);
nor U1221 (N_1221,N_1086,N_1085);
nand U1222 (N_1222,N_1046,N_1140);
or U1223 (N_1223,N_1077,N_1083);
or U1224 (N_1224,N_1003,N_1103);
nand U1225 (N_1225,N_1184,N_1165);
nand U1226 (N_1226,N_1132,N_1018);
xnor U1227 (N_1227,N_1117,N_1172);
or U1228 (N_1228,N_1029,N_1114);
nor U1229 (N_1229,N_1006,N_1045);
and U1230 (N_1230,N_1152,N_1062);
nand U1231 (N_1231,N_1043,N_1011);
and U1232 (N_1232,N_1134,N_1025);
or U1233 (N_1233,N_1119,N_1155);
or U1234 (N_1234,N_1164,N_1141);
nor U1235 (N_1235,N_1162,N_1113);
xor U1236 (N_1236,N_1054,N_1078);
nand U1237 (N_1237,N_1042,N_1049);
or U1238 (N_1238,N_1111,N_1059);
xnor U1239 (N_1239,N_1160,N_1190);
nand U1240 (N_1240,N_1001,N_1067);
xnor U1241 (N_1241,N_1074,N_1019);
and U1242 (N_1242,N_1060,N_1017);
or U1243 (N_1243,N_1136,N_1163);
xnor U1244 (N_1244,N_1153,N_1173);
nand U1245 (N_1245,N_1020,N_1000);
nand U1246 (N_1246,N_1158,N_1079);
nand U1247 (N_1247,N_1076,N_1154);
nand U1248 (N_1248,N_1058,N_1069);
xor U1249 (N_1249,N_1161,N_1186);
nor U1250 (N_1250,N_1068,N_1196);
nor U1251 (N_1251,N_1014,N_1167);
xnor U1252 (N_1252,N_1159,N_1093);
nor U1253 (N_1253,N_1035,N_1130);
nand U1254 (N_1254,N_1150,N_1108);
nor U1255 (N_1255,N_1071,N_1176);
or U1256 (N_1256,N_1090,N_1010);
and U1257 (N_1257,N_1129,N_1036);
nand U1258 (N_1258,N_1070,N_1116);
nor U1259 (N_1259,N_1121,N_1028);
or U1260 (N_1260,N_1110,N_1099);
and U1261 (N_1261,N_1144,N_1026);
nand U1262 (N_1262,N_1084,N_1107);
xnor U1263 (N_1263,N_1032,N_1021);
xnor U1264 (N_1264,N_1055,N_1008);
and U1265 (N_1265,N_1118,N_1131);
or U1266 (N_1266,N_1125,N_1175);
or U1267 (N_1267,N_1038,N_1115);
xor U1268 (N_1268,N_1098,N_1149);
nand U1269 (N_1269,N_1031,N_1195);
xor U1270 (N_1270,N_1181,N_1138);
and U1271 (N_1271,N_1166,N_1007);
xor U1272 (N_1272,N_1101,N_1199);
xor U1273 (N_1273,N_1015,N_1039);
and U1274 (N_1274,N_1096,N_1194);
nor U1275 (N_1275,N_1157,N_1002);
xnor U1276 (N_1276,N_1073,N_1094);
nand U1277 (N_1277,N_1064,N_1061);
nor U1278 (N_1278,N_1030,N_1081);
xnor U1279 (N_1279,N_1095,N_1109);
xnor U1280 (N_1280,N_1097,N_1034);
and U1281 (N_1281,N_1177,N_1072);
and U1282 (N_1282,N_1146,N_1137);
nand U1283 (N_1283,N_1024,N_1122);
or U1284 (N_1284,N_1040,N_1009);
or U1285 (N_1285,N_1050,N_1051);
or U1286 (N_1286,N_1087,N_1123);
nand U1287 (N_1287,N_1191,N_1124);
nor U1288 (N_1288,N_1120,N_1053);
nand U1289 (N_1289,N_1013,N_1126);
and U1290 (N_1290,N_1047,N_1189);
xnor U1291 (N_1291,N_1139,N_1066);
xnor U1292 (N_1292,N_1063,N_1075);
or U1293 (N_1293,N_1178,N_1088);
or U1294 (N_1294,N_1182,N_1127);
nand U1295 (N_1295,N_1151,N_1089);
nand U1296 (N_1296,N_1041,N_1048);
nand U1297 (N_1297,N_1193,N_1004);
and U1298 (N_1298,N_1145,N_1174);
xor U1299 (N_1299,N_1192,N_1133);
nor U1300 (N_1300,N_1170,N_1112);
and U1301 (N_1301,N_1037,N_1015);
and U1302 (N_1302,N_1037,N_1022);
nand U1303 (N_1303,N_1064,N_1175);
or U1304 (N_1304,N_1059,N_1032);
xnor U1305 (N_1305,N_1025,N_1167);
nor U1306 (N_1306,N_1172,N_1011);
nand U1307 (N_1307,N_1035,N_1101);
nand U1308 (N_1308,N_1131,N_1150);
nor U1309 (N_1309,N_1139,N_1076);
nand U1310 (N_1310,N_1169,N_1057);
or U1311 (N_1311,N_1041,N_1178);
or U1312 (N_1312,N_1089,N_1088);
nor U1313 (N_1313,N_1137,N_1033);
nand U1314 (N_1314,N_1187,N_1034);
nand U1315 (N_1315,N_1133,N_1083);
xor U1316 (N_1316,N_1135,N_1143);
nand U1317 (N_1317,N_1144,N_1117);
nor U1318 (N_1318,N_1198,N_1002);
or U1319 (N_1319,N_1050,N_1142);
xnor U1320 (N_1320,N_1101,N_1095);
and U1321 (N_1321,N_1057,N_1081);
and U1322 (N_1322,N_1123,N_1153);
xor U1323 (N_1323,N_1191,N_1059);
and U1324 (N_1324,N_1074,N_1006);
nor U1325 (N_1325,N_1130,N_1143);
xnor U1326 (N_1326,N_1185,N_1101);
xor U1327 (N_1327,N_1124,N_1056);
nor U1328 (N_1328,N_1133,N_1015);
and U1329 (N_1329,N_1047,N_1096);
and U1330 (N_1330,N_1082,N_1019);
nand U1331 (N_1331,N_1127,N_1060);
xnor U1332 (N_1332,N_1150,N_1140);
nor U1333 (N_1333,N_1068,N_1093);
xnor U1334 (N_1334,N_1081,N_1183);
xor U1335 (N_1335,N_1109,N_1132);
xnor U1336 (N_1336,N_1010,N_1074);
or U1337 (N_1337,N_1137,N_1091);
nand U1338 (N_1338,N_1173,N_1060);
or U1339 (N_1339,N_1092,N_1083);
nor U1340 (N_1340,N_1061,N_1091);
nor U1341 (N_1341,N_1120,N_1044);
or U1342 (N_1342,N_1131,N_1061);
nand U1343 (N_1343,N_1039,N_1147);
nand U1344 (N_1344,N_1130,N_1165);
nand U1345 (N_1345,N_1071,N_1081);
nor U1346 (N_1346,N_1008,N_1111);
nor U1347 (N_1347,N_1168,N_1106);
nand U1348 (N_1348,N_1032,N_1040);
nand U1349 (N_1349,N_1115,N_1078);
xnor U1350 (N_1350,N_1024,N_1043);
or U1351 (N_1351,N_1130,N_1175);
nor U1352 (N_1352,N_1078,N_1069);
nor U1353 (N_1353,N_1161,N_1061);
or U1354 (N_1354,N_1151,N_1116);
nor U1355 (N_1355,N_1138,N_1008);
xor U1356 (N_1356,N_1116,N_1139);
xor U1357 (N_1357,N_1048,N_1091);
xor U1358 (N_1358,N_1025,N_1147);
nand U1359 (N_1359,N_1173,N_1013);
xnor U1360 (N_1360,N_1155,N_1172);
or U1361 (N_1361,N_1162,N_1045);
xnor U1362 (N_1362,N_1108,N_1013);
nor U1363 (N_1363,N_1129,N_1034);
xor U1364 (N_1364,N_1053,N_1124);
or U1365 (N_1365,N_1170,N_1072);
xor U1366 (N_1366,N_1099,N_1057);
xnor U1367 (N_1367,N_1192,N_1039);
or U1368 (N_1368,N_1090,N_1026);
nand U1369 (N_1369,N_1131,N_1099);
or U1370 (N_1370,N_1097,N_1069);
and U1371 (N_1371,N_1147,N_1040);
nand U1372 (N_1372,N_1124,N_1059);
nand U1373 (N_1373,N_1161,N_1163);
xor U1374 (N_1374,N_1119,N_1017);
and U1375 (N_1375,N_1066,N_1026);
nand U1376 (N_1376,N_1068,N_1048);
and U1377 (N_1377,N_1192,N_1009);
or U1378 (N_1378,N_1027,N_1003);
nor U1379 (N_1379,N_1164,N_1182);
nand U1380 (N_1380,N_1021,N_1181);
nor U1381 (N_1381,N_1046,N_1101);
or U1382 (N_1382,N_1116,N_1077);
nand U1383 (N_1383,N_1116,N_1008);
and U1384 (N_1384,N_1047,N_1140);
or U1385 (N_1385,N_1119,N_1064);
and U1386 (N_1386,N_1074,N_1082);
nand U1387 (N_1387,N_1076,N_1156);
or U1388 (N_1388,N_1187,N_1143);
nor U1389 (N_1389,N_1027,N_1161);
xor U1390 (N_1390,N_1148,N_1031);
xor U1391 (N_1391,N_1122,N_1110);
and U1392 (N_1392,N_1079,N_1176);
and U1393 (N_1393,N_1147,N_1044);
or U1394 (N_1394,N_1128,N_1080);
nor U1395 (N_1395,N_1052,N_1087);
nor U1396 (N_1396,N_1022,N_1105);
nand U1397 (N_1397,N_1025,N_1132);
and U1398 (N_1398,N_1181,N_1103);
or U1399 (N_1399,N_1104,N_1102);
or U1400 (N_1400,N_1366,N_1303);
or U1401 (N_1401,N_1347,N_1221);
nand U1402 (N_1402,N_1282,N_1307);
nand U1403 (N_1403,N_1293,N_1243);
and U1404 (N_1404,N_1200,N_1277);
and U1405 (N_1405,N_1321,N_1320);
nand U1406 (N_1406,N_1270,N_1222);
xnor U1407 (N_1407,N_1244,N_1223);
nor U1408 (N_1408,N_1241,N_1345);
nand U1409 (N_1409,N_1383,N_1352);
or U1410 (N_1410,N_1279,N_1396);
nor U1411 (N_1411,N_1262,N_1297);
and U1412 (N_1412,N_1357,N_1249);
xor U1413 (N_1413,N_1387,N_1225);
and U1414 (N_1414,N_1254,N_1230);
nor U1415 (N_1415,N_1388,N_1274);
nor U1416 (N_1416,N_1360,N_1259);
or U1417 (N_1417,N_1286,N_1275);
nor U1418 (N_1418,N_1367,N_1340);
and U1419 (N_1419,N_1364,N_1215);
and U1420 (N_1420,N_1304,N_1228);
and U1421 (N_1421,N_1398,N_1229);
or U1422 (N_1422,N_1386,N_1336);
xnor U1423 (N_1423,N_1319,N_1240);
nand U1424 (N_1424,N_1231,N_1355);
nand U1425 (N_1425,N_1373,N_1338);
or U1426 (N_1426,N_1219,N_1264);
xnor U1427 (N_1427,N_1369,N_1202);
nor U1428 (N_1428,N_1385,N_1330);
xnor U1429 (N_1429,N_1327,N_1354);
xnor U1430 (N_1430,N_1343,N_1232);
nor U1431 (N_1431,N_1310,N_1276);
xor U1432 (N_1432,N_1337,N_1204);
xnor U1433 (N_1433,N_1271,N_1258);
and U1434 (N_1434,N_1392,N_1314);
nor U1435 (N_1435,N_1300,N_1236);
nand U1436 (N_1436,N_1322,N_1361);
nand U1437 (N_1437,N_1266,N_1227);
nor U1438 (N_1438,N_1280,N_1389);
nand U1439 (N_1439,N_1213,N_1305);
and U1440 (N_1440,N_1341,N_1207);
or U1441 (N_1441,N_1217,N_1390);
nand U1442 (N_1442,N_1237,N_1356);
xor U1443 (N_1443,N_1375,N_1203);
and U1444 (N_1444,N_1209,N_1292);
nand U1445 (N_1445,N_1278,N_1212);
nand U1446 (N_1446,N_1260,N_1285);
nand U1447 (N_1447,N_1291,N_1395);
xnor U1448 (N_1448,N_1290,N_1201);
nand U1449 (N_1449,N_1296,N_1288);
nand U1450 (N_1450,N_1211,N_1308);
nor U1451 (N_1451,N_1206,N_1214);
or U1452 (N_1452,N_1245,N_1272);
nand U1453 (N_1453,N_1318,N_1346);
nor U1454 (N_1454,N_1252,N_1391);
or U1455 (N_1455,N_1208,N_1316);
nand U1456 (N_1456,N_1309,N_1250);
and U1457 (N_1457,N_1265,N_1363);
or U1458 (N_1458,N_1205,N_1251);
xnor U1459 (N_1459,N_1339,N_1324);
nor U1460 (N_1460,N_1370,N_1323);
and U1461 (N_1461,N_1247,N_1353);
or U1462 (N_1462,N_1218,N_1326);
nand U1463 (N_1463,N_1382,N_1284);
xnor U1464 (N_1464,N_1331,N_1380);
xnor U1465 (N_1465,N_1216,N_1374);
nand U1466 (N_1466,N_1381,N_1253);
or U1467 (N_1467,N_1220,N_1301);
xor U1468 (N_1468,N_1394,N_1224);
and U1469 (N_1469,N_1298,N_1273);
xnor U1470 (N_1470,N_1295,N_1238);
nand U1471 (N_1471,N_1332,N_1317);
xnor U1472 (N_1472,N_1378,N_1350);
nor U1473 (N_1473,N_1239,N_1306);
nand U1474 (N_1474,N_1234,N_1334);
or U1475 (N_1475,N_1344,N_1248);
nand U1476 (N_1476,N_1311,N_1267);
nand U1477 (N_1477,N_1315,N_1377);
and U1478 (N_1478,N_1368,N_1342);
or U1479 (N_1479,N_1372,N_1287);
or U1480 (N_1480,N_1358,N_1329);
nor U1481 (N_1481,N_1283,N_1242);
or U1482 (N_1482,N_1365,N_1269);
or U1483 (N_1483,N_1299,N_1235);
xor U1484 (N_1484,N_1371,N_1379);
nor U1485 (N_1485,N_1263,N_1397);
xor U1486 (N_1486,N_1281,N_1257);
and U1487 (N_1487,N_1335,N_1325);
and U1488 (N_1488,N_1294,N_1268);
xnor U1489 (N_1489,N_1384,N_1328);
and U1490 (N_1490,N_1349,N_1362);
xor U1491 (N_1491,N_1313,N_1393);
xor U1492 (N_1492,N_1376,N_1359);
or U1493 (N_1493,N_1289,N_1351);
nand U1494 (N_1494,N_1399,N_1348);
xnor U1495 (N_1495,N_1261,N_1226);
or U1496 (N_1496,N_1302,N_1333);
nor U1497 (N_1497,N_1233,N_1256);
or U1498 (N_1498,N_1210,N_1312);
or U1499 (N_1499,N_1255,N_1246);
and U1500 (N_1500,N_1254,N_1277);
xnor U1501 (N_1501,N_1314,N_1264);
xor U1502 (N_1502,N_1325,N_1255);
xnor U1503 (N_1503,N_1258,N_1353);
xnor U1504 (N_1504,N_1341,N_1386);
xor U1505 (N_1505,N_1221,N_1220);
xnor U1506 (N_1506,N_1341,N_1354);
and U1507 (N_1507,N_1337,N_1269);
nor U1508 (N_1508,N_1384,N_1299);
nor U1509 (N_1509,N_1251,N_1338);
or U1510 (N_1510,N_1297,N_1311);
nand U1511 (N_1511,N_1212,N_1207);
xor U1512 (N_1512,N_1225,N_1311);
nand U1513 (N_1513,N_1252,N_1271);
or U1514 (N_1514,N_1271,N_1243);
or U1515 (N_1515,N_1202,N_1277);
nor U1516 (N_1516,N_1397,N_1288);
xnor U1517 (N_1517,N_1209,N_1205);
or U1518 (N_1518,N_1298,N_1377);
nand U1519 (N_1519,N_1377,N_1262);
and U1520 (N_1520,N_1271,N_1313);
or U1521 (N_1521,N_1386,N_1353);
xor U1522 (N_1522,N_1318,N_1259);
and U1523 (N_1523,N_1260,N_1247);
xor U1524 (N_1524,N_1242,N_1207);
xnor U1525 (N_1525,N_1260,N_1336);
nor U1526 (N_1526,N_1343,N_1339);
xnor U1527 (N_1527,N_1263,N_1224);
nand U1528 (N_1528,N_1361,N_1320);
nand U1529 (N_1529,N_1336,N_1318);
xnor U1530 (N_1530,N_1274,N_1202);
nor U1531 (N_1531,N_1258,N_1317);
nand U1532 (N_1532,N_1327,N_1363);
or U1533 (N_1533,N_1303,N_1339);
or U1534 (N_1534,N_1365,N_1332);
nor U1535 (N_1535,N_1326,N_1393);
and U1536 (N_1536,N_1382,N_1328);
or U1537 (N_1537,N_1262,N_1268);
or U1538 (N_1538,N_1315,N_1207);
nand U1539 (N_1539,N_1316,N_1320);
or U1540 (N_1540,N_1208,N_1342);
nand U1541 (N_1541,N_1237,N_1288);
nor U1542 (N_1542,N_1229,N_1385);
nand U1543 (N_1543,N_1202,N_1209);
xor U1544 (N_1544,N_1259,N_1261);
xnor U1545 (N_1545,N_1311,N_1212);
xor U1546 (N_1546,N_1303,N_1285);
and U1547 (N_1547,N_1222,N_1313);
xor U1548 (N_1548,N_1301,N_1256);
xnor U1549 (N_1549,N_1341,N_1398);
xnor U1550 (N_1550,N_1294,N_1266);
or U1551 (N_1551,N_1383,N_1355);
xor U1552 (N_1552,N_1309,N_1389);
and U1553 (N_1553,N_1346,N_1347);
xnor U1554 (N_1554,N_1245,N_1302);
nor U1555 (N_1555,N_1373,N_1309);
or U1556 (N_1556,N_1249,N_1393);
or U1557 (N_1557,N_1388,N_1370);
and U1558 (N_1558,N_1260,N_1328);
xnor U1559 (N_1559,N_1228,N_1330);
xor U1560 (N_1560,N_1255,N_1365);
xnor U1561 (N_1561,N_1244,N_1318);
nor U1562 (N_1562,N_1317,N_1218);
nand U1563 (N_1563,N_1307,N_1365);
nand U1564 (N_1564,N_1325,N_1252);
nor U1565 (N_1565,N_1213,N_1331);
and U1566 (N_1566,N_1255,N_1386);
and U1567 (N_1567,N_1345,N_1250);
or U1568 (N_1568,N_1306,N_1317);
xor U1569 (N_1569,N_1252,N_1256);
nand U1570 (N_1570,N_1328,N_1232);
and U1571 (N_1571,N_1287,N_1331);
and U1572 (N_1572,N_1205,N_1287);
or U1573 (N_1573,N_1366,N_1273);
or U1574 (N_1574,N_1370,N_1244);
nor U1575 (N_1575,N_1282,N_1236);
or U1576 (N_1576,N_1309,N_1200);
xor U1577 (N_1577,N_1389,N_1223);
or U1578 (N_1578,N_1355,N_1319);
xor U1579 (N_1579,N_1366,N_1327);
xor U1580 (N_1580,N_1212,N_1251);
nand U1581 (N_1581,N_1281,N_1348);
and U1582 (N_1582,N_1372,N_1344);
xnor U1583 (N_1583,N_1248,N_1289);
nand U1584 (N_1584,N_1318,N_1345);
xor U1585 (N_1585,N_1273,N_1325);
nand U1586 (N_1586,N_1304,N_1314);
and U1587 (N_1587,N_1211,N_1324);
xnor U1588 (N_1588,N_1384,N_1215);
or U1589 (N_1589,N_1203,N_1211);
xnor U1590 (N_1590,N_1296,N_1276);
nand U1591 (N_1591,N_1313,N_1378);
nand U1592 (N_1592,N_1222,N_1360);
nand U1593 (N_1593,N_1212,N_1303);
nand U1594 (N_1594,N_1275,N_1255);
nor U1595 (N_1595,N_1306,N_1226);
and U1596 (N_1596,N_1320,N_1257);
xor U1597 (N_1597,N_1374,N_1294);
and U1598 (N_1598,N_1288,N_1316);
xnor U1599 (N_1599,N_1235,N_1338);
and U1600 (N_1600,N_1564,N_1555);
or U1601 (N_1601,N_1401,N_1513);
and U1602 (N_1602,N_1484,N_1455);
and U1603 (N_1603,N_1549,N_1477);
nand U1604 (N_1604,N_1505,N_1404);
or U1605 (N_1605,N_1506,N_1454);
or U1606 (N_1606,N_1571,N_1527);
or U1607 (N_1607,N_1490,N_1433);
or U1608 (N_1608,N_1457,N_1532);
and U1609 (N_1609,N_1557,N_1551);
nand U1610 (N_1610,N_1517,N_1451);
nor U1611 (N_1611,N_1581,N_1406);
xnor U1612 (N_1612,N_1473,N_1594);
xnor U1613 (N_1613,N_1511,N_1592);
or U1614 (N_1614,N_1499,N_1576);
and U1615 (N_1615,N_1418,N_1461);
and U1616 (N_1616,N_1588,N_1493);
and U1617 (N_1617,N_1480,N_1482);
and U1618 (N_1618,N_1568,N_1421);
or U1619 (N_1619,N_1538,N_1509);
nor U1620 (N_1620,N_1546,N_1475);
xor U1621 (N_1621,N_1420,N_1472);
nor U1622 (N_1622,N_1528,N_1501);
or U1623 (N_1623,N_1437,N_1492);
and U1624 (N_1624,N_1452,N_1453);
and U1625 (N_1625,N_1467,N_1589);
and U1626 (N_1626,N_1500,N_1458);
nand U1627 (N_1627,N_1531,N_1518);
xnor U1628 (N_1628,N_1550,N_1577);
nor U1629 (N_1629,N_1495,N_1402);
nand U1630 (N_1630,N_1598,N_1560);
or U1631 (N_1631,N_1412,N_1439);
and U1632 (N_1632,N_1587,N_1488);
nand U1633 (N_1633,N_1425,N_1521);
nand U1634 (N_1634,N_1416,N_1471);
xor U1635 (N_1635,N_1438,N_1429);
xor U1636 (N_1636,N_1556,N_1444);
and U1637 (N_1637,N_1442,N_1573);
nor U1638 (N_1638,N_1515,N_1540);
nand U1639 (N_1639,N_1534,N_1574);
nand U1640 (N_1640,N_1408,N_1547);
xor U1641 (N_1641,N_1428,N_1462);
or U1642 (N_1642,N_1435,N_1507);
and U1643 (N_1643,N_1519,N_1504);
xor U1644 (N_1644,N_1431,N_1449);
nand U1645 (N_1645,N_1562,N_1566);
nand U1646 (N_1646,N_1464,N_1586);
or U1647 (N_1647,N_1569,N_1409);
and U1648 (N_1648,N_1403,N_1479);
nor U1649 (N_1649,N_1489,N_1502);
or U1650 (N_1650,N_1459,N_1456);
nand U1651 (N_1651,N_1539,N_1561);
nand U1652 (N_1652,N_1413,N_1470);
and U1653 (N_1653,N_1432,N_1526);
or U1654 (N_1654,N_1595,N_1423);
nand U1655 (N_1655,N_1494,N_1415);
nor U1656 (N_1656,N_1448,N_1434);
nor U1657 (N_1657,N_1422,N_1414);
nor U1658 (N_1658,N_1537,N_1520);
nand U1659 (N_1659,N_1536,N_1580);
or U1660 (N_1660,N_1447,N_1597);
xnor U1661 (N_1661,N_1446,N_1426);
nor U1662 (N_1662,N_1544,N_1584);
and U1663 (N_1663,N_1545,N_1559);
xnor U1664 (N_1664,N_1525,N_1483);
and U1665 (N_1665,N_1558,N_1567);
nor U1666 (N_1666,N_1563,N_1565);
and U1667 (N_1667,N_1548,N_1485);
and U1668 (N_1668,N_1440,N_1543);
or U1669 (N_1669,N_1582,N_1436);
nor U1670 (N_1670,N_1474,N_1405);
nand U1671 (N_1671,N_1512,N_1400);
xnor U1672 (N_1672,N_1496,N_1486);
nand U1673 (N_1673,N_1596,N_1530);
nor U1674 (N_1674,N_1572,N_1599);
xnor U1675 (N_1675,N_1578,N_1460);
and U1676 (N_1676,N_1575,N_1523);
nor U1677 (N_1677,N_1508,N_1553);
nor U1678 (N_1678,N_1554,N_1427);
nor U1679 (N_1679,N_1510,N_1443);
and U1680 (N_1680,N_1417,N_1516);
xor U1681 (N_1681,N_1579,N_1570);
nand U1682 (N_1682,N_1590,N_1491);
nand U1683 (N_1683,N_1465,N_1541);
nor U1684 (N_1684,N_1542,N_1552);
or U1685 (N_1685,N_1478,N_1468);
nor U1686 (N_1686,N_1411,N_1481);
and U1687 (N_1687,N_1524,N_1498);
xnor U1688 (N_1688,N_1476,N_1533);
or U1689 (N_1689,N_1535,N_1529);
nor U1690 (N_1690,N_1469,N_1583);
nor U1691 (N_1691,N_1591,N_1487);
nor U1692 (N_1692,N_1503,N_1497);
and U1693 (N_1693,N_1410,N_1466);
and U1694 (N_1694,N_1430,N_1463);
nand U1695 (N_1695,N_1424,N_1407);
nor U1696 (N_1696,N_1419,N_1445);
nand U1697 (N_1697,N_1585,N_1593);
xnor U1698 (N_1698,N_1522,N_1441);
nand U1699 (N_1699,N_1514,N_1450);
or U1700 (N_1700,N_1597,N_1536);
nand U1701 (N_1701,N_1409,N_1596);
xor U1702 (N_1702,N_1564,N_1562);
xnor U1703 (N_1703,N_1449,N_1480);
and U1704 (N_1704,N_1536,N_1469);
and U1705 (N_1705,N_1412,N_1512);
or U1706 (N_1706,N_1434,N_1422);
nand U1707 (N_1707,N_1488,N_1544);
or U1708 (N_1708,N_1401,N_1410);
xnor U1709 (N_1709,N_1501,N_1431);
nand U1710 (N_1710,N_1580,N_1529);
or U1711 (N_1711,N_1517,N_1481);
nand U1712 (N_1712,N_1592,N_1471);
nand U1713 (N_1713,N_1586,N_1500);
and U1714 (N_1714,N_1448,N_1552);
nor U1715 (N_1715,N_1407,N_1413);
nor U1716 (N_1716,N_1591,N_1511);
xnor U1717 (N_1717,N_1476,N_1546);
nor U1718 (N_1718,N_1563,N_1417);
nand U1719 (N_1719,N_1406,N_1477);
and U1720 (N_1720,N_1517,N_1582);
or U1721 (N_1721,N_1466,N_1475);
or U1722 (N_1722,N_1555,N_1489);
or U1723 (N_1723,N_1496,N_1420);
nand U1724 (N_1724,N_1503,N_1421);
and U1725 (N_1725,N_1444,N_1511);
xnor U1726 (N_1726,N_1553,N_1558);
nand U1727 (N_1727,N_1429,N_1480);
xor U1728 (N_1728,N_1535,N_1590);
or U1729 (N_1729,N_1491,N_1505);
xor U1730 (N_1730,N_1545,N_1599);
and U1731 (N_1731,N_1542,N_1596);
xnor U1732 (N_1732,N_1466,N_1596);
nand U1733 (N_1733,N_1531,N_1433);
nor U1734 (N_1734,N_1410,N_1583);
or U1735 (N_1735,N_1436,N_1411);
xor U1736 (N_1736,N_1595,N_1513);
nand U1737 (N_1737,N_1485,N_1512);
or U1738 (N_1738,N_1456,N_1495);
xor U1739 (N_1739,N_1472,N_1509);
xor U1740 (N_1740,N_1547,N_1574);
and U1741 (N_1741,N_1468,N_1534);
nor U1742 (N_1742,N_1580,N_1522);
or U1743 (N_1743,N_1508,N_1571);
or U1744 (N_1744,N_1423,N_1493);
nand U1745 (N_1745,N_1597,N_1571);
and U1746 (N_1746,N_1541,N_1430);
and U1747 (N_1747,N_1529,N_1403);
and U1748 (N_1748,N_1578,N_1441);
xnor U1749 (N_1749,N_1504,N_1522);
nor U1750 (N_1750,N_1458,N_1466);
or U1751 (N_1751,N_1574,N_1552);
and U1752 (N_1752,N_1492,N_1462);
xor U1753 (N_1753,N_1415,N_1477);
nor U1754 (N_1754,N_1476,N_1451);
nor U1755 (N_1755,N_1491,N_1565);
nor U1756 (N_1756,N_1504,N_1568);
nor U1757 (N_1757,N_1545,N_1525);
nand U1758 (N_1758,N_1584,N_1515);
nor U1759 (N_1759,N_1419,N_1537);
nand U1760 (N_1760,N_1592,N_1479);
and U1761 (N_1761,N_1542,N_1404);
xnor U1762 (N_1762,N_1575,N_1425);
nand U1763 (N_1763,N_1538,N_1569);
nand U1764 (N_1764,N_1577,N_1515);
and U1765 (N_1765,N_1409,N_1559);
and U1766 (N_1766,N_1427,N_1489);
and U1767 (N_1767,N_1464,N_1441);
nand U1768 (N_1768,N_1436,N_1469);
nor U1769 (N_1769,N_1504,N_1582);
or U1770 (N_1770,N_1510,N_1546);
nand U1771 (N_1771,N_1405,N_1559);
xnor U1772 (N_1772,N_1468,N_1583);
nand U1773 (N_1773,N_1512,N_1589);
or U1774 (N_1774,N_1594,N_1401);
nand U1775 (N_1775,N_1592,N_1578);
and U1776 (N_1776,N_1540,N_1422);
or U1777 (N_1777,N_1588,N_1474);
nor U1778 (N_1778,N_1591,N_1507);
xor U1779 (N_1779,N_1500,N_1406);
nand U1780 (N_1780,N_1429,N_1485);
nand U1781 (N_1781,N_1473,N_1460);
and U1782 (N_1782,N_1424,N_1483);
xor U1783 (N_1783,N_1589,N_1483);
and U1784 (N_1784,N_1591,N_1561);
and U1785 (N_1785,N_1461,N_1490);
xor U1786 (N_1786,N_1540,N_1579);
xnor U1787 (N_1787,N_1576,N_1509);
nor U1788 (N_1788,N_1584,N_1590);
nor U1789 (N_1789,N_1520,N_1585);
nor U1790 (N_1790,N_1596,N_1451);
nand U1791 (N_1791,N_1548,N_1470);
nor U1792 (N_1792,N_1593,N_1532);
or U1793 (N_1793,N_1445,N_1435);
and U1794 (N_1794,N_1596,N_1565);
nor U1795 (N_1795,N_1400,N_1473);
and U1796 (N_1796,N_1458,N_1503);
xnor U1797 (N_1797,N_1467,N_1537);
or U1798 (N_1798,N_1486,N_1466);
nand U1799 (N_1799,N_1502,N_1454);
or U1800 (N_1800,N_1650,N_1659);
nand U1801 (N_1801,N_1743,N_1782);
xnor U1802 (N_1802,N_1605,N_1786);
nor U1803 (N_1803,N_1711,N_1600);
and U1804 (N_1804,N_1716,N_1710);
or U1805 (N_1805,N_1696,N_1636);
nor U1806 (N_1806,N_1703,N_1758);
xor U1807 (N_1807,N_1756,N_1668);
nand U1808 (N_1808,N_1647,N_1734);
and U1809 (N_1809,N_1686,N_1671);
nand U1810 (N_1810,N_1601,N_1742);
and U1811 (N_1811,N_1737,N_1763);
xnor U1812 (N_1812,N_1673,N_1749);
nor U1813 (N_1813,N_1704,N_1660);
nor U1814 (N_1814,N_1765,N_1715);
or U1815 (N_1815,N_1757,N_1642);
nand U1816 (N_1816,N_1791,N_1717);
and U1817 (N_1817,N_1613,N_1744);
nor U1818 (N_1818,N_1700,N_1677);
nand U1819 (N_1819,N_1627,N_1759);
xor U1820 (N_1820,N_1665,N_1718);
nor U1821 (N_1821,N_1616,N_1643);
or U1822 (N_1822,N_1621,N_1609);
nor U1823 (N_1823,N_1730,N_1761);
nand U1824 (N_1824,N_1784,N_1767);
or U1825 (N_1825,N_1741,N_1688);
and U1826 (N_1826,N_1787,N_1721);
nand U1827 (N_1827,N_1745,N_1752);
and U1828 (N_1828,N_1632,N_1633);
or U1829 (N_1829,N_1682,N_1794);
nor U1830 (N_1830,N_1753,N_1653);
or U1831 (N_1831,N_1661,N_1729);
or U1832 (N_1832,N_1738,N_1691);
nand U1833 (N_1833,N_1768,N_1707);
nor U1834 (N_1834,N_1622,N_1610);
xnor U1835 (N_1835,N_1766,N_1614);
and U1836 (N_1836,N_1722,N_1676);
nor U1837 (N_1837,N_1771,N_1635);
nand U1838 (N_1838,N_1736,N_1777);
or U1839 (N_1839,N_1626,N_1618);
nand U1840 (N_1840,N_1663,N_1732);
nand U1841 (N_1841,N_1774,N_1685);
or U1842 (N_1842,N_1769,N_1712);
and U1843 (N_1843,N_1681,N_1735);
nor U1844 (N_1844,N_1683,N_1638);
or U1845 (N_1845,N_1629,N_1720);
or U1846 (N_1846,N_1666,N_1713);
nand U1847 (N_1847,N_1687,N_1706);
or U1848 (N_1848,N_1640,N_1695);
nand U1849 (N_1849,N_1624,N_1657);
xor U1850 (N_1850,N_1679,N_1669);
nor U1851 (N_1851,N_1760,N_1764);
or U1852 (N_1852,N_1772,N_1630);
nor U1853 (N_1853,N_1689,N_1724);
nor U1854 (N_1854,N_1776,N_1655);
nor U1855 (N_1855,N_1654,N_1723);
or U1856 (N_1856,N_1746,N_1781);
and U1857 (N_1857,N_1625,N_1641);
nand U1858 (N_1858,N_1697,N_1797);
nand U1859 (N_1859,N_1719,N_1708);
nor U1860 (N_1860,N_1615,N_1733);
or U1861 (N_1861,N_1634,N_1796);
or U1862 (N_1862,N_1652,N_1658);
or U1863 (N_1863,N_1762,N_1603);
or U1864 (N_1864,N_1608,N_1790);
and U1865 (N_1865,N_1645,N_1656);
or U1866 (N_1866,N_1779,N_1693);
xor U1867 (N_1867,N_1611,N_1792);
nand U1868 (N_1868,N_1714,N_1728);
nor U1869 (N_1869,N_1694,N_1788);
nor U1870 (N_1870,N_1754,N_1602);
nand U1871 (N_1871,N_1662,N_1678);
nor U1872 (N_1872,N_1675,N_1799);
nor U1873 (N_1873,N_1725,N_1664);
or U1874 (N_1874,N_1604,N_1698);
xnor U1875 (N_1875,N_1667,N_1619);
xor U1876 (N_1876,N_1637,N_1623);
or U1877 (N_1877,N_1607,N_1680);
or U1878 (N_1878,N_1684,N_1701);
nor U1879 (N_1879,N_1690,N_1778);
nor U1880 (N_1880,N_1702,N_1649);
xor U1881 (N_1881,N_1748,N_1651);
xnor U1882 (N_1882,N_1709,N_1648);
nor U1883 (N_1883,N_1795,N_1631);
and U1884 (N_1884,N_1793,N_1726);
nand U1885 (N_1885,N_1750,N_1670);
or U1886 (N_1886,N_1798,N_1699);
or U1887 (N_1887,N_1674,N_1639);
and U1888 (N_1888,N_1740,N_1780);
and U1889 (N_1889,N_1705,N_1739);
or U1890 (N_1890,N_1751,N_1755);
nand U1891 (N_1891,N_1773,N_1785);
or U1892 (N_1892,N_1617,N_1644);
and U1893 (N_1893,N_1775,N_1770);
and U1894 (N_1894,N_1646,N_1727);
nor U1895 (N_1895,N_1789,N_1620);
or U1896 (N_1896,N_1783,N_1731);
nor U1897 (N_1897,N_1672,N_1628);
and U1898 (N_1898,N_1606,N_1692);
or U1899 (N_1899,N_1747,N_1612);
nand U1900 (N_1900,N_1779,N_1794);
and U1901 (N_1901,N_1606,N_1695);
nor U1902 (N_1902,N_1622,N_1615);
nor U1903 (N_1903,N_1672,N_1731);
or U1904 (N_1904,N_1649,N_1634);
and U1905 (N_1905,N_1784,N_1696);
nor U1906 (N_1906,N_1749,N_1651);
nor U1907 (N_1907,N_1727,N_1656);
nor U1908 (N_1908,N_1679,N_1775);
or U1909 (N_1909,N_1781,N_1608);
or U1910 (N_1910,N_1691,N_1781);
and U1911 (N_1911,N_1733,N_1772);
nand U1912 (N_1912,N_1610,N_1715);
nor U1913 (N_1913,N_1678,N_1735);
nand U1914 (N_1914,N_1775,N_1761);
or U1915 (N_1915,N_1699,N_1787);
and U1916 (N_1916,N_1722,N_1769);
and U1917 (N_1917,N_1684,N_1768);
or U1918 (N_1918,N_1740,N_1654);
or U1919 (N_1919,N_1772,N_1631);
xor U1920 (N_1920,N_1745,N_1688);
nand U1921 (N_1921,N_1680,N_1726);
or U1922 (N_1922,N_1714,N_1671);
and U1923 (N_1923,N_1706,N_1669);
nor U1924 (N_1924,N_1768,N_1751);
or U1925 (N_1925,N_1689,N_1780);
or U1926 (N_1926,N_1610,N_1696);
nor U1927 (N_1927,N_1659,N_1767);
or U1928 (N_1928,N_1785,N_1721);
and U1929 (N_1929,N_1725,N_1710);
nand U1930 (N_1930,N_1669,N_1742);
nand U1931 (N_1931,N_1779,N_1703);
or U1932 (N_1932,N_1747,N_1791);
xor U1933 (N_1933,N_1623,N_1767);
or U1934 (N_1934,N_1753,N_1717);
or U1935 (N_1935,N_1686,N_1718);
xnor U1936 (N_1936,N_1771,N_1610);
xor U1937 (N_1937,N_1615,N_1772);
or U1938 (N_1938,N_1646,N_1767);
and U1939 (N_1939,N_1758,N_1741);
or U1940 (N_1940,N_1775,N_1712);
nor U1941 (N_1941,N_1641,N_1617);
or U1942 (N_1942,N_1628,N_1662);
nand U1943 (N_1943,N_1665,N_1714);
and U1944 (N_1944,N_1790,N_1764);
or U1945 (N_1945,N_1735,N_1601);
and U1946 (N_1946,N_1686,N_1682);
and U1947 (N_1947,N_1703,N_1687);
nor U1948 (N_1948,N_1643,N_1647);
nand U1949 (N_1949,N_1670,N_1613);
or U1950 (N_1950,N_1626,N_1762);
nand U1951 (N_1951,N_1634,N_1799);
nand U1952 (N_1952,N_1666,N_1688);
nand U1953 (N_1953,N_1788,N_1782);
and U1954 (N_1954,N_1705,N_1660);
or U1955 (N_1955,N_1672,N_1629);
nor U1956 (N_1956,N_1709,N_1690);
xnor U1957 (N_1957,N_1714,N_1716);
nor U1958 (N_1958,N_1721,N_1603);
xnor U1959 (N_1959,N_1653,N_1663);
nor U1960 (N_1960,N_1618,N_1739);
nand U1961 (N_1961,N_1779,N_1619);
nand U1962 (N_1962,N_1665,N_1634);
and U1963 (N_1963,N_1727,N_1623);
or U1964 (N_1964,N_1781,N_1792);
or U1965 (N_1965,N_1600,N_1605);
or U1966 (N_1966,N_1649,N_1693);
nor U1967 (N_1967,N_1676,N_1609);
or U1968 (N_1968,N_1698,N_1748);
and U1969 (N_1969,N_1787,N_1740);
nand U1970 (N_1970,N_1689,N_1669);
nor U1971 (N_1971,N_1693,N_1799);
and U1972 (N_1972,N_1642,N_1743);
xor U1973 (N_1973,N_1607,N_1769);
nand U1974 (N_1974,N_1793,N_1606);
and U1975 (N_1975,N_1682,N_1764);
xnor U1976 (N_1976,N_1720,N_1786);
and U1977 (N_1977,N_1691,N_1668);
or U1978 (N_1978,N_1797,N_1674);
nand U1979 (N_1979,N_1642,N_1680);
nor U1980 (N_1980,N_1609,N_1683);
and U1981 (N_1981,N_1778,N_1652);
or U1982 (N_1982,N_1790,N_1667);
xor U1983 (N_1983,N_1683,N_1604);
and U1984 (N_1984,N_1713,N_1659);
xor U1985 (N_1985,N_1724,N_1699);
nand U1986 (N_1986,N_1716,N_1641);
nand U1987 (N_1987,N_1744,N_1600);
or U1988 (N_1988,N_1702,N_1758);
nor U1989 (N_1989,N_1666,N_1789);
nand U1990 (N_1990,N_1704,N_1762);
nor U1991 (N_1991,N_1697,N_1617);
xor U1992 (N_1992,N_1772,N_1774);
nor U1993 (N_1993,N_1648,N_1606);
xor U1994 (N_1994,N_1605,N_1725);
xnor U1995 (N_1995,N_1704,N_1763);
and U1996 (N_1996,N_1612,N_1752);
nand U1997 (N_1997,N_1648,N_1793);
xnor U1998 (N_1998,N_1677,N_1646);
nand U1999 (N_1999,N_1682,N_1601);
and U2000 (N_2000,N_1861,N_1902);
nand U2001 (N_2001,N_1917,N_1903);
nor U2002 (N_2002,N_1932,N_1893);
or U2003 (N_2003,N_1975,N_1988);
nand U2004 (N_2004,N_1976,N_1986);
xor U2005 (N_2005,N_1947,N_1918);
nand U2006 (N_2006,N_1831,N_1995);
nand U2007 (N_2007,N_1821,N_1996);
nor U2008 (N_2008,N_1997,N_1973);
xnor U2009 (N_2009,N_1824,N_1966);
nor U2010 (N_2010,N_1803,N_1895);
xor U2011 (N_2011,N_1854,N_1907);
and U2012 (N_2012,N_1872,N_1925);
and U2013 (N_2013,N_1941,N_1874);
nor U2014 (N_2014,N_1804,N_1914);
or U2015 (N_2015,N_1823,N_1980);
nor U2016 (N_2016,N_1828,N_1969);
xor U2017 (N_2017,N_1919,N_1837);
nor U2018 (N_2018,N_1911,N_1838);
and U2019 (N_2019,N_1886,N_1816);
nor U2020 (N_2020,N_1952,N_1807);
xor U2021 (N_2021,N_1956,N_1910);
xor U2022 (N_2022,N_1999,N_1845);
nor U2023 (N_2023,N_1990,N_1938);
and U2024 (N_2024,N_1965,N_1891);
or U2025 (N_2025,N_1846,N_1819);
nand U2026 (N_2026,N_1987,N_1915);
nand U2027 (N_2027,N_1979,N_1818);
or U2028 (N_2028,N_1815,N_1964);
and U2029 (N_2029,N_1960,N_1805);
and U2030 (N_2030,N_1834,N_1924);
nand U2031 (N_2031,N_1898,N_1928);
and U2032 (N_2032,N_1870,N_1880);
and U2033 (N_2033,N_1878,N_1998);
or U2034 (N_2034,N_1901,N_1867);
and U2035 (N_2035,N_1904,N_1820);
xnor U2036 (N_2036,N_1847,N_1953);
or U2037 (N_2037,N_1936,N_1868);
xor U2038 (N_2038,N_1905,N_1929);
or U2039 (N_2039,N_1926,N_1993);
or U2040 (N_2040,N_1897,N_1800);
or U2041 (N_2041,N_1842,N_1857);
and U2042 (N_2042,N_1841,N_1963);
or U2043 (N_2043,N_1916,N_1927);
nor U2044 (N_2044,N_1801,N_1931);
and U2045 (N_2045,N_1866,N_1982);
nand U2046 (N_2046,N_1912,N_1812);
nor U2047 (N_2047,N_1942,N_1968);
nand U2048 (N_2048,N_1961,N_1978);
nand U2049 (N_2049,N_1962,N_1977);
nand U2050 (N_2050,N_1954,N_1922);
or U2051 (N_2051,N_1827,N_1970);
or U2052 (N_2052,N_1882,N_1894);
nand U2053 (N_2053,N_1948,N_1985);
nand U2054 (N_2054,N_1808,N_1810);
or U2055 (N_2055,N_1989,N_1983);
or U2056 (N_2056,N_1863,N_1865);
or U2057 (N_2057,N_1851,N_1935);
nor U2058 (N_2058,N_1848,N_1833);
or U2059 (N_2059,N_1850,N_1814);
xnor U2060 (N_2060,N_1809,N_1825);
or U2061 (N_2061,N_1829,N_1817);
nand U2062 (N_2062,N_1991,N_1885);
and U2063 (N_2063,N_1887,N_1855);
and U2064 (N_2064,N_1869,N_1873);
xor U2065 (N_2065,N_1945,N_1971);
or U2066 (N_2066,N_1860,N_1877);
nand U2067 (N_2067,N_1862,N_1864);
and U2068 (N_2068,N_1913,N_1967);
nor U2069 (N_2069,N_1889,N_1802);
or U2070 (N_2070,N_1974,N_1994);
and U2071 (N_2071,N_1881,N_1888);
nor U2072 (N_2072,N_1940,N_1899);
nand U2073 (N_2073,N_1875,N_1852);
and U2074 (N_2074,N_1871,N_1835);
or U2075 (N_2075,N_1951,N_1959);
or U2076 (N_2076,N_1984,N_1896);
nand U2077 (N_2077,N_1950,N_1900);
nor U2078 (N_2078,N_1843,N_1981);
nor U2079 (N_2079,N_1853,N_1858);
or U2080 (N_2080,N_1958,N_1906);
or U2081 (N_2081,N_1811,N_1884);
nor U2082 (N_2082,N_1859,N_1806);
nand U2083 (N_2083,N_1836,N_1933);
or U2084 (N_2084,N_1946,N_1923);
xnor U2085 (N_2085,N_1844,N_1957);
nand U2086 (N_2086,N_1949,N_1937);
or U2087 (N_2087,N_1934,N_1908);
or U2088 (N_2088,N_1892,N_1849);
xnor U2089 (N_2089,N_1822,N_1876);
or U2090 (N_2090,N_1909,N_1832);
nand U2091 (N_2091,N_1920,N_1890);
nor U2092 (N_2092,N_1944,N_1856);
nand U2093 (N_2093,N_1839,N_1992);
xor U2094 (N_2094,N_1930,N_1879);
nor U2095 (N_2095,N_1939,N_1972);
xnor U2096 (N_2096,N_1883,N_1813);
or U2097 (N_2097,N_1826,N_1921);
and U2098 (N_2098,N_1840,N_1830);
or U2099 (N_2099,N_1943,N_1955);
and U2100 (N_2100,N_1894,N_1965);
nand U2101 (N_2101,N_1918,N_1894);
xnor U2102 (N_2102,N_1882,N_1949);
and U2103 (N_2103,N_1989,N_1869);
nor U2104 (N_2104,N_1962,N_1920);
nand U2105 (N_2105,N_1969,N_1807);
xnor U2106 (N_2106,N_1961,N_1854);
nor U2107 (N_2107,N_1824,N_1909);
nor U2108 (N_2108,N_1947,N_1973);
xor U2109 (N_2109,N_1839,N_1901);
nor U2110 (N_2110,N_1845,N_1913);
and U2111 (N_2111,N_1942,N_1995);
nor U2112 (N_2112,N_1890,N_1810);
xnor U2113 (N_2113,N_1830,N_1960);
and U2114 (N_2114,N_1843,N_1848);
nand U2115 (N_2115,N_1933,N_1838);
or U2116 (N_2116,N_1918,N_1815);
and U2117 (N_2117,N_1904,N_1921);
nand U2118 (N_2118,N_1841,N_1978);
nor U2119 (N_2119,N_1834,N_1892);
nor U2120 (N_2120,N_1970,N_1972);
or U2121 (N_2121,N_1930,N_1815);
and U2122 (N_2122,N_1909,N_1950);
nand U2123 (N_2123,N_1960,N_1853);
nor U2124 (N_2124,N_1975,N_1813);
or U2125 (N_2125,N_1933,N_1837);
nand U2126 (N_2126,N_1846,N_1974);
or U2127 (N_2127,N_1902,N_1880);
or U2128 (N_2128,N_1920,N_1995);
and U2129 (N_2129,N_1956,N_1986);
or U2130 (N_2130,N_1877,N_1976);
xor U2131 (N_2131,N_1914,N_1831);
xnor U2132 (N_2132,N_1828,N_1940);
nor U2133 (N_2133,N_1922,N_1956);
xor U2134 (N_2134,N_1846,N_1892);
or U2135 (N_2135,N_1992,N_1844);
nor U2136 (N_2136,N_1941,N_1875);
xnor U2137 (N_2137,N_1950,N_1837);
nand U2138 (N_2138,N_1836,N_1887);
or U2139 (N_2139,N_1924,N_1930);
xor U2140 (N_2140,N_1800,N_1944);
nand U2141 (N_2141,N_1846,N_1903);
nand U2142 (N_2142,N_1953,N_1933);
and U2143 (N_2143,N_1975,N_1905);
and U2144 (N_2144,N_1948,N_1953);
nand U2145 (N_2145,N_1858,N_1922);
nand U2146 (N_2146,N_1879,N_1964);
nor U2147 (N_2147,N_1881,N_1821);
and U2148 (N_2148,N_1936,N_1900);
or U2149 (N_2149,N_1938,N_1826);
xnor U2150 (N_2150,N_1832,N_1923);
or U2151 (N_2151,N_1966,N_1906);
nor U2152 (N_2152,N_1862,N_1815);
or U2153 (N_2153,N_1890,N_1908);
nor U2154 (N_2154,N_1881,N_1896);
xor U2155 (N_2155,N_1883,N_1902);
and U2156 (N_2156,N_1991,N_1869);
or U2157 (N_2157,N_1856,N_1812);
nand U2158 (N_2158,N_1877,N_1959);
nor U2159 (N_2159,N_1953,N_1977);
nor U2160 (N_2160,N_1988,N_1923);
nand U2161 (N_2161,N_1866,N_1977);
or U2162 (N_2162,N_1822,N_1819);
nor U2163 (N_2163,N_1850,N_1965);
nand U2164 (N_2164,N_1916,N_1907);
xnor U2165 (N_2165,N_1962,N_1876);
nand U2166 (N_2166,N_1819,N_1947);
and U2167 (N_2167,N_1958,N_1909);
xor U2168 (N_2168,N_1827,N_1854);
and U2169 (N_2169,N_1852,N_1964);
and U2170 (N_2170,N_1836,N_1869);
xor U2171 (N_2171,N_1837,N_1833);
or U2172 (N_2172,N_1801,N_1873);
nand U2173 (N_2173,N_1996,N_1941);
xnor U2174 (N_2174,N_1858,N_1859);
nor U2175 (N_2175,N_1845,N_1994);
nand U2176 (N_2176,N_1959,N_1965);
or U2177 (N_2177,N_1836,N_1958);
xnor U2178 (N_2178,N_1860,N_1921);
xor U2179 (N_2179,N_1921,N_1932);
or U2180 (N_2180,N_1853,N_1865);
and U2181 (N_2181,N_1887,N_1992);
and U2182 (N_2182,N_1917,N_1969);
nor U2183 (N_2183,N_1821,N_1835);
xor U2184 (N_2184,N_1818,N_1835);
and U2185 (N_2185,N_1994,N_1929);
or U2186 (N_2186,N_1925,N_1873);
nand U2187 (N_2187,N_1829,N_1839);
nor U2188 (N_2188,N_1816,N_1826);
nand U2189 (N_2189,N_1988,N_1835);
and U2190 (N_2190,N_1868,N_1941);
or U2191 (N_2191,N_1899,N_1991);
xnor U2192 (N_2192,N_1812,N_1837);
xor U2193 (N_2193,N_1840,N_1855);
nor U2194 (N_2194,N_1976,N_1971);
and U2195 (N_2195,N_1864,N_1815);
or U2196 (N_2196,N_1854,N_1930);
nand U2197 (N_2197,N_1927,N_1923);
and U2198 (N_2198,N_1820,N_1884);
or U2199 (N_2199,N_1858,N_1925);
or U2200 (N_2200,N_2072,N_2156);
and U2201 (N_2201,N_2158,N_2135);
xnor U2202 (N_2202,N_2108,N_2065);
or U2203 (N_2203,N_2151,N_2020);
and U2204 (N_2204,N_2141,N_2129);
nand U2205 (N_2205,N_2057,N_2149);
xnor U2206 (N_2206,N_2138,N_2159);
nor U2207 (N_2207,N_2031,N_2030);
nand U2208 (N_2208,N_2021,N_2060);
nor U2209 (N_2209,N_2167,N_2093);
nand U2210 (N_2210,N_2062,N_2170);
xnor U2211 (N_2211,N_2115,N_2015);
nand U2212 (N_2212,N_2175,N_2082);
nand U2213 (N_2213,N_2024,N_2081);
and U2214 (N_2214,N_2016,N_2096);
and U2215 (N_2215,N_2127,N_2023);
nand U2216 (N_2216,N_2098,N_2056);
nor U2217 (N_2217,N_2122,N_2107);
or U2218 (N_2218,N_2095,N_2187);
xor U2219 (N_2219,N_2152,N_2042);
nand U2220 (N_2220,N_2181,N_2007);
nand U2221 (N_2221,N_2100,N_2010);
nand U2222 (N_2222,N_2079,N_2184);
nand U2223 (N_2223,N_2124,N_2077);
nand U2224 (N_2224,N_2088,N_2097);
nand U2225 (N_2225,N_2011,N_2087);
xnor U2226 (N_2226,N_2155,N_2191);
or U2227 (N_2227,N_2084,N_2103);
nor U2228 (N_2228,N_2171,N_2070);
xor U2229 (N_2229,N_2085,N_2118);
and U2230 (N_2230,N_2195,N_2133);
xor U2231 (N_2231,N_2044,N_2026);
or U2232 (N_2232,N_2075,N_2001);
or U2233 (N_2233,N_2199,N_2025);
or U2234 (N_2234,N_2153,N_2005);
xnor U2235 (N_2235,N_2182,N_2193);
nor U2236 (N_2236,N_2148,N_2033);
and U2237 (N_2237,N_2116,N_2035);
and U2238 (N_2238,N_2132,N_2045);
xnor U2239 (N_2239,N_2080,N_2014);
or U2240 (N_2240,N_2022,N_2120);
and U2241 (N_2241,N_2053,N_2058);
xor U2242 (N_2242,N_2198,N_2050);
nand U2243 (N_2243,N_2076,N_2163);
xor U2244 (N_2244,N_2018,N_2136);
nor U2245 (N_2245,N_2092,N_2183);
xor U2246 (N_2246,N_2131,N_2164);
nand U2247 (N_2247,N_2119,N_2172);
xor U2248 (N_2248,N_2089,N_2126);
or U2249 (N_2249,N_2109,N_2117);
and U2250 (N_2250,N_2146,N_2143);
nand U2251 (N_2251,N_2157,N_2196);
nand U2252 (N_2252,N_2192,N_2180);
nand U2253 (N_2253,N_2165,N_2166);
or U2254 (N_2254,N_2003,N_2168);
nand U2255 (N_2255,N_2017,N_2130);
xor U2256 (N_2256,N_2176,N_2197);
nor U2257 (N_2257,N_2036,N_2169);
nand U2258 (N_2258,N_2094,N_2038);
nand U2259 (N_2259,N_2002,N_2055);
or U2260 (N_2260,N_2178,N_2110);
nand U2261 (N_2261,N_2039,N_2012);
nand U2262 (N_2262,N_2008,N_2123);
and U2263 (N_2263,N_2029,N_2069);
nor U2264 (N_2264,N_2105,N_2140);
xnor U2265 (N_2265,N_2034,N_2071);
or U2266 (N_2266,N_2154,N_2162);
or U2267 (N_2267,N_2186,N_2037);
nand U2268 (N_2268,N_2090,N_2043);
nand U2269 (N_2269,N_2161,N_2142);
nand U2270 (N_2270,N_2004,N_2099);
nand U2271 (N_2271,N_2027,N_2013);
and U2272 (N_2272,N_2188,N_2179);
nand U2273 (N_2273,N_2106,N_2000);
and U2274 (N_2274,N_2063,N_2137);
xor U2275 (N_2275,N_2047,N_2125);
and U2276 (N_2276,N_2112,N_2113);
nor U2277 (N_2277,N_2121,N_2101);
xor U2278 (N_2278,N_2066,N_2068);
nand U2279 (N_2279,N_2194,N_2041);
or U2280 (N_2280,N_2078,N_2173);
or U2281 (N_2281,N_2073,N_2114);
nor U2282 (N_2282,N_2019,N_2185);
xor U2283 (N_2283,N_2177,N_2040);
or U2284 (N_2284,N_2052,N_2061);
nand U2285 (N_2285,N_2128,N_2150);
nor U2286 (N_2286,N_2086,N_2147);
and U2287 (N_2287,N_2111,N_2174);
nand U2288 (N_2288,N_2009,N_2102);
nor U2289 (N_2289,N_2059,N_2028);
or U2290 (N_2290,N_2074,N_2054);
and U2291 (N_2291,N_2083,N_2046);
nand U2292 (N_2292,N_2032,N_2104);
xor U2293 (N_2293,N_2160,N_2049);
and U2294 (N_2294,N_2189,N_2144);
or U2295 (N_2295,N_2145,N_2064);
nor U2296 (N_2296,N_2048,N_2190);
nand U2297 (N_2297,N_2067,N_2091);
or U2298 (N_2298,N_2139,N_2134);
nor U2299 (N_2299,N_2051,N_2006);
nand U2300 (N_2300,N_2155,N_2132);
nor U2301 (N_2301,N_2073,N_2063);
nor U2302 (N_2302,N_2125,N_2024);
xnor U2303 (N_2303,N_2157,N_2006);
xor U2304 (N_2304,N_2081,N_2073);
nand U2305 (N_2305,N_2184,N_2188);
and U2306 (N_2306,N_2188,N_2031);
nand U2307 (N_2307,N_2133,N_2120);
nand U2308 (N_2308,N_2043,N_2028);
nand U2309 (N_2309,N_2003,N_2114);
nor U2310 (N_2310,N_2164,N_2001);
nand U2311 (N_2311,N_2090,N_2027);
nand U2312 (N_2312,N_2189,N_2021);
and U2313 (N_2313,N_2136,N_2155);
xor U2314 (N_2314,N_2152,N_2122);
nor U2315 (N_2315,N_2160,N_2129);
nand U2316 (N_2316,N_2024,N_2195);
xor U2317 (N_2317,N_2034,N_2043);
nand U2318 (N_2318,N_2061,N_2080);
nor U2319 (N_2319,N_2193,N_2155);
xor U2320 (N_2320,N_2014,N_2198);
nand U2321 (N_2321,N_2030,N_2056);
nor U2322 (N_2322,N_2101,N_2134);
xor U2323 (N_2323,N_2073,N_2083);
or U2324 (N_2324,N_2176,N_2052);
or U2325 (N_2325,N_2154,N_2132);
and U2326 (N_2326,N_2049,N_2180);
or U2327 (N_2327,N_2158,N_2082);
xor U2328 (N_2328,N_2116,N_2155);
nand U2329 (N_2329,N_2046,N_2068);
xnor U2330 (N_2330,N_2060,N_2179);
or U2331 (N_2331,N_2095,N_2175);
and U2332 (N_2332,N_2154,N_2124);
and U2333 (N_2333,N_2109,N_2199);
or U2334 (N_2334,N_2159,N_2133);
nor U2335 (N_2335,N_2162,N_2199);
nand U2336 (N_2336,N_2071,N_2143);
nor U2337 (N_2337,N_2171,N_2010);
or U2338 (N_2338,N_2066,N_2152);
nand U2339 (N_2339,N_2010,N_2057);
xor U2340 (N_2340,N_2138,N_2095);
xnor U2341 (N_2341,N_2111,N_2142);
or U2342 (N_2342,N_2113,N_2177);
xor U2343 (N_2343,N_2115,N_2094);
nand U2344 (N_2344,N_2199,N_2185);
and U2345 (N_2345,N_2076,N_2089);
nor U2346 (N_2346,N_2194,N_2184);
nand U2347 (N_2347,N_2166,N_2102);
xor U2348 (N_2348,N_2023,N_2007);
or U2349 (N_2349,N_2094,N_2015);
xor U2350 (N_2350,N_2092,N_2041);
xnor U2351 (N_2351,N_2056,N_2145);
nand U2352 (N_2352,N_2137,N_2148);
or U2353 (N_2353,N_2003,N_2078);
nor U2354 (N_2354,N_2127,N_2064);
nand U2355 (N_2355,N_2075,N_2193);
nand U2356 (N_2356,N_2041,N_2095);
and U2357 (N_2357,N_2017,N_2007);
nand U2358 (N_2358,N_2121,N_2192);
nand U2359 (N_2359,N_2133,N_2132);
and U2360 (N_2360,N_2097,N_2111);
nand U2361 (N_2361,N_2123,N_2149);
xnor U2362 (N_2362,N_2068,N_2073);
nand U2363 (N_2363,N_2028,N_2109);
nor U2364 (N_2364,N_2086,N_2067);
nor U2365 (N_2365,N_2141,N_2048);
nand U2366 (N_2366,N_2038,N_2135);
nor U2367 (N_2367,N_2104,N_2004);
nor U2368 (N_2368,N_2112,N_2077);
and U2369 (N_2369,N_2023,N_2065);
nand U2370 (N_2370,N_2168,N_2057);
nor U2371 (N_2371,N_2012,N_2157);
xnor U2372 (N_2372,N_2066,N_2035);
nand U2373 (N_2373,N_2061,N_2097);
xor U2374 (N_2374,N_2113,N_2191);
or U2375 (N_2375,N_2124,N_2082);
and U2376 (N_2376,N_2060,N_2044);
nand U2377 (N_2377,N_2188,N_2051);
nor U2378 (N_2378,N_2026,N_2049);
or U2379 (N_2379,N_2021,N_2125);
nand U2380 (N_2380,N_2114,N_2159);
xnor U2381 (N_2381,N_2129,N_2029);
xnor U2382 (N_2382,N_2107,N_2177);
nor U2383 (N_2383,N_2117,N_2090);
nor U2384 (N_2384,N_2034,N_2119);
nor U2385 (N_2385,N_2062,N_2097);
and U2386 (N_2386,N_2071,N_2029);
or U2387 (N_2387,N_2193,N_2129);
or U2388 (N_2388,N_2141,N_2181);
xor U2389 (N_2389,N_2146,N_2121);
and U2390 (N_2390,N_2115,N_2187);
and U2391 (N_2391,N_2130,N_2106);
xor U2392 (N_2392,N_2153,N_2096);
nand U2393 (N_2393,N_2039,N_2050);
nand U2394 (N_2394,N_2120,N_2089);
xor U2395 (N_2395,N_2085,N_2026);
or U2396 (N_2396,N_2119,N_2037);
nor U2397 (N_2397,N_2049,N_2057);
and U2398 (N_2398,N_2181,N_2057);
nand U2399 (N_2399,N_2183,N_2051);
nor U2400 (N_2400,N_2301,N_2267);
nor U2401 (N_2401,N_2383,N_2264);
nand U2402 (N_2402,N_2266,N_2325);
xnor U2403 (N_2403,N_2307,N_2385);
and U2404 (N_2404,N_2349,N_2243);
and U2405 (N_2405,N_2255,N_2220);
and U2406 (N_2406,N_2276,N_2240);
or U2407 (N_2407,N_2358,N_2225);
nand U2408 (N_2408,N_2208,N_2369);
nor U2409 (N_2409,N_2226,N_2275);
and U2410 (N_2410,N_2363,N_2212);
nand U2411 (N_2411,N_2206,N_2234);
or U2412 (N_2412,N_2392,N_2277);
xnor U2413 (N_2413,N_2390,N_2273);
and U2414 (N_2414,N_2218,N_2354);
or U2415 (N_2415,N_2377,N_2305);
and U2416 (N_2416,N_2253,N_2360);
nand U2417 (N_2417,N_2394,N_2330);
nand U2418 (N_2418,N_2357,N_2319);
nand U2419 (N_2419,N_2329,N_2343);
nor U2420 (N_2420,N_2219,N_2346);
nand U2421 (N_2421,N_2335,N_2387);
nor U2422 (N_2422,N_2374,N_2283);
xnor U2423 (N_2423,N_2250,N_2202);
xnor U2424 (N_2424,N_2282,N_2322);
nor U2425 (N_2425,N_2396,N_2236);
nand U2426 (N_2426,N_2274,N_2367);
nand U2427 (N_2427,N_2316,N_2263);
and U2428 (N_2428,N_2365,N_2291);
xor U2429 (N_2429,N_2313,N_2362);
and U2430 (N_2430,N_2295,N_2359);
xor U2431 (N_2431,N_2303,N_2306);
and U2432 (N_2432,N_2389,N_2222);
or U2433 (N_2433,N_2397,N_2270);
xor U2434 (N_2434,N_2210,N_2217);
and U2435 (N_2435,N_2294,N_2355);
nand U2436 (N_2436,N_2381,N_2378);
nand U2437 (N_2437,N_2333,N_2249);
and U2438 (N_2438,N_2284,N_2371);
nor U2439 (N_2439,N_2379,N_2347);
or U2440 (N_2440,N_2399,N_2344);
nor U2441 (N_2441,N_2321,N_2289);
and U2442 (N_2442,N_2304,N_2233);
and U2443 (N_2443,N_2352,N_2293);
nor U2444 (N_2444,N_2292,N_2272);
nor U2445 (N_2445,N_2256,N_2311);
or U2446 (N_2446,N_2336,N_2258);
or U2447 (N_2447,N_2265,N_2364);
or U2448 (N_2448,N_2298,N_2315);
and U2449 (N_2449,N_2280,N_2310);
nor U2450 (N_2450,N_2224,N_2228);
xor U2451 (N_2451,N_2286,N_2260);
nand U2452 (N_2452,N_2238,N_2393);
and U2453 (N_2453,N_2327,N_2376);
and U2454 (N_2454,N_2351,N_2215);
xnor U2455 (N_2455,N_2262,N_2353);
xor U2456 (N_2456,N_2341,N_2302);
xnor U2457 (N_2457,N_2361,N_2342);
nor U2458 (N_2458,N_2388,N_2320);
xor U2459 (N_2459,N_2398,N_2259);
or U2460 (N_2460,N_2382,N_2391);
nand U2461 (N_2461,N_2334,N_2268);
and U2462 (N_2462,N_2247,N_2384);
nor U2463 (N_2463,N_2241,N_2296);
and U2464 (N_2464,N_2395,N_2242);
and U2465 (N_2465,N_2380,N_2257);
nand U2466 (N_2466,N_2309,N_2211);
nand U2467 (N_2467,N_2339,N_2245);
and U2468 (N_2468,N_2278,N_2223);
or U2469 (N_2469,N_2288,N_2231);
nor U2470 (N_2470,N_2230,N_2386);
and U2471 (N_2471,N_2297,N_2201);
xnor U2472 (N_2472,N_2200,N_2237);
xnor U2473 (N_2473,N_2299,N_2323);
nor U2474 (N_2474,N_2239,N_2205);
nor U2475 (N_2475,N_2269,N_2332);
or U2476 (N_2476,N_2350,N_2368);
or U2477 (N_2477,N_2232,N_2216);
nand U2478 (N_2478,N_2317,N_2300);
nand U2479 (N_2479,N_2235,N_2227);
nand U2480 (N_2480,N_2326,N_2328);
and U2481 (N_2481,N_2281,N_2366);
xnor U2482 (N_2482,N_2287,N_2221);
nor U2483 (N_2483,N_2254,N_2312);
nor U2484 (N_2484,N_2203,N_2340);
or U2485 (N_2485,N_2370,N_2348);
or U2486 (N_2486,N_2279,N_2290);
nand U2487 (N_2487,N_2356,N_2331);
nor U2488 (N_2488,N_2285,N_2324);
nand U2489 (N_2489,N_2261,N_2204);
or U2490 (N_2490,N_2244,N_2252);
xor U2491 (N_2491,N_2318,N_2251);
xnor U2492 (N_2492,N_2372,N_2308);
xor U2493 (N_2493,N_2214,N_2337);
xor U2494 (N_2494,N_2373,N_2209);
or U2495 (N_2495,N_2213,N_2248);
xor U2496 (N_2496,N_2338,N_2345);
or U2497 (N_2497,N_2375,N_2207);
and U2498 (N_2498,N_2271,N_2229);
and U2499 (N_2499,N_2314,N_2246);
xnor U2500 (N_2500,N_2313,N_2325);
nor U2501 (N_2501,N_2391,N_2276);
or U2502 (N_2502,N_2380,N_2251);
nor U2503 (N_2503,N_2248,N_2305);
xor U2504 (N_2504,N_2226,N_2205);
xnor U2505 (N_2505,N_2347,N_2389);
and U2506 (N_2506,N_2249,N_2270);
nor U2507 (N_2507,N_2391,N_2200);
nor U2508 (N_2508,N_2351,N_2352);
and U2509 (N_2509,N_2259,N_2225);
nor U2510 (N_2510,N_2221,N_2214);
nor U2511 (N_2511,N_2399,N_2231);
or U2512 (N_2512,N_2396,N_2321);
nand U2513 (N_2513,N_2208,N_2214);
nor U2514 (N_2514,N_2380,N_2356);
nor U2515 (N_2515,N_2286,N_2284);
xor U2516 (N_2516,N_2376,N_2340);
and U2517 (N_2517,N_2348,N_2295);
nand U2518 (N_2518,N_2383,N_2266);
or U2519 (N_2519,N_2342,N_2375);
and U2520 (N_2520,N_2281,N_2273);
xnor U2521 (N_2521,N_2278,N_2308);
xor U2522 (N_2522,N_2273,N_2234);
and U2523 (N_2523,N_2357,N_2362);
or U2524 (N_2524,N_2373,N_2357);
nor U2525 (N_2525,N_2295,N_2283);
nor U2526 (N_2526,N_2377,N_2225);
and U2527 (N_2527,N_2218,N_2272);
xnor U2528 (N_2528,N_2388,N_2386);
nand U2529 (N_2529,N_2220,N_2285);
xor U2530 (N_2530,N_2306,N_2382);
and U2531 (N_2531,N_2278,N_2345);
or U2532 (N_2532,N_2268,N_2220);
xor U2533 (N_2533,N_2390,N_2287);
or U2534 (N_2534,N_2266,N_2332);
nand U2535 (N_2535,N_2352,N_2230);
nor U2536 (N_2536,N_2229,N_2252);
nor U2537 (N_2537,N_2322,N_2230);
nor U2538 (N_2538,N_2345,N_2289);
xnor U2539 (N_2539,N_2352,N_2277);
xor U2540 (N_2540,N_2362,N_2277);
nor U2541 (N_2541,N_2370,N_2312);
xnor U2542 (N_2542,N_2314,N_2396);
nand U2543 (N_2543,N_2317,N_2233);
or U2544 (N_2544,N_2209,N_2252);
or U2545 (N_2545,N_2299,N_2284);
nor U2546 (N_2546,N_2213,N_2208);
and U2547 (N_2547,N_2389,N_2300);
xnor U2548 (N_2548,N_2284,N_2273);
or U2549 (N_2549,N_2221,N_2335);
or U2550 (N_2550,N_2284,N_2334);
and U2551 (N_2551,N_2254,N_2315);
and U2552 (N_2552,N_2229,N_2311);
and U2553 (N_2553,N_2329,N_2328);
xor U2554 (N_2554,N_2366,N_2219);
and U2555 (N_2555,N_2397,N_2366);
xor U2556 (N_2556,N_2353,N_2272);
nand U2557 (N_2557,N_2264,N_2260);
or U2558 (N_2558,N_2308,N_2384);
or U2559 (N_2559,N_2222,N_2398);
nand U2560 (N_2560,N_2316,N_2294);
or U2561 (N_2561,N_2351,N_2341);
nand U2562 (N_2562,N_2279,N_2261);
nor U2563 (N_2563,N_2218,N_2246);
xnor U2564 (N_2564,N_2238,N_2369);
and U2565 (N_2565,N_2376,N_2280);
and U2566 (N_2566,N_2320,N_2286);
nand U2567 (N_2567,N_2226,N_2290);
and U2568 (N_2568,N_2283,N_2342);
xor U2569 (N_2569,N_2285,N_2373);
and U2570 (N_2570,N_2387,N_2318);
or U2571 (N_2571,N_2361,N_2276);
xor U2572 (N_2572,N_2255,N_2246);
nor U2573 (N_2573,N_2243,N_2353);
or U2574 (N_2574,N_2266,N_2362);
nor U2575 (N_2575,N_2363,N_2347);
nand U2576 (N_2576,N_2215,N_2275);
nor U2577 (N_2577,N_2369,N_2298);
nand U2578 (N_2578,N_2276,N_2225);
or U2579 (N_2579,N_2375,N_2297);
xor U2580 (N_2580,N_2315,N_2324);
or U2581 (N_2581,N_2210,N_2250);
xnor U2582 (N_2582,N_2233,N_2236);
nand U2583 (N_2583,N_2269,N_2344);
xor U2584 (N_2584,N_2305,N_2239);
nor U2585 (N_2585,N_2212,N_2288);
nand U2586 (N_2586,N_2393,N_2260);
and U2587 (N_2587,N_2335,N_2319);
xnor U2588 (N_2588,N_2230,N_2329);
xor U2589 (N_2589,N_2260,N_2223);
nor U2590 (N_2590,N_2220,N_2385);
nor U2591 (N_2591,N_2377,N_2244);
and U2592 (N_2592,N_2208,N_2334);
nand U2593 (N_2593,N_2297,N_2292);
nor U2594 (N_2594,N_2295,N_2249);
or U2595 (N_2595,N_2265,N_2353);
or U2596 (N_2596,N_2336,N_2365);
xnor U2597 (N_2597,N_2316,N_2201);
or U2598 (N_2598,N_2360,N_2213);
xor U2599 (N_2599,N_2399,N_2224);
nor U2600 (N_2600,N_2482,N_2471);
nor U2601 (N_2601,N_2416,N_2515);
or U2602 (N_2602,N_2584,N_2583);
and U2603 (N_2603,N_2441,N_2594);
or U2604 (N_2604,N_2571,N_2585);
or U2605 (N_2605,N_2458,N_2563);
xnor U2606 (N_2606,N_2470,N_2581);
and U2607 (N_2607,N_2525,N_2503);
nand U2608 (N_2608,N_2550,N_2445);
nand U2609 (N_2609,N_2436,N_2549);
nand U2610 (N_2610,N_2444,N_2423);
or U2611 (N_2611,N_2454,N_2501);
and U2612 (N_2612,N_2415,N_2505);
xnor U2613 (N_2613,N_2517,N_2590);
nor U2614 (N_2614,N_2481,N_2464);
or U2615 (N_2615,N_2559,N_2476);
and U2616 (N_2616,N_2452,N_2430);
nor U2617 (N_2617,N_2534,N_2554);
and U2618 (N_2618,N_2480,N_2478);
nand U2619 (N_2619,N_2558,N_2544);
nor U2620 (N_2620,N_2440,N_2417);
or U2621 (N_2621,N_2443,N_2466);
and U2622 (N_2622,N_2492,N_2455);
nor U2623 (N_2623,N_2516,N_2493);
nor U2624 (N_2624,N_2530,N_2513);
or U2625 (N_2625,N_2403,N_2420);
nor U2626 (N_2626,N_2541,N_2487);
or U2627 (N_2627,N_2456,N_2461);
nor U2628 (N_2628,N_2555,N_2446);
nand U2629 (N_2629,N_2553,N_2514);
nand U2630 (N_2630,N_2404,N_2457);
or U2631 (N_2631,N_2485,N_2488);
nor U2632 (N_2632,N_2406,N_2546);
nand U2633 (N_2633,N_2483,N_2539);
nor U2634 (N_2634,N_2469,N_2599);
or U2635 (N_2635,N_2498,N_2477);
or U2636 (N_2636,N_2459,N_2576);
nand U2637 (N_2637,N_2465,N_2491);
and U2638 (N_2638,N_2543,N_2568);
and U2639 (N_2639,N_2591,N_2410);
or U2640 (N_2640,N_2588,N_2405);
and U2641 (N_2641,N_2523,N_2486);
nand U2642 (N_2642,N_2418,N_2527);
or U2643 (N_2643,N_2435,N_2460);
nand U2644 (N_2644,N_2518,N_2521);
or U2645 (N_2645,N_2542,N_2596);
nand U2646 (N_2646,N_2531,N_2421);
nor U2647 (N_2647,N_2507,N_2439);
nand U2648 (N_2648,N_2598,N_2448);
and U2649 (N_2649,N_2475,N_2575);
and U2650 (N_2650,N_2522,N_2556);
xor U2651 (N_2651,N_2536,N_2538);
nand U2652 (N_2652,N_2520,N_2597);
nor U2653 (N_2653,N_2533,N_2426);
nand U2654 (N_2654,N_2592,N_2562);
and U2655 (N_2655,N_2552,N_2508);
xnor U2656 (N_2656,N_2411,N_2472);
xnor U2657 (N_2657,N_2431,N_2506);
and U2658 (N_2658,N_2408,N_2565);
nor U2659 (N_2659,N_2422,N_2560);
or U2660 (N_2660,N_2499,N_2402);
nor U2661 (N_2661,N_2551,N_2494);
xor U2662 (N_2662,N_2548,N_2427);
nor U2663 (N_2663,N_2407,N_2529);
xor U2664 (N_2664,N_2409,N_2587);
xor U2665 (N_2665,N_2557,N_2489);
xor U2666 (N_2666,N_2526,N_2545);
nor U2667 (N_2667,N_2467,N_2569);
nand U2668 (N_2668,N_2442,N_2561);
nand U2669 (N_2669,N_2400,N_2462);
nor U2670 (N_2670,N_2474,N_2425);
and U2671 (N_2671,N_2484,N_2570);
nand U2672 (N_2672,N_2412,N_2589);
nor U2673 (N_2673,N_2429,N_2579);
xnor U2674 (N_2674,N_2500,N_2490);
xor U2675 (N_2675,N_2519,N_2453);
or U2676 (N_2676,N_2566,N_2509);
and U2677 (N_2677,N_2511,N_2413);
nor U2678 (N_2678,N_2547,N_2540);
xor U2679 (N_2679,N_2432,N_2473);
and U2680 (N_2680,N_2449,N_2578);
or U2681 (N_2681,N_2512,N_2468);
xnor U2682 (N_2682,N_2586,N_2535);
nor U2683 (N_2683,N_2414,N_2447);
xnor U2684 (N_2684,N_2577,N_2573);
nand U2685 (N_2685,N_2433,N_2450);
nor U2686 (N_2686,N_2567,N_2593);
and U2687 (N_2687,N_2463,N_2438);
or U2688 (N_2688,N_2532,N_2479);
nand U2689 (N_2689,N_2574,N_2497);
or U2690 (N_2690,N_2572,N_2401);
nor U2691 (N_2691,N_2528,N_2434);
or U2692 (N_2692,N_2595,N_2451);
or U2693 (N_2693,N_2495,N_2582);
or U2694 (N_2694,N_2496,N_2437);
xnor U2695 (N_2695,N_2504,N_2564);
nor U2696 (N_2696,N_2510,N_2580);
nor U2697 (N_2697,N_2524,N_2424);
xnor U2698 (N_2698,N_2428,N_2537);
or U2699 (N_2699,N_2502,N_2419);
nand U2700 (N_2700,N_2429,N_2521);
nand U2701 (N_2701,N_2496,N_2532);
and U2702 (N_2702,N_2598,N_2469);
or U2703 (N_2703,N_2585,N_2565);
nand U2704 (N_2704,N_2536,N_2441);
and U2705 (N_2705,N_2449,N_2440);
or U2706 (N_2706,N_2573,N_2525);
nor U2707 (N_2707,N_2507,N_2500);
or U2708 (N_2708,N_2510,N_2568);
nand U2709 (N_2709,N_2494,N_2525);
nor U2710 (N_2710,N_2543,N_2440);
and U2711 (N_2711,N_2567,N_2487);
nand U2712 (N_2712,N_2407,N_2419);
nor U2713 (N_2713,N_2517,N_2559);
xor U2714 (N_2714,N_2420,N_2411);
nand U2715 (N_2715,N_2563,N_2478);
and U2716 (N_2716,N_2574,N_2460);
nor U2717 (N_2717,N_2552,N_2405);
nor U2718 (N_2718,N_2459,N_2546);
and U2719 (N_2719,N_2421,N_2583);
nand U2720 (N_2720,N_2494,N_2427);
nand U2721 (N_2721,N_2493,N_2546);
nor U2722 (N_2722,N_2513,N_2562);
nand U2723 (N_2723,N_2584,N_2412);
xor U2724 (N_2724,N_2429,N_2587);
and U2725 (N_2725,N_2573,N_2550);
and U2726 (N_2726,N_2590,N_2528);
or U2727 (N_2727,N_2500,N_2438);
xor U2728 (N_2728,N_2431,N_2517);
nand U2729 (N_2729,N_2592,N_2517);
nand U2730 (N_2730,N_2443,N_2559);
nand U2731 (N_2731,N_2406,N_2467);
or U2732 (N_2732,N_2586,N_2590);
or U2733 (N_2733,N_2428,N_2518);
nor U2734 (N_2734,N_2511,N_2499);
and U2735 (N_2735,N_2409,N_2456);
or U2736 (N_2736,N_2588,N_2437);
or U2737 (N_2737,N_2558,N_2409);
or U2738 (N_2738,N_2525,N_2400);
xnor U2739 (N_2739,N_2529,N_2436);
or U2740 (N_2740,N_2423,N_2570);
and U2741 (N_2741,N_2578,N_2550);
and U2742 (N_2742,N_2446,N_2468);
xnor U2743 (N_2743,N_2598,N_2415);
nor U2744 (N_2744,N_2536,N_2558);
nand U2745 (N_2745,N_2410,N_2508);
and U2746 (N_2746,N_2569,N_2423);
and U2747 (N_2747,N_2427,N_2438);
and U2748 (N_2748,N_2429,N_2481);
nor U2749 (N_2749,N_2443,N_2497);
nor U2750 (N_2750,N_2472,N_2595);
xor U2751 (N_2751,N_2459,N_2578);
xor U2752 (N_2752,N_2461,N_2508);
nand U2753 (N_2753,N_2555,N_2523);
nor U2754 (N_2754,N_2572,N_2538);
or U2755 (N_2755,N_2486,N_2439);
xor U2756 (N_2756,N_2465,N_2577);
and U2757 (N_2757,N_2474,N_2401);
nand U2758 (N_2758,N_2537,N_2575);
xnor U2759 (N_2759,N_2497,N_2412);
xnor U2760 (N_2760,N_2475,N_2585);
nor U2761 (N_2761,N_2500,N_2475);
and U2762 (N_2762,N_2421,N_2576);
or U2763 (N_2763,N_2407,N_2425);
and U2764 (N_2764,N_2488,N_2533);
and U2765 (N_2765,N_2420,N_2493);
and U2766 (N_2766,N_2468,N_2522);
nand U2767 (N_2767,N_2534,N_2563);
and U2768 (N_2768,N_2477,N_2503);
nand U2769 (N_2769,N_2576,N_2519);
nor U2770 (N_2770,N_2470,N_2559);
nor U2771 (N_2771,N_2479,N_2551);
nand U2772 (N_2772,N_2546,N_2579);
nor U2773 (N_2773,N_2565,N_2550);
and U2774 (N_2774,N_2444,N_2577);
and U2775 (N_2775,N_2477,N_2412);
nor U2776 (N_2776,N_2422,N_2493);
nor U2777 (N_2777,N_2571,N_2466);
and U2778 (N_2778,N_2568,N_2582);
and U2779 (N_2779,N_2495,N_2516);
nand U2780 (N_2780,N_2503,N_2407);
xor U2781 (N_2781,N_2408,N_2529);
or U2782 (N_2782,N_2447,N_2452);
or U2783 (N_2783,N_2540,N_2582);
nor U2784 (N_2784,N_2581,N_2583);
or U2785 (N_2785,N_2537,N_2526);
or U2786 (N_2786,N_2589,N_2424);
nor U2787 (N_2787,N_2438,N_2498);
nand U2788 (N_2788,N_2422,N_2459);
xnor U2789 (N_2789,N_2547,N_2520);
and U2790 (N_2790,N_2561,N_2546);
and U2791 (N_2791,N_2515,N_2446);
nand U2792 (N_2792,N_2515,N_2473);
or U2793 (N_2793,N_2444,N_2589);
nand U2794 (N_2794,N_2580,N_2458);
and U2795 (N_2795,N_2445,N_2545);
nand U2796 (N_2796,N_2504,N_2452);
nand U2797 (N_2797,N_2569,N_2479);
xnor U2798 (N_2798,N_2492,N_2437);
nand U2799 (N_2799,N_2432,N_2581);
and U2800 (N_2800,N_2797,N_2783);
and U2801 (N_2801,N_2656,N_2666);
nand U2802 (N_2802,N_2628,N_2609);
nand U2803 (N_2803,N_2720,N_2678);
nand U2804 (N_2804,N_2690,N_2646);
or U2805 (N_2805,N_2695,N_2652);
nor U2806 (N_2806,N_2795,N_2698);
nor U2807 (N_2807,N_2703,N_2709);
nand U2808 (N_2808,N_2757,N_2626);
nand U2809 (N_2809,N_2710,N_2764);
xor U2810 (N_2810,N_2642,N_2779);
or U2811 (N_2811,N_2776,N_2692);
xor U2812 (N_2812,N_2699,N_2714);
nor U2813 (N_2813,N_2693,N_2706);
nand U2814 (N_2814,N_2772,N_2702);
and U2815 (N_2815,N_2665,N_2736);
and U2816 (N_2816,N_2613,N_2713);
nand U2817 (N_2817,N_2791,N_2653);
or U2818 (N_2818,N_2740,N_2634);
nand U2819 (N_2819,N_2615,N_2700);
or U2820 (N_2820,N_2681,N_2694);
nor U2821 (N_2821,N_2729,N_2605);
nor U2822 (N_2822,N_2667,N_2688);
nor U2823 (N_2823,N_2662,N_2600);
nand U2824 (N_2824,N_2773,N_2668);
and U2825 (N_2825,N_2731,N_2610);
or U2826 (N_2826,N_2601,N_2796);
or U2827 (N_2827,N_2670,N_2682);
nand U2828 (N_2828,N_2673,N_2753);
nor U2829 (N_2829,N_2739,N_2616);
nor U2830 (N_2830,N_2781,N_2606);
nand U2831 (N_2831,N_2743,N_2689);
or U2832 (N_2832,N_2683,N_2766);
nand U2833 (N_2833,N_2786,N_2798);
nor U2834 (N_2834,N_2684,N_2770);
nor U2835 (N_2835,N_2658,N_2633);
nor U2836 (N_2836,N_2602,N_2733);
and U2837 (N_2837,N_2734,N_2732);
or U2838 (N_2838,N_2614,N_2768);
xnor U2839 (N_2839,N_2696,N_2669);
xnor U2840 (N_2840,N_2782,N_2711);
and U2841 (N_2841,N_2793,N_2778);
and U2842 (N_2842,N_2659,N_2635);
xnor U2843 (N_2843,N_2771,N_2632);
and U2844 (N_2844,N_2763,N_2686);
and U2845 (N_2845,N_2620,N_2637);
nor U2846 (N_2846,N_2676,N_2608);
and U2847 (N_2847,N_2680,N_2742);
or U2848 (N_2848,N_2737,N_2691);
nor U2849 (N_2849,N_2640,N_2752);
nand U2850 (N_2850,N_2715,N_2780);
or U2851 (N_2851,N_2627,N_2760);
xor U2852 (N_2852,N_2738,N_2777);
nor U2853 (N_2853,N_2769,N_2744);
or U2854 (N_2854,N_2749,N_2708);
nor U2855 (N_2855,N_2761,N_2765);
nand U2856 (N_2856,N_2701,N_2716);
or U2857 (N_2857,N_2636,N_2799);
and U2858 (N_2858,N_2657,N_2607);
and U2859 (N_2859,N_2604,N_2622);
and U2860 (N_2860,N_2741,N_2671);
nand U2861 (N_2861,N_2748,N_2735);
and U2862 (N_2862,N_2723,N_2630);
xnor U2863 (N_2863,N_2655,N_2641);
and U2864 (N_2864,N_2730,N_2707);
nand U2865 (N_2865,N_2724,N_2697);
nand U2866 (N_2866,N_2767,N_2664);
and U2867 (N_2867,N_2750,N_2790);
xnor U2868 (N_2868,N_2648,N_2745);
nor U2869 (N_2869,N_2631,N_2754);
nor U2870 (N_2870,N_2687,N_2788);
nor U2871 (N_2871,N_2675,N_2746);
xor U2872 (N_2872,N_2677,N_2717);
or U2873 (N_2873,N_2785,N_2756);
or U2874 (N_2874,N_2705,N_2787);
or U2875 (N_2875,N_2712,N_2651);
or U2876 (N_2876,N_2645,N_2704);
nand U2877 (N_2877,N_2718,N_2794);
nand U2878 (N_2878,N_2726,N_2654);
or U2879 (N_2879,N_2751,N_2643);
xnor U2880 (N_2880,N_2629,N_2789);
nand U2881 (N_2881,N_2612,N_2638);
nand U2882 (N_2882,N_2617,N_2660);
nand U2883 (N_2883,N_2639,N_2625);
and U2884 (N_2884,N_2611,N_2647);
nand U2885 (N_2885,N_2762,N_2663);
xor U2886 (N_2886,N_2792,N_2685);
nor U2887 (N_2887,N_2722,N_2679);
nand U2888 (N_2888,N_2603,N_2624);
nor U2889 (N_2889,N_2619,N_2618);
nand U2890 (N_2890,N_2727,N_2747);
nand U2891 (N_2891,N_2725,N_2644);
nor U2892 (N_2892,N_2649,N_2721);
nand U2893 (N_2893,N_2621,N_2784);
and U2894 (N_2894,N_2623,N_2672);
or U2895 (N_2895,N_2775,N_2728);
nor U2896 (N_2896,N_2719,N_2650);
nand U2897 (N_2897,N_2661,N_2759);
xnor U2898 (N_2898,N_2774,N_2755);
or U2899 (N_2899,N_2674,N_2758);
or U2900 (N_2900,N_2698,N_2641);
and U2901 (N_2901,N_2743,N_2668);
nor U2902 (N_2902,N_2660,N_2702);
nor U2903 (N_2903,N_2626,N_2660);
xnor U2904 (N_2904,N_2682,N_2754);
or U2905 (N_2905,N_2713,N_2766);
and U2906 (N_2906,N_2780,N_2702);
and U2907 (N_2907,N_2689,N_2705);
nor U2908 (N_2908,N_2615,N_2740);
nor U2909 (N_2909,N_2621,N_2604);
nand U2910 (N_2910,N_2734,N_2767);
nor U2911 (N_2911,N_2710,N_2773);
and U2912 (N_2912,N_2734,N_2658);
nand U2913 (N_2913,N_2652,N_2688);
or U2914 (N_2914,N_2608,N_2786);
nor U2915 (N_2915,N_2772,N_2676);
or U2916 (N_2916,N_2664,N_2633);
or U2917 (N_2917,N_2610,N_2699);
nor U2918 (N_2918,N_2735,N_2676);
xor U2919 (N_2919,N_2725,N_2673);
or U2920 (N_2920,N_2699,N_2739);
or U2921 (N_2921,N_2714,N_2689);
nand U2922 (N_2922,N_2670,N_2769);
or U2923 (N_2923,N_2664,N_2787);
and U2924 (N_2924,N_2620,N_2621);
or U2925 (N_2925,N_2605,N_2727);
or U2926 (N_2926,N_2625,N_2739);
nor U2927 (N_2927,N_2605,N_2752);
nor U2928 (N_2928,N_2600,N_2709);
xnor U2929 (N_2929,N_2786,N_2793);
or U2930 (N_2930,N_2689,N_2731);
xnor U2931 (N_2931,N_2629,N_2754);
and U2932 (N_2932,N_2656,N_2751);
nand U2933 (N_2933,N_2700,N_2634);
nand U2934 (N_2934,N_2774,N_2706);
nand U2935 (N_2935,N_2666,N_2774);
nand U2936 (N_2936,N_2795,N_2745);
nand U2937 (N_2937,N_2613,N_2736);
and U2938 (N_2938,N_2645,N_2781);
nor U2939 (N_2939,N_2738,N_2639);
or U2940 (N_2940,N_2743,N_2661);
or U2941 (N_2941,N_2690,N_2798);
nor U2942 (N_2942,N_2604,N_2786);
nor U2943 (N_2943,N_2753,N_2623);
nor U2944 (N_2944,N_2727,N_2609);
and U2945 (N_2945,N_2707,N_2630);
or U2946 (N_2946,N_2683,N_2715);
xnor U2947 (N_2947,N_2689,N_2639);
or U2948 (N_2948,N_2714,N_2795);
xor U2949 (N_2949,N_2703,N_2698);
or U2950 (N_2950,N_2654,N_2776);
nand U2951 (N_2951,N_2642,N_2687);
nor U2952 (N_2952,N_2684,N_2741);
or U2953 (N_2953,N_2791,N_2755);
nor U2954 (N_2954,N_2677,N_2682);
or U2955 (N_2955,N_2741,N_2799);
nand U2956 (N_2956,N_2657,N_2709);
nor U2957 (N_2957,N_2702,N_2622);
nor U2958 (N_2958,N_2739,N_2711);
nor U2959 (N_2959,N_2720,N_2613);
xor U2960 (N_2960,N_2685,N_2670);
nand U2961 (N_2961,N_2723,N_2762);
nor U2962 (N_2962,N_2634,N_2647);
and U2963 (N_2963,N_2747,N_2795);
xor U2964 (N_2964,N_2779,N_2787);
or U2965 (N_2965,N_2681,N_2637);
nand U2966 (N_2966,N_2667,N_2732);
or U2967 (N_2967,N_2626,N_2662);
nor U2968 (N_2968,N_2780,N_2791);
or U2969 (N_2969,N_2663,N_2781);
nor U2970 (N_2970,N_2705,N_2603);
or U2971 (N_2971,N_2704,N_2600);
nand U2972 (N_2972,N_2773,N_2730);
or U2973 (N_2973,N_2712,N_2612);
and U2974 (N_2974,N_2744,N_2662);
xnor U2975 (N_2975,N_2745,N_2608);
nand U2976 (N_2976,N_2661,N_2793);
nor U2977 (N_2977,N_2748,N_2681);
nand U2978 (N_2978,N_2720,N_2679);
and U2979 (N_2979,N_2635,N_2668);
nand U2980 (N_2980,N_2794,N_2649);
and U2981 (N_2981,N_2686,N_2768);
and U2982 (N_2982,N_2764,N_2698);
nand U2983 (N_2983,N_2648,N_2783);
or U2984 (N_2984,N_2602,N_2663);
or U2985 (N_2985,N_2666,N_2668);
nor U2986 (N_2986,N_2752,N_2659);
nand U2987 (N_2987,N_2612,N_2649);
or U2988 (N_2988,N_2647,N_2610);
xnor U2989 (N_2989,N_2616,N_2667);
nor U2990 (N_2990,N_2655,N_2723);
nor U2991 (N_2991,N_2637,N_2652);
xnor U2992 (N_2992,N_2676,N_2763);
or U2993 (N_2993,N_2746,N_2792);
or U2994 (N_2994,N_2646,N_2783);
and U2995 (N_2995,N_2637,N_2788);
nand U2996 (N_2996,N_2757,N_2692);
xor U2997 (N_2997,N_2795,N_2690);
nor U2998 (N_2998,N_2705,N_2763);
nand U2999 (N_2999,N_2778,N_2619);
nand U3000 (N_3000,N_2985,N_2978);
xnor U3001 (N_3001,N_2938,N_2833);
and U3002 (N_3002,N_2964,N_2868);
and U3003 (N_3003,N_2840,N_2910);
or U3004 (N_3004,N_2902,N_2836);
and U3005 (N_3005,N_2980,N_2862);
and U3006 (N_3006,N_2829,N_2999);
nor U3007 (N_3007,N_2888,N_2929);
xnor U3008 (N_3008,N_2903,N_2965);
and U3009 (N_3009,N_2974,N_2822);
and U3010 (N_3010,N_2852,N_2951);
or U3011 (N_3011,N_2858,N_2960);
or U3012 (N_3012,N_2893,N_2823);
xnor U3013 (N_3013,N_2826,N_2989);
nor U3014 (N_3014,N_2934,N_2907);
xnor U3015 (N_3015,N_2804,N_2877);
or U3016 (N_3016,N_2975,N_2924);
nor U3017 (N_3017,N_2966,N_2825);
or U3018 (N_3018,N_2971,N_2871);
or U3019 (N_3019,N_2905,N_2896);
nand U3020 (N_3020,N_2820,N_2879);
and U3021 (N_3021,N_2914,N_2819);
or U3022 (N_3022,N_2842,N_2863);
and U3023 (N_3023,N_2854,N_2919);
xnor U3024 (N_3024,N_2956,N_2917);
xnor U3025 (N_3025,N_2901,N_2880);
nor U3026 (N_3026,N_2831,N_2932);
nor U3027 (N_3027,N_2913,N_2982);
or U3028 (N_3028,N_2894,N_2948);
xnor U3029 (N_3029,N_2887,N_2945);
nand U3030 (N_3030,N_2940,N_2898);
nor U3031 (N_3031,N_2860,N_2806);
nor U3032 (N_3032,N_2937,N_2832);
nand U3033 (N_3033,N_2963,N_2861);
and U3034 (N_3034,N_2911,N_2977);
nor U3035 (N_3035,N_2915,N_2931);
nor U3036 (N_3036,N_2816,N_2997);
xor U3037 (N_3037,N_2812,N_2983);
and U3038 (N_3038,N_2908,N_2996);
xor U3039 (N_3039,N_2800,N_2920);
xor U3040 (N_3040,N_2853,N_2817);
and U3041 (N_3041,N_2922,N_2950);
xnor U3042 (N_3042,N_2942,N_2838);
and U3043 (N_3043,N_2815,N_2890);
nand U3044 (N_3044,N_2998,N_2874);
xor U3045 (N_3045,N_2949,N_2885);
nor U3046 (N_3046,N_2866,N_2986);
nor U3047 (N_3047,N_2904,N_2830);
xnor U3048 (N_3048,N_2848,N_2962);
nand U3049 (N_3049,N_2878,N_2943);
and U3050 (N_3050,N_2850,N_2883);
and U3051 (N_3051,N_2992,N_2946);
or U3052 (N_3052,N_2809,N_2990);
or U3053 (N_3053,N_2995,N_2926);
and U3054 (N_3054,N_2906,N_2918);
and U3055 (N_3055,N_2813,N_2936);
and U3056 (N_3056,N_2882,N_2876);
nand U3057 (N_3057,N_2891,N_2835);
nor U3058 (N_3058,N_2856,N_2969);
nor U3059 (N_3059,N_2961,N_2972);
or U3060 (N_3060,N_2941,N_2981);
and U3061 (N_3061,N_2988,N_2839);
nand U3062 (N_3062,N_2851,N_2921);
and U3063 (N_3063,N_2807,N_2846);
nand U3064 (N_3064,N_2923,N_2959);
or U3065 (N_3065,N_2873,N_2803);
nor U3066 (N_3066,N_2827,N_2805);
nor U3067 (N_3067,N_2849,N_2864);
and U3068 (N_3068,N_2814,N_2994);
or U3069 (N_3069,N_2976,N_2821);
and U3070 (N_3070,N_2953,N_2955);
nand U3071 (N_3071,N_2867,N_2884);
and U3072 (N_3072,N_2824,N_2930);
nand U3073 (N_3073,N_2828,N_2895);
or U3074 (N_3074,N_2870,N_2810);
or U3075 (N_3075,N_2855,N_2909);
xor U3076 (N_3076,N_2841,N_2818);
nand U3077 (N_3077,N_2865,N_2916);
or U3078 (N_3078,N_2958,N_2881);
and U3079 (N_3079,N_2859,N_2875);
nand U3080 (N_3080,N_2927,N_2952);
nor U3081 (N_3081,N_2933,N_2808);
xor U3082 (N_3082,N_2947,N_2900);
nand U3083 (N_3083,N_2844,N_2837);
nor U3084 (N_3084,N_2811,N_2935);
and U3085 (N_3085,N_2892,N_2967);
or U3086 (N_3086,N_2993,N_2939);
nand U3087 (N_3087,N_2968,N_2843);
nor U3088 (N_3088,N_2845,N_2984);
nor U3089 (N_3089,N_2869,N_2987);
nor U3090 (N_3090,N_2991,N_2897);
xnor U3091 (N_3091,N_2802,N_2872);
xor U3092 (N_3092,N_2970,N_2834);
xor U3093 (N_3093,N_2899,N_2886);
xor U3094 (N_3094,N_2925,N_2973);
nand U3095 (N_3095,N_2857,N_2912);
and U3096 (N_3096,N_2944,N_2889);
and U3097 (N_3097,N_2957,N_2954);
or U3098 (N_3098,N_2928,N_2979);
or U3099 (N_3099,N_2847,N_2801);
or U3100 (N_3100,N_2923,N_2816);
or U3101 (N_3101,N_2999,N_2875);
xor U3102 (N_3102,N_2814,N_2999);
nand U3103 (N_3103,N_2963,N_2844);
or U3104 (N_3104,N_2893,N_2810);
or U3105 (N_3105,N_2942,N_2854);
nand U3106 (N_3106,N_2931,N_2949);
nor U3107 (N_3107,N_2967,N_2846);
and U3108 (N_3108,N_2911,N_2892);
xnor U3109 (N_3109,N_2996,N_2853);
nand U3110 (N_3110,N_2979,N_2937);
or U3111 (N_3111,N_2819,N_2814);
nand U3112 (N_3112,N_2829,N_2896);
nand U3113 (N_3113,N_2948,N_2957);
nor U3114 (N_3114,N_2968,N_2803);
or U3115 (N_3115,N_2933,N_2803);
or U3116 (N_3116,N_2836,N_2800);
and U3117 (N_3117,N_2966,N_2858);
nand U3118 (N_3118,N_2821,N_2910);
nor U3119 (N_3119,N_2812,N_2814);
and U3120 (N_3120,N_2822,N_2976);
or U3121 (N_3121,N_2875,N_2905);
nor U3122 (N_3122,N_2954,N_2850);
and U3123 (N_3123,N_2904,N_2818);
and U3124 (N_3124,N_2886,N_2991);
nor U3125 (N_3125,N_2813,N_2942);
nor U3126 (N_3126,N_2885,N_2824);
xor U3127 (N_3127,N_2943,N_2871);
nand U3128 (N_3128,N_2857,N_2974);
nand U3129 (N_3129,N_2960,N_2860);
nand U3130 (N_3130,N_2997,N_2941);
nand U3131 (N_3131,N_2819,N_2866);
nand U3132 (N_3132,N_2926,N_2908);
and U3133 (N_3133,N_2829,N_2872);
or U3134 (N_3134,N_2999,N_2958);
nor U3135 (N_3135,N_2967,N_2819);
or U3136 (N_3136,N_2930,N_2867);
xnor U3137 (N_3137,N_2808,N_2886);
xor U3138 (N_3138,N_2964,N_2938);
or U3139 (N_3139,N_2980,N_2935);
and U3140 (N_3140,N_2804,N_2879);
nor U3141 (N_3141,N_2937,N_2921);
xnor U3142 (N_3142,N_2810,N_2809);
xor U3143 (N_3143,N_2816,N_2968);
xor U3144 (N_3144,N_2934,N_2973);
xnor U3145 (N_3145,N_2980,N_2831);
nor U3146 (N_3146,N_2956,N_2875);
xor U3147 (N_3147,N_2954,N_2828);
nor U3148 (N_3148,N_2809,N_2925);
nor U3149 (N_3149,N_2828,N_2808);
nand U3150 (N_3150,N_2974,N_2986);
nand U3151 (N_3151,N_2908,N_2842);
xnor U3152 (N_3152,N_2959,N_2805);
xnor U3153 (N_3153,N_2942,N_2895);
and U3154 (N_3154,N_2818,N_2813);
or U3155 (N_3155,N_2894,N_2966);
nand U3156 (N_3156,N_2972,N_2864);
or U3157 (N_3157,N_2971,N_2820);
nor U3158 (N_3158,N_2813,N_2999);
nand U3159 (N_3159,N_2930,N_2964);
xor U3160 (N_3160,N_2830,N_2839);
and U3161 (N_3161,N_2943,N_2859);
xnor U3162 (N_3162,N_2962,N_2867);
nor U3163 (N_3163,N_2929,N_2871);
nand U3164 (N_3164,N_2942,N_2848);
xor U3165 (N_3165,N_2887,N_2849);
and U3166 (N_3166,N_2885,N_2875);
nand U3167 (N_3167,N_2888,N_2904);
or U3168 (N_3168,N_2850,N_2990);
nor U3169 (N_3169,N_2995,N_2855);
nor U3170 (N_3170,N_2971,N_2915);
or U3171 (N_3171,N_2887,N_2966);
nand U3172 (N_3172,N_2849,N_2861);
nor U3173 (N_3173,N_2911,N_2816);
nor U3174 (N_3174,N_2871,N_2964);
or U3175 (N_3175,N_2989,N_2832);
nand U3176 (N_3176,N_2995,N_2993);
xor U3177 (N_3177,N_2969,N_2885);
or U3178 (N_3178,N_2991,N_2954);
or U3179 (N_3179,N_2894,N_2863);
or U3180 (N_3180,N_2807,N_2968);
and U3181 (N_3181,N_2969,N_2813);
and U3182 (N_3182,N_2803,N_2892);
and U3183 (N_3183,N_2953,N_2829);
nand U3184 (N_3184,N_2918,N_2881);
and U3185 (N_3185,N_2890,N_2863);
nand U3186 (N_3186,N_2985,N_2972);
nor U3187 (N_3187,N_2964,N_2834);
xor U3188 (N_3188,N_2831,N_2978);
and U3189 (N_3189,N_2846,N_2836);
xor U3190 (N_3190,N_2980,N_2826);
nor U3191 (N_3191,N_2835,N_2833);
or U3192 (N_3192,N_2815,N_2839);
nand U3193 (N_3193,N_2950,N_2915);
nor U3194 (N_3194,N_2885,N_2814);
nor U3195 (N_3195,N_2982,N_2854);
and U3196 (N_3196,N_2929,N_2811);
xnor U3197 (N_3197,N_2976,N_2993);
nor U3198 (N_3198,N_2835,N_2927);
nor U3199 (N_3199,N_2840,N_2976);
nor U3200 (N_3200,N_3148,N_3177);
xnor U3201 (N_3201,N_3008,N_3184);
xor U3202 (N_3202,N_3039,N_3188);
xor U3203 (N_3203,N_3066,N_3053);
xor U3204 (N_3204,N_3116,N_3195);
and U3205 (N_3205,N_3046,N_3151);
and U3206 (N_3206,N_3145,N_3182);
or U3207 (N_3207,N_3098,N_3118);
nand U3208 (N_3208,N_3005,N_3189);
or U3209 (N_3209,N_3104,N_3120);
nor U3210 (N_3210,N_3006,N_3028);
and U3211 (N_3211,N_3001,N_3067);
and U3212 (N_3212,N_3150,N_3009);
or U3213 (N_3213,N_3147,N_3134);
and U3214 (N_3214,N_3157,N_3156);
or U3215 (N_3215,N_3024,N_3171);
xor U3216 (N_3216,N_3063,N_3136);
or U3217 (N_3217,N_3130,N_3004);
and U3218 (N_3218,N_3140,N_3115);
nand U3219 (N_3219,N_3198,N_3010);
xnor U3220 (N_3220,N_3146,N_3161);
and U3221 (N_3221,N_3026,N_3035);
or U3222 (N_3222,N_3091,N_3094);
xor U3223 (N_3223,N_3111,N_3129);
xor U3224 (N_3224,N_3190,N_3183);
xor U3225 (N_3225,N_3128,N_3057);
nand U3226 (N_3226,N_3126,N_3163);
or U3227 (N_3227,N_3034,N_3084);
or U3228 (N_3228,N_3194,N_3187);
and U3229 (N_3229,N_3139,N_3062);
xor U3230 (N_3230,N_3080,N_3032);
or U3231 (N_3231,N_3107,N_3090);
xnor U3232 (N_3232,N_3133,N_3162);
or U3233 (N_3233,N_3123,N_3119);
nand U3234 (N_3234,N_3153,N_3007);
and U3235 (N_3235,N_3054,N_3127);
and U3236 (N_3236,N_3180,N_3011);
nand U3237 (N_3237,N_3052,N_3160);
and U3238 (N_3238,N_3103,N_3099);
or U3239 (N_3239,N_3017,N_3154);
xor U3240 (N_3240,N_3113,N_3106);
nor U3241 (N_3241,N_3027,N_3138);
nor U3242 (N_3242,N_3131,N_3038);
or U3243 (N_3243,N_3045,N_3051);
xnor U3244 (N_3244,N_3020,N_3072);
or U3245 (N_3245,N_3108,N_3141);
or U3246 (N_3246,N_3077,N_3070);
or U3247 (N_3247,N_3081,N_3043);
nand U3248 (N_3248,N_3036,N_3093);
xor U3249 (N_3249,N_3117,N_3186);
nand U3250 (N_3250,N_3155,N_3199);
nor U3251 (N_3251,N_3073,N_3074);
xor U3252 (N_3252,N_3078,N_3029);
nor U3253 (N_3253,N_3076,N_3168);
and U3254 (N_3254,N_3065,N_3170);
nand U3255 (N_3255,N_3031,N_3089);
nand U3256 (N_3256,N_3149,N_3030);
or U3257 (N_3257,N_3064,N_3087);
and U3258 (N_3258,N_3164,N_3042);
and U3259 (N_3259,N_3105,N_3112);
nand U3260 (N_3260,N_3025,N_3176);
and U3261 (N_3261,N_3191,N_3092);
or U3262 (N_3262,N_3012,N_3100);
nor U3263 (N_3263,N_3000,N_3055);
or U3264 (N_3264,N_3037,N_3069);
or U3265 (N_3265,N_3060,N_3088);
nand U3266 (N_3266,N_3178,N_3173);
and U3267 (N_3267,N_3110,N_3049);
xor U3268 (N_3268,N_3068,N_3152);
or U3269 (N_3269,N_3058,N_3075);
and U3270 (N_3270,N_3014,N_3048);
or U3271 (N_3271,N_3079,N_3193);
xor U3272 (N_3272,N_3144,N_3158);
or U3273 (N_3273,N_3125,N_3083);
nor U3274 (N_3274,N_3015,N_3121);
and U3275 (N_3275,N_3085,N_3101);
and U3276 (N_3276,N_3135,N_3022);
xnor U3277 (N_3277,N_3102,N_3023);
and U3278 (N_3278,N_3095,N_3142);
nor U3279 (N_3279,N_3175,N_3050);
nor U3280 (N_3280,N_3021,N_3013);
and U3281 (N_3281,N_3061,N_3033);
or U3282 (N_3282,N_3174,N_3196);
xnor U3283 (N_3283,N_3003,N_3181);
nor U3284 (N_3284,N_3086,N_3002);
and U3285 (N_3285,N_3019,N_3018);
xnor U3286 (N_3286,N_3179,N_3109);
xor U3287 (N_3287,N_3114,N_3167);
xnor U3288 (N_3288,N_3082,N_3047);
nand U3289 (N_3289,N_3122,N_3172);
or U3290 (N_3290,N_3192,N_3071);
nor U3291 (N_3291,N_3132,N_3143);
and U3292 (N_3292,N_3040,N_3044);
xnor U3293 (N_3293,N_3137,N_3185);
nand U3294 (N_3294,N_3097,N_3041);
nor U3295 (N_3295,N_3059,N_3166);
xor U3296 (N_3296,N_3197,N_3169);
xnor U3297 (N_3297,N_3096,N_3165);
or U3298 (N_3298,N_3124,N_3016);
nor U3299 (N_3299,N_3159,N_3056);
or U3300 (N_3300,N_3158,N_3056);
and U3301 (N_3301,N_3010,N_3021);
nand U3302 (N_3302,N_3084,N_3080);
xor U3303 (N_3303,N_3071,N_3110);
nand U3304 (N_3304,N_3126,N_3189);
or U3305 (N_3305,N_3110,N_3074);
xnor U3306 (N_3306,N_3053,N_3092);
nor U3307 (N_3307,N_3155,N_3046);
or U3308 (N_3308,N_3171,N_3103);
nor U3309 (N_3309,N_3042,N_3064);
nor U3310 (N_3310,N_3043,N_3065);
nor U3311 (N_3311,N_3130,N_3027);
and U3312 (N_3312,N_3014,N_3184);
and U3313 (N_3313,N_3081,N_3024);
xor U3314 (N_3314,N_3019,N_3007);
xor U3315 (N_3315,N_3038,N_3072);
nand U3316 (N_3316,N_3010,N_3050);
nand U3317 (N_3317,N_3116,N_3075);
or U3318 (N_3318,N_3009,N_3142);
nand U3319 (N_3319,N_3054,N_3181);
and U3320 (N_3320,N_3012,N_3148);
and U3321 (N_3321,N_3097,N_3035);
nor U3322 (N_3322,N_3072,N_3160);
xor U3323 (N_3323,N_3066,N_3166);
xnor U3324 (N_3324,N_3054,N_3083);
nand U3325 (N_3325,N_3043,N_3097);
or U3326 (N_3326,N_3164,N_3189);
or U3327 (N_3327,N_3177,N_3019);
or U3328 (N_3328,N_3168,N_3077);
nand U3329 (N_3329,N_3108,N_3084);
xnor U3330 (N_3330,N_3028,N_3011);
and U3331 (N_3331,N_3084,N_3113);
and U3332 (N_3332,N_3115,N_3016);
xor U3333 (N_3333,N_3197,N_3012);
and U3334 (N_3334,N_3129,N_3071);
or U3335 (N_3335,N_3054,N_3086);
and U3336 (N_3336,N_3173,N_3053);
and U3337 (N_3337,N_3175,N_3038);
nor U3338 (N_3338,N_3125,N_3165);
nor U3339 (N_3339,N_3118,N_3184);
nor U3340 (N_3340,N_3014,N_3026);
and U3341 (N_3341,N_3199,N_3149);
or U3342 (N_3342,N_3011,N_3143);
or U3343 (N_3343,N_3193,N_3021);
xor U3344 (N_3344,N_3006,N_3115);
nor U3345 (N_3345,N_3029,N_3007);
xor U3346 (N_3346,N_3089,N_3191);
and U3347 (N_3347,N_3005,N_3017);
nor U3348 (N_3348,N_3089,N_3006);
nand U3349 (N_3349,N_3002,N_3159);
nor U3350 (N_3350,N_3154,N_3027);
and U3351 (N_3351,N_3152,N_3143);
and U3352 (N_3352,N_3016,N_3037);
nand U3353 (N_3353,N_3094,N_3098);
and U3354 (N_3354,N_3048,N_3031);
or U3355 (N_3355,N_3176,N_3158);
nor U3356 (N_3356,N_3162,N_3117);
xnor U3357 (N_3357,N_3070,N_3169);
xnor U3358 (N_3358,N_3106,N_3151);
nand U3359 (N_3359,N_3146,N_3087);
or U3360 (N_3360,N_3028,N_3035);
nand U3361 (N_3361,N_3054,N_3007);
nor U3362 (N_3362,N_3173,N_3032);
or U3363 (N_3363,N_3192,N_3093);
or U3364 (N_3364,N_3039,N_3165);
or U3365 (N_3365,N_3143,N_3190);
nand U3366 (N_3366,N_3114,N_3000);
nor U3367 (N_3367,N_3145,N_3172);
xor U3368 (N_3368,N_3043,N_3067);
or U3369 (N_3369,N_3144,N_3113);
nor U3370 (N_3370,N_3052,N_3189);
nor U3371 (N_3371,N_3035,N_3073);
and U3372 (N_3372,N_3190,N_3174);
or U3373 (N_3373,N_3082,N_3150);
nor U3374 (N_3374,N_3115,N_3017);
nor U3375 (N_3375,N_3040,N_3089);
or U3376 (N_3376,N_3088,N_3137);
or U3377 (N_3377,N_3104,N_3174);
nand U3378 (N_3378,N_3113,N_3120);
nor U3379 (N_3379,N_3084,N_3104);
xnor U3380 (N_3380,N_3014,N_3086);
xnor U3381 (N_3381,N_3025,N_3191);
nand U3382 (N_3382,N_3119,N_3147);
or U3383 (N_3383,N_3008,N_3074);
nor U3384 (N_3384,N_3077,N_3033);
or U3385 (N_3385,N_3023,N_3049);
xnor U3386 (N_3386,N_3025,N_3189);
xnor U3387 (N_3387,N_3126,N_3025);
xnor U3388 (N_3388,N_3096,N_3142);
nand U3389 (N_3389,N_3010,N_3178);
or U3390 (N_3390,N_3149,N_3182);
or U3391 (N_3391,N_3016,N_3174);
or U3392 (N_3392,N_3160,N_3115);
nor U3393 (N_3393,N_3038,N_3198);
and U3394 (N_3394,N_3127,N_3145);
or U3395 (N_3395,N_3154,N_3022);
or U3396 (N_3396,N_3119,N_3042);
nand U3397 (N_3397,N_3151,N_3077);
and U3398 (N_3398,N_3109,N_3071);
nand U3399 (N_3399,N_3026,N_3158);
nand U3400 (N_3400,N_3343,N_3338);
nand U3401 (N_3401,N_3298,N_3375);
nand U3402 (N_3402,N_3267,N_3384);
xor U3403 (N_3403,N_3236,N_3296);
or U3404 (N_3404,N_3370,N_3399);
and U3405 (N_3405,N_3253,N_3320);
and U3406 (N_3406,N_3348,N_3259);
nor U3407 (N_3407,N_3265,N_3380);
nand U3408 (N_3408,N_3212,N_3349);
and U3409 (N_3409,N_3252,N_3364);
nand U3410 (N_3410,N_3302,N_3392);
nand U3411 (N_3411,N_3240,N_3334);
and U3412 (N_3412,N_3255,N_3374);
or U3413 (N_3413,N_3365,N_3331);
and U3414 (N_3414,N_3368,N_3237);
and U3415 (N_3415,N_3280,N_3247);
xor U3416 (N_3416,N_3225,N_3321);
and U3417 (N_3417,N_3394,N_3272);
and U3418 (N_3418,N_3254,N_3397);
nand U3419 (N_3419,N_3391,N_3290);
or U3420 (N_3420,N_3309,N_3224);
xor U3421 (N_3421,N_3233,N_3200);
and U3422 (N_3422,N_3382,N_3221);
xor U3423 (N_3423,N_3330,N_3390);
nand U3424 (N_3424,N_3208,N_3281);
xor U3425 (N_3425,N_3304,N_3317);
and U3426 (N_3426,N_3250,N_3377);
nand U3427 (N_3427,N_3319,N_3305);
xnor U3428 (N_3428,N_3363,N_3273);
xor U3429 (N_3429,N_3307,N_3354);
xnor U3430 (N_3430,N_3369,N_3387);
nand U3431 (N_3431,N_3228,N_3249);
xor U3432 (N_3432,N_3270,N_3258);
nor U3433 (N_3433,N_3293,N_3206);
and U3434 (N_3434,N_3203,N_3341);
nand U3435 (N_3435,N_3395,N_3220);
nand U3436 (N_3436,N_3332,N_3367);
nor U3437 (N_3437,N_3314,N_3300);
nor U3438 (N_3438,N_3299,N_3371);
xnor U3439 (N_3439,N_3276,N_3231);
nor U3440 (N_3440,N_3386,N_3342);
or U3441 (N_3441,N_3323,N_3204);
or U3442 (N_3442,N_3336,N_3283);
and U3443 (N_3443,N_3269,N_3398);
or U3444 (N_3444,N_3337,N_3216);
nand U3445 (N_3445,N_3211,N_3285);
xnor U3446 (N_3446,N_3286,N_3308);
nor U3447 (N_3447,N_3227,N_3361);
or U3448 (N_3448,N_3243,N_3388);
and U3449 (N_3449,N_3260,N_3262);
nand U3450 (N_3450,N_3318,N_3263);
or U3451 (N_3451,N_3282,N_3297);
nor U3452 (N_3452,N_3385,N_3213);
nand U3453 (N_3453,N_3215,N_3292);
nor U3454 (N_3454,N_3324,N_3275);
and U3455 (N_3455,N_3289,N_3376);
and U3456 (N_3456,N_3316,N_3222);
nand U3457 (N_3457,N_3242,N_3329);
nand U3458 (N_3458,N_3335,N_3294);
xnor U3459 (N_3459,N_3383,N_3295);
nand U3460 (N_3460,N_3372,N_3381);
xnor U3461 (N_3461,N_3312,N_3353);
xor U3462 (N_3462,N_3346,N_3347);
and U3463 (N_3463,N_3340,N_3345);
nand U3464 (N_3464,N_3244,N_3248);
nand U3465 (N_3465,N_3378,N_3325);
nand U3466 (N_3466,N_3328,N_3358);
and U3467 (N_3467,N_3210,N_3360);
nor U3468 (N_3468,N_3226,N_3322);
nor U3469 (N_3469,N_3251,N_3207);
nor U3470 (N_3470,N_3355,N_3327);
xor U3471 (N_3471,N_3303,N_3396);
and U3472 (N_3472,N_3389,N_3271);
or U3473 (N_3473,N_3218,N_3239);
nand U3474 (N_3474,N_3326,N_3266);
and U3475 (N_3475,N_3274,N_3278);
nor U3476 (N_3476,N_3201,N_3356);
nand U3477 (N_3477,N_3202,N_3279);
nor U3478 (N_3478,N_3234,N_3223);
nand U3479 (N_3479,N_3287,N_3351);
nor U3480 (N_3480,N_3291,N_3238);
and U3481 (N_3481,N_3288,N_3229);
xnor U3482 (N_3482,N_3393,N_3339);
and U3483 (N_3483,N_3209,N_3357);
and U3484 (N_3484,N_3352,N_3235);
nand U3485 (N_3485,N_3313,N_3362);
and U3486 (N_3486,N_3217,N_3344);
nor U3487 (N_3487,N_3214,N_3315);
or U3488 (N_3488,N_3261,N_3257);
nor U3489 (N_3489,N_3350,N_3306);
and U3490 (N_3490,N_3256,N_3232);
or U3491 (N_3491,N_3301,N_3311);
xnor U3492 (N_3492,N_3277,N_3359);
or U3493 (N_3493,N_3205,N_3245);
nand U3494 (N_3494,N_3230,N_3284);
xnor U3495 (N_3495,N_3264,N_3219);
xnor U3496 (N_3496,N_3379,N_3268);
xor U3497 (N_3497,N_3366,N_3373);
or U3498 (N_3498,N_3246,N_3241);
nand U3499 (N_3499,N_3310,N_3333);
nor U3500 (N_3500,N_3375,N_3367);
and U3501 (N_3501,N_3396,N_3353);
xor U3502 (N_3502,N_3317,N_3203);
xnor U3503 (N_3503,N_3296,N_3373);
and U3504 (N_3504,N_3205,N_3223);
or U3505 (N_3505,N_3389,N_3337);
or U3506 (N_3506,N_3254,N_3290);
nor U3507 (N_3507,N_3396,N_3376);
nor U3508 (N_3508,N_3246,N_3373);
xor U3509 (N_3509,N_3375,N_3335);
nor U3510 (N_3510,N_3289,N_3385);
nand U3511 (N_3511,N_3280,N_3316);
nand U3512 (N_3512,N_3289,N_3340);
xor U3513 (N_3513,N_3276,N_3380);
or U3514 (N_3514,N_3247,N_3329);
or U3515 (N_3515,N_3215,N_3226);
or U3516 (N_3516,N_3344,N_3362);
xor U3517 (N_3517,N_3222,N_3257);
nor U3518 (N_3518,N_3277,N_3311);
nor U3519 (N_3519,N_3236,N_3374);
xor U3520 (N_3520,N_3200,N_3324);
or U3521 (N_3521,N_3310,N_3336);
and U3522 (N_3522,N_3210,N_3272);
nand U3523 (N_3523,N_3354,N_3235);
nand U3524 (N_3524,N_3387,N_3258);
xor U3525 (N_3525,N_3398,N_3359);
nand U3526 (N_3526,N_3216,N_3228);
xor U3527 (N_3527,N_3243,N_3396);
and U3528 (N_3528,N_3275,N_3302);
xnor U3529 (N_3529,N_3211,N_3359);
nand U3530 (N_3530,N_3285,N_3230);
nor U3531 (N_3531,N_3250,N_3230);
or U3532 (N_3532,N_3217,N_3249);
and U3533 (N_3533,N_3350,N_3318);
nand U3534 (N_3534,N_3211,N_3245);
and U3535 (N_3535,N_3268,N_3341);
or U3536 (N_3536,N_3259,N_3285);
xor U3537 (N_3537,N_3203,N_3342);
xor U3538 (N_3538,N_3291,N_3258);
nand U3539 (N_3539,N_3254,N_3387);
and U3540 (N_3540,N_3395,N_3206);
and U3541 (N_3541,N_3230,N_3346);
or U3542 (N_3542,N_3284,N_3254);
nor U3543 (N_3543,N_3269,N_3291);
and U3544 (N_3544,N_3206,N_3235);
and U3545 (N_3545,N_3242,N_3234);
or U3546 (N_3546,N_3339,N_3277);
xor U3547 (N_3547,N_3308,N_3331);
or U3548 (N_3548,N_3308,N_3200);
xor U3549 (N_3549,N_3325,N_3360);
nor U3550 (N_3550,N_3348,N_3275);
nand U3551 (N_3551,N_3260,N_3355);
xor U3552 (N_3552,N_3313,N_3220);
and U3553 (N_3553,N_3390,N_3206);
xnor U3554 (N_3554,N_3394,N_3312);
or U3555 (N_3555,N_3295,N_3240);
nor U3556 (N_3556,N_3277,N_3237);
xor U3557 (N_3557,N_3215,N_3240);
nand U3558 (N_3558,N_3384,N_3221);
nor U3559 (N_3559,N_3278,N_3347);
and U3560 (N_3560,N_3212,N_3248);
nor U3561 (N_3561,N_3255,N_3206);
and U3562 (N_3562,N_3344,N_3213);
and U3563 (N_3563,N_3247,N_3372);
xor U3564 (N_3564,N_3214,N_3342);
nor U3565 (N_3565,N_3223,N_3208);
or U3566 (N_3566,N_3260,N_3331);
nor U3567 (N_3567,N_3218,N_3396);
nor U3568 (N_3568,N_3393,N_3371);
or U3569 (N_3569,N_3350,N_3241);
and U3570 (N_3570,N_3324,N_3316);
nand U3571 (N_3571,N_3387,N_3352);
or U3572 (N_3572,N_3398,N_3303);
or U3573 (N_3573,N_3343,N_3228);
and U3574 (N_3574,N_3291,N_3263);
or U3575 (N_3575,N_3283,N_3264);
and U3576 (N_3576,N_3347,N_3314);
nor U3577 (N_3577,N_3309,N_3239);
or U3578 (N_3578,N_3286,N_3293);
nor U3579 (N_3579,N_3326,N_3366);
nand U3580 (N_3580,N_3302,N_3339);
xor U3581 (N_3581,N_3257,N_3329);
or U3582 (N_3582,N_3229,N_3262);
nand U3583 (N_3583,N_3361,N_3375);
xor U3584 (N_3584,N_3352,N_3295);
xor U3585 (N_3585,N_3380,N_3362);
xnor U3586 (N_3586,N_3319,N_3294);
xor U3587 (N_3587,N_3211,N_3393);
nand U3588 (N_3588,N_3349,N_3354);
or U3589 (N_3589,N_3380,N_3352);
nand U3590 (N_3590,N_3367,N_3296);
and U3591 (N_3591,N_3352,N_3336);
and U3592 (N_3592,N_3295,N_3213);
and U3593 (N_3593,N_3386,N_3216);
or U3594 (N_3594,N_3399,N_3277);
or U3595 (N_3595,N_3373,N_3234);
or U3596 (N_3596,N_3359,N_3268);
or U3597 (N_3597,N_3340,N_3300);
nor U3598 (N_3598,N_3373,N_3342);
or U3599 (N_3599,N_3258,N_3360);
xor U3600 (N_3600,N_3458,N_3497);
nand U3601 (N_3601,N_3435,N_3569);
nand U3602 (N_3602,N_3496,N_3570);
and U3603 (N_3603,N_3445,N_3457);
and U3604 (N_3604,N_3577,N_3464);
or U3605 (N_3605,N_3410,N_3551);
nand U3606 (N_3606,N_3425,N_3519);
nand U3607 (N_3607,N_3557,N_3532);
or U3608 (N_3608,N_3523,N_3545);
and U3609 (N_3609,N_3586,N_3503);
xor U3610 (N_3610,N_3494,N_3585);
nor U3611 (N_3611,N_3488,N_3543);
and U3612 (N_3612,N_3486,N_3429);
nand U3613 (N_3613,N_3453,N_3472);
or U3614 (N_3614,N_3546,N_3579);
or U3615 (N_3615,N_3414,N_3454);
and U3616 (N_3616,N_3555,N_3487);
nand U3617 (N_3617,N_3516,N_3491);
nor U3618 (N_3618,N_3599,N_3483);
nor U3619 (N_3619,N_3449,N_3447);
nand U3620 (N_3620,N_3561,N_3473);
or U3621 (N_3621,N_3430,N_3404);
and U3622 (N_3622,N_3448,N_3530);
xor U3623 (N_3623,N_3506,N_3493);
xor U3624 (N_3624,N_3580,N_3427);
nand U3625 (N_3625,N_3535,N_3542);
and U3626 (N_3626,N_3584,N_3596);
nand U3627 (N_3627,N_3463,N_3411);
nor U3628 (N_3628,N_3508,N_3574);
and U3629 (N_3629,N_3556,N_3538);
and U3630 (N_3630,N_3597,N_3451);
xnor U3631 (N_3631,N_3564,N_3568);
nand U3632 (N_3632,N_3499,N_3573);
and U3633 (N_3633,N_3548,N_3438);
xor U3634 (N_3634,N_3423,N_3459);
nor U3635 (N_3635,N_3510,N_3527);
nand U3636 (N_3636,N_3419,N_3431);
and U3637 (N_3637,N_3460,N_3504);
xnor U3638 (N_3638,N_3592,N_3441);
or U3639 (N_3639,N_3469,N_3582);
or U3640 (N_3640,N_3501,N_3528);
or U3641 (N_3641,N_3518,N_3541);
xnor U3642 (N_3642,N_3439,N_3511);
nor U3643 (N_3643,N_3442,N_3540);
nor U3644 (N_3644,N_3547,N_3426);
or U3645 (N_3645,N_3558,N_3544);
nand U3646 (N_3646,N_3515,N_3509);
or U3647 (N_3647,N_3594,N_3481);
nand U3648 (N_3648,N_3524,N_3461);
nor U3649 (N_3649,N_3467,N_3480);
nor U3650 (N_3650,N_3406,N_3575);
and U3651 (N_3651,N_3578,N_3581);
nor U3652 (N_3652,N_3420,N_3479);
xor U3653 (N_3653,N_3571,N_3462);
xnor U3654 (N_3654,N_3492,N_3450);
or U3655 (N_3655,N_3514,N_3475);
or U3656 (N_3656,N_3466,N_3428);
and U3657 (N_3657,N_3500,N_3553);
nor U3658 (N_3658,N_3520,N_3489);
nor U3659 (N_3659,N_3440,N_3560);
xor U3660 (N_3660,N_3407,N_3482);
or U3661 (N_3661,N_3405,N_3531);
xor U3662 (N_3662,N_3495,N_3408);
or U3663 (N_3663,N_3583,N_3416);
and U3664 (N_3664,N_3550,N_3456);
or U3665 (N_3665,N_3563,N_3415);
and U3666 (N_3666,N_3598,N_3572);
nand U3667 (N_3667,N_3477,N_3517);
xor U3668 (N_3668,N_3562,N_3554);
nand U3669 (N_3669,N_3507,N_3436);
or U3670 (N_3670,N_3455,N_3513);
nor U3671 (N_3671,N_3422,N_3444);
xor U3672 (N_3672,N_3476,N_3537);
or U3673 (N_3673,N_3433,N_3589);
or U3674 (N_3674,N_3446,N_3403);
xnor U3675 (N_3675,N_3409,N_3521);
and U3676 (N_3676,N_3402,N_3529);
nand U3677 (N_3677,N_3595,N_3502);
or U3678 (N_3678,N_3443,N_3418);
xnor U3679 (N_3679,N_3490,N_3432);
nand U3680 (N_3680,N_3434,N_3452);
and U3681 (N_3681,N_3485,N_3401);
or U3682 (N_3682,N_3424,N_3421);
or U3683 (N_3683,N_3471,N_3522);
nor U3684 (N_3684,N_3549,N_3512);
and U3685 (N_3685,N_3565,N_3474);
or U3686 (N_3686,N_3470,N_3400);
xnor U3687 (N_3687,N_3526,N_3536);
and U3688 (N_3688,N_3525,N_3534);
nand U3689 (N_3689,N_3539,N_3593);
nand U3690 (N_3690,N_3588,N_3566);
and U3691 (N_3691,N_3590,N_3567);
nor U3692 (N_3692,N_3412,N_3591);
nor U3693 (N_3693,N_3484,N_3559);
and U3694 (N_3694,N_3437,N_3478);
or U3695 (N_3695,N_3465,N_3533);
nand U3696 (N_3696,N_3417,N_3576);
nand U3697 (N_3697,N_3552,N_3413);
or U3698 (N_3698,N_3468,N_3587);
xnor U3699 (N_3699,N_3498,N_3505);
or U3700 (N_3700,N_3472,N_3569);
and U3701 (N_3701,N_3425,N_3484);
nor U3702 (N_3702,N_3489,N_3479);
nor U3703 (N_3703,N_3512,N_3480);
or U3704 (N_3704,N_3407,N_3450);
and U3705 (N_3705,N_3465,N_3583);
or U3706 (N_3706,N_3546,N_3437);
and U3707 (N_3707,N_3538,N_3420);
and U3708 (N_3708,N_3508,N_3547);
or U3709 (N_3709,N_3500,N_3501);
nand U3710 (N_3710,N_3445,N_3464);
xnor U3711 (N_3711,N_3411,N_3414);
nor U3712 (N_3712,N_3412,N_3573);
nand U3713 (N_3713,N_3522,N_3538);
xor U3714 (N_3714,N_3424,N_3439);
nand U3715 (N_3715,N_3526,N_3437);
xor U3716 (N_3716,N_3452,N_3498);
nor U3717 (N_3717,N_3571,N_3565);
or U3718 (N_3718,N_3438,N_3485);
xor U3719 (N_3719,N_3509,N_3574);
xor U3720 (N_3720,N_3418,N_3455);
xor U3721 (N_3721,N_3495,N_3567);
nand U3722 (N_3722,N_3554,N_3527);
nor U3723 (N_3723,N_3463,N_3465);
nand U3724 (N_3724,N_3580,N_3495);
or U3725 (N_3725,N_3570,N_3482);
and U3726 (N_3726,N_3414,N_3593);
or U3727 (N_3727,N_3518,N_3463);
xor U3728 (N_3728,N_3512,N_3474);
and U3729 (N_3729,N_3421,N_3587);
nor U3730 (N_3730,N_3485,N_3578);
nand U3731 (N_3731,N_3418,N_3436);
or U3732 (N_3732,N_3534,N_3488);
xnor U3733 (N_3733,N_3567,N_3458);
nor U3734 (N_3734,N_3492,N_3556);
xnor U3735 (N_3735,N_3448,N_3465);
nand U3736 (N_3736,N_3476,N_3406);
nand U3737 (N_3737,N_3531,N_3503);
or U3738 (N_3738,N_3412,N_3442);
or U3739 (N_3739,N_3493,N_3452);
xnor U3740 (N_3740,N_3487,N_3413);
and U3741 (N_3741,N_3496,N_3468);
or U3742 (N_3742,N_3563,N_3568);
xor U3743 (N_3743,N_3498,N_3507);
xnor U3744 (N_3744,N_3551,N_3515);
or U3745 (N_3745,N_3425,N_3555);
and U3746 (N_3746,N_3425,N_3485);
nand U3747 (N_3747,N_3407,N_3578);
xor U3748 (N_3748,N_3479,N_3417);
or U3749 (N_3749,N_3500,N_3416);
nand U3750 (N_3750,N_3469,N_3423);
and U3751 (N_3751,N_3500,N_3496);
nand U3752 (N_3752,N_3481,N_3512);
xor U3753 (N_3753,N_3557,N_3468);
or U3754 (N_3754,N_3595,N_3559);
xnor U3755 (N_3755,N_3565,N_3456);
nand U3756 (N_3756,N_3441,N_3447);
xor U3757 (N_3757,N_3586,N_3595);
nand U3758 (N_3758,N_3573,N_3572);
nor U3759 (N_3759,N_3440,N_3439);
or U3760 (N_3760,N_3539,N_3521);
and U3761 (N_3761,N_3450,N_3453);
and U3762 (N_3762,N_3435,N_3502);
nor U3763 (N_3763,N_3472,N_3484);
nor U3764 (N_3764,N_3577,N_3485);
xnor U3765 (N_3765,N_3495,N_3477);
or U3766 (N_3766,N_3408,N_3528);
xnor U3767 (N_3767,N_3469,N_3435);
nor U3768 (N_3768,N_3549,N_3557);
or U3769 (N_3769,N_3407,N_3543);
nand U3770 (N_3770,N_3486,N_3488);
and U3771 (N_3771,N_3513,N_3568);
xor U3772 (N_3772,N_3462,N_3524);
or U3773 (N_3773,N_3445,N_3585);
or U3774 (N_3774,N_3401,N_3507);
and U3775 (N_3775,N_3567,N_3528);
nor U3776 (N_3776,N_3537,N_3454);
nand U3777 (N_3777,N_3579,N_3444);
nor U3778 (N_3778,N_3436,N_3569);
xor U3779 (N_3779,N_3598,N_3463);
and U3780 (N_3780,N_3568,N_3473);
and U3781 (N_3781,N_3462,N_3527);
nand U3782 (N_3782,N_3465,N_3510);
xnor U3783 (N_3783,N_3472,N_3574);
or U3784 (N_3784,N_3494,N_3459);
and U3785 (N_3785,N_3535,N_3599);
nor U3786 (N_3786,N_3497,N_3558);
nor U3787 (N_3787,N_3596,N_3495);
xnor U3788 (N_3788,N_3443,N_3469);
xor U3789 (N_3789,N_3541,N_3547);
xor U3790 (N_3790,N_3407,N_3441);
xor U3791 (N_3791,N_3430,N_3580);
or U3792 (N_3792,N_3589,N_3492);
nand U3793 (N_3793,N_3453,N_3433);
and U3794 (N_3794,N_3459,N_3475);
and U3795 (N_3795,N_3569,N_3504);
and U3796 (N_3796,N_3555,N_3556);
xnor U3797 (N_3797,N_3462,N_3400);
xnor U3798 (N_3798,N_3449,N_3517);
nand U3799 (N_3799,N_3429,N_3500);
nand U3800 (N_3800,N_3796,N_3656);
xor U3801 (N_3801,N_3610,N_3682);
and U3802 (N_3802,N_3670,N_3630);
xnor U3803 (N_3803,N_3750,N_3709);
or U3804 (N_3804,N_3737,N_3754);
xnor U3805 (N_3805,N_3713,N_3600);
nor U3806 (N_3806,N_3767,N_3793);
nor U3807 (N_3807,N_3690,N_3757);
xnor U3808 (N_3808,N_3685,N_3627);
and U3809 (N_3809,N_3786,N_3747);
or U3810 (N_3810,N_3671,N_3677);
nand U3811 (N_3811,N_3738,N_3647);
xnor U3812 (N_3812,N_3740,N_3790);
nor U3813 (N_3813,N_3604,N_3650);
nor U3814 (N_3814,N_3691,N_3640);
nor U3815 (N_3815,N_3621,N_3632);
xnor U3816 (N_3816,N_3628,N_3624);
nor U3817 (N_3817,N_3755,N_3783);
nand U3818 (N_3818,N_3602,N_3605);
and U3819 (N_3819,N_3657,N_3689);
or U3820 (N_3820,N_3639,N_3648);
nand U3821 (N_3821,N_3743,N_3629);
or U3822 (N_3822,N_3751,N_3649);
nand U3823 (N_3823,N_3718,N_3787);
nor U3824 (N_3824,N_3728,N_3601);
nor U3825 (N_3825,N_3616,N_3715);
nor U3826 (N_3826,N_3724,N_3712);
nand U3827 (N_3827,N_3635,N_3717);
xor U3828 (N_3828,N_3725,N_3700);
or U3829 (N_3829,N_3739,N_3703);
nand U3830 (N_3830,N_3668,N_3766);
nand U3831 (N_3831,N_3694,N_3683);
and U3832 (N_3832,N_3731,N_3723);
xnor U3833 (N_3833,N_3768,N_3654);
nand U3834 (N_3834,N_3704,N_3662);
nor U3835 (N_3835,N_3660,N_3637);
nand U3836 (N_3836,N_3765,N_3698);
or U3837 (N_3837,N_3669,N_3675);
or U3838 (N_3838,N_3772,N_3607);
xnor U3839 (N_3839,N_3617,N_3777);
xor U3840 (N_3840,N_3779,N_3618);
nor U3841 (N_3841,N_3612,N_3642);
nand U3842 (N_3842,N_3705,N_3778);
nand U3843 (N_3843,N_3692,N_3614);
xor U3844 (N_3844,N_3638,N_3644);
nand U3845 (N_3845,N_3730,N_3633);
nor U3846 (N_3846,N_3702,N_3696);
xor U3847 (N_3847,N_3665,N_3761);
xnor U3848 (N_3848,N_3716,N_3780);
and U3849 (N_3849,N_3746,N_3655);
nand U3850 (N_3850,N_3646,N_3661);
nor U3851 (N_3851,N_3726,N_3678);
or U3852 (N_3852,N_3613,N_3736);
and U3853 (N_3853,N_3688,N_3720);
or U3854 (N_3854,N_3667,N_3734);
or U3855 (N_3855,N_3773,N_3606);
nor U3856 (N_3856,N_3697,N_3721);
xor U3857 (N_3857,N_3745,N_3785);
and U3858 (N_3858,N_3684,N_3770);
nor U3859 (N_3859,N_3760,N_3615);
nand U3860 (N_3860,N_3681,N_3753);
nand U3861 (N_3861,N_3792,N_3699);
nor U3862 (N_3862,N_3774,N_3788);
nand U3863 (N_3863,N_3622,N_3664);
nor U3864 (N_3864,N_3722,N_3749);
and U3865 (N_3865,N_3626,N_3714);
xor U3866 (N_3866,N_3625,N_3789);
nand U3867 (N_3867,N_3659,N_3676);
nor U3868 (N_3868,N_3641,N_3769);
and U3869 (N_3869,N_3758,N_3651);
xor U3870 (N_3870,N_3762,N_3794);
xnor U3871 (N_3871,N_3708,N_3666);
nor U3872 (N_3872,N_3631,N_3686);
nand U3873 (N_3873,N_3775,N_3735);
nand U3874 (N_3874,N_3742,N_3680);
nand U3875 (N_3875,N_3727,N_3782);
nor U3876 (N_3876,N_3764,N_3781);
and U3877 (N_3877,N_3784,N_3791);
and U3878 (N_3878,N_3609,N_3658);
nor U3879 (N_3879,N_3759,N_3672);
nand U3880 (N_3880,N_3763,N_3673);
or U3881 (N_3881,N_3797,N_3643);
xor U3882 (N_3882,N_3674,N_3620);
nand U3883 (N_3883,N_3798,N_3776);
nand U3884 (N_3884,N_3795,N_3756);
nand U3885 (N_3885,N_3711,N_3706);
or U3886 (N_3886,N_3663,N_3653);
xnor U3887 (N_3887,N_3771,N_3799);
nand U3888 (N_3888,N_3733,N_3693);
nand U3889 (N_3889,N_3611,N_3701);
nand U3890 (N_3890,N_3707,N_3634);
or U3891 (N_3891,N_3748,N_3623);
xor U3892 (N_3892,N_3710,N_3687);
and U3893 (N_3893,N_3603,N_3636);
and U3894 (N_3894,N_3619,N_3645);
nor U3895 (N_3895,N_3652,N_3744);
or U3896 (N_3896,N_3679,N_3752);
xnor U3897 (N_3897,N_3719,N_3608);
and U3898 (N_3898,N_3732,N_3695);
or U3899 (N_3899,N_3741,N_3729);
nand U3900 (N_3900,N_3618,N_3770);
xnor U3901 (N_3901,N_3716,N_3603);
nor U3902 (N_3902,N_3733,N_3750);
nand U3903 (N_3903,N_3645,N_3793);
nand U3904 (N_3904,N_3724,N_3658);
nand U3905 (N_3905,N_3673,N_3728);
nand U3906 (N_3906,N_3773,N_3793);
and U3907 (N_3907,N_3718,N_3625);
nand U3908 (N_3908,N_3636,N_3673);
nor U3909 (N_3909,N_3720,N_3695);
or U3910 (N_3910,N_3694,N_3743);
nor U3911 (N_3911,N_3667,N_3636);
nand U3912 (N_3912,N_3703,N_3673);
nand U3913 (N_3913,N_3605,N_3796);
or U3914 (N_3914,N_3780,N_3751);
xor U3915 (N_3915,N_3616,N_3790);
and U3916 (N_3916,N_3711,N_3798);
and U3917 (N_3917,N_3653,N_3778);
nand U3918 (N_3918,N_3611,N_3685);
or U3919 (N_3919,N_3691,N_3754);
nand U3920 (N_3920,N_3655,N_3636);
and U3921 (N_3921,N_3644,N_3721);
xor U3922 (N_3922,N_3755,N_3797);
or U3923 (N_3923,N_3626,N_3610);
xor U3924 (N_3924,N_3642,N_3671);
or U3925 (N_3925,N_3621,N_3792);
and U3926 (N_3926,N_3717,N_3689);
xor U3927 (N_3927,N_3677,N_3689);
nand U3928 (N_3928,N_3789,N_3749);
nor U3929 (N_3929,N_3737,N_3735);
nand U3930 (N_3930,N_3792,N_3601);
or U3931 (N_3931,N_3686,N_3601);
and U3932 (N_3932,N_3757,N_3760);
nand U3933 (N_3933,N_3756,N_3669);
xor U3934 (N_3934,N_3614,N_3706);
nand U3935 (N_3935,N_3759,N_3750);
xor U3936 (N_3936,N_3763,N_3601);
and U3937 (N_3937,N_3717,N_3779);
or U3938 (N_3938,N_3632,N_3799);
or U3939 (N_3939,N_3766,N_3672);
nor U3940 (N_3940,N_3600,N_3654);
nand U3941 (N_3941,N_3777,N_3655);
nand U3942 (N_3942,N_3633,N_3733);
and U3943 (N_3943,N_3678,N_3634);
xnor U3944 (N_3944,N_3679,N_3709);
xnor U3945 (N_3945,N_3603,N_3660);
nand U3946 (N_3946,N_3681,N_3704);
nand U3947 (N_3947,N_3799,N_3631);
nor U3948 (N_3948,N_3620,N_3677);
nand U3949 (N_3949,N_3709,N_3632);
or U3950 (N_3950,N_3612,N_3737);
and U3951 (N_3951,N_3662,N_3700);
and U3952 (N_3952,N_3619,N_3780);
nor U3953 (N_3953,N_3738,N_3798);
nor U3954 (N_3954,N_3639,N_3756);
nand U3955 (N_3955,N_3786,N_3797);
and U3956 (N_3956,N_3640,N_3683);
nor U3957 (N_3957,N_3689,N_3675);
nand U3958 (N_3958,N_3720,N_3714);
or U3959 (N_3959,N_3637,N_3738);
or U3960 (N_3960,N_3620,N_3612);
nor U3961 (N_3961,N_3751,N_3636);
or U3962 (N_3962,N_3710,N_3780);
xor U3963 (N_3963,N_3706,N_3612);
nand U3964 (N_3964,N_3643,N_3682);
xor U3965 (N_3965,N_3756,N_3658);
xor U3966 (N_3966,N_3641,N_3730);
or U3967 (N_3967,N_3610,N_3671);
or U3968 (N_3968,N_3640,N_3607);
nand U3969 (N_3969,N_3702,N_3716);
and U3970 (N_3970,N_3733,N_3771);
xor U3971 (N_3971,N_3742,N_3789);
xor U3972 (N_3972,N_3627,N_3638);
or U3973 (N_3973,N_3763,N_3742);
and U3974 (N_3974,N_3675,N_3756);
nor U3975 (N_3975,N_3692,N_3605);
nor U3976 (N_3976,N_3628,N_3689);
nor U3977 (N_3977,N_3738,N_3795);
nand U3978 (N_3978,N_3606,N_3669);
nand U3979 (N_3979,N_3628,N_3616);
nand U3980 (N_3980,N_3796,N_3664);
and U3981 (N_3981,N_3746,N_3672);
nand U3982 (N_3982,N_3682,N_3750);
and U3983 (N_3983,N_3637,N_3723);
xnor U3984 (N_3984,N_3756,N_3742);
and U3985 (N_3985,N_3721,N_3655);
and U3986 (N_3986,N_3795,N_3629);
and U3987 (N_3987,N_3740,N_3681);
and U3988 (N_3988,N_3652,N_3726);
nor U3989 (N_3989,N_3662,N_3600);
nand U3990 (N_3990,N_3781,N_3686);
xnor U3991 (N_3991,N_3677,N_3663);
xor U3992 (N_3992,N_3662,N_3661);
or U3993 (N_3993,N_3639,N_3792);
xnor U3994 (N_3994,N_3722,N_3799);
nor U3995 (N_3995,N_3769,N_3669);
xor U3996 (N_3996,N_3777,N_3761);
and U3997 (N_3997,N_3758,N_3603);
or U3998 (N_3998,N_3634,N_3735);
and U3999 (N_3999,N_3718,N_3626);
xor U4000 (N_4000,N_3965,N_3951);
nand U4001 (N_4001,N_3801,N_3881);
or U4002 (N_4002,N_3889,N_3960);
xnor U4003 (N_4003,N_3824,N_3908);
nand U4004 (N_4004,N_3933,N_3875);
or U4005 (N_4005,N_3934,N_3911);
nand U4006 (N_4006,N_3978,N_3859);
and U4007 (N_4007,N_3809,N_3868);
and U4008 (N_4008,N_3973,N_3822);
xor U4009 (N_4009,N_3854,N_3969);
nand U4010 (N_4010,N_3986,N_3953);
nor U4011 (N_4011,N_3983,N_3853);
xnor U4012 (N_4012,N_3925,N_3929);
and U4013 (N_4013,N_3846,N_3865);
xor U4014 (N_4014,N_3860,N_3998);
nor U4015 (N_4015,N_3936,N_3807);
nand U4016 (N_4016,N_3917,N_3818);
and U4017 (N_4017,N_3898,N_3841);
or U4018 (N_4018,N_3836,N_3872);
nor U4019 (N_4019,N_3930,N_3894);
nor U4020 (N_4020,N_3977,N_3959);
and U4021 (N_4021,N_3989,N_3949);
or U4022 (N_4022,N_3913,N_3842);
and U4023 (N_4023,N_3849,N_3827);
nand U4024 (N_4024,N_3931,N_3902);
xor U4025 (N_4025,N_3855,N_3935);
xnor U4026 (N_4026,N_3851,N_3915);
and U4027 (N_4027,N_3961,N_3800);
nand U4028 (N_4028,N_3834,N_3967);
nand U4029 (N_4029,N_3999,N_3987);
nand U4030 (N_4030,N_3957,N_3912);
nand U4031 (N_4031,N_3985,N_3924);
or U4032 (N_4032,N_3907,N_3815);
xnor U4033 (N_4033,N_3821,N_3992);
nand U4034 (N_4034,N_3848,N_3877);
nor U4035 (N_4035,N_3988,N_3937);
nor U4036 (N_4036,N_3995,N_3997);
and U4037 (N_4037,N_3927,N_3814);
nor U4038 (N_4038,N_3845,N_3941);
nor U4039 (N_4039,N_3910,N_3825);
or U4040 (N_4040,N_3950,N_3900);
nor U4041 (N_4041,N_3954,N_3944);
nor U4042 (N_4042,N_3904,N_3883);
nand U4043 (N_4043,N_3873,N_3952);
or U4044 (N_4044,N_3896,N_3867);
xor U4045 (N_4045,N_3939,N_3837);
or U4046 (N_4046,N_3990,N_3823);
and U4047 (N_4047,N_3886,N_3878);
or U4048 (N_4048,N_3938,N_3905);
nand U4049 (N_4049,N_3962,N_3948);
xor U4050 (N_4050,N_3892,N_3832);
or U4051 (N_4051,N_3893,N_3861);
nor U4052 (N_4052,N_3901,N_3979);
or U4053 (N_4053,N_3811,N_3890);
or U4054 (N_4054,N_3947,N_3819);
or U4055 (N_4055,N_3816,N_3850);
nand U4056 (N_4056,N_3866,N_3820);
nor U4057 (N_4057,N_3870,N_3888);
and U4058 (N_4058,N_3928,N_3970);
nand U4059 (N_4059,N_3817,N_3926);
or U4060 (N_4060,N_3826,N_3980);
nand U4061 (N_4061,N_3812,N_3974);
nand U4062 (N_4062,N_3810,N_3991);
xor U4063 (N_4063,N_3981,N_3887);
nor U4064 (N_4064,N_3879,N_3876);
and U4065 (N_4065,N_3895,N_3920);
or U4066 (N_4066,N_3963,N_3994);
nor U4067 (N_4067,N_3828,N_3996);
nand U4068 (N_4068,N_3806,N_3964);
nand U4069 (N_4069,N_3869,N_3943);
and U4070 (N_4070,N_3802,N_3839);
nor U4071 (N_4071,N_3899,N_3966);
xnor U4072 (N_4072,N_3813,N_3840);
and U4073 (N_4073,N_3946,N_3982);
and U4074 (N_4074,N_3847,N_3916);
nor U4075 (N_4075,N_3808,N_3830);
nor U4076 (N_4076,N_3906,N_3968);
nor U4077 (N_4077,N_3958,N_3897);
nand U4078 (N_4078,N_3831,N_3923);
xor U4079 (N_4079,N_3956,N_3844);
nand U4080 (N_4080,N_3803,N_3976);
xnor U4081 (N_4081,N_3903,N_3922);
and U4082 (N_4082,N_3843,N_3863);
nand U4083 (N_4083,N_3993,N_3805);
and U4084 (N_4084,N_3880,N_3884);
or U4085 (N_4085,N_3909,N_3857);
or U4086 (N_4086,N_3891,N_3856);
nor U4087 (N_4087,N_3829,N_3804);
xnor U4088 (N_4088,N_3835,N_3862);
and U4089 (N_4089,N_3932,N_3885);
xor U4090 (N_4090,N_3971,N_3914);
and U4091 (N_4091,N_3874,N_3919);
and U4092 (N_4092,N_3882,N_3852);
nand U4093 (N_4093,N_3838,N_3864);
nand U4094 (N_4094,N_3940,N_3833);
nand U4095 (N_4095,N_3955,N_3858);
nor U4096 (N_4096,N_3942,N_3975);
xor U4097 (N_4097,N_3984,N_3921);
nand U4098 (N_4098,N_3918,N_3945);
or U4099 (N_4099,N_3871,N_3972);
nor U4100 (N_4100,N_3967,N_3851);
nor U4101 (N_4101,N_3853,N_3931);
nor U4102 (N_4102,N_3835,N_3853);
nand U4103 (N_4103,N_3983,N_3957);
nand U4104 (N_4104,N_3894,N_3847);
or U4105 (N_4105,N_3904,N_3995);
xnor U4106 (N_4106,N_3905,N_3822);
xor U4107 (N_4107,N_3903,N_3829);
and U4108 (N_4108,N_3945,N_3968);
or U4109 (N_4109,N_3824,N_3843);
or U4110 (N_4110,N_3927,N_3987);
nor U4111 (N_4111,N_3928,N_3864);
nor U4112 (N_4112,N_3896,N_3984);
or U4113 (N_4113,N_3944,N_3899);
xnor U4114 (N_4114,N_3885,N_3959);
nor U4115 (N_4115,N_3972,N_3844);
nand U4116 (N_4116,N_3887,N_3870);
nand U4117 (N_4117,N_3968,N_3865);
and U4118 (N_4118,N_3923,N_3808);
xnor U4119 (N_4119,N_3895,N_3808);
nor U4120 (N_4120,N_3995,N_3972);
or U4121 (N_4121,N_3986,N_3838);
nand U4122 (N_4122,N_3840,N_3870);
and U4123 (N_4123,N_3913,N_3815);
nand U4124 (N_4124,N_3857,N_3901);
xor U4125 (N_4125,N_3809,N_3829);
nand U4126 (N_4126,N_3942,N_3820);
and U4127 (N_4127,N_3837,N_3908);
nand U4128 (N_4128,N_3997,N_3883);
xor U4129 (N_4129,N_3834,N_3857);
nor U4130 (N_4130,N_3889,N_3831);
xor U4131 (N_4131,N_3940,N_3992);
and U4132 (N_4132,N_3933,N_3809);
or U4133 (N_4133,N_3860,N_3922);
nand U4134 (N_4134,N_3925,N_3948);
or U4135 (N_4135,N_3973,N_3886);
nand U4136 (N_4136,N_3988,N_3883);
nor U4137 (N_4137,N_3882,N_3924);
xnor U4138 (N_4138,N_3976,N_3955);
and U4139 (N_4139,N_3897,N_3908);
nand U4140 (N_4140,N_3844,N_3906);
nand U4141 (N_4141,N_3844,N_3974);
or U4142 (N_4142,N_3880,N_3945);
or U4143 (N_4143,N_3976,N_3812);
nor U4144 (N_4144,N_3828,N_3907);
or U4145 (N_4145,N_3848,N_3940);
xor U4146 (N_4146,N_3871,N_3903);
xor U4147 (N_4147,N_3825,N_3924);
or U4148 (N_4148,N_3964,N_3952);
xor U4149 (N_4149,N_3815,N_3869);
or U4150 (N_4150,N_3882,N_3825);
nand U4151 (N_4151,N_3962,N_3869);
nand U4152 (N_4152,N_3940,N_3965);
nor U4153 (N_4153,N_3833,N_3947);
xor U4154 (N_4154,N_3976,N_3871);
nand U4155 (N_4155,N_3893,N_3840);
or U4156 (N_4156,N_3999,N_3918);
nand U4157 (N_4157,N_3895,N_3917);
nand U4158 (N_4158,N_3848,N_3800);
nand U4159 (N_4159,N_3945,N_3972);
nor U4160 (N_4160,N_3963,N_3860);
nor U4161 (N_4161,N_3828,N_3875);
xor U4162 (N_4162,N_3800,N_3913);
nand U4163 (N_4163,N_3864,N_3903);
nand U4164 (N_4164,N_3973,N_3810);
xor U4165 (N_4165,N_3911,N_3980);
and U4166 (N_4166,N_3999,N_3948);
nand U4167 (N_4167,N_3842,N_3810);
and U4168 (N_4168,N_3964,N_3975);
nor U4169 (N_4169,N_3957,N_3942);
xor U4170 (N_4170,N_3816,N_3854);
nand U4171 (N_4171,N_3861,N_3989);
nand U4172 (N_4172,N_3876,N_3945);
or U4173 (N_4173,N_3986,N_3891);
nor U4174 (N_4174,N_3846,N_3849);
and U4175 (N_4175,N_3955,N_3971);
nand U4176 (N_4176,N_3956,N_3916);
or U4177 (N_4177,N_3820,N_3835);
xnor U4178 (N_4178,N_3946,N_3999);
xnor U4179 (N_4179,N_3863,N_3821);
xor U4180 (N_4180,N_3812,N_3860);
xor U4181 (N_4181,N_3905,N_3831);
nand U4182 (N_4182,N_3987,N_3852);
nand U4183 (N_4183,N_3991,N_3802);
xor U4184 (N_4184,N_3841,N_3883);
xor U4185 (N_4185,N_3963,N_3851);
nor U4186 (N_4186,N_3820,N_3890);
nand U4187 (N_4187,N_3918,N_3964);
nand U4188 (N_4188,N_3866,N_3867);
xnor U4189 (N_4189,N_3815,N_3943);
xnor U4190 (N_4190,N_3936,N_3834);
nand U4191 (N_4191,N_3914,N_3896);
or U4192 (N_4192,N_3905,N_3878);
nor U4193 (N_4193,N_3840,N_3803);
xnor U4194 (N_4194,N_3908,N_3875);
and U4195 (N_4195,N_3901,N_3883);
nor U4196 (N_4196,N_3895,N_3991);
nand U4197 (N_4197,N_3803,N_3925);
nor U4198 (N_4198,N_3873,N_3895);
nand U4199 (N_4199,N_3990,N_3982);
nor U4200 (N_4200,N_4181,N_4086);
or U4201 (N_4201,N_4040,N_4136);
xnor U4202 (N_4202,N_4074,N_4122);
and U4203 (N_4203,N_4082,N_4045);
and U4204 (N_4204,N_4053,N_4035);
nor U4205 (N_4205,N_4002,N_4048);
nor U4206 (N_4206,N_4070,N_4016);
nand U4207 (N_4207,N_4155,N_4011);
nor U4208 (N_4208,N_4167,N_4096);
nand U4209 (N_4209,N_4064,N_4071);
and U4210 (N_4210,N_4001,N_4139);
and U4211 (N_4211,N_4063,N_4125);
nand U4212 (N_4212,N_4158,N_4196);
nand U4213 (N_4213,N_4033,N_4104);
or U4214 (N_4214,N_4147,N_4187);
or U4215 (N_4215,N_4089,N_4198);
xor U4216 (N_4216,N_4107,N_4188);
and U4217 (N_4217,N_4007,N_4084);
nand U4218 (N_4218,N_4050,N_4156);
or U4219 (N_4219,N_4020,N_4174);
nand U4220 (N_4220,N_4129,N_4140);
xnor U4221 (N_4221,N_4003,N_4058);
xor U4222 (N_4222,N_4061,N_4093);
or U4223 (N_4223,N_4010,N_4013);
xnor U4224 (N_4224,N_4005,N_4173);
nand U4225 (N_4225,N_4037,N_4166);
xor U4226 (N_4226,N_4014,N_4118);
xnor U4227 (N_4227,N_4103,N_4057);
or U4228 (N_4228,N_4132,N_4094);
and U4229 (N_4229,N_4112,N_4163);
or U4230 (N_4230,N_4062,N_4119);
and U4231 (N_4231,N_4006,N_4030);
nor U4232 (N_4232,N_4000,N_4021);
and U4233 (N_4233,N_4032,N_4012);
nand U4234 (N_4234,N_4152,N_4161);
or U4235 (N_4235,N_4175,N_4191);
nand U4236 (N_4236,N_4085,N_4179);
nand U4237 (N_4237,N_4009,N_4049);
nor U4238 (N_4238,N_4115,N_4121);
xor U4239 (N_4239,N_4076,N_4072);
nand U4240 (N_4240,N_4075,N_4060);
or U4241 (N_4241,N_4029,N_4113);
and U4242 (N_4242,N_4059,N_4176);
nor U4243 (N_4243,N_4055,N_4039);
and U4244 (N_4244,N_4168,N_4068);
or U4245 (N_4245,N_4131,N_4151);
nor U4246 (N_4246,N_4098,N_4124);
or U4247 (N_4247,N_4114,N_4034);
nor U4248 (N_4248,N_4066,N_4024);
xnor U4249 (N_4249,N_4194,N_4189);
and U4250 (N_4250,N_4195,N_4190);
nor U4251 (N_4251,N_4197,N_4022);
xor U4252 (N_4252,N_4038,N_4133);
and U4253 (N_4253,N_4182,N_4044);
nand U4254 (N_4254,N_4088,N_4144);
nand U4255 (N_4255,N_4169,N_4192);
nor U4256 (N_4256,N_4162,N_4036);
nor U4257 (N_4257,N_4123,N_4092);
and U4258 (N_4258,N_4047,N_4023);
nor U4259 (N_4259,N_4081,N_4046);
and U4260 (N_4260,N_4160,N_4141);
nor U4261 (N_4261,N_4065,N_4083);
and U4262 (N_4262,N_4165,N_4159);
nor U4263 (N_4263,N_4116,N_4134);
or U4264 (N_4264,N_4177,N_4199);
and U4265 (N_4265,N_4130,N_4157);
nand U4266 (N_4266,N_4041,N_4051);
and U4267 (N_4267,N_4079,N_4106);
and U4268 (N_4268,N_4017,N_4073);
and U4269 (N_4269,N_4031,N_4137);
or U4270 (N_4270,N_4052,N_4126);
nor U4271 (N_4271,N_4067,N_4111);
nor U4272 (N_4272,N_4100,N_4145);
and U4273 (N_4273,N_4056,N_4018);
nand U4274 (N_4274,N_4043,N_4095);
and U4275 (N_4275,N_4180,N_4091);
xor U4276 (N_4276,N_4110,N_4148);
and U4277 (N_4277,N_4120,N_4186);
xnor U4278 (N_4278,N_4008,N_4069);
xor U4279 (N_4279,N_4019,N_4109);
and U4280 (N_4280,N_4185,N_4153);
nor U4281 (N_4281,N_4117,N_4170);
or U4282 (N_4282,N_4183,N_4150);
and U4283 (N_4283,N_4078,N_4077);
or U4284 (N_4284,N_4135,N_4090);
or U4285 (N_4285,N_4127,N_4154);
nand U4286 (N_4286,N_4101,N_4138);
nor U4287 (N_4287,N_4128,N_4143);
and U4288 (N_4288,N_4028,N_4164);
xnor U4289 (N_4289,N_4054,N_4099);
nand U4290 (N_4290,N_4080,N_4097);
or U4291 (N_4291,N_4193,N_4026);
nand U4292 (N_4292,N_4172,N_4142);
and U4293 (N_4293,N_4171,N_4184);
and U4294 (N_4294,N_4178,N_4015);
nand U4295 (N_4295,N_4025,N_4042);
nor U4296 (N_4296,N_4146,N_4102);
or U4297 (N_4297,N_4149,N_4004);
and U4298 (N_4298,N_4108,N_4027);
nand U4299 (N_4299,N_4087,N_4105);
xor U4300 (N_4300,N_4194,N_4185);
xnor U4301 (N_4301,N_4066,N_4087);
or U4302 (N_4302,N_4040,N_4067);
or U4303 (N_4303,N_4171,N_4067);
nand U4304 (N_4304,N_4088,N_4093);
or U4305 (N_4305,N_4097,N_4067);
nand U4306 (N_4306,N_4076,N_4086);
xnor U4307 (N_4307,N_4104,N_4198);
and U4308 (N_4308,N_4174,N_4080);
and U4309 (N_4309,N_4197,N_4113);
nor U4310 (N_4310,N_4171,N_4049);
xor U4311 (N_4311,N_4026,N_4157);
xor U4312 (N_4312,N_4032,N_4121);
or U4313 (N_4313,N_4015,N_4117);
nand U4314 (N_4314,N_4124,N_4028);
nor U4315 (N_4315,N_4036,N_4079);
nand U4316 (N_4316,N_4161,N_4071);
or U4317 (N_4317,N_4119,N_4190);
nand U4318 (N_4318,N_4019,N_4104);
or U4319 (N_4319,N_4020,N_4001);
nor U4320 (N_4320,N_4169,N_4007);
or U4321 (N_4321,N_4130,N_4052);
xnor U4322 (N_4322,N_4088,N_4103);
nand U4323 (N_4323,N_4196,N_4044);
nand U4324 (N_4324,N_4139,N_4190);
nor U4325 (N_4325,N_4004,N_4114);
and U4326 (N_4326,N_4189,N_4092);
or U4327 (N_4327,N_4171,N_4092);
xor U4328 (N_4328,N_4190,N_4188);
and U4329 (N_4329,N_4006,N_4053);
xor U4330 (N_4330,N_4191,N_4015);
and U4331 (N_4331,N_4125,N_4088);
xnor U4332 (N_4332,N_4004,N_4152);
and U4333 (N_4333,N_4071,N_4085);
or U4334 (N_4334,N_4089,N_4125);
and U4335 (N_4335,N_4037,N_4143);
and U4336 (N_4336,N_4118,N_4092);
nor U4337 (N_4337,N_4166,N_4025);
and U4338 (N_4338,N_4005,N_4130);
nand U4339 (N_4339,N_4117,N_4024);
or U4340 (N_4340,N_4080,N_4066);
xnor U4341 (N_4341,N_4167,N_4089);
nand U4342 (N_4342,N_4066,N_4147);
nand U4343 (N_4343,N_4132,N_4095);
or U4344 (N_4344,N_4193,N_4118);
or U4345 (N_4345,N_4149,N_4019);
or U4346 (N_4346,N_4191,N_4195);
nor U4347 (N_4347,N_4106,N_4059);
and U4348 (N_4348,N_4109,N_4097);
nor U4349 (N_4349,N_4112,N_4086);
xor U4350 (N_4350,N_4057,N_4027);
xnor U4351 (N_4351,N_4101,N_4109);
xnor U4352 (N_4352,N_4016,N_4037);
and U4353 (N_4353,N_4010,N_4133);
nor U4354 (N_4354,N_4147,N_4102);
nor U4355 (N_4355,N_4171,N_4101);
xor U4356 (N_4356,N_4099,N_4066);
xnor U4357 (N_4357,N_4060,N_4144);
and U4358 (N_4358,N_4029,N_4103);
xnor U4359 (N_4359,N_4120,N_4177);
nand U4360 (N_4360,N_4170,N_4181);
nor U4361 (N_4361,N_4106,N_4050);
or U4362 (N_4362,N_4185,N_4029);
nand U4363 (N_4363,N_4036,N_4161);
and U4364 (N_4364,N_4167,N_4036);
or U4365 (N_4365,N_4164,N_4009);
xor U4366 (N_4366,N_4070,N_4154);
xor U4367 (N_4367,N_4073,N_4009);
or U4368 (N_4368,N_4033,N_4170);
nand U4369 (N_4369,N_4066,N_4161);
or U4370 (N_4370,N_4065,N_4022);
nand U4371 (N_4371,N_4023,N_4061);
nand U4372 (N_4372,N_4111,N_4169);
or U4373 (N_4373,N_4025,N_4083);
and U4374 (N_4374,N_4043,N_4071);
nand U4375 (N_4375,N_4014,N_4057);
and U4376 (N_4376,N_4023,N_4182);
xor U4377 (N_4377,N_4060,N_4031);
nor U4378 (N_4378,N_4185,N_4073);
or U4379 (N_4379,N_4091,N_4012);
or U4380 (N_4380,N_4178,N_4018);
nor U4381 (N_4381,N_4147,N_4091);
nor U4382 (N_4382,N_4058,N_4181);
nor U4383 (N_4383,N_4034,N_4105);
or U4384 (N_4384,N_4078,N_4022);
xor U4385 (N_4385,N_4033,N_4101);
xor U4386 (N_4386,N_4107,N_4040);
or U4387 (N_4387,N_4109,N_4037);
nor U4388 (N_4388,N_4046,N_4087);
xor U4389 (N_4389,N_4069,N_4174);
nand U4390 (N_4390,N_4153,N_4026);
xor U4391 (N_4391,N_4102,N_4028);
nor U4392 (N_4392,N_4066,N_4046);
xor U4393 (N_4393,N_4169,N_4103);
and U4394 (N_4394,N_4085,N_4093);
nor U4395 (N_4395,N_4157,N_4165);
xnor U4396 (N_4396,N_4152,N_4185);
and U4397 (N_4397,N_4078,N_4198);
xnor U4398 (N_4398,N_4085,N_4083);
nand U4399 (N_4399,N_4119,N_4045);
or U4400 (N_4400,N_4321,N_4396);
xor U4401 (N_4401,N_4279,N_4201);
nand U4402 (N_4402,N_4397,N_4374);
xor U4403 (N_4403,N_4338,N_4282);
xor U4404 (N_4404,N_4209,N_4270);
nor U4405 (N_4405,N_4277,N_4356);
nor U4406 (N_4406,N_4389,N_4248);
nand U4407 (N_4407,N_4293,N_4238);
nand U4408 (N_4408,N_4269,N_4202);
nor U4409 (N_4409,N_4342,N_4292);
or U4410 (N_4410,N_4243,N_4272);
and U4411 (N_4411,N_4365,N_4263);
nand U4412 (N_4412,N_4325,N_4284);
nand U4413 (N_4413,N_4247,N_4380);
nand U4414 (N_4414,N_4215,N_4262);
nor U4415 (N_4415,N_4239,N_4391);
and U4416 (N_4416,N_4367,N_4312);
nor U4417 (N_4417,N_4348,N_4289);
or U4418 (N_4418,N_4395,N_4265);
nor U4419 (N_4419,N_4343,N_4291);
or U4420 (N_4420,N_4274,N_4366);
or U4421 (N_4421,N_4317,N_4359);
nor U4422 (N_4422,N_4370,N_4223);
or U4423 (N_4423,N_4300,N_4288);
and U4424 (N_4424,N_4252,N_4222);
nor U4425 (N_4425,N_4382,N_4254);
or U4426 (N_4426,N_4392,N_4332);
xor U4427 (N_4427,N_4286,N_4226);
and U4428 (N_4428,N_4221,N_4232);
nor U4429 (N_4429,N_4257,N_4258);
or U4430 (N_4430,N_4361,N_4281);
xor U4431 (N_4431,N_4245,N_4302);
and U4432 (N_4432,N_4358,N_4373);
and U4433 (N_4433,N_4255,N_4377);
nand U4434 (N_4434,N_4339,N_4384);
xnor U4435 (N_4435,N_4346,N_4309);
or U4436 (N_4436,N_4360,N_4335);
xnor U4437 (N_4437,N_4313,N_4208);
or U4438 (N_4438,N_4331,N_4318);
xnor U4439 (N_4439,N_4350,N_4319);
or U4440 (N_4440,N_4344,N_4271);
or U4441 (N_4441,N_4285,N_4362);
nand U4442 (N_4442,N_4204,N_4236);
xor U4443 (N_4443,N_4212,N_4235);
or U4444 (N_4444,N_4294,N_4320);
nand U4445 (N_4445,N_4234,N_4357);
nor U4446 (N_4446,N_4267,N_4328);
nand U4447 (N_4447,N_4301,N_4227);
xnor U4448 (N_4448,N_4347,N_4295);
or U4449 (N_4449,N_4379,N_4203);
nor U4450 (N_4450,N_4371,N_4375);
xor U4451 (N_4451,N_4399,N_4364);
xnor U4452 (N_4452,N_4290,N_4388);
or U4453 (N_4453,N_4322,N_4207);
xnor U4454 (N_4454,N_4349,N_4308);
and U4455 (N_4455,N_4230,N_4278);
nand U4456 (N_4456,N_4369,N_4345);
nand U4457 (N_4457,N_4326,N_4363);
or U4458 (N_4458,N_4376,N_4217);
or U4459 (N_4459,N_4219,N_4250);
nor U4460 (N_4460,N_4336,N_4303);
and U4461 (N_4461,N_4228,N_4280);
or U4462 (N_4462,N_4244,N_4283);
nand U4463 (N_4463,N_4225,N_4206);
nor U4464 (N_4464,N_4275,N_4394);
or U4465 (N_4465,N_4390,N_4211);
xnor U4466 (N_4466,N_4372,N_4261);
and U4467 (N_4467,N_4315,N_4220);
or U4468 (N_4468,N_4256,N_4340);
nand U4469 (N_4469,N_4299,N_4341);
xor U4470 (N_4470,N_4200,N_4378);
nor U4471 (N_4471,N_4398,N_4205);
xnor U4472 (N_4472,N_4337,N_4264);
or U4473 (N_4473,N_4314,N_4296);
or U4474 (N_4474,N_4324,N_4229);
nand U4475 (N_4475,N_4354,N_4237);
nor U4476 (N_4476,N_4249,N_4316);
xor U4477 (N_4477,N_4306,N_4297);
and U4478 (N_4478,N_4353,N_4246);
or U4479 (N_4479,N_4351,N_4276);
and U4480 (N_4480,N_4233,N_4210);
nand U4481 (N_4481,N_4214,N_4330);
and U4482 (N_4482,N_4329,N_4273);
nand U4483 (N_4483,N_4304,N_4393);
nand U4484 (N_4484,N_4386,N_4307);
or U4485 (N_4485,N_4352,N_4241);
nand U4486 (N_4486,N_4218,N_4355);
or U4487 (N_4487,N_4287,N_4213);
and U4488 (N_4488,N_4251,N_4333);
and U4489 (N_4489,N_4334,N_4240);
nor U4490 (N_4490,N_4242,N_4385);
nand U4491 (N_4491,N_4383,N_4298);
xor U4492 (N_4492,N_4216,N_4266);
and U4493 (N_4493,N_4311,N_4310);
nand U4494 (N_4494,N_4231,N_4268);
and U4495 (N_4495,N_4305,N_4224);
or U4496 (N_4496,N_4327,N_4323);
nand U4497 (N_4497,N_4260,N_4387);
xnor U4498 (N_4498,N_4381,N_4259);
xnor U4499 (N_4499,N_4368,N_4253);
or U4500 (N_4500,N_4265,N_4239);
nand U4501 (N_4501,N_4259,N_4377);
or U4502 (N_4502,N_4220,N_4248);
nand U4503 (N_4503,N_4289,N_4394);
nand U4504 (N_4504,N_4215,N_4348);
and U4505 (N_4505,N_4340,N_4249);
nor U4506 (N_4506,N_4327,N_4229);
xnor U4507 (N_4507,N_4204,N_4271);
nor U4508 (N_4508,N_4345,N_4301);
nand U4509 (N_4509,N_4238,N_4274);
nand U4510 (N_4510,N_4229,N_4345);
and U4511 (N_4511,N_4357,N_4350);
or U4512 (N_4512,N_4343,N_4339);
or U4513 (N_4513,N_4269,N_4280);
nor U4514 (N_4514,N_4251,N_4342);
and U4515 (N_4515,N_4220,N_4209);
xor U4516 (N_4516,N_4317,N_4213);
nand U4517 (N_4517,N_4325,N_4346);
and U4518 (N_4518,N_4395,N_4378);
nand U4519 (N_4519,N_4372,N_4380);
or U4520 (N_4520,N_4296,N_4227);
xor U4521 (N_4521,N_4378,N_4278);
xnor U4522 (N_4522,N_4295,N_4289);
xnor U4523 (N_4523,N_4295,N_4390);
nor U4524 (N_4524,N_4259,N_4362);
nor U4525 (N_4525,N_4228,N_4267);
xnor U4526 (N_4526,N_4230,N_4284);
xor U4527 (N_4527,N_4346,N_4289);
or U4528 (N_4528,N_4262,N_4237);
or U4529 (N_4529,N_4242,N_4232);
or U4530 (N_4530,N_4347,N_4232);
xnor U4531 (N_4531,N_4266,N_4268);
nor U4532 (N_4532,N_4397,N_4354);
nor U4533 (N_4533,N_4213,N_4228);
nor U4534 (N_4534,N_4315,N_4337);
nand U4535 (N_4535,N_4307,N_4374);
and U4536 (N_4536,N_4203,N_4302);
xnor U4537 (N_4537,N_4209,N_4295);
and U4538 (N_4538,N_4289,N_4385);
and U4539 (N_4539,N_4374,N_4294);
or U4540 (N_4540,N_4245,N_4237);
xnor U4541 (N_4541,N_4288,N_4398);
xnor U4542 (N_4542,N_4200,N_4246);
nor U4543 (N_4543,N_4210,N_4258);
nor U4544 (N_4544,N_4253,N_4243);
nand U4545 (N_4545,N_4212,N_4277);
nor U4546 (N_4546,N_4350,N_4370);
nand U4547 (N_4547,N_4254,N_4223);
or U4548 (N_4548,N_4267,N_4220);
and U4549 (N_4549,N_4325,N_4337);
nor U4550 (N_4550,N_4394,N_4231);
or U4551 (N_4551,N_4395,N_4376);
nor U4552 (N_4552,N_4255,N_4390);
nand U4553 (N_4553,N_4387,N_4381);
nor U4554 (N_4554,N_4325,N_4254);
xnor U4555 (N_4555,N_4265,N_4202);
xor U4556 (N_4556,N_4273,N_4359);
nor U4557 (N_4557,N_4399,N_4271);
nand U4558 (N_4558,N_4338,N_4290);
nor U4559 (N_4559,N_4318,N_4367);
xnor U4560 (N_4560,N_4328,N_4314);
nor U4561 (N_4561,N_4397,N_4310);
and U4562 (N_4562,N_4328,N_4222);
or U4563 (N_4563,N_4337,N_4336);
or U4564 (N_4564,N_4251,N_4374);
or U4565 (N_4565,N_4237,N_4398);
nand U4566 (N_4566,N_4369,N_4215);
xor U4567 (N_4567,N_4330,N_4315);
and U4568 (N_4568,N_4365,N_4236);
nor U4569 (N_4569,N_4240,N_4329);
nor U4570 (N_4570,N_4261,N_4285);
and U4571 (N_4571,N_4224,N_4230);
nand U4572 (N_4572,N_4369,N_4327);
nand U4573 (N_4573,N_4392,N_4242);
xor U4574 (N_4574,N_4295,N_4217);
and U4575 (N_4575,N_4281,N_4385);
xor U4576 (N_4576,N_4287,N_4301);
or U4577 (N_4577,N_4232,N_4310);
nand U4578 (N_4578,N_4296,N_4341);
and U4579 (N_4579,N_4325,N_4361);
xor U4580 (N_4580,N_4236,N_4306);
or U4581 (N_4581,N_4254,N_4336);
and U4582 (N_4582,N_4390,N_4294);
and U4583 (N_4583,N_4333,N_4309);
nand U4584 (N_4584,N_4242,N_4231);
nand U4585 (N_4585,N_4245,N_4247);
or U4586 (N_4586,N_4336,N_4387);
or U4587 (N_4587,N_4253,N_4286);
nand U4588 (N_4588,N_4355,N_4389);
nand U4589 (N_4589,N_4297,N_4386);
nand U4590 (N_4590,N_4263,N_4252);
xnor U4591 (N_4591,N_4392,N_4256);
and U4592 (N_4592,N_4259,N_4241);
and U4593 (N_4593,N_4368,N_4353);
nor U4594 (N_4594,N_4376,N_4270);
nor U4595 (N_4595,N_4224,N_4257);
nand U4596 (N_4596,N_4267,N_4362);
nor U4597 (N_4597,N_4378,N_4262);
and U4598 (N_4598,N_4271,N_4374);
nor U4599 (N_4599,N_4269,N_4394);
xor U4600 (N_4600,N_4567,N_4445);
xor U4601 (N_4601,N_4588,N_4486);
and U4602 (N_4602,N_4419,N_4585);
xor U4603 (N_4603,N_4519,N_4430);
or U4604 (N_4604,N_4540,N_4403);
nor U4605 (N_4605,N_4539,N_4418);
nand U4606 (N_4606,N_4554,N_4425);
nand U4607 (N_4607,N_4458,N_4504);
nand U4608 (N_4608,N_4479,N_4562);
xnor U4609 (N_4609,N_4571,N_4447);
or U4610 (N_4610,N_4513,N_4484);
nor U4611 (N_4611,N_4532,N_4498);
nor U4612 (N_4612,N_4517,N_4493);
nand U4613 (N_4613,N_4515,N_4564);
nor U4614 (N_4614,N_4597,N_4443);
or U4615 (N_4615,N_4481,N_4521);
or U4616 (N_4616,N_4457,N_4590);
nor U4617 (N_4617,N_4553,N_4424);
nor U4618 (N_4618,N_4546,N_4409);
xor U4619 (N_4619,N_4527,N_4506);
and U4620 (N_4620,N_4428,N_4501);
and U4621 (N_4621,N_4496,N_4435);
or U4622 (N_4622,N_4483,N_4412);
nor U4623 (N_4623,N_4512,N_4491);
nor U4624 (N_4624,N_4534,N_4531);
xnor U4625 (N_4625,N_4505,N_4509);
nand U4626 (N_4626,N_4520,N_4561);
nor U4627 (N_4627,N_4456,N_4488);
or U4628 (N_4628,N_4475,N_4441);
xnor U4629 (N_4629,N_4576,N_4402);
xor U4630 (N_4630,N_4548,N_4551);
nor U4631 (N_4631,N_4433,N_4538);
and U4632 (N_4632,N_4480,N_4469);
nor U4633 (N_4633,N_4558,N_4490);
nand U4634 (N_4634,N_4477,N_4439);
nor U4635 (N_4635,N_4500,N_4522);
or U4636 (N_4636,N_4568,N_4463);
or U4637 (N_4637,N_4448,N_4593);
nand U4638 (N_4638,N_4495,N_4560);
nor U4639 (N_4639,N_4579,N_4533);
xnor U4640 (N_4640,N_4503,N_4452);
nand U4641 (N_4641,N_4599,N_4494);
and U4642 (N_4642,N_4537,N_4415);
nor U4643 (N_4643,N_4474,N_4581);
or U4644 (N_4644,N_4596,N_4575);
or U4645 (N_4645,N_4563,N_4423);
nor U4646 (N_4646,N_4440,N_4427);
nor U4647 (N_4647,N_4482,N_4587);
nand U4648 (N_4648,N_4489,N_4438);
nand U4649 (N_4649,N_4595,N_4429);
xnor U4650 (N_4650,N_4492,N_4454);
nor U4651 (N_4651,N_4478,N_4459);
or U4652 (N_4652,N_4507,N_4449);
xor U4653 (N_4653,N_4572,N_4543);
nand U4654 (N_4654,N_4465,N_4455);
and U4655 (N_4655,N_4528,N_4530);
and U4656 (N_4656,N_4514,N_4557);
or U4657 (N_4657,N_4591,N_4437);
xor U4658 (N_4658,N_4464,N_4404);
nor U4659 (N_4659,N_4542,N_4446);
xnor U4660 (N_4660,N_4422,N_4594);
xnor U4661 (N_4661,N_4434,N_4566);
nand U4662 (N_4662,N_4555,N_4516);
nor U4663 (N_4663,N_4547,N_4578);
nand U4664 (N_4664,N_4436,N_4577);
or U4665 (N_4665,N_4545,N_4414);
nand U4666 (N_4666,N_4518,N_4476);
and U4667 (N_4667,N_4401,N_4541);
nand U4668 (N_4668,N_4485,N_4400);
and U4669 (N_4669,N_4544,N_4450);
or U4670 (N_4670,N_4471,N_4451);
nor U4671 (N_4671,N_4470,N_4411);
xor U4672 (N_4672,N_4405,N_4598);
nand U4673 (N_4673,N_4473,N_4549);
xor U4674 (N_4674,N_4559,N_4406);
and U4675 (N_4675,N_4552,N_4573);
and U4676 (N_4676,N_4460,N_4453);
nand U4677 (N_4677,N_4580,N_4535);
nand U4678 (N_4678,N_4583,N_4442);
nand U4679 (N_4679,N_4508,N_4466);
or U4680 (N_4680,N_4550,N_4586);
and U4681 (N_4681,N_4497,N_4420);
xnor U4682 (N_4682,N_4582,N_4467);
and U4683 (N_4683,N_4556,N_4461);
or U4684 (N_4684,N_4421,N_4413);
or U4685 (N_4685,N_4417,N_4407);
and U4686 (N_4686,N_4523,N_4536);
nand U4687 (N_4687,N_4499,N_4526);
nor U4688 (N_4688,N_4444,N_4589);
or U4689 (N_4689,N_4592,N_4511);
nor U4690 (N_4690,N_4525,N_4524);
xor U4691 (N_4691,N_4408,N_4529);
or U4692 (N_4692,N_4410,N_4565);
nand U4693 (N_4693,N_4510,N_4584);
or U4694 (N_4694,N_4569,N_4574);
and U4695 (N_4695,N_4416,N_4462);
or U4696 (N_4696,N_4468,N_4487);
xor U4697 (N_4697,N_4426,N_4432);
nor U4698 (N_4698,N_4502,N_4431);
and U4699 (N_4699,N_4472,N_4570);
or U4700 (N_4700,N_4566,N_4536);
nor U4701 (N_4701,N_4564,N_4450);
nor U4702 (N_4702,N_4403,N_4567);
nor U4703 (N_4703,N_4596,N_4534);
and U4704 (N_4704,N_4552,N_4551);
xnor U4705 (N_4705,N_4407,N_4566);
nor U4706 (N_4706,N_4507,N_4470);
nor U4707 (N_4707,N_4449,N_4576);
nor U4708 (N_4708,N_4536,N_4535);
and U4709 (N_4709,N_4509,N_4450);
xnor U4710 (N_4710,N_4492,N_4409);
or U4711 (N_4711,N_4582,N_4580);
or U4712 (N_4712,N_4510,N_4570);
nor U4713 (N_4713,N_4482,N_4526);
or U4714 (N_4714,N_4494,N_4440);
or U4715 (N_4715,N_4591,N_4521);
or U4716 (N_4716,N_4439,N_4571);
nor U4717 (N_4717,N_4429,N_4517);
or U4718 (N_4718,N_4561,N_4491);
nand U4719 (N_4719,N_4597,N_4591);
or U4720 (N_4720,N_4455,N_4566);
or U4721 (N_4721,N_4594,N_4450);
nand U4722 (N_4722,N_4487,N_4493);
xor U4723 (N_4723,N_4413,N_4529);
xor U4724 (N_4724,N_4464,N_4508);
nor U4725 (N_4725,N_4444,N_4542);
or U4726 (N_4726,N_4488,N_4515);
nand U4727 (N_4727,N_4549,N_4572);
nor U4728 (N_4728,N_4447,N_4544);
or U4729 (N_4729,N_4528,N_4452);
nor U4730 (N_4730,N_4507,N_4428);
and U4731 (N_4731,N_4595,N_4527);
nor U4732 (N_4732,N_4481,N_4453);
xor U4733 (N_4733,N_4551,N_4555);
or U4734 (N_4734,N_4453,N_4593);
nor U4735 (N_4735,N_4488,N_4411);
nand U4736 (N_4736,N_4587,N_4540);
or U4737 (N_4737,N_4404,N_4420);
nand U4738 (N_4738,N_4404,N_4430);
and U4739 (N_4739,N_4425,N_4469);
nand U4740 (N_4740,N_4542,N_4484);
or U4741 (N_4741,N_4589,N_4508);
and U4742 (N_4742,N_4439,N_4525);
nor U4743 (N_4743,N_4506,N_4541);
nor U4744 (N_4744,N_4423,N_4586);
xor U4745 (N_4745,N_4475,N_4478);
xnor U4746 (N_4746,N_4411,N_4422);
or U4747 (N_4747,N_4572,N_4442);
nor U4748 (N_4748,N_4453,N_4410);
or U4749 (N_4749,N_4459,N_4429);
nor U4750 (N_4750,N_4436,N_4491);
nand U4751 (N_4751,N_4546,N_4439);
or U4752 (N_4752,N_4592,N_4572);
or U4753 (N_4753,N_4538,N_4421);
or U4754 (N_4754,N_4539,N_4570);
or U4755 (N_4755,N_4541,N_4402);
and U4756 (N_4756,N_4526,N_4427);
xnor U4757 (N_4757,N_4491,N_4435);
and U4758 (N_4758,N_4434,N_4486);
or U4759 (N_4759,N_4559,N_4487);
nor U4760 (N_4760,N_4408,N_4463);
nand U4761 (N_4761,N_4482,N_4530);
nand U4762 (N_4762,N_4508,N_4580);
and U4763 (N_4763,N_4533,N_4564);
or U4764 (N_4764,N_4506,N_4531);
nand U4765 (N_4765,N_4551,N_4569);
xor U4766 (N_4766,N_4474,N_4582);
and U4767 (N_4767,N_4452,N_4521);
or U4768 (N_4768,N_4415,N_4533);
or U4769 (N_4769,N_4467,N_4577);
or U4770 (N_4770,N_4534,N_4406);
nor U4771 (N_4771,N_4569,N_4589);
xnor U4772 (N_4772,N_4523,N_4572);
xor U4773 (N_4773,N_4430,N_4423);
xnor U4774 (N_4774,N_4408,N_4413);
and U4775 (N_4775,N_4464,N_4474);
and U4776 (N_4776,N_4507,N_4405);
or U4777 (N_4777,N_4532,N_4453);
or U4778 (N_4778,N_4521,N_4514);
nand U4779 (N_4779,N_4496,N_4448);
xnor U4780 (N_4780,N_4558,N_4420);
xor U4781 (N_4781,N_4470,N_4519);
and U4782 (N_4782,N_4574,N_4524);
xor U4783 (N_4783,N_4525,N_4417);
nand U4784 (N_4784,N_4562,N_4518);
nor U4785 (N_4785,N_4519,N_4521);
nor U4786 (N_4786,N_4477,N_4456);
nand U4787 (N_4787,N_4544,N_4474);
xnor U4788 (N_4788,N_4458,N_4597);
nor U4789 (N_4789,N_4476,N_4517);
nand U4790 (N_4790,N_4572,N_4520);
nand U4791 (N_4791,N_4573,N_4592);
and U4792 (N_4792,N_4501,N_4527);
nand U4793 (N_4793,N_4491,N_4477);
xnor U4794 (N_4794,N_4505,N_4500);
and U4795 (N_4795,N_4584,N_4534);
nor U4796 (N_4796,N_4524,N_4482);
and U4797 (N_4797,N_4484,N_4501);
or U4798 (N_4798,N_4439,N_4461);
or U4799 (N_4799,N_4531,N_4567);
nand U4800 (N_4800,N_4710,N_4605);
and U4801 (N_4801,N_4781,N_4727);
xor U4802 (N_4802,N_4657,N_4646);
xor U4803 (N_4803,N_4742,N_4728);
or U4804 (N_4804,N_4725,N_4741);
nand U4805 (N_4805,N_4723,N_4622);
and U4806 (N_4806,N_4667,N_4771);
nor U4807 (N_4807,N_4706,N_4733);
nor U4808 (N_4808,N_4719,N_4743);
nor U4809 (N_4809,N_4798,N_4778);
xor U4810 (N_4810,N_4751,N_4775);
or U4811 (N_4811,N_4624,N_4626);
nand U4812 (N_4812,N_4793,N_4707);
xnor U4813 (N_4813,N_4752,N_4668);
and U4814 (N_4814,N_4740,N_4628);
nor U4815 (N_4815,N_4696,N_4653);
and U4816 (N_4816,N_4658,N_4656);
and U4817 (N_4817,N_4690,N_4625);
or U4818 (N_4818,N_4747,N_4693);
nor U4819 (N_4819,N_4699,N_4673);
and U4820 (N_4820,N_4601,N_4744);
or U4821 (N_4821,N_4615,N_4670);
nor U4822 (N_4822,N_4634,N_4722);
xnor U4823 (N_4823,N_4730,N_4799);
xor U4824 (N_4824,N_4791,N_4619);
xor U4825 (N_4825,N_4650,N_4678);
nor U4826 (N_4826,N_4633,N_4635);
nand U4827 (N_4827,N_4623,N_4754);
nor U4828 (N_4828,N_4756,N_4684);
or U4829 (N_4829,N_4685,N_4738);
nor U4830 (N_4830,N_4726,N_4702);
and U4831 (N_4831,N_4765,N_4636);
xnor U4832 (N_4832,N_4796,N_4716);
or U4833 (N_4833,N_4618,N_4651);
nor U4834 (N_4834,N_4704,N_4645);
xnor U4835 (N_4835,N_4682,N_4613);
or U4836 (N_4836,N_4715,N_4637);
nand U4837 (N_4837,N_4647,N_4611);
nand U4838 (N_4838,N_4768,N_4773);
and U4839 (N_4839,N_4680,N_4753);
and U4840 (N_4840,N_4664,N_4714);
nor U4841 (N_4841,N_4770,N_4705);
xor U4842 (N_4842,N_4772,N_4708);
nor U4843 (N_4843,N_4787,N_4679);
xnor U4844 (N_4844,N_4766,N_4709);
or U4845 (N_4845,N_4736,N_4717);
nor U4846 (N_4846,N_4639,N_4612);
and U4847 (N_4847,N_4698,N_4759);
xor U4848 (N_4848,N_4602,N_4688);
nor U4849 (N_4849,N_4607,N_4786);
and U4850 (N_4850,N_4643,N_4780);
nor U4851 (N_4851,N_4711,N_4674);
or U4852 (N_4852,N_4692,N_4750);
and U4853 (N_4853,N_4671,N_4764);
or U4854 (N_4854,N_4649,N_4795);
nor U4855 (N_4855,N_4642,N_4660);
xnor U4856 (N_4856,N_4757,N_4669);
or U4857 (N_4857,N_4659,N_4779);
or U4858 (N_4858,N_4703,N_4640);
and U4859 (N_4859,N_4789,N_4629);
xnor U4860 (N_4860,N_4769,N_4737);
nor U4861 (N_4861,N_4617,N_4675);
or U4862 (N_4862,N_4755,N_4713);
nor U4863 (N_4863,N_4631,N_4712);
and U4864 (N_4864,N_4638,N_4666);
or U4865 (N_4865,N_4724,N_4630);
and U4866 (N_4866,N_4784,N_4677);
xnor U4867 (N_4867,N_4762,N_4739);
and U4868 (N_4868,N_4608,N_4600);
xor U4869 (N_4869,N_4610,N_4697);
nor U4870 (N_4870,N_4603,N_4641);
nand U4871 (N_4871,N_4687,N_4721);
nor U4872 (N_4872,N_4783,N_4788);
and U4873 (N_4873,N_4665,N_4694);
nand U4874 (N_4874,N_4606,N_4689);
nand U4875 (N_4875,N_4662,N_4661);
and U4876 (N_4876,N_4609,N_4621);
nand U4877 (N_4877,N_4734,N_4760);
nand U4878 (N_4878,N_4748,N_4763);
and U4879 (N_4879,N_4720,N_4681);
or U4880 (N_4880,N_4700,N_4676);
or U4881 (N_4881,N_4735,N_4745);
and U4882 (N_4882,N_4691,N_4655);
or U4883 (N_4883,N_4732,N_4774);
and U4884 (N_4884,N_4644,N_4663);
or U4885 (N_4885,N_4652,N_4782);
nand U4886 (N_4886,N_4614,N_4746);
xor U4887 (N_4887,N_4654,N_4718);
or U4888 (N_4888,N_4797,N_4776);
nand U4889 (N_4889,N_4632,N_4785);
xor U4890 (N_4890,N_4767,N_4627);
nor U4891 (N_4891,N_4686,N_4648);
or U4892 (N_4892,N_4792,N_4790);
nor U4893 (N_4893,N_4695,N_4731);
or U4894 (N_4894,N_4701,N_4620);
nand U4895 (N_4895,N_4604,N_4616);
xnor U4896 (N_4896,N_4683,N_4672);
and U4897 (N_4897,N_4777,N_4729);
nor U4898 (N_4898,N_4749,N_4758);
nor U4899 (N_4899,N_4794,N_4761);
and U4900 (N_4900,N_4613,N_4798);
nor U4901 (N_4901,N_4726,N_4636);
and U4902 (N_4902,N_4717,N_4701);
nor U4903 (N_4903,N_4754,N_4693);
nor U4904 (N_4904,N_4705,N_4716);
xor U4905 (N_4905,N_4768,N_4695);
xor U4906 (N_4906,N_4670,N_4668);
nor U4907 (N_4907,N_4647,N_4767);
and U4908 (N_4908,N_4791,N_4772);
xnor U4909 (N_4909,N_4703,N_4621);
and U4910 (N_4910,N_4662,N_4645);
and U4911 (N_4911,N_4657,N_4699);
or U4912 (N_4912,N_4667,N_4610);
nor U4913 (N_4913,N_4769,N_4700);
xnor U4914 (N_4914,N_4625,N_4733);
and U4915 (N_4915,N_4794,N_4726);
and U4916 (N_4916,N_4677,N_4680);
and U4917 (N_4917,N_4720,N_4699);
or U4918 (N_4918,N_4704,N_4746);
nand U4919 (N_4919,N_4691,N_4663);
or U4920 (N_4920,N_4627,N_4787);
or U4921 (N_4921,N_4635,N_4662);
xor U4922 (N_4922,N_4656,N_4716);
nand U4923 (N_4923,N_4758,N_4700);
xor U4924 (N_4924,N_4746,N_4650);
nand U4925 (N_4925,N_4683,N_4747);
nor U4926 (N_4926,N_4791,N_4656);
nand U4927 (N_4927,N_4627,N_4706);
or U4928 (N_4928,N_4761,N_4627);
and U4929 (N_4929,N_4781,N_4739);
nand U4930 (N_4930,N_4745,N_4639);
xnor U4931 (N_4931,N_4607,N_4763);
xnor U4932 (N_4932,N_4765,N_4617);
or U4933 (N_4933,N_4637,N_4681);
nor U4934 (N_4934,N_4764,N_4688);
xor U4935 (N_4935,N_4678,N_4753);
nor U4936 (N_4936,N_4679,N_4715);
nor U4937 (N_4937,N_4689,N_4766);
xnor U4938 (N_4938,N_4689,N_4605);
xnor U4939 (N_4939,N_4722,N_4625);
nor U4940 (N_4940,N_4718,N_4769);
xor U4941 (N_4941,N_4679,N_4766);
and U4942 (N_4942,N_4648,N_4717);
xnor U4943 (N_4943,N_4641,N_4767);
xor U4944 (N_4944,N_4644,N_4752);
nand U4945 (N_4945,N_4657,N_4729);
xor U4946 (N_4946,N_4677,N_4715);
nor U4947 (N_4947,N_4798,N_4736);
nand U4948 (N_4948,N_4712,N_4681);
or U4949 (N_4949,N_4748,N_4636);
nor U4950 (N_4950,N_4782,N_4649);
nor U4951 (N_4951,N_4724,N_4735);
and U4952 (N_4952,N_4726,N_4704);
nand U4953 (N_4953,N_4739,N_4610);
nor U4954 (N_4954,N_4773,N_4737);
nand U4955 (N_4955,N_4685,N_4684);
and U4956 (N_4956,N_4750,N_4736);
nand U4957 (N_4957,N_4656,N_4644);
nor U4958 (N_4958,N_4779,N_4752);
or U4959 (N_4959,N_4688,N_4711);
nand U4960 (N_4960,N_4687,N_4745);
xnor U4961 (N_4961,N_4753,N_4621);
nor U4962 (N_4962,N_4783,N_4753);
nand U4963 (N_4963,N_4643,N_4753);
or U4964 (N_4964,N_4712,N_4786);
xnor U4965 (N_4965,N_4779,N_4782);
or U4966 (N_4966,N_4684,N_4617);
and U4967 (N_4967,N_4710,N_4793);
nor U4968 (N_4968,N_4717,N_4693);
nor U4969 (N_4969,N_4729,N_4717);
nand U4970 (N_4970,N_4715,N_4707);
nand U4971 (N_4971,N_4760,N_4773);
or U4972 (N_4972,N_4662,N_4782);
xnor U4973 (N_4973,N_4683,N_4682);
nand U4974 (N_4974,N_4729,N_4759);
or U4975 (N_4975,N_4693,N_4629);
nand U4976 (N_4976,N_4751,N_4794);
nand U4977 (N_4977,N_4764,N_4784);
or U4978 (N_4978,N_4736,N_4710);
or U4979 (N_4979,N_4700,N_4793);
or U4980 (N_4980,N_4758,N_4772);
nand U4981 (N_4981,N_4618,N_4703);
and U4982 (N_4982,N_4698,N_4699);
nor U4983 (N_4983,N_4716,N_4626);
and U4984 (N_4984,N_4615,N_4656);
nand U4985 (N_4985,N_4683,N_4692);
and U4986 (N_4986,N_4664,N_4798);
and U4987 (N_4987,N_4744,N_4713);
xnor U4988 (N_4988,N_4730,N_4703);
or U4989 (N_4989,N_4735,N_4730);
or U4990 (N_4990,N_4792,N_4756);
and U4991 (N_4991,N_4796,N_4774);
nand U4992 (N_4992,N_4720,N_4630);
or U4993 (N_4993,N_4782,N_4640);
nor U4994 (N_4994,N_4631,N_4671);
and U4995 (N_4995,N_4651,N_4661);
nor U4996 (N_4996,N_4768,N_4732);
nor U4997 (N_4997,N_4728,N_4720);
or U4998 (N_4998,N_4780,N_4708);
nand U4999 (N_4999,N_4771,N_4622);
nand U5000 (N_5000,N_4872,N_4918);
nand U5001 (N_5001,N_4861,N_4889);
and U5002 (N_5002,N_4909,N_4848);
and U5003 (N_5003,N_4945,N_4956);
nand U5004 (N_5004,N_4953,N_4813);
xnor U5005 (N_5005,N_4951,N_4862);
xnor U5006 (N_5006,N_4850,N_4892);
nand U5007 (N_5007,N_4943,N_4901);
or U5008 (N_5008,N_4845,N_4841);
nand U5009 (N_5009,N_4912,N_4973);
and U5010 (N_5010,N_4883,N_4990);
or U5011 (N_5011,N_4869,N_4890);
and U5012 (N_5012,N_4871,N_4975);
or U5013 (N_5013,N_4969,N_4941);
xnor U5014 (N_5014,N_4991,N_4961);
xnor U5015 (N_5015,N_4919,N_4838);
nand U5016 (N_5016,N_4930,N_4939);
and U5017 (N_5017,N_4824,N_4966);
nor U5018 (N_5018,N_4825,N_4856);
or U5019 (N_5019,N_4834,N_4952);
xor U5020 (N_5020,N_4979,N_4882);
nor U5021 (N_5021,N_4935,N_4873);
nor U5022 (N_5022,N_4819,N_4926);
or U5023 (N_5023,N_4829,N_4881);
nand U5024 (N_5024,N_4996,N_4895);
or U5025 (N_5025,N_4851,N_4947);
nand U5026 (N_5026,N_4923,N_4921);
and U5027 (N_5027,N_4839,N_4807);
or U5028 (N_5028,N_4927,N_4978);
or U5029 (N_5029,N_4897,N_4955);
or U5030 (N_5030,N_4844,N_4899);
and U5031 (N_5031,N_4977,N_4828);
xnor U5032 (N_5032,N_4863,N_4925);
and U5033 (N_5033,N_4976,N_4870);
nor U5034 (N_5034,N_4864,N_4866);
xnor U5035 (N_5035,N_4910,N_4971);
or U5036 (N_5036,N_4960,N_4997);
xor U5037 (N_5037,N_4994,N_4988);
or U5038 (N_5038,N_4815,N_4808);
xor U5039 (N_5039,N_4974,N_4984);
xnor U5040 (N_5040,N_4833,N_4893);
and U5041 (N_5041,N_4809,N_4868);
nand U5042 (N_5042,N_4993,N_4888);
nand U5043 (N_5043,N_4922,N_4820);
xnor U5044 (N_5044,N_4878,N_4875);
and U5045 (N_5045,N_4906,N_4818);
nand U5046 (N_5046,N_4936,N_4934);
nor U5047 (N_5047,N_4831,N_4902);
nor U5048 (N_5048,N_4987,N_4985);
xor U5049 (N_5049,N_4814,N_4886);
nor U5050 (N_5050,N_4836,N_4865);
and U5051 (N_5051,N_4822,N_4887);
or U5052 (N_5052,N_4900,N_4913);
xor U5053 (N_5053,N_4964,N_4933);
xnor U5054 (N_5054,N_4903,N_4931);
or U5055 (N_5055,N_4908,N_4803);
and U5056 (N_5056,N_4959,N_4884);
or U5057 (N_5057,N_4904,N_4920);
and U5058 (N_5058,N_4894,N_4891);
or U5059 (N_5059,N_4837,N_4911);
and U5060 (N_5060,N_4957,N_4802);
nand U5061 (N_5061,N_4958,N_4847);
or U5062 (N_5062,N_4898,N_4948);
nor U5063 (N_5063,N_4924,N_4981);
and U5064 (N_5064,N_4998,N_4980);
nor U5065 (N_5065,N_4995,N_4929);
or U5066 (N_5066,N_4972,N_4867);
nor U5067 (N_5067,N_4907,N_4982);
or U5068 (N_5068,N_4846,N_4821);
xnor U5069 (N_5069,N_4858,N_4855);
or U5070 (N_5070,N_4876,N_4812);
or U5071 (N_5071,N_4810,N_4874);
xnor U5072 (N_5072,N_4963,N_4938);
nand U5073 (N_5073,N_4949,N_4860);
nand U5074 (N_5074,N_4970,N_4852);
nor U5075 (N_5075,N_4999,N_4857);
nand U5076 (N_5076,N_4849,N_4896);
or U5077 (N_5077,N_4986,N_4937);
and U5078 (N_5078,N_4917,N_4811);
and U5079 (N_5079,N_4940,N_4968);
nor U5080 (N_5080,N_4905,N_4805);
nand U5081 (N_5081,N_4880,N_4801);
nor U5082 (N_5082,N_4826,N_4954);
nor U5083 (N_5083,N_4944,N_4832);
xor U5084 (N_5084,N_4827,N_4804);
xor U5085 (N_5085,N_4840,N_4853);
xnor U5086 (N_5086,N_4835,N_4946);
nand U5087 (N_5087,N_4989,N_4817);
or U5088 (N_5088,N_4950,N_4806);
xor U5089 (N_5089,N_4877,N_4830);
nand U5090 (N_5090,N_4965,N_4916);
xnor U5091 (N_5091,N_4859,N_4962);
or U5092 (N_5092,N_4800,N_4823);
and U5093 (N_5093,N_4843,N_4879);
xor U5094 (N_5094,N_4942,N_4967);
nand U5095 (N_5095,N_4992,N_4914);
nor U5096 (N_5096,N_4915,N_4983);
and U5097 (N_5097,N_4854,N_4816);
nor U5098 (N_5098,N_4842,N_4932);
and U5099 (N_5099,N_4928,N_4885);
or U5100 (N_5100,N_4923,N_4894);
or U5101 (N_5101,N_4803,N_4876);
or U5102 (N_5102,N_4894,N_4916);
nand U5103 (N_5103,N_4906,N_4932);
nand U5104 (N_5104,N_4873,N_4823);
nand U5105 (N_5105,N_4893,N_4880);
nand U5106 (N_5106,N_4822,N_4832);
and U5107 (N_5107,N_4945,N_4855);
nand U5108 (N_5108,N_4822,N_4989);
or U5109 (N_5109,N_4862,N_4988);
or U5110 (N_5110,N_4998,N_4863);
xnor U5111 (N_5111,N_4862,N_4866);
or U5112 (N_5112,N_4922,N_4906);
xor U5113 (N_5113,N_4946,N_4888);
and U5114 (N_5114,N_4991,N_4833);
nand U5115 (N_5115,N_4830,N_4963);
nor U5116 (N_5116,N_4893,N_4836);
xnor U5117 (N_5117,N_4937,N_4824);
xnor U5118 (N_5118,N_4840,N_4850);
nor U5119 (N_5119,N_4821,N_4844);
or U5120 (N_5120,N_4945,N_4952);
and U5121 (N_5121,N_4912,N_4975);
xnor U5122 (N_5122,N_4802,N_4955);
and U5123 (N_5123,N_4844,N_4895);
xor U5124 (N_5124,N_4993,N_4970);
and U5125 (N_5125,N_4965,N_4966);
and U5126 (N_5126,N_4816,N_4934);
and U5127 (N_5127,N_4882,N_4932);
nand U5128 (N_5128,N_4978,N_4881);
nor U5129 (N_5129,N_4986,N_4951);
nand U5130 (N_5130,N_4830,N_4857);
nor U5131 (N_5131,N_4896,N_4860);
or U5132 (N_5132,N_4916,N_4881);
xnor U5133 (N_5133,N_4854,N_4856);
xnor U5134 (N_5134,N_4850,N_4813);
nand U5135 (N_5135,N_4824,N_4835);
nand U5136 (N_5136,N_4887,N_4976);
nor U5137 (N_5137,N_4974,N_4944);
xor U5138 (N_5138,N_4815,N_4912);
or U5139 (N_5139,N_4861,N_4846);
or U5140 (N_5140,N_4834,N_4939);
nor U5141 (N_5141,N_4936,N_4997);
nor U5142 (N_5142,N_4927,N_4906);
nor U5143 (N_5143,N_4982,N_4963);
xor U5144 (N_5144,N_4928,N_4949);
nand U5145 (N_5145,N_4866,N_4998);
nand U5146 (N_5146,N_4885,N_4851);
nor U5147 (N_5147,N_4870,N_4848);
xor U5148 (N_5148,N_4857,N_4859);
and U5149 (N_5149,N_4990,N_4922);
xnor U5150 (N_5150,N_4985,N_4855);
or U5151 (N_5151,N_4853,N_4950);
and U5152 (N_5152,N_4977,N_4953);
and U5153 (N_5153,N_4984,N_4822);
nor U5154 (N_5154,N_4976,N_4990);
nor U5155 (N_5155,N_4837,N_4930);
nor U5156 (N_5156,N_4955,N_4924);
nor U5157 (N_5157,N_4844,N_4936);
nand U5158 (N_5158,N_4813,N_4886);
nor U5159 (N_5159,N_4950,N_4885);
and U5160 (N_5160,N_4887,N_4985);
nor U5161 (N_5161,N_4894,N_4818);
xnor U5162 (N_5162,N_4973,N_4892);
or U5163 (N_5163,N_4971,N_4889);
or U5164 (N_5164,N_4996,N_4814);
or U5165 (N_5165,N_4963,N_4846);
and U5166 (N_5166,N_4987,N_4850);
and U5167 (N_5167,N_4816,N_4975);
nand U5168 (N_5168,N_4986,N_4815);
nor U5169 (N_5169,N_4965,N_4957);
nand U5170 (N_5170,N_4955,N_4882);
nor U5171 (N_5171,N_4868,N_4826);
or U5172 (N_5172,N_4848,N_4888);
or U5173 (N_5173,N_4994,N_4841);
nand U5174 (N_5174,N_4918,N_4967);
and U5175 (N_5175,N_4804,N_4819);
nor U5176 (N_5176,N_4982,N_4991);
and U5177 (N_5177,N_4812,N_4874);
nor U5178 (N_5178,N_4962,N_4991);
xor U5179 (N_5179,N_4919,N_4894);
nor U5180 (N_5180,N_4802,N_4905);
nand U5181 (N_5181,N_4979,N_4802);
and U5182 (N_5182,N_4982,N_4972);
or U5183 (N_5183,N_4920,N_4878);
or U5184 (N_5184,N_4963,N_4900);
nand U5185 (N_5185,N_4850,N_4980);
and U5186 (N_5186,N_4968,N_4817);
and U5187 (N_5187,N_4819,N_4999);
nand U5188 (N_5188,N_4840,N_4921);
nand U5189 (N_5189,N_4807,N_4911);
and U5190 (N_5190,N_4982,N_4931);
nand U5191 (N_5191,N_4887,N_4948);
or U5192 (N_5192,N_4876,N_4841);
nand U5193 (N_5193,N_4922,N_4800);
nand U5194 (N_5194,N_4971,N_4961);
xnor U5195 (N_5195,N_4854,N_4861);
xor U5196 (N_5196,N_4851,N_4825);
nor U5197 (N_5197,N_4819,N_4874);
xor U5198 (N_5198,N_4846,N_4822);
nand U5199 (N_5199,N_4989,N_4948);
xor U5200 (N_5200,N_5089,N_5195);
or U5201 (N_5201,N_5051,N_5039);
nor U5202 (N_5202,N_5119,N_5109);
nand U5203 (N_5203,N_5099,N_5002);
and U5204 (N_5204,N_5163,N_5075);
or U5205 (N_5205,N_5032,N_5025);
nand U5206 (N_5206,N_5033,N_5056);
and U5207 (N_5207,N_5014,N_5031);
and U5208 (N_5208,N_5132,N_5057);
or U5209 (N_5209,N_5147,N_5084);
and U5210 (N_5210,N_5193,N_5097);
and U5211 (N_5211,N_5146,N_5116);
nand U5212 (N_5212,N_5092,N_5093);
xor U5213 (N_5213,N_5111,N_5198);
xnor U5214 (N_5214,N_5159,N_5066);
and U5215 (N_5215,N_5169,N_5192);
and U5216 (N_5216,N_5167,N_5096);
nand U5217 (N_5217,N_5076,N_5113);
nand U5218 (N_5218,N_5182,N_5095);
nand U5219 (N_5219,N_5052,N_5110);
xor U5220 (N_5220,N_5134,N_5070);
nor U5221 (N_5221,N_5187,N_5024);
nand U5222 (N_5222,N_5157,N_5004);
and U5223 (N_5223,N_5180,N_5103);
or U5224 (N_5224,N_5101,N_5141);
xor U5225 (N_5225,N_5068,N_5127);
xor U5226 (N_5226,N_5078,N_5177);
xor U5227 (N_5227,N_5139,N_5009);
or U5228 (N_5228,N_5011,N_5108);
or U5229 (N_5229,N_5144,N_5044);
and U5230 (N_5230,N_5081,N_5067);
nor U5231 (N_5231,N_5140,N_5152);
or U5232 (N_5232,N_5080,N_5054);
nor U5233 (N_5233,N_5120,N_5038);
nand U5234 (N_5234,N_5016,N_5199);
and U5235 (N_5235,N_5077,N_5050);
or U5236 (N_5236,N_5015,N_5189);
xnor U5237 (N_5237,N_5150,N_5118);
or U5238 (N_5238,N_5171,N_5100);
and U5239 (N_5239,N_5007,N_5043);
or U5240 (N_5240,N_5073,N_5188);
or U5241 (N_5241,N_5164,N_5129);
and U5242 (N_5242,N_5185,N_5102);
nand U5243 (N_5243,N_5172,N_5020);
xor U5244 (N_5244,N_5161,N_5123);
nor U5245 (N_5245,N_5088,N_5142);
xnor U5246 (N_5246,N_5065,N_5005);
and U5247 (N_5247,N_5155,N_5055);
xnor U5248 (N_5248,N_5196,N_5174);
or U5249 (N_5249,N_5178,N_5106);
nand U5250 (N_5250,N_5160,N_5154);
or U5251 (N_5251,N_5197,N_5026);
and U5252 (N_5252,N_5045,N_5069);
nor U5253 (N_5253,N_5194,N_5037);
xor U5254 (N_5254,N_5156,N_5184);
and U5255 (N_5255,N_5071,N_5115);
or U5256 (N_5256,N_5166,N_5013);
and U5257 (N_5257,N_5105,N_5162);
and U5258 (N_5258,N_5074,N_5165);
or U5259 (N_5259,N_5030,N_5090);
nor U5260 (N_5260,N_5112,N_5006);
nand U5261 (N_5261,N_5186,N_5125);
nand U5262 (N_5262,N_5191,N_5021);
nand U5263 (N_5263,N_5094,N_5135);
nor U5264 (N_5264,N_5079,N_5183);
nand U5265 (N_5265,N_5131,N_5104);
or U5266 (N_5266,N_5136,N_5022);
or U5267 (N_5267,N_5017,N_5107);
and U5268 (N_5268,N_5048,N_5176);
or U5269 (N_5269,N_5148,N_5042);
xnor U5270 (N_5270,N_5060,N_5058);
nand U5271 (N_5271,N_5029,N_5190);
or U5272 (N_5272,N_5168,N_5072);
and U5273 (N_5273,N_5010,N_5046);
and U5274 (N_5274,N_5098,N_5061);
nand U5275 (N_5275,N_5018,N_5138);
xnor U5276 (N_5276,N_5003,N_5179);
and U5277 (N_5277,N_5158,N_5137);
nor U5278 (N_5278,N_5000,N_5181);
nand U5279 (N_5279,N_5064,N_5151);
and U5280 (N_5280,N_5083,N_5114);
or U5281 (N_5281,N_5041,N_5028);
nor U5282 (N_5282,N_5133,N_5059);
or U5283 (N_5283,N_5036,N_5082);
nand U5284 (N_5284,N_5173,N_5170);
or U5285 (N_5285,N_5040,N_5047);
or U5286 (N_5286,N_5035,N_5086);
nor U5287 (N_5287,N_5012,N_5001);
nor U5288 (N_5288,N_5145,N_5053);
nand U5289 (N_5289,N_5049,N_5034);
nor U5290 (N_5290,N_5085,N_5019);
and U5291 (N_5291,N_5117,N_5124);
xnor U5292 (N_5292,N_5153,N_5149);
xor U5293 (N_5293,N_5063,N_5008);
nand U5294 (N_5294,N_5062,N_5128);
or U5295 (N_5295,N_5027,N_5122);
and U5296 (N_5296,N_5175,N_5143);
nand U5297 (N_5297,N_5091,N_5023);
and U5298 (N_5298,N_5126,N_5121);
xnor U5299 (N_5299,N_5130,N_5087);
and U5300 (N_5300,N_5039,N_5101);
and U5301 (N_5301,N_5143,N_5073);
nor U5302 (N_5302,N_5039,N_5002);
nor U5303 (N_5303,N_5087,N_5044);
xor U5304 (N_5304,N_5160,N_5018);
or U5305 (N_5305,N_5196,N_5140);
xor U5306 (N_5306,N_5126,N_5178);
nand U5307 (N_5307,N_5020,N_5098);
or U5308 (N_5308,N_5171,N_5073);
and U5309 (N_5309,N_5086,N_5198);
xor U5310 (N_5310,N_5180,N_5126);
nand U5311 (N_5311,N_5116,N_5045);
or U5312 (N_5312,N_5113,N_5107);
and U5313 (N_5313,N_5152,N_5172);
nand U5314 (N_5314,N_5025,N_5144);
and U5315 (N_5315,N_5133,N_5017);
xor U5316 (N_5316,N_5012,N_5000);
nor U5317 (N_5317,N_5112,N_5167);
and U5318 (N_5318,N_5163,N_5143);
xnor U5319 (N_5319,N_5184,N_5043);
or U5320 (N_5320,N_5017,N_5159);
and U5321 (N_5321,N_5023,N_5064);
nand U5322 (N_5322,N_5008,N_5073);
nor U5323 (N_5323,N_5001,N_5152);
nand U5324 (N_5324,N_5177,N_5002);
xor U5325 (N_5325,N_5184,N_5122);
nor U5326 (N_5326,N_5132,N_5148);
or U5327 (N_5327,N_5179,N_5000);
and U5328 (N_5328,N_5118,N_5124);
nand U5329 (N_5329,N_5005,N_5082);
nor U5330 (N_5330,N_5110,N_5089);
nor U5331 (N_5331,N_5063,N_5068);
and U5332 (N_5332,N_5147,N_5030);
and U5333 (N_5333,N_5163,N_5127);
nand U5334 (N_5334,N_5147,N_5102);
nand U5335 (N_5335,N_5093,N_5191);
xnor U5336 (N_5336,N_5146,N_5111);
xnor U5337 (N_5337,N_5080,N_5183);
xor U5338 (N_5338,N_5058,N_5054);
nand U5339 (N_5339,N_5023,N_5038);
xnor U5340 (N_5340,N_5063,N_5012);
nand U5341 (N_5341,N_5080,N_5171);
xor U5342 (N_5342,N_5184,N_5196);
xor U5343 (N_5343,N_5048,N_5164);
or U5344 (N_5344,N_5040,N_5182);
xor U5345 (N_5345,N_5157,N_5028);
nand U5346 (N_5346,N_5026,N_5013);
and U5347 (N_5347,N_5102,N_5152);
nand U5348 (N_5348,N_5043,N_5029);
xor U5349 (N_5349,N_5169,N_5052);
nand U5350 (N_5350,N_5198,N_5109);
nand U5351 (N_5351,N_5177,N_5058);
nor U5352 (N_5352,N_5122,N_5035);
and U5353 (N_5353,N_5159,N_5045);
nor U5354 (N_5354,N_5015,N_5009);
and U5355 (N_5355,N_5112,N_5081);
or U5356 (N_5356,N_5078,N_5035);
nand U5357 (N_5357,N_5135,N_5014);
nor U5358 (N_5358,N_5156,N_5100);
xor U5359 (N_5359,N_5060,N_5050);
xor U5360 (N_5360,N_5090,N_5017);
nor U5361 (N_5361,N_5188,N_5032);
nand U5362 (N_5362,N_5110,N_5072);
and U5363 (N_5363,N_5061,N_5066);
nor U5364 (N_5364,N_5188,N_5119);
xnor U5365 (N_5365,N_5159,N_5172);
nand U5366 (N_5366,N_5001,N_5149);
nand U5367 (N_5367,N_5128,N_5046);
or U5368 (N_5368,N_5146,N_5035);
or U5369 (N_5369,N_5098,N_5114);
nand U5370 (N_5370,N_5029,N_5191);
xnor U5371 (N_5371,N_5169,N_5101);
nor U5372 (N_5372,N_5143,N_5070);
and U5373 (N_5373,N_5106,N_5175);
xnor U5374 (N_5374,N_5128,N_5095);
or U5375 (N_5375,N_5092,N_5066);
xor U5376 (N_5376,N_5170,N_5039);
nor U5377 (N_5377,N_5166,N_5045);
and U5378 (N_5378,N_5033,N_5064);
or U5379 (N_5379,N_5123,N_5163);
nand U5380 (N_5380,N_5060,N_5155);
nand U5381 (N_5381,N_5169,N_5050);
nor U5382 (N_5382,N_5112,N_5169);
xor U5383 (N_5383,N_5128,N_5189);
and U5384 (N_5384,N_5094,N_5063);
and U5385 (N_5385,N_5124,N_5137);
nand U5386 (N_5386,N_5030,N_5131);
nor U5387 (N_5387,N_5132,N_5077);
and U5388 (N_5388,N_5033,N_5155);
nor U5389 (N_5389,N_5002,N_5194);
or U5390 (N_5390,N_5102,N_5170);
nand U5391 (N_5391,N_5059,N_5015);
nand U5392 (N_5392,N_5138,N_5188);
xor U5393 (N_5393,N_5143,N_5047);
nand U5394 (N_5394,N_5014,N_5002);
nor U5395 (N_5395,N_5169,N_5095);
xnor U5396 (N_5396,N_5010,N_5186);
and U5397 (N_5397,N_5126,N_5140);
nand U5398 (N_5398,N_5073,N_5009);
nand U5399 (N_5399,N_5124,N_5086);
nand U5400 (N_5400,N_5329,N_5243);
xor U5401 (N_5401,N_5246,N_5396);
nor U5402 (N_5402,N_5267,N_5251);
nor U5403 (N_5403,N_5372,N_5303);
xnor U5404 (N_5404,N_5290,N_5315);
nand U5405 (N_5405,N_5257,N_5256);
nand U5406 (N_5406,N_5254,N_5284);
nand U5407 (N_5407,N_5362,N_5203);
nand U5408 (N_5408,N_5331,N_5278);
and U5409 (N_5409,N_5320,N_5347);
or U5410 (N_5410,N_5299,N_5212);
xor U5411 (N_5411,N_5272,N_5361);
or U5412 (N_5412,N_5206,N_5217);
and U5413 (N_5413,N_5306,N_5348);
xor U5414 (N_5414,N_5374,N_5244);
nand U5415 (N_5415,N_5264,N_5281);
xor U5416 (N_5416,N_5317,N_5345);
nor U5417 (N_5417,N_5273,N_5210);
or U5418 (N_5418,N_5357,N_5369);
or U5419 (N_5419,N_5350,N_5380);
nand U5420 (N_5420,N_5352,N_5245);
nor U5421 (N_5421,N_5226,N_5346);
or U5422 (N_5422,N_5259,N_5287);
or U5423 (N_5423,N_5309,N_5354);
nor U5424 (N_5424,N_5343,N_5231);
and U5425 (N_5425,N_5392,N_5397);
xor U5426 (N_5426,N_5227,N_5393);
and U5427 (N_5427,N_5219,N_5384);
and U5428 (N_5428,N_5330,N_5216);
or U5429 (N_5429,N_5253,N_5266);
nor U5430 (N_5430,N_5292,N_5319);
xor U5431 (N_5431,N_5230,N_5201);
or U5432 (N_5432,N_5218,N_5356);
nor U5433 (N_5433,N_5252,N_5239);
nor U5434 (N_5434,N_5242,N_5341);
nor U5435 (N_5435,N_5235,N_5258);
xor U5436 (N_5436,N_5214,N_5205);
nor U5437 (N_5437,N_5285,N_5291);
nor U5438 (N_5438,N_5234,N_5316);
xor U5439 (N_5439,N_5351,N_5282);
or U5440 (N_5440,N_5237,N_5376);
xor U5441 (N_5441,N_5274,N_5333);
and U5442 (N_5442,N_5387,N_5289);
or U5443 (N_5443,N_5334,N_5233);
nand U5444 (N_5444,N_5308,N_5338);
and U5445 (N_5445,N_5304,N_5342);
and U5446 (N_5446,N_5224,N_5359);
nand U5447 (N_5447,N_5337,N_5377);
xor U5448 (N_5448,N_5204,N_5339);
or U5449 (N_5449,N_5215,N_5307);
nand U5450 (N_5450,N_5335,N_5247);
nor U5451 (N_5451,N_5365,N_5325);
and U5452 (N_5452,N_5298,N_5379);
nand U5453 (N_5453,N_5232,N_5209);
nor U5454 (N_5454,N_5288,N_5375);
and U5455 (N_5455,N_5248,N_5225);
xor U5456 (N_5456,N_5395,N_5312);
or U5457 (N_5457,N_5213,N_5263);
nand U5458 (N_5458,N_5321,N_5344);
and U5459 (N_5459,N_5240,N_5295);
xor U5460 (N_5460,N_5367,N_5336);
nor U5461 (N_5461,N_5260,N_5378);
and U5462 (N_5462,N_5360,N_5318);
nand U5463 (N_5463,N_5301,N_5355);
nor U5464 (N_5464,N_5200,N_5328);
or U5465 (N_5465,N_5271,N_5277);
and U5466 (N_5466,N_5324,N_5388);
xnor U5467 (N_5467,N_5364,N_5279);
xnor U5468 (N_5468,N_5368,N_5383);
xor U5469 (N_5469,N_5283,N_5373);
nor U5470 (N_5470,N_5314,N_5391);
xor U5471 (N_5471,N_5386,N_5313);
nand U5472 (N_5472,N_5323,N_5382);
and U5473 (N_5473,N_5269,N_5221);
nor U5474 (N_5474,N_5322,N_5332);
nor U5475 (N_5475,N_5394,N_5363);
or U5476 (N_5476,N_5202,N_5340);
nand U5477 (N_5477,N_5265,N_5236);
xor U5478 (N_5478,N_5276,N_5370);
or U5479 (N_5479,N_5229,N_5327);
or U5480 (N_5480,N_5261,N_5249);
nor U5481 (N_5481,N_5385,N_5223);
nor U5482 (N_5482,N_5353,N_5228);
nand U5483 (N_5483,N_5297,N_5311);
nor U5484 (N_5484,N_5305,N_5207);
xnor U5485 (N_5485,N_5366,N_5241);
and U5486 (N_5486,N_5296,N_5371);
xnor U5487 (N_5487,N_5280,N_5390);
and U5488 (N_5488,N_5220,N_5208);
nand U5489 (N_5489,N_5222,N_5250);
or U5490 (N_5490,N_5255,N_5294);
nor U5491 (N_5491,N_5310,N_5286);
and U5492 (N_5492,N_5268,N_5389);
and U5493 (N_5493,N_5300,N_5211);
nand U5494 (N_5494,N_5275,N_5238);
nor U5495 (N_5495,N_5270,N_5349);
nor U5496 (N_5496,N_5398,N_5293);
nor U5497 (N_5497,N_5326,N_5358);
nor U5498 (N_5498,N_5381,N_5262);
nor U5499 (N_5499,N_5399,N_5302);
and U5500 (N_5500,N_5305,N_5283);
and U5501 (N_5501,N_5234,N_5305);
and U5502 (N_5502,N_5344,N_5342);
nand U5503 (N_5503,N_5385,N_5209);
xor U5504 (N_5504,N_5376,N_5377);
and U5505 (N_5505,N_5377,N_5219);
nor U5506 (N_5506,N_5378,N_5216);
nand U5507 (N_5507,N_5333,N_5247);
and U5508 (N_5508,N_5211,N_5356);
nand U5509 (N_5509,N_5283,N_5279);
and U5510 (N_5510,N_5312,N_5227);
or U5511 (N_5511,N_5234,N_5378);
and U5512 (N_5512,N_5348,N_5233);
or U5513 (N_5513,N_5303,N_5311);
nor U5514 (N_5514,N_5207,N_5365);
and U5515 (N_5515,N_5395,N_5335);
xnor U5516 (N_5516,N_5383,N_5205);
xnor U5517 (N_5517,N_5298,N_5234);
xor U5518 (N_5518,N_5394,N_5278);
xor U5519 (N_5519,N_5283,N_5246);
nand U5520 (N_5520,N_5281,N_5300);
or U5521 (N_5521,N_5391,N_5341);
nor U5522 (N_5522,N_5377,N_5293);
nand U5523 (N_5523,N_5380,N_5246);
and U5524 (N_5524,N_5356,N_5399);
and U5525 (N_5525,N_5371,N_5282);
nand U5526 (N_5526,N_5267,N_5327);
and U5527 (N_5527,N_5343,N_5331);
or U5528 (N_5528,N_5211,N_5354);
or U5529 (N_5529,N_5315,N_5397);
or U5530 (N_5530,N_5388,N_5237);
nor U5531 (N_5531,N_5259,N_5206);
or U5532 (N_5532,N_5361,N_5344);
nand U5533 (N_5533,N_5332,N_5283);
nor U5534 (N_5534,N_5319,N_5318);
xnor U5535 (N_5535,N_5369,N_5332);
xor U5536 (N_5536,N_5297,N_5385);
nand U5537 (N_5537,N_5214,N_5392);
nor U5538 (N_5538,N_5372,N_5219);
or U5539 (N_5539,N_5265,N_5250);
or U5540 (N_5540,N_5351,N_5239);
and U5541 (N_5541,N_5339,N_5322);
or U5542 (N_5542,N_5208,N_5224);
or U5543 (N_5543,N_5308,N_5378);
nand U5544 (N_5544,N_5222,N_5288);
xnor U5545 (N_5545,N_5395,N_5393);
xor U5546 (N_5546,N_5328,N_5235);
nand U5547 (N_5547,N_5300,N_5222);
or U5548 (N_5548,N_5335,N_5380);
xor U5549 (N_5549,N_5223,N_5251);
or U5550 (N_5550,N_5209,N_5308);
nand U5551 (N_5551,N_5204,N_5284);
and U5552 (N_5552,N_5374,N_5216);
and U5553 (N_5553,N_5218,N_5267);
and U5554 (N_5554,N_5306,N_5304);
and U5555 (N_5555,N_5329,N_5291);
xor U5556 (N_5556,N_5273,N_5346);
or U5557 (N_5557,N_5230,N_5316);
nor U5558 (N_5558,N_5383,N_5255);
nor U5559 (N_5559,N_5208,N_5338);
or U5560 (N_5560,N_5317,N_5289);
nor U5561 (N_5561,N_5310,N_5248);
and U5562 (N_5562,N_5203,N_5271);
xnor U5563 (N_5563,N_5331,N_5313);
nor U5564 (N_5564,N_5284,N_5378);
and U5565 (N_5565,N_5224,N_5331);
nor U5566 (N_5566,N_5350,N_5249);
nand U5567 (N_5567,N_5201,N_5284);
nand U5568 (N_5568,N_5203,N_5352);
and U5569 (N_5569,N_5322,N_5214);
nor U5570 (N_5570,N_5263,N_5279);
nand U5571 (N_5571,N_5323,N_5259);
nor U5572 (N_5572,N_5330,N_5242);
xor U5573 (N_5573,N_5392,N_5323);
xor U5574 (N_5574,N_5277,N_5273);
xor U5575 (N_5575,N_5235,N_5294);
and U5576 (N_5576,N_5329,N_5206);
nor U5577 (N_5577,N_5246,N_5244);
nand U5578 (N_5578,N_5350,N_5371);
xor U5579 (N_5579,N_5219,N_5255);
and U5580 (N_5580,N_5278,N_5322);
nand U5581 (N_5581,N_5327,N_5370);
nand U5582 (N_5582,N_5334,N_5208);
nor U5583 (N_5583,N_5374,N_5220);
xnor U5584 (N_5584,N_5318,N_5251);
or U5585 (N_5585,N_5293,N_5301);
or U5586 (N_5586,N_5352,N_5207);
nand U5587 (N_5587,N_5249,N_5304);
nand U5588 (N_5588,N_5269,N_5351);
or U5589 (N_5589,N_5331,N_5238);
nor U5590 (N_5590,N_5397,N_5391);
and U5591 (N_5591,N_5289,N_5260);
and U5592 (N_5592,N_5233,N_5264);
and U5593 (N_5593,N_5367,N_5208);
xor U5594 (N_5594,N_5328,N_5275);
nand U5595 (N_5595,N_5213,N_5377);
or U5596 (N_5596,N_5233,N_5265);
nand U5597 (N_5597,N_5333,N_5272);
or U5598 (N_5598,N_5227,N_5371);
or U5599 (N_5599,N_5338,N_5287);
xor U5600 (N_5600,N_5596,N_5494);
nand U5601 (N_5601,N_5584,N_5525);
or U5602 (N_5602,N_5522,N_5472);
nand U5603 (N_5603,N_5561,N_5559);
xnor U5604 (N_5604,N_5565,N_5538);
or U5605 (N_5605,N_5488,N_5449);
nand U5606 (N_5606,N_5463,N_5482);
nand U5607 (N_5607,N_5420,N_5465);
nand U5608 (N_5608,N_5597,N_5572);
nand U5609 (N_5609,N_5564,N_5544);
nand U5610 (N_5610,N_5513,N_5576);
xnor U5611 (N_5611,N_5400,N_5578);
and U5612 (N_5612,N_5523,N_5454);
xor U5613 (N_5613,N_5451,N_5466);
xor U5614 (N_5614,N_5432,N_5534);
or U5615 (N_5615,N_5441,N_5456);
nand U5616 (N_5616,N_5434,N_5548);
xor U5617 (N_5617,N_5598,N_5536);
xor U5618 (N_5618,N_5521,N_5438);
and U5619 (N_5619,N_5563,N_5497);
xnor U5620 (N_5620,N_5457,N_5545);
xor U5621 (N_5621,N_5413,N_5433);
nand U5622 (N_5622,N_5590,N_5549);
or U5623 (N_5623,N_5539,N_5542);
xor U5624 (N_5624,N_5450,N_5473);
and U5625 (N_5625,N_5593,N_5510);
xnor U5626 (N_5626,N_5547,N_5444);
xnor U5627 (N_5627,N_5502,N_5503);
or U5628 (N_5628,N_5531,N_5505);
nor U5629 (N_5629,N_5574,N_5546);
and U5630 (N_5630,N_5486,N_5589);
and U5631 (N_5631,N_5526,N_5557);
xnor U5632 (N_5632,N_5512,N_5582);
nand U5633 (N_5633,N_5422,N_5567);
xor U5634 (N_5634,N_5493,N_5445);
and U5635 (N_5635,N_5550,N_5571);
nand U5636 (N_5636,N_5515,N_5417);
nor U5637 (N_5637,N_5517,N_5479);
nand U5638 (N_5638,N_5411,N_5415);
nand U5639 (N_5639,N_5579,N_5528);
and U5640 (N_5640,N_5460,N_5423);
nor U5641 (N_5641,N_5407,N_5462);
nand U5642 (N_5642,N_5431,N_5455);
nor U5643 (N_5643,N_5474,N_5524);
and U5644 (N_5644,N_5595,N_5496);
and U5645 (N_5645,N_5527,N_5405);
nand U5646 (N_5646,N_5583,N_5554);
or U5647 (N_5647,N_5558,N_5489);
xor U5648 (N_5648,N_5537,N_5458);
nor U5649 (N_5649,N_5436,N_5587);
nand U5650 (N_5650,N_5467,N_5425);
nor U5651 (N_5651,N_5498,N_5448);
nor U5652 (N_5652,N_5439,N_5483);
or U5653 (N_5653,N_5470,N_5430);
nand U5654 (N_5654,N_5453,N_5581);
xor U5655 (N_5655,N_5573,N_5452);
and U5656 (N_5656,N_5532,N_5553);
or U5657 (N_5657,N_5428,N_5530);
and U5658 (N_5658,N_5508,N_5469);
or U5659 (N_5659,N_5492,N_5447);
xnor U5660 (N_5660,N_5588,N_5477);
nand U5661 (N_5661,N_5418,N_5491);
nor U5662 (N_5662,N_5519,N_5426);
and U5663 (N_5663,N_5437,N_5419);
and U5664 (N_5664,N_5499,N_5461);
nand U5665 (N_5665,N_5484,N_5520);
nor U5666 (N_5666,N_5516,N_5446);
or U5667 (N_5667,N_5468,N_5506);
nor U5668 (N_5668,N_5464,N_5481);
xor U5669 (N_5669,N_5569,N_5408);
or U5670 (N_5670,N_5504,N_5487);
nor U5671 (N_5671,N_5560,N_5566);
and U5672 (N_5672,N_5443,N_5476);
nand U5673 (N_5673,N_5551,N_5570);
nand U5674 (N_5674,N_5577,N_5592);
xnor U5675 (N_5675,N_5495,N_5403);
nor U5676 (N_5676,N_5540,N_5594);
nor U5677 (N_5677,N_5401,N_5591);
nand U5678 (N_5678,N_5555,N_5406);
nand U5679 (N_5679,N_5529,N_5518);
or U5680 (N_5680,N_5424,N_5404);
xor U5681 (N_5681,N_5599,N_5440);
nor U5682 (N_5682,N_5427,N_5478);
xnor U5683 (N_5683,N_5507,N_5414);
or U5684 (N_5684,N_5533,N_5575);
xor U5685 (N_5685,N_5442,N_5500);
nand U5686 (N_5686,N_5562,N_5421);
nand U5687 (N_5687,N_5552,N_5543);
nor U5688 (N_5688,N_5514,N_5416);
and U5689 (N_5689,N_5568,N_5535);
or U5690 (N_5690,N_5471,N_5429);
nand U5691 (N_5691,N_5480,N_5501);
and U5692 (N_5692,N_5475,N_5586);
and U5693 (N_5693,N_5409,N_5485);
and U5694 (N_5694,N_5541,N_5459);
and U5695 (N_5695,N_5511,N_5435);
nor U5696 (N_5696,N_5556,N_5402);
nor U5697 (N_5697,N_5585,N_5412);
nor U5698 (N_5698,N_5490,N_5410);
and U5699 (N_5699,N_5580,N_5509);
nand U5700 (N_5700,N_5439,N_5426);
xor U5701 (N_5701,N_5485,N_5569);
xor U5702 (N_5702,N_5575,N_5453);
nand U5703 (N_5703,N_5572,N_5411);
nand U5704 (N_5704,N_5549,N_5543);
nand U5705 (N_5705,N_5499,N_5501);
or U5706 (N_5706,N_5414,N_5532);
xor U5707 (N_5707,N_5438,N_5454);
and U5708 (N_5708,N_5541,N_5585);
and U5709 (N_5709,N_5443,N_5558);
nor U5710 (N_5710,N_5590,N_5430);
and U5711 (N_5711,N_5570,N_5568);
nand U5712 (N_5712,N_5465,N_5502);
xnor U5713 (N_5713,N_5485,N_5598);
nand U5714 (N_5714,N_5444,N_5520);
xnor U5715 (N_5715,N_5449,N_5505);
nor U5716 (N_5716,N_5568,N_5431);
or U5717 (N_5717,N_5477,N_5531);
or U5718 (N_5718,N_5564,N_5437);
and U5719 (N_5719,N_5553,N_5559);
xor U5720 (N_5720,N_5493,N_5500);
nand U5721 (N_5721,N_5420,N_5433);
and U5722 (N_5722,N_5412,N_5508);
nand U5723 (N_5723,N_5541,N_5429);
or U5724 (N_5724,N_5464,N_5492);
nor U5725 (N_5725,N_5466,N_5544);
xor U5726 (N_5726,N_5451,N_5462);
nand U5727 (N_5727,N_5534,N_5478);
xnor U5728 (N_5728,N_5474,N_5559);
nor U5729 (N_5729,N_5458,N_5529);
nand U5730 (N_5730,N_5422,N_5544);
and U5731 (N_5731,N_5449,N_5461);
and U5732 (N_5732,N_5463,N_5429);
nor U5733 (N_5733,N_5423,N_5546);
or U5734 (N_5734,N_5554,N_5512);
nand U5735 (N_5735,N_5571,N_5486);
nor U5736 (N_5736,N_5598,N_5427);
and U5737 (N_5737,N_5420,N_5498);
and U5738 (N_5738,N_5581,N_5403);
nand U5739 (N_5739,N_5596,N_5570);
xor U5740 (N_5740,N_5456,N_5516);
or U5741 (N_5741,N_5502,N_5559);
xor U5742 (N_5742,N_5551,N_5505);
or U5743 (N_5743,N_5514,N_5597);
nand U5744 (N_5744,N_5498,N_5432);
nor U5745 (N_5745,N_5593,N_5442);
or U5746 (N_5746,N_5406,N_5419);
or U5747 (N_5747,N_5435,N_5481);
and U5748 (N_5748,N_5424,N_5595);
nand U5749 (N_5749,N_5457,N_5535);
nor U5750 (N_5750,N_5479,N_5529);
nor U5751 (N_5751,N_5591,N_5534);
xnor U5752 (N_5752,N_5563,N_5532);
nor U5753 (N_5753,N_5495,N_5446);
xor U5754 (N_5754,N_5536,N_5400);
xor U5755 (N_5755,N_5493,N_5590);
and U5756 (N_5756,N_5589,N_5507);
or U5757 (N_5757,N_5413,N_5594);
nand U5758 (N_5758,N_5568,N_5527);
nor U5759 (N_5759,N_5471,N_5587);
nor U5760 (N_5760,N_5580,N_5568);
nand U5761 (N_5761,N_5505,N_5578);
xnor U5762 (N_5762,N_5451,N_5537);
xnor U5763 (N_5763,N_5498,N_5419);
and U5764 (N_5764,N_5566,N_5402);
nor U5765 (N_5765,N_5478,N_5506);
or U5766 (N_5766,N_5542,N_5516);
nand U5767 (N_5767,N_5449,N_5586);
and U5768 (N_5768,N_5512,N_5499);
xor U5769 (N_5769,N_5446,N_5417);
and U5770 (N_5770,N_5412,N_5545);
and U5771 (N_5771,N_5591,N_5537);
xnor U5772 (N_5772,N_5547,N_5542);
nand U5773 (N_5773,N_5510,N_5414);
and U5774 (N_5774,N_5494,N_5476);
or U5775 (N_5775,N_5446,N_5527);
xnor U5776 (N_5776,N_5479,N_5485);
and U5777 (N_5777,N_5480,N_5496);
and U5778 (N_5778,N_5596,N_5527);
nand U5779 (N_5779,N_5471,N_5561);
or U5780 (N_5780,N_5470,N_5462);
xor U5781 (N_5781,N_5544,N_5537);
and U5782 (N_5782,N_5592,N_5421);
or U5783 (N_5783,N_5542,N_5412);
and U5784 (N_5784,N_5497,N_5489);
or U5785 (N_5785,N_5546,N_5590);
xnor U5786 (N_5786,N_5501,N_5536);
nor U5787 (N_5787,N_5405,N_5449);
xnor U5788 (N_5788,N_5581,N_5438);
xor U5789 (N_5789,N_5432,N_5417);
nand U5790 (N_5790,N_5420,N_5432);
nor U5791 (N_5791,N_5514,N_5463);
or U5792 (N_5792,N_5483,N_5570);
nor U5793 (N_5793,N_5432,N_5512);
or U5794 (N_5794,N_5532,N_5484);
nor U5795 (N_5795,N_5460,N_5527);
nor U5796 (N_5796,N_5588,N_5432);
nand U5797 (N_5797,N_5483,N_5487);
nor U5798 (N_5798,N_5414,N_5503);
nor U5799 (N_5799,N_5420,N_5533);
and U5800 (N_5800,N_5793,N_5683);
nand U5801 (N_5801,N_5764,N_5750);
nand U5802 (N_5802,N_5763,N_5719);
and U5803 (N_5803,N_5725,N_5731);
xor U5804 (N_5804,N_5738,N_5672);
and U5805 (N_5805,N_5762,N_5674);
nor U5806 (N_5806,N_5675,N_5688);
xnor U5807 (N_5807,N_5723,N_5693);
nand U5808 (N_5808,N_5716,N_5780);
or U5809 (N_5809,N_5798,N_5709);
and U5810 (N_5810,N_5778,N_5757);
or U5811 (N_5811,N_5603,N_5734);
or U5812 (N_5812,N_5752,N_5666);
nor U5813 (N_5813,N_5681,N_5652);
nand U5814 (N_5814,N_5664,N_5728);
xnor U5815 (N_5815,N_5729,N_5651);
or U5816 (N_5816,N_5690,N_5673);
xor U5817 (N_5817,N_5724,N_5604);
or U5818 (N_5818,N_5749,N_5602);
nand U5819 (N_5819,N_5637,N_5670);
or U5820 (N_5820,N_5617,N_5715);
or U5821 (N_5821,N_5711,N_5665);
or U5822 (N_5822,N_5772,N_5643);
or U5823 (N_5823,N_5792,N_5649);
nand U5824 (N_5824,N_5741,N_5684);
nor U5825 (N_5825,N_5620,N_5691);
nand U5826 (N_5826,N_5783,N_5625);
and U5827 (N_5827,N_5735,N_5739);
nand U5828 (N_5828,N_5694,N_5708);
and U5829 (N_5829,N_5775,N_5621);
and U5830 (N_5830,N_5767,N_5689);
and U5831 (N_5831,N_5636,N_5782);
or U5832 (N_5832,N_5785,N_5787);
and U5833 (N_5833,N_5795,N_5663);
or U5834 (N_5834,N_5722,N_5732);
and U5835 (N_5835,N_5700,N_5765);
xnor U5836 (N_5836,N_5650,N_5642);
nor U5837 (N_5837,N_5677,N_5610);
or U5838 (N_5838,N_5756,N_5622);
and U5839 (N_5839,N_5769,N_5768);
and U5840 (N_5840,N_5737,N_5605);
or U5841 (N_5841,N_5705,N_5601);
nand U5842 (N_5842,N_5744,N_5669);
nand U5843 (N_5843,N_5755,N_5624);
xor U5844 (N_5844,N_5773,N_5678);
xnor U5845 (N_5845,N_5745,N_5698);
nand U5846 (N_5846,N_5632,N_5779);
or U5847 (N_5847,N_5611,N_5799);
xnor U5848 (N_5848,N_5613,N_5760);
xnor U5849 (N_5849,N_5609,N_5746);
and U5850 (N_5850,N_5742,N_5692);
and U5851 (N_5851,N_5781,N_5615);
and U5852 (N_5852,N_5623,N_5655);
nand U5853 (N_5853,N_5616,N_5704);
nor U5854 (N_5854,N_5702,N_5656);
and U5855 (N_5855,N_5612,N_5628);
or U5856 (N_5856,N_5777,N_5796);
nand U5857 (N_5857,N_5730,N_5696);
xnor U5858 (N_5858,N_5639,N_5659);
or U5859 (N_5859,N_5784,N_5627);
or U5860 (N_5860,N_5759,N_5654);
and U5861 (N_5861,N_5638,N_5667);
nor U5862 (N_5862,N_5606,N_5747);
nand U5863 (N_5863,N_5758,N_5647);
and U5864 (N_5864,N_5706,N_5736);
and U5865 (N_5865,N_5646,N_5657);
and U5866 (N_5866,N_5774,N_5600);
nand U5867 (N_5867,N_5653,N_5680);
xor U5868 (N_5868,N_5714,N_5713);
nor U5869 (N_5869,N_5771,N_5712);
and U5870 (N_5870,N_5607,N_5676);
and U5871 (N_5871,N_5721,N_5633);
nor U5872 (N_5872,N_5645,N_5644);
and U5873 (N_5873,N_5770,N_5641);
nand U5874 (N_5874,N_5751,N_5658);
or U5875 (N_5875,N_5686,N_5640);
xor U5876 (N_5876,N_5614,N_5662);
or U5877 (N_5877,N_5766,N_5697);
nor U5878 (N_5878,N_5797,N_5733);
and U5879 (N_5879,N_5740,N_5743);
nor U5880 (N_5880,N_5786,N_5695);
or U5881 (N_5881,N_5791,N_5608);
or U5882 (N_5882,N_5776,N_5753);
nand U5883 (N_5883,N_5629,N_5619);
and U5884 (N_5884,N_5754,N_5788);
or U5885 (N_5885,N_5790,N_5661);
and U5886 (N_5886,N_5685,N_5727);
nand U5887 (N_5887,N_5789,N_5630);
xnor U5888 (N_5888,N_5761,N_5794);
nand U5889 (N_5889,N_5726,N_5748);
and U5890 (N_5890,N_5699,N_5710);
nor U5891 (N_5891,N_5717,N_5648);
xor U5892 (N_5892,N_5660,N_5679);
and U5893 (N_5893,N_5720,N_5626);
nor U5894 (N_5894,N_5671,N_5631);
nor U5895 (N_5895,N_5635,N_5701);
nand U5896 (N_5896,N_5668,N_5618);
and U5897 (N_5897,N_5687,N_5703);
or U5898 (N_5898,N_5718,N_5634);
and U5899 (N_5899,N_5707,N_5682);
nor U5900 (N_5900,N_5761,N_5726);
xnor U5901 (N_5901,N_5631,N_5724);
xnor U5902 (N_5902,N_5743,N_5764);
nand U5903 (N_5903,N_5682,N_5646);
nand U5904 (N_5904,N_5634,N_5702);
nor U5905 (N_5905,N_5662,N_5789);
nor U5906 (N_5906,N_5629,N_5753);
nor U5907 (N_5907,N_5641,N_5745);
or U5908 (N_5908,N_5672,N_5754);
nand U5909 (N_5909,N_5752,N_5709);
and U5910 (N_5910,N_5658,N_5737);
or U5911 (N_5911,N_5713,N_5720);
nor U5912 (N_5912,N_5702,N_5757);
xor U5913 (N_5913,N_5725,N_5611);
nand U5914 (N_5914,N_5716,N_5712);
and U5915 (N_5915,N_5614,N_5619);
nand U5916 (N_5916,N_5680,N_5719);
xor U5917 (N_5917,N_5669,N_5746);
and U5918 (N_5918,N_5681,N_5600);
or U5919 (N_5919,N_5620,N_5669);
xor U5920 (N_5920,N_5765,N_5607);
xor U5921 (N_5921,N_5670,N_5638);
xor U5922 (N_5922,N_5650,N_5790);
nand U5923 (N_5923,N_5690,N_5798);
xor U5924 (N_5924,N_5782,N_5734);
and U5925 (N_5925,N_5712,N_5626);
xnor U5926 (N_5926,N_5789,N_5626);
and U5927 (N_5927,N_5788,N_5609);
nand U5928 (N_5928,N_5642,N_5745);
xor U5929 (N_5929,N_5740,N_5790);
or U5930 (N_5930,N_5711,N_5725);
nand U5931 (N_5931,N_5790,N_5709);
nor U5932 (N_5932,N_5713,N_5780);
xor U5933 (N_5933,N_5696,N_5695);
or U5934 (N_5934,N_5619,N_5738);
nand U5935 (N_5935,N_5688,N_5683);
xor U5936 (N_5936,N_5752,N_5773);
or U5937 (N_5937,N_5609,N_5678);
nor U5938 (N_5938,N_5734,N_5605);
xor U5939 (N_5939,N_5737,N_5773);
or U5940 (N_5940,N_5730,N_5775);
and U5941 (N_5941,N_5670,N_5730);
nor U5942 (N_5942,N_5655,N_5650);
nand U5943 (N_5943,N_5760,N_5605);
and U5944 (N_5944,N_5725,N_5691);
or U5945 (N_5945,N_5669,N_5732);
nand U5946 (N_5946,N_5613,N_5680);
and U5947 (N_5947,N_5717,N_5796);
and U5948 (N_5948,N_5799,N_5698);
and U5949 (N_5949,N_5637,N_5656);
and U5950 (N_5950,N_5653,N_5671);
nor U5951 (N_5951,N_5705,N_5736);
nor U5952 (N_5952,N_5729,N_5776);
xor U5953 (N_5953,N_5609,N_5785);
and U5954 (N_5954,N_5765,N_5693);
xor U5955 (N_5955,N_5677,N_5711);
or U5956 (N_5956,N_5652,N_5653);
and U5957 (N_5957,N_5777,N_5624);
or U5958 (N_5958,N_5766,N_5674);
nand U5959 (N_5959,N_5711,N_5650);
or U5960 (N_5960,N_5691,N_5601);
and U5961 (N_5961,N_5602,N_5629);
or U5962 (N_5962,N_5729,N_5649);
xor U5963 (N_5963,N_5684,N_5685);
nand U5964 (N_5964,N_5751,N_5713);
nor U5965 (N_5965,N_5697,N_5688);
nand U5966 (N_5966,N_5758,N_5685);
or U5967 (N_5967,N_5634,N_5733);
or U5968 (N_5968,N_5795,N_5696);
nand U5969 (N_5969,N_5655,N_5661);
and U5970 (N_5970,N_5788,N_5657);
xnor U5971 (N_5971,N_5635,N_5667);
nor U5972 (N_5972,N_5744,N_5703);
xor U5973 (N_5973,N_5645,N_5678);
or U5974 (N_5974,N_5705,N_5609);
and U5975 (N_5975,N_5622,N_5694);
nor U5976 (N_5976,N_5704,N_5641);
nand U5977 (N_5977,N_5613,N_5676);
and U5978 (N_5978,N_5726,N_5796);
or U5979 (N_5979,N_5716,N_5709);
and U5980 (N_5980,N_5746,N_5734);
nor U5981 (N_5981,N_5659,N_5705);
xor U5982 (N_5982,N_5709,N_5726);
nand U5983 (N_5983,N_5785,N_5769);
or U5984 (N_5984,N_5701,N_5741);
or U5985 (N_5985,N_5787,N_5792);
nand U5986 (N_5986,N_5665,N_5725);
and U5987 (N_5987,N_5776,N_5653);
nand U5988 (N_5988,N_5668,N_5761);
or U5989 (N_5989,N_5716,N_5738);
xnor U5990 (N_5990,N_5783,N_5686);
or U5991 (N_5991,N_5767,N_5683);
or U5992 (N_5992,N_5779,N_5777);
or U5993 (N_5993,N_5699,N_5687);
and U5994 (N_5994,N_5716,N_5748);
nor U5995 (N_5995,N_5797,N_5627);
nand U5996 (N_5996,N_5670,N_5643);
nand U5997 (N_5997,N_5734,N_5790);
nor U5998 (N_5998,N_5755,N_5785);
nor U5999 (N_5999,N_5633,N_5698);
nand U6000 (N_6000,N_5841,N_5983);
nor U6001 (N_6001,N_5846,N_5889);
and U6002 (N_6002,N_5862,N_5850);
xnor U6003 (N_6003,N_5927,N_5806);
or U6004 (N_6004,N_5988,N_5972);
and U6005 (N_6005,N_5948,N_5808);
and U6006 (N_6006,N_5879,N_5935);
nand U6007 (N_6007,N_5807,N_5981);
or U6008 (N_6008,N_5857,N_5893);
nand U6009 (N_6009,N_5804,N_5837);
or U6010 (N_6010,N_5887,N_5845);
nand U6011 (N_6011,N_5928,N_5914);
nand U6012 (N_6012,N_5951,N_5913);
xor U6013 (N_6013,N_5884,N_5836);
nor U6014 (N_6014,N_5949,N_5847);
nand U6015 (N_6015,N_5896,N_5819);
nor U6016 (N_6016,N_5980,N_5805);
or U6017 (N_6017,N_5973,N_5921);
nand U6018 (N_6018,N_5829,N_5865);
nor U6019 (N_6019,N_5801,N_5894);
nor U6020 (N_6020,N_5968,N_5957);
nand U6021 (N_6021,N_5833,N_5956);
nor U6022 (N_6022,N_5892,N_5964);
or U6023 (N_6023,N_5946,N_5963);
nand U6024 (N_6024,N_5938,N_5978);
nand U6025 (N_6025,N_5838,N_5975);
nor U6026 (N_6026,N_5891,N_5911);
xor U6027 (N_6027,N_5835,N_5965);
or U6028 (N_6028,N_5851,N_5912);
nor U6029 (N_6029,N_5967,N_5942);
xor U6030 (N_6030,N_5877,N_5936);
and U6031 (N_6031,N_5955,N_5998);
xor U6032 (N_6032,N_5849,N_5809);
nand U6033 (N_6033,N_5864,N_5999);
or U6034 (N_6034,N_5867,N_5823);
xnor U6035 (N_6035,N_5944,N_5947);
nor U6036 (N_6036,N_5876,N_5843);
or U6037 (N_6037,N_5868,N_5922);
or U6038 (N_6038,N_5923,N_5901);
or U6039 (N_6039,N_5918,N_5994);
xor U6040 (N_6040,N_5989,N_5910);
or U6041 (N_6041,N_5869,N_5916);
or U6042 (N_6042,N_5858,N_5840);
and U6043 (N_6043,N_5834,N_5990);
and U6044 (N_6044,N_5900,N_5976);
xor U6045 (N_6045,N_5822,N_5888);
xnor U6046 (N_6046,N_5943,N_5954);
nand U6047 (N_6047,N_5908,N_5812);
nor U6048 (N_6048,N_5969,N_5826);
nand U6049 (N_6049,N_5919,N_5930);
nand U6050 (N_6050,N_5926,N_5933);
xor U6051 (N_6051,N_5952,N_5945);
and U6052 (N_6052,N_5830,N_5881);
or U6053 (N_6053,N_5971,N_5953);
nand U6054 (N_6054,N_5813,N_5905);
nor U6055 (N_6055,N_5871,N_5863);
nand U6056 (N_6056,N_5992,N_5842);
xor U6057 (N_6057,N_5902,N_5925);
xor U6058 (N_6058,N_5950,N_5873);
xor U6059 (N_6059,N_5825,N_5960);
nand U6060 (N_6060,N_5985,N_5939);
xnor U6061 (N_6061,N_5997,N_5872);
xor U6062 (N_6062,N_5931,N_5984);
xor U6063 (N_6063,N_5929,N_5866);
or U6064 (N_6064,N_5800,N_5816);
nand U6065 (N_6065,N_5920,N_5870);
nand U6066 (N_6066,N_5970,N_5828);
nor U6067 (N_6067,N_5979,N_5906);
nor U6068 (N_6068,N_5909,N_5993);
and U6069 (N_6069,N_5853,N_5839);
nor U6070 (N_6070,N_5995,N_5982);
nor U6071 (N_6071,N_5855,N_5860);
or U6072 (N_6072,N_5821,N_5915);
nor U6073 (N_6073,N_5861,N_5885);
xor U6074 (N_6074,N_5882,N_5924);
nor U6075 (N_6075,N_5974,N_5904);
xnor U6076 (N_6076,N_5811,N_5886);
or U6077 (N_6077,N_5987,N_5977);
or U6078 (N_6078,N_5880,N_5820);
and U6079 (N_6079,N_5890,N_5898);
nor U6080 (N_6080,N_5824,N_5934);
nand U6081 (N_6081,N_5844,N_5831);
or U6082 (N_6082,N_5961,N_5996);
xor U6083 (N_6083,N_5827,N_5940);
or U6084 (N_6084,N_5895,N_5917);
and U6085 (N_6085,N_5854,N_5832);
nor U6086 (N_6086,N_5959,N_5802);
or U6087 (N_6087,N_5899,N_5818);
nand U6088 (N_6088,N_5897,N_5932);
and U6089 (N_6089,N_5803,N_5883);
nand U6090 (N_6090,N_5814,N_5848);
and U6091 (N_6091,N_5817,N_5941);
nand U6092 (N_6092,N_5958,N_5859);
nor U6093 (N_6093,N_5878,N_5815);
or U6094 (N_6094,N_5903,N_5875);
nor U6095 (N_6095,N_5856,N_5907);
and U6096 (N_6096,N_5962,N_5810);
or U6097 (N_6097,N_5852,N_5874);
or U6098 (N_6098,N_5991,N_5986);
nand U6099 (N_6099,N_5937,N_5966);
nand U6100 (N_6100,N_5920,N_5959);
nor U6101 (N_6101,N_5949,N_5812);
nand U6102 (N_6102,N_5905,N_5961);
and U6103 (N_6103,N_5806,N_5997);
xnor U6104 (N_6104,N_5976,N_5927);
nand U6105 (N_6105,N_5914,N_5805);
or U6106 (N_6106,N_5856,N_5936);
nand U6107 (N_6107,N_5907,N_5989);
nand U6108 (N_6108,N_5952,N_5803);
xor U6109 (N_6109,N_5832,N_5839);
nor U6110 (N_6110,N_5828,N_5897);
and U6111 (N_6111,N_5922,N_5949);
or U6112 (N_6112,N_5912,N_5894);
nand U6113 (N_6113,N_5998,N_5968);
or U6114 (N_6114,N_5952,N_5959);
nand U6115 (N_6115,N_5932,N_5998);
and U6116 (N_6116,N_5865,N_5815);
or U6117 (N_6117,N_5991,N_5956);
xnor U6118 (N_6118,N_5956,N_5880);
nand U6119 (N_6119,N_5980,N_5876);
xnor U6120 (N_6120,N_5900,N_5951);
nor U6121 (N_6121,N_5889,N_5897);
nand U6122 (N_6122,N_5942,N_5846);
and U6123 (N_6123,N_5939,N_5903);
xor U6124 (N_6124,N_5897,N_5847);
nand U6125 (N_6125,N_5919,N_5970);
nor U6126 (N_6126,N_5980,N_5822);
nand U6127 (N_6127,N_5924,N_5890);
and U6128 (N_6128,N_5839,N_5961);
or U6129 (N_6129,N_5979,N_5887);
nor U6130 (N_6130,N_5889,N_5864);
or U6131 (N_6131,N_5892,N_5884);
or U6132 (N_6132,N_5854,N_5991);
and U6133 (N_6133,N_5930,N_5980);
nand U6134 (N_6134,N_5805,N_5873);
or U6135 (N_6135,N_5966,N_5861);
or U6136 (N_6136,N_5924,N_5817);
nand U6137 (N_6137,N_5866,N_5998);
xnor U6138 (N_6138,N_5910,N_5949);
or U6139 (N_6139,N_5981,N_5833);
or U6140 (N_6140,N_5973,N_5882);
or U6141 (N_6141,N_5838,N_5899);
nor U6142 (N_6142,N_5841,N_5820);
nand U6143 (N_6143,N_5959,N_5921);
nor U6144 (N_6144,N_5901,N_5965);
and U6145 (N_6145,N_5966,N_5948);
xnor U6146 (N_6146,N_5964,N_5957);
nor U6147 (N_6147,N_5939,N_5861);
and U6148 (N_6148,N_5997,N_5903);
nand U6149 (N_6149,N_5887,N_5848);
nor U6150 (N_6150,N_5899,N_5918);
nor U6151 (N_6151,N_5962,N_5928);
nor U6152 (N_6152,N_5954,N_5941);
or U6153 (N_6153,N_5857,N_5888);
nand U6154 (N_6154,N_5903,N_5959);
or U6155 (N_6155,N_5829,N_5961);
or U6156 (N_6156,N_5849,N_5828);
and U6157 (N_6157,N_5851,N_5850);
nor U6158 (N_6158,N_5960,N_5970);
and U6159 (N_6159,N_5914,N_5867);
xnor U6160 (N_6160,N_5937,N_5862);
nor U6161 (N_6161,N_5955,N_5824);
nor U6162 (N_6162,N_5921,N_5877);
or U6163 (N_6163,N_5902,N_5966);
xnor U6164 (N_6164,N_5981,N_5871);
xor U6165 (N_6165,N_5901,N_5912);
nor U6166 (N_6166,N_5902,N_5884);
nand U6167 (N_6167,N_5929,N_5937);
and U6168 (N_6168,N_5813,N_5852);
xnor U6169 (N_6169,N_5854,N_5855);
or U6170 (N_6170,N_5881,N_5842);
xnor U6171 (N_6171,N_5913,N_5833);
xor U6172 (N_6172,N_5832,N_5961);
or U6173 (N_6173,N_5890,N_5823);
or U6174 (N_6174,N_5945,N_5811);
nand U6175 (N_6175,N_5825,N_5999);
nand U6176 (N_6176,N_5812,N_5828);
nor U6177 (N_6177,N_5901,N_5928);
and U6178 (N_6178,N_5955,N_5963);
xnor U6179 (N_6179,N_5952,N_5812);
nor U6180 (N_6180,N_5871,N_5854);
and U6181 (N_6181,N_5966,N_5873);
nor U6182 (N_6182,N_5834,N_5805);
nand U6183 (N_6183,N_5980,N_5935);
nand U6184 (N_6184,N_5854,N_5918);
and U6185 (N_6185,N_5890,N_5960);
nor U6186 (N_6186,N_5839,N_5884);
xor U6187 (N_6187,N_5913,N_5814);
nand U6188 (N_6188,N_5985,N_5854);
or U6189 (N_6189,N_5953,N_5821);
nor U6190 (N_6190,N_5839,N_5860);
or U6191 (N_6191,N_5905,N_5895);
or U6192 (N_6192,N_5873,N_5942);
nand U6193 (N_6193,N_5849,N_5874);
nand U6194 (N_6194,N_5802,N_5945);
xor U6195 (N_6195,N_5886,N_5909);
nand U6196 (N_6196,N_5922,N_5852);
and U6197 (N_6197,N_5881,N_5998);
xnor U6198 (N_6198,N_5838,N_5833);
nand U6199 (N_6199,N_5922,N_5820);
xor U6200 (N_6200,N_6076,N_6084);
xnor U6201 (N_6201,N_6056,N_6174);
nor U6202 (N_6202,N_6196,N_6189);
nand U6203 (N_6203,N_6141,N_6022);
nor U6204 (N_6204,N_6015,N_6170);
or U6205 (N_6205,N_6191,N_6146);
nand U6206 (N_6206,N_6098,N_6023);
nor U6207 (N_6207,N_6100,N_6178);
nand U6208 (N_6208,N_6094,N_6061);
and U6209 (N_6209,N_6008,N_6129);
xnor U6210 (N_6210,N_6135,N_6122);
nand U6211 (N_6211,N_6077,N_6085);
nand U6212 (N_6212,N_6165,N_6169);
and U6213 (N_6213,N_6025,N_6046);
or U6214 (N_6214,N_6075,N_6168);
and U6215 (N_6215,N_6137,N_6062);
xor U6216 (N_6216,N_6043,N_6116);
nor U6217 (N_6217,N_6186,N_6029);
xor U6218 (N_6218,N_6158,N_6014);
nor U6219 (N_6219,N_6037,N_6193);
and U6220 (N_6220,N_6059,N_6065);
nor U6221 (N_6221,N_6074,N_6149);
and U6222 (N_6222,N_6195,N_6063);
nand U6223 (N_6223,N_6090,N_6053);
nor U6224 (N_6224,N_6071,N_6048);
nor U6225 (N_6225,N_6114,N_6028);
nand U6226 (N_6226,N_6128,N_6067);
and U6227 (N_6227,N_6087,N_6181);
xnor U6228 (N_6228,N_6013,N_6017);
nor U6229 (N_6229,N_6197,N_6187);
or U6230 (N_6230,N_6134,N_6182);
nand U6231 (N_6231,N_6180,N_6138);
nor U6232 (N_6232,N_6069,N_6111);
and U6233 (N_6233,N_6064,N_6119);
nand U6234 (N_6234,N_6002,N_6167);
or U6235 (N_6235,N_6035,N_6089);
nand U6236 (N_6236,N_6120,N_6072);
nor U6237 (N_6237,N_6096,N_6131);
nor U6238 (N_6238,N_6162,N_6007);
xnor U6239 (N_6239,N_6026,N_6126);
or U6240 (N_6240,N_6109,N_6052);
or U6241 (N_6241,N_6051,N_6117);
nand U6242 (N_6242,N_6018,N_6107);
and U6243 (N_6243,N_6112,N_6038);
and U6244 (N_6244,N_6054,N_6009);
nor U6245 (N_6245,N_6095,N_6148);
nor U6246 (N_6246,N_6130,N_6024);
nor U6247 (N_6247,N_6097,N_6171);
and U6248 (N_6248,N_6124,N_6034);
or U6249 (N_6249,N_6042,N_6190);
nand U6250 (N_6250,N_6088,N_6123);
xnor U6251 (N_6251,N_6152,N_6093);
xnor U6252 (N_6252,N_6155,N_6082);
and U6253 (N_6253,N_6176,N_6183);
and U6254 (N_6254,N_6006,N_6143);
nor U6255 (N_6255,N_6102,N_6081);
nor U6256 (N_6256,N_6091,N_6060);
or U6257 (N_6257,N_6140,N_6184);
nand U6258 (N_6258,N_6055,N_6106);
or U6259 (N_6259,N_6033,N_6080);
nand U6260 (N_6260,N_6086,N_6147);
nand U6261 (N_6261,N_6113,N_6150);
xnor U6262 (N_6262,N_6153,N_6172);
nor U6263 (N_6263,N_6031,N_6011);
nand U6264 (N_6264,N_6010,N_6066);
nand U6265 (N_6265,N_6045,N_6103);
or U6266 (N_6266,N_6099,N_6125);
xor U6267 (N_6267,N_6020,N_6157);
nand U6268 (N_6268,N_6040,N_6199);
and U6269 (N_6269,N_6049,N_6027);
xnor U6270 (N_6270,N_6078,N_6001);
nor U6271 (N_6271,N_6012,N_6164);
xor U6272 (N_6272,N_6121,N_6083);
nand U6273 (N_6273,N_6163,N_6047);
and U6274 (N_6274,N_6005,N_6050);
nor U6275 (N_6275,N_6173,N_6188);
nor U6276 (N_6276,N_6144,N_6185);
or U6277 (N_6277,N_6036,N_6104);
nand U6278 (N_6278,N_6068,N_6079);
xor U6279 (N_6279,N_6108,N_6105);
nor U6280 (N_6280,N_6154,N_6156);
xnor U6281 (N_6281,N_6016,N_6132);
xor U6282 (N_6282,N_6041,N_6057);
nand U6283 (N_6283,N_6070,N_6003);
or U6284 (N_6284,N_6160,N_6118);
and U6285 (N_6285,N_6159,N_6194);
nor U6286 (N_6286,N_6039,N_6030);
or U6287 (N_6287,N_6115,N_6139);
or U6288 (N_6288,N_6145,N_6175);
and U6289 (N_6289,N_6110,N_6058);
and U6290 (N_6290,N_6151,N_6101);
or U6291 (N_6291,N_6004,N_6161);
or U6292 (N_6292,N_6166,N_6127);
or U6293 (N_6293,N_6192,N_6021);
or U6294 (N_6294,N_6136,N_6000);
xor U6295 (N_6295,N_6179,N_6198);
nor U6296 (N_6296,N_6092,N_6073);
xor U6297 (N_6297,N_6142,N_6177);
nand U6298 (N_6298,N_6044,N_6019);
nand U6299 (N_6299,N_6032,N_6133);
xnor U6300 (N_6300,N_6049,N_6100);
xor U6301 (N_6301,N_6029,N_6001);
or U6302 (N_6302,N_6121,N_6140);
nor U6303 (N_6303,N_6047,N_6003);
xor U6304 (N_6304,N_6032,N_6037);
nand U6305 (N_6305,N_6128,N_6171);
or U6306 (N_6306,N_6073,N_6066);
or U6307 (N_6307,N_6125,N_6161);
nand U6308 (N_6308,N_6076,N_6157);
nor U6309 (N_6309,N_6093,N_6083);
and U6310 (N_6310,N_6122,N_6173);
nor U6311 (N_6311,N_6185,N_6072);
nor U6312 (N_6312,N_6049,N_6112);
xor U6313 (N_6313,N_6131,N_6090);
and U6314 (N_6314,N_6192,N_6077);
or U6315 (N_6315,N_6071,N_6178);
or U6316 (N_6316,N_6001,N_6162);
or U6317 (N_6317,N_6026,N_6051);
and U6318 (N_6318,N_6077,N_6056);
nor U6319 (N_6319,N_6101,N_6014);
or U6320 (N_6320,N_6035,N_6028);
xor U6321 (N_6321,N_6126,N_6098);
and U6322 (N_6322,N_6076,N_6096);
nand U6323 (N_6323,N_6029,N_6070);
or U6324 (N_6324,N_6134,N_6090);
nor U6325 (N_6325,N_6022,N_6165);
nand U6326 (N_6326,N_6035,N_6068);
and U6327 (N_6327,N_6062,N_6047);
xnor U6328 (N_6328,N_6155,N_6075);
nor U6329 (N_6329,N_6100,N_6155);
xor U6330 (N_6330,N_6098,N_6143);
and U6331 (N_6331,N_6158,N_6139);
nor U6332 (N_6332,N_6127,N_6154);
nor U6333 (N_6333,N_6174,N_6089);
nor U6334 (N_6334,N_6145,N_6064);
nor U6335 (N_6335,N_6117,N_6071);
nor U6336 (N_6336,N_6015,N_6199);
or U6337 (N_6337,N_6185,N_6019);
or U6338 (N_6338,N_6023,N_6137);
xor U6339 (N_6339,N_6141,N_6119);
xor U6340 (N_6340,N_6116,N_6145);
nor U6341 (N_6341,N_6016,N_6107);
nand U6342 (N_6342,N_6187,N_6037);
xor U6343 (N_6343,N_6157,N_6032);
nor U6344 (N_6344,N_6077,N_6031);
and U6345 (N_6345,N_6199,N_6165);
xor U6346 (N_6346,N_6168,N_6026);
and U6347 (N_6347,N_6137,N_6172);
nand U6348 (N_6348,N_6183,N_6049);
and U6349 (N_6349,N_6055,N_6199);
and U6350 (N_6350,N_6119,N_6038);
xnor U6351 (N_6351,N_6054,N_6095);
xor U6352 (N_6352,N_6003,N_6129);
and U6353 (N_6353,N_6003,N_6106);
xnor U6354 (N_6354,N_6055,N_6029);
and U6355 (N_6355,N_6111,N_6193);
or U6356 (N_6356,N_6174,N_6176);
xor U6357 (N_6357,N_6109,N_6169);
nor U6358 (N_6358,N_6146,N_6155);
or U6359 (N_6359,N_6019,N_6094);
or U6360 (N_6360,N_6176,N_6119);
nand U6361 (N_6361,N_6199,N_6181);
nor U6362 (N_6362,N_6073,N_6061);
nor U6363 (N_6363,N_6146,N_6090);
or U6364 (N_6364,N_6124,N_6183);
nand U6365 (N_6365,N_6020,N_6171);
nand U6366 (N_6366,N_6005,N_6041);
and U6367 (N_6367,N_6027,N_6026);
nand U6368 (N_6368,N_6059,N_6082);
xnor U6369 (N_6369,N_6050,N_6091);
or U6370 (N_6370,N_6040,N_6075);
xor U6371 (N_6371,N_6014,N_6174);
and U6372 (N_6372,N_6100,N_6084);
or U6373 (N_6373,N_6114,N_6151);
xor U6374 (N_6374,N_6193,N_6165);
and U6375 (N_6375,N_6035,N_6041);
or U6376 (N_6376,N_6097,N_6194);
nand U6377 (N_6377,N_6039,N_6197);
xnor U6378 (N_6378,N_6041,N_6143);
nor U6379 (N_6379,N_6025,N_6049);
and U6380 (N_6380,N_6168,N_6166);
or U6381 (N_6381,N_6062,N_6078);
nor U6382 (N_6382,N_6155,N_6152);
xnor U6383 (N_6383,N_6081,N_6030);
nand U6384 (N_6384,N_6146,N_6118);
xnor U6385 (N_6385,N_6033,N_6087);
nor U6386 (N_6386,N_6063,N_6161);
or U6387 (N_6387,N_6182,N_6106);
nor U6388 (N_6388,N_6111,N_6136);
and U6389 (N_6389,N_6076,N_6027);
nand U6390 (N_6390,N_6065,N_6080);
nand U6391 (N_6391,N_6038,N_6140);
nand U6392 (N_6392,N_6003,N_6074);
xor U6393 (N_6393,N_6173,N_6170);
or U6394 (N_6394,N_6065,N_6119);
nand U6395 (N_6395,N_6004,N_6072);
or U6396 (N_6396,N_6068,N_6029);
xnor U6397 (N_6397,N_6008,N_6022);
and U6398 (N_6398,N_6010,N_6118);
xnor U6399 (N_6399,N_6185,N_6007);
and U6400 (N_6400,N_6247,N_6266);
nor U6401 (N_6401,N_6383,N_6245);
or U6402 (N_6402,N_6293,N_6224);
and U6403 (N_6403,N_6390,N_6315);
and U6404 (N_6404,N_6254,N_6201);
and U6405 (N_6405,N_6292,N_6208);
nand U6406 (N_6406,N_6327,N_6377);
nand U6407 (N_6407,N_6299,N_6213);
or U6408 (N_6408,N_6338,N_6361);
nand U6409 (N_6409,N_6270,N_6303);
or U6410 (N_6410,N_6207,N_6221);
xnor U6411 (N_6411,N_6263,N_6230);
or U6412 (N_6412,N_6310,N_6272);
nand U6413 (N_6413,N_6333,N_6211);
nor U6414 (N_6414,N_6283,N_6260);
xor U6415 (N_6415,N_6284,N_6243);
or U6416 (N_6416,N_6236,N_6366);
nand U6417 (N_6417,N_6351,N_6205);
or U6418 (N_6418,N_6250,N_6295);
or U6419 (N_6419,N_6352,N_6334);
or U6420 (N_6420,N_6273,N_6244);
xnor U6421 (N_6421,N_6335,N_6340);
nand U6422 (N_6422,N_6281,N_6350);
or U6423 (N_6423,N_6306,N_6395);
xnor U6424 (N_6424,N_6368,N_6380);
nor U6425 (N_6425,N_6242,N_6268);
nor U6426 (N_6426,N_6277,N_6210);
and U6427 (N_6427,N_6288,N_6328);
or U6428 (N_6428,N_6233,N_6339);
xor U6429 (N_6429,N_6342,N_6323);
or U6430 (N_6430,N_6290,N_6349);
nor U6431 (N_6431,N_6389,N_6225);
and U6432 (N_6432,N_6382,N_6379);
xnor U6433 (N_6433,N_6325,N_6316);
and U6434 (N_6434,N_6364,N_6397);
or U6435 (N_6435,N_6394,N_6219);
and U6436 (N_6436,N_6354,N_6256);
and U6437 (N_6437,N_6291,N_6238);
nor U6438 (N_6438,N_6276,N_6232);
and U6439 (N_6439,N_6375,N_6248);
xor U6440 (N_6440,N_6320,N_6304);
nand U6441 (N_6441,N_6282,N_6367);
nand U6442 (N_6442,N_6302,N_6384);
and U6443 (N_6443,N_6330,N_6278);
or U6444 (N_6444,N_6312,N_6259);
nor U6445 (N_6445,N_6345,N_6216);
or U6446 (N_6446,N_6285,N_6241);
nor U6447 (N_6447,N_6381,N_6309);
xor U6448 (N_6448,N_6212,N_6321);
and U6449 (N_6449,N_6300,N_6324);
nand U6450 (N_6450,N_6275,N_6329);
nor U6451 (N_6451,N_6264,N_6296);
or U6452 (N_6452,N_6279,N_6344);
nor U6453 (N_6453,N_6267,N_6217);
nor U6454 (N_6454,N_6200,N_6258);
nor U6455 (N_6455,N_6398,N_6249);
nor U6456 (N_6456,N_6369,N_6360);
nor U6457 (N_6457,N_6255,N_6286);
and U6458 (N_6458,N_6239,N_6331);
and U6459 (N_6459,N_6374,N_6376);
nor U6460 (N_6460,N_6246,N_6388);
and U6461 (N_6461,N_6308,N_6265);
xor U6462 (N_6462,N_6240,N_6372);
nor U6463 (N_6463,N_6347,N_6362);
nor U6464 (N_6464,N_6203,N_6378);
and U6465 (N_6465,N_6237,N_6346);
or U6466 (N_6466,N_6271,N_6348);
or U6467 (N_6467,N_6298,N_6357);
or U6468 (N_6468,N_6214,N_6355);
xor U6469 (N_6469,N_6391,N_6253);
nand U6470 (N_6470,N_6294,N_6385);
nand U6471 (N_6471,N_6204,N_6341);
xor U6472 (N_6472,N_6222,N_6274);
nand U6473 (N_6473,N_6363,N_6257);
or U6474 (N_6474,N_6371,N_6359);
nor U6475 (N_6475,N_6336,N_6392);
nor U6476 (N_6476,N_6234,N_6218);
and U6477 (N_6477,N_6206,N_6301);
xor U6478 (N_6478,N_6317,N_6319);
nand U6479 (N_6479,N_6365,N_6227);
nor U6480 (N_6480,N_6370,N_6373);
nor U6481 (N_6481,N_6215,N_6202);
or U6482 (N_6482,N_6314,N_6280);
and U6483 (N_6483,N_6386,N_6251);
nand U6484 (N_6484,N_6289,N_6262);
and U6485 (N_6485,N_6343,N_6318);
and U6486 (N_6486,N_6356,N_6220);
nand U6487 (N_6487,N_6223,N_6393);
nand U6488 (N_6488,N_6387,N_6209);
xnor U6489 (N_6489,N_6322,N_6261);
nand U6490 (N_6490,N_6287,N_6297);
xor U6491 (N_6491,N_6311,N_6228);
xnor U6492 (N_6492,N_6326,N_6353);
or U6493 (N_6493,N_6252,N_6332);
and U6494 (N_6494,N_6396,N_6226);
or U6495 (N_6495,N_6307,N_6231);
and U6496 (N_6496,N_6399,N_6269);
xor U6497 (N_6497,N_6305,N_6235);
nand U6498 (N_6498,N_6313,N_6229);
xor U6499 (N_6499,N_6358,N_6337);
nor U6500 (N_6500,N_6237,N_6286);
nor U6501 (N_6501,N_6381,N_6216);
xor U6502 (N_6502,N_6384,N_6334);
or U6503 (N_6503,N_6345,N_6244);
nor U6504 (N_6504,N_6328,N_6253);
nand U6505 (N_6505,N_6309,N_6258);
xor U6506 (N_6506,N_6233,N_6235);
nor U6507 (N_6507,N_6290,N_6227);
xor U6508 (N_6508,N_6238,N_6342);
nor U6509 (N_6509,N_6329,N_6387);
xor U6510 (N_6510,N_6203,N_6389);
nor U6511 (N_6511,N_6286,N_6270);
and U6512 (N_6512,N_6373,N_6290);
xnor U6513 (N_6513,N_6270,N_6232);
xnor U6514 (N_6514,N_6319,N_6210);
nand U6515 (N_6515,N_6309,N_6358);
or U6516 (N_6516,N_6260,N_6201);
nand U6517 (N_6517,N_6241,N_6245);
nand U6518 (N_6518,N_6218,N_6391);
and U6519 (N_6519,N_6260,N_6248);
or U6520 (N_6520,N_6332,N_6393);
and U6521 (N_6521,N_6334,N_6389);
nand U6522 (N_6522,N_6245,N_6313);
nor U6523 (N_6523,N_6271,N_6399);
nor U6524 (N_6524,N_6316,N_6372);
xor U6525 (N_6525,N_6384,N_6325);
nor U6526 (N_6526,N_6280,N_6209);
or U6527 (N_6527,N_6364,N_6382);
xor U6528 (N_6528,N_6201,N_6353);
nand U6529 (N_6529,N_6317,N_6320);
nand U6530 (N_6530,N_6200,N_6342);
nand U6531 (N_6531,N_6366,N_6206);
and U6532 (N_6532,N_6335,N_6331);
or U6533 (N_6533,N_6291,N_6273);
or U6534 (N_6534,N_6248,N_6340);
nand U6535 (N_6535,N_6279,N_6365);
xnor U6536 (N_6536,N_6224,N_6221);
nand U6537 (N_6537,N_6372,N_6264);
or U6538 (N_6538,N_6382,N_6308);
xnor U6539 (N_6539,N_6259,N_6279);
nor U6540 (N_6540,N_6289,N_6337);
xor U6541 (N_6541,N_6363,N_6289);
nor U6542 (N_6542,N_6213,N_6395);
and U6543 (N_6543,N_6288,N_6373);
nor U6544 (N_6544,N_6393,N_6293);
or U6545 (N_6545,N_6228,N_6209);
nor U6546 (N_6546,N_6320,N_6213);
or U6547 (N_6547,N_6348,N_6217);
xnor U6548 (N_6548,N_6335,N_6321);
and U6549 (N_6549,N_6398,N_6295);
and U6550 (N_6550,N_6372,N_6330);
and U6551 (N_6551,N_6200,N_6305);
and U6552 (N_6552,N_6359,N_6386);
xor U6553 (N_6553,N_6230,N_6312);
nand U6554 (N_6554,N_6208,N_6211);
nor U6555 (N_6555,N_6232,N_6339);
nand U6556 (N_6556,N_6395,N_6232);
nand U6557 (N_6557,N_6335,N_6231);
nor U6558 (N_6558,N_6209,N_6248);
nor U6559 (N_6559,N_6386,N_6367);
nor U6560 (N_6560,N_6301,N_6287);
and U6561 (N_6561,N_6205,N_6385);
xnor U6562 (N_6562,N_6215,N_6228);
nand U6563 (N_6563,N_6343,N_6223);
nand U6564 (N_6564,N_6392,N_6240);
or U6565 (N_6565,N_6233,N_6216);
nor U6566 (N_6566,N_6298,N_6208);
or U6567 (N_6567,N_6305,N_6342);
xor U6568 (N_6568,N_6318,N_6379);
nor U6569 (N_6569,N_6293,N_6225);
and U6570 (N_6570,N_6267,N_6334);
nor U6571 (N_6571,N_6343,N_6358);
nand U6572 (N_6572,N_6238,N_6220);
xnor U6573 (N_6573,N_6273,N_6296);
xnor U6574 (N_6574,N_6337,N_6225);
xor U6575 (N_6575,N_6218,N_6281);
nor U6576 (N_6576,N_6321,N_6207);
nor U6577 (N_6577,N_6291,N_6241);
or U6578 (N_6578,N_6228,N_6323);
nand U6579 (N_6579,N_6389,N_6297);
nand U6580 (N_6580,N_6223,N_6263);
and U6581 (N_6581,N_6333,N_6392);
nor U6582 (N_6582,N_6258,N_6332);
nor U6583 (N_6583,N_6369,N_6201);
xor U6584 (N_6584,N_6298,N_6334);
xnor U6585 (N_6585,N_6317,N_6237);
xor U6586 (N_6586,N_6205,N_6391);
or U6587 (N_6587,N_6262,N_6395);
and U6588 (N_6588,N_6376,N_6395);
nor U6589 (N_6589,N_6344,N_6224);
xnor U6590 (N_6590,N_6244,N_6240);
xnor U6591 (N_6591,N_6389,N_6308);
nor U6592 (N_6592,N_6326,N_6242);
and U6593 (N_6593,N_6382,N_6315);
xnor U6594 (N_6594,N_6304,N_6262);
nor U6595 (N_6595,N_6329,N_6213);
or U6596 (N_6596,N_6307,N_6344);
nor U6597 (N_6597,N_6331,N_6351);
and U6598 (N_6598,N_6287,N_6398);
nand U6599 (N_6599,N_6281,N_6370);
xor U6600 (N_6600,N_6483,N_6413);
or U6601 (N_6601,N_6482,N_6594);
nand U6602 (N_6602,N_6530,N_6465);
nand U6603 (N_6603,N_6432,N_6584);
xnor U6604 (N_6604,N_6533,N_6480);
nand U6605 (N_6605,N_6405,N_6433);
xnor U6606 (N_6606,N_6516,N_6559);
or U6607 (N_6607,N_6403,N_6458);
nand U6608 (N_6608,N_6415,N_6464);
nor U6609 (N_6609,N_6474,N_6579);
or U6610 (N_6610,N_6434,N_6498);
xnor U6611 (N_6611,N_6492,N_6538);
and U6612 (N_6612,N_6549,N_6410);
xor U6613 (N_6613,N_6572,N_6451);
and U6614 (N_6614,N_6588,N_6449);
nor U6615 (N_6615,N_6472,N_6519);
nand U6616 (N_6616,N_6551,N_6445);
xor U6617 (N_6617,N_6528,N_6564);
nor U6618 (N_6618,N_6543,N_6456);
and U6619 (N_6619,N_6556,N_6406);
nand U6620 (N_6620,N_6489,N_6475);
xor U6621 (N_6621,N_6504,N_6425);
nor U6622 (N_6622,N_6452,N_6505);
or U6623 (N_6623,N_6502,N_6487);
or U6624 (N_6624,N_6422,N_6414);
xnor U6625 (N_6625,N_6591,N_6524);
xor U6626 (N_6626,N_6440,N_6486);
nand U6627 (N_6627,N_6478,N_6525);
nor U6628 (N_6628,N_6523,N_6575);
xnor U6629 (N_6629,N_6419,N_6454);
and U6630 (N_6630,N_6548,N_6597);
and U6631 (N_6631,N_6539,N_6471);
or U6632 (N_6632,N_6411,N_6560);
or U6633 (N_6633,N_6412,N_6569);
nand U6634 (N_6634,N_6435,N_6553);
and U6635 (N_6635,N_6490,N_6552);
and U6636 (N_6636,N_6598,N_6563);
or U6637 (N_6637,N_6583,N_6596);
nand U6638 (N_6638,N_6473,N_6402);
and U6639 (N_6639,N_6541,N_6550);
nor U6640 (N_6640,N_6485,N_6461);
nand U6641 (N_6641,N_6476,N_6593);
xnor U6642 (N_6642,N_6501,N_6418);
nand U6643 (N_6643,N_6580,N_6439);
or U6644 (N_6644,N_6488,N_6511);
or U6645 (N_6645,N_6423,N_6540);
xor U6646 (N_6646,N_6460,N_6508);
or U6647 (N_6647,N_6582,N_6522);
or U6648 (N_6648,N_6484,N_6459);
and U6649 (N_6649,N_6562,N_6577);
nor U6650 (N_6650,N_6586,N_6437);
or U6651 (N_6651,N_6436,N_6529);
nand U6652 (N_6652,N_6576,N_6441);
xnor U6653 (N_6653,N_6444,N_6520);
nor U6654 (N_6654,N_6470,N_6431);
xnor U6655 (N_6655,N_6536,N_6408);
nor U6656 (N_6656,N_6566,N_6503);
nand U6657 (N_6657,N_6493,N_6455);
or U6658 (N_6658,N_6450,N_6587);
nand U6659 (N_6659,N_6547,N_6494);
nand U6660 (N_6660,N_6578,N_6416);
xnor U6661 (N_6661,N_6526,N_6507);
nand U6662 (N_6662,N_6527,N_6442);
or U6663 (N_6663,N_6573,N_6409);
and U6664 (N_6664,N_6546,N_6554);
nor U6665 (N_6665,N_6570,N_6429);
or U6666 (N_6666,N_6430,N_6438);
xnor U6667 (N_6667,N_6500,N_6532);
or U6668 (N_6668,N_6407,N_6595);
xnor U6669 (N_6669,N_6447,N_6581);
or U6670 (N_6670,N_6495,N_6426);
nand U6671 (N_6671,N_6427,N_6443);
nand U6672 (N_6672,N_6448,N_6514);
xor U6673 (N_6673,N_6469,N_6534);
nor U6674 (N_6674,N_6515,N_6571);
or U6675 (N_6675,N_6420,N_6557);
nor U6676 (N_6676,N_6499,N_6497);
and U6677 (N_6677,N_6404,N_6599);
nor U6678 (N_6678,N_6424,N_6555);
and U6679 (N_6679,N_6463,N_6521);
xnor U6680 (N_6680,N_6446,N_6561);
nand U6681 (N_6681,N_6558,N_6481);
and U6682 (N_6682,N_6589,N_6535);
nand U6683 (N_6683,N_6590,N_6531);
nand U6684 (N_6684,N_6510,N_6467);
nor U6685 (N_6685,N_6453,N_6428);
nor U6686 (N_6686,N_6567,N_6506);
and U6687 (N_6687,N_6468,N_6457);
nor U6688 (N_6688,N_6544,N_6574);
and U6689 (N_6689,N_6509,N_6417);
nand U6690 (N_6690,N_6421,N_6496);
and U6691 (N_6691,N_6513,N_6517);
or U6692 (N_6692,N_6479,N_6565);
nand U6693 (N_6693,N_6462,N_6545);
xor U6694 (N_6694,N_6512,N_6537);
xnor U6695 (N_6695,N_6518,N_6491);
xnor U6696 (N_6696,N_6477,N_6585);
or U6697 (N_6697,N_6592,N_6401);
nand U6698 (N_6698,N_6400,N_6466);
and U6699 (N_6699,N_6542,N_6568);
and U6700 (N_6700,N_6425,N_6548);
nand U6701 (N_6701,N_6542,N_6563);
or U6702 (N_6702,N_6578,N_6556);
nor U6703 (N_6703,N_6513,N_6563);
xor U6704 (N_6704,N_6409,N_6599);
or U6705 (N_6705,N_6455,N_6536);
xor U6706 (N_6706,N_6464,N_6587);
nor U6707 (N_6707,N_6491,N_6586);
xnor U6708 (N_6708,N_6413,N_6571);
nor U6709 (N_6709,N_6411,N_6441);
xnor U6710 (N_6710,N_6460,N_6439);
nand U6711 (N_6711,N_6531,N_6452);
and U6712 (N_6712,N_6436,N_6446);
xor U6713 (N_6713,N_6435,N_6457);
and U6714 (N_6714,N_6571,N_6551);
or U6715 (N_6715,N_6472,N_6475);
and U6716 (N_6716,N_6542,N_6521);
and U6717 (N_6717,N_6483,N_6579);
or U6718 (N_6718,N_6493,N_6523);
and U6719 (N_6719,N_6406,N_6460);
nor U6720 (N_6720,N_6497,N_6417);
and U6721 (N_6721,N_6405,N_6560);
nor U6722 (N_6722,N_6530,N_6459);
or U6723 (N_6723,N_6401,N_6555);
nor U6724 (N_6724,N_6481,N_6429);
nor U6725 (N_6725,N_6441,N_6490);
xor U6726 (N_6726,N_6501,N_6406);
xnor U6727 (N_6727,N_6567,N_6511);
nor U6728 (N_6728,N_6453,N_6403);
or U6729 (N_6729,N_6417,N_6456);
nand U6730 (N_6730,N_6456,N_6548);
xnor U6731 (N_6731,N_6463,N_6433);
nor U6732 (N_6732,N_6557,N_6527);
nand U6733 (N_6733,N_6488,N_6438);
nand U6734 (N_6734,N_6559,N_6457);
and U6735 (N_6735,N_6579,N_6561);
nand U6736 (N_6736,N_6507,N_6560);
nand U6737 (N_6737,N_6435,N_6597);
and U6738 (N_6738,N_6447,N_6414);
xnor U6739 (N_6739,N_6529,N_6432);
and U6740 (N_6740,N_6440,N_6444);
nor U6741 (N_6741,N_6516,N_6407);
nor U6742 (N_6742,N_6498,N_6520);
and U6743 (N_6743,N_6523,N_6459);
nor U6744 (N_6744,N_6428,N_6486);
or U6745 (N_6745,N_6541,N_6478);
xnor U6746 (N_6746,N_6467,N_6533);
xnor U6747 (N_6747,N_6490,N_6497);
or U6748 (N_6748,N_6496,N_6520);
xnor U6749 (N_6749,N_6489,N_6446);
xnor U6750 (N_6750,N_6402,N_6438);
nor U6751 (N_6751,N_6416,N_6525);
or U6752 (N_6752,N_6597,N_6537);
or U6753 (N_6753,N_6447,N_6566);
or U6754 (N_6754,N_6556,N_6427);
or U6755 (N_6755,N_6507,N_6512);
nand U6756 (N_6756,N_6598,N_6526);
and U6757 (N_6757,N_6542,N_6467);
or U6758 (N_6758,N_6492,N_6481);
nand U6759 (N_6759,N_6503,N_6431);
and U6760 (N_6760,N_6533,N_6462);
xor U6761 (N_6761,N_6445,N_6510);
xor U6762 (N_6762,N_6518,N_6413);
nor U6763 (N_6763,N_6436,N_6434);
and U6764 (N_6764,N_6514,N_6547);
nand U6765 (N_6765,N_6497,N_6481);
nand U6766 (N_6766,N_6466,N_6470);
xnor U6767 (N_6767,N_6474,N_6595);
xor U6768 (N_6768,N_6557,N_6435);
nor U6769 (N_6769,N_6578,N_6519);
nand U6770 (N_6770,N_6559,N_6597);
xnor U6771 (N_6771,N_6499,N_6522);
and U6772 (N_6772,N_6502,N_6407);
and U6773 (N_6773,N_6512,N_6562);
xor U6774 (N_6774,N_6575,N_6440);
or U6775 (N_6775,N_6480,N_6548);
nor U6776 (N_6776,N_6499,N_6527);
or U6777 (N_6777,N_6518,N_6568);
nor U6778 (N_6778,N_6413,N_6512);
xnor U6779 (N_6779,N_6512,N_6528);
nor U6780 (N_6780,N_6584,N_6458);
nor U6781 (N_6781,N_6438,N_6523);
xnor U6782 (N_6782,N_6413,N_6412);
and U6783 (N_6783,N_6576,N_6466);
and U6784 (N_6784,N_6488,N_6424);
or U6785 (N_6785,N_6532,N_6592);
and U6786 (N_6786,N_6545,N_6558);
and U6787 (N_6787,N_6520,N_6421);
nand U6788 (N_6788,N_6458,N_6594);
xnor U6789 (N_6789,N_6482,N_6422);
xnor U6790 (N_6790,N_6469,N_6559);
xor U6791 (N_6791,N_6462,N_6472);
or U6792 (N_6792,N_6428,N_6591);
or U6793 (N_6793,N_6431,N_6465);
nor U6794 (N_6794,N_6570,N_6478);
nor U6795 (N_6795,N_6551,N_6580);
and U6796 (N_6796,N_6578,N_6516);
nor U6797 (N_6797,N_6467,N_6505);
nor U6798 (N_6798,N_6452,N_6584);
and U6799 (N_6799,N_6518,N_6532);
nor U6800 (N_6800,N_6657,N_6733);
nor U6801 (N_6801,N_6723,N_6751);
and U6802 (N_6802,N_6650,N_6702);
nor U6803 (N_6803,N_6628,N_6765);
nor U6804 (N_6804,N_6739,N_6799);
xor U6805 (N_6805,N_6688,N_6617);
xnor U6806 (N_6806,N_6687,N_6796);
nand U6807 (N_6807,N_6649,N_6759);
nor U6808 (N_6808,N_6616,N_6745);
and U6809 (N_6809,N_6662,N_6797);
and U6810 (N_6810,N_6760,N_6756);
nand U6811 (N_6811,N_6712,N_6608);
and U6812 (N_6812,N_6707,N_6681);
and U6813 (N_6813,N_6658,N_6684);
nand U6814 (N_6814,N_6782,N_6647);
nor U6815 (N_6815,N_6746,N_6631);
or U6816 (N_6816,N_6655,N_6734);
xnor U6817 (N_6817,N_6675,N_6638);
nand U6818 (N_6818,N_6741,N_6784);
and U6819 (N_6819,N_6632,N_6667);
or U6820 (N_6820,N_6715,N_6742);
nor U6821 (N_6821,N_6641,N_6607);
nor U6822 (N_6822,N_6754,N_6798);
xnor U6823 (N_6823,N_6708,N_6661);
xor U6824 (N_6824,N_6781,N_6749);
nor U6825 (N_6825,N_6753,N_6726);
nand U6826 (N_6826,N_6648,N_6697);
nor U6827 (N_6827,N_6785,N_6652);
nor U6828 (N_6828,N_6772,N_6627);
xor U6829 (N_6829,N_6762,N_6664);
xor U6830 (N_6830,N_6757,N_6716);
nand U6831 (N_6831,N_6724,N_6699);
xor U6832 (N_6832,N_6748,N_6651);
xnor U6833 (N_6833,N_6621,N_6659);
nand U6834 (N_6834,N_6791,N_6710);
and U6835 (N_6835,N_6663,N_6635);
or U6836 (N_6836,N_6686,N_6605);
xnor U6837 (N_6837,N_6705,N_6680);
xnor U6838 (N_6838,N_6611,N_6717);
nor U6839 (N_6839,N_6674,N_6771);
nand U6840 (N_6840,N_6603,N_6630);
xor U6841 (N_6841,N_6792,N_6685);
xnor U6842 (N_6842,N_6747,N_6735);
or U6843 (N_6843,N_6613,N_6618);
and U6844 (N_6844,N_6728,N_6677);
or U6845 (N_6845,N_6768,N_6634);
nand U6846 (N_6846,N_6718,N_6755);
or U6847 (N_6847,N_6633,N_6714);
xor U6848 (N_6848,N_6640,N_6767);
nand U6849 (N_6849,N_6720,N_6642);
xnor U6850 (N_6850,N_6673,N_6614);
nor U6851 (N_6851,N_6601,N_6722);
xnor U6852 (N_6852,N_6622,N_6758);
xnor U6853 (N_6853,N_6615,N_6620);
nor U6854 (N_6854,N_6619,N_6653);
nor U6855 (N_6855,N_6654,N_6743);
nand U6856 (N_6856,N_6610,N_6786);
nor U6857 (N_6857,N_6612,N_6636);
and U6858 (N_6858,N_6692,N_6668);
nand U6859 (N_6859,N_6740,N_6725);
or U6860 (N_6860,N_6670,N_6766);
nor U6861 (N_6861,N_6689,N_6776);
nor U6862 (N_6862,N_6693,N_6721);
nand U6863 (N_6863,N_6671,N_6779);
or U6864 (N_6864,N_6626,N_6676);
nor U6865 (N_6865,N_6698,N_6682);
or U6866 (N_6866,N_6645,N_6625);
and U6867 (N_6867,N_6732,N_6701);
nor U6868 (N_6868,N_6709,N_6623);
or U6869 (N_6869,N_6719,N_6775);
or U6870 (N_6870,N_6790,N_6744);
nand U6871 (N_6871,N_6665,N_6777);
and U6872 (N_6872,N_6644,N_6787);
nand U6873 (N_6873,N_6602,N_6696);
and U6874 (N_6874,N_6700,N_6660);
or U6875 (N_6875,N_6773,N_6624);
nor U6876 (N_6876,N_6761,N_6679);
xnor U6877 (N_6877,N_6704,N_6774);
or U6878 (N_6878,N_6770,N_6783);
nand U6879 (N_6879,N_6637,N_6795);
or U6880 (N_6880,N_6666,N_6794);
nor U6881 (N_6881,N_6727,N_6690);
nand U6882 (N_6882,N_6778,N_6750);
and U6883 (N_6883,N_6646,N_6695);
xnor U6884 (N_6884,N_6793,N_6738);
nor U6885 (N_6885,N_6669,N_6694);
nand U6886 (N_6886,N_6683,N_6606);
and U6887 (N_6887,N_6730,N_6656);
and U6888 (N_6888,N_6609,N_6769);
nor U6889 (N_6889,N_6604,N_6752);
or U6890 (N_6890,N_6789,N_6788);
nand U6891 (N_6891,N_6729,N_6672);
or U6892 (N_6892,N_6639,N_6763);
and U6893 (N_6893,N_6600,N_6736);
or U6894 (N_6894,N_6711,N_6780);
xor U6895 (N_6895,N_6678,N_6703);
and U6896 (N_6896,N_6706,N_6731);
and U6897 (N_6897,N_6691,N_6713);
and U6898 (N_6898,N_6764,N_6629);
nor U6899 (N_6899,N_6737,N_6643);
nor U6900 (N_6900,N_6681,N_6679);
xor U6901 (N_6901,N_6627,N_6662);
and U6902 (N_6902,N_6788,N_6717);
nor U6903 (N_6903,N_6616,N_6767);
nor U6904 (N_6904,N_6623,N_6627);
nor U6905 (N_6905,N_6721,N_6646);
and U6906 (N_6906,N_6774,N_6640);
or U6907 (N_6907,N_6699,N_6777);
xnor U6908 (N_6908,N_6756,N_6687);
or U6909 (N_6909,N_6626,N_6610);
or U6910 (N_6910,N_6702,N_6610);
nor U6911 (N_6911,N_6796,N_6677);
nand U6912 (N_6912,N_6709,N_6696);
and U6913 (N_6913,N_6722,N_6718);
nor U6914 (N_6914,N_6659,N_6736);
nand U6915 (N_6915,N_6746,N_6799);
nor U6916 (N_6916,N_6676,N_6654);
nor U6917 (N_6917,N_6777,N_6728);
nor U6918 (N_6918,N_6633,N_6661);
nand U6919 (N_6919,N_6670,N_6679);
nand U6920 (N_6920,N_6689,N_6649);
or U6921 (N_6921,N_6790,N_6722);
nand U6922 (N_6922,N_6682,N_6794);
xor U6923 (N_6923,N_6693,N_6764);
nand U6924 (N_6924,N_6600,N_6712);
or U6925 (N_6925,N_6653,N_6734);
xor U6926 (N_6926,N_6605,N_6704);
and U6927 (N_6927,N_6723,N_6795);
and U6928 (N_6928,N_6620,N_6781);
xnor U6929 (N_6929,N_6622,N_6791);
and U6930 (N_6930,N_6771,N_6727);
nand U6931 (N_6931,N_6609,N_6797);
or U6932 (N_6932,N_6713,N_6741);
nand U6933 (N_6933,N_6732,N_6753);
xor U6934 (N_6934,N_6650,N_6653);
nand U6935 (N_6935,N_6730,N_6714);
nor U6936 (N_6936,N_6679,N_6684);
and U6937 (N_6937,N_6738,N_6771);
xnor U6938 (N_6938,N_6686,N_6726);
or U6939 (N_6939,N_6656,N_6719);
xnor U6940 (N_6940,N_6630,N_6789);
xnor U6941 (N_6941,N_6665,N_6787);
nor U6942 (N_6942,N_6615,N_6749);
xnor U6943 (N_6943,N_6799,N_6642);
nand U6944 (N_6944,N_6793,N_6715);
or U6945 (N_6945,N_6780,N_6742);
nand U6946 (N_6946,N_6629,N_6757);
and U6947 (N_6947,N_6712,N_6634);
or U6948 (N_6948,N_6791,N_6784);
or U6949 (N_6949,N_6788,N_6644);
nor U6950 (N_6950,N_6625,N_6797);
nand U6951 (N_6951,N_6725,N_6793);
nand U6952 (N_6952,N_6669,N_6701);
or U6953 (N_6953,N_6790,N_6646);
or U6954 (N_6954,N_6752,N_6631);
or U6955 (N_6955,N_6602,N_6725);
xor U6956 (N_6956,N_6772,N_6622);
xnor U6957 (N_6957,N_6761,N_6777);
xor U6958 (N_6958,N_6694,N_6662);
or U6959 (N_6959,N_6677,N_6616);
nand U6960 (N_6960,N_6724,N_6649);
nand U6961 (N_6961,N_6758,N_6713);
or U6962 (N_6962,N_6723,N_6618);
or U6963 (N_6963,N_6776,N_6662);
and U6964 (N_6964,N_6730,N_6695);
nand U6965 (N_6965,N_6734,N_6779);
nor U6966 (N_6966,N_6642,N_6738);
or U6967 (N_6967,N_6649,N_6616);
nor U6968 (N_6968,N_6795,N_6772);
or U6969 (N_6969,N_6728,N_6624);
nand U6970 (N_6970,N_6760,N_6691);
xor U6971 (N_6971,N_6617,N_6672);
nor U6972 (N_6972,N_6723,N_6690);
or U6973 (N_6973,N_6608,N_6698);
nand U6974 (N_6974,N_6770,N_6644);
nand U6975 (N_6975,N_6733,N_6748);
xnor U6976 (N_6976,N_6724,N_6745);
and U6977 (N_6977,N_6743,N_6676);
xnor U6978 (N_6978,N_6772,N_6667);
and U6979 (N_6979,N_6757,N_6670);
nand U6980 (N_6980,N_6678,N_6708);
and U6981 (N_6981,N_6742,N_6702);
or U6982 (N_6982,N_6686,N_6700);
nand U6983 (N_6983,N_6644,N_6696);
and U6984 (N_6984,N_6725,N_6677);
xor U6985 (N_6985,N_6637,N_6653);
nor U6986 (N_6986,N_6749,N_6760);
xnor U6987 (N_6987,N_6612,N_6601);
nor U6988 (N_6988,N_6707,N_6797);
and U6989 (N_6989,N_6617,N_6722);
or U6990 (N_6990,N_6776,N_6744);
nor U6991 (N_6991,N_6607,N_6700);
xnor U6992 (N_6992,N_6604,N_6732);
xor U6993 (N_6993,N_6701,N_6672);
nor U6994 (N_6994,N_6631,N_6729);
nand U6995 (N_6995,N_6757,N_6621);
nor U6996 (N_6996,N_6791,N_6769);
nand U6997 (N_6997,N_6707,N_6720);
and U6998 (N_6998,N_6700,N_6690);
nand U6999 (N_6999,N_6619,N_6723);
nor U7000 (N_7000,N_6908,N_6943);
or U7001 (N_7001,N_6932,N_6935);
and U7002 (N_7002,N_6844,N_6802);
or U7003 (N_7003,N_6832,N_6942);
and U7004 (N_7004,N_6882,N_6886);
or U7005 (N_7005,N_6930,N_6818);
xor U7006 (N_7006,N_6973,N_6907);
nand U7007 (N_7007,N_6968,N_6974);
nand U7008 (N_7008,N_6814,N_6888);
nor U7009 (N_7009,N_6835,N_6890);
or U7010 (N_7010,N_6828,N_6895);
or U7011 (N_7011,N_6813,N_6855);
xnor U7012 (N_7012,N_6846,N_6961);
xor U7013 (N_7013,N_6876,N_6823);
nand U7014 (N_7014,N_6868,N_6898);
nor U7015 (N_7015,N_6880,N_6812);
and U7016 (N_7016,N_6983,N_6904);
and U7017 (N_7017,N_6897,N_6951);
nand U7018 (N_7018,N_6856,N_6808);
nand U7019 (N_7019,N_6970,N_6892);
nand U7020 (N_7020,N_6825,N_6874);
nor U7021 (N_7021,N_6990,N_6857);
and U7022 (N_7022,N_6900,N_6864);
nor U7023 (N_7023,N_6928,N_6944);
and U7024 (N_7024,N_6909,N_6964);
xnor U7025 (N_7025,N_6849,N_6853);
or U7026 (N_7026,N_6946,N_6960);
or U7027 (N_7027,N_6836,N_6877);
and U7028 (N_7028,N_6981,N_6803);
or U7029 (N_7029,N_6972,N_6914);
nand U7030 (N_7030,N_6933,N_6843);
xor U7031 (N_7031,N_6851,N_6881);
xnor U7032 (N_7032,N_6822,N_6854);
xnor U7033 (N_7033,N_6865,N_6919);
and U7034 (N_7034,N_6869,N_6940);
nand U7035 (N_7035,N_6873,N_6826);
nor U7036 (N_7036,N_6924,N_6871);
xor U7037 (N_7037,N_6998,N_6905);
nand U7038 (N_7038,N_6954,N_6986);
nand U7039 (N_7039,N_6840,N_6920);
or U7040 (N_7040,N_6820,N_6947);
xnor U7041 (N_7041,N_6830,N_6827);
and U7042 (N_7042,N_6922,N_6936);
nor U7043 (N_7043,N_6982,N_6884);
nand U7044 (N_7044,N_6941,N_6889);
nor U7045 (N_7045,N_6957,N_6817);
nand U7046 (N_7046,N_6875,N_6956);
nor U7047 (N_7047,N_6848,N_6985);
and U7048 (N_7048,N_6939,N_6952);
xnor U7049 (N_7049,N_6816,N_6883);
nand U7050 (N_7050,N_6979,N_6821);
xor U7051 (N_7051,N_6894,N_6870);
or U7052 (N_7052,N_6804,N_6850);
nand U7053 (N_7053,N_6991,N_6842);
xnor U7054 (N_7054,N_6831,N_6847);
nand U7055 (N_7055,N_6863,N_6980);
and U7056 (N_7056,N_6993,N_6858);
nand U7057 (N_7057,N_6997,N_6915);
nor U7058 (N_7058,N_6971,N_6838);
nand U7059 (N_7059,N_6806,N_6859);
and U7060 (N_7060,N_6934,N_6965);
nand U7061 (N_7061,N_6910,N_6977);
or U7062 (N_7062,N_6837,N_6824);
nor U7063 (N_7063,N_6921,N_6926);
xnor U7064 (N_7064,N_6902,N_6992);
or U7065 (N_7065,N_6862,N_6945);
and U7066 (N_7066,N_6999,N_6962);
nand U7067 (N_7067,N_6931,N_6949);
xor U7068 (N_7068,N_6887,N_6987);
and U7069 (N_7069,N_6903,N_6927);
or U7070 (N_7070,N_6938,N_6805);
and U7071 (N_7071,N_6948,N_6912);
or U7072 (N_7072,N_6872,N_6845);
and U7073 (N_7073,N_6801,N_6807);
nand U7074 (N_7074,N_6811,N_6959);
and U7075 (N_7075,N_6878,N_6815);
or U7076 (N_7076,N_6899,N_6833);
and U7077 (N_7077,N_6913,N_6906);
nand U7078 (N_7078,N_6963,N_6839);
nand U7079 (N_7079,N_6891,N_6867);
nor U7080 (N_7080,N_6879,N_6953);
and U7081 (N_7081,N_6955,N_6969);
xor U7082 (N_7082,N_6809,N_6925);
nor U7083 (N_7083,N_6916,N_6994);
nor U7084 (N_7084,N_6917,N_6988);
nor U7085 (N_7085,N_6901,N_6911);
or U7086 (N_7086,N_6958,N_6885);
xnor U7087 (N_7087,N_6810,N_6841);
nor U7088 (N_7088,N_6918,N_6995);
xor U7089 (N_7089,N_6967,N_6950);
xor U7090 (N_7090,N_6937,N_6800);
nor U7091 (N_7091,N_6866,N_6984);
xnor U7092 (N_7092,N_6975,N_6829);
xnor U7093 (N_7093,N_6989,N_6976);
and U7094 (N_7094,N_6929,N_6819);
nor U7095 (N_7095,N_6966,N_6861);
nor U7096 (N_7096,N_6852,N_6923);
nor U7097 (N_7097,N_6996,N_6896);
nand U7098 (N_7098,N_6893,N_6978);
and U7099 (N_7099,N_6860,N_6834);
nand U7100 (N_7100,N_6925,N_6845);
or U7101 (N_7101,N_6923,N_6837);
nand U7102 (N_7102,N_6882,N_6880);
or U7103 (N_7103,N_6844,N_6872);
and U7104 (N_7104,N_6988,N_6990);
nand U7105 (N_7105,N_6977,N_6840);
nand U7106 (N_7106,N_6911,N_6924);
xnor U7107 (N_7107,N_6859,N_6813);
xnor U7108 (N_7108,N_6927,N_6823);
and U7109 (N_7109,N_6806,N_6974);
xor U7110 (N_7110,N_6857,N_6861);
xnor U7111 (N_7111,N_6971,N_6956);
or U7112 (N_7112,N_6873,N_6879);
or U7113 (N_7113,N_6975,N_6910);
nand U7114 (N_7114,N_6850,N_6960);
xnor U7115 (N_7115,N_6919,N_6991);
nand U7116 (N_7116,N_6969,N_6930);
nand U7117 (N_7117,N_6834,N_6964);
nor U7118 (N_7118,N_6991,N_6802);
nor U7119 (N_7119,N_6944,N_6848);
nor U7120 (N_7120,N_6977,N_6986);
or U7121 (N_7121,N_6981,N_6993);
nor U7122 (N_7122,N_6951,N_6881);
and U7123 (N_7123,N_6939,N_6918);
xor U7124 (N_7124,N_6836,N_6825);
nor U7125 (N_7125,N_6910,N_6805);
nand U7126 (N_7126,N_6947,N_6928);
nor U7127 (N_7127,N_6885,N_6856);
xor U7128 (N_7128,N_6802,N_6821);
xor U7129 (N_7129,N_6976,N_6880);
or U7130 (N_7130,N_6854,N_6954);
xor U7131 (N_7131,N_6943,N_6869);
xor U7132 (N_7132,N_6918,N_6985);
or U7133 (N_7133,N_6820,N_6955);
nand U7134 (N_7134,N_6964,N_6994);
xnor U7135 (N_7135,N_6912,N_6866);
xor U7136 (N_7136,N_6815,N_6860);
nor U7137 (N_7137,N_6869,N_6977);
and U7138 (N_7138,N_6904,N_6839);
nor U7139 (N_7139,N_6971,N_6865);
and U7140 (N_7140,N_6896,N_6999);
nor U7141 (N_7141,N_6802,N_6831);
and U7142 (N_7142,N_6959,N_6898);
nand U7143 (N_7143,N_6898,N_6994);
nor U7144 (N_7144,N_6880,N_6974);
nor U7145 (N_7145,N_6980,N_6829);
and U7146 (N_7146,N_6844,N_6812);
xnor U7147 (N_7147,N_6983,N_6876);
and U7148 (N_7148,N_6901,N_6919);
and U7149 (N_7149,N_6895,N_6919);
and U7150 (N_7150,N_6913,N_6986);
nand U7151 (N_7151,N_6990,N_6925);
nand U7152 (N_7152,N_6801,N_6953);
xor U7153 (N_7153,N_6977,N_6873);
or U7154 (N_7154,N_6985,N_6849);
nor U7155 (N_7155,N_6874,N_6991);
nand U7156 (N_7156,N_6809,N_6957);
nand U7157 (N_7157,N_6967,N_6821);
or U7158 (N_7158,N_6977,N_6865);
nand U7159 (N_7159,N_6893,N_6952);
nand U7160 (N_7160,N_6805,N_6897);
nand U7161 (N_7161,N_6937,N_6964);
or U7162 (N_7162,N_6943,N_6892);
or U7163 (N_7163,N_6945,N_6871);
or U7164 (N_7164,N_6979,N_6922);
and U7165 (N_7165,N_6989,N_6981);
nor U7166 (N_7166,N_6934,N_6919);
and U7167 (N_7167,N_6896,N_6957);
or U7168 (N_7168,N_6891,N_6914);
nand U7169 (N_7169,N_6951,N_6966);
nor U7170 (N_7170,N_6858,N_6950);
and U7171 (N_7171,N_6915,N_6926);
or U7172 (N_7172,N_6879,N_6821);
or U7173 (N_7173,N_6899,N_6944);
or U7174 (N_7174,N_6993,N_6958);
or U7175 (N_7175,N_6825,N_6808);
xor U7176 (N_7176,N_6983,N_6988);
or U7177 (N_7177,N_6874,N_6998);
and U7178 (N_7178,N_6926,N_6938);
nand U7179 (N_7179,N_6847,N_6913);
or U7180 (N_7180,N_6964,N_6873);
and U7181 (N_7181,N_6809,N_6982);
and U7182 (N_7182,N_6883,N_6878);
and U7183 (N_7183,N_6926,N_6858);
xnor U7184 (N_7184,N_6836,N_6968);
nand U7185 (N_7185,N_6822,N_6825);
nor U7186 (N_7186,N_6893,N_6841);
nand U7187 (N_7187,N_6876,N_6841);
nor U7188 (N_7188,N_6802,N_6944);
nand U7189 (N_7189,N_6855,N_6922);
nor U7190 (N_7190,N_6894,N_6966);
or U7191 (N_7191,N_6900,N_6944);
nor U7192 (N_7192,N_6854,N_6967);
and U7193 (N_7193,N_6987,N_6957);
xor U7194 (N_7194,N_6843,N_6900);
xnor U7195 (N_7195,N_6856,N_6932);
nand U7196 (N_7196,N_6993,N_6840);
nand U7197 (N_7197,N_6952,N_6840);
and U7198 (N_7198,N_6816,N_6839);
or U7199 (N_7199,N_6941,N_6817);
xor U7200 (N_7200,N_7033,N_7188);
nor U7201 (N_7201,N_7183,N_7105);
and U7202 (N_7202,N_7161,N_7182);
nand U7203 (N_7203,N_7057,N_7142);
nor U7204 (N_7204,N_7081,N_7041);
and U7205 (N_7205,N_7151,N_7150);
nand U7206 (N_7206,N_7080,N_7038);
xor U7207 (N_7207,N_7186,N_7199);
nor U7208 (N_7208,N_7140,N_7058);
nand U7209 (N_7209,N_7174,N_7021);
nand U7210 (N_7210,N_7144,N_7157);
nor U7211 (N_7211,N_7027,N_7138);
and U7212 (N_7212,N_7035,N_7141);
nand U7213 (N_7213,N_7082,N_7015);
nor U7214 (N_7214,N_7064,N_7034);
or U7215 (N_7215,N_7184,N_7069);
and U7216 (N_7216,N_7098,N_7145);
nand U7217 (N_7217,N_7131,N_7028);
and U7218 (N_7218,N_7167,N_7114);
xor U7219 (N_7219,N_7147,N_7133);
and U7220 (N_7220,N_7165,N_7037);
and U7221 (N_7221,N_7053,N_7120);
xnor U7222 (N_7222,N_7065,N_7036);
nand U7223 (N_7223,N_7198,N_7177);
or U7224 (N_7224,N_7126,N_7139);
nand U7225 (N_7225,N_7024,N_7054);
or U7226 (N_7226,N_7003,N_7005);
or U7227 (N_7227,N_7169,N_7099);
xor U7228 (N_7228,N_7078,N_7159);
nor U7229 (N_7229,N_7012,N_7103);
nor U7230 (N_7230,N_7046,N_7136);
nand U7231 (N_7231,N_7008,N_7000);
and U7232 (N_7232,N_7032,N_7158);
nand U7233 (N_7233,N_7062,N_7152);
nor U7234 (N_7234,N_7134,N_7087);
xor U7235 (N_7235,N_7178,N_7044);
xnor U7236 (N_7236,N_7197,N_7085);
nand U7237 (N_7237,N_7059,N_7102);
and U7238 (N_7238,N_7045,N_7084);
nor U7239 (N_7239,N_7052,N_7164);
nand U7240 (N_7240,N_7115,N_7173);
nand U7241 (N_7241,N_7089,N_7129);
or U7242 (N_7242,N_7043,N_7092);
nand U7243 (N_7243,N_7106,N_7190);
or U7244 (N_7244,N_7018,N_7117);
and U7245 (N_7245,N_7020,N_7125);
xor U7246 (N_7246,N_7193,N_7124);
and U7247 (N_7247,N_7192,N_7181);
nor U7248 (N_7248,N_7088,N_7154);
or U7249 (N_7249,N_7104,N_7191);
nand U7250 (N_7250,N_7042,N_7146);
xnor U7251 (N_7251,N_7055,N_7016);
nand U7252 (N_7252,N_7163,N_7132);
or U7253 (N_7253,N_7073,N_7030);
or U7254 (N_7254,N_7079,N_7072);
xnor U7255 (N_7255,N_7056,N_7155);
nand U7256 (N_7256,N_7090,N_7110);
nor U7257 (N_7257,N_7007,N_7180);
nor U7258 (N_7258,N_7001,N_7091);
nor U7259 (N_7259,N_7060,N_7009);
nand U7260 (N_7260,N_7121,N_7017);
or U7261 (N_7261,N_7113,N_7185);
or U7262 (N_7262,N_7066,N_7168);
and U7263 (N_7263,N_7026,N_7101);
nor U7264 (N_7264,N_7179,N_7112);
or U7265 (N_7265,N_7172,N_7109);
xor U7266 (N_7266,N_7076,N_7040);
and U7267 (N_7267,N_7166,N_7122);
or U7268 (N_7268,N_7135,N_7029);
nand U7269 (N_7269,N_7019,N_7127);
and U7270 (N_7270,N_7097,N_7194);
nor U7271 (N_7271,N_7070,N_7108);
or U7272 (N_7272,N_7077,N_7118);
and U7273 (N_7273,N_7011,N_7086);
nor U7274 (N_7274,N_7075,N_7068);
and U7275 (N_7275,N_7010,N_7196);
nor U7276 (N_7276,N_7187,N_7153);
or U7277 (N_7277,N_7100,N_7130);
xnor U7278 (N_7278,N_7061,N_7049);
or U7279 (N_7279,N_7031,N_7047);
nand U7280 (N_7280,N_7143,N_7048);
nand U7281 (N_7281,N_7002,N_7006);
xor U7282 (N_7282,N_7170,N_7083);
or U7283 (N_7283,N_7175,N_7013);
nand U7284 (N_7284,N_7111,N_7171);
xnor U7285 (N_7285,N_7063,N_7160);
and U7286 (N_7286,N_7039,N_7074);
and U7287 (N_7287,N_7050,N_7123);
xor U7288 (N_7288,N_7119,N_7116);
and U7289 (N_7289,N_7162,N_7095);
nand U7290 (N_7290,N_7094,N_7176);
or U7291 (N_7291,N_7137,N_7051);
or U7292 (N_7292,N_7096,N_7195);
nor U7293 (N_7293,N_7189,N_7071);
nand U7294 (N_7294,N_7149,N_7004);
nand U7295 (N_7295,N_7156,N_7067);
or U7296 (N_7296,N_7093,N_7128);
xor U7297 (N_7297,N_7014,N_7148);
and U7298 (N_7298,N_7023,N_7025);
or U7299 (N_7299,N_7022,N_7107);
nand U7300 (N_7300,N_7031,N_7194);
nor U7301 (N_7301,N_7027,N_7157);
or U7302 (N_7302,N_7105,N_7018);
xor U7303 (N_7303,N_7152,N_7078);
and U7304 (N_7304,N_7109,N_7080);
xnor U7305 (N_7305,N_7158,N_7152);
or U7306 (N_7306,N_7070,N_7085);
or U7307 (N_7307,N_7059,N_7041);
nor U7308 (N_7308,N_7113,N_7164);
nand U7309 (N_7309,N_7031,N_7141);
xor U7310 (N_7310,N_7167,N_7127);
or U7311 (N_7311,N_7178,N_7022);
or U7312 (N_7312,N_7068,N_7198);
and U7313 (N_7313,N_7027,N_7137);
nor U7314 (N_7314,N_7004,N_7168);
nand U7315 (N_7315,N_7070,N_7101);
nand U7316 (N_7316,N_7068,N_7087);
nand U7317 (N_7317,N_7129,N_7111);
nor U7318 (N_7318,N_7025,N_7062);
and U7319 (N_7319,N_7083,N_7019);
and U7320 (N_7320,N_7052,N_7076);
xnor U7321 (N_7321,N_7038,N_7088);
nand U7322 (N_7322,N_7070,N_7136);
nor U7323 (N_7323,N_7069,N_7074);
and U7324 (N_7324,N_7124,N_7137);
nand U7325 (N_7325,N_7081,N_7072);
xnor U7326 (N_7326,N_7147,N_7172);
or U7327 (N_7327,N_7158,N_7094);
nand U7328 (N_7328,N_7111,N_7183);
nand U7329 (N_7329,N_7022,N_7196);
nand U7330 (N_7330,N_7041,N_7060);
and U7331 (N_7331,N_7005,N_7127);
xor U7332 (N_7332,N_7045,N_7074);
nand U7333 (N_7333,N_7111,N_7177);
or U7334 (N_7334,N_7117,N_7186);
nor U7335 (N_7335,N_7105,N_7164);
and U7336 (N_7336,N_7190,N_7103);
or U7337 (N_7337,N_7029,N_7121);
xnor U7338 (N_7338,N_7139,N_7093);
nand U7339 (N_7339,N_7116,N_7067);
xnor U7340 (N_7340,N_7060,N_7138);
xor U7341 (N_7341,N_7152,N_7034);
nand U7342 (N_7342,N_7160,N_7131);
nand U7343 (N_7343,N_7076,N_7069);
and U7344 (N_7344,N_7038,N_7132);
and U7345 (N_7345,N_7090,N_7041);
or U7346 (N_7346,N_7067,N_7163);
or U7347 (N_7347,N_7047,N_7173);
and U7348 (N_7348,N_7166,N_7119);
or U7349 (N_7349,N_7124,N_7153);
xnor U7350 (N_7350,N_7155,N_7043);
nor U7351 (N_7351,N_7094,N_7165);
nor U7352 (N_7352,N_7180,N_7153);
nor U7353 (N_7353,N_7086,N_7198);
nor U7354 (N_7354,N_7051,N_7135);
nand U7355 (N_7355,N_7066,N_7018);
or U7356 (N_7356,N_7062,N_7082);
nand U7357 (N_7357,N_7175,N_7071);
nor U7358 (N_7358,N_7002,N_7140);
or U7359 (N_7359,N_7072,N_7155);
or U7360 (N_7360,N_7051,N_7151);
or U7361 (N_7361,N_7106,N_7178);
xnor U7362 (N_7362,N_7107,N_7019);
nand U7363 (N_7363,N_7185,N_7082);
and U7364 (N_7364,N_7093,N_7145);
or U7365 (N_7365,N_7109,N_7161);
nand U7366 (N_7366,N_7180,N_7102);
or U7367 (N_7367,N_7082,N_7038);
nor U7368 (N_7368,N_7067,N_7084);
nor U7369 (N_7369,N_7059,N_7185);
and U7370 (N_7370,N_7041,N_7113);
nor U7371 (N_7371,N_7080,N_7162);
and U7372 (N_7372,N_7178,N_7063);
and U7373 (N_7373,N_7014,N_7008);
nand U7374 (N_7374,N_7172,N_7022);
and U7375 (N_7375,N_7080,N_7012);
nor U7376 (N_7376,N_7049,N_7110);
nand U7377 (N_7377,N_7020,N_7086);
nand U7378 (N_7378,N_7174,N_7023);
and U7379 (N_7379,N_7044,N_7114);
nand U7380 (N_7380,N_7061,N_7088);
and U7381 (N_7381,N_7140,N_7087);
xnor U7382 (N_7382,N_7020,N_7071);
nor U7383 (N_7383,N_7045,N_7003);
or U7384 (N_7384,N_7169,N_7160);
nor U7385 (N_7385,N_7126,N_7009);
and U7386 (N_7386,N_7112,N_7195);
nand U7387 (N_7387,N_7005,N_7144);
and U7388 (N_7388,N_7001,N_7022);
or U7389 (N_7389,N_7168,N_7056);
xor U7390 (N_7390,N_7025,N_7159);
nor U7391 (N_7391,N_7091,N_7108);
xnor U7392 (N_7392,N_7086,N_7032);
and U7393 (N_7393,N_7185,N_7195);
or U7394 (N_7394,N_7080,N_7196);
nand U7395 (N_7395,N_7093,N_7184);
and U7396 (N_7396,N_7118,N_7008);
nor U7397 (N_7397,N_7199,N_7100);
nand U7398 (N_7398,N_7137,N_7118);
or U7399 (N_7399,N_7145,N_7157);
nand U7400 (N_7400,N_7241,N_7204);
or U7401 (N_7401,N_7356,N_7247);
xnor U7402 (N_7402,N_7390,N_7245);
and U7403 (N_7403,N_7220,N_7304);
and U7404 (N_7404,N_7354,N_7372);
xor U7405 (N_7405,N_7327,N_7377);
xnor U7406 (N_7406,N_7339,N_7328);
nor U7407 (N_7407,N_7225,N_7258);
and U7408 (N_7408,N_7305,N_7342);
xnor U7409 (N_7409,N_7300,N_7265);
nand U7410 (N_7410,N_7209,N_7289);
nand U7411 (N_7411,N_7272,N_7357);
xnor U7412 (N_7412,N_7333,N_7249);
nand U7413 (N_7413,N_7313,N_7279);
and U7414 (N_7414,N_7207,N_7299);
nand U7415 (N_7415,N_7324,N_7373);
or U7416 (N_7416,N_7212,N_7215);
and U7417 (N_7417,N_7365,N_7214);
and U7418 (N_7418,N_7321,N_7332);
xor U7419 (N_7419,N_7283,N_7338);
and U7420 (N_7420,N_7329,N_7281);
xor U7421 (N_7421,N_7227,N_7392);
xnor U7422 (N_7422,N_7246,N_7353);
nor U7423 (N_7423,N_7294,N_7259);
xnor U7424 (N_7424,N_7396,N_7226);
and U7425 (N_7425,N_7287,N_7255);
xor U7426 (N_7426,N_7383,N_7382);
xnor U7427 (N_7427,N_7296,N_7271);
nor U7428 (N_7428,N_7203,N_7317);
and U7429 (N_7429,N_7222,N_7312);
nor U7430 (N_7430,N_7274,N_7376);
and U7431 (N_7431,N_7297,N_7244);
nor U7432 (N_7432,N_7242,N_7253);
and U7433 (N_7433,N_7231,N_7284);
xnor U7434 (N_7434,N_7369,N_7293);
nor U7435 (N_7435,N_7268,N_7266);
and U7436 (N_7436,N_7224,N_7316);
nor U7437 (N_7437,N_7308,N_7387);
or U7438 (N_7438,N_7210,N_7320);
xor U7439 (N_7439,N_7219,N_7366);
xor U7440 (N_7440,N_7334,N_7206);
or U7441 (N_7441,N_7282,N_7398);
or U7442 (N_7442,N_7200,N_7311);
nand U7443 (N_7443,N_7368,N_7309);
nor U7444 (N_7444,N_7236,N_7234);
xnor U7445 (N_7445,N_7323,N_7218);
nand U7446 (N_7446,N_7389,N_7391);
or U7447 (N_7447,N_7348,N_7257);
or U7448 (N_7448,N_7292,N_7388);
xnor U7449 (N_7449,N_7288,N_7330);
or U7450 (N_7450,N_7341,N_7201);
and U7451 (N_7451,N_7270,N_7276);
xor U7452 (N_7452,N_7263,N_7352);
xnor U7453 (N_7453,N_7307,N_7298);
nand U7454 (N_7454,N_7223,N_7326);
and U7455 (N_7455,N_7264,N_7290);
and U7456 (N_7456,N_7250,N_7248);
nand U7457 (N_7457,N_7230,N_7379);
and U7458 (N_7458,N_7331,N_7394);
and U7459 (N_7459,N_7310,N_7256);
or U7460 (N_7460,N_7252,N_7285);
nand U7461 (N_7461,N_7280,N_7397);
and U7462 (N_7462,N_7378,N_7233);
and U7463 (N_7463,N_7343,N_7208);
or U7464 (N_7464,N_7291,N_7375);
or U7465 (N_7465,N_7360,N_7239);
and U7466 (N_7466,N_7277,N_7351);
or U7467 (N_7467,N_7361,N_7371);
and U7468 (N_7468,N_7229,N_7314);
nand U7469 (N_7469,N_7350,N_7337);
or U7470 (N_7470,N_7240,N_7303);
xnor U7471 (N_7471,N_7355,N_7254);
xnor U7472 (N_7472,N_7243,N_7370);
nor U7473 (N_7473,N_7367,N_7381);
nand U7474 (N_7474,N_7217,N_7260);
or U7475 (N_7475,N_7399,N_7349);
xor U7476 (N_7476,N_7295,N_7275);
or U7477 (N_7477,N_7344,N_7267);
and U7478 (N_7478,N_7213,N_7318);
xnor U7479 (N_7479,N_7359,N_7380);
nor U7480 (N_7480,N_7232,N_7335);
or U7481 (N_7481,N_7235,N_7364);
or U7482 (N_7482,N_7319,N_7238);
or U7483 (N_7483,N_7386,N_7322);
nor U7484 (N_7484,N_7385,N_7315);
xor U7485 (N_7485,N_7261,N_7269);
xnor U7486 (N_7486,N_7325,N_7395);
xnor U7487 (N_7487,N_7345,N_7216);
nor U7488 (N_7488,N_7262,N_7384);
nand U7489 (N_7489,N_7346,N_7362);
xnor U7490 (N_7490,N_7302,N_7374);
nor U7491 (N_7491,N_7221,N_7347);
xor U7492 (N_7492,N_7336,N_7273);
nor U7493 (N_7493,N_7251,N_7393);
nor U7494 (N_7494,N_7363,N_7202);
or U7495 (N_7495,N_7211,N_7278);
nand U7496 (N_7496,N_7306,N_7358);
and U7497 (N_7497,N_7228,N_7237);
and U7498 (N_7498,N_7286,N_7340);
nor U7499 (N_7499,N_7301,N_7205);
xnor U7500 (N_7500,N_7343,N_7217);
xor U7501 (N_7501,N_7267,N_7210);
nand U7502 (N_7502,N_7383,N_7290);
nor U7503 (N_7503,N_7279,N_7301);
nand U7504 (N_7504,N_7233,N_7324);
nand U7505 (N_7505,N_7220,N_7360);
xnor U7506 (N_7506,N_7305,N_7364);
or U7507 (N_7507,N_7283,N_7382);
nand U7508 (N_7508,N_7289,N_7269);
xor U7509 (N_7509,N_7385,N_7391);
nand U7510 (N_7510,N_7232,N_7364);
xor U7511 (N_7511,N_7256,N_7284);
nand U7512 (N_7512,N_7292,N_7389);
nor U7513 (N_7513,N_7309,N_7218);
xor U7514 (N_7514,N_7328,N_7358);
xnor U7515 (N_7515,N_7271,N_7255);
xor U7516 (N_7516,N_7201,N_7355);
xnor U7517 (N_7517,N_7276,N_7324);
and U7518 (N_7518,N_7232,N_7382);
nand U7519 (N_7519,N_7261,N_7297);
and U7520 (N_7520,N_7285,N_7352);
and U7521 (N_7521,N_7260,N_7238);
xnor U7522 (N_7522,N_7336,N_7309);
nor U7523 (N_7523,N_7235,N_7282);
or U7524 (N_7524,N_7248,N_7319);
xnor U7525 (N_7525,N_7295,N_7261);
and U7526 (N_7526,N_7275,N_7302);
xnor U7527 (N_7527,N_7213,N_7316);
and U7528 (N_7528,N_7278,N_7294);
nor U7529 (N_7529,N_7200,N_7324);
or U7530 (N_7530,N_7245,N_7392);
and U7531 (N_7531,N_7380,N_7230);
nand U7532 (N_7532,N_7232,N_7381);
or U7533 (N_7533,N_7355,N_7206);
xor U7534 (N_7534,N_7306,N_7391);
xnor U7535 (N_7535,N_7324,N_7307);
nand U7536 (N_7536,N_7355,N_7228);
nor U7537 (N_7537,N_7295,N_7233);
and U7538 (N_7538,N_7218,N_7228);
and U7539 (N_7539,N_7236,N_7360);
and U7540 (N_7540,N_7254,N_7357);
nor U7541 (N_7541,N_7312,N_7226);
xnor U7542 (N_7542,N_7361,N_7342);
and U7543 (N_7543,N_7243,N_7271);
xnor U7544 (N_7544,N_7302,N_7360);
nand U7545 (N_7545,N_7367,N_7307);
and U7546 (N_7546,N_7302,N_7350);
nand U7547 (N_7547,N_7377,N_7227);
or U7548 (N_7548,N_7315,N_7266);
nor U7549 (N_7549,N_7335,N_7276);
or U7550 (N_7550,N_7272,N_7244);
xor U7551 (N_7551,N_7205,N_7293);
xor U7552 (N_7552,N_7337,N_7255);
or U7553 (N_7553,N_7210,N_7340);
nand U7554 (N_7554,N_7214,N_7250);
xnor U7555 (N_7555,N_7271,N_7258);
xor U7556 (N_7556,N_7388,N_7298);
nand U7557 (N_7557,N_7247,N_7289);
nand U7558 (N_7558,N_7351,N_7391);
nor U7559 (N_7559,N_7346,N_7308);
xor U7560 (N_7560,N_7223,N_7267);
xnor U7561 (N_7561,N_7389,N_7311);
xor U7562 (N_7562,N_7370,N_7275);
and U7563 (N_7563,N_7327,N_7312);
xor U7564 (N_7564,N_7354,N_7259);
and U7565 (N_7565,N_7285,N_7241);
and U7566 (N_7566,N_7368,N_7333);
or U7567 (N_7567,N_7353,N_7213);
nand U7568 (N_7568,N_7247,N_7358);
nand U7569 (N_7569,N_7326,N_7262);
nor U7570 (N_7570,N_7291,N_7264);
xnor U7571 (N_7571,N_7259,N_7303);
xor U7572 (N_7572,N_7289,N_7339);
nor U7573 (N_7573,N_7200,N_7341);
and U7574 (N_7574,N_7305,N_7373);
or U7575 (N_7575,N_7233,N_7247);
nand U7576 (N_7576,N_7306,N_7399);
or U7577 (N_7577,N_7324,N_7331);
nor U7578 (N_7578,N_7284,N_7342);
xnor U7579 (N_7579,N_7360,N_7366);
nand U7580 (N_7580,N_7306,N_7225);
nand U7581 (N_7581,N_7375,N_7201);
or U7582 (N_7582,N_7220,N_7278);
nand U7583 (N_7583,N_7369,N_7211);
or U7584 (N_7584,N_7302,N_7306);
nor U7585 (N_7585,N_7305,N_7237);
or U7586 (N_7586,N_7375,N_7357);
nor U7587 (N_7587,N_7292,N_7350);
or U7588 (N_7588,N_7382,N_7314);
nand U7589 (N_7589,N_7209,N_7372);
or U7590 (N_7590,N_7384,N_7382);
xor U7591 (N_7591,N_7208,N_7231);
nand U7592 (N_7592,N_7291,N_7398);
nand U7593 (N_7593,N_7358,N_7322);
or U7594 (N_7594,N_7334,N_7346);
nor U7595 (N_7595,N_7365,N_7213);
xor U7596 (N_7596,N_7201,N_7347);
nor U7597 (N_7597,N_7253,N_7218);
nand U7598 (N_7598,N_7316,N_7246);
xor U7599 (N_7599,N_7234,N_7274);
and U7600 (N_7600,N_7570,N_7452);
and U7601 (N_7601,N_7578,N_7530);
xor U7602 (N_7602,N_7457,N_7552);
nor U7603 (N_7603,N_7463,N_7567);
and U7604 (N_7604,N_7556,N_7403);
nand U7605 (N_7605,N_7467,N_7401);
nor U7606 (N_7606,N_7468,N_7541);
nand U7607 (N_7607,N_7524,N_7559);
nor U7608 (N_7608,N_7532,N_7430);
or U7609 (N_7609,N_7549,N_7590);
xnor U7610 (N_7610,N_7526,N_7425);
or U7611 (N_7611,N_7507,N_7479);
and U7612 (N_7612,N_7472,N_7485);
xnor U7613 (N_7613,N_7565,N_7400);
nor U7614 (N_7614,N_7522,N_7572);
nor U7615 (N_7615,N_7412,N_7505);
or U7616 (N_7616,N_7529,N_7514);
nor U7617 (N_7617,N_7551,N_7455);
and U7618 (N_7618,N_7475,N_7406);
nor U7619 (N_7619,N_7451,N_7482);
xor U7620 (N_7620,N_7435,N_7465);
and U7621 (N_7621,N_7418,N_7486);
nand U7622 (N_7622,N_7594,N_7553);
and U7623 (N_7623,N_7424,N_7518);
and U7624 (N_7624,N_7433,N_7434);
nor U7625 (N_7625,N_7577,N_7423);
nor U7626 (N_7626,N_7404,N_7510);
nor U7627 (N_7627,N_7477,N_7444);
or U7628 (N_7628,N_7422,N_7471);
xor U7629 (N_7629,N_7414,N_7428);
or U7630 (N_7630,N_7473,N_7438);
nand U7631 (N_7631,N_7508,N_7499);
or U7632 (N_7632,N_7536,N_7589);
or U7633 (N_7633,N_7576,N_7421);
xnor U7634 (N_7634,N_7580,N_7408);
and U7635 (N_7635,N_7446,N_7546);
or U7636 (N_7636,N_7597,N_7497);
nor U7637 (N_7637,N_7441,N_7521);
nand U7638 (N_7638,N_7439,N_7448);
nor U7639 (N_7639,N_7450,N_7511);
nor U7640 (N_7640,N_7484,N_7598);
or U7641 (N_7641,N_7466,N_7407);
xnor U7642 (N_7642,N_7456,N_7458);
xor U7643 (N_7643,N_7402,N_7564);
xnor U7644 (N_7644,N_7527,N_7409);
nand U7645 (N_7645,N_7431,N_7550);
and U7646 (N_7646,N_7461,N_7520);
nor U7647 (N_7647,N_7554,N_7493);
nor U7648 (N_7648,N_7437,N_7464);
xnor U7649 (N_7649,N_7506,N_7585);
and U7650 (N_7650,N_7539,N_7442);
and U7651 (N_7651,N_7426,N_7503);
or U7652 (N_7652,N_7574,N_7540);
and U7653 (N_7653,N_7481,N_7583);
xnor U7654 (N_7654,N_7447,N_7413);
nor U7655 (N_7655,N_7538,N_7531);
nand U7656 (N_7656,N_7462,N_7449);
or U7657 (N_7657,N_7525,N_7591);
xor U7658 (N_7658,N_7480,N_7443);
xor U7659 (N_7659,N_7488,N_7533);
nor U7660 (N_7660,N_7557,N_7561);
and U7661 (N_7661,N_7411,N_7483);
xnor U7662 (N_7662,N_7596,N_7560);
nand U7663 (N_7663,N_7592,N_7445);
or U7664 (N_7664,N_7440,N_7500);
xnor U7665 (N_7665,N_7582,N_7573);
nor U7666 (N_7666,N_7568,N_7581);
and U7667 (N_7667,N_7460,N_7545);
or U7668 (N_7668,N_7535,N_7588);
or U7669 (N_7669,N_7586,N_7566);
nand U7670 (N_7670,N_7436,N_7575);
nor U7671 (N_7671,N_7415,N_7593);
nand U7672 (N_7672,N_7512,N_7495);
nand U7673 (N_7673,N_7476,N_7502);
nand U7674 (N_7674,N_7547,N_7478);
nand U7675 (N_7675,N_7490,N_7469);
and U7676 (N_7676,N_7489,N_7416);
xnor U7677 (N_7677,N_7548,N_7509);
and U7678 (N_7678,N_7420,N_7494);
xor U7679 (N_7679,N_7544,N_7519);
xnor U7680 (N_7680,N_7487,N_7579);
nand U7681 (N_7681,N_7537,N_7405);
nand U7682 (N_7682,N_7584,N_7558);
or U7683 (N_7683,N_7474,N_7496);
or U7684 (N_7684,N_7599,N_7595);
xor U7685 (N_7685,N_7513,N_7543);
nor U7686 (N_7686,N_7501,N_7498);
xnor U7687 (N_7687,N_7504,N_7517);
nor U7688 (N_7688,N_7562,N_7571);
nand U7689 (N_7689,N_7470,N_7587);
nand U7690 (N_7690,N_7563,N_7542);
nand U7691 (N_7691,N_7419,N_7516);
or U7692 (N_7692,N_7429,N_7523);
and U7693 (N_7693,N_7427,N_7453);
or U7694 (N_7694,N_7454,N_7417);
or U7695 (N_7695,N_7410,N_7432);
xnor U7696 (N_7696,N_7491,N_7459);
nand U7697 (N_7697,N_7534,N_7555);
or U7698 (N_7698,N_7492,N_7569);
nor U7699 (N_7699,N_7528,N_7515);
xor U7700 (N_7700,N_7582,N_7425);
and U7701 (N_7701,N_7557,N_7401);
nand U7702 (N_7702,N_7521,N_7492);
or U7703 (N_7703,N_7414,N_7418);
or U7704 (N_7704,N_7576,N_7484);
xor U7705 (N_7705,N_7497,N_7456);
and U7706 (N_7706,N_7524,N_7428);
and U7707 (N_7707,N_7448,N_7491);
nand U7708 (N_7708,N_7521,N_7517);
or U7709 (N_7709,N_7579,N_7407);
nand U7710 (N_7710,N_7443,N_7427);
xnor U7711 (N_7711,N_7596,N_7499);
xor U7712 (N_7712,N_7575,N_7535);
and U7713 (N_7713,N_7466,N_7468);
or U7714 (N_7714,N_7488,N_7509);
nand U7715 (N_7715,N_7510,N_7586);
nor U7716 (N_7716,N_7465,N_7471);
and U7717 (N_7717,N_7505,N_7477);
nand U7718 (N_7718,N_7471,N_7584);
or U7719 (N_7719,N_7557,N_7552);
and U7720 (N_7720,N_7597,N_7536);
nor U7721 (N_7721,N_7413,N_7539);
or U7722 (N_7722,N_7426,N_7479);
and U7723 (N_7723,N_7434,N_7474);
nand U7724 (N_7724,N_7435,N_7558);
and U7725 (N_7725,N_7536,N_7566);
nand U7726 (N_7726,N_7506,N_7494);
nor U7727 (N_7727,N_7482,N_7543);
or U7728 (N_7728,N_7585,N_7587);
nor U7729 (N_7729,N_7445,N_7546);
or U7730 (N_7730,N_7485,N_7482);
and U7731 (N_7731,N_7548,N_7572);
xnor U7732 (N_7732,N_7567,N_7432);
or U7733 (N_7733,N_7533,N_7411);
and U7734 (N_7734,N_7586,N_7526);
xnor U7735 (N_7735,N_7526,N_7470);
nor U7736 (N_7736,N_7595,N_7452);
nand U7737 (N_7737,N_7579,N_7590);
and U7738 (N_7738,N_7551,N_7428);
nor U7739 (N_7739,N_7560,N_7514);
and U7740 (N_7740,N_7530,N_7532);
nand U7741 (N_7741,N_7413,N_7452);
or U7742 (N_7742,N_7498,N_7421);
and U7743 (N_7743,N_7561,N_7547);
and U7744 (N_7744,N_7524,N_7508);
and U7745 (N_7745,N_7551,N_7486);
nand U7746 (N_7746,N_7473,N_7421);
xnor U7747 (N_7747,N_7474,N_7467);
nor U7748 (N_7748,N_7414,N_7457);
xnor U7749 (N_7749,N_7496,N_7596);
nand U7750 (N_7750,N_7420,N_7525);
and U7751 (N_7751,N_7523,N_7533);
nor U7752 (N_7752,N_7483,N_7488);
nand U7753 (N_7753,N_7527,N_7569);
xnor U7754 (N_7754,N_7513,N_7554);
and U7755 (N_7755,N_7439,N_7572);
or U7756 (N_7756,N_7580,N_7586);
or U7757 (N_7757,N_7449,N_7416);
or U7758 (N_7758,N_7423,N_7415);
xnor U7759 (N_7759,N_7586,N_7438);
nor U7760 (N_7760,N_7441,N_7572);
nor U7761 (N_7761,N_7411,N_7580);
nor U7762 (N_7762,N_7499,N_7517);
and U7763 (N_7763,N_7539,N_7573);
and U7764 (N_7764,N_7546,N_7419);
nor U7765 (N_7765,N_7416,N_7470);
nand U7766 (N_7766,N_7404,N_7572);
xor U7767 (N_7767,N_7536,N_7434);
xnor U7768 (N_7768,N_7527,N_7561);
xnor U7769 (N_7769,N_7461,N_7578);
nor U7770 (N_7770,N_7584,N_7484);
nand U7771 (N_7771,N_7521,N_7481);
nand U7772 (N_7772,N_7408,N_7577);
xor U7773 (N_7773,N_7482,N_7471);
xor U7774 (N_7774,N_7414,N_7477);
nand U7775 (N_7775,N_7578,N_7586);
or U7776 (N_7776,N_7538,N_7507);
and U7777 (N_7777,N_7524,N_7452);
and U7778 (N_7778,N_7478,N_7488);
and U7779 (N_7779,N_7407,N_7595);
nor U7780 (N_7780,N_7469,N_7509);
and U7781 (N_7781,N_7422,N_7587);
or U7782 (N_7782,N_7466,N_7517);
and U7783 (N_7783,N_7425,N_7400);
nor U7784 (N_7784,N_7434,N_7578);
nor U7785 (N_7785,N_7448,N_7513);
nand U7786 (N_7786,N_7419,N_7529);
nor U7787 (N_7787,N_7434,N_7544);
xor U7788 (N_7788,N_7571,N_7538);
or U7789 (N_7789,N_7435,N_7417);
or U7790 (N_7790,N_7492,N_7413);
nor U7791 (N_7791,N_7442,N_7481);
nor U7792 (N_7792,N_7503,N_7475);
nor U7793 (N_7793,N_7507,N_7401);
nand U7794 (N_7794,N_7488,N_7489);
and U7795 (N_7795,N_7431,N_7422);
or U7796 (N_7796,N_7433,N_7457);
nand U7797 (N_7797,N_7534,N_7585);
nand U7798 (N_7798,N_7588,N_7407);
nor U7799 (N_7799,N_7534,N_7511);
nor U7800 (N_7800,N_7720,N_7759);
or U7801 (N_7801,N_7733,N_7792);
and U7802 (N_7802,N_7724,N_7743);
or U7803 (N_7803,N_7663,N_7612);
nor U7804 (N_7804,N_7646,N_7639);
nor U7805 (N_7805,N_7603,N_7637);
and U7806 (N_7806,N_7633,N_7678);
nand U7807 (N_7807,N_7699,N_7607);
and U7808 (N_7808,N_7734,N_7601);
nor U7809 (N_7809,N_7651,N_7757);
nor U7810 (N_7810,N_7706,N_7708);
and U7811 (N_7811,N_7779,N_7789);
and U7812 (N_7812,N_7608,N_7731);
and U7813 (N_7813,N_7600,N_7751);
xnor U7814 (N_7814,N_7632,N_7655);
xor U7815 (N_7815,N_7658,N_7659);
nand U7816 (N_7816,N_7625,N_7614);
nand U7817 (N_7817,N_7747,N_7719);
nand U7818 (N_7818,N_7705,N_7652);
nand U7819 (N_7819,N_7752,N_7618);
nor U7820 (N_7820,N_7628,N_7643);
nor U7821 (N_7821,N_7764,N_7664);
and U7822 (N_7822,N_7777,N_7716);
and U7823 (N_7823,N_7741,N_7626);
and U7824 (N_7824,N_7799,N_7616);
nor U7825 (N_7825,N_7718,N_7620);
and U7826 (N_7826,N_7797,N_7790);
xor U7827 (N_7827,N_7670,N_7684);
xor U7828 (N_7828,N_7647,N_7700);
xor U7829 (N_7829,N_7665,N_7730);
or U7830 (N_7830,N_7693,N_7673);
xnor U7831 (N_7831,N_7694,N_7770);
or U7832 (N_7832,N_7662,N_7675);
and U7833 (N_7833,N_7640,N_7740);
xnor U7834 (N_7834,N_7713,N_7727);
and U7835 (N_7835,N_7689,N_7763);
and U7836 (N_7836,N_7735,N_7660);
nand U7837 (N_7837,N_7645,N_7692);
or U7838 (N_7838,N_7690,N_7648);
xor U7839 (N_7839,N_7709,N_7602);
or U7840 (N_7840,N_7666,N_7776);
nor U7841 (N_7841,N_7609,N_7787);
xnor U7842 (N_7842,N_7773,N_7712);
or U7843 (N_7843,N_7744,N_7795);
nand U7844 (N_7844,N_7676,N_7615);
nor U7845 (N_7845,N_7624,N_7742);
xor U7846 (N_7846,N_7768,N_7688);
xnor U7847 (N_7847,N_7653,N_7685);
and U7848 (N_7848,N_7736,N_7729);
nand U7849 (N_7849,N_7704,N_7610);
xor U7850 (N_7850,N_7707,N_7630);
nand U7851 (N_7851,N_7657,N_7749);
nor U7852 (N_7852,N_7739,N_7765);
xor U7853 (N_7853,N_7782,N_7635);
xnor U7854 (N_7854,N_7780,N_7754);
xor U7855 (N_7855,N_7769,N_7771);
nand U7856 (N_7856,N_7617,N_7629);
and U7857 (N_7857,N_7737,N_7745);
and U7858 (N_7858,N_7621,N_7654);
xor U7859 (N_7859,N_7756,N_7672);
or U7860 (N_7860,N_7796,N_7669);
and U7861 (N_7861,N_7748,N_7622);
xor U7862 (N_7862,N_7679,N_7717);
or U7863 (N_7863,N_7696,N_7793);
xor U7864 (N_7864,N_7762,N_7686);
nand U7865 (N_7865,N_7746,N_7605);
and U7866 (N_7866,N_7691,N_7604);
xor U7867 (N_7867,N_7683,N_7725);
nand U7868 (N_7868,N_7619,N_7766);
and U7869 (N_7869,N_7650,N_7750);
and U7870 (N_7870,N_7606,N_7671);
xor U7871 (N_7871,N_7634,N_7695);
or U7872 (N_7872,N_7714,N_7698);
xor U7873 (N_7873,N_7775,N_7703);
nor U7874 (N_7874,N_7641,N_7668);
or U7875 (N_7875,N_7761,N_7631);
or U7876 (N_7876,N_7794,N_7656);
xor U7877 (N_7877,N_7627,N_7661);
nand U7878 (N_7878,N_7710,N_7723);
nor U7879 (N_7879,N_7636,N_7774);
or U7880 (N_7880,N_7702,N_7638);
or U7881 (N_7881,N_7791,N_7649);
xnor U7882 (N_7882,N_7785,N_7786);
xnor U7883 (N_7883,N_7611,N_7778);
or U7884 (N_7884,N_7798,N_7728);
and U7885 (N_7885,N_7758,N_7667);
and U7886 (N_7886,N_7755,N_7760);
nand U7887 (N_7887,N_7781,N_7697);
and U7888 (N_7888,N_7623,N_7642);
or U7889 (N_7889,N_7644,N_7732);
nor U7890 (N_7890,N_7767,N_7715);
or U7891 (N_7891,N_7681,N_7701);
or U7892 (N_7892,N_7721,N_7711);
xnor U7893 (N_7893,N_7726,N_7677);
nand U7894 (N_7894,N_7753,N_7687);
xnor U7895 (N_7895,N_7674,N_7613);
or U7896 (N_7896,N_7680,N_7784);
or U7897 (N_7897,N_7772,N_7783);
nand U7898 (N_7898,N_7722,N_7788);
and U7899 (N_7899,N_7738,N_7682);
nor U7900 (N_7900,N_7784,N_7643);
and U7901 (N_7901,N_7744,N_7710);
nand U7902 (N_7902,N_7766,N_7719);
nand U7903 (N_7903,N_7656,N_7797);
xnor U7904 (N_7904,N_7746,N_7652);
nand U7905 (N_7905,N_7709,N_7738);
xnor U7906 (N_7906,N_7691,N_7694);
and U7907 (N_7907,N_7751,N_7745);
nor U7908 (N_7908,N_7663,N_7790);
nand U7909 (N_7909,N_7772,N_7668);
xnor U7910 (N_7910,N_7630,N_7660);
nor U7911 (N_7911,N_7655,N_7609);
nor U7912 (N_7912,N_7760,N_7667);
and U7913 (N_7913,N_7711,N_7661);
nand U7914 (N_7914,N_7710,N_7679);
or U7915 (N_7915,N_7657,N_7714);
nand U7916 (N_7916,N_7749,N_7736);
or U7917 (N_7917,N_7614,N_7754);
xnor U7918 (N_7918,N_7736,N_7647);
nand U7919 (N_7919,N_7705,N_7747);
or U7920 (N_7920,N_7604,N_7638);
nand U7921 (N_7921,N_7724,N_7649);
nor U7922 (N_7922,N_7732,N_7609);
and U7923 (N_7923,N_7606,N_7600);
and U7924 (N_7924,N_7620,N_7701);
xnor U7925 (N_7925,N_7705,N_7690);
xnor U7926 (N_7926,N_7661,N_7710);
or U7927 (N_7927,N_7699,N_7615);
nor U7928 (N_7928,N_7769,N_7693);
and U7929 (N_7929,N_7654,N_7671);
nand U7930 (N_7930,N_7697,N_7714);
xnor U7931 (N_7931,N_7656,N_7662);
nor U7932 (N_7932,N_7610,N_7638);
or U7933 (N_7933,N_7753,N_7673);
nand U7934 (N_7934,N_7697,N_7756);
or U7935 (N_7935,N_7799,N_7674);
and U7936 (N_7936,N_7725,N_7736);
nor U7937 (N_7937,N_7728,N_7738);
or U7938 (N_7938,N_7600,N_7676);
and U7939 (N_7939,N_7633,N_7645);
or U7940 (N_7940,N_7710,N_7609);
nand U7941 (N_7941,N_7785,N_7653);
or U7942 (N_7942,N_7654,N_7658);
xor U7943 (N_7943,N_7604,N_7655);
and U7944 (N_7944,N_7686,N_7656);
nor U7945 (N_7945,N_7640,N_7701);
nor U7946 (N_7946,N_7738,N_7639);
xor U7947 (N_7947,N_7693,N_7715);
xnor U7948 (N_7948,N_7770,N_7673);
and U7949 (N_7949,N_7716,N_7739);
nand U7950 (N_7950,N_7715,N_7620);
nor U7951 (N_7951,N_7668,N_7700);
nor U7952 (N_7952,N_7739,N_7605);
nor U7953 (N_7953,N_7616,N_7755);
nand U7954 (N_7954,N_7714,N_7792);
xnor U7955 (N_7955,N_7739,N_7761);
nor U7956 (N_7956,N_7697,N_7613);
and U7957 (N_7957,N_7618,N_7677);
or U7958 (N_7958,N_7706,N_7731);
nand U7959 (N_7959,N_7611,N_7731);
or U7960 (N_7960,N_7650,N_7715);
nand U7961 (N_7961,N_7620,N_7776);
and U7962 (N_7962,N_7609,N_7678);
nor U7963 (N_7963,N_7644,N_7631);
xnor U7964 (N_7964,N_7720,N_7628);
or U7965 (N_7965,N_7616,N_7700);
nand U7966 (N_7966,N_7676,N_7683);
or U7967 (N_7967,N_7793,N_7695);
or U7968 (N_7968,N_7684,N_7713);
and U7969 (N_7969,N_7659,N_7667);
nand U7970 (N_7970,N_7680,N_7684);
xnor U7971 (N_7971,N_7758,N_7762);
nand U7972 (N_7972,N_7621,N_7750);
nor U7973 (N_7973,N_7678,N_7617);
nor U7974 (N_7974,N_7679,N_7758);
xor U7975 (N_7975,N_7779,N_7727);
or U7976 (N_7976,N_7679,N_7623);
xor U7977 (N_7977,N_7749,N_7672);
or U7978 (N_7978,N_7767,N_7730);
nor U7979 (N_7979,N_7701,N_7784);
nor U7980 (N_7980,N_7747,N_7678);
or U7981 (N_7981,N_7793,N_7682);
xnor U7982 (N_7982,N_7693,N_7742);
and U7983 (N_7983,N_7727,N_7610);
nand U7984 (N_7984,N_7619,N_7775);
or U7985 (N_7985,N_7639,N_7725);
and U7986 (N_7986,N_7783,N_7794);
xor U7987 (N_7987,N_7755,N_7719);
xnor U7988 (N_7988,N_7738,N_7768);
or U7989 (N_7989,N_7782,N_7686);
xnor U7990 (N_7990,N_7793,N_7652);
xnor U7991 (N_7991,N_7731,N_7632);
nor U7992 (N_7992,N_7724,N_7799);
nand U7993 (N_7993,N_7732,N_7651);
nor U7994 (N_7994,N_7697,N_7674);
and U7995 (N_7995,N_7703,N_7660);
nand U7996 (N_7996,N_7799,N_7691);
xor U7997 (N_7997,N_7645,N_7663);
and U7998 (N_7998,N_7773,N_7600);
nand U7999 (N_7999,N_7666,N_7785);
xor U8000 (N_8000,N_7871,N_7832);
xor U8001 (N_8001,N_7951,N_7931);
or U8002 (N_8002,N_7963,N_7894);
and U8003 (N_8003,N_7998,N_7848);
nand U8004 (N_8004,N_7861,N_7926);
and U8005 (N_8005,N_7827,N_7818);
and U8006 (N_8006,N_7888,N_7845);
nand U8007 (N_8007,N_7941,N_7828);
nor U8008 (N_8008,N_7834,N_7810);
nand U8009 (N_8009,N_7809,N_7918);
or U8010 (N_8010,N_7944,N_7911);
nand U8011 (N_8011,N_7876,N_7983);
or U8012 (N_8012,N_7844,N_7856);
nand U8013 (N_8013,N_7982,N_7804);
or U8014 (N_8014,N_7959,N_7936);
and U8015 (N_8015,N_7921,N_7993);
or U8016 (N_8016,N_7900,N_7867);
nor U8017 (N_8017,N_7912,N_7905);
nand U8018 (N_8018,N_7830,N_7873);
nor U8019 (N_8019,N_7831,N_7952);
nor U8020 (N_8020,N_7978,N_7863);
nor U8021 (N_8021,N_7837,N_7977);
xnor U8022 (N_8022,N_7817,N_7899);
or U8023 (N_8023,N_7914,N_7940);
nand U8024 (N_8024,N_7806,N_7891);
and U8025 (N_8025,N_7976,N_7996);
or U8026 (N_8026,N_7821,N_7961);
or U8027 (N_8027,N_7992,N_7955);
nand U8028 (N_8028,N_7934,N_7859);
nand U8029 (N_8029,N_7960,N_7954);
nand U8030 (N_8030,N_7853,N_7864);
xor U8031 (N_8031,N_7924,N_7858);
xnor U8032 (N_8032,N_7917,N_7964);
xor U8033 (N_8033,N_7816,N_7895);
nor U8034 (N_8034,N_7813,N_7836);
xor U8035 (N_8035,N_7915,N_7985);
and U8036 (N_8036,N_7820,N_7957);
or U8037 (N_8037,N_7865,N_7807);
and U8038 (N_8038,N_7969,N_7984);
nor U8039 (N_8039,N_7814,N_7930);
nor U8040 (N_8040,N_7842,N_7889);
or U8041 (N_8041,N_7851,N_7862);
nor U8042 (N_8042,N_7805,N_7822);
nand U8043 (N_8043,N_7800,N_7945);
xnor U8044 (N_8044,N_7972,N_7875);
nor U8045 (N_8045,N_7995,N_7947);
nand U8046 (N_8046,N_7812,N_7970);
and U8047 (N_8047,N_7843,N_7835);
nand U8048 (N_8048,N_7950,N_7896);
xnor U8049 (N_8049,N_7932,N_7923);
nand U8050 (N_8050,N_7901,N_7823);
xor U8051 (N_8051,N_7883,N_7933);
nor U8052 (N_8052,N_7819,N_7973);
xor U8053 (N_8053,N_7815,N_7987);
and U8054 (N_8054,N_7904,N_7881);
nor U8055 (N_8055,N_7868,N_7927);
nand U8056 (N_8056,N_7946,N_7880);
nor U8057 (N_8057,N_7890,N_7850);
nor U8058 (N_8058,N_7878,N_7886);
xnor U8059 (N_8059,N_7965,N_7884);
nor U8060 (N_8060,N_7903,N_7866);
nand U8061 (N_8061,N_7909,N_7980);
xnor U8062 (N_8062,N_7919,N_7989);
and U8063 (N_8063,N_7833,N_7887);
and U8064 (N_8064,N_7879,N_7847);
or U8065 (N_8065,N_7824,N_7852);
or U8066 (N_8066,N_7801,N_7898);
nor U8067 (N_8067,N_7966,N_7829);
or U8068 (N_8068,N_7808,N_7962);
or U8069 (N_8069,N_7874,N_7907);
xor U8070 (N_8070,N_7953,N_7988);
nor U8071 (N_8071,N_7803,N_7839);
xnor U8072 (N_8072,N_7811,N_7975);
nand U8073 (N_8073,N_7929,N_7882);
or U8074 (N_8074,N_7892,N_7870);
or U8075 (N_8075,N_7956,N_7916);
and U8076 (N_8076,N_7877,N_7981);
or U8077 (N_8077,N_7872,N_7840);
or U8078 (N_8078,N_7854,N_7857);
and U8079 (N_8079,N_7860,N_7999);
xor U8080 (N_8080,N_7910,N_7968);
or U8081 (N_8081,N_7974,N_7920);
and U8082 (N_8082,N_7825,N_7826);
nor U8083 (N_8083,N_7846,N_7958);
xnor U8084 (N_8084,N_7885,N_7928);
nand U8085 (N_8085,N_7942,N_7948);
or U8086 (N_8086,N_7849,N_7925);
or U8087 (N_8087,N_7971,N_7935);
or U8088 (N_8088,N_7841,N_7838);
and U8089 (N_8089,N_7949,N_7937);
nor U8090 (N_8090,N_7938,N_7997);
xnor U8091 (N_8091,N_7943,N_7994);
nand U8092 (N_8092,N_7897,N_7802);
xnor U8093 (N_8093,N_7990,N_7979);
nand U8094 (N_8094,N_7967,N_7906);
nand U8095 (N_8095,N_7939,N_7902);
and U8096 (N_8096,N_7986,N_7869);
and U8097 (N_8097,N_7913,N_7991);
and U8098 (N_8098,N_7855,N_7893);
nand U8099 (N_8099,N_7922,N_7908);
or U8100 (N_8100,N_7822,N_7945);
nand U8101 (N_8101,N_7872,N_7967);
nand U8102 (N_8102,N_7961,N_7893);
and U8103 (N_8103,N_7900,N_7973);
nor U8104 (N_8104,N_7809,N_7853);
or U8105 (N_8105,N_7835,N_7966);
nand U8106 (N_8106,N_7988,N_7968);
and U8107 (N_8107,N_7871,N_7990);
nand U8108 (N_8108,N_7808,N_7925);
or U8109 (N_8109,N_7998,N_7974);
nand U8110 (N_8110,N_7876,N_7877);
and U8111 (N_8111,N_7969,N_7958);
xnor U8112 (N_8112,N_7927,N_7970);
and U8113 (N_8113,N_7992,N_7968);
nand U8114 (N_8114,N_7831,N_7950);
nand U8115 (N_8115,N_7993,N_7900);
nor U8116 (N_8116,N_7807,N_7864);
xor U8117 (N_8117,N_7929,N_7928);
or U8118 (N_8118,N_7917,N_7952);
nor U8119 (N_8119,N_7998,N_7900);
nor U8120 (N_8120,N_7840,N_7800);
nand U8121 (N_8121,N_7981,N_7940);
or U8122 (N_8122,N_7992,N_7970);
xor U8123 (N_8123,N_7941,N_7976);
nand U8124 (N_8124,N_7924,N_7893);
or U8125 (N_8125,N_7906,N_7894);
and U8126 (N_8126,N_7898,N_7969);
and U8127 (N_8127,N_7855,N_7901);
and U8128 (N_8128,N_7857,N_7826);
and U8129 (N_8129,N_7857,N_7824);
and U8130 (N_8130,N_7896,N_7901);
nor U8131 (N_8131,N_7953,N_7926);
nand U8132 (N_8132,N_7859,N_7995);
nand U8133 (N_8133,N_7878,N_7833);
nand U8134 (N_8134,N_7833,N_7877);
xor U8135 (N_8135,N_7961,N_7813);
and U8136 (N_8136,N_7978,N_7892);
nor U8137 (N_8137,N_7995,N_7887);
xnor U8138 (N_8138,N_7882,N_7873);
nand U8139 (N_8139,N_7979,N_7837);
nand U8140 (N_8140,N_7801,N_7936);
xor U8141 (N_8141,N_7950,N_7952);
and U8142 (N_8142,N_7986,N_7987);
and U8143 (N_8143,N_7968,N_7999);
or U8144 (N_8144,N_7953,N_7848);
or U8145 (N_8145,N_7968,N_7912);
or U8146 (N_8146,N_7992,N_7890);
nand U8147 (N_8147,N_7818,N_7803);
or U8148 (N_8148,N_7985,N_7823);
nor U8149 (N_8149,N_7812,N_7901);
nor U8150 (N_8150,N_7826,N_7967);
and U8151 (N_8151,N_7891,N_7818);
nand U8152 (N_8152,N_7919,N_7813);
nor U8153 (N_8153,N_7864,N_7898);
or U8154 (N_8154,N_7836,N_7889);
xnor U8155 (N_8155,N_7850,N_7901);
nor U8156 (N_8156,N_7891,N_7999);
and U8157 (N_8157,N_7929,N_7998);
nand U8158 (N_8158,N_7931,N_7882);
xnor U8159 (N_8159,N_7881,N_7820);
nand U8160 (N_8160,N_7935,N_7929);
xor U8161 (N_8161,N_7811,N_7889);
nor U8162 (N_8162,N_7863,N_7942);
and U8163 (N_8163,N_7864,N_7892);
nand U8164 (N_8164,N_7946,N_7918);
nand U8165 (N_8165,N_7932,N_7805);
and U8166 (N_8166,N_7974,N_7990);
xor U8167 (N_8167,N_7957,N_7942);
xnor U8168 (N_8168,N_7825,N_7814);
and U8169 (N_8169,N_7898,N_7845);
nand U8170 (N_8170,N_7897,N_7916);
nand U8171 (N_8171,N_7802,N_7893);
xor U8172 (N_8172,N_7962,N_7908);
xnor U8173 (N_8173,N_7893,N_7878);
and U8174 (N_8174,N_7974,N_7897);
nor U8175 (N_8175,N_7999,N_7959);
xor U8176 (N_8176,N_7811,N_7862);
or U8177 (N_8177,N_7914,N_7899);
nand U8178 (N_8178,N_7861,N_7822);
nand U8179 (N_8179,N_7831,N_7917);
nand U8180 (N_8180,N_7971,N_7932);
xor U8181 (N_8181,N_7803,N_7978);
nor U8182 (N_8182,N_7911,N_7848);
xor U8183 (N_8183,N_7841,N_7899);
nand U8184 (N_8184,N_7935,N_7995);
or U8185 (N_8185,N_7821,N_7931);
and U8186 (N_8186,N_7999,N_7950);
nor U8187 (N_8187,N_7866,N_7963);
nor U8188 (N_8188,N_7988,N_7803);
and U8189 (N_8189,N_7835,N_7804);
nor U8190 (N_8190,N_7976,N_7914);
nor U8191 (N_8191,N_7920,N_7993);
or U8192 (N_8192,N_7959,N_7848);
or U8193 (N_8193,N_7963,N_7868);
xnor U8194 (N_8194,N_7915,N_7839);
xor U8195 (N_8195,N_7916,N_7963);
nor U8196 (N_8196,N_7882,N_7828);
and U8197 (N_8197,N_7958,N_7861);
nor U8198 (N_8198,N_7822,N_7887);
nand U8199 (N_8199,N_7866,N_7853);
nand U8200 (N_8200,N_8058,N_8003);
and U8201 (N_8201,N_8054,N_8066);
and U8202 (N_8202,N_8132,N_8126);
nand U8203 (N_8203,N_8074,N_8043);
xnor U8204 (N_8204,N_8124,N_8158);
nand U8205 (N_8205,N_8071,N_8161);
or U8206 (N_8206,N_8045,N_8186);
or U8207 (N_8207,N_8151,N_8052);
nor U8208 (N_8208,N_8051,N_8187);
xnor U8209 (N_8209,N_8137,N_8025);
xnor U8210 (N_8210,N_8024,N_8094);
xor U8211 (N_8211,N_8072,N_8114);
nor U8212 (N_8212,N_8033,N_8093);
and U8213 (N_8213,N_8073,N_8050);
xnor U8214 (N_8214,N_8148,N_8039);
nand U8215 (N_8215,N_8133,N_8192);
nor U8216 (N_8216,N_8145,N_8027);
nor U8217 (N_8217,N_8057,N_8170);
xor U8218 (N_8218,N_8061,N_8163);
and U8219 (N_8219,N_8108,N_8087);
or U8220 (N_8220,N_8085,N_8152);
nand U8221 (N_8221,N_8125,N_8078);
and U8222 (N_8222,N_8171,N_8041);
nor U8223 (N_8223,N_8008,N_8032);
nand U8224 (N_8224,N_8119,N_8062);
nor U8225 (N_8225,N_8035,N_8101);
xor U8226 (N_8226,N_8079,N_8194);
nor U8227 (N_8227,N_8029,N_8009);
xnor U8228 (N_8228,N_8019,N_8026);
xor U8229 (N_8229,N_8042,N_8056);
nor U8230 (N_8230,N_8000,N_8038);
xnor U8231 (N_8231,N_8179,N_8030);
or U8232 (N_8232,N_8060,N_8135);
xnor U8233 (N_8233,N_8011,N_8083);
xor U8234 (N_8234,N_8034,N_8165);
nand U8235 (N_8235,N_8059,N_8031);
or U8236 (N_8236,N_8118,N_8105);
or U8237 (N_8237,N_8096,N_8067);
nor U8238 (N_8238,N_8064,N_8107);
xnor U8239 (N_8239,N_8013,N_8082);
nor U8240 (N_8240,N_8015,N_8049);
nor U8241 (N_8241,N_8070,N_8053);
nand U8242 (N_8242,N_8127,N_8117);
nand U8243 (N_8243,N_8182,N_8189);
or U8244 (N_8244,N_8111,N_8097);
nor U8245 (N_8245,N_8121,N_8084);
xnor U8246 (N_8246,N_8017,N_8153);
xnor U8247 (N_8247,N_8142,N_8081);
nor U8248 (N_8248,N_8103,N_8007);
nor U8249 (N_8249,N_8088,N_8065);
nand U8250 (N_8250,N_8167,N_8014);
or U8251 (N_8251,N_8131,N_8147);
xnor U8252 (N_8252,N_8091,N_8173);
or U8253 (N_8253,N_8004,N_8010);
and U8254 (N_8254,N_8149,N_8089);
nor U8255 (N_8255,N_8047,N_8068);
nor U8256 (N_8256,N_8143,N_8018);
and U8257 (N_8257,N_8016,N_8184);
xor U8258 (N_8258,N_8168,N_8012);
or U8259 (N_8259,N_8037,N_8005);
nand U8260 (N_8260,N_8198,N_8176);
nand U8261 (N_8261,N_8048,N_8040);
or U8262 (N_8262,N_8075,N_8046);
nand U8263 (N_8263,N_8191,N_8138);
nor U8264 (N_8264,N_8196,N_8112);
nand U8265 (N_8265,N_8095,N_8110);
nand U8266 (N_8266,N_8104,N_8020);
or U8267 (N_8267,N_8130,N_8139);
nand U8268 (N_8268,N_8174,N_8063);
and U8269 (N_8269,N_8092,N_8156);
or U8270 (N_8270,N_8193,N_8006);
or U8271 (N_8271,N_8023,N_8159);
nand U8272 (N_8272,N_8106,N_8122);
xor U8273 (N_8273,N_8120,N_8141);
and U8274 (N_8274,N_8188,N_8195);
and U8275 (N_8275,N_8144,N_8166);
nor U8276 (N_8276,N_8100,N_8164);
and U8277 (N_8277,N_8022,N_8146);
or U8278 (N_8278,N_8197,N_8183);
nor U8279 (N_8279,N_8177,N_8116);
and U8280 (N_8280,N_8113,N_8134);
xor U8281 (N_8281,N_8109,N_8128);
nor U8282 (N_8282,N_8178,N_8199);
and U8283 (N_8283,N_8140,N_8080);
and U8284 (N_8284,N_8077,N_8123);
xor U8285 (N_8285,N_8028,N_8169);
and U8286 (N_8286,N_8172,N_8154);
nand U8287 (N_8287,N_8160,N_8102);
and U8288 (N_8288,N_8021,N_8175);
xnor U8289 (N_8289,N_8099,N_8001);
nor U8290 (N_8290,N_8086,N_8044);
nor U8291 (N_8291,N_8162,N_8185);
xor U8292 (N_8292,N_8129,N_8069);
xnor U8293 (N_8293,N_8076,N_8181);
and U8294 (N_8294,N_8090,N_8036);
xnor U8295 (N_8295,N_8098,N_8002);
and U8296 (N_8296,N_8136,N_8190);
or U8297 (N_8297,N_8115,N_8155);
xnor U8298 (N_8298,N_8180,N_8157);
xor U8299 (N_8299,N_8055,N_8150);
nor U8300 (N_8300,N_8125,N_8031);
or U8301 (N_8301,N_8152,N_8022);
and U8302 (N_8302,N_8118,N_8141);
nor U8303 (N_8303,N_8095,N_8041);
xnor U8304 (N_8304,N_8164,N_8114);
or U8305 (N_8305,N_8040,N_8078);
and U8306 (N_8306,N_8173,N_8088);
nor U8307 (N_8307,N_8121,N_8012);
xnor U8308 (N_8308,N_8053,N_8164);
nor U8309 (N_8309,N_8041,N_8188);
nand U8310 (N_8310,N_8075,N_8065);
xnor U8311 (N_8311,N_8122,N_8173);
or U8312 (N_8312,N_8049,N_8181);
xor U8313 (N_8313,N_8136,N_8057);
nand U8314 (N_8314,N_8083,N_8050);
nor U8315 (N_8315,N_8139,N_8105);
or U8316 (N_8316,N_8146,N_8031);
xnor U8317 (N_8317,N_8122,N_8035);
nor U8318 (N_8318,N_8025,N_8099);
nand U8319 (N_8319,N_8114,N_8119);
and U8320 (N_8320,N_8027,N_8013);
xor U8321 (N_8321,N_8150,N_8186);
nand U8322 (N_8322,N_8104,N_8158);
nand U8323 (N_8323,N_8020,N_8030);
and U8324 (N_8324,N_8051,N_8033);
or U8325 (N_8325,N_8024,N_8025);
nand U8326 (N_8326,N_8068,N_8077);
or U8327 (N_8327,N_8176,N_8061);
or U8328 (N_8328,N_8098,N_8119);
xor U8329 (N_8329,N_8080,N_8177);
nand U8330 (N_8330,N_8192,N_8198);
or U8331 (N_8331,N_8130,N_8022);
or U8332 (N_8332,N_8089,N_8016);
xor U8333 (N_8333,N_8001,N_8110);
or U8334 (N_8334,N_8049,N_8190);
xor U8335 (N_8335,N_8177,N_8141);
and U8336 (N_8336,N_8185,N_8055);
xnor U8337 (N_8337,N_8194,N_8131);
nand U8338 (N_8338,N_8084,N_8073);
nand U8339 (N_8339,N_8060,N_8103);
nor U8340 (N_8340,N_8142,N_8132);
xnor U8341 (N_8341,N_8105,N_8087);
xor U8342 (N_8342,N_8183,N_8114);
nor U8343 (N_8343,N_8090,N_8078);
xnor U8344 (N_8344,N_8056,N_8068);
nor U8345 (N_8345,N_8066,N_8183);
nand U8346 (N_8346,N_8020,N_8058);
nand U8347 (N_8347,N_8111,N_8100);
xor U8348 (N_8348,N_8175,N_8103);
nand U8349 (N_8349,N_8057,N_8116);
xnor U8350 (N_8350,N_8102,N_8149);
nor U8351 (N_8351,N_8131,N_8197);
nand U8352 (N_8352,N_8099,N_8029);
or U8353 (N_8353,N_8133,N_8149);
and U8354 (N_8354,N_8128,N_8075);
or U8355 (N_8355,N_8042,N_8125);
nor U8356 (N_8356,N_8032,N_8095);
nand U8357 (N_8357,N_8183,N_8173);
nand U8358 (N_8358,N_8147,N_8084);
and U8359 (N_8359,N_8006,N_8074);
and U8360 (N_8360,N_8098,N_8021);
and U8361 (N_8361,N_8031,N_8194);
nor U8362 (N_8362,N_8062,N_8163);
nor U8363 (N_8363,N_8195,N_8077);
or U8364 (N_8364,N_8135,N_8167);
and U8365 (N_8365,N_8194,N_8119);
or U8366 (N_8366,N_8011,N_8136);
xor U8367 (N_8367,N_8181,N_8158);
xor U8368 (N_8368,N_8135,N_8081);
nor U8369 (N_8369,N_8194,N_8029);
or U8370 (N_8370,N_8110,N_8054);
nand U8371 (N_8371,N_8167,N_8093);
and U8372 (N_8372,N_8153,N_8085);
nand U8373 (N_8373,N_8072,N_8018);
nand U8374 (N_8374,N_8109,N_8047);
nor U8375 (N_8375,N_8070,N_8057);
or U8376 (N_8376,N_8081,N_8195);
nor U8377 (N_8377,N_8027,N_8098);
nand U8378 (N_8378,N_8172,N_8185);
and U8379 (N_8379,N_8033,N_8198);
or U8380 (N_8380,N_8044,N_8149);
nor U8381 (N_8381,N_8195,N_8068);
or U8382 (N_8382,N_8146,N_8108);
and U8383 (N_8383,N_8161,N_8099);
or U8384 (N_8384,N_8052,N_8118);
nor U8385 (N_8385,N_8004,N_8183);
or U8386 (N_8386,N_8018,N_8181);
or U8387 (N_8387,N_8058,N_8061);
or U8388 (N_8388,N_8031,N_8171);
nand U8389 (N_8389,N_8145,N_8063);
nand U8390 (N_8390,N_8017,N_8025);
xor U8391 (N_8391,N_8196,N_8109);
or U8392 (N_8392,N_8098,N_8062);
nand U8393 (N_8393,N_8159,N_8018);
or U8394 (N_8394,N_8008,N_8001);
nand U8395 (N_8395,N_8082,N_8072);
xor U8396 (N_8396,N_8187,N_8181);
and U8397 (N_8397,N_8068,N_8105);
nand U8398 (N_8398,N_8154,N_8115);
nand U8399 (N_8399,N_8022,N_8123);
nand U8400 (N_8400,N_8278,N_8333);
or U8401 (N_8401,N_8318,N_8398);
nand U8402 (N_8402,N_8277,N_8220);
or U8403 (N_8403,N_8250,N_8249);
nor U8404 (N_8404,N_8326,N_8216);
xnor U8405 (N_8405,N_8205,N_8311);
or U8406 (N_8406,N_8351,N_8359);
or U8407 (N_8407,N_8372,N_8337);
xor U8408 (N_8408,N_8236,N_8252);
and U8409 (N_8409,N_8273,N_8322);
and U8410 (N_8410,N_8212,N_8263);
or U8411 (N_8411,N_8226,N_8234);
xnor U8412 (N_8412,N_8284,N_8366);
or U8413 (N_8413,N_8339,N_8321);
nor U8414 (N_8414,N_8374,N_8268);
and U8415 (N_8415,N_8244,N_8243);
xnor U8416 (N_8416,N_8315,N_8264);
xnor U8417 (N_8417,N_8207,N_8358);
and U8418 (N_8418,N_8383,N_8300);
nand U8419 (N_8419,N_8390,N_8281);
xnor U8420 (N_8420,N_8309,N_8221);
nor U8421 (N_8421,N_8200,N_8202);
nand U8422 (N_8422,N_8285,N_8320);
nor U8423 (N_8423,N_8265,N_8381);
and U8424 (N_8424,N_8299,N_8267);
xor U8425 (N_8425,N_8266,N_8363);
xor U8426 (N_8426,N_8314,N_8257);
or U8427 (N_8427,N_8334,N_8251);
or U8428 (N_8428,N_8338,N_8356);
nand U8429 (N_8429,N_8229,N_8335);
xnor U8430 (N_8430,N_8203,N_8352);
or U8431 (N_8431,N_8384,N_8382);
or U8432 (N_8432,N_8237,N_8349);
or U8433 (N_8433,N_8376,N_8293);
and U8434 (N_8434,N_8368,N_8310);
and U8435 (N_8435,N_8369,N_8396);
or U8436 (N_8436,N_8253,N_8294);
and U8437 (N_8437,N_8217,N_8282);
and U8438 (N_8438,N_8354,N_8258);
nand U8439 (N_8439,N_8271,N_8370);
xor U8440 (N_8440,N_8213,N_8204);
xor U8441 (N_8441,N_8377,N_8323);
and U8442 (N_8442,N_8317,N_8331);
or U8443 (N_8443,N_8342,N_8329);
nand U8444 (N_8444,N_8245,N_8241);
xor U8445 (N_8445,N_8242,N_8259);
nor U8446 (N_8446,N_8324,N_8288);
nor U8447 (N_8447,N_8301,N_8228);
and U8448 (N_8448,N_8392,N_8319);
or U8449 (N_8449,N_8270,N_8256);
nor U8450 (N_8450,N_8308,N_8227);
xnor U8451 (N_8451,N_8223,N_8387);
xor U8452 (N_8452,N_8378,N_8214);
nor U8453 (N_8453,N_8313,N_8375);
nand U8454 (N_8454,N_8208,N_8344);
and U8455 (N_8455,N_8373,N_8275);
nand U8456 (N_8456,N_8395,N_8232);
nand U8457 (N_8457,N_8303,N_8312);
nor U8458 (N_8458,N_8291,N_8283);
or U8459 (N_8459,N_8385,N_8371);
nor U8460 (N_8460,N_8348,N_8260);
xnor U8461 (N_8461,N_8238,N_8388);
or U8462 (N_8462,N_8287,N_8389);
or U8463 (N_8463,N_8233,N_8350);
nor U8464 (N_8464,N_8231,N_8330);
and U8465 (N_8465,N_8347,N_8296);
and U8466 (N_8466,N_8279,N_8362);
nor U8467 (N_8467,N_8316,N_8379);
nand U8468 (N_8468,N_8255,N_8248);
nand U8469 (N_8469,N_8261,N_8399);
nor U8470 (N_8470,N_8391,N_8292);
or U8471 (N_8471,N_8295,N_8346);
and U8472 (N_8472,N_8218,N_8235);
and U8473 (N_8473,N_8201,N_8225);
and U8474 (N_8474,N_8355,N_8336);
nand U8475 (N_8475,N_8290,N_8345);
and U8476 (N_8476,N_8397,N_8274);
xor U8477 (N_8477,N_8247,N_8210);
and U8478 (N_8478,N_8304,N_8340);
nand U8479 (N_8479,N_8215,N_8298);
or U8480 (N_8480,N_8219,N_8367);
or U8481 (N_8481,N_8280,N_8286);
nand U8482 (N_8482,N_8246,N_8297);
and U8483 (N_8483,N_8305,N_8341);
nand U8484 (N_8484,N_8254,N_8240);
xor U8485 (N_8485,N_8272,N_8209);
nand U8486 (N_8486,N_8307,N_8325);
xnor U8487 (N_8487,N_8364,N_8386);
nor U8488 (N_8488,N_8230,N_8211);
xor U8489 (N_8489,N_8327,N_8206);
nand U8490 (N_8490,N_8224,N_8262);
nor U8491 (N_8491,N_8380,N_8306);
xor U8492 (N_8492,N_8357,N_8394);
xor U8493 (N_8493,N_8343,N_8302);
nand U8494 (N_8494,N_8332,N_8269);
xor U8495 (N_8495,N_8353,N_8361);
xnor U8496 (N_8496,N_8289,N_8393);
or U8497 (N_8497,N_8360,N_8276);
xor U8498 (N_8498,N_8365,N_8222);
or U8499 (N_8499,N_8239,N_8328);
or U8500 (N_8500,N_8345,N_8217);
or U8501 (N_8501,N_8271,N_8303);
xnor U8502 (N_8502,N_8209,N_8268);
and U8503 (N_8503,N_8364,N_8323);
and U8504 (N_8504,N_8275,N_8394);
xnor U8505 (N_8505,N_8315,N_8292);
xnor U8506 (N_8506,N_8256,N_8346);
nor U8507 (N_8507,N_8351,N_8376);
or U8508 (N_8508,N_8249,N_8240);
or U8509 (N_8509,N_8346,N_8282);
nand U8510 (N_8510,N_8281,N_8209);
nor U8511 (N_8511,N_8210,N_8331);
nor U8512 (N_8512,N_8398,N_8265);
nor U8513 (N_8513,N_8217,N_8386);
xor U8514 (N_8514,N_8377,N_8249);
and U8515 (N_8515,N_8251,N_8352);
nand U8516 (N_8516,N_8256,N_8357);
nand U8517 (N_8517,N_8326,N_8354);
nand U8518 (N_8518,N_8377,N_8356);
nand U8519 (N_8519,N_8367,N_8350);
or U8520 (N_8520,N_8235,N_8300);
or U8521 (N_8521,N_8287,N_8266);
nand U8522 (N_8522,N_8398,N_8235);
and U8523 (N_8523,N_8317,N_8225);
nor U8524 (N_8524,N_8289,N_8226);
and U8525 (N_8525,N_8350,N_8272);
or U8526 (N_8526,N_8375,N_8211);
nand U8527 (N_8527,N_8380,N_8207);
nand U8528 (N_8528,N_8300,N_8347);
nand U8529 (N_8529,N_8267,N_8214);
nand U8530 (N_8530,N_8235,N_8279);
nor U8531 (N_8531,N_8224,N_8351);
or U8532 (N_8532,N_8370,N_8309);
nand U8533 (N_8533,N_8304,N_8279);
and U8534 (N_8534,N_8361,N_8203);
nand U8535 (N_8535,N_8244,N_8340);
nand U8536 (N_8536,N_8251,N_8212);
nor U8537 (N_8537,N_8245,N_8350);
nand U8538 (N_8538,N_8312,N_8358);
and U8539 (N_8539,N_8399,N_8305);
xor U8540 (N_8540,N_8337,N_8284);
nand U8541 (N_8541,N_8342,N_8343);
or U8542 (N_8542,N_8369,N_8296);
xnor U8543 (N_8543,N_8377,N_8257);
nor U8544 (N_8544,N_8271,N_8264);
nor U8545 (N_8545,N_8341,N_8308);
nand U8546 (N_8546,N_8349,N_8336);
nand U8547 (N_8547,N_8266,N_8389);
and U8548 (N_8548,N_8305,N_8226);
or U8549 (N_8549,N_8216,N_8292);
xnor U8550 (N_8550,N_8263,N_8334);
nor U8551 (N_8551,N_8333,N_8244);
nor U8552 (N_8552,N_8396,N_8338);
and U8553 (N_8553,N_8200,N_8208);
nand U8554 (N_8554,N_8333,N_8239);
nand U8555 (N_8555,N_8348,N_8264);
nand U8556 (N_8556,N_8324,N_8228);
nand U8557 (N_8557,N_8214,N_8218);
xor U8558 (N_8558,N_8331,N_8308);
xnor U8559 (N_8559,N_8334,N_8390);
nand U8560 (N_8560,N_8382,N_8398);
nand U8561 (N_8561,N_8362,N_8308);
nand U8562 (N_8562,N_8394,N_8347);
or U8563 (N_8563,N_8282,N_8213);
nand U8564 (N_8564,N_8395,N_8265);
xnor U8565 (N_8565,N_8301,N_8353);
nor U8566 (N_8566,N_8244,N_8397);
xnor U8567 (N_8567,N_8269,N_8228);
nand U8568 (N_8568,N_8282,N_8326);
nand U8569 (N_8569,N_8319,N_8311);
nand U8570 (N_8570,N_8336,N_8251);
xnor U8571 (N_8571,N_8211,N_8241);
and U8572 (N_8572,N_8318,N_8391);
nand U8573 (N_8573,N_8263,N_8241);
nand U8574 (N_8574,N_8356,N_8271);
or U8575 (N_8575,N_8381,N_8274);
xor U8576 (N_8576,N_8348,N_8214);
nor U8577 (N_8577,N_8282,N_8397);
or U8578 (N_8578,N_8267,N_8303);
or U8579 (N_8579,N_8316,N_8206);
or U8580 (N_8580,N_8338,N_8287);
and U8581 (N_8581,N_8399,N_8308);
nand U8582 (N_8582,N_8252,N_8338);
and U8583 (N_8583,N_8374,N_8217);
or U8584 (N_8584,N_8251,N_8392);
nor U8585 (N_8585,N_8247,N_8282);
nand U8586 (N_8586,N_8368,N_8325);
nand U8587 (N_8587,N_8288,N_8326);
and U8588 (N_8588,N_8378,N_8207);
nor U8589 (N_8589,N_8385,N_8351);
and U8590 (N_8590,N_8307,N_8340);
nor U8591 (N_8591,N_8210,N_8216);
and U8592 (N_8592,N_8232,N_8237);
or U8593 (N_8593,N_8397,N_8327);
xnor U8594 (N_8594,N_8326,N_8342);
and U8595 (N_8595,N_8303,N_8250);
nand U8596 (N_8596,N_8211,N_8343);
xor U8597 (N_8597,N_8304,N_8365);
nand U8598 (N_8598,N_8318,N_8213);
nand U8599 (N_8599,N_8398,N_8310);
nand U8600 (N_8600,N_8595,N_8568);
nor U8601 (N_8601,N_8548,N_8419);
or U8602 (N_8602,N_8530,N_8430);
or U8603 (N_8603,N_8450,N_8539);
or U8604 (N_8604,N_8563,N_8451);
nand U8605 (N_8605,N_8432,N_8458);
nor U8606 (N_8606,N_8513,N_8526);
nor U8607 (N_8607,N_8538,N_8436);
nor U8608 (N_8608,N_8414,N_8581);
nor U8609 (N_8609,N_8543,N_8582);
nand U8610 (N_8610,N_8492,N_8479);
nor U8611 (N_8611,N_8402,N_8422);
and U8612 (N_8612,N_8462,N_8577);
xnor U8613 (N_8613,N_8592,N_8567);
and U8614 (N_8614,N_8481,N_8516);
and U8615 (N_8615,N_8437,N_8590);
nor U8616 (N_8616,N_8456,N_8566);
and U8617 (N_8617,N_8535,N_8413);
or U8618 (N_8618,N_8557,N_8598);
or U8619 (N_8619,N_8453,N_8517);
nand U8620 (N_8620,N_8427,N_8527);
or U8621 (N_8621,N_8501,N_8507);
or U8622 (N_8622,N_8429,N_8586);
xor U8623 (N_8623,N_8589,N_8541);
nand U8624 (N_8624,N_8572,N_8417);
or U8625 (N_8625,N_8404,N_8476);
xor U8626 (N_8626,N_8468,N_8489);
and U8627 (N_8627,N_8485,N_8502);
and U8628 (N_8628,N_8483,N_8559);
nor U8629 (N_8629,N_8534,N_8529);
or U8630 (N_8630,N_8552,N_8521);
nand U8631 (N_8631,N_8486,N_8519);
and U8632 (N_8632,N_8425,N_8440);
or U8633 (N_8633,N_8588,N_8421);
nand U8634 (N_8634,N_8447,N_8444);
nand U8635 (N_8635,N_8474,N_8593);
nor U8636 (N_8636,N_8464,N_8499);
xor U8637 (N_8637,N_8438,N_8509);
xor U8638 (N_8638,N_8573,N_8504);
nand U8639 (N_8639,N_8431,N_8463);
or U8640 (N_8640,N_8599,N_8518);
or U8641 (N_8641,N_8545,N_8547);
nand U8642 (N_8642,N_8415,N_8574);
xnor U8643 (N_8643,N_8571,N_8555);
and U8644 (N_8644,N_8569,N_8418);
or U8645 (N_8645,N_8410,N_8487);
nor U8646 (N_8646,N_8411,N_8452);
and U8647 (N_8647,N_8470,N_8523);
or U8648 (N_8648,N_8484,N_8578);
xor U8649 (N_8649,N_8554,N_8493);
or U8650 (N_8650,N_8442,N_8550);
nand U8651 (N_8651,N_8473,N_8565);
nand U8652 (N_8652,N_8400,N_8505);
nand U8653 (N_8653,N_8512,N_8457);
or U8654 (N_8654,N_8405,N_8584);
and U8655 (N_8655,N_8575,N_8401);
xor U8656 (N_8656,N_8537,N_8594);
and U8657 (N_8657,N_8403,N_8449);
xnor U8658 (N_8658,N_8477,N_8446);
or U8659 (N_8659,N_8585,N_8524);
nor U8660 (N_8660,N_8570,N_8556);
and U8661 (N_8661,N_8542,N_8471);
xor U8662 (N_8662,N_8511,N_8433);
nand U8663 (N_8663,N_8435,N_8472);
nor U8664 (N_8664,N_8407,N_8455);
nor U8665 (N_8665,N_8461,N_8416);
xnor U8666 (N_8666,N_8424,N_8439);
nand U8667 (N_8667,N_8597,N_8490);
nor U8668 (N_8668,N_8443,N_8448);
xor U8669 (N_8669,N_8494,N_8583);
or U8670 (N_8670,N_8531,N_8459);
xnor U8671 (N_8671,N_8469,N_8500);
nand U8672 (N_8672,N_8467,N_8525);
xnor U8673 (N_8673,N_8482,N_8576);
nand U8674 (N_8674,N_8426,N_8551);
nand U8675 (N_8675,N_8591,N_8408);
nor U8676 (N_8676,N_8522,N_8561);
nor U8677 (N_8677,N_8497,N_8549);
nor U8678 (N_8678,N_8478,N_8434);
or U8679 (N_8679,N_8558,N_8560);
nand U8680 (N_8680,N_8506,N_8587);
nand U8681 (N_8681,N_8515,N_8428);
nand U8682 (N_8682,N_8495,N_8553);
nand U8683 (N_8683,N_8533,N_8445);
nand U8684 (N_8684,N_8536,N_8514);
nor U8685 (N_8685,N_8475,N_8488);
nand U8686 (N_8686,N_8544,N_8496);
or U8687 (N_8687,N_8406,N_8579);
xor U8688 (N_8688,N_8532,N_8546);
and U8689 (N_8689,N_8454,N_8409);
or U8690 (N_8690,N_8460,N_8503);
nand U8691 (N_8691,N_8466,N_8564);
xor U8692 (N_8692,N_8510,N_8520);
nand U8693 (N_8693,N_8596,N_8423);
and U8694 (N_8694,N_8498,N_8540);
xnor U8695 (N_8695,N_8465,N_8420);
or U8696 (N_8696,N_8491,N_8528);
nand U8697 (N_8697,N_8508,N_8441);
or U8698 (N_8698,N_8412,N_8580);
or U8699 (N_8699,N_8480,N_8562);
nand U8700 (N_8700,N_8511,N_8451);
nor U8701 (N_8701,N_8492,N_8547);
nand U8702 (N_8702,N_8537,N_8447);
and U8703 (N_8703,N_8417,N_8592);
or U8704 (N_8704,N_8511,N_8480);
xor U8705 (N_8705,N_8466,N_8573);
and U8706 (N_8706,N_8503,N_8559);
nand U8707 (N_8707,N_8592,N_8518);
nand U8708 (N_8708,N_8520,N_8581);
nand U8709 (N_8709,N_8437,N_8404);
nor U8710 (N_8710,N_8539,N_8542);
nand U8711 (N_8711,N_8523,N_8511);
and U8712 (N_8712,N_8475,N_8473);
xor U8713 (N_8713,N_8408,N_8551);
nand U8714 (N_8714,N_8515,N_8452);
or U8715 (N_8715,N_8486,N_8502);
nand U8716 (N_8716,N_8463,N_8400);
nand U8717 (N_8717,N_8599,N_8545);
or U8718 (N_8718,N_8512,N_8502);
nor U8719 (N_8719,N_8414,N_8400);
nor U8720 (N_8720,N_8514,N_8459);
or U8721 (N_8721,N_8472,N_8449);
xor U8722 (N_8722,N_8506,N_8533);
xor U8723 (N_8723,N_8452,N_8513);
nand U8724 (N_8724,N_8479,N_8584);
nand U8725 (N_8725,N_8558,N_8420);
nor U8726 (N_8726,N_8450,N_8581);
and U8727 (N_8727,N_8418,N_8553);
and U8728 (N_8728,N_8526,N_8596);
and U8729 (N_8729,N_8527,N_8420);
and U8730 (N_8730,N_8552,N_8569);
or U8731 (N_8731,N_8527,N_8599);
nand U8732 (N_8732,N_8472,N_8415);
nor U8733 (N_8733,N_8490,N_8582);
nor U8734 (N_8734,N_8532,N_8562);
xor U8735 (N_8735,N_8509,N_8490);
nor U8736 (N_8736,N_8572,N_8489);
and U8737 (N_8737,N_8589,N_8432);
xor U8738 (N_8738,N_8556,N_8528);
nand U8739 (N_8739,N_8568,N_8486);
or U8740 (N_8740,N_8516,N_8526);
or U8741 (N_8741,N_8514,N_8584);
nor U8742 (N_8742,N_8459,N_8543);
and U8743 (N_8743,N_8518,N_8550);
or U8744 (N_8744,N_8409,N_8464);
nor U8745 (N_8745,N_8492,N_8549);
and U8746 (N_8746,N_8591,N_8422);
xor U8747 (N_8747,N_8588,N_8556);
or U8748 (N_8748,N_8557,N_8596);
xor U8749 (N_8749,N_8428,N_8434);
and U8750 (N_8750,N_8475,N_8460);
and U8751 (N_8751,N_8483,N_8445);
xor U8752 (N_8752,N_8507,N_8514);
nand U8753 (N_8753,N_8450,N_8438);
and U8754 (N_8754,N_8595,N_8522);
or U8755 (N_8755,N_8469,N_8580);
xor U8756 (N_8756,N_8582,N_8484);
or U8757 (N_8757,N_8542,N_8488);
xnor U8758 (N_8758,N_8575,N_8420);
nand U8759 (N_8759,N_8409,N_8439);
xor U8760 (N_8760,N_8413,N_8591);
xor U8761 (N_8761,N_8448,N_8498);
xor U8762 (N_8762,N_8429,N_8452);
and U8763 (N_8763,N_8560,N_8481);
xnor U8764 (N_8764,N_8447,N_8588);
nor U8765 (N_8765,N_8487,N_8419);
or U8766 (N_8766,N_8405,N_8501);
xnor U8767 (N_8767,N_8518,N_8519);
nor U8768 (N_8768,N_8468,N_8528);
and U8769 (N_8769,N_8472,N_8574);
nand U8770 (N_8770,N_8537,N_8496);
nor U8771 (N_8771,N_8503,N_8525);
or U8772 (N_8772,N_8531,N_8599);
nor U8773 (N_8773,N_8430,N_8489);
xor U8774 (N_8774,N_8582,N_8488);
xor U8775 (N_8775,N_8422,N_8421);
and U8776 (N_8776,N_8404,N_8533);
nor U8777 (N_8777,N_8475,N_8410);
or U8778 (N_8778,N_8578,N_8433);
nor U8779 (N_8779,N_8557,N_8489);
and U8780 (N_8780,N_8543,N_8554);
or U8781 (N_8781,N_8405,N_8436);
nor U8782 (N_8782,N_8599,N_8540);
and U8783 (N_8783,N_8553,N_8584);
nand U8784 (N_8784,N_8415,N_8411);
nand U8785 (N_8785,N_8496,N_8524);
nand U8786 (N_8786,N_8434,N_8505);
and U8787 (N_8787,N_8582,N_8585);
or U8788 (N_8788,N_8578,N_8517);
nor U8789 (N_8789,N_8541,N_8567);
and U8790 (N_8790,N_8488,N_8409);
nand U8791 (N_8791,N_8564,N_8489);
nor U8792 (N_8792,N_8520,N_8463);
or U8793 (N_8793,N_8420,N_8455);
xor U8794 (N_8794,N_8548,N_8569);
xnor U8795 (N_8795,N_8514,N_8474);
and U8796 (N_8796,N_8511,N_8522);
xnor U8797 (N_8797,N_8471,N_8531);
nand U8798 (N_8798,N_8490,N_8481);
nor U8799 (N_8799,N_8523,N_8447);
nor U8800 (N_8800,N_8697,N_8714);
nor U8801 (N_8801,N_8759,N_8626);
nor U8802 (N_8802,N_8689,N_8706);
or U8803 (N_8803,N_8730,N_8771);
or U8804 (N_8804,N_8653,N_8671);
and U8805 (N_8805,N_8734,N_8708);
and U8806 (N_8806,N_8655,N_8633);
xnor U8807 (N_8807,N_8642,N_8761);
or U8808 (N_8808,N_8647,N_8636);
or U8809 (N_8809,N_8776,N_8618);
nor U8810 (N_8810,N_8783,N_8792);
nor U8811 (N_8811,N_8693,N_8742);
nor U8812 (N_8812,N_8721,N_8681);
nand U8813 (N_8813,N_8602,N_8641);
and U8814 (N_8814,N_8621,N_8627);
nand U8815 (N_8815,N_8796,N_8749);
or U8816 (N_8816,N_8649,N_8700);
nand U8817 (N_8817,N_8748,N_8637);
or U8818 (N_8818,N_8798,N_8613);
and U8819 (N_8819,N_8600,N_8604);
nor U8820 (N_8820,N_8767,N_8654);
or U8821 (N_8821,N_8608,N_8793);
xnor U8822 (N_8822,N_8664,N_8659);
nand U8823 (N_8823,N_8666,N_8678);
nor U8824 (N_8824,N_8747,N_8797);
nand U8825 (N_8825,N_8732,N_8780);
or U8826 (N_8826,N_8754,N_8769);
or U8827 (N_8827,N_8687,N_8603);
nor U8828 (N_8828,N_8625,N_8745);
and U8829 (N_8829,N_8778,N_8795);
xnor U8830 (N_8830,N_8652,N_8645);
and U8831 (N_8831,N_8648,N_8752);
and U8832 (N_8832,N_8683,N_8741);
nor U8833 (N_8833,N_8668,N_8644);
xnor U8834 (N_8834,N_8782,N_8725);
or U8835 (N_8835,N_8722,N_8619);
nand U8836 (N_8836,N_8672,N_8764);
nor U8837 (N_8837,N_8794,N_8766);
and U8838 (N_8838,N_8727,N_8660);
or U8839 (N_8839,N_8770,N_8674);
and U8840 (N_8840,N_8682,N_8643);
nand U8841 (N_8841,N_8785,N_8777);
and U8842 (N_8842,N_8779,N_8605);
xnor U8843 (N_8843,N_8699,N_8616);
nand U8844 (N_8844,N_8787,N_8650);
nor U8845 (N_8845,N_8784,N_8629);
nor U8846 (N_8846,N_8713,N_8612);
nor U8847 (N_8847,N_8673,N_8753);
nand U8848 (N_8848,N_8694,N_8737);
nand U8849 (N_8849,N_8726,N_8635);
and U8850 (N_8850,N_8601,N_8698);
xnor U8851 (N_8851,N_8617,N_8679);
or U8852 (N_8852,N_8788,N_8661);
xnor U8853 (N_8853,N_8718,N_8738);
and U8854 (N_8854,N_8606,N_8663);
and U8855 (N_8855,N_8733,N_8758);
nor U8856 (N_8856,N_8670,N_8773);
nor U8857 (N_8857,N_8765,N_8715);
nor U8858 (N_8858,N_8712,N_8786);
or U8859 (N_8859,N_8760,N_8640);
xor U8860 (N_8860,N_8638,N_8763);
xor U8861 (N_8861,N_8790,N_8609);
xor U8862 (N_8862,N_8744,N_8724);
or U8863 (N_8863,N_8688,N_8658);
xor U8864 (N_8864,N_8675,N_8729);
and U8865 (N_8865,N_8702,N_8762);
or U8866 (N_8866,N_8680,N_8791);
and U8867 (N_8867,N_8781,N_8768);
xor U8868 (N_8868,N_8720,N_8711);
nand U8869 (N_8869,N_8611,N_8685);
and U8870 (N_8870,N_8705,N_8707);
xor U8871 (N_8871,N_8716,N_8622);
nor U8872 (N_8872,N_8614,N_8701);
and U8873 (N_8873,N_8620,N_8686);
and U8874 (N_8874,N_8667,N_8676);
and U8875 (N_8875,N_8775,N_8631);
nor U8876 (N_8876,N_8799,N_8703);
nand U8877 (N_8877,N_8607,N_8624);
and U8878 (N_8878,N_8639,N_8630);
nor U8879 (N_8879,N_8665,N_8657);
nand U8880 (N_8880,N_8634,N_8756);
and U8881 (N_8881,N_8740,N_8750);
nor U8882 (N_8882,N_8628,N_8755);
nand U8883 (N_8883,N_8695,N_8704);
xor U8884 (N_8884,N_8610,N_8774);
nand U8885 (N_8885,N_8736,N_8692);
nand U8886 (N_8886,N_8757,N_8651);
nand U8887 (N_8887,N_8728,N_8710);
xnor U8888 (N_8888,N_8615,N_8656);
or U8889 (N_8889,N_8731,N_8662);
and U8890 (N_8890,N_8669,N_8646);
and U8891 (N_8891,N_8789,N_8719);
nor U8892 (N_8892,N_8677,N_8623);
nor U8893 (N_8893,N_8632,N_8746);
nor U8894 (N_8894,N_8691,N_8709);
nor U8895 (N_8895,N_8751,N_8743);
or U8896 (N_8896,N_8739,N_8684);
nor U8897 (N_8897,N_8696,N_8690);
or U8898 (N_8898,N_8723,N_8717);
xnor U8899 (N_8899,N_8735,N_8772);
nand U8900 (N_8900,N_8734,N_8682);
xnor U8901 (N_8901,N_8631,N_8627);
xnor U8902 (N_8902,N_8658,N_8619);
nand U8903 (N_8903,N_8682,N_8787);
xor U8904 (N_8904,N_8757,N_8769);
or U8905 (N_8905,N_8636,N_8721);
and U8906 (N_8906,N_8748,N_8675);
and U8907 (N_8907,N_8649,N_8633);
nand U8908 (N_8908,N_8789,N_8620);
xor U8909 (N_8909,N_8630,N_8772);
or U8910 (N_8910,N_8697,N_8706);
xor U8911 (N_8911,N_8663,N_8646);
nor U8912 (N_8912,N_8615,N_8737);
xnor U8913 (N_8913,N_8620,N_8795);
nor U8914 (N_8914,N_8665,N_8776);
and U8915 (N_8915,N_8756,N_8717);
nor U8916 (N_8916,N_8746,N_8694);
xnor U8917 (N_8917,N_8666,N_8611);
and U8918 (N_8918,N_8655,N_8739);
nor U8919 (N_8919,N_8731,N_8656);
xnor U8920 (N_8920,N_8739,N_8746);
xor U8921 (N_8921,N_8760,N_8653);
and U8922 (N_8922,N_8739,N_8740);
nor U8923 (N_8923,N_8792,N_8692);
and U8924 (N_8924,N_8600,N_8675);
nor U8925 (N_8925,N_8777,N_8746);
nand U8926 (N_8926,N_8611,N_8799);
or U8927 (N_8927,N_8621,N_8605);
nor U8928 (N_8928,N_8683,N_8771);
and U8929 (N_8929,N_8687,N_8753);
nand U8930 (N_8930,N_8645,N_8619);
xor U8931 (N_8931,N_8645,N_8690);
xor U8932 (N_8932,N_8782,N_8664);
nor U8933 (N_8933,N_8617,N_8626);
and U8934 (N_8934,N_8650,N_8729);
xor U8935 (N_8935,N_8709,N_8719);
nor U8936 (N_8936,N_8729,N_8703);
xor U8937 (N_8937,N_8617,N_8619);
nor U8938 (N_8938,N_8774,N_8639);
nand U8939 (N_8939,N_8618,N_8682);
or U8940 (N_8940,N_8645,N_8720);
or U8941 (N_8941,N_8755,N_8688);
and U8942 (N_8942,N_8648,N_8613);
and U8943 (N_8943,N_8686,N_8749);
or U8944 (N_8944,N_8781,N_8732);
xnor U8945 (N_8945,N_8747,N_8631);
and U8946 (N_8946,N_8697,N_8783);
xor U8947 (N_8947,N_8669,N_8715);
or U8948 (N_8948,N_8756,N_8722);
nand U8949 (N_8949,N_8752,N_8661);
and U8950 (N_8950,N_8624,N_8664);
xnor U8951 (N_8951,N_8730,N_8601);
nand U8952 (N_8952,N_8664,N_8715);
xor U8953 (N_8953,N_8684,N_8704);
nand U8954 (N_8954,N_8700,N_8708);
nor U8955 (N_8955,N_8644,N_8685);
or U8956 (N_8956,N_8765,N_8730);
or U8957 (N_8957,N_8747,N_8717);
and U8958 (N_8958,N_8779,N_8645);
or U8959 (N_8959,N_8612,N_8651);
nor U8960 (N_8960,N_8648,N_8626);
or U8961 (N_8961,N_8725,N_8608);
xnor U8962 (N_8962,N_8613,N_8607);
nor U8963 (N_8963,N_8671,N_8649);
and U8964 (N_8964,N_8632,N_8608);
or U8965 (N_8965,N_8656,N_8643);
nor U8966 (N_8966,N_8610,N_8793);
and U8967 (N_8967,N_8638,N_8688);
xor U8968 (N_8968,N_8766,N_8747);
nand U8969 (N_8969,N_8681,N_8620);
and U8970 (N_8970,N_8751,N_8614);
nand U8971 (N_8971,N_8722,N_8784);
xor U8972 (N_8972,N_8771,N_8666);
nor U8973 (N_8973,N_8609,N_8606);
xnor U8974 (N_8974,N_8758,N_8602);
nor U8975 (N_8975,N_8762,N_8631);
and U8976 (N_8976,N_8669,N_8733);
or U8977 (N_8977,N_8782,N_8766);
or U8978 (N_8978,N_8675,N_8750);
or U8979 (N_8979,N_8692,N_8719);
or U8980 (N_8980,N_8702,N_8691);
nand U8981 (N_8981,N_8772,N_8682);
and U8982 (N_8982,N_8733,N_8773);
and U8983 (N_8983,N_8798,N_8695);
xnor U8984 (N_8984,N_8618,N_8677);
xor U8985 (N_8985,N_8641,N_8723);
xnor U8986 (N_8986,N_8723,N_8636);
nand U8987 (N_8987,N_8764,N_8696);
and U8988 (N_8988,N_8794,N_8710);
nor U8989 (N_8989,N_8671,N_8687);
nand U8990 (N_8990,N_8724,N_8601);
and U8991 (N_8991,N_8636,N_8712);
nand U8992 (N_8992,N_8657,N_8770);
nor U8993 (N_8993,N_8680,N_8671);
xor U8994 (N_8994,N_8792,N_8789);
xnor U8995 (N_8995,N_8758,N_8694);
xor U8996 (N_8996,N_8618,N_8741);
and U8997 (N_8997,N_8799,N_8644);
and U8998 (N_8998,N_8673,N_8762);
nor U8999 (N_8999,N_8738,N_8715);
or U9000 (N_9000,N_8923,N_8895);
xnor U9001 (N_9001,N_8842,N_8935);
nand U9002 (N_9002,N_8902,N_8900);
or U9003 (N_9003,N_8963,N_8953);
and U9004 (N_9004,N_8985,N_8858);
or U9005 (N_9005,N_8885,N_8814);
and U9006 (N_9006,N_8947,N_8987);
nor U9007 (N_9007,N_8825,N_8944);
and U9008 (N_9008,N_8862,N_8971);
nor U9009 (N_9009,N_8955,N_8848);
nand U9010 (N_9010,N_8886,N_8838);
and U9011 (N_9011,N_8928,N_8986);
and U9012 (N_9012,N_8847,N_8998);
nor U9013 (N_9013,N_8929,N_8918);
nand U9014 (N_9014,N_8989,N_8994);
nor U9015 (N_9015,N_8818,N_8832);
xnor U9016 (N_9016,N_8835,N_8908);
nand U9017 (N_9017,N_8959,N_8840);
and U9018 (N_9018,N_8804,N_8965);
and U9019 (N_9019,N_8888,N_8952);
or U9020 (N_9020,N_8917,N_8864);
nand U9021 (N_9021,N_8871,N_8878);
nor U9022 (N_9022,N_8823,N_8803);
xnor U9023 (N_9023,N_8837,N_8933);
nand U9024 (N_9024,N_8974,N_8833);
or U9025 (N_9025,N_8925,N_8802);
nor U9026 (N_9026,N_8907,N_8932);
nand U9027 (N_9027,N_8868,N_8873);
nand U9028 (N_9028,N_8915,N_8817);
nand U9029 (N_9029,N_8827,N_8831);
or U9030 (N_9030,N_8820,N_8949);
nor U9031 (N_9031,N_8958,N_8887);
and U9032 (N_9032,N_8863,N_8811);
or U9033 (N_9033,N_8897,N_8903);
or U9034 (N_9034,N_8984,N_8910);
nand U9035 (N_9035,N_8957,N_8881);
and U9036 (N_9036,N_8853,N_8800);
xnor U9037 (N_9037,N_8939,N_8828);
nor U9038 (N_9038,N_8934,N_8836);
xor U9039 (N_9039,N_8826,N_8941);
nand U9040 (N_9040,N_8927,N_8812);
nor U9041 (N_9041,N_8936,N_8877);
xnor U9042 (N_9042,N_8816,N_8909);
nor U9043 (N_9043,N_8970,N_8824);
or U9044 (N_9044,N_8942,N_8951);
nand U9045 (N_9045,N_8839,N_8968);
or U9046 (N_9046,N_8901,N_8852);
and U9047 (N_9047,N_8866,N_8843);
and U9048 (N_9048,N_8892,N_8992);
xnor U9049 (N_9049,N_8899,N_8830);
xor U9050 (N_9050,N_8937,N_8930);
nand U9051 (N_9051,N_8972,N_8884);
xnor U9052 (N_9052,N_8977,N_8962);
or U9053 (N_9053,N_8996,N_8813);
and U9054 (N_9054,N_8912,N_8846);
and U9055 (N_9055,N_8880,N_8919);
or U9056 (N_9056,N_8995,N_8938);
nand U9057 (N_9057,N_8926,N_8964);
and U9058 (N_9058,N_8834,N_8980);
and U9059 (N_9059,N_8879,N_8898);
and U9060 (N_9060,N_8896,N_8991);
nand U9061 (N_9061,N_8809,N_8854);
nand U9062 (N_9062,N_8969,N_8867);
nor U9063 (N_9063,N_8876,N_8806);
nor U9064 (N_9064,N_8882,N_8967);
and U9065 (N_9065,N_8870,N_8821);
xor U9066 (N_9066,N_8875,N_8889);
xor U9067 (N_9067,N_8861,N_8801);
nand U9068 (N_9068,N_8819,N_8851);
or U9069 (N_9069,N_8855,N_8931);
and U9070 (N_9070,N_8924,N_8921);
nand U9071 (N_9071,N_8990,N_8805);
nor U9072 (N_9072,N_8913,N_8943);
nor U9073 (N_9073,N_8906,N_8905);
nor U9074 (N_9074,N_8954,N_8960);
xnor U9075 (N_9075,N_8883,N_8856);
or U9076 (N_9076,N_8844,N_8916);
nand U9077 (N_9077,N_8982,N_8865);
and U9078 (N_9078,N_8845,N_8914);
nor U9079 (N_9079,N_8822,N_8860);
or U9080 (N_9080,N_8872,N_8891);
and U9081 (N_9081,N_8966,N_8922);
xnor U9082 (N_9082,N_8940,N_8979);
nand U9083 (N_9083,N_8874,N_8945);
nor U9084 (N_9084,N_8850,N_8807);
nand U9085 (N_9085,N_8904,N_8841);
and U9086 (N_9086,N_8894,N_8869);
xnor U9087 (N_9087,N_8810,N_8956);
or U9088 (N_9088,N_8849,N_8859);
xor U9089 (N_9089,N_8893,N_8961);
xnor U9090 (N_9090,N_8920,N_8993);
xor U9091 (N_9091,N_8978,N_8911);
or U9092 (N_9092,N_8857,N_8815);
nor U9093 (N_9093,N_8808,N_8950);
or U9094 (N_9094,N_8999,N_8890);
nand U9095 (N_9095,N_8988,N_8983);
or U9096 (N_9096,N_8829,N_8981);
and U9097 (N_9097,N_8948,N_8975);
and U9098 (N_9098,N_8976,N_8946);
nor U9099 (N_9099,N_8997,N_8973);
nand U9100 (N_9100,N_8830,N_8926);
nor U9101 (N_9101,N_8879,N_8956);
or U9102 (N_9102,N_8873,N_8882);
xnor U9103 (N_9103,N_8981,N_8817);
nand U9104 (N_9104,N_8850,N_8919);
nor U9105 (N_9105,N_8829,N_8943);
nand U9106 (N_9106,N_8867,N_8887);
or U9107 (N_9107,N_8928,N_8904);
and U9108 (N_9108,N_8933,N_8841);
or U9109 (N_9109,N_8841,N_8949);
or U9110 (N_9110,N_8907,N_8837);
and U9111 (N_9111,N_8913,N_8885);
xor U9112 (N_9112,N_8836,N_8809);
or U9113 (N_9113,N_8930,N_8890);
or U9114 (N_9114,N_8893,N_8937);
nor U9115 (N_9115,N_8845,N_8939);
or U9116 (N_9116,N_8946,N_8859);
nand U9117 (N_9117,N_8912,N_8998);
nor U9118 (N_9118,N_8946,N_8894);
nor U9119 (N_9119,N_8939,N_8974);
nand U9120 (N_9120,N_8851,N_8986);
and U9121 (N_9121,N_8889,N_8814);
or U9122 (N_9122,N_8955,N_8907);
nand U9123 (N_9123,N_8977,N_8890);
xnor U9124 (N_9124,N_8907,N_8893);
xor U9125 (N_9125,N_8976,N_8977);
nor U9126 (N_9126,N_8870,N_8860);
nand U9127 (N_9127,N_8984,N_8806);
or U9128 (N_9128,N_8900,N_8891);
and U9129 (N_9129,N_8981,N_8877);
or U9130 (N_9130,N_8932,N_8995);
nor U9131 (N_9131,N_8818,N_8983);
or U9132 (N_9132,N_8975,N_8879);
or U9133 (N_9133,N_8879,N_8955);
and U9134 (N_9134,N_8981,N_8896);
or U9135 (N_9135,N_8885,N_8904);
xor U9136 (N_9136,N_8924,N_8944);
nor U9137 (N_9137,N_8898,N_8984);
and U9138 (N_9138,N_8996,N_8923);
nor U9139 (N_9139,N_8941,N_8969);
and U9140 (N_9140,N_8808,N_8846);
nand U9141 (N_9141,N_8808,N_8969);
nand U9142 (N_9142,N_8833,N_8839);
xor U9143 (N_9143,N_8801,N_8804);
nand U9144 (N_9144,N_8809,N_8943);
xnor U9145 (N_9145,N_8858,N_8882);
xor U9146 (N_9146,N_8989,N_8934);
nor U9147 (N_9147,N_8980,N_8923);
xnor U9148 (N_9148,N_8932,N_8841);
nor U9149 (N_9149,N_8950,N_8979);
nand U9150 (N_9150,N_8884,N_8805);
xor U9151 (N_9151,N_8828,N_8876);
nor U9152 (N_9152,N_8996,N_8938);
nor U9153 (N_9153,N_8975,N_8929);
or U9154 (N_9154,N_8926,N_8810);
or U9155 (N_9155,N_8933,N_8863);
nor U9156 (N_9156,N_8849,N_8906);
xor U9157 (N_9157,N_8983,N_8845);
nand U9158 (N_9158,N_8868,N_8883);
nand U9159 (N_9159,N_8885,N_8983);
nor U9160 (N_9160,N_8875,N_8974);
nand U9161 (N_9161,N_8893,N_8934);
nor U9162 (N_9162,N_8925,N_8824);
nand U9163 (N_9163,N_8815,N_8984);
nor U9164 (N_9164,N_8930,N_8970);
or U9165 (N_9165,N_8806,N_8923);
xnor U9166 (N_9166,N_8987,N_8830);
xnor U9167 (N_9167,N_8814,N_8983);
and U9168 (N_9168,N_8969,N_8985);
or U9169 (N_9169,N_8923,N_8833);
nor U9170 (N_9170,N_8956,N_8811);
and U9171 (N_9171,N_8982,N_8950);
nand U9172 (N_9172,N_8815,N_8905);
nand U9173 (N_9173,N_8935,N_8837);
xor U9174 (N_9174,N_8827,N_8986);
and U9175 (N_9175,N_8856,N_8891);
xnor U9176 (N_9176,N_8885,N_8851);
nor U9177 (N_9177,N_8887,N_8871);
and U9178 (N_9178,N_8941,N_8824);
or U9179 (N_9179,N_8881,N_8982);
xnor U9180 (N_9180,N_8917,N_8814);
or U9181 (N_9181,N_8853,N_8820);
nand U9182 (N_9182,N_8908,N_8937);
or U9183 (N_9183,N_8893,N_8849);
nor U9184 (N_9184,N_8970,N_8943);
or U9185 (N_9185,N_8912,N_8887);
or U9186 (N_9186,N_8886,N_8978);
nand U9187 (N_9187,N_8956,N_8817);
nor U9188 (N_9188,N_8848,N_8898);
nand U9189 (N_9189,N_8948,N_8969);
nand U9190 (N_9190,N_8993,N_8952);
nor U9191 (N_9191,N_8855,N_8995);
nand U9192 (N_9192,N_8969,N_8874);
or U9193 (N_9193,N_8914,N_8894);
xor U9194 (N_9194,N_8950,N_8895);
or U9195 (N_9195,N_8946,N_8804);
nand U9196 (N_9196,N_8947,N_8812);
or U9197 (N_9197,N_8981,N_8949);
or U9198 (N_9198,N_8842,N_8899);
and U9199 (N_9199,N_8899,N_8948);
nor U9200 (N_9200,N_9147,N_9118);
or U9201 (N_9201,N_9101,N_9045);
nor U9202 (N_9202,N_9098,N_9005);
nand U9203 (N_9203,N_9164,N_9003);
or U9204 (N_9204,N_9057,N_9157);
xor U9205 (N_9205,N_9084,N_9117);
nor U9206 (N_9206,N_9167,N_9053);
or U9207 (N_9207,N_9100,N_9188);
and U9208 (N_9208,N_9006,N_9081);
and U9209 (N_9209,N_9044,N_9055);
or U9210 (N_9210,N_9011,N_9136);
xor U9211 (N_9211,N_9022,N_9114);
and U9212 (N_9212,N_9054,N_9048);
xnor U9213 (N_9213,N_9033,N_9073);
or U9214 (N_9214,N_9079,N_9018);
nand U9215 (N_9215,N_9028,N_9189);
nand U9216 (N_9216,N_9001,N_9181);
xnor U9217 (N_9217,N_9056,N_9177);
or U9218 (N_9218,N_9088,N_9155);
xor U9219 (N_9219,N_9130,N_9038);
nor U9220 (N_9220,N_9183,N_9091);
nand U9221 (N_9221,N_9036,N_9134);
xnor U9222 (N_9222,N_9162,N_9035);
nor U9223 (N_9223,N_9043,N_9042);
nand U9224 (N_9224,N_9106,N_9166);
or U9225 (N_9225,N_9170,N_9026);
nor U9226 (N_9226,N_9129,N_9111);
and U9227 (N_9227,N_9014,N_9058);
nor U9228 (N_9228,N_9143,N_9175);
nand U9229 (N_9229,N_9063,N_9027);
nor U9230 (N_9230,N_9163,N_9105);
and U9231 (N_9231,N_9000,N_9116);
xor U9232 (N_9232,N_9065,N_9094);
or U9233 (N_9233,N_9191,N_9152);
xnor U9234 (N_9234,N_9107,N_9103);
nor U9235 (N_9235,N_9127,N_9110);
nand U9236 (N_9236,N_9034,N_9082);
and U9237 (N_9237,N_9086,N_9156);
xnor U9238 (N_9238,N_9004,N_9146);
xnor U9239 (N_9239,N_9122,N_9153);
xnor U9240 (N_9240,N_9049,N_9019);
xnor U9241 (N_9241,N_9184,N_9171);
nor U9242 (N_9242,N_9062,N_9090);
nor U9243 (N_9243,N_9140,N_9132);
or U9244 (N_9244,N_9097,N_9104);
nor U9245 (N_9245,N_9083,N_9197);
nor U9246 (N_9246,N_9023,N_9198);
nand U9247 (N_9247,N_9076,N_9180);
and U9248 (N_9248,N_9072,N_9135);
and U9249 (N_9249,N_9121,N_9150);
nand U9250 (N_9250,N_9138,N_9069);
xor U9251 (N_9251,N_9031,N_9050);
nand U9252 (N_9252,N_9078,N_9002);
or U9253 (N_9253,N_9040,N_9039);
nand U9254 (N_9254,N_9025,N_9179);
nand U9255 (N_9255,N_9182,N_9099);
or U9256 (N_9256,N_9151,N_9187);
or U9257 (N_9257,N_9161,N_9010);
xor U9258 (N_9258,N_9037,N_9144);
or U9259 (N_9259,N_9199,N_9194);
or U9260 (N_9260,N_9158,N_9108);
nand U9261 (N_9261,N_9046,N_9115);
xor U9262 (N_9262,N_9133,N_9172);
or U9263 (N_9263,N_9169,N_9120);
nand U9264 (N_9264,N_9074,N_9052);
and U9265 (N_9265,N_9007,N_9148);
xnor U9266 (N_9266,N_9080,N_9092);
nor U9267 (N_9267,N_9087,N_9142);
xnor U9268 (N_9268,N_9176,N_9095);
xor U9269 (N_9269,N_9126,N_9112);
nand U9270 (N_9270,N_9016,N_9013);
nor U9271 (N_9271,N_9173,N_9195);
nor U9272 (N_9272,N_9124,N_9119);
and U9273 (N_9273,N_9051,N_9185);
and U9274 (N_9274,N_9030,N_9141);
xor U9275 (N_9275,N_9070,N_9160);
xor U9276 (N_9276,N_9123,N_9113);
nor U9277 (N_9277,N_9024,N_9017);
nor U9278 (N_9278,N_9061,N_9096);
nor U9279 (N_9279,N_9165,N_9125);
xor U9280 (N_9280,N_9077,N_9159);
nand U9281 (N_9281,N_9139,N_9029);
and U9282 (N_9282,N_9066,N_9102);
nand U9283 (N_9283,N_9093,N_9145);
or U9284 (N_9284,N_9196,N_9012);
xor U9285 (N_9285,N_9041,N_9168);
and U9286 (N_9286,N_9109,N_9060);
nand U9287 (N_9287,N_9075,N_9193);
xnor U9288 (N_9288,N_9071,N_9021);
xnor U9289 (N_9289,N_9089,N_9015);
nand U9290 (N_9290,N_9067,N_9178);
nor U9291 (N_9291,N_9032,N_9008);
nor U9292 (N_9292,N_9059,N_9131);
or U9293 (N_9293,N_9064,N_9020);
and U9294 (N_9294,N_9137,N_9149);
or U9295 (N_9295,N_9186,N_9068);
or U9296 (N_9296,N_9154,N_9009);
and U9297 (N_9297,N_9128,N_9192);
and U9298 (N_9298,N_9190,N_9047);
or U9299 (N_9299,N_9174,N_9085);
nand U9300 (N_9300,N_9184,N_9186);
nand U9301 (N_9301,N_9086,N_9061);
xor U9302 (N_9302,N_9017,N_9000);
nand U9303 (N_9303,N_9143,N_9044);
nor U9304 (N_9304,N_9134,N_9100);
or U9305 (N_9305,N_9026,N_9188);
nand U9306 (N_9306,N_9072,N_9087);
xor U9307 (N_9307,N_9106,N_9141);
and U9308 (N_9308,N_9130,N_9058);
nor U9309 (N_9309,N_9129,N_9136);
xnor U9310 (N_9310,N_9077,N_9130);
nor U9311 (N_9311,N_9065,N_9158);
nand U9312 (N_9312,N_9039,N_9126);
or U9313 (N_9313,N_9144,N_9148);
or U9314 (N_9314,N_9048,N_9179);
nand U9315 (N_9315,N_9134,N_9142);
nand U9316 (N_9316,N_9043,N_9105);
and U9317 (N_9317,N_9015,N_9194);
nor U9318 (N_9318,N_9174,N_9177);
xnor U9319 (N_9319,N_9096,N_9015);
xor U9320 (N_9320,N_9137,N_9040);
xnor U9321 (N_9321,N_9141,N_9028);
xor U9322 (N_9322,N_9059,N_9160);
nor U9323 (N_9323,N_9109,N_9081);
nor U9324 (N_9324,N_9195,N_9034);
nand U9325 (N_9325,N_9000,N_9018);
and U9326 (N_9326,N_9152,N_9017);
nand U9327 (N_9327,N_9054,N_9192);
nor U9328 (N_9328,N_9090,N_9155);
or U9329 (N_9329,N_9142,N_9032);
nor U9330 (N_9330,N_9148,N_9015);
or U9331 (N_9331,N_9143,N_9107);
nand U9332 (N_9332,N_9006,N_9107);
nand U9333 (N_9333,N_9030,N_9032);
and U9334 (N_9334,N_9168,N_9142);
or U9335 (N_9335,N_9067,N_9086);
nand U9336 (N_9336,N_9013,N_9009);
nor U9337 (N_9337,N_9192,N_9115);
nor U9338 (N_9338,N_9061,N_9177);
and U9339 (N_9339,N_9165,N_9099);
and U9340 (N_9340,N_9006,N_9188);
xor U9341 (N_9341,N_9199,N_9156);
nor U9342 (N_9342,N_9160,N_9004);
nand U9343 (N_9343,N_9135,N_9077);
and U9344 (N_9344,N_9183,N_9146);
nor U9345 (N_9345,N_9150,N_9030);
xnor U9346 (N_9346,N_9068,N_9141);
nor U9347 (N_9347,N_9102,N_9046);
xnor U9348 (N_9348,N_9130,N_9013);
xnor U9349 (N_9349,N_9057,N_9024);
or U9350 (N_9350,N_9176,N_9112);
nand U9351 (N_9351,N_9063,N_9002);
nor U9352 (N_9352,N_9035,N_9078);
nand U9353 (N_9353,N_9006,N_9073);
and U9354 (N_9354,N_9042,N_9031);
xor U9355 (N_9355,N_9122,N_9009);
nor U9356 (N_9356,N_9165,N_9114);
xnor U9357 (N_9357,N_9111,N_9117);
nand U9358 (N_9358,N_9081,N_9070);
and U9359 (N_9359,N_9134,N_9172);
and U9360 (N_9360,N_9044,N_9172);
or U9361 (N_9361,N_9085,N_9189);
nor U9362 (N_9362,N_9169,N_9041);
or U9363 (N_9363,N_9136,N_9089);
nor U9364 (N_9364,N_9171,N_9127);
nor U9365 (N_9365,N_9053,N_9060);
xnor U9366 (N_9366,N_9190,N_9144);
or U9367 (N_9367,N_9160,N_9086);
and U9368 (N_9368,N_9069,N_9025);
nand U9369 (N_9369,N_9173,N_9153);
nand U9370 (N_9370,N_9108,N_9010);
or U9371 (N_9371,N_9064,N_9002);
or U9372 (N_9372,N_9120,N_9078);
xnor U9373 (N_9373,N_9169,N_9123);
xor U9374 (N_9374,N_9034,N_9146);
and U9375 (N_9375,N_9132,N_9151);
or U9376 (N_9376,N_9021,N_9063);
or U9377 (N_9377,N_9110,N_9019);
and U9378 (N_9378,N_9142,N_9198);
xnor U9379 (N_9379,N_9199,N_9162);
xor U9380 (N_9380,N_9147,N_9072);
xnor U9381 (N_9381,N_9174,N_9031);
nor U9382 (N_9382,N_9086,N_9105);
nand U9383 (N_9383,N_9116,N_9081);
and U9384 (N_9384,N_9112,N_9148);
nor U9385 (N_9385,N_9151,N_9143);
or U9386 (N_9386,N_9162,N_9148);
and U9387 (N_9387,N_9157,N_9172);
and U9388 (N_9388,N_9176,N_9052);
nor U9389 (N_9389,N_9033,N_9013);
nand U9390 (N_9390,N_9100,N_9042);
or U9391 (N_9391,N_9031,N_9182);
or U9392 (N_9392,N_9008,N_9114);
nand U9393 (N_9393,N_9095,N_9154);
or U9394 (N_9394,N_9160,N_9192);
nor U9395 (N_9395,N_9061,N_9126);
and U9396 (N_9396,N_9171,N_9117);
and U9397 (N_9397,N_9140,N_9150);
xnor U9398 (N_9398,N_9168,N_9178);
xnor U9399 (N_9399,N_9080,N_9005);
or U9400 (N_9400,N_9346,N_9265);
xnor U9401 (N_9401,N_9247,N_9275);
or U9402 (N_9402,N_9330,N_9369);
nand U9403 (N_9403,N_9260,N_9373);
xnor U9404 (N_9404,N_9240,N_9288);
or U9405 (N_9405,N_9376,N_9339);
nand U9406 (N_9406,N_9372,N_9331);
nand U9407 (N_9407,N_9203,N_9221);
nor U9408 (N_9408,N_9209,N_9284);
xor U9409 (N_9409,N_9223,N_9202);
or U9410 (N_9410,N_9338,N_9348);
nand U9411 (N_9411,N_9263,N_9388);
and U9412 (N_9412,N_9345,N_9311);
nand U9413 (N_9413,N_9321,N_9305);
xnor U9414 (N_9414,N_9279,N_9313);
xor U9415 (N_9415,N_9341,N_9237);
or U9416 (N_9416,N_9258,N_9241);
and U9417 (N_9417,N_9361,N_9296);
nor U9418 (N_9418,N_9262,N_9363);
or U9419 (N_9419,N_9201,N_9266);
nor U9420 (N_9420,N_9366,N_9350);
or U9421 (N_9421,N_9278,N_9355);
nor U9422 (N_9422,N_9302,N_9328);
nand U9423 (N_9423,N_9390,N_9292);
and U9424 (N_9424,N_9300,N_9234);
and U9425 (N_9425,N_9259,N_9364);
or U9426 (N_9426,N_9378,N_9236);
nor U9427 (N_9427,N_9282,N_9204);
or U9428 (N_9428,N_9213,N_9243);
xor U9429 (N_9429,N_9285,N_9324);
nand U9430 (N_9430,N_9271,N_9316);
and U9431 (N_9431,N_9309,N_9360);
or U9432 (N_9432,N_9224,N_9342);
xor U9433 (N_9433,N_9347,N_9280);
xor U9434 (N_9434,N_9248,N_9233);
or U9435 (N_9435,N_9289,N_9381);
nor U9436 (N_9436,N_9244,N_9225);
nor U9437 (N_9437,N_9398,N_9270);
and U9438 (N_9438,N_9367,N_9255);
nand U9439 (N_9439,N_9303,N_9337);
nand U9440 (N_9440,N_9229,N_9357);
and U9441 (N_9441,N_9205,N_9326);
xor U9442 (N_9442,N_9294,N_9394);
or U9443 (N_9443,N_9343,N_9396);
nand U9444 (N_9444,N_9232,N_9252);
xnor U9445 (N_9445,N_9293,N_9272);
xor U9446 (N_9446,N_9214,N_9317);
nand U9447 (N_9447,N_9217,N_9297);
xnor U9448 (N_9448,N_9315,N_9267);
nor U9449 (N_9449,N_9371,N_9249);
and U9450 (N_9450,N_9256,N_9384);
nand U9451 (N_9451,N_9274,N_9399);
nor U9452 (N_9452,N_9298,N_9264);
xor U9453 (N_9453,N_9310,N_9322);
xor U9454 (N_9454,N_9242,N_9349);
nor U9455 (N_9455,N_9352,N_9395);
or U9456 (N_9456,N_9304,N_9218);
or U9457 (N_9457,N_9253,N_9333);
or U9458 (N_9458,N_9210,N_9319);
or U9459 (N_9459,N_9336,N_9392);
xor U9460 (N_9460,N_9382,N_9239);
xnor U9461 (N_9461,N_9375,N_9314);
nand U9462 (N_9462,N_9312,N_9358);
xnor U9463 (N_9463,N_9273,N_9261);
or U9464 (N_9464,N_9226,N_9318);
and U9465 (N_9465,N_9320,N_9301);
nor U9466 (N_9466,N_9238,N_9389);
nor U9467 (N_9467,N_9215,N_9329);
nor U9468 (N_9468,N_9377,N_9332);
xor U9469 (N_9469,N_9380,N_9283);
or U9470 (N_9470,N_9359,N_9212);
and U9471 (N_9471,N_9277,N_9379);
xor U9472 (N_9472,N_9220,N_9368);
nand U9473 (N_9473,N_9351,N_9386);
and U9474 (N_9474,N_9340,N_9397);
nand U9475 (N_9475,N_9335,N_9208);
or U9476 (N_9476,N_9344,N_9286);
or U9477 (N_9477,N_9334,N_9268);
or U9478 (N_9478,N_9353,N_9354);
or U9479 (N_9479,N_9287,N_9323);
xor U9480 (N_9480,N_9254,N_9306);
or U9481 (N_9481,N_9276,N_9269);
nor U9482 (N_9482,N_9230,N_9281);
xnor U9483 (N_9483,N_9290,N_9391);
nand U9484 (N_9484,N_9299,N_9370);
xnor U9485 (N_9485,N_9257,N_9291);
and U9486 (N_9486,N_9251,N_9206);
nand U9487 (N_9487,N_9308,N_9362);
nand U9488 (N_9488,N_9365,N_9200);
and U9489 (N_9489,N_9211,N_9325);
or U9490 (N_9490,N_9246,N_9219);
nand U9491 (N_9491,N_9207,N_9216);
or U9492 (N_9492,N_9228,N_9356);
and U9493 (N_9493,N_9387,N_9383);
xnor U9494 (N_9494,N_9245,N_9250);
nand U9495 (N_9495,N_9295,N_9327);
nor U9496 (N_9496,N_9374,N_9235);
nand U9497 (N_9497,N_9227,N_9231);
and U9498 (N_9498,N_9393,N_9307);
nor U9499 (N_9499,N_9385,N_9222);
nor U9500 (N_9500,N_9296,N_9297);
or U9501 (N_9501,N_9291,N_9383);
or U9502 (N_9502,N_9318,N_9355);
xnor U9503 (N_9503,N_9267,N_9230);
nand U9504 (N_9504,N_9365,N_9243);
or U9505 (N_9505,N_9274,N_9322);
or U9506 (N_9506,N_9243,N_9237);
nor U9507 (N_9507,N_9372,N_9222);
nand U9508 (N_9508,N_9279,N_9241);
or U9509 (N_9509,N_9391,N_9250);
nand U9510 (N_9510,N_9250,N_9370);
nand U9511 (N_9511,N_9216,N_9394);
nor U9512 (N_9512,N_9303,N_9240);
xor U9513 (N_9513,N_9290,N_9361);
and U9514 (N_9514,N_9231,N_9336);
and U9515 (N_9515,N_9293,N_9241);
and U9516 (N_9516,N_9345,N_9396);
or U9517 (N_9517,N_9347,N_9228);
nand U9518 (N_9518,N_9234,N_9355);
and U9519 (N_9519,N_9322,N_9243);
or U9520 (N_9520,N_9378,N_9314);
nor U9521 (N_9521,N_9207,N_9282);
nand U9522 (N_9522,N_9315,N_9387);
nor U9523 (N_9523,N_9282,N_9382);
and U9524 (N_9524,N_9200,N_9281);
xnor U9525 (N_9525,N_9228,N_9327);
xor U9526 (N_9526,N_9317,N_9249);
and U9527 (N_9527,N_9270,N_9342);
and U9528 (N_9528,N_9282,N_9317);
xnor U9529 (N_9529,N_9280,N_9211);
and U9530 (N_9530,N_9200,N_9322);
nand U9531 (N_9531,N_9361,N_9284);
nand U9532 (N_9532,N_9294,N_9304);
and U9533 (N_9533,N_9272,N_9247);
and U9534 (N_9534,N_9200,N_9391);
nor U9535 (N_9535,N_9381,N_9246);
and U9536 (N_9536,N_9366,N_9226);
or U9537 (N_9537,N_9302,N_9296);
and U9538 (N_9538,N_9283,N_9303);
xnor U9539 (N_9539,N_9240,N_9376);
or U9540 (N_9540,N_9201,N_9221);
xnor U9541 (N_9541,N_9292,N_9256);
xnor U9542 (N_9542,N_9226,N_9372);
nand U9543 (N_9543,N_9324,N_9244);
and U9544 (N_9544,N_9230,N_9237);
and U9545 (N_9545,N_9215,N_9216);
nor U9546 (N_9546,N_9367,N_9257);
and U9547 (N_9547,N_9296,N_9352);
and U9548 (N_9548,N_9272,N_9211);
xnor U9549 (N_9549,N_9367,N_9290);
nand U9550 (N_9550,N_9270,N_9332);
nor U9551 (N_9551,N_9330,N_9382);
xnor U9552 (N_9552,N_9233,N_9224);
nand U9553 (N_9553,N_9308,N_9216);
nor U9554 (N_9554,N_9320,N_9305);
nand U9555 (N_9555,N_9384,N_9241);
xor U9556 (N_9556,N_9261,N_9333);
and U9557 (N_9557,N_9351,N_9233);
nand U9558 (N_9558,N_9297,N_9346);
xor U9559 (N_9559,N_9374,N_9344);
xor U9560 (N_9560,N_9215,N_9287);
nor U9561 (N_9561,N_9358,N_9213);
nand U9562 (N_9562,N_9344,N_9281);
xor U9563 (N_9563,N_9312,N_9304);
xor U9564 (N_9564,N_9205,N_9257);
and U9565 (N_9565,N_9308,N_9363);
nor U9566 (N_9566,N_9260,N_9202);
or U9567 (N_9567,N_9208,N_9273);
nor U9568 (N_9568,N_9369,N_9301);
xor U9569 (N_9569,N_9288,N_9390);
and U9570 (N_9570,N_9278,N_9299);
and U9571 (N_9571,N_9378,N_9367);
nand U9572 (N_9572,N_9330,N_9392);
nor U9573 (N_9573,N_9253,N_9216);
or U9574 (N_9574,N_9235,N_9216);
xnor U9575 (N_9575,N_9211,N_9344);
or U9576 (N_9576,N_9393,N_9264);
or U9577 (N_9577,N_9338,N_9243);
nand U9578 (N_9578,N_9272,N_9373);
and U9579 (N_9579,N_9377,N_9208);
nor U9580 (N_9580,N_9309,N_9333);
xor U9581 (N_9581,N_9292,N_9388);
nor U9582 (N_9582,N_9264,N_9259);
xnor U9583 (N_9583,N_9369,N_9345);
nand U9584 (N_9584,N_9361,N_9242);
or U9585 (N_9585,N_9398,N_9344);
nand U9586 (N_9586,N_9399,N_9365);
and U9587 (N_9587,N_9373,N_9381);
and U9588 (N_9588,N_9366,N_9269);
or U9589 (N_9589,N_9283,N_9370);
nand U9590 (N_9590,N_9329,N_9300);
nor U9591 (N_9591,N_9376,N_9344);
xnor U9592 (N_9592,N_9318,N_9373);
and U9593 (N_9593,N_9365,N_9381);
and U9594 (N_9594,N_9397,N_9241);
or U9595 (N_9595,N_9376,N_9224);
nand U9596 (N_9596,N_9263,N_9367);
or U9597 (N_9597,N_9394,N_9276);
xnor U9598 (N_9598,N_9348,N_9263);
nand U9599 (N_9599,N_9355,N_9367);
xnor U9600 (N_9600,N_9541,N_9423);
or U9601 (N_9601,N_9491,N_9436);
nor U9602 (N_9602,N_9478,N_9463);
xnor U9603 (N_9603,N_9557,N_9555);
or U9604 (N_9604,N_9475,N_9570);
nor U9605 (N_9605,N_9418,N_9453);
xor U9606 (N_9606,N_9554,N_9432);
nor U9607 (N_9607,N_9558,N_9486);
xor U9608 (N_9608,N_9568,N_9477);
nand U9609 (N_9609,N_9429,N_9580);
and U9610 (N_9610,N_9550,N_9565);
nor U9611 (N_9611,N_9579,N_9575);
xor U9612 (N_9612,N_9513,N_9566);
and U9613 (N_9613,N_9467,N_9439);
xnor U9614 (N_9614,N_9598,N_9562);
xor U9615 (N_9615,N_9595,N_9523);
or U9616 (N_9616,N_9407,N_9404);
and U9617 (N_9617,N_9574,N_9531);
or U9618 (N_9618,N_9470,N_9548);
and U9619 (N_9619,N_9573,N_9560);
or U9620 (N_9620,N_9485,N_9444);
or U9621 (N_9621,N_9545,N_9414);
nand U9622 (N_9622,N_9515,N_9505);
or U9623 (N_9623,N_9532,N_9497);
and U9624 (N_9624,N_9488,N_9447);
xor U9625 (N_9625,N_9421,N_9521);
nor U9626 (N_9626,N_9489,N_9484);
xor U9627 (N_9627,N_9587,N_9535);
nor U9628 (N_9628,N_9435,N_9469);
or U9629 (N_9629,N_9425,N_9437);
nand U9630 (N_9630,N_9519,N_9449);
and U9631 (N_9631,N_9563,N_9594);
nor U9632 (N_9632,N_9460,N_9508);
and U9633 (N_9633,N_9529,N_9415);
nand U9634 (N_9634,N_9542,N_9520);
nor U9635 (N_9635,N_9517,N_9401);
nand U9636 (N_9636,N_9472,N_9493);
nor U9637 (N_9637,N_9585,N_9504);
xnor U9638 (N_9638,N_9501,N_9589);
and U9639 (N_9639,N_9537,N_9487);
nand U9640 (N_9640,N_9583,N_9496);
and U9641 (N_9641,N_9443,N_9567);
nand U9642 (N_9642,N_9446,N_9546);
nor U9643 (N_9643,N_9581,N_9556);
and U9644 (N_9644,N_9534,N_9528);
or U9645 (N_9645,N_9416,N_9473);
and U9646 (N_9646,N_9438,N_9572);
and U9647 (N_9647,N_9576,N_9405);
or U9648 (N_9648,N_9547,N_9474);
xor U9649 (N_9649,N_9413,N_9549);
or U9650 (N_9650,N_9507,N_9403);
nand U9651 (N_9651,N_9494,N_9522);
xor U9652 (N_9652,N_9536,N_9559);
xor U9653 (N_9653,N_9586,N_9509);
nor U9654 (N_9654,N_9540,N_9527);
or U9655 (N_9655,N_9482,N_9569);
nand U9656 (N_9656,N_9420,N_9483);
xor U9657 (N_9657,N_9433,N_9476);
nor U9658 (N_9658,N_9406,N_9578);
xnor U9659 (N_9659,N_9490,N_9454);
or U9660 (N_9660,N_9465,N_9468);
xnor U9661 (N_9661,N_9526,N_9597);
or U9662 (N_9662,N_9599,N_9458);
nand U9663 (N_9663,N_9440,N_9577);
or U9664 (N_9664,N_9448,N_9512);
nand U9665 (N_9665,N_9495,N_9492);
xor U9666 (N_9666,N_9464,N_9408);
nand U9667 (N_9667,N_9503,N_9410);
and U9668 (N_9668,N_9400,N_9419);
nand U9669 (N_9669,N_9596,N_9498);
and U9670 (N_9670,N_9462,N_9452);
nand U9671 (N_9671,N_9481,N_9430);
and U9672 (N_9672,N_9480,N_9431);
nor U9673 (N_9673,N_9561,N_9466);
or U9674 (N_9674,N_9530,N_9525);
nand U9675 (N_9675,N_9409,N_9538);
nand U9676 (N_9676,N_9424,N_9551);
xor U9677 (N_9677,N_9434,N_9412);
or U9678 (N_9678,N_9422,N_9506);
nor U9679 (N_9679,N_9499,N_9402);
nand U9680 (N_9680,N_9428,N_9450);
nand U9681 (N_9681,N_9455,N_9461);
xor U9682 (N_9682,N_9427,N_9442);
and U9683 (N_9683,N_9411,N_9510);
or U9684 (N_9684,N_9518,N_9553);
or U9685 (N_9685,N_9524,N_9592);
and U9686 (N_9686,N_9544,N_9533);
nor U9687 (N_9687,N_9582,N_9502);
nand U9688 (N_9688,N_9459,N_9426);
nand U9689 (N_9689,N_9471,N_9516);
xor U9690 (N_9690,N_9500,N_9417);
nand U9691 (N_9691,N_9552,N_9584);
or U9692 (N_9692,N_9590,N_9445);
nand U9693 (N_9693,N_9514,N_9593);
or U9694 (N_9694,N_9564,N_9451);
and U9695 (N_9695,N_9479,N_9588);
nand U9696 (N_9696,N_9539,N_9457);
xnor U9697 (N_9697,N_9571,N_9456);
nand U9698 (N_9698,N_9441,N_9511);
and U9699 (N_9699,N_9591,N_9543);
or U9700 (N_9700,N_9495,N_9597);
xnor U9701 (N_9701,N_9536,N_9475);
nand U9702 (N_9702,N_9470,N_9593);
or U9703 (N_9703,N_9476,N_9557);
or U9704 (N_9704,N_9599,N_9591);
xnor U9705 (N_9705,N_9516,N_9442);
xnor U9706 (N_9706,N_9456,N_9581);
or U9707 (N_9707,N_9407,N_9440);
nor U9708 (N_9708,N_9579,N_9448);
xnor U9709 (N_9709,N_9450,N_9472);
xor U9710 (N_9710,N_9573,N_9435);
and U9711 (N_9711,N_9536,N_9425);
and U9712 (N_9712,N_9496,N_9501);
xnor U9713 (N_9713,N_9538,N_9492);
or U9714 (N_9714,N_9419,N_9422);
nor U9715 (N_9715,N_9568,N_9427);
nor U9716 (N_9716,N_9452,N_9581);
xnor U9717 (N_9717,N_9502,N_9495);
nor U9718 (N_9718,N_9502,N_9404);
and U9719 (N_9719,N_9426,N_9407);
nand U9720 (N_9720,N_9579,N_9576);
nor U9721 (N_9721,N_9565,N_9512);
or U9722 (N_9722,N_9410,N_9485);
or U9723 (N_9723,N_9505,N_9417);
nand U9724 (N_9724,N_9567,N_9440);
xnor U9725 (N_9725,N_9496,N_9447);
and U9726 (N_9726,N_9459,N_9507);
xor U9727 (N_9727,N_9468,N_9474);
and U9728 (N_9728,N_9584,N_9402);
xnor U9729 (N_9729,N_9440,N_9582);
or U9730 (N_9730,N_9406,N_9455);
nand U9731 (N_9731,N_9458,N_9428);
nand U9732 (N_9732,N_9552,N_9430);
and U9733 (N_9733,N_9431,N_9580);
nand U9734 (N_9734,N_9547,N_9500);
nand U9735 (N_9735,N_9461,N_9491);
and U9736 (N_9736,N_9421,N_9432);
nor U9737 (N_9737,N_9591,N_9447);
or U9738 (N_9738,N_9413,N_9485);
nand U9739 (N_9739,N_9593,N_9534);
nor U9740 (N_9740,N_9443,N_9539);
or U9741 (N_9741,N_9563,N_9573);
xor U9742 (N_9742,N_9501,N_9541);
or U9743 (N_9743,N_9502,N_9432);
nor U9744 (N_9744,N_9423,N_9584);
and U9745 (N_9745,N_9480,N_9435);
nor U9746 (N_9746,N_9459,N_9521);
xnor U9747 (N_9747,N_9451,N_9593);
and U9748 (N_9748,N_9452,N_9573);
or U9749 (N_9749,N_9556,N_9465);
and U9750 (N_9750,N_9412,N_9452);
nand U9751 (N_9751,N_9558,N_9408);
nand U9752 (N_9752,N_9447,N_9592);
nor U9753 (N_9753,N_9591,N_9518);
or U9754 (N_9754,N_9507,N_9543);
and U9755 (N_9755,N_9532,N_9402);
nor U9756 (N_9756,N_9503,N_9477);
xnor U9757 (N_9757,N_9431,N_9513);
or U9758 (N_9758,N_9537,N_9574);
xor U9759 (N_9759,N_9557,N_9505);
and U9760 (N_9760,N_9581,N_9477);
and U9761 (N_9761,N_9580,N_9518);
and U9762 (N_9762,N_9430,N_9487);
nand U9763 (N_9763,N_9535,N_9550);
and U9764 (N_9764,N_9504,N_9587);
or U9765 (N_9765,N_9574,N_9495);
nand U9766 (N_9766,N_9502,N_9523);
nand U9767 (N_9767,N_9514,N_9478);
nand U9768 (N_9768,N_9450,N_9452);
nor U9769 (N_9769,N_9512,N_9549);
nor U9770 (N_9770,N_9404,N_9558);
nand U9771 (N_9771,N_9585,N_9445);
nor U9772 (N_9772,N_9574,N_9526);
nand U9773 (N_9773,N_9506,N_9468);
and U9774 (N_9774,N_9453,N_9591);
xor U9775 (N_9775,N_9411,N_9483);
or U9776 (N_9776,N_9565,N_9509);
nor U9777 (N_9777,N_9430,N_9453);
nor U9778 (N_9778,N_9560,N_9473);
and U9779 (N_9779,N_9405,N_9527);
xnor U9780 (N_9780,N_9529,N_9596);
xor U9781 (N_9781,N_9535,N_9554);
nand U9782 (N_9782,N_9420,N_9523);
and U9783 (N_9783,N_9512,N_9455);
nand U9784 (N_9784,N_9511,N_9599);
nor U9785 (N_9785,N_9472,N_9571);
nand U9786 (N_9786,N_9447,N_9578);
xor U9787 (N_9787,N_9473,N_9567);
nor U9788 (N_9788,N_9581,N_9406);
and U9789 (N_9789,N_9581,N_9589);
nand U9790 (N_9790,N_9489,N_9495);
xnor U9791 (N_9791,N_9583,N_9412);
nor U9792 (N_9792,N_9550,N_9525);
or U9793 (N_9793,N_9516,N_9548);
nor U9794 (N_9794,N_9448,N_9569);
xnor U9795 (N_9795,N_9449,N_9541);
xnor U9796 (N_9796,N_9463,N_9453);
and U9797 (N_9797,N_9488,N_9495);
xor U9798 (N_9798,N_9452,N_9488);
or U9799 (N_9799,N_9435,N_9562);
nor U9800 (N_9800,N_9791,N_9764);
nor U9801 (N_9801,N_9797,N_9731);
and U9802 (N_9802,N_9648,N_9641);
nor U9803 (N_9803,N_9605,N_9734);
or U9804 (N_9804,N_9735,N_9742);
or U9805 (N_9805,N_9726,N_9795);
xnor U9806 (N_9806,N_9668,N_9620);
xnor U9807 (N_9807,N_9732,N_9689);
or U9808 (N_9808,N_9697,N_9761);
or U9809 (N_9809,N_9792,N_9747);
and U9810 (N_9810,N_9753,N_9757);
nor U9811 (N_9811,N_9671,N_9690);
nor U9812 (N_9812,N_9681,N_9642);
or U9813 (N_9813,N_9781,N_9750);
nor U9814 (N_9814,N_9717,N_9619);
nor U9815 (N_9815,N_9686,N_9646);
nand U9816 (N_9816,N_9656,N_9624);
and U9817 (N_9817,N_9688,N_9607);
nand U9818 (N_9818,N_9775,N_9730);
or U9819 (N_9819,N_9739,N_9674);
nand U9820 (N_9820,N_9774,N_9770);
nand U9821 (N_9821,N_9756,N_9768);
and U9822 (N_9822,N_9632,N_9719);
and U9823 (N_9823,N_9702,N_9673);
xor U9824 (N_9824,N_9704,N_9758);
xnor U9825 (N_9825,N_9694,N_9603);
and U9826 (N_9826,N_9787,N_9779);
nor U9827 (N_9827,N_9691,N_9773);
and U9828 (N_9828,N_9728,N_9696);
nand U9829 (N_9829,N_9666,N_9749);
or U9830 (N_9830,N_9615,N_9617);
xor U9831 (N_9831,N_9755,N_9789);
and U9832 (N_9832,N_9608,N_9633);
or U9833 (N_9833,N_9647,N_9752);
or U9834 (N_9834,N_9796,N_9723);
and U9835 (N_9835,N_9629,N_9780);
xor U9836 (N_9836,N_9606,N_9659);
nor U9837 (N_9837,N_9713,N_9751);
nor U9838 (N_9838,N_9613,N_9655);
nand U9839 (N_9839,N_9746,N_9675);
nand U9840 (N_9840,N_9604,N_9700);
xnor U9841 (N_9841,N_9651,N_9790);
xnor U9842 (N_9842,N_9721,N_9762);
and U9843 (N_9843,N_9712,N_9602);
or U9844 (N_9844,N_9616,N_9733);
xor U9845 (N_9845,N_9765,N_9623);
nor U9846 (N_9846,N_9766,N_9782);
nand U9847 (N_9847,N_9711,N_9705);
or U9848 (N_9848,N_9706,N_9715);
xor U9849 (N_9849,N_9683,N_9708);
xor U9850 (N_9850,N_9612,N_9718);
xor U9851 (N_9851,N_9664,N_9658);
and U9852 (N_9852,N_9710,N_9628);
nor U9853 (N_9853,N_9667,N_9625);
or U9854 (N_9854,N_9654,N_9622);
or U9855 (N_9855,N_9741,N_9669);
or U9856 (N_9856,N_9737,N_9794);
or U9857 (N_9857,N_9660,N_9631);
xnor U9858 (N_9858,N_9693,N_9639);
nand U9859 (N_9859,N_9670,N_9745);
xor U9860 (N_9860,N_9600,N_9784);
nand U9861 (N_9861,N_9677,N_9614);
nand U9862 (N_9862,N_9634,N_9759);
and U9863 (N_9863,N_9799,N_9783);
nor U9864 (N_9864,N_9662,N_9687);
and U9865 (N_9865,N_9692,N_9618);
or U9866 (N_9866,N_9786,N_9767);
nand U9867 (N_9867,N_9740,N_9645);
xnor U9868 (N_9868,N_9772,N_9672);
nand U9869 (N_9869,N_9725,N_9743);
and U9870 (N_9870,N_9744,N_9709);
or U9871 (N_9871,N_9778,N_9650);
and U9872 (N_9872,N_9601,N_9678);
and U9873 (N_9873,N_9714,N_9630);
and U9874 (N_9874,N_9682,N_9727);
nor U9875 (N_9875,N_9754,N_9638);
nand U9876 (N_9876,N_9769,N_9729);
or U9877 (N_9877,N_9676,N_9738);
xnor U9878 (N_9878,N_9643,N_9626);
nor U9879 (N_9879,N_9707,N_9665);
and U9880 (N_9880,N_9637,N_9777);
nand U9881 (N_9881,N_9621,N_9640);
or U9882 (N_9882,N_9657,N_9722);
nor U9883 (N_9883,N_9771,N_9798);
and U9884 (N_9884,N_9699,N_9701);
nand U9885 (N_9885,N_9627,N_9685);
and U9886 (N_9886,N_9649,N_9793);
and U9887 (N_9887,N_9661,N_9748);
nand U9888 (N_9888,N_9788,N_9776);
nand U9889 (N_9889,N_9684,N_9644);
nor U9890 (N_9890,N_9636,N_9736);
nor U9891 (N_9891,N_9680,N_9652);
nor U9892 (N_9892,N_9724,N_9720);
nor U9893 (N_9893,N_9611,N_9663);
or U9894 (N_9894,N_9695,N_9653);
xnor U9895 (N_9895,N_9760,N_9785);
or U9896 (N_9896,N_9763,N_9679);
nor U9897 (N_9897,N_9610,N_9703);
and U9898 (N_9898,N_9698,N_9635);
and U9899 (N_9899,N_9609,N_9716);
nor U9900 (N_9900,N_9637,N_9790);
nor U9901 (N_9901,N_9669,N_9695);
xnor U9902 (N_9902,N_9639,N_9654);
and U9903 (N_9903,N_9683,N_9795);
xnor U9904 (N_9904,N_9693,N_9617);
nor U9905 (N_9905,N_9727,N_9683);
or U9906 (N_9906,N_9686,N_9713);
or U9907 (N_9907,N_9605,N_9613);
nor U9908 (N_9908,N_9645,N_9642);
or U9909 (N_9909,N_9675,N_9767);
or U9910 (N_9910,N_9658,N_9722);
nand U9911 (N_9911,N_9761,N_9719);
or U9912 (N_9912,N_9699,N_9673);
nand U9913 (N_9913,N_9611,N_9617);
nor U9914 (N_9914,N_9796,N_9795);
nor U9915 (N_9915,N_9628,N_9773);
and U9916 (N_9916,N_9663,N_9604);
nor U9917 (N_9917,N_9647,N_9729);
xor U9918 (N_9918,N_9737,N_9627);
xnor U9919 (N_9919,N_9755,N_9647);
or U9920 (N_9920,N_9753,N_9619);
and U9921 (N_9921,N_9703,N_9768);
and U9922 (N_9922,N_9631,N_9610);
and U9923 (N_9923,N_9612,N_9660);
or U9924 (N_9924,N_9754,N_9685);
nand U9925 (N_9925,N_9712,N_9653);
xor U9926 (N_9926,N_9612,N_9636);
xnor U9927 (N_9927,N_9775,N_9734);
nand U9928 (N_9928,N_9758,N_9712);
xor U9929 (N_9929,N_9652,N_9670);
nand U9930 (N_9930,N_9683,N_9601);
or U9931 (N_9931,N_9792,N_9727);
xnor U9932 (N_9932,N_9788,N_9767);
nor U9933 (N_9933,N_9681,N_9641);
xor U9934 (N_9934,N_9604,N_9708);
nor U9935 (N_9935,N_9681,N_9784);
or U9936 (N_9936,N_9775,N_9749);
nand U9937 (N_9937,N_9612,N_9613);
or U9938 (N_9938,N_9692,N_9608);
and U9939 (N_9939,N_9702,N_9792);
nor U9940 (N_9940,N_9768,N_9689);
or U9941 (N_9941,N_9774,N_9763);
and U9942 (N_9942,N_9765,N_9785);
and U9943 (N_9943,N_9738,N_9769);
nand U9944 (N_9944,N_9609,N_9606);
nor U9945 (N_9945,N_9710,N_9745);
and U9946 (N_9946,N_9631,N_9654);
nand U9947 (N_9947,N_9755,N_9698);
xnor U9948 (N_9948,N_9762,N_9608);
nand U9949 (N_9949,N_9732,N_9773);
xnor U9950 (N_9950,N_9603,N_9739);
or U9951 (N_9951,N_9649,N_9736);
nor U9952 (N_9952,N_9712,N_9609);
nand U9953 (N_9953,N_9691,N_9697);
xor U9954 (N_9954,N_9639,N_9730);
xor U9955 (N_9955,N_9679,N_9611);
xor U9956 (N_9956,N_9686,N_9761);
xnor U9957 (N_9957,N_9744,N_9710);
nor U9958 (N_9958,N_9635,N_9626);
nand U9959 (N_9959,N_9606,N_9690);
nand U9960 (N_9960,N_9702,N_9727);
or U9961 (N_9961,N_9713,N_9645);
or U9962 (N_9962,N_9696,N_9708);
nor U9963 (N_9963,N_9764,N_9699);
nand U9964 (N_9964,N_9724,N_9754);
and U9965 (N_9965,N_9785,N_9708);
nand U9966 (N_9966,N_9741,N_9697);
or U9967 (N_9967,N_9785,N_9791);
nor U9968 (N_9968,N_9623,N_9769);
nor U9969 (N_9969,N_9657,N_9691);
xnor U9970 (N_9970,N_9776,N_9750);
nor U9971 (N_9971,N_9715,N_9752);
and U9972 (N_9972,N_9648,N_9710);
xor U9973 (N_9973,N_9754,N_9788);
and U9974 (N_9974,N_9631,N_9745);
xnor U9975 (N_9975,N_9758,N_9759);
nor U9976 (N_9976,N_9637,N_9766);
nor U9977 (N_9977,N_9767,N_9676);
or U9978 (N_9978,N_9737,N_9731);
and U9979 (N_9979,N_9737,N_9666);
nand U9980 (N_9980,N_9636,N_9719);
or U9981 (N_9981,N_9629,N_9662);
or U9982 (N_9982,N_9709,N_9604);
and U9983 (N_9983,N_9757,N_9642);
nor U9984 (N_9984,N_9749,N_9716);
or U9985 (N_9985,N_9716,N_9701);
and U9986 (N_9986,N_9639,N_9688);
nand U9987 (N_9987,N_9766,N_9651);
and U9988 (N_9988,N_9690,N_9712);
nand U9989 (N_9989,N_9656,N_9740);
nand U9990 (N_9990,N_9720,N_9607);
or U9991 (N_9991,N_9695,N_9612);
nor U9992 (N_9992,N_9752,N_9604);
xnor U9993 (N_9993,N_9623,N_9686);
xnor U9994 (N_9994,N_9629,N_9745);
nand U9995 (N_9995,N_9782,N_9795);
and U9996 (N_9996,N_9770,N_9666);
nor U9997 (N_9997,N_9672,N_9798);
nand U9998 (N_9998,N_9660,N_9697);
and U9999 (N_9999,N_9749,N_9771);
and UO_0 (O_0,N_9901,N_9964);
nand UO_1 (O_1,N_9881,N_9891);
and UO_2 (O_2,N_9999,N_9963);
and UO_3 (O_3,N_9951,N_9924);
and UO_4 (O_4,N_9867,N_9852);
and UO_5 (O_5,N_9941,N_9853);
and UO_6 (O_6,N_9961,N_9956);
nor UO_7 (O_7,N_9871,N_9811);
or UO_8 (O_8,N_9994,N_9893);
nand UO_9 (O_9,N_9940,N_9854);
or UO_10 (O_10,N_9882,N_9886);
or UO_11 (O_11,N_9874,N_9906);
and UO_12 (O_12,N_9947,N_9974);
nor UO_13 (O_13,N_9997,N_9932);
xor UO_14 (O_14,N_9814,N_9816);
nand UO_15 (O_15,N_9821,N_9897);
xor UO_16 (O_16,N_9800,N_9838);
nand UO_17 (O_17,N_9885,N_9898);
nor UO_18 (O_18,N_9972,N_9860);
nor UO_19 (O_19,N_9894,N_9960);
nand UO_20 (O_20,N_9808,N_9984);
nand UO_21 (O_21,N_9950,N_9824);
and UO_22 (O_22,N_9848,N_9958);
and UO_23 (O_23,N_9929,N_9919);
and UO_24 (O_24,N_9959,N_9869);
xnor UO_25 (O_25,N_9986,N_9985);
nand UO_26 (O_26,N_9827,N_9813);
or UO_27 (O_27,N_9903,N_9968);
or UO_28 (O_28,N_9908,N_9802);
nor UO_29 (O_29,N_9832,N_9948);
nand UO_30 (O_30,N_9916,N_9954);
and UO_31 (O_31,N_9868,N_9938);
and UO_32 (O_32,N_9945,N_9846);
nor UO_33 (O_33,N_9815,N_9939);
or UO_34 (O_34,N_9884,N_9933);
nor UO_35 (O_35,N_9879,N_9805);
nand UO_36 (O_36,N_9942,N_9944);
nor UO_37 (O_37,N_9988,N_9996);
and UO_38 (O_38,N_9807,N_9831);
xor UO_39 (O_39,N_9973,N_9880);
and UO_40 (O_40,N_9820,N_9979);
or UO_41 (O_41,N_9842,N_9856);
nor UO_42 (O_42,N_9981,N_9989);
xnor UO_43 (O_43,N_9978,N_9900);
nand UO_44 (O_44,N_9928,N_9822);
or UO_45 (O_45,N_9966,N_9876);
nor UO_46 (O_46,N_9943,N_9965);
nor UO_47 (O_47,N_9930,N_9847);
and UO_48 (O_48,N_9825,N_9819);
or UO_49 (O_49,N_9836,N_9833);
and UO_50 (O_50,N_9845,N_9803);
and UO_51 (O_51,N_9912,N_9926);
or UO_52 (O_52,N_9922,N_9976);
and UO_53 (O_53,N_9877,N_9980);
or UO_54 (O_54,N_9883,N_9895);
xnor UO_55 (O_55,N_9840,N_9872);
nand UO_56 (O_56,N_9826,N_9862);
and UO_57 (O_57,N_9873,N_9914);
nor UO_58 (O_58,N_9917,N_9993);
and UO_59 (O_59,N_9849,N_9946);
nand UO_60 (O_60,N_9804,N_9896);
xnor UO_61 (O_61,N_9935,N_9987);
or UO_62 (O_62,N_9920,N_9957);
xor UO_63 (O_63,N_9844,N_9817);
nor UO_64 (O_64,N_9982,N_9823);
and UO_65 (O_65,N_9955,N_9887);
nand UO_66 (O_66,N_9855,N_9969);
xor UO_67 (O_67,N_9962,N_9991);
nor UO_68 (O_68,N_9904,N_9801);
nor UO_69 (O_69,N_9859,N_9971);
nand UO_70 (O_70,N_9875,N_9810);
nor UO_71 (O_71,N_9857,N_9902);
nor UO_72 (O_72,N_9931,N_9861);
nor UO_73 (O_73,N_9936,N_9841);
nor UO_74 (O_74,N_9890,N_9878);
nor UO_75 (O_75,N_9866,N_9835);
nand UO_76 (O_76,N_9915,N_9850);
xnor UO_77 (O_77,N_9925,N_9907);
xor UO_78 (O_78,N_9809,N_9843);
nand UO_79 (O_79,N_9911,N_9863);
xor UO_80 (O_80,N_9864,N_9828);
and UO_81 (O_81,N_9953,N_9905);
nand UO_82 (O_82,N_9921,N_9913);
or UO_83 (O_83,N_9909,N_9806);
nor UO_84 (O_84,N_9858,N_9927);
nand UO_85 (O_85,N_9834,N_9983);
and UO_86 (O_86,N_9998,N_9934);
and UO_87 (O_87,N_9918,N_9990);
and UO_88 (O_88,N_9865,N_9952);
or UO_89 (O_89,N_9812,N_9830);
xor UO_90 (O_90,N_9837,N_9829);
nand UO_91 (O_91,N_9967,N_9851);
nor UO_92 (O_92,N_9995,N_9937);
xnor UO_93 (O_93,N_9839,N_9818);
nor UO_94 (O_94,N_9977,N_9910);
or UO_95 (O_95,N_9949,N_9899);
nor UO_96 (O_96,N_9888,N_9975);
nor UO_97 (O_97,N_9889,N_9870);
and UO_98 (O_98,N_9992,N_9970);
and UO_99 (O_99,N_9923,N_9892);
nand UO_100 (O_100,N_9978,N_9995);
or UO_101 (O_101,N_9865,N_9823);
xnor UO_102 (O_102,N_9807,N_9808);
or UO_103 (O_103,N_9964,N_9878);
xor UO_104 (O_104,N_9833,N_9911);
and UO_105 (O_105,N_9918,N_9881);
nand UO_106 (O_106,N_9875,N_9905);
nor UO_107 (O_107,N_9988,N_9875);
xnor UO_108 (O_108,N_9892,N_9904);
or UO_109 (O_109,N_9944,N_9858);
and UO_110 (O_110,N_9999,N_9987);
nand UO_111 (O_111,N_9830,N_9963);
nand UO_112 (O_112,N_9987,N_9885);
xnor UO_113 (O_113,N_9909,N_9982);
and UO_114 (O_114,N_9837,N_9900);
and UO_115 (O_115,N_9921,N_9931);
xor UO_116 (O_116,N_9901,N_9874);
nand UO_117 (O_117,N_9950,N_9821);
nand UO_118 (O_118,N_9869,N_9926);
xnor UO_119 (O_119,N_9828,N_9938);
xnor UO_120 (O_120,N_9827,N_9834);
and UO_121 (O_121,N_9967,N_9884);
xnor UO_122 (O_122,N_9854,N_9809);
nand UO_123 (O_123,N_9819,N_9998);
or UO_124 (O_124,N_9849,N_9882);
nor UO_125 (O_125,N_9842,N_9812);
xor UO_126 (O_126,N_9904,N_9848);
and UO_127 (O_127,N_9811,N_9961);
and UO_128 (O_128,N_9947,N_9951);
xor UO_129 (O_129,N_9964,N_9856);
nor UO_130 (O_130,N_9914,N_9925);
or UO_131 (O_131,N_9915,N_9985);
and UO_132 (O_132,N_9951,N_9864);
nand UO_133 (O_133,N_9898,N_9887);
and UO_134 (O_134,N_9972,N_9884);
or UO_135 (O_135,N_9949,N_9955);
nor UO_136 (O_136,N_9958,N_9982);
xnor UO_137 (O_137,N_9810,N_9833);
and UO_138 (O_138,N_9862,N_9917);
nor UO_139 (O_139,N_9870,N_9938);
xnor UO_140 (O_140,N_9943,N_9907);
nor UO_141 (O_141,N_9910,N_9952);
xnor UO_142 (O_142,N_9929,N_9816);
nand UO_143 (O_143,N_9996,N_9858);
or UO_144 (O_144,N_9927,N_9848);
nor UO_145 (O_145,N_9979,N_9848);
nand UO_146 (O_146,N_9902,N_9900);
xnor UO_147 (O_147,N_9962,N_9813);
and UO_148 (O_148,N_9930,N_9992);
or UO_149 (O_149,N_9887,N_9872);
nor UO_150 (O_150,N_9802,N_9831);
or UO_151 (O_151,N_9892,N_9950);
nand UO_152 (O_152,N_9974,N_9829);
or UO_153 (O_153,N_9821,N_9869);
and UO_154 (O_154,N_9877,N_9909);
nor UO_155 (O_155,N_9883,N_9830);
and UO_156 (O_156,N_9894,N_9906);
or UO_157 (O_157,N_9946,N_9902);
xor UO_158 (O_158,N_9962,N_9865);
nand UO_159 (O_159,N_9808,N_9943);
nor UO_160 (O_160,N_9889,N_9853);
xor UO_161 (O_161,N_9896,N_9933);
and UO_162 (O_162,N_9849,N_9886);
xnor UO_163 (O_163,N_9952,N_9854);
and UO_164 (O_164,N_9918,N_9953);
or UO_165 (O_165,N_9889,N_9838);
xor UO_166 (O_166,N_9944,N_9892);
and UO_167 (O_167,N_9886,N_9974);
nand UO_168 (O_168,N_9922,N_9944);
nor UO_169 (O_169,N_9835,N_9818);
or UO_170 (O_170,N_9862,N_9803);
nand UO_171 (O_171,N_9926,N_9881);
or UO_172 (O_172,N_9849,N_9892);
nand UO_173 (O_173,N_9933,N_9815);
and UO_174 (O_174,N_9840,N_9973);
and UO_175 (O_175,N_9959,N_9979);
and UO_176 (O_176,N_9825,N_9959);
xor UO_177 (O_177,N_9914,N_9867);
nand UO_178 (O_178,N_9830,N_9910);
xor UO_179 (O_179,N_9855,N_9973);
and UO_180 (O_180,N_9801,N_9806);
and UO_181 (O_181,N_9858,N_9982);
nor UO_182 (O_182,N_9809,N_9862);
and UO_183 (O_183,N_9945,N_9922);
xnor UO_184 (O_184,N_9823,N_9805);
xor UO_185 (O_185,N_9813,N_9897);
xnor UO_186 (O_186,N_9967,N_9951);
or UO_187 (O_187,N_9887,N_9875);
or UO_188 (O_188,N_9816,N_9967);
and UO_189 (O_189,N_9947,N_9980);
xnor UO_190 (O_190,N_9986,N_9804);
xor UO_191 (O_191,N_9816,N_9855);
nor UO_192 (O_192,N_9901,N_9880);
nand UO_193 (O_193,N_9978,N_9839);
nor UO_194 (O_194,N_9872,N_9976);
nand UO_195 (O_195,N_9862,N_9913);
nand UO_196 (O_196,N_9828,N_9883);
or UO_197 (O_197,N_9948,N_9813);
nand UO_198 (O_198,N_9896,N_9818);
xnor UO_199 (O_199,N_9907,N_9962);
nor UO_200 (O_200,N_9972,N_9953);
nor UO_201 (O_201,N_9946,N_9988);
nand UO_202 (O_202,N_9935,N_9835);
nor UO_203 (O_203,N_9984,N_9842);
xnor UO_204 (O_204,N_9905,N_9874);
or UO_205 (O_205,N_9907,N_9847);
nand UO_206 (O_206,N_9984,N_9936);
and UO_207 (O_207,N_9810,N_9921);
xnor UO_208 (O_208,N_9811,N_9905);
and UO_209 (O_209,N_9858,N_9868);
and UO_210 (O_210,N_9915,N_9802);
nor UO_211 (O_211,N_9939,N_9851);
nor UO_212 (O_212,N_9844,N_9804);
xnor UO_213 (O_213,N_9964,N_9831);
or UO_214 (O_214,N_9982,N_9971);
and UO_215 (O_215,N_9930,N_9851);
nand UO_216 (O_216,N_9982,N_9981);
nand UO_217 (O_217,N_9829,N_9969);
nand UO_218 (O_218,N_9917,N_9821);
nor UO_219 (O_219,N_9801,N_9941);
nor UO_220 (O_220,N_9905,N_9817);
xor UO_221 (O_221,N_9882,N_9858);
or UO_222 (O_222,N_9822,N_9976);
and UO_223 (O_223,N_9903,N_9854);
and UO_224 (O_224,N_9805,N_9854);
nand UO_225 (O_225,N_9947,N_9854);
or UO_226 (O_226,N_9960,N_9927);
or UO_227 (O_227,N_9846,N_9898);
nand UO_228 (O_228,N_9819,N_9981);
xnor UO_229 (O_229,N_9850,N_9808);
and UO_230 (O_230,N_9926,N_9813);
xnor UO_231 (O_231,N_9965,N_9981);
and UO_232 (O_232,N_9815,N_9872);
nor UO_233 (O_233,N_9920,N_9963);
or UO_234 (O_234,N_9802,N_9969);
nand UO_235 (O_235,N_9950,N_9875);
or UO_236 (O_236,N_9911,N_9875);
xnor UO_237 (O_237,N_9805,N_9960);
and UO_238 (O_238,N_9805,N_9871);
or UO_239 (O_239,N_9959,N_9983);
xor UO_240 (O_240,N_9974,N_9875);
nor UO_241 (O_241,N_9902,N_9896);
nor UO_242 (O_242,N_9914,N_9833);
xor UO_243 (O_243,N_9891,N_9928);
and UO_244 (O_244,N_9981,N_9815);
nand UO_245 (O_245,N_9832,N_9860);
xor UO_246 (O_246,N_9892,N_9957);
or UO_247 (O_247,N_9932,N_9886);
nor UO_248 (O_248,N_9979,N_9994);
xnor UO_249 (O_249,N_9981,N_9952);
nand UO_250 (O_250,N_9858,N_9957);
or UO_251 (O_251,N_9877,N_9821);
or UO_252 (O_252,N_9830,N_9926);
nor UO_253 (O_253,N_9906,N_9873);
and UO_254 (O_254,N_9824,N_9811);
and UO_255 (O_255,N_9904,N_9930);
xor UO_256 (O_256,N_9910,N_9863);
nand UO_257 (O_257,N_9812,N_9858);
xor UO_258 (O_258,N_9955,N_9993);
xnor UO_259 (O_259,N_9907,N_9909);
or UO_260 (O_260,N_9918,N_9986);
nor UO_261 (O_261,N_9989,N_9958);
or UO_262 (O_262,N_9832,N_9853);
xnor UO_263 (O_263,N_9924,N_9930);
nand UO_264 (O_264,N_9871,N_9823);
and UO_265 (O_265,N_9984,N_9822);
xor UO_266 (O_266,N_9897,N_9984);
and UO_267 (O_267,N_9845,N_9974);
nand UO_268 (O_268,N_9951,N_9956);
nand UO_269 (O_269,N_9848,N_9903);
nand UO_270 (O_270,N_9958,N_9829);
or UO_271 (O_271,N_9845,N_9848);
nand UO_272 (O_272,N_9869,N_9947);
nor UO_273 (O_273,N_9944,N_9856);
xor UO_274 (O_274,N_9834,N_9992);
and UO_275 (O_275,N_9996,N_9820);
nor UO_276 (O_276,N_9833,N_9873);
xor UO_277 (O_277,N_9884,N_9878);
and UO_278 (O_278,N_9861,N_9954);
xnor UO_279 (O_279,N_9866,N_9928);
nor UO_280 (O_280,N_9952,N_9885);
xor UO_281 (O_281,N_9852,N_9993);
nor UO_282 (O_282,N_9917,N_9909);
xnor UO_283 (O_283,N_9934,N_9825);
nand UO_284 (O_284,N_9878,N_9936);
and UO_285 (O_285,N_9871,N_9909);
and UO_286 (O_286,N_9849,N_9975);
nand UO_287 (O_287,N_9983,N_9993);
nand UO_288 (O_288,N_9934,N_9840);
nor UO_289 (O_289,N_9857,N_9957);
and UO_290 (O_290,N_9966,N_9889);
nand UO_291 (O_291,N_9933,N_9873);
and UO_292 (O_292,N_9964,N_9809);
nor UO_293 (O_293,N_9835,N_9884);
xor UO_294 (O_294,N_9845,N_9892);
xor UO_295 (O_295,N_9989,N_9939);
nand UO_296 (O_296,N_9907,N_9804);
xnor UO_297 (O_297,N_9904,N_9818);
nand UO_298 (O_298,N_9926,N_9852);
and UO_299 (O_299,N_9842,N_9823);
xnor UO_300 (O_300,N_9953,N_9995);
and UO_301 (O_301,N_9874,N_9971);
nand UO_302 (O_302,N_9817,N_9867);
nand UO_303 (O_303,N_9853,N_9904);
or UO_304 (O_304,N_9921,N_9814);
nor UO_305 (O_305,N_9856,N_9839);
nor UO_306 (O_306,N_9930,N_9868);
or UO_307 (O_307,N_9961,N_9986);
nor UO_308 (O_308,N_9804,N_9973);
xor UO_309 (O_309,N_9861,N_9884);
xnor UO_310 (O_310,N_9963,N_9953);
nand UO_311 (O_311,N_9985,N_9874);
nand UO_312 (O_312,N_9938,N_9926);
nor UO_313 (O_313,N_9895,N_9947);
nand UO_314 (O_314,N_9938,N_9931);
xnor UO_315 (O_315,N_9857,N_9958);
or UO_316 (O_316,N_9957,N_9846);
nor UO_317 (O_317,N_9808,N_9804);
or UO_318 (O_318,N_9941,N_9986);
or UO_319 (O_319,N_9803,N_9987);
nand UO_320 (O_320,N_9879,N_9895);
nor UO_321 (O_321,N_9867,N_9883);
and UO_322 (O_322,N_9990,N_9923);
or UO_323 (O_323,N_9998,N_9883);
nor UO_324 (O_324,N_9804,N_9966);
nand UO_325 (O_325,N_9848,N_9896);
and UO_326 (O_326,N_9939,N_9909);
or UO_327 (O_327,N_9936,N_9858);
nand UO_328 (O_328,N_9830,N_9870);
nor UO_329 (O_329,N_9956,N_9869);
or UO_330 (O_330,N_9978,N_9880);
and UO_331 (O_331,N_9829,N_9840);
and UO_332 (O_332,N_9972,N_9859);
nand UO_333 (O_333,N_9933,N_9934);
or UO_334 (O_334,N_9892,N_9862);
or UO_335 (O_335,N_9846,N_9961);
nor UO_336 (O_336,N_9862,N_9848);
xor UO_337 (O_337,N_9870,N_9898);
nand UO_338 (O_338,N_9812,N_9815);
and UO_339 (O_339,N_9907,N_9828);
nor UO_340 (O_340,N_9916,N_9800);
and UO_341 (O_341,N_9903,N_9822);
or UO_342 (O_342,N_9994,N_9998);
nand UO_343 (O_343,N_9953,N_9944);
nor UO_344 (O_344,N_9804,N_9829);
and UO_345 (O_345,N_9805,N_9915);
nor UO_346 (O_346,N_9999,N_9949);
xor UO_347 (O_347,N_9847,N_9926);
and UO_348 (O_348,N_9879,N_9802);
nand UO_349 (O_349,N_9998,N_9924);
nand UO_350 (O_350,N_9892,N_9866);
or UO_351 (O_351,N_9841,N_9819);
nand UO_352 (O_352,N_9993,N_9801);
and UO_353 (O_353,N_9979,N_9884);
nand UO_354 (O_354,N_9812,N_9926);
or UO_355 (O_355,N_9814,N_9920);
nand UO_356 (O_356,N_9878,N_9821);
nand UO_357 (O_357,N_9840,N_9814);
or UO_358 (O_358,N_9954,N_9975);
xnor UO_359 (O_359,N_9867,N_9920);
and UO_360 (O_360,N_9949,N_9948);
or UO_361 (O_361,N_9892,N_9821);
and UO_362 (O_362,N_9809,N_9900);
nor UO_363 (O_363,N_9962,N_9978);
and UO_364 (O_364,N_9860,N_9891);
nor UO_365 (O_365,N_9809,N_9810);
or UO_366 (O_366,N_9976,N_9873);
nand UO_367 (O_367,N_9842,N_9923);
xnor UO_368 (O_368,N_9943,N_9902);
or UO_369 (O_369,N_9815,N_9816);
xnor UO_370 (O_370,N_9886,N_9860);
nand UO_371 (O_371,N_9990,N_9921);
nor UO_372 (O_372,N_9832,N_9917);
nor UO_373 (O_373,N_9917,N_9962);
xnor UO_374 (O_374,N_9962,N_9941);
nor UO_375 (O_375,N_9974,N_9901);
nand UO_376 (O_376,N_9950,N_9991);
nor UO_377 (O_377,N_9907,N_9844);
and UO_378 (O_378,N_9804,N_9988);
xor UO_379 (O_379,N_9867,N_9845);
and UO_380 (O_380,N_9878,N_9875);
nor UO_381 (O_381,N_9836,N_9989);
or UO_382 (O_382,N_9931,N_9849);
nor UO_383 (O_383,N_9919,N_9968);
nand UO_384 (O_384,N_9917,N_9930);
nand UO_385 (O_385,N_9883,N_9832);
nand UO_386 (O_386,N_9813,N_9801);
xnor UO_387 (O_387,N_9952,N_9973);
xnor UO_388 (O_388,N_9858,N_9833);
nor UO_389 (O_389,N_9940,N_9857);
or UO_390 (O_390,N_9978,N_9845);
xor UO_391 (O_391,N_9910,N_9844);
xnor UO_392 (O_392,N_9902,N_9986);
nor UO_393 (O_393,N_9996,N_9971);
or UO_394 (O_394,N_9867,N_9826);
nand UO_395 (O_395,N_9994,N_9914);
and UO_396 (O_396,N_9874,N_9904);
nor UO_397 (O_397,N_9862,N_9967);
xor UO_398 (O_398,N_9886,N_9884);
or UO_399 (O_399,N_9966,N_9963);
and UO_400 (O_400,N_9870,N_9811);
or UO_401 (O_401,N_9932,N_9953);
nor UO_402 (O_402,N_9922,N_9908);
or UO_403 (O_403,N_9965,N_9827);
nand UO_404 (O_404,N_9960,N_9833);
and UO_405 (O_405,N_9970,N_9891);
nand UO_406 (O_406,N_9872,N_9908);
xnor UO_407 (O_407,N_9902,N_9973);
or UO_408 (O_408,N_9911,N_9902);
or UO_409 (O_409,N_9895,N_9901);
and UO_410 (O_410,N_9827,N_9993);
xnor UO_411 (O_411,N_9885,N_9886);
nand UO_412 (O_412,N_9846,N_9946);
nor UO_413 (O_413,N_9935,N_9963);
or UO_414 (O_414,N_9807,N_9948);
and UO_415 (O_415,N_9876,N_9963);
nand UO_416 (O_416,N_9984,N_9899);
xnor UO_417 (O_417,N_9921,N_9881);
nor UO_418 (O_418,N_9847,N_9941);
or UO_419 (O_419,N_9930,N_9873);
or UO_420 (O_420,N_9862,N_9878);
and UO_421 (O_421,N_9803,N_9814);
and UO_422 (O_422,N_9931,N_9886);
nand UO_423 (O_423,N_9828,N_9926);
or UO_424 (O_424,N_9880,N_9967);
or UO_425 (O_425,N_9872,N_9813);
or UO_426 (O_426,N_9954,N_9823);
xor UO_427 (O_427,N_9866,N_9952);
or UO_428 (O_428,N_9870,N_9914);
and UO_429 (O_429,N_9994,N_9879);
or UO_430 (O_430,N_9848,N_9886);
xor UO_431 (O_431,N_9841,N_9933);
or UO_432 (O_432,N_9965,N_9948);
and UO_433 (O_433,N_9948,N_9946);
nand UO_434 (O_434,N_9816,N_9840);
xnor UO_435 (O_435,N_9902,N_9907);
and UO_436 (O_436,N_9963,N_9977);
or UO_437 (O_437,N_9902,N_9858);
xnor UO_438 (O_438,N_9860,N_9893);
xor UO_439 (O_439,N_9991,N_9826);
and UO_440 (O_440,N_9882,N_9817);
or UO_441 (O_441,N_9932,N_9893);
nand UO_442 (O_442,N_9935,N_9979);
nand UO_443 (O_443,N_9917,N_9890);
nand UO_444 (O_444,N_9933,N_9883);
nor UO_445 (O_445,N_9805,N_9838);
or UO_446 (O_446,N_9874,N_9984);
nor UO_447 (O_447,N_9856,N_9920);
nor UO_448 (O_448,N_9958,N_9813);
and UO_449 (O_449,N_9957,N_9826);
nand UO_450 (O_450,N_9911,N_9846);
xnor UO_451 (O_451,N_9983,N_9936);
nor UO_452 (O_452,N_9863,N_9871);
nor UO_453 (O_453,N_9825,N_9975);
and UO_454 (O_454,N_9988,N_9838);
nor UO_455 (O_455,N_9830,N_9904);
and UO_456 (O_456,N_9924,N_9912);
xnor UO_457 (O_457,N_9862,N_9965);
and UO_458 (O_458,N_9956,N_9885);
and UO_459 (O_459,N_9853,N_9918);
or UO_460 (O_460,N_9867,N_9981);
nor UO_461 (O_461,N_9829,N_9930);
xor UO_462 (O_462,N_9825,N_9869);
and UO_463 (O_463,N_9804,N_9952);
or UO_464 (O_464,N_9822,N_9847);
nor UO_465 (O_465,N_9989,N_9946);
nor UO_466 (O_466,N_9812,N_9981);
xor UO_467 (O_467,N_9895,N_9991);
nand UO_468 (O_468,N_9880,N_9990);
and UO_469 (O_469,N_9832,N_9890);
or UO_470 (O_470,N_9934,N_9956);
nand UO_471 (O_471,N_9871,N_9870);
or UO_472 (O_472,N_9977,N_9927);
nor UO_473 (O_473,N_9926,N_9832);
nor UO_474 (O_474,N_9924,N_9836);
nand UO_475 (O_475,N_9952,N_9899);
xnor UO_476 (O_476,N_9917,N_9829);
or UO_477 (O_477,N_9981,N_9825);
and UO_478 (O_478,N_9844,N_9954);
nand UO_479 (O_479,N_9864,N_9905);
or UO_480 (O_480,N_9983,N_9986);
xnor UO_481 (O_481,N_9811,N_9862);
xor UO_482 (O_482,N_9890,N_9857);
nor UO_483 (O_483,N_9951,N_9870);
xor UO_484 (O_484,N_9997,N_9887);
nor UO_485 (O_485,N_9908,N_9962);
xnor UO_486 (O_486,N_9943,N_9937);
xnor UO_487 (O_487,N_9974,N_9820);
xnor UO_488 (O_488,N_9918,N_9875);
nand UO_489 (O_489,N_9842,N_9944);
and UO_490 (O_490,N_9948,N_9887);
and UO_491 (O_491,N_9839,N_9964);
nand UO_492 (O_492,N_9904,N_9915);
nand UO_493 (O_493,N_9964,N_9880);
and UO_494 (O_494,N_9921,N_9973);
and UO_495 (O_495,N_9860,N_9840);
or UO_496 (O_496,N_9800,N_9942);
or UO_497 (O_497,N_9856,N_9890);
nand UO_498 (O_498,N_9941,N_9837);
and UO_499 (O_499,N_9999,N_9821);
or UO_500 (O_500,N_9878,N_9990);
and UO_501 (O_501,N_9891,N_9802);
nor UO_502 (O_502,N_9991,N_9840);
or UO_503 (O_503,N_9960,N_9971);
nor UO_504 (O_504,N_9814,N_9939);
nor UO_505 (O_505,N_9965,N_9936);
xnor UO_506 (O_506,N_9868,N_9873);
and UO_507 (O_507,N_9909,N_9966);
nor UO_508 (O_508,N_9853,N_9969);
xor UO_509 (O_509,N_9962,N_9975);
nand UO_510 (O_510,N_9920,N_9828);
and UO_511 (O_511,N_9832,N_9964);
and UO_512 (O_512,N_9952,N_9963);
nor UO_513 (O_513,N_9901,N_9980);
nand UO_514 (O_514,N_9940,N_9946);
nand UO_515 (O_515,N_9862,N_9963);
nor UO_516 (O_516,N_9961,N_9997);
nor UO_517 (O_517,N_9957,N_9939);
nand UO_518 (O_518,N_9801,N_9893);
or UO_519 (O_519,N_9828,N_9955);
and UO_520 (O_520,N_9904,N_9881);
and UO_521 (O_521,N_9869,N_9816);
nor UO_522 (O_522,N_9954,N_9857);
nand UO_523 (O_523,N_9811,N_9904);
nor UO_524 (O_524,N_9969,N_9974);
and UO_525 (O_525,N_9938,N_9913);
nand UO_526 (O_526,N_9974,N_9801);
or UO_527 (O_527,N_9900,N_9894);
and UO_528 (O_528,N_9995,N_9879);
nor UO_529 (O_529,N_9806,N_9981);
xor UO_530 (O_530,N_9845,N_9969);
nor UO_531 (O_531,N_9827,N_9829);
and UO_532 (O_532,N_9955,N_9990);
xnor UO_533 (O_533,N_9895,N_9833);
xor UO_534 (O_534,N_9815,N_9889);
nand UO_535 (O_535,N_9830,N_9932);
and UO_536 (O_536,N_9853,N_9830);
and UO_537 (O_537,N_9840,N_9952);
nor UO_538 (O_538,N_9916,N_9858);
and UO_539 (O_539,N_9809,N_9954);
nand UO_540 (O_540,N_9863,N_9948);
nand UO_541 (O_541,N_9864,N_9843);
nor UO_542 (O_542,N_9917,N_9933);
nor UO_543 (O_543,N_9889,N_9994);
and UO_544 (O_544,N_9919,N_9974);
nor UO_545 (O_545,N_9831,N_9848);
xor UO_546 (O_546,N_9922,N_9936);
or UO_547 (O_547,N_9926,N_9862);
xor UO_548 (O_548,N_9908,N_9900);
xor UO_549 (O_549,N_9891,N_9911);
nand UO_550 (O_550,N_9855,N_9905);
nor UO_551 (O_551,N_9801,N_9986);
nor UO_552 (O_552,N_9881,N_9808);
nand UO_553 (O_553,N_9912,N_9835);
nor UO_554 (O_554,N_9942,N_9935);
xor UO_555 (O_555,N_9895,N_9967);
and UO_556 (O_556,N_9857,N_9880);
nand UO_557 (O_557,N_9806,N_9982);
nor UO_558 (O_558,N_9850,N_9977);
or UO_559 (O_559,N_9975,N_9944);
nand UO_560 (O_560,N_9876,N_9827);
nor UO_561 (O_561,N_9855,N_9953);
nor UO_562 (O_562,N_9906,N_9845);
nand UO_563 (O_563,N_9975,N_9832);
and UO_564 (O_564,N_9856,N_9819);
nor UO_565 (O_565,N_9834,N_9923);
nand UO_566 (O_566,N_9886,N_9955);
nor UO_567 (O_567,N_9939,N_9846);
and UO_568 (O_568,N_9940,N_9981);
or UO_569 (O_569,N_9980,N_9886);
nand UO_570 (O_570,N_9870,N_9952);
xnor UO_571 (O_571,N_9814,N_9894);
or UO_572 (O_572,N_9837,N_9817);
xnor UO_573 (O_573,N_9986,N_9845);
xnor UO_574 (O_574,N_9855,N_9866);
nand UO_575 (O_575,N_9820,N_9873);
xnor UO_576 (O_576,N_9934,N_9845);
nand UO_577 (O_577,N_9925,N_9885);
or UO_578 (O_578,N_9960,N_9822);
xor UO_579 (O_579,N_9952,N_9929);
and UO_580 (O_580,N_9967,N_9905);
nor UO_581 (O_581,N_9849,N_9862);
nand UO_582 (O_582,N_9946,N_9947);
nand UO_583 (O_583,N_9941,N_9973);
nand UO_584 (O_584,N_9950,N_9804);
xnor UO_585 (O_585,N_9845,N_9999);
and UO_586 (O_586,N_9810,N_9918);
xnor UO_587 (O_587,N_9966,N_9954);
nand UO_588 (O_588,N_9918,N_9978);
nor UO_589 (O_589,N_9943,N_9893);
nor UO_590 (O_590,N_9850,N_9828);
and UO_591 (O_591,N_9925,N_9986);
xor UO_592 (O_592,N_9990,N_9847);
or UO_593 (O_593,N_9898,N_9955);
nand UO_594 (O_594,N_9836,N_9840);
nor UO_595 (O_595,N_9858,N_9913);
nor UO_596 (O_596,N_9980,N_9844);
or UO_597 (O_597,N_9995,N_9949);
nand UO_598 (O_598,N_9975,N_9865);
nand UO_599 (O_599,N_9889,N_9876);
nand UO_600 (O_600,N_9812,N_9896);
or UO_601 (O_601,N_9888,N_9822);
nand UO_602 (O_602,N_9807,N_9883);
xnor UO_603 (O_603,N_9913,N_9875);
or UO_604 (O_604,N_9856,N_9961);
xnor UO_605 (O_605,N_9836,N_9912);
xor UO_606 (O_606,N_9994,N_9924);
or UO_607 (O_607,N_9844,N_9918);
and UO_608 (O_608,N_9981,N_9820);
and UO_609 (O_609,N_9800,N_9876);
nor UO_610 (O_610,N_9858,N_9947);
nand UO_611 (O_611,N_9968,N_9879);
nor UO_612 (O_612,N_9852,N_9919);
or UO_613 (O_613,N_9908,N_9974);
nor UO_614 (O_614,N_9875,N_9899);
nand UO_615 (O_615,N_9896,N_9837);
nand UO_616 (O_616,N_9943,N_9868);
and UO_617 (O_617,N_9996,N_9935);
nor UO_618 (O_618,N_9831,N_9961);
nand UO_619 (O_619,N_9912,N_9820);
nor UO_620 (O_620,N_9955,N_9925);
or UO_621 (O_621,N_9818,N_9962);
and UO_622 (O_622,N_9893,N_9914);
xor UO_623 (O_623,N_9840,N_9970);
or UO_624 (O_624,N_9856,N_9923);
nor UO_625 (O_625,N_9909,N_9838);
and UO_626 (O_626,N_9887,N_9846);
and UO_627 (O_627,N_9994,N_9930);
nor UO_628 (O_628,N_9885,N_9838);
or UO_629 (O_629,N_9976,N_9929);
nand UO_630 (O_630,N_9903,N_9948);
nor UO_631 (O_631,N_9835,N_9821);
xnor UO_632 (O_632,N_9984,N_9977);
nand UO_633 (O_633,N_9900,N_9838);
xnor UO_634 (O_634,N_9841,N_9818);
and UO_635 (O_635,N_9876,N_9847);
xnor UO_636 (O_636,N_9954,N_9930);
nand UO_637 (O_637,N_9975,N_9848);
nand UO_638 (O_638,N_9867,N_9830);
or UO_639 (O_639,N_9922,N_9960);
and UO_640 (O_640,N_9899,N_9995);
or UO_641 (O_641,N_9929,N_9989);
nand UO_642 (O_642,N_9875,N_9965);
nand UO_643 (O_643,N_9960,N_9820);
nand UO_644 (O_644,N_9843,N_9831);
nor UO_645 (O_645,N_9854,N_9850);
and UO_646 (O_646,N_9835,N_9915);
xor UO_647 (O_647,N_9977,N_9806);
or UO_648 (O_648,N_9818,N_9837);
or UO_649 (O_649,N_9857,N_9825);
and UO_650 (O_650,N_9850,N_9884);
xor UO_651 (O_651,N_9806,N_9983);
nand UO_652 (O_652,N_9990,N_9943);
nor UO_653 (O_653,N_9863,N_9912);
and UO_654 (O_654,N_9869,N_9925);
xor UO_655 (O_655,N_9906,N_9996);
or UO_656 (O_656,N_9944,N_9815);
nand UO_657 (O_657,N_9918,N_9965);
nor UO_658 (O_658,N_9927,N_9943);
or UO_659 (O_659,N_9867,N_9828);
nor UO_660 (O_660,N_9829,N_9927);
and UO_661 (O_661,N_9896,N_9956);
xnor UO_662 (O_662,N_9873,N_9977);
or UO_663 (O_663,N_9995,N_9938);
or UO_664 (O_664,N_9843,N_9847);
or UO_665 (O_665,N_9862,N_9843);
and UO_666 (O_666,N_9849,N_9891);
nand UO_667 (O_667,N_9935,N_9853);
xor UO_668 (O_668,N_9901,N_9931);
xor UO_669 (O_669,N_9950,N_9976);
xor UO_670 (O_670,N_9996,N_9907);
nor UO_671 (O_671,N_9904,N_9868);
or UO_672 (O_672,N_9952,N_9894);
nand UO_673 (O_673,N_9822,N_9897);
nor UO_674 (O_674,N_9914,N_9986);
or UO_675 (O_675,N_9974,N_9967);
nor UO_676 (O_676,N_9911,N_9964);
nor UO_677 (O_677,N_9878,N_9928);
xor UO_678 (O_678,N_9999,N_9842);
xnor UO_679 (O_679,N_9897,N_9847);
nor UO_680 (O_680,N_9917,N_9898);
nor UO_681 (O_681,N_9863,N_9919);
nor UO_682 (O_682,N_9848,N_9952);
xor UO_683 (O_683,N_9837,N_9800);
nand UO_684 (O_684,N_9838,N_9946);
xnor UO_685 (O_685,N_9969,N_9905);
xor UO_686 (O_686,N_9978,N_9965);
or UO_687 (O_687,N_9857,N_9897);
or UO_688 (O_688,N_9913,N_9838);
nand UO_689 (O_689,N_9833,N_9812);
xnor UO_690 (O_690,N_9868,N_9988);
xnor UO_691 (O_691,N_9965,N_9892);
nor UO_692 (O_692,N_9815,N_9923);
and UO_693 (O_693,N_9899,N_9832);
or UO_694 (O_694,N_9801,N_9970);
nor UO_695 (O_695,N_9936,N_9874);
nor UO_696 (O_696,N_9899,N_9908);
nand UO_697 (O_697,N_9800,N_9899);
nor UO_698 (O_698,N_9960,N_9964);
nor UO_699 (O_699,N_9855,N_9823);
and UO_700 (O_700,N_9966,N_9829);
xor UO_701 (O_701,N_9867,N_9868);
xnor UO_702 (O_702,N_9829,N_9801);
or UO_703 (O_703,N_9948,N_9872);
nand UO_704 (O_704,N_9842,N_9929);
nand UO_705 (O_705,N_9971,N_9938);
and UO_706 (O_706,N_9943,N_9968);
nor UO_707 (O_707,N_9951,N_9843);
and UO_708 (O_708,N_9920,N_9823);
nor UO_709 (O_709,N_9971,N_9955);
and UO_710 (O_710,N_9887,N_9843);
xnor UO_711 (O_711,N_9832,N_9881);
nand UO_712 (O_712,N_9961,N_9828);
xnor UO_713 (O_713,N_9904,N_9836);
nand UO_714 (O_714,N_9946,N_9866);
xor UO_715 (O_715,N_9925,N_9827);
and UO_716 (O_716,N_9857,N_9997);
and UO_717 (O_717,N_9997,N_9941);
and UO_718 (O_718,N_9951,N_9913);
or UO_719 (O_719,N_9834,N_9857);
nor UO_720 (O_720,N_9929,N_9801);
or UO_721 (O_721,N_9804,N_9971);
nand UO_722 (O_722,N_9826,N_9903);
xnor UO_723 (O_723,N_9812,N_9898);
or UO_724 (O_724,N_9938,N_9891);
xnor UO_725 (O_725,N_9843,N_9852);
xor UO_726 (O_726,N_9984,N_9870);
xor UO_727 (O_727,N_9884,N_9806);
and UO_728 (O_728,N_9829,N_9897);
nor UO_729 (O_729,N_9908,N_9927);
and UO_730 (O_730,N_9878,N_9958);
or UO_731 (O_731,N_9800,N_9917);
xor UO_732 (O_732,N_9885,N_9875);
nor UO_733 (O_733,N_9820,N_9806);
nand UO_734 (O_734,N_9949,N_9903);
nor UO_735 (O_735,N_9899,N_9999);
and UO_736 (O_736,N_9848,N_9840);
xnor UO_737 (O_737,N_9892,N_9909);
and UO_738 (O_738,N_9971,N_9818);
nor UO_739 (O_739,N_9937,N_9834);
nor UO_740 (O_740,N_9870,N_9850);
xor UO_741 (O_741,N_9958,N_9904);
or UO_742 (O_742,N_9831,N_9821);
and UO_743 (O_743,N_9991,N_9944);
and UO_744 (O_744,N_9903,N_9995);
nand UO_745 (O_745,N_9909,N_9927);
nor UO_746 (O_746,N_9830,N_9806);
xor UO_747 (O_747,N_9883,N_9902);
nand UO_748 (O_748,N_9937,N_9855);
or UO_749 (O_749,N_9846,N_9830);
and UO_750 (O_750,N_9955,N_9808);
xnor UO_751 (O_751,N_9822,N_9881);
nand UO_752 (O_752,N_9954,N_9805);
nor UO_753 (O_753,N_9903,N_9878);
xor UO_754 (O_754,N_9815,N_9857);
or UO_755 (O_755,N_9939,N_9949);
xor UO_756 (O_756,N_9968,N_9888);
xnor UO_757 (O_757,N_9986,N_9892);
nor UO_758 (O_758,N_9847,N_9840);
xor UO_759 (O_759,N_9991,N_9837);
nand UO_760 (O_760,N_9885,N_9884);
or UO_761 (O_761,N_9991,N_9934);
nor UO_762 (O_762,N_9841,N_9815);
nor UO_763 (O_763,N_9878,N_9851);
nor UO_764 (O_764,N_9868,N_9955);
and UO_765 (O_765,N_9812,N_9839);
nor UO_766 (O_766,N_9890,N_9990);
nor UO_767 (O_767,N_9887,N_9892);
nand UO_768 (O_768,N_9965,N_9959);
nor UO_769 (O_769,N_9950,N_9888);
nand UO_770 (O_770,N_9967,N_9920);
nand UO_771 (O_771,N_9903,N_9924);
xor UO_772 (O_772,N_9924,N_9895);
xnor UO_773 (O_773,N_9995,N_9887);
or UO_774 (O_774,N_9837,N_9884);
nand UO_775 (O_775,N_9834,N_9917);
or UO_776 (O_776,N_9837,N_9894);
nand UO_777 (O_777,N_9805,N_9815);
xnor UO_778 (O_778,N_9892,N_9813);
and UO_779 (O_779,N_9980,N_9907);
xor UO_780 (O_780,N_9894,N_9918);
xor UO_781 (O_781,N_9834,N_9803);
xnor UO_782 (O_782,N_9884,N_9946);
nor UO_783 (O_783,N_9950,N_9935);
xor UO_784 (O_784,N_9861,N_9838);
and UO_785 (O_785,N_9847,N_9934);
or UO_786 (O_786,N_9949,N_9828);
nand UO_787 (O_787,N_9891,N_9838);
or UO_788 (O_788,N_9880,N_9887);
and UO_789 (O_789,N_9919,N_9803);
nand UO_790 (O_790,N_9982,N_9865);
nand UO_791 (O_791,N_9888,N_9813);
xnor UO_792 (O_792,N_9859,N_9835);
nand UO_793 (O_793,N_9947,N_9993);
nor UO_794 (O_794,N_9982,N_9991);
and UO_795 (O_795,N_9983,N_9962);
xnor UO_796 (O_796,N_9801,N_9821);
or UO_797 (O_797,N_9908,N_9966);
nor UO_798 (O_798,N_9973,N_9836);
and UO_799 (O_799,N_9877,N_9932);
or UO_800 (O_800,N_9886,N_9893);
or UO_801 (O_801,N_9957,N_9909);
nor UO_802 (O_802,N_9815,N_9947);
nor UO_803 (O_803,N_9878,N_9930);
or UO_804 (O_804,N_9956,N_9901);
and UO_805 (O_805,N_9803,N_9846);
xor UO_806 (O_806,N_9904,N_9936);
and UO_807 (O_807,N_9889,N_9942);
xor UO_808 (O_808,N_9920,N_9927);
nand UO_809 (O_809,N_9806,N_9802);
or UO_810 (O_810,N_9855,N_9925);
and UO_811 (O_811,N_9800,N_9877);
nor UO_812 (O_812,N_9830,N_9985);
nand UO_813 (O_813,N_9975,N_9906);
xor UO_814 (O_814,N_9927,N_9823);
xor UO_815 (O_815,N_9813,N_9981);
or UO_816 (O_816,N_9823,N_9993);
nor UO_817 (O_817,N_9936,N_9952);
xor UO_818 (O_818,N_9815,N_9806);
nand UO_819 (O_819,N_9936,N_9941);
nand UO_820 (O_820,N_9835,N_9869);
or UO_821 (O_821,N_9970,N_9931);
xnor UO_822 (O_822,N_9868,N_9848);
nor UO_823 (O_823,N_9908,N_9977);
or UO_824 (O_824,N_9831,N_9994);
or UO_825 (O_825,N_9951,N_9848);
or UO_826 (O_826,N_9976,N_9889);
and UO_827 (O_827,N_9958,N_9834);
xnor UO_828 (O_828,N_9933,N_9859);
nand UO_829 (O_829,N_9820,N_9983);
xnor UO_830 (O_830,N_9872,N_9899);
and UO_831 (O_831,N_9819,N_9839);
nand UO_832 (O_832,N_9826,N_9887);
and UO_833 (O_833,N_9842,N_9858);
or UO_834 (O_834,N_9818,N_9845);
nor UO_835 (O_835,N_9923,N_9882);
xnor UO_836 (O_836,N_9803,N_9907);
and UO_837 (O_837,N_9859,N_9951);
nor UO_838 (O_838,N_9903,N_9933);
or UO_839 (O_839,N_9988,N_9858);
and UO_840 (O_840,N_9886,N_9814);
nand UO_841 (O_841,N_9829,N_9952);
and UO_842 (O_842,N_9855,N_9892);
nor UO_843 (O_843,N_9950,N_9984);
and UO_844 (O_844,N_9983,N_9991);
nor UO_845 (O_845,N_9921,N_9831);
and UO_846 (O_846,N_9838,N_9977);
xor UO_847 (O_847,N_9818,N_9875);
nor UO_848 (O_848,N_9815,N_9824);
or UO_849 (O_849,N_9935,N_9818);
nor UO_850 (O_850,N_9974,N_9873);
or UO_851 (O_851,N_9887,N_9847);
nand UO_852 (O_852,N_9968,N_9908);
and UO_853 (O_853,N_9961,N_9908);
nor UO_854 (O_854,N_9994,N_9997);
nor UO_855 (O_855,N_9982,N_9825);
or UO_856 (O_856,N_9952,N_9992);
nand UO_857 (O_857,N_9875,N_9908);
or UO_858 (O_858,N_9919,N_9995);
or UO_859 (O_859,N_9936,N_9906);
or UO_860 (O_860,N_9982,N_9812);
nor UO_861 (O_861,N_9955,N_9961);
and UO_862 (O_862,N_9977,N_9855);
xor UO_863 (O_863,N_9964,N_9812);
nand UO_864 (O_864,N_9935,N_9898);
or UO_865 (O_865,N_9844,N_9953);
nor UO_866 (O_866,N_9914,N_9935);
or UO_867 (O_867,N_9846,N_9884);
nand UO_868 (O_868,N_9883,N_9931);
xor UO_869 (O_869,N_9910,N_9914);
and UO_870 (O_870,N_9942,N_9961);
and UO_871 (O_871,N_9880,N_9810);
nor UO_872 (O_872,N_9995,N_9924);
nand UO_873 (O_873,N_9828,N_9927);
or UO_874 (O_874,N_9972,N_9841);
and UO_875 (O_875,N_9833,N_9887);
nor UO_876 (O_876,N_9860,N_9943);
nor UO_877 (O_877,N_9838,N_9881);
nor UO_878 (O_878,N_9837,N_9863);
xor UO_879 (O_879,N_9812,N_9861);
nor UO_880 (O_880,N_9980,N_9847);
or UO_881 (O_881,N_9937,N_9896);
or UO_882 (O_882,N_9900,N_9988);
and UO_883 (O_883,N_9875,N_9872);
nand UO_884 (O_884,N_9812,N_9999);
and UO_885 (O_885,N_9851,N_9877);
and UO_886 (O_886,N_9900,N_9923);
and UO_887 (O_887,N_9854,N_9971);
or UO_888 (O_888,N_9839,N_9958);
or UO_889 (O_889,N_9911,N_9835);
and UO_890 (O_890,N_9831,N_9864);
nand UO_891 (O_891,N_9890,N_9930);
nand UO_892 (O_892,N_9913,N_9857);
nor UO_893 (O_893,N_9995,N_9943);
xnor UO_894 (O_894,N_9826,N_9975);
nand UO_895 (O_895,N_9813,N_9889);
or UO_896 (O_896,N_9976,N_9860);
and UO_897 (O_897,N_9837,N_9848);
or UO_898 (O_898,N_9860,N_9956);
xnor UO_899 (O_899,N_9929,N_9834);
xnor UO_900 (O_900,N_9839,N_9920);
nor UO_901 (O_901,N_9995,N_9980);
nor UO_902 (O_902,N_9824,N_9934);
nand UO_903 (O_903,N_9960,N_9967);
and UO_904 (O_904,N_9864,N_9915);
nand UO_905 (O_905,N_9942,N_9909);
nor UO_906 (O_906,N_9865,N_9972);
xor UO_907 (O_907,N_9941,N_9811);
xnor UO_908 (O_908,N_9944,N_9831);
or UO_909 (O_909,N_9997,N_9899);
or UO_910 (O_910,N_9802,N_9884);
and UO_911 (O_911,N_9906,N_9898);
xor UO_912 (O_912,N_9832,N_9983);
nand UO_913 (O_913,N_9872,N_9878);
or UO_914 (O_914,N_9823,N_9849);
nand UO_915 (O_915,N_9956,N_9886);
nor UO_916 (O_916,N_9850,N_9887);
nor UO_917 (O_917,N_9990,N_9962);
xnor UO_918 (O_918,N_9824,N_9914);
nor UO_919 (O_919,N_9854,N_9835);
xnor UO_920 (O_920,N_9810,N_9879);
nor UO_921 (O_921,N_9992,N_9936);
or UO_922 (O_922,N_9901,N_9816);
nor UO_923 (O_923,N_9943,N_9852);
nand UO_924 (O_924,N_9930,N_9974);
and UO_925 (O_925,N_9925,N_9848);
nand UO_926 (O_926,N_9932,N_9990);
xor UO_927 (O_927,N_9927,N_9957);
nor UO_928 (O_928,N_9964,N_9817);
nand UO_929 (O_929,N_9865,N_9918);
nor UO_930 (O_930,N_9884,N_9866);
nand UO_931 (O_931,N_9973,N_9978);
xor UO_932 (O_932,N_9914,N_9835);
nor UO_933 (O_933,N_9888,N_9959);
xor UO_934 (O_934,N_9869,N_9908);
or UO_935 (O_935,N_9842,N_9866);
and UO_936 (O_936,N_9966,N_9946);
xnor UO_937 (O_937,N_9946,N_9919);
nor UO_938 (O_938,N_9917,N_9841);
and UO_939 (O_939,N_9857,N_9922);
nor UO_940 (O_940,N_9834,N_9915);
and UO_941 (O_941,N_9829,N_9871);
or UO_942 (O_942,N_9872,N_9913);
nand UO_943 (O_943,N_9821,N_9966);
or UO_944 (O_944,N_9850,N_9868);
nand UO_945 (O_945,N_9886,N_9824);
nor UO_946 (O_946,N_9814,N_9969);
nand UO_947 (O_947,N_9858,N_9918);
nor UO_948 (O_948,N_9953,N_9997);
nand UO_949 (O_949,N_9891,N_9997);
or UO_950 (O_950,N_9834,N_9822);
and UO_951 (O_951,N_9846,N_9879);
xnor UO_952 (O_952,N_9817,N_9842);
nand UO_953 (O_953,N_9876,N_9804);
nor UO_954 (O_954,N_9927,N_9889);
or UO_955 (O_955,N_9822,N_9883);
or UO_956 (O_956,N_9964,N_9894);
or UO_957 (O_957,N_9809,N_9831);
nand UO_958 (O_958,N_9914,N_9827);
nand UO_959 (O_959,N_9987,N_9973);
nor UO_960 (O_960,N_9849,N_9820);
and UO_961 (O_961,N_9972,N_9905);
or UO_962 (O_962,N_9820,N_9956);
or UO_963 (O_963,N_9912,N_9882);
and UO_964 (O_964,N_9889,N_9879);
nor UO_965 (O_965,N_9831,N_9878);
and UO_966 (O_966,N_9918,N_9956);
or UO_967 (O_967,N_9958,N_9860);
nor UO_968 (O_968,N_9969,N_9811);
nand UO_969 (O_969,N_9901,N_9841);
nor UO_970 (O_970,N_9920,N_9883);
or UO_971 (O_971,N_9901,N_9876);
or UO_972 (O_972,N_9869,N_9811);
and UO_973 (O_973,N_9975,N_9928);
nand UO_974 (O_974,N_9932,N_9801);
nor UO_975 (O_975,N_9923,N_9938);
and UO_976 (O_976,N_9854,N_9818);
nand UO_977 (O_977,N_9803,N_9832);
xor UO_978 (O_978,N_9998,N_9800);
nand UO_979 (O_979,N_9895,N_9897);
and UO_980 (O_980,N_9940,N_9886);
xnor UO_981 (O_981,N_9903,N_9939);
nand UO_982 (O_982,N_9824,N_9879);
nand UO_983 (O_983,N_9871,N_9804);
nand UO_984 (O_984,N_9917,N_9997);
nor UO_985 (O_985,N_9920,N_9954);
nor UO_986 (O_986,N_9961,N_9851);
nand UO_987 (O_987,N_9896,N_9872);
nand UO_988 (O_988,N_9834,N_9840);
nor UO_989 (O_989,N_9986,N_9999);
and UO_990 (O_990,N_9839,N_9859);
or UO_991 (O_991,N_9909,N_9945);
nand UO_992 (O_992,N_9931,N_9803);
and UO_993 (O_993,N_9905,N_9949);
nor UO_994 (O_994,N_9887,N_9842);
xnor UO_995 (O_995,N_9944,N_9804);
xnor UO_996 (O_996,N_9834,N_9843);
xor UO_997 (O_997,N_9980,N_9915);
nor UO_998 (O_998,N_9949,N_9804);
xnor UO_999 (O_999,N_9817,N_9955);
nand UO_1000 (O_1000,N_9956,N_9841);
xor UO_1001 (O_1001,N_9853,N_9927);
and UO_1002 (O_1002,N_9863,N_9880);
xor UO_1003 (O_1003,N_9890,N_9863);
xnor UO_1004 (O_1004,N_9809,N_9807);
xnor UO_1005 (O_1005,N_9984,N_9812);
or UO_1006 (O_1006,N_9823,N_9868);
nor UO_1007 (O_1007,N_9865,N_9886);
nor UO_1008 (O_1008,N_9884,N_9862);
nor UO_1009 (O_1009,N_9984,N_9853);
or UO_1010 (O_1010,N_9967,N_9879);
xnor UO_1011 (O_1011,N_9930,N_9900);
nand UO_1012 (O_1012,N_9816,N_9968);
and UO_1013 (O_1013,N_9828,N_9837);
and UO_1014 (O_1014,N_9971,N_9909);
nor UO_1015 (O_1015,N_9912,N_9885);
nand UO_1016 (O_1016,N_9989,N_9969);
nor UO_1017 (O_1017,N_9858,N_9870);
xnor UO_1018 (O_1018,N_9845,N_9879);
nor UO_1019 (O_1019,N_9852,N_9908);
nand UO_1020 (O_1020,N_9937,N_9830);
nor UO_1021 (O_1021,N_9919,N_9808);
or UO_1022 (O_1022,N_9879,N_9886);
xor UO_1023 (O_1023,N_9841,N_9837);
nand UO_1024 (O_1024,N_9939,N_9826);
xor UO_1025 (O_1025,N_9942,N_9989);
nor UO_1026 (O_1026,N_9985,N_9980);
nor UO_1027 (O_1027,N_9923,N_9854);
nor UO_1028 (O_1028,N_9897,N_9842);
xor UO_1029 (O_1029,N_9863,N_9865);
and UO_1030 (O_1030,N_9980,N_9822);
or UO_1031 (O_1031,N_9964,N_9969);
or UO_1032 (O_1032,N_9988,N_9932);
xnor UO_1033 (O_1033,N_9834,N_9971);
xor UO_1034 (O_1034,N_9873,N_9965);
nand UO_1035 (O_1035,N_9963,N_9946);
xor UO_1036 (O_1036,N_9813,N_9938);
nand UO_1037 (O_1037,N_9972,N_9821);
nor UO_1038 (O_1038,N_9956,N_9965);
and UO_1039 (O_1039,N_9871,N_9993);
nand UO_1040 (O_1040,N_9873,N_9981);
nand UO_1041 (O_1041,N_9874,N_9800);
nor UO_1042 (O_1042,N_9814,N_9878);
xor UO_1043 (O_1043,N_9934,N_9897);
nor UO_1044 (O_1044,N_9847,N_9905);
nor UO_1045 (O_1045,N_9949,N_9922);
or UO_1046 (O_1046,N_9854,N_9994);
nor UO_1047 (O_1047,N_9896,N_9905);
or UO_1048 (O_1048,N_9806,N_9991);
nor UO_1049 (O_1049,N_9933,N_9988);
or UO_1050 (O_1050,N_9926,N_9986);
nand UO_1051 (O_1051,N_9930,N_9918);
and UO_1052 (O_1052,N_9863,N_9963);
nand UO_1053 (O_1053,N_9860,N_9836);
xor UO_1054 (O_1054,N_9922,N_9891);
nand UO_1055 (O_1055,N_9800,N_9875);
and UO_1056 (O_1056,N_9960,N_9885);
or UO_1057 (O_1057,N_9940,N_9903);
or UO_1058 (O_1058,N_9986,N_9963);
nor UO_1059 (O_1059,N_9851,N_9974);
xnor UO_1060 (O_1060,N_9986,N_9995);
or UO_1061 (O_1061,N_9865,N_9984);
and UO_1062 (O_1062,N_9878,N_9933);
xor UO_1063 (O_1063,N_9972,N_9941);
nor UO_1064 (O_1064,N_9901,N_9848);
or UO_1065 (O_1065,N_9994,N_9825);
nor UO_1066 (O_1066,N_9981,N_9829);
and UO_1067 (O_1067,N_9835,N_9971);
xor UO_1068 (O_1068,N_9950,N_9800);
nand UO_1069 (O_1069,N_9953,N_9852);
xnor UO_1070 (O_1070,N_9814,N_9883);
nor UO_1071 (O_1071,N_9801,N_9906);
or UO_1072 (O_1072,N_9894,N_9956);
xor UO_1073 (O_1073,N_9805,N_9863);
or UO_1074 (O_1074,N_9886,N_9970);
and UO_1075 (O_1075,N_9884,N_9934);
nand UO_1076 (O_1076,N_9901,N_9808);
xor UO_1077 (O_1077,N_9940,N_9825);
or UO_1078 (O_1078,N_9910,N_9866);
and UO_1079 (O_1079,N_9843,N_9990);
xnor UO_1080 (O_1080,N_9909,N_9873);
nand UO_1081 (O_1081,N_9934,N_9849);
nand UO_1082 (O_1082,N_9935,N_9837);
nand UO_1083 (O_1083,N_9933,N_9997);
or UO_1084 (O_1084,N_9848,N_9964);
nand UO_1085 (O_1085,N_9840,N_9911);
xnor UO_1086 (O_1086,N_9846,N_9917);
or UO_1087 (O_1087,N_9860,N_9930);
xnor UO_1088 (O_1088,N_9942,N_9918);
nor UO_1089 (O_1089,N_9827,N_9944);
or UO_1090 (O_1090,N_9963,N_9821);
nand UO_1091 (O_1091,N_9921,N_9897);
xor UO_1092 (O_1092,N_9984,N_9807);
xnor UO_1093 (O_1093,N_9812,N_9994);
xor UO_1094 (O_1094,N_9883,N_9910);
nand UO_1095 (O_1095,N_9803,N_9817);
nor UO_1096 (O_1096,N_9957,N_9972);
or UO_1097 (O_1097,N_9878,N_9829);
and UO_1098 (O_1098,N_9861,N_9902);
xor UO_1099 (O_1099,N_9994,N_9833);
and UO_1100 (O_1100,N_9944,N_9970);
and UO_1101 (O_1101,N_9916,N_9880);
nor UO_1102 (O_1102,N_9958,N_9852);
nand UO_1103 (O_1103,N_9842,N_9822);
nor UO_1104 (O_1104,N_9840,N_9871);
and UO_1105 (O_1105,N_9968,N_9858);
nor UO_1106 (O_1106,N_9993,N_9838);
nand UO_1107 (O_1107,N_9833,N_9973);
or UO_1108 (O_1108,N_9826,N_9983);
nor UO_1109 (O_1109,N_9972,N_9834);
or UO_1110 (O_1110,N_9971,N_9936);
or UO_1111 (O_1111,N_9993,N_9894);
nand UO_1112 (O_1112,N_9835,N_9814);
nand UO_1113 (O_1113,N_9983,N_9904);
or UO_1114 (O_1114,N_9821,N_9953);
or UO_1115 (O_1115,N_9877,N_9848);
nor UO_1116 (O_1116,N_9966,N_9994);
nor UO_1117 (O_1117,N_9990,N_9860);
nand UO_1118 (O_1118,N_9982,N_9844);
nand UO_1119 (O_1119,N_9855,N_9820);
xnor UO_1120 (O_1120,N_9910,N_9865);
xor UO_1121 (O_1121,N_9879,N_9933);
or UO_1122 (O_1122,N_9972,N_9993);
nand UO_1123 (O_1123,N_9899,N_9940);
and UO_1124 (O_1124,N_9913,N_9897);
nand UO_1125 (O_1125,N_9836,N_9842);
nor UO_1126 (O_1126,N_9977,N_9988);
and UO_1127 (O_1127,N_9827,N_9901);
nor UO_1128 (O_1128,N_9940,N_9879);
or UO_1129 (O_1129,N_9944,N_9809);
nor UO_1130 (O_1130,N_9994,N_9947);
nor UO_1131 (O_1131,N_9805,N_9989);
nand UO_1132 (O_1132,N_9904,N_9914);
nand UO_1133 (O_1133,N_9983,N_9813);
nor UO_1134 (O_1134,N_9909,N_9801);
nand UO_1135 (O_1135,N_9948,N_9861);
or UO_1136 (O_1136,N_9879,N_9937);
or UO_1137 (O_1137,N_9895,N_9893);
nor UO_1138 (O_1138,N_9900,N_9881);
nand UO_1139 (O_1139,N_9845,N_9870);
nand UO_1140 (O_1140,N_9821,N_9887);
or UO_1141 (O_1141,N_9898,N_9852);
nand UO_1142 (O_1142,N_9874,N_9969);
xnor UO_1143 (O_1143,N_9804,N_9893);
xor UO_1144 (O_1144,N_9886,N_9877);
and UO_1145 (O_1145,N_9836,N_9919);
xnor UO_1146 (O_1146,N_9816,N_9943);
nor UO_1147 (O_1147,N_9813,N_9809);
or UO_1148 (O_1148,N_9995,N_9841);
nand UO_1149 (O_1149,N_9921,N_9841);
nand UO_1150 (O_1150,N_9816,N_9818);
and UO_1151 (O_1151,N_9926,N_9944);
xor UO_1152 (O_1152,N_9979,N_9827);
nor UO_1153 (O_1153,N_9920,N_9899);
nor UO_1154 (O_1154,N_9811,N_9984);
and UO_1155 (O_1155,N_9813,N_9840);
or UO_1156 (O_1156,N_9836,N_9903);
and UO_1157 (O_1157,N_9977,N_9818);
nand UO_1158 (O_1158,N_9824,N_9917);
and UO_1159 (O_1159,N_9818,N_9849);
and UO_1160 (O_1160,N_9823,N_9912);
nand UO_1161 (O_1161,N_9999,N_9944);
and UO_1162 (O_1162,N_9895,N_9965);
nand UO_1163 (O_1163,N_9873,N_9851);
xor UO_1164 (O_1164,N_9958,N_9833);
xnor UO_1165 (O_1165,N_9952,N_9851);
and UO_1166 (O_1166,N_9913,N_9883);
and UO_1167 (O_1167,N_9952,N_9930);
and UO_1168 (O_1168,N_9980,N_9938);
xor UO_1169 (O_1169,N_9965,N_9879);
xnor UO_1170 (O_1170,N_9941,N_9905);
or UO_1171 (O_1171,N_9889,N_9921);
or UO_1172 (O_1172,N_9830,N_9851);
nand UO_1173 (O_1173,N_9963,N_9940);
or UO_1174 (O_1174,N_9944,N_9980);
nand UO_1175 (O_1175,N_9860,N_9848);
xnor UO_1176 (O_1176,N_9863,N_9958);
xor UO_1177 (O_1177,N_9999,N_9826);
and UO_1178 (O_1178,N_9992,N_9883);
xor UO_1179 (O_1179,N_9904,N_9841);
nor UO_1180 (O_1180,N_9804,N_9912);
and UO_1181 (O_1181,N_9845,N_9832);
and UO_1182 (O_1182,N_9993,N_9954);
or UO_1183 (O_1183,N_9843,N_9928);
nor UO_1184 (O_1184,N_9966,N_9935);
xnor UO_1185 (O_1185,N_9818,N_9914);
xnor UO_1186 (O_1186,N_9942,N_9845);
xnor UO_1187 (O_1187,N_9871,N_9878);
and UO_1188 (O_1188,N_9838,N_9942);
nand UO_1189 (O_1189,N_9951,N_9994);
nor UO_1190 (O_1190,N_9948,N_9855);
nand UO_1191 (O_1191,N_9930,N_9911);
nor UO_1192 (O_1192,N_9984,N_9806);
nor UO_1193 (O_1193,N_9847,N_9995);
and UO_1194 (O_1194,N_9939,N_9908);
or UO_1195 (O_1195,N_9864,N_9821);
and UO_1196 (O_1196,N_9973,N_9955);
nand UO_1197 (O_1197,N_9827,N_9954);
nand UO_1198 (O_1198,N_9955,N_9934);
nand UO_1199 (O_1199,N_9938,N_9893);
nand UO_1200 (O_1200,N_9950,N_9955);
xor UO_1201 (O_1201,N_9940,N_9993);
nand UO_1202 (O_1202,N_9918,N_9912);
nand UO_1203 (O_1203,N_9900,N_9861);
and UO_1204 (O_1204,N_9860,N_9959);
nand UO_1205 (O_1205,N_9964,N_9982);
nand UO_1206 (O_1206,N_9935,N_9940);
xor UO_1207 (O_1207,N_9849,N_9898);
nand UO_1208 (O_1208,N_9941,N_9886);
and UO_1209 (O_1209,N_9808,N_9835);
nand UO_1210 (O_1210,N_9844,N_9864);
nor UO_1211 (O_1211,N_9967,N_9938);
and UO_1212 (O_1212,N_9910,N_9818);
nor UO_1213 (O_1213,N_9820,N_9881);
and UO_1214 (O_1214,N_9901,N_9983);
xnor UO_1215 (O_1215,N_9828,N_9921);
or UO_1216 (O_1216,N_9918,N_9982);
nor UO_1217 (O_1217,N_9999,N_9848);
nor UO_1218 (O_1218,N_9964,N_9873);
nor UO_1219 (O_1219,N_9977,N_9986);
xnor UO_1220 (O_1220,N_9863,N_9997);
nand UO_1221 (O_1221,N_9905,N_9912);
nand UO_1222 (O_1222,N_9818,N_9916);
xor UO_1223 (O_1223,N_9868,N_9900);
or UO_1224 (O_1224,N_9937,N_9911);
xor UO_1225 (O_1225,N_9997,N_9851);
xnor UO_1226 (O_1226,N_9948,N_9805);
and UO_1227 (O_1227,N_9905,N_9868);
nor UO_1228 (O_1228,N_9857,N_9858);
or UO_1229 (O_1229,N_9948,N_9822);
and UO_1230 (O_1230,N_9880,N_9853);
xnor UO_1231 (O_1231,N_9968,N_9904);
or UO_1232 (O_1232,N_9817,N_9982);
or UO_1233 (O_1233,N_9916,N_9805);
nor UO_1234 (O_1234,N_9880,N_9975);
and UO_1235 (O_1235,N_9826,N_9850);
xor UO_1236 (O_1236,N_9901,N_9914);
nand UO_1237 (O_1237,N_9932,N_9840);
nor UO_1238 (O_1238,N_9813,N_9905);
or UO_1239 (O_1239,N_9970,N_9928);
and UO_1240 (O_1240,N_9961,N_9805);
and UO_1241 (O_1241,N_9938,N_9856);
or UO_1242 (O_1242,N_9864,N_9908);
xor UO_1243 (O_1243,N_9865,N_9983);
xor UO_1244 (O_1244,N_9870,N_9837);
xor UO_1245 (O_1245,N_9913,N_9918);
nand UO_1246 (O_1246,N_9923,N_9976);
and UO_1247 (O_1247,N_9876,N_9971);
xor UO_1248 (O_1248,N_9856,N_9992);
xor UO_1249 (O_1249,N_9867,N_9838);
or UO_1250 (O_1250,N_9983,N_9920);
or UO_1251 (O_1251,N_9873,N_9925);
or UO_1252 (O_1252,N_9803,N_9805);
and UO_1253 (O_1253,N_9839,N_9929);
nand UO_1254 (O_1254,N_9941,N_9918);
and UO_1255 (O_1255,N_9875,N_9980);
or UO_1256 (O_1256,N_9808,N_9938);
and UO_1257 (O_1257,N_9912,N_9906);
xnor UO_1258 (O_1258,N_9992,N_9977);
or UO_1259 (O_1259,N_9854,N_9817);
or UO_1260 (O_1260,N_9979,N_9898);
xor UO_1261 (O_1261,N_9916,N_9933);
and UO_1262 (O_1262,N_9945,N_9812);
or UO_1263 (O_1263,N_9881,N_9889);
nand UO_1264 (O_1264,N_9990,N_9846);
and UO_1265 (O_1265,N_9895,N_9971);
nor UO_1266 (O_1266,N_9853,N_9910);
nand UO_1267 (O_1267,N_9991,N_9906);
nand UO_1268 (O_1268,N_9820,N_9986);
nand UO_1269 (O_1269,N_9877,N_9872);
and UO_1270 (O_1270,N_9865,N_9988);
nand UO_1271 (O_1271,N_9805,N_9858);
nand UO_1272 (O_1272,N_9844,N_9833);
and UO_1273 (O_1273,N_9916,N_9882);
and UO_1274 (O_1274,N_9956,N_9988);
or UO_1275 (O_1275,N_9935,N_9825);
or UO_1276 (O_1276,N_9806,N_9879);
nor UO_1277 (O_1277,N_9929,N_9835);
or UO_1278 (O_1278,N_9877,N_9891);
nand UO_1279 (O_1279,N_9972,N_9906);
or UO_1280 (O_1280,N_9817,N_9841);
or UO_1281 (O_1281,N_9911,N_9836);
and UO_1282 (O_1282,N_9812,N_9957);
and UO_1283 (O_1283,N_9973,N_9931);
nor UO_1284 (O_1284,N_9935,N_9976);
nor UO_1285 (O_1285,N_9960,N_9916);
or UO_1286 (O_1286,N_9880,N_9837);
xnor UO_1287 (O_1287,N_9993,N_9976);
nand UO_1288 (O_1288,N_9970,N_9908);
and UO_1289 (O_1289,N_9965,N_9902);
nand UO_1290 (O_1290,N_9822,N_9981);
or UO_1291 (O_1291,N_9901,N_9990);
nor UO_1292 (O_1292,N_9852,N_9951);
or UO_1293 (O_1293,N_9966,N_9808);
xnor UO_1294 (O_1294,N_9994,N_9828);
xnor UO_1295 (O_1295,N_9855,N_9966);
and UO_1296 (O_1296,N_9834,N_9975);
nand UO_1297 (O_1297,N_9878,N_9943);
nand UO_1298 (O_1298,N_9828,N_9930);
nand UO_1299 (O_1299,N_9813,N_9869);
xor UO_1300 (O_1300,N_9908,N_9954);
nand UO_1301 (O_1301,N_9906,N_9988);
nor UO_1302 (O_1302,N_9982,N_9979);
nor UO_1303 (O_1303,N_9829,N_9914);
xor UO_1304 (O_1304,N_9893,N_9946);
nand UO_1305 (O_1305,N_9852,N_9978);
nand UO_1306 (O_1306,N_9967,N_9906);
nand UO_1307 (O_1307,N_9977,N_9882);
nand UO_1308 (O_1308,N_9841,N_9970);
and UO_1309 (O_1309,N_9877,N_9971);
or UO_1310 (O_1310,N_9822,N_9846);
xor UO_1311 (O_1311,N_9946,N_9939);
xor UO_1312 (O_1312,N_9968,N_9892);
or UO_1313 (O_1313,N_9966,N_9879);
nor UO_1314 (O_1314,N_9958,N_9844);
nor UO_1315 (O_1315,N_9896,N_9852);
or UO_1316 (O_1316,N_9990,N_9961);
or UO_1317 (O_1317,N_9847,N_9986);
nand UO_1318 (O_1318,N_9893,N_9810);
nor UO_1319 (O_1319,N_9867,N_9894);
nand UO_1320 (O_1320,N_9951,N_9908);
and UO_1321 (O_1321,N_9841,N_9908);
nand UO_1322 (O_1322,N_9968,N_9813);
or UO_1323 (O_1323,N_9918,N_9961);
and UO_1324 (O_1324,N_9986,N_9934);
nand UO_1325 (O_1325,N_9999,N_9898);
nor UO_1326 (O_1326,N_9808,N_9957);
nand UO_1327 (O_1327,N_9942,N_9893);
or UO_1328 (O_1328,N_9882,N_9853);
xnor UO_1329 (O_1329,N_9827,N_9932);
nand UO_1330 (O_1330,N_9954,N_9892);
and UO_1331 (O_1331,N_9878,N_9942);
xor UO_1332 (O_1332,N_9889,N_9969);
nand UO_1333 (O_1333,N_9854,N_9915);
nor UO_1334 (O_1334,N_9876,N_9845);
nor UO_1335 (O_1335,N_9946,N_9858);
and UO_1336 (O_1336,N_9893,N_9858);
and UO_1337 (O_1337,N_9854,N_9916);
nor UO_1338 (O_1338,N_9898,N_9959);
xnor UO_1339 (O_1339,N_9823,N_9837);
and UO_1340 (O_1340,N_9881,N_9898);
nand UO_1341 (O_1341,N_9965,N_9946);
or UO_1342 (O_1342,N_9890,N_9933);
or UO_1343 (O_1343,N_9933,N_9839);
and UO_1344 (O_1344,N_9994,N_9907);
or UO_1345 (O_1345,N_9889,N_9964);
xnor UO_1346 (O_1346,N_9936,N_9994);
nor UO_1347 (O_1347,N_9838,N_9844);
nand UO_1348 (O_1348,N_9902,N_9985);
and UO_1349 (O_1349,N_9960,N_9802);
nor UO_1350 (O_1350,N_9864,N_9863);
nor UO_1351 (O_1351,N_9803,N_9903);
nor UO_1352 (O_1352,N_9809,N_9994);
and UO_1353 (O_1353,N_9910,N_9934);
and UO_1354 (O_1354,N_9978,N_9873);
nand UO_1355 (O_1355,N_9977,N_9909);
nand UO_1356 (O_1356,N_9910,N_9955);
and UO_1357 (O_1357,N_9952,N_9935);
nand UO_1358 (O_1358,N_9869,N_9915);
nor UO_1359 (O_1359,N_9919,N_9905);
nor UO_1360 (O_1360,N_9939,N_9852);
or UO_1361 (O_1361,N_9805,N_9821);
xnor UO_1362 (O_1362,N_9956,N_9891);
nor UO_1363 (O_1363,N_9998,N_9847);
and UO_1364 (O_1364,N_9815,N_9800);
or UO_1365 (O_1365,N_9979,N_9860);
nand UO_1366 (O_1366,N_9891,N_9831);
xor UO_1367 (O_1367,N_9816,N_9916);
and UO_1368 (O_1368,N_9818,N_9921);
and UO_1369 (O_1369,N_9899,N_9969);
and UO_1370 (O_1370,N_9804,N_9965);
xor UO_1371 (O_1371,N_9844,N_9926);
and UO_1372 (O_1372,N_9860,N_9994);
and UO_1373 (O_1373,N_9810,N_9876);
nor UO_1374 (O_1374,N_9913,N_9911);
and UO_1375 (O_1375,N_9840,N_9827);
nor UO_1376 (O_1376,N_9941,N_9875);
or UO_1377 (O_1377,N_9853,N_9922);
nand UO_1378 (O_1378,N_9910,N_9857);
xor UO_1379 (O_1379,N_9934,N_9866);
xor UO_1380 (O_1380,N_9914,N_9929);
nor UO_1381 (O_1381,N_9900,N_9832);
or UO_1382 (O_1382,N_9912,N_9943);
nor UO_1383 (O_1383,N_9848,N_9878);
nor UO_1384 (O_1384,N_9978,N_9811);
or UO_1385 (O_1385,N_9899,N_9968);
nand UO_1386 (O_1386,N_9974,N_9803);
nand UO_1387 (O_1387,N_9878,N_9912);
or UO_1388 (O_1388,N_9865,N_9960);
and UO_1389 (O_1389,N_9927,N_9821);
nand UO_1390 (O_1390,N_9877,N_9934);
xnor UO_1391 (O_1391,N_9881,N_9836);
xnor UO_1392 (O_1392,N_9812,N_9910);
xnor UO_1393 (O_1393,N_9917,N_9805);
and UO_1394 (O_1394,N_9882,N_9883);
or UO_1395 (O_1395,N_9944,N_9905);
nand UO_1396 (O_1396,N_9931,N_9800);
nand UO_1397 (O_1397,N_9835,N_9907);
nor UO_1398 (O_1398,N_9908,N_9933);
xor UO_1399 (O_1399,N_9971,N_9972);
nor UO_1400 (O_1400,N_9984,N_9889);
xnor UO_1401 (O_1401,N_9829,N_9854);
or UO_1402 (O_1402,N_9800,N_9983);
and UO_1403 (O_1403,N_9809,N_9986);
or UO_1404 (O_1404,N_9856,N_9864);
nor UO_1405 (O_1405,N_9961,N_9943);
and UO_1406 (O_1406,N_9921,N_9907);
nand UO_1407 (O_1407,N_9897,N_9942);
nand UO_1408 (O_1408,N_9974,N_9983);
nand UO_1409 (O_1409,N_9963,N_9879);
nand UO_1410 (O_1410,N_9935,N_9859);
nand UO_1411 (O_1411,N_9977,N_9919);
nand UO_1412 (O_1412,N_9893,N_9829);
or UO_1413 (O_1413,N_9849,N_9904);
or UO_1414 (O_1414,N_9871,N_9819);
and UO_1415 (O_1415,N_9861,N_9879);
xor UO_1416 (O_1416,N_9912,N_9989);
or UO_1417 (O_1417,N_9926,N_9877);
and UO_1418 (O_1418,N_9938,N_9950);
xnor UO_1419 (O_1419,N_9850,N_9839);
nand UO_1420 (O_1420,N_9854,N_9977);
xnor UO_1421 (O_1421,N_9933,N_9907);
nor UO_1422 (O_1422,N_9828,N_9954);
or UO_1423 (O_1423,N_9850,N_9849);
and UO_1424 (O_1424,N_9892,N_9943);
and UO_1425 (O_1425,N_9860,N_9904);
nand UO_1426 (O_1426,N_9839,N_9995);
nor UO_1427 (O_1427,N_9980,N_9969);
and UO_1428 (O_1428,N_9952,N_9800);
nor UO_1429 (O_1429,N_9827,N_9910);
xnor UO_1430 (O_1430,N_9973,N_9887);
or UO_1431 (O_1431,N_9958,N_9940);
and UO_1432 (O_1432,N_9830,N_9960);
nand UO_1433 (O_1433,N_9838,N_9829);
xor UO_1434 (O_1434,N_9868,N_9928);
nor UO_1435 (O_1435,N_9943,N_9933);
and UO_1436 (O_1436,N_9885,N_9822);
xnor UO_1437 (O_1437,N_9901,N_9856);
and UO_1438 (O_1438,N_9846,N_9986);
xor UO_1439 (O_1439,N_9953,N_9870);
xnor UO_1440 (O_1440,N_9817,N_9918);
or UO_1441 (O_1441,N_9869,N_9822);
nor UO_1442 (O_1442,N_9951,N_9891);
nor UO_1443 (O_1443,N_9933,N_9809);
xor UO_1444 (O_1444,N_9892,N_9941);
nand UO_1445 (O_1445,N_9946,N_9921);
xnor UO_1446 (O_1446,N_9869,N_9901);
nor UO_1447 (O_1447,N_9813,N_9878);
or UO_1448 (O_1448,N_9960,N_9849);
or UO_1449 (O_1449,N_9962,N_9828);
and UO_1450 (O_1450,N_9831,N_9977);
xor UO_1451 (O_1451,N_9801,N_9955);
nand UO_1452 (O_1452,N_9945,N_9819);
or UO_1453 (O_1453,N_9832,N_9858);
xor UO_1454 (O_1454,N_9969,N_9973);
nand UO_1455 (O_1455,N_9839,N_9976);
nor UO_1456 (O_1456,N_9913,N_9977);
nand UO_1457 (O_1457,N_9985,N_9872);
or UO_1458 (O_1458,N_9889,N_9823);
xnor UO_1459 (O_1459,N_9963,N_9961);
nand UO_1460 (O_1460,N_9940,N_9847);
and UO_1461 (O_1461,N_9808,N_9886);
and UO_1462 (O_1462,N_9927,N_9822);
xor UO_1463 (O_1463,N_9927,N_9993);
xnor UO_1464 (O_1464,N_9936,N_9963);
xor UO_1465 (O_1465,N_9826,N_9836);
or UO_1466 (O_1466,N_9996,N_9866);
nand UO_1467 (O_1467,N_9816,N_9842);
nor UO_1468 (O_1468,N_9838,N_9998);
nor UO_1469 (O_1469,N_9920,N_9908);
nor UO_1470 (O_1470,N_9820,N_9972);
nand UO_1471 (O_1471,N_9816,N_9930);
nor UO_1472 (O_1472,N_9983,N_9926);
xor UO_1473 (O_1473,N_9914,N_9981);
nand UO_1474 (O_1474,N_9886,N_9992);
nor UO_1475 (O_1475,N_9994,N_9993);
or UO_1476 (O_1476,N_9937,N_9970);
and UO_1477 (O_1477,N_9962,N_9909);
nand UO_1478 (O_1478,N_9924,N_9817);
nor UO_1479 (O_1479,N_9877,N_9860);
and UO_1480 (O_1480,N_9801,N_9877);
nor UO_1481 (O_1481,N_9871,N_9872);
nand UO_1482 (O_1482,N_9865,N_9946);
and UO_1483 (O_1483,N_9857,N_9967);
and UO_1484 (O_1484,N_9857,N_9911);
or UO_1485 (O_1485,N_9867,N_9880);
nand UO_1486 (O_1486,N_9999,N_9844);
nor UO_1487 (O_1487,N_9842,N_9851);
nor UO_1488 (O_1488,N_9956,N_9912);
nor UO_1489 (O_1489,N_9937,N_9861);
or UO_1490 (O_1490,N_9899,N_9898);
or UO_1491 (O_1491,N_9891,N_9917);
nor UO_1492 (O_1492,N_9987,N_9992);
or UO_1493 (O_1493,N_9918,N_9920);
or UO_1494 (O_1494,N_9955,N_9869);
or UO_1495 (O_1495,N_9906,N_9856);
or UO_1496 (O_1496,N_9869,N_9997);
and UO_1497 (O_1497,N_9939,N_9913);
nand UO_1498 (O_1498,N_9811,N_9903);
nor UO_1499 (O_1499,N_9931,N_9897);
endmodule