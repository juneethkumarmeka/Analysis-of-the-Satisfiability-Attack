module basic_1500_15000_2000_100_levels_5xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nor U0 (N_0,In_743,In_521);
or U1 (N_1,In_876,In_62);
and U2 (N_2,In_657,In_52);
or U3 (N_3,In_1214,In_1318);
nand U4 (N_4,In_680,In_1361);
or U5 (N_5,In_1401,In_1362);
and U6 (N_6,In_385,In_764);
or U7 (N_7,In_503,In_854);
nand U8 (N_8,In_140,In_419);
xor U9 (N_9,In_287,In_1018);
xnor U10 (N_10,In_429,In_294);
nand U11 (N_11,In_1356,In_1269);
or U12 (N_12,In_967,In_1475);
nand U13 (N_13,In_247,In_783);
nand U14 (N_14,In_1164,In_72);
or U15 (N_15,In_1021,In_1186);
or U16 (N_16,In_964,In_1173);
or U17 (N_17,In_932,In_891);
nor U18 (N_18,In_953,In_453);
nand U19 (N_19,In_102,In_421);
nand U20 (N_20,In_499,In_966);
nand U21 (N_21,In_1313,In_674);
or U22 (N_22,In_1266,In_442);
nor U23 (N_23,In_1322,In_1245);
or U24 (N_24,In_726,In_1357);
and U25 (N_25,In_951,In_904);
and U26 (N_26,In_1092,In_469);
and U27 (N_27,In_661,In_666);
nor U28 (N_28,In_1123,In_1295);
nor U29 (N_29,In_1177,In_393);
xnor U30 (N_30,In_578,In_775);
nand U31 (N_31,In_769,In_56);
or U32 (N_32,In_173,In_166);
nand U33 (N_33,In_1010,In_980);
xor U34 (N_34,In_1126,In_88);
xnor U35 (N_35,In_472,In_747);
nor U36 (N_36,In_284,In_12);
or U37 (N_37,In_878,In_1335);
nand U38 (N_38,In_283,In_136);
nor U39 (N_39,In_383,In_1296);
and U40 (N_40,In_706,In_68);
and U41 (N_41,In_778,In_709);
and U42 (N_42,In_201,In_150);
nor U43 (N_43,In_780,In_896);
and U44 (N_44,In_466,In_1047);
or U45 (N_45,In_800,In_1168);
or U46 (N_46,In_722,In_330);
nand U47 (N_47,In_221,In_1455);
and U48 (N_48,In_853,In_464);
and U49 (N_49,In_347,In_683);
or U50 (N_50,In_1308,In_1);
and U51 (N_51,In_749,In_779);
and U52 (N_52,In_888,In_1145);
nor U53 (N_53,In_649,In_546);
and U54 (N_54,In_1138,In_757);
xnor U55 (N_55,In_881,In_282);
and U56 (N_56,In_887,In_1017);
nand U57 (N_57,In_1349,In_1074);
nor U58 (N_58,In_416,In_296);
nor U59 (N_59,In_720,In_1370);
and U60 (N_60,In_1206,In_101);
and U61 (N_61,In_149,In_627);
or U62 (N_62,In_1024,In_831);
or U63 (N_63,In_1449,In_804);
nand U64 (N_64,In_1107,In_653);
nand U65 (N_65,In_1013,In_332);
xor U66 (N_66,In_1140,In_885);
xnor U67 (N_67,In_1089,In_1417);
and U68 (N_68,In_1456,In_406);
and U69 (N_69,In_890,In_847);
nor U70 (N_70,In_353,In_801);
nor U71 (N_71,In_679,In_1108);
or U72 (N_72,In_1135,In_690);
xnor U73 (N_73,In_83,In_937);
nand U74 (N_74,In_1000,In_312);
nand U75 (N_75,In_174,In_835);
and U76 (N_76,In_130,In_281);
or U77 (N_77,In_197,In_672);
nor U78 (N_78,In_1427,In_467);
nand U79 (N_79,In_104,In_940);
nor U80 (N_80,In_1451,In_923);
xnor U81 (N_81,In_1376,In_868);
nor U82 (N_82,In_1262,In_1007);
or U83 (N_83,In_16,In_367);
nor U84 (N_84,In_1345,In_208);
and U85 (N_85,In_148,In_756);
nor U86 (N_86,In_1191,In_1154);
or U87 (N_87,In_376,In_298);
nor U88 (N_88,In_1174,In_1129);
and U89 (N_89,In_697,In_1254);
nor U90 (N_90,In_603,In_508);
or U91 (N_91,In_1205,In_1180);
and U92 (N_92,In_209,In_817);
xnor U93 (N_93,In_1088,In_850);
and U94 (N_94,In_46,In_1213);
xnor U95 (N_95,In_1044,In_1436);
nand U96 (N_96,In_326,In_109);
or U97 (N_97,In_211,In_218);
nand U98 (N_98,In_1187,In_788);
or U99 (N_99,In_699,In_658);
nor U100 (N_100,In_1265,In_580);
nor U101 (N_101,In_856,In_1453);
and U102 (N_102,In_321,In_1033);
nor U103 (N_103,In_1330,In_646);
nor U104 (N_104,In_1151,In_561);
and U105 (N_105,In_242,In_1182);
nor U106 (N_106,In_773,In_1144);
and U107 (N_107,In_115,In_436);
and U108 (N_108,In_1442,In_586);
nand U109 (N_109,In_1250,In_414);
nand U110 (N_110,In_1257,In_498);
and U111 (N_111,In_39,In_1172);
nor U112 (N_112,In_620,In_734);
nor U113 (N_113,In_23,In_1067);
nor U114 (N_114,In_316,In_3);
nor U115 (N_115,In_714,In_176);
nand U116 (N_116,In_1090,In_848);
nand U117 (N_117,In_1333,In_202);
or U118 (N_118,In_1227,In_1353);
xor U119 (N_119,In_269,In_231);
and U120 (N_120,In_1200,In_65);
nand U121 (N_121,In_698,In_403);
nand U122 (N_122,In_640,In_1190);
nand U123 (N_123,In_259,In_609);
nor U124 (N_124,In_573,In_771);
xnor U125 (N_125,In_270,In_628);
nand U126 (N_126,In_1378,In_372);
and U127 (N_127,In_359,In_1400);
or U128 (N_128,In_1328,In_205);
nand U129 (N_129,In_1368,In_1251);
nor U130 (N_130,In_420,In_217);
nor U131 (N_131,In_753,In_648);
or U132 (N_132,In_559,In_1188);
nor U133 (N_133,In_632,In_802);
nor U134 (N_134,In_76,In_1043);
and U135 (N_135,In_1408,In_1022);
and U136 (N_136,In_501,In_103);
or U137 (N_137,In_132,In_664);
or U138 (N_138,In_1252,In_688);
or U139 (N_139,In_1359,In_1127);
or U140 (N_140,In_568,In_796);
xor U141 (N_141,In_1087,In_1425);
nand U142 (N_142,In_789,In_1344);
and U143 (N_143,In_790,In_486);
or U144 (N_144,In_67,In_1136);
or U145 (N_145,In_1419,In_1426);
xnor U146 (N_146,In_551,In_234);
and U147 (N_147,In_1494,In_500);
nand U148 (N_148,In_1149,In_575);
or U149 (N_149,In_1041,In_765);
nand U150 (N_150,In_708,In_825);
nand U151 (N_151,In_4,In_1054);
nand U152 (N_152,In_970,In_671);
nand U153 (N_153,In_556,In_1342);
nor U154 (N_154,In_1462,N_99);
and U155 (N_155,In_812,In_643);
nand U156 (N_156,In_553,In_1255);
nand U157 (N_157,In_1194,In_1207);
nor U158 (N_158,In_867,In_922);
and U159 (N_159,In_363,In_1263);
nor U160 (N_160,In_668,In_273);
nor U161 (N_161,In_418,In_328);
xor U162 (N_162,In_502,N_133);
nand U163 (N_163,In_1066,In_1236);
nand U164 (N_164,In_1230,In_380);
or U165 (N_165,N_33,In_725);
nand U166 (N_166,In_879,In_96);
nor U167 (N_167,In_1304,In_261);
or U168 (N_168,In_331,In_1120);
xnor U169 (N_169,In_151,In_134);
or U170 (N_170,In_934,In_564);
and U171 (N_171,In_641,In_48);
or U172 (N_172,In_950,In_249);
nand U173 (N_173,In_1413,In_837);
nand U174 (N_174,In_1051,In_1146);
nand U175 (N_175,In_358,In_1373);
xnor U176 (N_176,In_1100,In_346);
xor U177 (N_177,In_1038,N_117);
nor U178 (N_178,In_991,In_244);
xnor U179 (N_179,In_1139,In_1472);
nand U180 (N_180,In_1468,In_523);
or U181 (N_181,In_689,In_718);
nand U182 (N_182,In_1485,In_1109);
or U183 (N_183,N_115,In_110);
nand U184 (N_184,In_514,In_100);
or U185 (N_185,In_29,In_184);
nor U186 (N_186,In_1256,In_577);
and U187 (N_187,In_1389,In_1032);
nand U188 (N_188,In_986,In_732);
and U189 (N_189,In_1477,In_260);
and U190 (N_190,In_836,In_622);
and U191 (N_191,In_144,In_105);
nor U192 (N_192,In_167,In_1011);
nand U193 (N_193,In_864,In_1244);
and U194 (N_194,In_624,In_996);
or U195 (N_195,In_1170,In_285);
xor U196 (N_196,In_869,In_1461);
or U197 (N_197,N_84,In_49);
nor U198 (N_198,In_735,N_102);
nand U199 (N_199,In_919,In_988);
and U200 (N_200,In_254,In_621);
or U201 (N_201,In_485,In_264);
xor U202 (N_202,In_567,In_159);
or U203 (N_203,In_785,In_1490);
xor U204 (N_204,In_112,In_1240);
xnor U205 (N_205,In_552,In_341);
nand U206 (N_206,In_345,In_871);
nor U207 (N_207,N_121,In_1082);
and U208 (N_208,In_895,In_659);
or U209 (N_209,In_713,In_1492);
and U210 (N_210,N_2,In_1476);
or U211 (N_211,In_400,In_1081);
or U212 (N_212,In_1185,In_163);
and U213 (N_213,In_894,N_147);
and U214 (N_214,N_32,In_536);
and U215 (N_215,In_118,In_1059);
nor U216 (N_216,In_228,In_252);
nor U217 (N_217,In_1445,In_379);
and U218 (N_218,In_517,In_1099);
or U219 (N_219,In_1212,In_1249);
nor U220 (N_220,N_52,In_458);
or U221 (N_221,In_1105,In_1029);
or U222 (N_222,N_111,N_127);
or U223 (N_223,N_69,N_83);
or U224 (N_224,In_288,In_731);
xor U225 (N_225,In_1235,In_815);
nor U226 (N_226,In_350,In_1034);
nand U227 (N_227,N_50,In_19);
and U228 (N_228,In_1294,In_484);
nand U229 (N_229,In_912,In_1379);
or U230 (N_230,In_447,In_87);
xor U231 (N_231,In_1117,In_1314);
nand U232 (N_232,In_647,N_38);
and U233 (N_233,In_1222,In_1438);
and U234 (N_234,In_576,N_73);
and U235 (N_235,N_48,In_560);
or U236 (N_236,In_1118,In_1480);
and U237 (N_237,In_1474,In_750);
nor U238 (N_238,In_129,In_926);
and U239 (N_239,In_843,In_1365);
or U240 (N_240,N_88,In_617);
or U241 (N_241,In_7,N_100);
and U242 (N_242,In_791,In_1452);
and U243 (N_243,In_160,N_80);
and U244 (N_244,In_89,In_444);
nor U245 (N_245,N_3,In_670);
or U246 (N_246,In_1458,In_510);
xor U247 (N_247,In_550,In_557);
and U248 (N_248,N_81,In_1454);
and U249 (N_249,In_1246,In_1479);
and U250 (N_250,In_687,In_207);
and U251 (N_251,In_98,N_27);
xnor U252 (N_252,N_65,N_4);
nor U253 (N_253,In_137,In_531);
xor U254 (N_254,In_369,In_248);
xor U255 (N_255,In_566,In_188);
nor U256 (N_256,In_1042,In_1299);
and U257 (N_257,N_47,In_995);
nor U258 (N_258,In_1096,In_1289);
and U259 (N_259,In_494,In_997);
nand U260 (N_260,In_973,In_535);
nand U261 (N_261,In_1157,In_862);
nand U262 (N_262,In_389,In_156);
or U263 (N_263,In_602,N_57);
nand U264 (N_264,In_475,In_682);
nor U265 (N_265,N_20,In_763);
and U266 (N_266,In_133,In_549);
nand U267 (N_267,In_968,In_607);
nand U268 (N_268,In_1460,In_117);
xnor U269 (N_269,In_183,In_1061);
nor U270 (N_270,In_318,In_1422);
and U271 (N_271,In_435,In_241);
nor U272 (N_272,In_366,In_53);
or U273 (N_273,In_827,In_1290);
nand U274 (N_274,In_972,In_1390);
or U275 (N_275,In_1130,In_1234);
nand U276 (N_276,In_1360,In_1152);
nor U277 (N_277,In_652,In_374);
or U278 (N_278,In_925,In_1469);
nor U279 (N_279,In_1473,In_761);
or U280 (N_280,In_776,In_373);
nand U281 (N_281,In_349,In_1448);
nor U282 (N_282,In_1424,In_784);
or U283 (N_283,In_1163,In_844);
and U284 (N_284,In_356,In_597);
or U285 (N_285,N_17,In_955);
or U286 (N_286,In_1093,In_64);
nand U287 (N_287,In_1094,In_1411);
or U288 (N_288,In_268,N_140);
or U289 (N_289,In_1006,In_439);
nor U290 (N_290,In_1482,In_1325);
or U291 (N_291,In_1332,In_518);
xor U292 (N_292,In_936,N_35);
or U293 (N_293,In_25,In_703);
nand U294 (N_294,In_1288,In_1125);
and U295 (N_295,N_16,In_1431);
nor U296 (N_296,In_198,In_942);
and U297 (N_297,N_7,In_1220);
nor U298 (N_298,N_122,In_604);
and U299 (N_299,In_277,In_711);
nand U300 (N_300,In_1057,N_139);
nor U301 (N_301,In_2,N_10);
and U302 (N_302,In_644,In_135);
and U303 (N_303,In_220,In_459);
or U304 (N_304,In_1056,In_94);
nand U305 (N_305,In_443,In_673);
nor U306 (N_306,N_152,In_1040);
xor U307 (N_307,N_55,In_548);
nand U308 (N_308,N_298,In_1119);
or U309 (N_309,In_1339,In_292);
nand U310 (N_310,In_1225,In_924);
or U311 (N_311,In_120,In_212);
or U312 (N_312,N_186,In_745);
and U313 (N_313,N_0,In_5);
nand U314 (N_314,In_766,In_1046);
or U315 (N_315,In_782,N_40);
nor U316 (N_316,In_61,In_478);
nand U317 (N_317,N_295,In_626);
or U318 (N_318,In_1440,N_285);
and U319 (N_319,In_1439,In_1496);
nand U320 (N_320,In_1278,In_1297);
nand U321 (N_321,In_900,In_194);
nor U322 (N_322,In_306,In_1277);
or U323 (N_323,In_1283,In_998);
xor U324 (N_324,In_1147,In_897);
nand U325 (N_325,N_184,N_199);
nand U326 (N_326,In_22,In_170);
or U327 (N_327,In_1323,In_266);
xnor U328 (N_328,In_147,In_1403);
nor U329 (N_329,In_1023,N_213);
and U330 (N_330,In_291,In_931);
nor U331 (N_331,In_1176,In_127);
nor U332 (N_332,In_267,N_231);
xor U333 (N_333,N_209,In_313);
nand U334 (N_334,In_781,In_1383);
or U335 (N_335,In_85,In_1048);
or U336 (N_336,N_204,In_615);
nand U337 (N_337,In_1459,In_816);
nand U338 (N_338,In_1050,In_477);
or U339 (N_339,In_655,In_10);
and U340 (N_340,N_205,N_86);
or U341 (N_341,N_246,N_120);
or U342 (N_342,In_1215,In_141);
or U343 (N_343,In_883,N_60);
and U344 (N_344,N_243,In_1415);
or U345 (N_345,In_841,N_141);
nand U346 (N_346,In_155,In_99);
and U347 (N_347,In_1124,N_206);
and U348 (N_348,In_901,N_62);
or U349 (N_349,In_606,N_31);
and U350 (N_350,In_920,In_855);
or U351 (N_351,In_397,In_872);
nor U352 (N_352,In_1301,In_1343);
and U353 (N_353,N_91,N_43);
and U354 (N_354,In_1003,In_44);
or U355 (N_355,In_333,In_344);
or U356 (N_356,In_335,In_1113);
xor U357 (N_357,In_537,N_39);
nand U358 (N_358,In_975,In_402);
nand U359 (N_359,N_167,In_1329);
and U360 (N_360,In_742,In_1259);
or U361 (N_361,In_128,In_235);
and U362 (N_362,In_834,In_365);
xnor U363 (N_363,In_272,In_424);
or U364 (N_364,N_106,In_941);
nand U365 (N_365,In_1060,N_242);
nand U366 (N_366,In_808,In_196);
nor U367 (N_367,In_905,In_90);
nand U368 (N_368,In_1310,In_1470);
nor U369 (N_369,N_168,In_907);
nor U370 (N_370,In_707,N_198);
or U371 (N_371,In_222,In_810);
nor U372 (N_372,N_128,In_1219);
nand U373 (N_373,In_210,In_1027);
or U374 (N_374,In_752,N_113);
and U375 (N_375,N_296,N_76);
nand U376 (N_376,In_1097,N_225);
and U377 (N_377,In_487,In_81);
or U378 (N_378,In_1084,N_175);
and U379 (N_379,N_176,In_987);
and U380 (N_380,In_465,N_241);
or U381 (N_381,In_431,N_182);
and U382 (N_382,In_343,In_55);
and U383 (N_383,In_600,In_1443);
and U384 (N_384,N_131,N_34);
nor U385 (N_385,In_86,In_172);
nand U386 (N_386,In_915,In_1467);
nand U387 (N_387,N_44,In_1291);
or U388 (N_388,In_84,In_1016);
and U389 (N_389,N_247,In_1364);
nor U390 (N_390,N_187,N_282);
nor U391 (N_391,In_73,In_1020);
or U392 (N_392,N_269,N_258);
or U393 (N_393,In_542,In_1354);
and U394 (N_394,In_9,In_1076);
nor U395 (N_395,In_1211,In_1327);
or U396 (N_396,N_66,In_1055);
nand U397 (N_397,In_1101,N_41);
and U398 (N_398,In_239,In_1111);
and U399 (N_399,N_159,In_114);
or U400 (N_400,In_719,N_260);
nor U401 (N_401,N_163,In_329);
nand U402 (N_402,N_179,N_275);
and U403 (N_403,In_1384,In_1104);
nand U404 (N_404,In_433,In_463);
and U405 (N_405,In_880,In_271);
or U406 (N_406,N_279,In_662);
nor U407 (N_407,In_645,In_1167);
and U408 (N_408,In_840,In_1495);
or U409 (N_409,In_608,In_911);
and U410 (N_410,N_264,In_1324);
or U411 (N_411,In_605,In_512);
or U412 (N_412,In_1128,In_390);
or U413 (N_413,N_137,In_1435);
nand U414 (N_414,In_432,In_1395);
and U415 (N_415,In_1183,N_263);
or U416 (N_416,In_663,In_651);
nor U417 (N_417,In_947,In_1068);
xnor U418 (N_418,In_1150,In_60);
nand U419 (N_419,In_164,N_70);
and U420 (N_420,In_1375,In_1447);
nand U421 (N_421,In_1137,In_434);
and U422 (N_422,In_59,In_1199);
nand U423 (N_423,In_741,In_1483);
xor U424 (N_424,In_1285,N_249);
nand U425 (N_425,In_301,In_587);
or U426 (N_426,In_38,In_1002);
or U427 (N_427,N_145,In_91);
nand U428 (N_428,In_1450,In_1209);
nand U429 (N_429,In_473,In_1337);
nand U430 (N_430,In_253,In_1039);
and U431 (N_431,In_8,N_112);
nor U432 (N_432,N_94,In_794);
xnor U433 (N_433,In_1171,In_1160);
xor U434 (N_434,In_863,In_152);
or U435 (N_435,In_1035,In_305);
xor U436 (N_436,In_1233,In_1487);
nand U437 (N_437,In_1280,In_943);
nand U438 (N_438,In_460,In_1189);
or U439 (N_439,In_496,In_770);
or U440 (N_440,In_1115,In_165);
or U441 (N_441,In_650,In_1303);
nand U442 (N_442,In_838,N_23);
and U443 (N_443,In_1274,N_172);
or U444 (N_444,N_107,In_807);
nand U445 (N_445,In_963,N_259);
nor U446 (N_446,N_236,N_132);
and U447 (N_447,In_178,In_866);
or U448 (N_448,In_1197,In_738);
nor U449 (N_449,In_540,In_952);
and U450 (N_450,In_143,In_162);
and U451 (N_451,N_381,N_437);
and U452 (N_452,N_90,In_612);
and U453 (N_453,In_1228,In_1005);
nand U454 (N_454,In_992,In_1428);
nand U455 (N_455,In_513,N_419);
nand U456 (N_456,In_1025,In_1009);
xor U457 (N_457,In_633,N_146);
and U458 (N_458,In_740,In_286);
nand U459 (N_459,In_1481,N_110);
nand U460 (N_460,N_347,In_492);
and U461 (N_461,In_192,In_596);
xnor U462 (N_462,In_14,N_191);
nor U463 (N_463,N_245,In_322);
nand U464 (N_464,In_497,In_851);
nor U465 (N_465,In_978,N_125);
nand U466 (N_466,N_5,In_569);
and U467 (N_467,N_166,In_1391);
and U468 (N_468,In_1366,In_910);
nand U469 (N_469,In_1272,In_594);
nor U470 (N_470,In_1471,In_1317);
or U471 (N_471,In_1078,N_373);
nor U472 (N_472,In_616,N_324);
nand U473 (N_473,N_216,In_956);
or U474 (N_474,N_331,N_287);
nor U475 (N_475,N_162,In_0);
nor U476 (N_476,In_462,In_693);
xnor U477 (N_477,In_495,N_330);
and U478 (N_478,In_1142,In_1374);
nand U479 (N_479,In_185,In_1224);
nand U480 (N_480,N_371,In_1371);
and U481 (N_481,In_727,In_859);
nor U482 (N_482,In_797,In_715);
or U483 (N_483,In_43,In_598);
and U484 (N_484,N_424,N_385);
nor U485 (N_485,In_1316,N_15);
nor U486 (N_486,In_425,In_1385);
nand U487 (N_487,In_723,In_13);
xor U488 (N_488,In_18,In_186);
or U489 (N_489,In_527,In_255);
nand U490 (N_490,In_1292,In_1457);
xor U491 (N_491,In_1004,In_1193);
nand U492 (N_492,In_1159,In_1261);
and U493 (N_493,In_793,N_395);
or U494 (N_494,N_273,In_232);
or U495 (N_495,In_32,In_528);
and U496 (N_496,N_157,N_443);
or U497 (N_497,In_69,N_297);
and U498 (N_498,In_928,In_696);
or U499 (N_499,In_1381,In_490);
xnor U500 (N_500,In_290,In_489);
nor U501 (N_501,N_332,N_194);
or U502 (N_502,In_33,In_455);
or U503 (N_503,N_343,N_440);
or U504 (N_504,In_507,In_11);
or U505 (N_505,In_1305,In_78);
and U506 (N_506,N_328,In_1407);
nor U507 (N_507,In_480,In_417);
and U508 (N_508,N_217,N_300);
and U509 (N_509,In_169,N_228);
nor U510 (N_510,In_977,In_565);
xnor U511 (N_511,In_42,In_1247);
nor U512 (N_512,In_1437,In_82);
nor U513 (N_513,N_290,In_229);
and U514 (N_514,N_447,N_292);
nor U515 (N_515,N_359,In_119);
xor U516 (N_516,In_562,In_906);
xor U517 (N_517,N_352,In_430);
or U518 (N_518,In_1367,N_9);
nand U519 (N_519,N_432,N_160);
and U520 (N_520,In_860,In_538);
and U521 (N_521,In_71,In_539);
nor U522 (N_522,N_302,In_1380);
or U523 (N_523,N_6,N_362);
nand U524 (N_524,N_267,N_394);
or U525 (N_525,N_377,In_334);
nor U526 (N_526,N_82,In_427);
nor U527 (N_527,In_1045,N_403);
or U528 (N_528,In_929,In_468);
and U529 (N_529,In_168,In_1393);
and U530 (N_530,In_1065,In_957);
nor U531 (N_531,In_17,N_315);
nand U532 (N_532,In_230,In_660);
nor U533 (N_533,In_476,N_402);
nor U534 (N_534,N_372,In_945);
or U535 (N_535,N_200,In_1114);
nor U536 (N_536,N_418,In_805);
nand U537 (N_537,In_1275,N_354);
and U538 (N_538,In_364,In_1484);
xor U539 (N_539,In_97,In_409);
and U540 (N_540,N_341,N_303);
nand U541 (N_541,N_234,N_349);
and U542 (N_542,N_374,In_310);
nor U543 (N_543,In_927,In_833);
nor U544 (N_544,In_407,In_1226);
nand U545 (N_545,In_767,N_215);
nor U546 (N_546,N_18,In_1031);
nor U547 (N_547,In_35,N_210);
or U548 (N_548,In_1208,In_522);
nor U549 (N_549,In_1198,N_433);
nor U550 (N_550,In_75,N_277);
xor U551 (N_551,In_1012,In_107);
nor U552 (N_552,In_351,N_64);
or U553 (N_553,In_451,In_438);
and U554 (N_554,N_138,In_1264);
and U555 (N_555,N_427,In_106);
xor U556 (N_556,N_316,In_1112);
nor U557 (N_557,In_1015,N_322);
and U558 (N_558,In_591,In_1169);
nor U559 (N_559,In_1077,In_257);
and U560 (N_560,In_180,In_909);
or U561 (N_561,In_839,In_200);
or U562 (N_562,In_1217,N_229);
nand U563 (N_563,In_30,N_158);
nor U564 (N_564,In_541,In_762);
or U565 (N_565,N_226,In_199);
nand U566 (N_566,N_12,N_161);
or U567 (N_567,In_579,N_196);
nand U568 (N_568,In_274,In_1306);
nand U569 (N_569,In_275,N_101);
nor U570 (N_570,N_75,N_29);
nand U571 (N_571,In_1410,N_108);
xnor U572 (N_572,N_299,In_1095);
nand U573 (N_573,In_470,In_471);
xnor U574 (N_574,In_792,N_365);
nand U575 (N_575,In_1086,In_108);
or U576 (N_576,In_171,N_250);
and U577 (N_577,In_1486,In_898);
nand U578 (N_578,In_935,In_593);
nand U579 (N_579,In_946,In_319);
nand U580 (N_580,In_307,In_563);
xor U581 (N_581,In_361,In_803);
or U582 (N_582,In_930,In_532);
nor U583 (N_583,N_239,In_362);
or U584 (N_584,In_758,In_70);
and U585 (N_585,N_380,N_388);
or U586 (N_586,In_40,In_819);
or U587 (N_587,In_694,In_1465);
nor U588 (N_588,N_291,N_181);
nor U589 (N_589,N_183,In_145);
xnor U590 (N_590,N_435,In_1062);
nand U591 (N_591,N_230,In_384);
nor U592 (N_592,In_822,In_293);
xor U593 (N_593,In_125,N_411);
or U594 (N_594,In_1196,N_237);
nand U595 (N_595,In_408,In_405);
nor U596 (N_596,In_34,In_1350);
nand U597 (N_597,In_618,N_136);
nand U598 (N_598,N_389,In_1229);
nor U599 (N_599,In_875,N_68);
nor U600 (N_600,N_547,N_221);
and U601 (N_601,In_122,In_74);
nor U602 (N_602,In_625,N_310);
or U603 (N_603,In_692,N_536);
nand U604 (N_604,N_407,N_335);
nand U605 (N_605,N_268,N_375);
nand U606 (N_606,N_207,N_189);
nor U607 (N_607,In_669,N_492);
nand U608 (N_608,N_114,N_558);
xnor U609 (N_609,In_423,In_1241);
nor U610 (N_610,N_289,N_565);
nor U611 (N_611,In_642,In_882);
or U612 (N_612,In_1153,N_567);
nor U613 (N_613,In_1239,N_382);
nand U614 (N_614,N_451,N_284);
and U615 (N_615,In_327,N_219);
and U616 (N_616,In_1499,In_1434);
and U617 (N_617,In_243,In_1334);
nor U618 (N_618,N_311,N_363);
and U619 (N_619,In_256,In_386);
nand U620 (N_620,In_760,In_1319);
or U621 (N_621,In_969,N_497);
xor U622 (N_622,In_1072,N_42);
or U623 (N_623,In_354,In_751);
nor U624 (N_624,In_382,In_404);
nand U625 (N_625,N_317,In_474);
and U626 (N_626,In_411,N_599);
and U627 (N_627,N_461,In_154);
nand U628 (N_628,N_553,In_1414);
nor U629 (N_629,N_591,N_423);
and U630 (N_630,In_238,In_504);
nor U631 (N_631,In_1070,In_983);
nand U632 (N_632,N_11,N_563);
and U633 (N_633,In_398,In_994);
or U634 (N_634,N_482,N_539);
xnor U635 (N_635,N_270,In_1053);
and U636 (N_636,In_1347,N_252);
and U637 (N_637,In_1348,N_178);
nor U638 (N_638,In_1260,In_481);
nand U639 (N_639,In_1276,N_401);
nor U640 (N_640,In_336,In_280);
and U641 (N_641,In_619,In_993);
or U642 (N_642,N_550,N_329);
nand U643 (N_643,N_484,N_489);
or U644 (N_644,N_448,In_739);
and U645 (N_645,In_811,N_306);
nand U646 (N_646,In_63,N_36);
or U647 (N_647,N_254,In_1273);
and U648 (N_648,In_1158,In_1079);
or U649 (N_649,N_473,In_1243);
or U650 (N_650,In_639,N_124);
nor U651 (N_651,N_544,In_1358);
nor U652 (N_652,In_1444,In_823);
and U653 (N_653,In_555,N_262);
or U654 (N_654,In_746,N_276);
xnor U655 (N_655,In_700,N_151);
and U656 (N_656,N_548,In_1210);
xnor U657 (N_657,In_37,N_513);
nor U658 (N_658,N_415,In_1201);
or U659 (N_659,In_355,N_323);
nor U660 (N_660,In_111,In_1133);
or U661 (N_661,N_422,N_579);
nor U662 (N_662,In_426,N_540);
nand U663 (N_663,In_729,N_528);
nor U664 (N_664,N_449,N_552);
nor U665 (N_665,In_954,In_873);
or U666 (N_666,In_158,In_1179);
xnor U667 (N_667,In_1464,N_595);
or U668 (N_668,In_636,N_201);
nor U669 (N_669,In_412,N_8);
xnor U670 (N_670,In_131,In_558);
nand U671 (N_671,N_171,In_748);
nand U672 (N_672,In_717,In_916);
or U673 (N_673,N_265,N_420);
or U674 (N_674,N_174,In_1204);
and U675 (N_675,N_467,In_638);
nor U676 (N_676,In_1184,N_63);
nand U677 (N_677,In_554,In_227);
or U678 (N_678,N_24,N_154);
and U679 (N_679,In_338,In_917);
and U680 (N_680,N_144,N_37);
or U681 (N_681,N_490,In_437);
nand U682 (N_682,N_462,N_592);
or U683 (N_683,In_695,N_436);
nand U684 (N_684,N_468,In_744);
or U685 (N_685,N_390,In_204);
nor U686 (N_686,In_299,In_153);
and U687 (N_687,N_118,N_193);
and U688 (N_688,N_488,In_572);
nand U689 (N_689,N_368,In_944);
and U690 (N_690,In_31,In_157);
or U691 (N_691,N_498,N_309);
nand U692 (N_692,In_889,N_379);
and U693 (N_693,N_572,In_1369);
nand U694 (N_694,N_77,N_214);
nor U695 (N_695,N_584,In_701);
nand U696 (N_696,N_529,In_315);
nand U697 (N_697,N_103,In_1143);
and U698 (N_698,In_918,In_214);
and U699 (N_699,N_405,In_1221);
or U700 (N_700,N_491,In_656);
nand U701 (N_701,In_1309,N_535);
or U702 (N_702,N_348,In_206);
nor U703 (N_703,In_1298,In_721);
nor U704 (N_704,In_445,In_939);
nor U705 (N_705,In_733,In_585);
nand U706 (N_706,In_824,N_190);
or U707 (N_707,In_516,N_526);
nand U708 (N_708,N_203,N_409);
or U709 (N_709,N_180,In_1058);
nand U710 (N_710,N_126,N_367);
or U711 (N_711,In_381,In_786);
nand U712 (N_712,In_1489,In_985);
nor U713 (N_713,In_1155,N_266);
nor U714 (N_714,In_399,In_1267);
and U715 (N_715,In_1141,N_165);
nor U716 (N_716,In_36,In_213);
nand U717 (N_717,N_472,N_487);
nand U718 (N_718,In_505,In_1271);
nand U719 (N_719,N_590,In_736);
nor U720 (N_720,N_514,In_378);
nand U721 (N_721,N_397,In_80);
and U722 (N_722,In_441,N_517);
and U723 (N_723,In_1331,In_1091);
nor U724 (N_724,N_286,In_422);
and U725 (N_725,In_415,In_547);
or U726 (N_726,N_408,N_294);
and U727 (N_727,In_1253,In_26);
or U728 (N_728,In_1203,N_51);
nand U729 (N_729,N_392,In_893);
or U730 (N_730,N_594,N_522);
nor U731 (N_731,N_557,In_236);
and U732 (N_732,In_892,In_686);
and U733 (N_733,N_28,N_134);
nor U734 (N_734,In_1232,In_601);
nand U735 (N_735,In_1463,N_314);
and U736 (N_736,N_393,In_308);
xor U737 (N_737,N_25,N_97);
or U738 (N_738,In_339,N_465);
nand U739 (N_739,In_377,In_303);
nor U740 (N_740,N_197,In_325);
nor U741 (N_741,N_235,N_321);
or U742 (N_742,In_181,N_466);
and U743 (N_743,In_1433,In_1404);
nand U744 (N_744,N_391,In_195);
or U745 (N_745,In_1423,In_730);
nor U746 (N_746,In_66,N_356);
nand U747 (N_747,N_586,N_22);
and U748 (N_748,In_126,N_504);
nor U749 (N_749,In_123,N_326);
and U750 (N_750,In_1302,N_633);
and U751 (N_751,N_412,N_571);
xor U752 (N_752,In_678,N_608);
or U753 (N_753,In_681,N_580);
and U754 (N_754,In_665,N_621);
nor U755 (N_755,In_1008,N_105);
nor U756 (N_756,N_361,In_614);
nor U757 (N_757,In_799,N_334);
and U758 (N_758,In_1181,In_121);
or U759 (N_759,N_610,N_566);
or U760 (N_760,N_494,N_747);
xor U761 (N_761,In_21,In_47);
nor U762 (N_762,In_676,In_187);
and U763 (N_763,N_554,In_352);
and U764 (N_764,In_410,N_720);
nor U765 (N_765,In_1387,N_177);
and U766 (N_766,N_96,N_616);
and U767 (N_767,In_58,N_631);
and U768 (N_768,N_512,In_534);
or U769 (N_769,N_202,N_278);
nand U770 (N_770,In_1355,N_446);
nor U771 (N_771,N_426,N_665);
and U772 (N_772,N_589,N_525);
xnor U773 (N_773,N_721,N_503);
nor U774 (N_774,N_684,In_388);
nor U775 (N_775,In_842,In_886);
nor U776 (N_776,N_675,In_832);
and U777 (N_777,N_305,N_453);
nand U778 (N_778,In_454,N_723);
or U779 (N_779,N_351,N_21);
and U780 (N_780,N_92,N_562);
and U781 (N_781,In_1340,In_1397);
or U782 (N_782,In_795,N_640);
xor U783 (N_783,N_486,N_342);
xor U784 (N_784,In_874,In_999);
or U785 (N_785,In_1311,In_1498);
nand U786 (N_786,In_1372,N_312);
and U787 (N_787,In_1409,In_483);
nand U788 (N_788,N_333,N_188);
or U789 (N_789,N_232,N_337);
nand U790 (N_790,N_716,In_1320);
nand U791 (N_791,In_337,N_516);
nand U792 (N_792,In_599,N_639);
and U793 (N_793,N_735,N_581);
nor U794 (N_794,In_54,In_138);
and U795 (N_795,In_1287,In_1493);
or U796 (N_796,N_744,N_450);
and U797 (N_797,In_1430,N_671);
nand U798 (N_798,N_685,In_759);
or U799 (N_799,N_135,N_95);
xor U800 (N_800,In_1216,In_1248);
nor U801 (N_801,N_169,In_401);
or U802 (N_802,In_396,N_588);
or U803 (N_803,N_666,In_1121);
or U804 (N_804,In_395,In_768);
nor U805 (N_805,In_984,In_716);
or U806 (N_806,N_561,N_731);
nand U807 (N_807,N_612,In_1218);
nor U808 (N_808,In_961,N_615);
or U809 (N_809,In_246,N_680);
nor U810 (N_810,In_821,N_664);
nor U811 (N_811,N_709,In_971);
or U812 (N_812,In_1069,N_656);
or U813 (N_813,N_509,N_726);
nand U814 (N_814,N_220,In_755);
xnor U815 (N_815,In_903,In_820);
or U816 (N_816,In_1175,In_798);
and U817 (N_817,N_474,N_620);
or U818 (N_818,N_143,In_311);
nand U819 (N_819,N_150,In_1382);
nand U820 (N_820,In_1402,In_1166);
nand U821 (N_821,In_529,N_281);
or U822 (N_822,N_72,N_541);
nor U823 (N_823,N_406,N_614);
and U824 (N_824,N_224,In_962);
nand U825 (N_825,N_734,In_1073);
xor U826 (N_826,N_698,In_479);
nor U827 (N_827,N_477,In_613);
nand U828 (N_828,N_123,N_736);
nor U829 (N_829,N_386,In_704);
and U830 (N_830,N_78,In_737);
or U831 (N_831,N_722,In_146);
nor U832 (N_832,In_846,N_71);
nand U833 (N_833,In_1284,N_549);
or U834 (N_834,N_304,N_223);
and U835 (N_835,In_520,N_650);
xor U836 (N_836,N_699,N_587);
nor U837 (N_837,N_543,N_670);
or U838 (N_838,N_538,N_520);
or U839 (N_839,In_829,In_1116);
nor U840 (N_840,N_510,In_899);
nor U841 (N_841,In_215,N_164);
or U842 (N_842,In_190,In_493);
nand U843 (N_843,In_1052,N_274);
nor U844 (N_844,In_877,In_818);
nand U845 (N_845,In_1085,In_193);
and U846 (N_846,N_398,In_1336);
nand U847 (N_847,In_225,N_149);
nand U848 (N_848,In_27,In_251);
and U849 (N_849,N_641,In_6);
and U850 (N_850,N_280,N_690);
and U851 (N_851,N_607,N_238);
and U852 (N_852,N_611,N_469);
nand U853 (N_853,In_324,In_45);
and U854 (N_854,N_674,In_809);
or U855 (N_855,In_958,In_428);
and U856 (N_856,N_49,N_609);
or U857 (N_857,In_724,N_527);
nor U858 (N_858,In_51,In_1075);
nor U859 (N_859,N_575,N_669);
or U860 (N_860,N_556,N_227);
or U861 (N_861,N_574,In_960);
xnor U862 (N_862,In_1441,N_626);
nor U863 (N_863,In_1037,In_348);
or U864 (N_864,In_685,N_702);
nor U865 (N_865,N_597,N_53);
nor U866 (N_866,In_279,N_643);
xor U867 (N_867,In_371,N_26);
nand U868 (N_868,In_921,In_340);
and U869 (N_869,In_113,In_849);
or U870 (N_870,N_678,N_628);
or U871 (N_871,In_634,N_459);
nand U872 (N_872,N_596,N_687);
nor U873 (N_873,In_691,N_648);
and U874 (N_874,In_884,N_658);
and U875 (N_875,N_30,In_223);
nand U876 (N_876,In_456,N_463);
and U877 (N_877,In_630,In_1326);
or U878 (N_878,In_448,N_619);
nand U879 (N_879,In_309,In_1049);
nand U880 (N_880,In_1019,N_248);
nor U881 (N_881,N_724,N_480);
and U882 (N_882,In_1281,In_77);
and U883 (N_883,In_828,In_574);
nand U884 (N_884,N_627,N_630);
nor U885 (N_885,In_1488,N_708);
nor U886 (N_886,In_1392,N_364);
and U887 (N_887,N_502,N_98);
or U888 (N_888,N_668,N_559);
nor U889 (N_889,N_142,N_695);
or U890 (N_890,N_104,In_511);
nand U891 (N_891,N_271,N_478);
nor U892 (N_892,In_570,In_1338);
or U893 (N_893,In_237,N_518);
nor U894 (N_894,In_304,In_440);
nor U895 (N_895,N_470,N_404);
or U896 (N_896,In_830,In_582);
nor U897 (N_897,In_584,In_654);
nor U898 (N_898,N_729,In_1478);
nor U899 (N_899,N_336,N_749);
nand U900 (N_900,N_500,N_679);
and U901 (N_901,N_773,N_256);
and U902 (N_902,N_681,N_795);
or U903 (N_903,N_456,In_583);
or U904 (N_904,N_764,N_807);
or U905 (N_905,N_383,N_645);
or U906 (N_906,In_482,N_399);
nor U907 (N_907,In_1399,In_1030);
nand U908 (N_908,N_318,In_1134);
nand U909 (N_909,In_265,In_1098);
nand U910 (N_910,N_706,N_842);
nand U911 (N_911,N_780,N_651);
nand U912 (N_912,N_109,In_1466);
nor U913 (N_913,N_776,In_667);
and U914 (N_914,In_588,N_476);
nor U915 (N_915,In_391,N_868);
xnor U916 (N_916,N_173,In_913);
or U917 (N_917,In_387,N_576);
and U918 (N_918,N_600,N_796);
and U919 (N_919,N_14,N_293);
or U920 (N_920,In_452,In_728);
nor U921 (N_921,N_93,N_786);
or U922 (N_922,N_434,N_784);
and U923 (N_923,In_631,In_857);
and U924 (N_924,N_717,N_551);
or U925 (N_925,In_675,N_703);
or U926 (N_926,N_378,N_659);
nand U927 (N_927,N_387,In_1351);
and U928 (N_928,N_624,N_755);
xor U929 (N_929,N_632,N_622);
nand U930 (N_930,N_761,In_1386);
nor U931 (N_931,N_346,N_417);
and U932 (N_932,N_806,N_787);
or U933 (N_933,N_560,In_865);
nor U934 (N_934,In_224,N_148);
and U935 (N_935,In_754,N_898);
and U936 (N_936,N_483,N_676);
and U937 (N_937,In_1238,In_1268);
nor U938 (N_938,N_818,In_509);
nor U939 (N_939,In_1282,In_488);
nor U940 (N_940,In_858,N_763);
nand U941 (N_941,N_775,N_153);
xor U942 (N_942,N_507,N_876);
and U943 (N_943,N_745,N_774);
xnor U944 (N_944,In_976,In_24);
nand U945 (N_945,N_211,N_766);
or U946 (N_946,N_710,In_590);
nor U947 (N_947,In_814,N_861);
or U948 (N_948,N_800,In_806);
nor U949 (N_949,N_886,In_1110);
and U950 (N_950,In_1300,N_694);
nand U951 (N_951,N_129,N_56);
nor U952 (N_952,N_689,N_801);
nand U953 (N_953,In_342,N_445);
nand U954 (N_954,In_289,In_491);
and U955 (N_955,N_825,N_441);
nor U956 (N_956,N_74,In_1398);
nand U957 (N_957,N_396,In_705);
and U958 (N_958,In_1279,N_212);
nor U959 (N_959,In_203,In_360);
or U960 (N_960,In_845,N_475);
or U961 (N_961,In_959,N_416);
and U962 (N_962,In_1237,In_1036);
nand U963 (N_963,N_244,In_93);
xor U964 (N_964,N_358,In_461);
and U965 (N_965,In_595,N_869);
nor U966 (N_966,N_357,N_578);
xnor U967 (N_967,N_485,In_1064);
nor U968 (N_968,N_251,In_1258);
or U969 (N_969,N_170,N_573);
and U970 (N_970,In_1102,N_704);
or U971 (N_971,N_852,N_524);
nor U972 (N_972,N_428,In_1148);
nor U973 (N_973,N_46,In_1132);
or U974 (N_974,N_442,In_1446);
nor U975 (N_975,In_317,N_888);
nand U976 (N_976,N_883,N_58);
nor U977 (N_977,N_431,N_570);
or U978 (N_978,In_870,N_771);
nand U979 (N_979,N_617,In_20);
or U980 (N_980,In_949,N_344);
and U981 (N_981,N_835,N_629);
and U982 (N_982,N_733,N_425);
and U983 (N_983,N_283,N_828);
xor U984 (N_984,In_1223,N_832);
nand U985 (N_985,N_682,N_863);
nor U986 (N_986,N_732,N_833);
nor U987 (N_987,In_1307,N_85);
nand U988 (N_988,In_179,N_634);
or U989 (N_989,N_452,N_683);
nand U990 (N_990,In_1028,In_50);
or U991 (N_991,In_15,N_877);
and U992 (N_992,In_1162,N_802);
nand U993 (N_993,In_948,N_255);
or U994 (N_994,In_1231,N_790);
nor U995 (N_995,N_301,N_779);
nand U996 (N_996,N_530,N_635);
nand U997 (N_997,N_192,N_455);
nor U998 (N_998,N_583,N_663);
nor U999 (N_999,N_421,N_677);
nand U1000 (N_1000,In_1156,N_499);
or U1001 (N_1001,N_569,N_233);
nor U1002 (N_1002,N_728,In_965);
and U1003 (N_1003,In_989,In_543);
xnor U1004 (N_1004,N_748,N_654);
nor U1005 (N_1005,N_743,N_815);
or U1006 (N_1006,N_534,N_384);
nand U1007 (N_1007,N_819,In_263);
or U1008 (N_1008,In_981,In_175);
xnor U1009 (N_1009,N_531,N_444);
nand U1010 (N_1010,N_827,N_846);
and U1011 (N_1011,N_762,In_258);
or U1012 (N_1012,In_1405,N_156);
or U1013 (N_1013,N_785,N_638);
or U1014 (N_1014,N_899,N_889);
or U1015 (N_1015,N_691,N_759);
nor U1016 (N_1016,N_878,N_655);
or U1017 (N_1017,N_61,N_400);
and U1018 (N_1018,N_798,N_697);
xnor U1019 (N_1019,N_320,N_839);
nand U1020 (N_1020,N_606,In_526);
or U1021 (N_1021,In_592,N_841);
and U1022 (N_1022,N_692,N_519);
nor U1023 (N_1023,In_1131,N_873);
and U1024 (N_1024,N_884,In_506);
or U1025 (N_1025,In_116,In_1346);
or U1026 (N_1026,In_1396,N_521);
and U1027 (N_1027,In_1001,N_714);
and U1028 (N_1028,N_894,In_1106);
or U1029 (N_1029,N_185,N_804);
nand U1030 (N_1030,N_119,N_642);
nand U1031 (N_1031,N_660,In_297);
and U1032 (N_1032,N_811,N_816);
or U1033 (N_1033,N_783,N_19);
or U1034 (N_1034,N_662,N_657);
nor U1035 (N_1035,N_870,N_719);
nand U1036 (N_1036,N_338,In_233);
or U1037 (N_1037,In_1341,N_858);
nand U1038 (N_1038,N_871,N_546);
xnor U1039 (N_1039,N_765,N_67);
nor U1040 (N_1040,N_810,In_990);
and U1041 (N_1041,N_817,In_772);
and U1042 (N_1042,N_496,N_895);
and U1043 (N_1043,In_1026,N_715);
nand U1044 (N_1044,N_727,In_1321);
and U1045 (N_1045,N_848,N_822);
nor U1046 (N_1046,N_644,N_701);
nand U1047 (N_1047,In_278,N_360);
and U1048 (N_1048,N_872,N_647);
nand U1049 (N_1049,In_1242,N_797);
nor U1050 (N_1050,N_952,N_885);
nand U1051 (N_1051,In_1377,N_998);
and U1052 (N_1052,In_623,N_957);
nor U1053 (N_1053,N_340,N_753);
or U1054 (N_1054,N_844,In_710);
nand U1055 (N_1055,N_880,In_702);
or U1056 (N_1056,N_917,In_530);
xor U1057 (N_1057,N_950,N_881);
nor U1058 (N_1058,In_226,In_28);
nand U1059 (N_1059,N_1025,N_713);
xnor U1060 (N_1060,N_792,N_661);
nand U1061 (N_1061,In_1103,In_57);
nor U1062 (N_1062,N_904,N_954);
nor U1063 (N_1063,N_934,In_1192);
xor U1064 (N_1064,N_1026,N_637);
xnor U1065 (N_1065,N_931,N_533);
nand U1066 (N_1066,N_686,In_139);
nand U1067 (N_1067,N_457,N_376);
nand U1068 (N_1068,N_820,N_413);
or U1069 (N_1069,N_307,N_834);
nor U1070 (N_1070,In_1014,N_195);
nor U1071 (N_1071,N_922,N_946);
nand U1072 (N_1072,N_936,N_438);
nor U1073 (N_1073,N_602,N_410);
or U1074 (N_1074,N_454,N_926);
or U1075 (N_1075,In_375,N_439);
nand U1076 (N_1076,N_515,N_981);
and U1077 (N_1077,In_1432,N_1024);
nor U1078 (N_1078,N_996,N_837);
nand U1079 (N_1079,N_985,N_1035);
and U1080 (N_1080,N_741,N_577);
nand U1081 (N_1081,N_501,N_912);
nand U1082 (N_1082,N_59,In_394);
and U1083 (N_1083,N_782,N_896);
nand U1084 (N_1084,N_707,N_928);
and U1085 (N_1085,N_933,N_943);
and U1086 (N_1086,N_840,In_1293);
nand U1087 (N_1087,N_636,N_1000);
or U1088 (N_1088,N_938,In_124);
and U1089 (N_1089,N_969,In_449);
nor U1090 (N_1090,N_738,N_958);
nor U1091 (N_1091,N_979,N_1002);
xnor U1092 (N_1092,N_508,N_856);
or U1093 (N_1093,N_672,In_320);
and U1094 (N_1094,N_962,N_845);
or U1095 (N_1095,N_920,N_1027);
nor U1096 (N_1096,N_949,N_992);
nor U1097 (N_1097,N_1003,N_867);
nor U1098 (N_1098,N_471,N_812);
xnor U1099 (N_1099,N_924,N_1012);
xnor U1100 (N_1100,N_854,N_1031);
or U1101 (N_1101,N_940,N_625);
xor U1102 (N_1102,N_711,N_523);
nor U1103 (N_1103,N_582,N_1001);
or U1104 (N_1104,N_866,N_972);
or U1105 (N_1105,N_887,N_980);
nor U1106 (N_1106,N_652,N_1005);
nand U1107 (N_1107,N_313,N_350);
and U1108 (N_1108,N_921,N_853);
and U1109 (N_1109,N_930,N_1019);
and U1110 (N_1110,N_805,N_705);
or U1111 (N_1111,N_623,N_688);
or U1112 (N_1112,N_953,N_902);
and U1113 (N_1113,N_857,N_13);
nand U1114 (N_1114,In_813,N_1015);
and U1115 (N_1115,N_1009,N_730);
xor U1116 (N_1116,In_1122,N_564);
nor U1117 (N_1117,N_925,N_532);
or U1118 (N_1118,In_1394,N_585);
or U1119 (N_1119,N_754,N_944);
xor U1120 (N_1120,N_909,In_262);
xor U1121 (N_1121,N_222,N_988);
nand U1122 (N_1122,N_1033,N_1018);
and U1123 (N_1123,N_89,N_1032);
and U1124 (N_1124,N_948,N_725);
and U1125 (N_1125,In_1406,In_276);
and U1126 (N_1126,N_505,N_907);
and U1127 (N_1127,In_41,N_1048);
nand U1128 (N_1128,In_611,N_956);
nor U1129 (N_1129,In_852,N_667);
nand U1130 (N_1130,In_524,N_1043);
nor U1131 (N_1131,N_967,In_684);
nor U1132 (N_1132,N_777,In_1312);
and U1133 (N_1133,N_911,N_843);
nor U1134 (N_1134,N_1034,N_770);
nand U1135 (N_1135,N_814,N_272);
or U1136 (N_1136,In_908,N_568);
xnor U1137 (N_1137,In_525,N_966);
nand U1138 (N_1138,N_353,In_323);
and U1139 (N_1139,N_1008,N_369);
or U1140 (N_1140,In_519,N_1047);
xor U1141 (N_1141,N_808,N_208);
nand U1142 (N_1142,N_995,In_1421);
nand U1143 (N_1143,In_545,N_850);
or U1144 (N_1144,N_976,In_1497);
nand U1145 (N_1145,N_824,In_1202);
nor U1146 (N_1146,N_493,N_900);
nand U1147 (N_1147,N_891,N_1042);
nand U1148 (N_1148,In_1429,In_635);
nand U1149 (N_1149,In_777,N_851);
or U1150 (N_1150,In_933,N_829);
or U1151 (N_1151,N_693,N_430);
or U1152 (N_1152,N_1046,In_295);
nand U1153 (N_1153,N_989,In_1063);
and U1154 (N_1154,N_155,N_862);
nand U1155 (N_1155,In_182,N_860);
or U1156 (N_1156,N_937,In_1195);
and U1157 (N_1157,In_1363,In_974);
nand U1158 (N_1158,In_177,N_984);
and U1159 (N_1159,In_240,N_1010);
or U1160 (N_1160,N_1,In_245);
and U1161 (N_1161,N_506,N_945);
nor U1162 (N_1162,N_414,N_757);
and U1163 (N_1163,N_849,N_345);
nor U1164 (N_1164,N_673,N_756);
and U1165 (N_1165,N_879,N_601);
nand U1166 (N_1166,N_935,N_982);
nand U1167 (N_1167,In_314,N_54);
nor U1168 (N_1168,In_571,N_751);
or U1169 (N_1169,N_964,N_1045);
nor U1170 (N_1170,In_1315,N_997);
and U1171 (N_1171,In_300,N_990);
nand U1172 (N_1172,In_446,N_830);
nor U1173 (N_1173,N_1007,N_882);
or U1174 (N_1174,N_618,N_960);
or U1175 (N_1175,In_370,N_1023);
or U1176 (N_1176,N_865,N_768);
nor U1177 (N_1177,N_932,N_646);
xnor U1178 (N_1178,N_999,In_1071);
xnor U1179 (N_1179,N_905,In_189);
or U1180 (N_1180,N_604,N_823);
nand U1181 (N_1181,In_610,N_965);
nor U1182 (N_1182,In_92,In_581);
xnor U1183 (N_1183,In_302,N_951);
nand U1184 (N_1184,N_130,N_87);
nor U1185 (N_1185,N_803,N_893);
or U1186 (N_1186,N_460,N_1020);
nand U1187 (N_1187,N_1039,N_973);
nor U1188 (N_1188,N_355,N_1016);
or U1189 (N_1189,N_772,In_1420);
nor U1190 (N_1190,N_919,In_191);
or U1191 (N_1191,In_1083,In_712);
xnor U1192 (N_1192,In_1416,N_327);
nand U1193 (N_1193,N_511,N_901);
nor U1194 (N_1194,In_914,N_791);
xor U1195 (N_1195,N_993,N_45);
nor U1196 (N_1196,In_216,N_1011);
nor U1197 (N_1197,N_913,N_847);
and U1198 (N_1198,N_261,In_219);
nand U1199 (N_1199,N_739,N_696);
nor U1200 (N_1200,N_366,N_875);
nor U1201 (N_1201,In_357,N_1179);
nand U1202 (N_1202,In_637,N_1036);
or U1203 (N_1203,N_1104,N_859);
nand U1204 (N_1204,In_1352,N_1195);
and U1205 (N_1205,N_1068,N_1162);
nor U1206 (N_1206,In_861,N_1189);
or U1207 (N_1207,N_929,N_1148);
or U1208 (N_1208,N_1143,N_1102);
nand U1209 (N_1209,N_1071,N_370);
nand U1210 (N_1210,N_1052,N_781);
nand U1211 (N_1211,N_1166,In_392);
or U1212 (N_1212,N_1180,N_1076);
nor U1213 (N_1213,N_1028,N_240);
or U1214 (N_1214,N_481,N_1181);
nand U1215 (N_1215,N_923,N_742);
or U1216 (N_1216,N_325,N_1135);
and U1217 (N_1217,N_1191,N_1146);
and U1218 (N_1218,N_1099,N_1004);
or U1219 (N_1219,N_542,N_1139);
and U1220 (N_1220,N_939,N_1108);
or U1221 (N_1221,N_218,N_740);
or U1222 (N_1222,N_1066,N_752);
or U1223 (N_1223,N_963,N_603);
and U1224 (N_1224,In_79,N_1138);
and U1225 (N_1225,N_653,N_1137);
or U1226 (N_1226,N_1160,N_1176);
and U1227 (N_1227,N_1065,N_1058);
or U1228 (N_1228,N_1072,N_1140);
nand U1229 (N_1229,N_1167,N_918);
and U1230 (N_1230,N_1122,N_1119);
nor U1231 (N_1231,N_1163,N_1054);
nor U1232 (N_1232,N_1030,N_718);
and U1233 (N_1233,N_1165,N_864);
nor U1234 (N_1234,N_1013,N_1044);
nor U1235 (N_1235,N_1190,N_288);
and U1236 (N_1236,N_1116,N_1183);
or U1237 (N_1237,N_1129,N_737);
nand U1238 (N_1238,N_1182,N_1061);
and U1239 (N_1239,N_1117,N_1093);
nor U1240 (N_1240,N_1040,N_1062);
or U1241 (N_1241,N_789,N_1142);
nor U1242 (N_1242,N_1106,N_1115);
and U1243 (N_1243,N_1050,N_793);
xor U1244 (N_1244,In_1165,N_1098);
nand U1245 (N_1245,N_1006,N_1056);
nor U1246 (N_1246,N_1080,In_979);
nand U1247 (N_1247,N_339,N_1092);
nand U1248 (N_1248,N_1085,In_250);
or U1249 (N_1249,N_1114,N_1152);
nand U1250 (N_1250,N_836,N_545);
and U1251 (N_1251,N_941,N_1113);
nand U1252 (N_1252,In_457,N_1073);
or U1253 (N_1253,N_1055,N_1121);
or U1254 (N_1254,N_942,N_458);
nor U1255 (N_1255,N_1168,In_1178);
and U1256 (N_1256,N_1087,N_1170);
nor U1257 (N_1257,N_1083,N_914);
nand U1258 (N_1258,N_1090,N_1173);
and U1259 (N_1259,N_1118,N_1164);
nand U1260 (N_1260,N_947,N_1038);
and U1261 (N_1261,In_787,N_910);
nand U1262 (N_1262,N_1144,N_1123);
and U1263 (N_1263,N_794,N_1089);
nand U1264 (N_1264,N_1074,N_769);
or U1265 (N_1265,N_1174,N_788);
or U1266 (N_1266,In_533,N_1064);
and U1267 (N_1267,N_1125,N_1069);
nand U1268 (N_1268,N_977,N_955);
xnor U1269 (N_1269,N_903,N_1141);
nor U1270 (N_1270,N_1021,N_874);
or U1271 (N_1271,N_927,In_982);
or U1272 (N_1272,N_1091,N_1197);
nor U1273 (N_1273,N_1094,N_1156);
or U1274 (N_1274,N_712,N_1103);
nor U1275 (N_1275,N_1101,N_1126);
nor U1276 (N_1276,N_1084,N_1149);
or U1277 (N_1277,N_1133,N_1041);
and U1278 (N_1278,In_1270,N_308);
nand U1279 (N_1279,N_319,N_1014);
or U1280 (N_1280,N_1186,N_987);
nand U1281 (N_1281,N_1131,In_142);
xnor U1282 (N_1282,In_677,N_1081);
and U1283 (N_1283,N_1063,N_1086);
xnor U1284 (N_1284,N_968,N_1198);
or U1285 (N_1285,N_1109,In_450);
or U1286 (N_1286,N_1188,In_1491);
and U1287 (N_1287,N_1192,In_515);
nor U1288 (N_1288,N_464,N_897);
or U1289 (N_1289,N_1096,N_1107);
or U1290 (N_1290,In_1286,N_983);
and U1291 (N_1291,N_975,N_1151);
and U1292 (N_1292,N_906,N_1185);
or U1293 (N_1293,N_826,In_1418);
nor U1294 (N_1294,N_974,N_1057);
nor U1295 (N_1295,In_1388,N_1017);
nand U1296 (N_1296,N_750,N_1171);
nor U1297 (N_1297,In_1080,N_1078);
or U1298 (N_1298,N_778,In_368);
nand U1299 (N_1299,N_649,N_961);
and U1300 (N_1300,N_746,In_938);
nor U1301 (N_1301,N_79,N_1105);
nor U1302 (N_1302,N_1077,N_1124);
nor U1303 (N_1303,N_555,In_826);
and U1304 (N_1304,N_1029,N_890);
nand U1305 (N_1305,N_855,N_1155);
xor U1306 (N_1306,In_544,N_613);
or U1307 (N_1307,N_1169,N_971);
or U1308 (N_1308,N_1053,N_799);
nor U1309 (N_1309,N_1158,N_1095);
or U1310 (N_1310,N_479,N_813);
nor U1311 (N_1311,N_1134,N_986);
or U1312 (N_1312,N_1111,N_767);
or U1313 (N_1313,N_605,N_959);
or U1314 (N_1314,N_760,N_991);
nand U1315 (N_1315,N_593,N_1128);
xor U1316 (N_1316,N_1059,N_253);
nor U1317 (N_1317,N_1097,N_970);
and U1318 (N_1318,N_1196,N_1070);
or U1319 (N_1319,N_838,N_908);
or U1320 (N_1320,In_1412,N_978);
and U1321 (N_1321,In_774,N_1136);
nand U1322 (N_1322,In_589,N_598);
nor U1323 (N_1323,N_1145,N_1037);
nand U1324 (N_1324,In_161,N_1177);
nand U1325 (N_1325,N_1120,N_1199);
or U1326 (N_1326,N_1172,N_1079);
nor U1327 (N_1327,N_1154,N_821);
or U1328 (N_1328,N_1110,N_1147);
nand U1329 (N_1329,N_1130,N_1112);
nor U1330 (N_1330,N_1075,N_1194);
xor U1331 (N_1331,In_1161,N_1067);
nand U1332 (N_1332,N_1187,N_537);
and U1333 (N_1333,In_629,N_700);
nor U1334 (N_1334,N_1127,N_1193);
and U1335 (N_1335,N_915,N_495);
xnor U1336 (N_1336,N_1132,In_902);
nor U1337 (N_1337,N_1100,N_916);
or U1338 (N_1338,N_1184,N_1150);
xnor U1339 (N_1339,N_1088,N_1175);
xor U1340 (N_1340,N_1082,In_413);
nor U1341 (N_1341,N_257,N_1051);
and U1342 (N_1342,N_1159,N_758);
and U1343 (N_1343,N_809,N_1060);
or U1344 (N_1344,N_892,N_1022);
or U1345 (N_1345,N_116,N_831);
or U1346 (N_1346,In_95,N_429);
nor U1347 (N_1347,N_1161,N_1178);
nand U1348 (N_1348,N_994,N_1049);
or U1349 (N_1349,N_1157,N_1153);
nand U1350 (N_1350,N_1283,N_1338);
nand U1351 (N_1351,N_1343,N_1211);
or U1352 (N_1352,N_1323,N_1251);
xor U1353 (N_1353,N_1330,N_1302);
and U1354 (N_1354,N_1296,N_1337);
or U1355 (N_1355,N_1230,N_1280);
or U1356 (N_1356,N_1274,N_1348);
and U1357 (N_1357,N_1332,N_1317);
or U1358 (N_1358,N_1247,N_1218);
nand U1359 (N_1359,N_1267,N_1282);
and U1360 (N_1360,N_1324,N_1221);
or U1361 (N_1361,N_1266,N_1208);
nor U1362 (N_1362,N_1308,N_1312);
nand U1363 (N_1363,N_1292,N_1232);
xnor U1364 (N_1364,N_1273,N_1210);
nand U1365 (N_1365,N_1320,N_1314);
or U1366 (N_1366,N_1249,N_1303);
nor U1367 (N_1367,N_1297,N_1217);
and U1368 (N_1368,N_1268,N_1220);
and U1369 (N_1369,N_1206,N_1225);
or U1370 (N_1370,N_1200,N_1226);
nand U1371 (N_1371,N_1339,N_1284);
nor U1372 (N_1372,N_1287,N_1325);
nand U1373 (N_1373,N_1240,N_1311);
and U1374 (N_1374,N_1347,N_1349);
and U1375 (N_1375,N_1345,N_1275);
nor U1376 (N_1376,N_1258,N_1334);
nand U1377 (N_1377,N_1246,N_1300);
nand U1378 (N_1378,N_1279,N_1257);
and U1379 (N_1379,N_1335,N_1340);
nor U1380 (N_1380,N_1262,N_1252);
nand U1381 (N_1381,N_1305,N_1256);
or U1382 (N_1382,N_1322,N_1254);
or U1383 (N_1383,N_1212,N_1329);
nor U1384 (N_1384,N_1316,N_1239);
or U1385 (N_1385,N_1234,N_1313);
nor U1386 (N_1386,N_1259,N_1301);
nor U1387 (N_1387,N_1319,N_1253);
nor U1388 (N_1388,N_1318,N_1326);
nor U1389 (N_1389,N_1214,N_1299);
or U1390 (N_1390,N_1237,N_1242);
nand U1391 (N_1391,N_1204,N_1207);
or U1392 (N_1392,N_1269,N_1255);
xnor U1393 (N_1393,N_1346,N_1272);
and U1394 (N_1394,N_1294,N_1264);
nor U1395 (N_1395,N_1244,N_1304);
and U1396 (N_1396,N_1223,N_1222);
nor U1397 (N_1397,N_1298,N_1321);
or U1398 (N_1398,N_1243,N_1216);
or U1399 (N_1399,N_1209,N_1236);
and U1400 (N_1400,N_1270,N_1307);
nor U1401 (N_1401,N_1306,N_1290);
nor U1402 (N_1402,N_1228,N_1245);
nor U1403 (N_1403,N_1227,N_1202);
nand U1404 (N_1404,N_1213,N_1342);
or U1405 (N_1405,N_1344,N_1215);
nand U1406 (N_1406,N_1285,N_1263);
and U1407 (N_1407,N_1289,N_1241);
nand U1408 (N_1408,N_1315,N_1295);
and U1409 (N_1409,N_1231,N_1260);
nor U1410 (N_1410,N_1205,N_1278);
xor U1411 (N_1411,N_1201,N_1271);
nand U1412 (N_1412,N_1291,N_1276);
nor U1413 (N_1413,N_1250,N_1286);
and U1414 (N_1414,N_1265,N_1277);
or U1415 (N_1415,N_1261,N_1341);
and U1416 (N_1416,N_1331,N_1328);
nand U1417 (N_1417,N_1235,N_1229);
xnor U1418 (N_1418,N_1293,N_1333);
nand U1419 (N_1419,N_1336,N_1233);
nor U1420 (N_1420,N_1327,N_1219);
xnor U1421 (N_1421,N_1281,N_1238);
nor U1422 (N_1422,N_1288,N_1310);
or U1423 (N_1423,N_1203,N_1224);
and U1424 (N_1424,N_1248,N_1309);
or U1425 (N_1425,N_1223,N_1325);
nor U1426 (N_1426,N_1310,N_1248);
xnor U1427 (N_1427,N_1210,N_1308);
or U1428 (N_1428,N_1248,N_1244);
nor U1429 (N_1429,N_1347,N_1265);
and U1430 (N_1430,N_1336,N_1310);
nor U1431 (N_1431,N_1282,N_1266);
xor U1432 (N_1432,N_1339,N_1293);
xnor U1433 (N_1433,N_1240,N_1283);
nand U1434 (N_1434,N_1246,N_1264);
nor U1435 (N_1435,N_1268,N_1272);
xor U1436 (N_1436,N_1270,N_1300);
and U1437 (N_1437,N_1264,N_1289);
and U1438 (N_1438,N_1288,N_1325);
nand U1439 (N_1439,N_1328,N_1225);
nor U1440 (N_1440,N_1207,N_1235);
and U1441 (N_1441,N_1231,N_1253);
xnor U1442 (N_1442,N_1256,N_1334);
and U1443 (N_1443,N_1305,N_1316);
nand U1444 (N_1444,N_1203,N_1291);
or U1445 (N_1445,N_1309,N_1232);
and U1446 (N_1446,N_1341,N_1245);
nand U1447 (N_1447,N_1228,N_1316);
xnor U1448 (N_1448,N_1343,N_1262);
nand U1449 (N_1449,N_1332,N_1212);
nand U1450 (N_1450,N_1312,N_1331);
or U1451 (N_1451,N_1316,N_1331);
nand U1452 (N_1452,N_1329,N_1345);
or U1453 (N_1453,N_1235,N_1264);
and U1454 (N_1454,N_1248,N_1335);
nor U1455 (N_1455,N_1211,N_1253);
nand U1456 (N_1456,N_1250,N_1253);
xnor U1457 (N_1457,N_1274,N_1289);
or U1458 (N_1458,N_1297,N_1310);
and U1459 (N_1459,N_1297,N_1295);
or U1460 (N_1460,N_1326,N_1299);
and U1461 (N_1461,N_1279,N_1243);
or U1462 (N_1462,N_1319,N_1223);
xnor U1463 (N_1463,N_1346,N_1320);
nand U1464 (N_1464,N_1201,N_1266);
xor U1465 (N_1465,N_1223,N_1349);
and U1466 (N_1466,N_1305,N_1308);
and U1467 (N_1467,N_1324,N_1201);
nand U1468 (N_1468,N_1265,N_1250);
or U1469 (N_1469,N_1342,N_1239);
nand U1470 (N_1470,N_1348,N_1223);
nor U1471 (N_1471,N_1225,N_1271);
nand U1472 (N_1472,N_1222,N_1261);
and U1473 (N_1473,N_1236,N_1229);
and U1474 (N_1474,N_1217,N_1233);
nand U1475 (N_1475,N_1227,N_1327);
nand U1476 (N_1476,N_1292,N_1322);
and U1477 (N_1477,N_1276,N_1349);
nor U1478 (N_1478,N_1311,N_1343);
xor U1479 (N_1479,N_1268,N_1277);
nand U1480 (N_1480,N_1315,N_1259);
nor U1481 (N_1481,N_1222,N_1226);
nand U1482 (N_1482,N_1299,N_1247);
and U1483 (N_1483,N_1316,N_1282);
nand U1484 (N_1484,N_1250,N_1312);
nor U1485 (N_1485,N_1209,N_1278);
or U1486 (N_1486,N_1299,N_1349);
nand U1487 (N_1487,N_1272,N_1293);
nor U1488 (N_1488,N_1326,N_1256);
or U1489 (N_1489,N_1244,N_1208);
nor U1490 (N_1490,N_1279,N_1230);
and U1491 (N_1491,N_1324,N_1339);
or U1492 (N_1492,N_1327,N_1264);
or U1493 (N_1493,N_1285,N_1259);
or U1494 (N_1494,N_1315,N_1327);
nor U1495 (N_1495,N_1245,N_1312);
nor U1496 (N_1496,N_1306,N_1276);
nand U1497 (N_1497,N_1243,N_1319);
and U1498 (N_1498,N_1328,N_1263);
xor U1499 (N_1499,N_1275,N_1268);
or U1500 (N_1500,N_1353,N_1486);
or U1501 (N_1501,N_1405,N_1466);
and U1502 (N_1502,N_1433,N_1452);
nor U1503 (N_1503,N_1432,N_1465);
or U1504 (N_1504,N_1361,N_1412);
nor U1505 (N_1505,N_1386,N_1495);
and U1506 (N_1506,N_1396,N_1484);
or U1507 (N_1507,N_1477,N_1395);
or U1508 (N_1508,N_1382,N_1402);
nand U1509 (N_1509,N_1365,N_1446);
and U1510 (N_1510,N_1410,N_1483);
nand U1511 (N_1511,N_1419,N_1479);
or U1512 (N_1512,N_1444,N_1398);
xnor U1513 (N_1513,N_1371,N_1494);
and U1514 (N_1514,N_1490,N_1457);
nand U1515 (N_1515,N_1438,N_1380);
nor U1516 (N_1516,N_1439,N_1397);
or U1517 (N_1517,N_1389,N_1392);
and U1518 (N_1518,N_1497,N_1451);
and U1519 (N_1519,N_1403,N_1492);
nand U1520 (N_1520,N_1478,N_1453);
xnor U1521 (N_1521,N_1414,N_1373);
xnor U1522 (N_1522,N_1499,N_1454);
nand U1523 (N_1523,N_1370,N_1469);
or U1524 (N_1524,N_1377,N_1471);
nor U1525 (N_1525,N_1393,N_1426);
or U1526 (N_1526,N_1378,N_1442);
or U1527 (N_1527,N_1475,N_1434);
xor U1528 (N_1528,N_1359,N_1430);
nand U1529 (N_1529,N_1358,N_1464);
and U1530 (N_1530,N_1468,N_1421);
nand U1531 (N_1531,N_1493,N_1472);
and U1532 (N_1532,N_1379,N_1470);
or U1533 (N_1533,N_1456,N_1422);
or U1534 (N_1534,N_1424,N_1401);
nand U1535 (N_1535,N_1372,N_1394);
or U1536 (N_1536,N_1431,N_1498);
nor U1537 (N_1537,N_1409,N_1443);
nand U1538 (N_1538,N_1447,N_1404);
nand U1539 (N_1539,N_1399,N_1363);
nand U1540 (N_1540,N_1485,N_1351);
nor U1541 (N_1541,N_1460,N_1428);
and U1542 (N_1542,N_1435,N_1445);
nor U1543 (N_1543,N_1381,N_1437);
and U1544 (N_1544,N_1385,N_1436);
and U1545 (N_1545,N_1491,N_1376);
and U1546 (N_1546,N_1406,N_1391);
nand U1547 (N_1547,N_1407,N_1416);
nor U1548 (N_1548,N_1367,N_1476);
and U1549 (N_1549,N_1408,N_1368);
xnor U1550 (N_1550,N_1427,N_1496);
nor U1551 (N_1551,N_1458,N_1352);
or U1552 (N_1552,N_1388,N_1449);
or U1553 (N_1553,N_1417,N_1357);
or U1554 (N_1554,N_1450,N_1369);
nand U1555 (N_1555,N_1481,N_1425);
and U1556 (N_1556,N_1448,N_1441);
xor U1557 (N_1557,N_1423,N_1488);
nor U1558 (N_1558,N_1487,N_1354);
nand U1559 (N_1559,N_1366,N_1387);
or U1560 (N_1560,N_1411,N_1473);
or U1561 (N_1561,N_1415,N_1429);
nand U1562 (N_1562,N_1350,N_1420);
or U1563 (N_1563,N_1384,N_1440);
nand U1564 (N_1564,N_1360,N_1455);
and U1565 (N_1565,N_1474,N_1459);
or U1566 (N_1566,N_1482,N_1462);
and U1567 (N_1567,N_1413,N_1362);
nor U1568 (N_1568,N_1418,N_1489);
and U1569 (N_1569,N_1355,N_1356);
xnor U1570 (N_1570,N_1461,N_1374);
nand U1571 (N_1571,N_1480,N_1390);
and U1572 (N_1572,N_1400,N_1383);
nand U1573 (N_1573,N_1364,N_1463);
and U1574 (N_1574,N_1375,N_1467);
nand U1575 (N_1575,N_1408,N_1358);
nor U1576 (N_1576,N_1496,N_1443);
and U1577 (N_1577,N_1467,N_1452);
or U1578 (N_1578,N_1421,N_1448);
nand U1579 (N_1579,N_1406,N_1433);
nand U1580 (N_1580,N_1451,N_1362);
nand U1581 (N_1581,N_1446,N_1387);
or U1582 (N_1582,N_1453,N_1473);
and U1583 (N_1583,N_1358,N_1352);
nor U1584 (N_1584,N_1409,N_1370);
nand U1585 (N_1585,N_1358,N_1486);
or U1586 (N_1586,N_1497,N_1429);
or U1587 (N_1587,N_1437,N_1492);
nand U1588 (N_1588,N_1384,N_1419);
nor U1589 (N_1589,N_1497,N_1404);
xnor U1590 (N_1590,N_1416,N_1399);
and U1591 (N_1591,N_1398,N_1408);
or U1592 (N_1592,N_1381,N_1435);
and U1593 (N_1593,N_1490,N_1439);
nand U1594 (N_1594,N_1361,N_1374);
and U1595 (N_1595,N_1458,N_1478);
or U1596 (N_1596,N_1443,N_1441);
or U1597 (N_1597,N_1411,N_1420);
and U1598 (N_1598,N_1482,N_1479);
and U1599 (N_1599,N_1450,N_1396);
nor U1600 (N_1600,N_1461,N_1455);
or U1601 (N_1601,N_1359,N_1355);
and U1602 (N_1602,N_1456,N_1406);
or U1603 (N_1603,N_1485,N_1458);
and U1604 (N_1604,N_1490,N_1418);
or U1605 (N_1605,N_1361,N_1435);
or U1606 (N_1606,N_1423,N_1416);
nand U1607 (N_1607,N_1393,N_1403);
or U1608 (N_1608,N_1427,N_1389);
nand U1609 (N_1609,N_1456,N_1452);
and U1610 (N_1610,N_1430,N_1389);
and U1611 (N_1611,N_1379,N_1444);
nor U1612 (N_1612,N_1382,N_1488);
or U1613 (N_1613,N_1463,N_1397);
nand U1614 (N_1614,N_1390,N_1384);
nand U1615 (N_1615,N_1451,N_1454);
nor U1616 (N_1616,N_1495,N_1494);
nor U1617 (N_1617,N_1486,N_1455);
nand U1618 (N_1618,N_1476,N_1412);
nor U1619 (N_1619,N_1395,N_1405);
and U1620 (N_1620,N_1370,N_1435);
or U1621 (N_1621,N_1402,N_1388);
xnor U1622 (N_1622,N_1475,N_1497);
and U1623 (N_1623,N_1451,N_1495);
and U1624 (N_1624,N_1456,N_1421);
and U1625 (N_1625,N_1424,N_1421);
or U1626 (N_1626,N_1362,N_1393);
nor U1627 (N_1627,N_1441,N_1425);
nor U1628 (N_1628,N_1491,N_1461);
nor U1629 (N_1629,N_1414,N_1449);
nor U1630 (N_1630,N_1463,N_1438);
xnor U1631 (N_1631,N_1408,N_1350);
or U1632 (N_1632,N_1475,N_1468);
and U1633 (N_1633,N_1371,N_1409);
xor U1634 (N_1634,N_1386,N_1477);
nor U1635 (N_1635,N_1359,N_1399);
xor U1636 (N_1636,N_1356,N_1485);
and U1637 (N_1637,N_1473,N_1360);
nor U1638 (N_1638,N_1403,N_1396);
xor U1639 (N_1639,N_1499,N_1398);
and U1640 (N_1640,N_1413,N_1442);
xor U1641 (N_1641,N_1465,N_1488);
xnor U1642 (N_1642,N_1375,N_1358);
and U1643 (N_1643,N_1409,N_1430);
and U1644 (N_1644,N_1387,N_1423);
and U1645 (N_1645,N_1421,N_1455);
and U1646 (N_1646,N_1453,N_1376);
or U1647 (N_1647,N_1366,N_1483);
and U1648 (N_1648,N_1437,N_1404);
xnor U1649 (N_1649,N_1471,N_1459);
or U1650 (N_1650,N_1533,N_1575);
and U1651 (N_1651,N_1553,N_1615);
or U1652 (N_1652,N_1585,N_1521);
nand U1653 (N_1653,N_1621,N_1646);
nand U1654 (N_1654,N_1578,N_1562);
nor U1655 (N_1655,N_1563,N_1513);
or U1656 (N_1656,N_1571,N_1532);
and U1657 (N_1657,N_1576,N_1580);
or U1658 (N_1658,N_1544,N_1638);
or U1659 (N_1659,N_1589,N_1614);
or U1660 (N_1660,N_1510,N_1545);
xor U1661 (N_1661,N_1500,N_1611);
and U1662 (N_1662,N_1600,N_1535);
nor U1663 (N_1663,N_1503,N_1507);
and U1664 (N_1664,N_1523,N_1622);
nor U1665 (N_1665,N_1573,N_1601);
nand U1666 (N_1666,N_1514,N_1531);
nand U1667 (N_1667,N_1527,N_1548);
nor U1668 (N_1668,N_1570,N_1592);
nor U1669 (N_1669,N_1616,N_1577);
and U1670 (N_1670,N_1591,N_1643);
nand U1671 (N_1671,N_1529,N_1590);
nor U1672 (N_1672,N_1582,N_1517);
xor U1673 (N_1673,N_1624,N_1550);
nor U1674 (N_1674,N_1647,N_1557);
nor U1675 (N_1675,N_1645,N_1649);
xnor U1676 (N_1676,N_1520,N_1603);
and U1677 (N_1677,N_1609,N_1560);
and U1678 (N_1678,N_1596,N_1509);
xnor U1679 (N_1679,N_1594,N_1623);
xnor U1680 (N_1680,N_1620,N_1551);
xnor U1681 (N_1681,N_1519,N_1628);
or U1682 (N_1682,N_1642,N_1542);
and U1683 (N_1683,N_1584,N_1602);
and U1684 (N_1684,N_1512,N_1636);
nor U1685 (N_1685,N_1581,N_1648);
or U1686 (N_1686,N_1511,N_1608);
nor U1687 (N_1687,N_1554,N_1605);
and U1688 (N_1688,N_1518,N_1536);
or U1689 (N_1689,N_1565,N_1644);
or U1690 (N_1690,N_1552,N_1639);
nor U1691 (N_1691,N_1569,N_1549);
and U1692 (N_1692,N_1593,N_1528);
nand U1693 (N_1693,N_1606,N_1618);
or U1694 (N_1694,N_1502,N_1556);
and U1695 (N_1695,N_1564,N_1522);
nor U1696 (N_1696,N_1588,N_1540);
nor U1697 (N_1697,N_1561,N_1579);
or U1698 (N_1698,N_1567,N_1506);
nor U1699 (N_1699,N_1516,N_1629);
nor U1700 (N_1700,N_1526,N_1558);
xnor U1701 (N_1701,N_1515,N_1604);
nor U1702 (N_1702,N_1612,N_1597);
nor U1703 (N_1703,N_1599,N_1534);
nor U1704 (N_1704,N_1587,N_1505);
nand U1705 (N_1705,N_1555,N_1640);
and U1706 (N_1706,N_1619,N_1627);
nand U1707 (N_1707,N_1617,N_1607);
or U1708 (N_1708,N_1610,N_1574);
nor U1709 (N_1709,N_1625,N_1632);
or U1710 (N_1710,N_1631,N_1630);
and U1711 (N_1711,N_1635,N_1537);
or U1712 (N_1712,N_1501,N_1566);
and U1713 (N_1713,N_1586,N_1539);
nand U1714 (N_1714,N_1525,N_1572);
or U1715 (N_1715,N_1508,N_1541);
and U1716 (N_1716,N_1530,N_1626);
and U1717 (N_1717,N_1546,N_1568);
nand U1718 (N_1718,N_1524,N_1641);
xnor U1719 (N_1719,N_1637,N_1547);
nand U1720 (N_1720,N_1633,N_1634);
and U1721 (N_1721,N_1595,N_1598);
nor U1722 (N_1722,N_1538,N_1504);
and U1723 (N_1723,N_1613,N_1559);
nand U1724 (N_1724,N_1583,N_1543);
nand U1725 (N_1725,N_1534,N_1648);
or U1726 (N_1726,N_1586,N_1584);
xor U1727 (N_1727,N_1527,N_1576);
nand U1728 (N_1728,N_1513,N_1510);
or U1729 (N_1729,N_1597,N_1574);
or U1730 (N_1730,N_1584,N_1547);
or U1731 (N_1731,N_1509,N_1612);
nand U1732 (N_1732,N_1500,N_1608);
and U1733 (N_1733,N_1566,N_1633);
and U1734 (N_1734,N_1588,N_1574);
or U1735 (N_1735,N_1606,N_1631);
nand U1736 (N_1736,N_1592,N_1617);
nor U1737 (N_1737,N_1518,N_1602);
nand U1738 (N_1738,N_1516,N_1564);
and U1739 (N_1739,N_1538,N_1516);
and U1740 (N_1740,N_1601,N_1626);
xnor U1741 (N_1741,N_1512,N_1612);
and U1742 (N_1742,N_1629,N_1551);
nor U1743 (N_1743,N_1596,N_1558);
and U1744 (N_1744,N_1555,N_1506);
and U1745 (N_1745,N_1616,N_1606);
nor U1746 (N_1746,N_1644,N_1541);
or U1747 (N_1747,N_1607,N_1586);
and U1748 (N_1748,N_1537,N_1642);
nor U1749 (N_1749,N_1620,N_1642);
and U1750 (N_1750,N_1603,N_1565);
nand U1751 (N_1751,N_1642,N_1611);
nand U1752 (N_1752,N_1622,N_1571);
nand U1753 (N_1753,N_1536,N_1508);
nand U1754 (N_1754,N_1527,N_1512);
nor U1755 (N_1755,N_1512,N_1611);
xor U1756 (N_1756,N_1549,N_1591);
and U1757 (N_1757,N_1640,N_1641);
nor U1758 (N_1758,N_1565,N_1619);
nand U1759 (N_1759,N_1576,N_1629);
or U1760 (N_1760,N_1510,N_1570);
nor U1761 (N_1761,N_1617,N_1568);
or U1762 (N_1762,N_1638,N_1581);
xnor U1763 (N_1763,N_1510,N_1532);
nand U1764 (N_1764,N_1560,N_1638);
nor U1765 (N_1765,N_1570,N_1551);
or U1766 (N_1766,N_1554,N_1557);
nor U1767 (N_1767,N_1567,N_1517);
xnor U1768 (N_1768,N_1622,N_1588);
and U1769 (N_1769,N_1501,N_1596);
xor U1770 (N_1770,N_1536,N_1530);
or U1771 (N_1771,N_1527,N_1595);
or U1772 (N_1772,N_1510,N_1500);
and U1773 (N_1773,N_1548,N_1618);
and U1774 (N_1774,N_1576,N_1604);
and U1775 (N_1775,N_1520,N_1518);
nand U1776 (N_1776,N_1595,N_1554);
and U1777 (N_1777,N_1635,N_1541);
nor U1778 (N_1778,N_1571,N_1646);
and U1779 (N_1779,N_1642,N_1505);
and U1780 (N_1780,N_1612,N_1555);
nand U1781 (N_1781,N_1500,N_1555);
or U1782 (N_1782,N_1523,N_1518);
nand U1783 (N_1783,N_1646,N_1565);
and U1784 (N_1784,N_1505,N_1533);
nor U1785 (N_1785,N_1531,N_1630);
nand U1786 (N_1786,N_1536,N_1550);
nor U1787 (N_1787,N_1604,N_1582);
nor U1788 (N_1788,N_1638,N_1636);
or U1789 (N_1789,N_1516,N_1643);
xor U1790 (N_1790,N_1546,N_1553);
or U1791 (N_1791,N_1555,N_1619);
and U1792 (N_1792,N_1614,N_1543);
xor U1793 (N_1793,N_1626,N_1522);
and U1794 (N_1794,N_1532,N_1528);
and U1795 (N_1795,N_1505,N_1544);
nand U1796 (N_1796,N_1573,N_1643);
xor U1797 (N_1797,N_1621,N_1600);
nor U1798 (N_1798,N_1626,N_1553);
or U1799 (N_1799,N_1645,N_1504);
nand U1800 (N_1800,N_1790,N_1770);
or U1801 (N_1801,N_1666,N_1748);
nor U1802 (N_1802,N_1654,N_1676);
nor U1803 (N_1803,N_1672,N_1723);
nand U1804 (N_1804,N_1677,N_1711);
or U1805 (N_1805,N_1709,N_1678);
and U1806 (N_1806,N_1651,N_1701);
or U1807 (N_1807,N_1784,N_1653);
xor U1808 (N_1808,N_1766,N_1732);
or U1809 (N_1809,N_1716,N_1727);
nand U1810 (N_1810,N_1776,N_1684);
nor U1811 (N_1811,N_1661,N_1664);
nor U1812 (N_1812,N_1745,N_1688);
or U1813 (N_1813,N_1662,N_1760);
or U1814 (N_1814,N_1699,N_1793);
xor U1815 (N_1815,N_1756,N_1740);
nor U1816 (N_1816,N_1722,N_1799);
nand U1817 (N_1817,N_1791,N_1786);
nor U1818 (N_1818,N_1752,N_1663);
xor U1819 (N_1819,N_1702,N_1704);
or U1820 (N_1820,N_1725,N_1751);
and U1821 (N_1821,N_1767,N_1665);
and U1822 (N_1822,N_1796,N_1650);
or U1823 (N_1823,N_1734,N_1771);
xnor U1824 (N_1824,N_1658,N_1785);
and U1825 (N_1825,N_1772,N_1675);
nand U1826 (N_1826,N_1765,N_1724);
or U1827 (N_1827,N_1679,N_1660);
nand U1828 (N_1828,N_1690,N_1763);
and U1829 (N_1829,N_1652,N_1680);
xor U1830 (N_1830,N_1782,N_1657);
or U1831 (N_1831,N_1753,N_1671);
and U1832 (N_1832,N_1698,N_1747);
nor U1833 (N_1833,N_1700,N_1741);
nor U1834 (N_1834,N_1674,N_1774);
xnor U1835 (N_1835,N_1707,N_1768);
or U1836 (N_1836,N_1778,N_1797);
and U1837 (N_1837,N_1746,N_1764);
xnor U1838 (N_1838,N_1757,N_1750);
nor U1839 (N_1839,N_1773,N_1742);
nor U1840 (N_1840,N_1758,N_1695);
or U1841 (N_1841,N_1736,N_1726);
and U1842 (N_1842,N_1743,N_1744);
nand U1843 (N_1843,N_1681,N_1720);
nor U1844 (N_1844,N_1769,N_1731);
or U1845 (N_1845,N_1655,N_1728);
xor U1846 (N_1846,N_1656,N_1794);
or U1847 (N_1847,N_1761,N_1669);
nand U1848 (N_1848,N_1738,N_1682);
xor U1849 (N_1849,N_1670,N_1789);
or U1850 (N_1850,N_1715,N_1783);
nor U1851 (N_1851,N_1696,N_1667);
nand U1852 (N_1852,N_1710,N_1692);
nand U1853 (N_1853,N_1693,N_1755);
and U1854 (N_1854,N_1714,N_1686);
nand U1855 (N_1855,N_1735,N_1729);
and U1856 (N_1856,N_1718,N_1779);
and U1857 (N_1857,N_1717,N_1798);
or U1858 (N_1858,N_1687,N_1759);
and U1859 (N_1859,N_1705,N_1713);
xor U1860 (N_1860,N_1703,N_1788);
nand U1861 (N_1861,N_1712,N_1780);
and U1862 (N_1862,N_1787,N_1683);
nand U1863 (N_1863,N_1708,N_1721);
nor U1864 (N_1864,N_1792,N_1781);
and U1865 (N_1865,N_1775,N_1685);
or U1866 (N_1866,N_1697,N_1739);
and U1867 (N_1867,N_1673,N_1694);
nand U1868 (N_1868,N_1795,N_1749);
and U1869 (N_1869,N_1706,N_1719);
and U1870 (N_1870,N_1668,N_1754);
and U1871 (N_1871,N_1733,N_1762);
and U1872 (N_1872,N_1689,N_1777);
and U1873 (N_1873,N_1730,N_1659);
nand U1874 (N_1874,N_1737,N_1691);
and U1875 (N_1875,N_1653,N_1765);
nand U1876 (N_1876,N_1737,N_1762);
and U1877 (N_1877,N_1729,N_1650);
or U1878 (N_1878,N_1690,N_1746);
or U1879 (N_1879,N_1698,N_1756);
xnor U1880 (N_1880,N_1651,N_1655);
nor U1881 (N_1881,N_1695,N_1748);
xnor U1882 (N_1882,N_1777,N_1725);
nand U1883 (N_1883,N_1679,N_1739);
and U1884 (N_1884,N_1782,N_1734);
nor U1885 (N_1885,N_1725,N_1664);
xor U1886 (N_1886,N_1660,N_1667);
or U1887 (N_1887,N_1783,N_1697);
and U1888 (N_1888,N_1721,N_1722);
and U1889 (N_1889,N_1795,N_1715);
xor U1890 (N_1890,N_1744,N_1714);
or U1891 (N_1891,N_1753,N_1665);
and U1892 (N_1892,N_1689,N_1671);
nor U1893 (N_1893,N_1787,N_1797);
or U1894 (N_1894,N_1659,N_1664);
nor U1895 (N_1895,N_1688,N_1659);
and U1896 (N_1896,N_1674,N_1762);
nor U1897 (N_1897,N_1771,N_1744);
and U1898 (N_1898,N_1673,N_1736);
nor U1899 (N_1899,N_1776,N_1722);
or U1900 (N_1900,N_1683,N_1742);
xnor U1901 (N_1901,N_1780,N_1697);
and U1902 (N_1902,N_1665,N_1719);
or U1903 (N_1903,N_1702,N_1662);
nor U1904 (N_1904,N_1763,N_1683);
nor U1905 (N_1905,N_1773,N_1689);
nor U1906 (N_1906,N_1747,N_1655);
nor U1907 (N_1907,N_1670,N_1779);
nor U1908 (N_1908,N_1716,N_1778);
or U1909 (N_1909,N_1676,N_1660);
or U1910 (N_1910,N_1652,N_1660);
nor U1911 (N_1911,N_1696,N_1713);
or U1912 (N_1912,N_1747,N_1777);
xnor U1913 (N_1913,N_1738,N_1781);
and U1914 (N_1914,N_1661,N_1744);
nor U1915 (N_1915,N_1783,N_1655);
or U1916 (N_1916,N_1658,N_1751);
and U1917 (N_1917,N_1652,N_1786);
nand U1918 (N_1918,N_1702,N_1747);
nor U1919 (N_1919,N_1797,N_1691);
nor U1920 (N_1920,N_1676,N_1695);
and U1921 (N_1921,N_1652,N_1764);
and U1922 (N_1922,N_1667,N_1754);
or U1923 (N_1923,N_1772,N_1673);
nand U1924 (N_1924,N_1776,N_1693);
or U1925 (N_1925,N_1720,N_1717);
nor U1926 (N_1926,N_1672,N_1761);
or U1927 (N_1927,N_1731,N_1683);
nor U1928 (N_1928,N_1741,N_1789);
nor U1929 (N_1929,N_1752,N_1739);
and U1930 (N_1930,N_1724,N_1688);
and U1931 (N_1931,N_1698,N_1683);
nor U1932 (N_1932,N_1717,N_1759);
and U1933 (N_1933,N_1754,N_1685);
or U1934 (N_1934,N_1716,N_1678);
or U1935 (N_1935,N_1797,N_1700);
nand U1936 (N_1936,N_1772,N_1752);
and U1937 (N_1937,N_1746,N_1731);
nor U1938 (N_1938,N_1735,N_1654);
nor U1939 (N_1939,N_1737,N_1683);
and U1940 (N_1940,N_1778,N_1682);
nand U1941 (N_1941,N_1685,N_1672);
and U1942 (N_1942,N_1653,N_1731);
or U1943 (N_1943,N_1777,N_1683);
nor U1944 (N_1944,N_1796,N_1673);
nor U1945 (N_1945,N_1785,N_1679);
or U1946 (N_1946,N_1749,N_1705);
nor U1947 (N_1947,N_1794,N_1677);
and U1948 (N_1948,N_1708,N_1662);
nor U1949 (N_1949,N_1799,N_1778);
and U1950 (N_1950,N_1865,N_1921);
or U1951 (N_1951,N_1856,N_1909);
xor U1952 (N_1952,N_1900,N_1934);
nor U1953 (N_1953,N_1875,N_1833);
or U1954 (N_1954,N_1845,N_1828);
and U1955 (N_1955,N_1882,N_1940);
xor U1956 (N_1956,N_1835,N_1864);
and U1957 (N_1957,N_1808,N_1832);
or U1958 (N_1958,N_1945,N_1894);
nand U1959 (N_1959,N_1830,N_1823);
xnor U1960 (N_1960,N_1863,N_1884);
or U1961 (N_1961,N_1922,N_1820);
nor U1962 (N_1962,N_1851,N_1804);
nand U1963 (N_1963,N_1919,N_1885);
xnor U1964 (N_1964,N_1888,N_1946);
or U1965 (N_1965,N_1893,N_1916);
or U1966 (N_1966,N_1839,N_1889);
nor U1967 (N_1967,N_1924,N_1825);
nand U1968 (N_1968,N_1930,N_1834);
nor U1969 (N_1969,N_1866,N_1812);
nor U1970 (N_1970,N_1891,N_1817);
xor U1971 (N_1971,N_1936,N_1905);
or U1972 (N_1972,N_1932,N_1898);
and U1973 (N_1973,N_1813,N_1824);
xnor U1974 (N_1974,N_1901,N_1841);
nand U1975 (N_1975,N_1897,N_1926);
nand U1976 (N_1976,N_1896,N_1819);
and U1977 (N_1977,N_1861,N_1822);
nand U1978 (N_1978,N_1915,N_1874);
or U1979 (N_1979,N_1800,N_1847);
xnor U1980 (N_1980,N_1801,N_1899);
nor U1981 (N_1981,N_1869,N_1802);
nor U1982 (N_1982,N_1876,N_1877);
nor U1983 (N_1983,N_1938,N_1911);
nor U1984 (N_1984,N_1842,N_1829);
nor U1985 (N_1985,N_1929,N_1852);
and U1986 (N_1986,N_1872,N_1859);
nor U1987 (N_1987,N_1886,N_1927);
and U1988 (N_1988,N_1943,N_1868);
nor U1989 (N_1989,N_1907,N_1844);
and U1990 (N_1990,N_1879,N_1933);
nand U1991 (N_1991,N_1806,N_1913);
or U1992 (N_1992,N_1878,N_1807);
xnor U1993 (N_1993,N_1949,N_1903);
nor U1994 (N_1994,N_1848,N_1892);
and U1995 (N_1995,N_1850,N_1826);
xor U1996 (N_1996,N_1912,N_1805);
or U1997 (N_1997,N_1858,N_1937);
and U1998 (N_1998,N_1855,N_1908);
nand U1999 (N_1999,N_1871,N_1918);
or U2000 (N_2000,N_1810,N_1941);
nor U2001 (N_2001,N_1931,N_1860);
nand U2002 (N_2002,N_1920,N_1942);
nor U2003 (N_2003,N_1948,N_1935);
nand U2004 (N_2004,N_1890,N_1947);
or U2005 (N_2005,N_1838,N_1803);
nor U2006 (N_2006,N_1906,N_1818);
nor U2007 (N_2007,N_1923,N_1914);
nor U2008 (N_2008,N_1846,N_1836);
or U2009 (N_2009,N_1811,N_1925);
or U2010 (N_2010,N_1881,N_1867);
nand U2011 (N_2011,N_1870,N_1862);
xnor U2012 (N_2012,N_1944,N_1857);
or U2013 (N_2013,N_1939,N_1904);
nand U2014 (N_2014,N_1821,N_1849);
nor U2015 (N_2015,N_1809,N_1814);
nor U2016 (N_2016,N_1895,N_1816);
nand U2017 (N_2017,N_1831,N_1815);
nand U2018 (N_2018,N_1887,N_1854);
and U2019 (N_2019,N_1880,N_1873);
or U2020 (N_2020,N_1917,N_1827);
or U2021 (N_2021,N_1853,N_1902);
nand U2022 (N_2022,N_1840,N_1883);
nand U2023 (N_2023,N_1910,N_1837);
nor U2024 (N_2024,N_1928,N_1843);
or U2025 (N_2025,N_1872,N_1854);
nor U2026 (N_2026,N_1819,N_1825);
and U2027 (N_2027,N_1825,N_1886);
nor U2028 (N_2028,N_1926,N_1938);
nor U2029 (N_2029,N_1860,N_1834);
nand U2030 (N_2030,N_1875,N_1863);
xnor U2031 (N_2031,N_1808,N_1852);
or U2032 (N_2032,N_1921,N_1815);
nor U2033 (N_2033,N_1809,N_1856);
and U2034 (N_2034,N_1807,N_1873);
or U2035 (N_2035,N_1850,N_1906);
and U2036 (N_2036,N_1864,N_1926);
nor U2037 (N_2037,N_1884,N_1878);
and U2038 (N_2038,N_1936,N_1877);
xnor U2039 (N_2039,N_1901,N_1940);
nand U2040 (N_2040,N_1870,N_1944);
and U2041 (N_2041,N_1920,N_1947);
nor U2042 (N_2042,N_1801,N_1904);
nand U2043 (N_2043,N_1820,N_1940);
nor U2044 (N_2044,N_1921,N_1948);
nor U2045 (N_2045,N_1853,N_1834);
nand U2046 (N_2046,N_1905,N_1890);
nor U2047 (N_2047,N_1807,N_1919);
nand U2048 (N_2048,N_1927,N_1870);
xnor U2049 (N_2049,N_1895,N_1890);
nor U2050 (N_2050,N_1921,N_1820);
nor U2051 (N_2051,N_1844,N_1897);
nor U2052 (N_2052,N_1909,N_1885);
nor U2053 (N_2053,N_1851,N_1827);
or U2054 (N_2054,N_1919,N_1882);
or U2055 (N_2055,N_1810,N_1895);
and U2056 (N_2056,N_1805,N_1808);
or U2057 (N_2057,N_1800,N_1892);
and U2058 (N_2058,N_1925,N_1924);
and U2059 (N_2059,N_1823,N_1842);
or U2060 (N_2060,N_1893,N_1897);
and U2061 (N_2061,N_1835,N_1833);
and U2062 (N_2062,N_1838,N_1836);
nor U2063 (N_2063,N_1872,N_1921);
or U2064 (N_2064,N_1827,N_1812);
and U2065 (N_2065,N_1847,N_1920);
nor U2066 (N_2066,N_1815,N_1868);
nor U2067 (N_2067,N_1855,N_1854);
and U2068 (N_2068,N_1888,N_1835);
or U2069 (N_2069,N_1835,N_1871);
nor U2070 (N_2070,N_1808,N_1896);
nand U2071 (N_2071,N_1913,N_1948);
nand U2072 (N_2072,N_1813,N_1944);
nor U2073 (N_2073,N_1833,N_1925);
and U2074 (N_2074,N_1847,N_1894);
nand U2075 (N_2075,N_1850,N_1830);
nor U2076 (N_2076,N_1848,N_1883);
or U2077 (N_2077,N_1829,N_1838);
and U2078 (N_2078,N_1873,N_1898);
or U2079 (N_2079,N_1829,N_1892);
nor U2080 (N_2080,N_1820,N_1816);
nor U2081 (N_2081,N_1936,N_1851);
nor U2082 (N_2082,N_1858,N_1805);
nand U2083 (N_2083,N_1824,N_1800);
and U2084 (N_2084,N_1822,N_1867);
and U2085 (N_2085,N_1868,N_1856);
xor U2086 (N_2086,N_1876,N_1896);
nand U2087 (N_2087,N_1870,N_1949);
or U2088 (N_2088,N_1902,N_1903);
or U2089 (N_2089,N_1868,N_1885);
or U2090 (N_2090,N_1904,N_1814);
xor U2091 (N_2091,N_1907,N_1817);
nor U2092 (N_2092,N_1852,N_1937);
and U2093 (N_2093,N_1843,N_1852);
nand U2094 (N_2094,N_1855,N_1897);
and U2095 (N_2095,N_1820,N_1813);
and U2096 (N_2096,N_1806,N_1847);
or U2097 (N_2097,N_1824,N_1873);
nand U2098 (N_2098,N_1816,N_1892);
or U2099 (N_2099,N_1808,N_1899);
and U2100 (N_2100,N_2008,N_2095);
nand U2101 (N_2101,N_2005,N_2062);
or U2102 (N_2102,N_2020,N_1995);
and U2103 (N_2103,N_2001,N_2033);
and U2104 (N_2104,N_1956,N_2056);
xor U2105 (N_2105,N_2026,N_1951);
xnor U2106 (N_2106,N_2073,N_2039);
nor U2107 (N_2107,N_2072,N_2058);
or U2108 (N_2108,N_2040,N_2034);
or U2109 (N_2109,N_2091,N_2070);
nor U2110 (N_2110,N_2088,N_2043);
nor U2111 (N_2111,N_2049,N_2065);
and U2112 (N_2112,N_1968,N_2094);
nor U2113 (N_2113,N_2032,N_1992);
nand U2114 (N_2114,N_2060,N_1990);
nand U2115 (N_2115,N_2059,N_2052);
or U2116 (N_2116,N_2096,N_1982);
and U2117 (N_2117,N_2006,N_2086);
or U2118 (N_2118,N_1981,N_2081);
nor U2119 (N_2119,N_2079,N_1999);
or U2120 (N_2120,N_1994,N_1973);
nand U2121 (N_2121,N_1996,N_2093);
nor U2122 (N_2122,N_2099,N_2046);
or U2123 (N_2123,N_1967,N_1997);
nor U2124 (N_2124,N_2068,N_2044);
or U2125 (N_2125,N_2022,N_2004);
or U2126 (N_2126,N_1972,N_1966);
or U2127 (N_2127,N_1983,N_2063);
nand U2128 (N_2128,N_1952,N_2031);
nand U2129 (N_2129,N_2083,N_1993);
or U2130 (N_2130,N_2097,N_2007);
nor U2131 (N_2131,N_2051,N_2077);
and U2132 (N_2132,N_2038,N_1955);
and U2133 (N_2133,N_1961,N_2017);
nor U2134 (N_2134,N_2054,N_2011);
and U2135 (N_2135,N_1985,N_2015);
or U2136 (N_2136,N_1991,N_2071);
or U2137 (N_2137,N_2069,N_2089);
and U2138 (N_2138,N_2057,N_2024);
nor U2139 (N_2139,N_2041,N_2002);
and U2140 (N_2140,N_1969,N_2053);
and U2141 (N_2141,N_1980,N_1964);
or U2142 (N_2142,N_1988,N_2076);
or U2143 (N_2143,N_2010,N_1987);
and U2144 (N_2144,N_2085,N_2090);
nor U2145 (N_2145,N_2025,N_2080);
and U2146 (N_2146,N_1962,N_2087);
and U2147 (N_2147,N_1963,N_2028);
nand U2148 (N_2148,N_2014,N_2078);
or U2149 (N_2149,N_1975,N_1998);
nor U2150 (N_2150,N_1984,N_1957);
nand U2151 (N_2151,N_1959,N_1950);
and U2152 (N_2152,N_2055,N_2018);
nor U2153 (N_2153,N_1986,N_2019);
nor U2154 (N_2154,N_2064,N_1978);
nor U2155 (N_2155,N_2016,N_1953);
and U2156 (N_2156,N_1974,N_2009);
and U2157 (N_2157,N_1965,N_1960);
or U2158 (N_2158,N_2030,N_2027);
or U2159 (N_2159,N_1989,N_1976);
and U2160 (N_2160,N_2084,N_1977);
nand U2161 (N_2161,N_2047,N_2000);
nor U2162 (N_2162,N_2012,N_1971);
nand U2163 (N_2163,N_2050,N_2067);
nor U2164 (N_2164,N_2036,N_2042);
and U2165 (N_2165,N_1979,N_2029);
nor U2166 (N_2166,N_2023,N_2048);
or U2167 (N_2167,N_2021,N_1970);
xnor U2168 (N_2168,N_2075,N_2045);
or U2169 (N_2169,N_2082,N_2037);
or U2170 (N_2170,N_2035,N_2066);
and U2171 (N_2171,N_2098,N_2061);
and U2172 (N_2172,N_2013,N_2092);
or U2173 (N_2173,N_1958,N_2074);
nor U2174 (N_2174,N_2003,N_1954);
and U2175 (N_2175,N_2047,N_1988);
or U2176 (N_2176,N_2077,N_2003);
or U2177 (N_2177,N_2052,N_2027);
nand U2178 (N_2178,N_2035,N_2067);
and U2179 (N_2179,N_2096,N_2099);
and U2180 (N_2180,N_2096,N_1962);
nor U2181 (N_2181,N_2035,N_2038);
nor U2182 (N_2182,N_2078,N_2030);
nand U2183 (N_2183,N_2079,N_1976);
xnor U2184 (N_2184,N_1986,N_2083);
nand U2185 (N_2185,N_2069,N_2075);
nor U2186 (N_2186,N_2030,N_1974);
or U2187 (N_2187,N_2073,N_2086);
nor U2188 (N_2188,N_2098,N_2004);
xnor U2189 (N_2189,N_2089,N_2088);
nand U2190 (N_2190,N_1956,N_2096);
nand U2191 (N_2191,N_2073,N_2076);
and U2192 (N_2192,N_2002,N_2056);
nand U2193 (N_2193,N_1962,N_1993);
nand U2194 (N_2194,N_2025,N_2017);
nand U2195 (N_2195,N_2054,N_2016);
or U2196 (N_2196,N_1979,N_2065);
or U2197 (N_2197,N_1997,N_2005);
nand U2198 (N_2198,N_2018,N_2090);
nand U2199 (N_2199,N_2049,N_2068);
nor U2200 (N_2200,N_2001,N_2027);
nor U2201 (N_2201,N_2014,N_2061);
nor U2202 (N_2202,N_1977,N_2065);
or U2203 (N_2203,N_2065,N_2066);
or U2204 (N_2204,N_2051,N_1966);
nand U2205 (N_2205,N_1963,N_2069);
nor U2206 (N_2206,N_2000,N_1958);
nand U2207 (N_2207,N_2046,N_2063);
xor U2208 (N_2208,N_2073,N_2080);
nor U2209 (N_2209,N_1958,N_1959);
nor U2210 (N_2210,N_1969,N_2004);
nor U2211 (N_2211,N_2014,N_1984);
and U2212 (N_2212,N_1952,N_2070);
or U2213 (N_2213,N_1999,N_2092);
nor U2214 (N_2214,N_2062,N_1975);
and U2215 (N_2215,N_2043,N_2070);
or U2216 (N_2216,N_2083,N_1958);
nor U2217 (N_2217,N_1975,N_1986);
and U2218 (N_2218,N_2078,N_1973);
and U2219 (N_2219,N_1996,N_2051);
nor U2220 (N_2220,N_2082,N_2065);
nor U2221 (N_2221,N_1955,N_1958);
or U2222 (N_2222,N_2028,N_2083);
nand U2223 (N_2223,N_2068,N_1999);
xor U2224 (N_2224,N_2003,N_2079);
nor U2225 (N_2225,N_1972,N_1995);
nand U2226 (N_2226,N_2065,N_2048);
or U2227 (N_2227,N_1999,N_2013);
nand U2228 (N_2228,N_2019,N_2009);
or U2229 (N_2229,N_1950,N_2023);
nand U2230 (N_2230,N_2014,N_1977);
or U2231 (N_2231,N_1957,N_2013);
nand U2232 (N_2232,N_2093,N_2040);
and U2233 (N_2233,N_2037,N_1985);
and U2234 (N_2234,N_2090,N_2020);
nand U2235 (N_2235,N_1991,N_1967);
nand U2236 (N_2236,N_2078,N_2076);
and U2237 (N_2237,N_2085,N_2053);
nor U2238 (N_2238,N_1994,N_2001);
nand U2239 (N_2239,N_1959,N_1973);
nor U2240 (N_2240,N_2043,N_2023);
or U2241 (N_2241,N_2005,N_2001);
nor U2242 (N_2242,N_2094,N_2075);
xor U2243 (N_2243,N_2066,N_2008);
and U2244 (N_2244,N_1982,N_1966);
or U2245 (N_2245,N_1994,N_2039);
xnor U2246 (N_2246,N_1951,N_2085);
xor U2247 (N_2247,N_2037,N_1981);
or U2248 (N_2248,N_2017,N_2057);
nor U2249 (N_2249,N_1972,N_1961);
nor U2250 (N_2250,N_2181,N_2145);
and U2251 (N_2251,N_2171,N_2180);
or U2252 (N_2252,N_2189,N_2245);
nor U2253 (N_2253,N_2210,N_2163);
nor U2254 (N_2254,N_2108,N_2187);
and U2255 (N_2255,N_2223,N_2191);
nor U2256 (N_2256,N_2235,N_2219);
nand U2257 (N_2257,N_2208,N_2209);
xnor U2258 (N_2258,N_2200,N_2192);
and U2259 (N_2259,N_2213,N_2150);
nor U2260 (N_2260,N_2199,N_2122);
nor U2261 (N_2261,N_2131,N_2128);
nor U2262 (N_2262,N_2142,N_2153);
and U2263 (N_2263,N_2207,N_2143);
and U2264 (N_2264,N_2240,N_2120);
and U2265 (N_2265,N_2100,N_2173);
and U2266 (N_2266,N_2165,N_2156);
nand U2267 (N_2267,N_2129,N_2149);
nor U2268 (N_2268,N_2184,N_2157);
or U2269 (N_2269,N_2111,N_2215);
and U2270 (N_2270,N_2204,N_2241);
and U2271 (N_2271,N_2117,N_2104);
nor U2272 (N_2272,N_2162,N_2221);
nand U2273 (N_2273,N_2196,N_2238);
or U2274 (N_2274,N_2179,N_2211);
nor U2275 (N_2275,N_2225,N_2178);
nor U2276 (N_2276,N_2110,N_2228);
or U2277 (N_2277,N_2114,N_2166);
nand U2278 (N_2278,N_2194,N_2105);
nor U2279 (N_2279,N_2161,N_2107);
nand U2280 (N_2280,N_2169,N_2116);
nand U2281 (N_2281,N_2140,N_2198);
nand U2282 (N_2282,N_2119,N_2126);
nor U2283 (N_2283,N_2172,N_2231);
nand U2284 (N_2284,N_2170,N_2133);
or U2285 (N_2285,N_2159,N_2203);
nor U2286 (N_2286,N_2185,N_2168);
nor U2287 (N_2287,N_2227,N_2109);
or U2288 (N_2288,N_2103,N_2249);
nor U2289 (N_2289,N_2148,N_2236);
nand U2290 (N_2290,N_2222,N_2234);
and U2291 (N_2291,N_2136,N_2121);
nor U2292 (N_2292,N_2127,N_2246);
or U2293 (N_2293,N_2195,N_2124);
and U2294 (N_2294,N_2160,N_2212);
xor U2295 (N_2295,N_2229,N_2239);
or U2296 (N_2296,N_2154,N_2233);
xor U2297 (N_2297,N_2248,N_2147);
or U2298 (N_2298,N_2144,N_2216);
or U2299 (N_2299,N_2183,N_2242);
nor U2300 (N_2300,N_2243,N_2202);
and U2301 (N_2301,N_2175,N_2167);
xnor U2302 (N_2302,N_2177,N_2125);
nand U2303 (N_2303,N_2188,N_2206);
or U2304 (N_2304,N_2138,N_2220);
or U2305 (N_2305,N_2135,N_2218);
nor U2306 (N_2306,N_2123,N_2232);
xor U2307 (N_2307,N_2230,N_2139);
nor U2308 (N_2308,N_2112,N_2158);
nand U2309 (N_2309,N_2151,N_2134);
nand U2310 (N_2310,N_2113,N_2190);
nand U2311 (N_2311,N_2182,N_2155);
or U2312 (N_2312,N_2176,N_2106);
or U2313 (N_2313,N_2137,N_2247);
nand U2314 (N_2314,N_2201,N_2174);
and U2315 (N_2315,N_2226,N_2152);
xnor U2316 (N_2316,N_2237,N_2141);
or U2317 (N_2317,N_2130,N_2164);
and U2318 (N_2318,N_2244,N_2146);
or U2319 (N_2319,N_2217,N_2193);
nor U2320 (N_2320,N_2115,N_2132);
and U2321 (N_2321,N_2224,N_2214);
nand U2322 (N_2322,N_2101,N_2118);
and U2323 (N_2323,N_2186,N_2102);
or U2324 (N_2324,N_2197,N_2205);
nor U2325 (N_2325,N_2112,N_2101);
or U2326 (N_2326,N_2104,N_2231);
or U2327 (N_2327,N_2228,N_2179);
and U2328 (N_2328,N_2173,N_2247);
or U2329 (N_2329,N_2182,N_2163);
nor U2330 (N_2330,N_2132,N_2221);
or U2331 (N_2331,N_2110,N_2118);
nor U2332 (N_2332,N_2196,N_2197);
or U2333 (N_2333,N_2149,N_2183);
and U2334 (N_2334,N_2235,N_2185);
nand U2335 (N_2335,N_2108,N_2214);
and U2336 (N_2336,N_2156,N_2174);
or U2337 (N_2337,N_2165,N_2215);
or U2338 (N_2338,N_2109,N_2138);
and U2339 (N_2339,N_2162,N_2204);
xnor U2340 (N_2340,N_2249,N_2153);
and U2341 (N_2341,N_2178,N_2131);
nor U2342 (N_2342,N_2120,N_2133);
and U2343 (N_2343,N_2244,N_2178);
and U2344 (N_2344,N_2190,N_2180);
and U2345 (N_2345,N_2102,N_2158);
nand U2346 (N_2346,N_2208,N_2113);
nand U2347 (N_2347,N_2168,N_2153);
and U2348 (N_2348,N_2137,N_2120);
xor U2349 (N_2349,N_2188,N_2237);
xor U2350 (N_2350,N_2150,N_2161);
and U2351 (N_2351,N_2136,N_2217);
nand U2352 (N_2352,N_2127,N_2215);
and U2353 (N_2353,N_2155,N_2156);
nor U2354 (N_2354,N_2158,N_2223);
nand U2355 (N_2355,N_2124,N_2114);
and U2356 (N_2356,N_2144,N_2163);
nor U2357 (N_2357,N_2125,N_2208);
nand U2358 (N_2358,N_2207,N_2125);
xnor U2359 (N_2359,N_2148,N_2103);
and U2360 (N_2360,N_2187,N_2110);
nand U2361 (N_2361,N_2214,N_2173);
or U2362 (N_2362,N_2171,N_2123);
or U2363 (N_2363,N_2156,N_2169);
and U2364 (N_2364,N_2132,N_2189);
xor U2365 (N_2365,N_2209,N_2247);
nand U2366 (N_2366,N_2120,N_2198);
nor U2367 (N_2367,N_2243,N_2234);
or U2368 (N_2368,N_2134,N_2121);
and U2369 (N_2369,N_2159,N_2112);
nor U2370 (N_2370,N_2153,N_2141);
and U2371 (N_2371,N_2171,N_2170);
xnor U2372 (N_2372,N_2189,N_2249);
or U2373 (N_2373,N_2219,N_2137);
nor U2374 (N_2374,N_2147,N_2201);
nand U2375 (N_2375,N_2235,N_2125);
nor U2376 (N_2376,N_2222,N_2157);
nand U2377 (N_2377,N_2141,N_2232);
and U2378 (N_2378,N_2138,N_2201);
nor U2379 (N_2379,N_2201,N_2207);
nor U2380 (N_2380,N_2168,N_2209);
or U2381 (N_2381,N_2230,N_2203);
or U2382 (N_2382,N_2189,N_2211);
and U2383 (N_2383,N_2242,N_2195);
or U2384 (N_2384,N_2112,N_2134);
nand U2385 (N_2385,N_2125,N_2145);
or U2386 (N_2386,N_2227,N_2102);
and U2387 (N_2387,N_2143,N_2155);
nor U2388 (N_2388,N_2205,N_2151);
nor U2389 (N_2389,N_2158,N_2180);
and U2390 (N_2390,N_2241,N_2186);
and U2391 (N_2391,N_2103,N_2113);
nor U2392 (N_2392,N_2217,N_2206);
nor U2393 (N_2393,N_2108,N_2126);
xor U2394 (N_2394,N_2191,N_2239);
xnor U2395 (N_2395,N_2141,N_2221);
nand U2396 (N_2396,N_2244,N_2110);
nand U2397 (N_2397,N_2154,N_2105);
and U2398 (N_2398,N_2143,N_2177);
nor U2399 (N_2399,N_2104,N_2189);
and U2400 (N_2400,N_2272,N_2290);
xor U2401 (N_2401,N_2307,N_2334);
nor U2402 (N_2402,N_2319,N_2295);
and U2403 (N_2403,N_2308,N_2380);
or U2404 (N_2404,N_2331,N_2310);
nor U2405 (N_2405,N_2268,N_2372);
nand U2406 (N_2406,N_2366,N_2258);
nor U2407 (N_2407,N_2320,N_2293);
and U2408 (N_2408,N_2377,N_2316);
and U2409 (N_2409,N_2285,N_2361);
and U2410 (N_2410,N_2332,N_2301);
or U2411 (N_2411,N_2254,N_2311);
nor U2412 (N_2412,N_2282,N_2363);
or U2413 (N_2413,N_2382,N_2271);
nor U2414 (N_2414,N_2291,N_2390);
and U2415 (N_2415,N_2396,N_2330);
and U2416 (N_2416,N_2300,N_2348);
nor U2417 (N_2417,N_2356,N_2274);
nand U2418 (N_2418,N_2284,N_2283);
nand U2419 (N_2419,N_2385,N_2278);
nor U2420 (N_2420,N_2297,N_2384);
or U2421 (N_2421,N_2350,N_2399);
xor U2422 (N_2422,N_2263,N_2364);
nand U2423 (N_2423,N_2376,N_2323);
and U2424 (N_2424,N_2303,N_2352);
nor U2425 (N_2425,N_2309,N_2342);
or U2426 (N_2426,N_2313,N_2355);
and U2427 (N_2427,N_2336,N_2260);
nand U2428 (N_2428,N_2280,N_2373);
nor U2429 (N_2429,N_2386,N_2314);
and U2430 (N_2430,N_2353,N_2279);
xor U2431 (N_2431,N_2252,N_2333);
or U2432 (N_2432,N_2292,N_2339);
nand U2433 (N_2433,N_2289,N_2251);
nor U2434 (N_2434,N_2287,N_2337);
nor U2435 (N_2435,N_2349,N_2360);
xnor U2436 (N_2436,N_2265,N_2322);
nand U2437 (N_2437,N_2304,N_2288);
or U2438 (N_2438,N_2388,N_2312);
and U2439 (N_2439,N_2398,N_2344);
xor U2440 (N_2440,N_2394,N_2347);
nor U2441 (N_2441,N_2362,N_2383);
nand U2442 (N_2442,N_2298,N_2275);
or U2443 (N_2443,N_2253,N_2392);
nor U2444 (N_2444,N_2302,N_2257);
nor U2445 (N_2445,N_2286,N_2374);
nor U2446 (N_2446,N_2299,N_2341);
or U2447 (N_2447,N_2294,N_2357);
nor U2448 (N_2448,N_2327,N_2395);
and U2449 (N_2449,N_2378,N_2318);
and U2450 (N_2450,N_2250,N_2375);
nor U2451 (N_2451,N_2305,N_2325);
and U2452 (N_2452,N_2264,N_2351);
xor U2453 (N_2453,N_2259,N_2358);
nand U2454 (N_2454,N_2370,N_2321);
nor U2455 (N_2455,N_2381,N_2393);
nor U2456 (N_2456,N_2340,N_2389);
and U2457 (N_2457,N_2315,N_2379);
and U2458 (N_2458,N_2371,N_2369);
or U2459 (N_2459,N_2269,N_2267);
or U2460 (N_2460,N_2338,N_2368);
nor U2461 (N_2461,N_2277,N_2270);
nand U2462 (N_2462,N_2328,N_2281);
nor U2463 (N_2463,N_2335,N_2354);
or U2464 (N_2464,N_2306,N_2345);
nand U2465 (N_2465,N_2343,N_2367);
and U2466 (N_2466,N_2346,N_2326);
and U2467 (N_2467,N_2387,N_2324);
nor U2468 (N_2468,N_2317,N_2276);
nor U2469 (N_2469,N_2262,N_2266);
nor U2470 (N_2470,N_2365,N_2391);
nand U2471 (N_2471,N_2256,N_2359);
nand U2472 (N_2472,N_2296,N_2255);
nor U2473 (N_2473,N_2273,N_2329);
nand U2474 (N_2474,N_2397,N_2261);
xnor U2475 (N_2475,N_2306,N_2292);
or U2476 (N_2476,N_2390,N_2267);
or U2477 (N_2477,N_2322,N_2348);
nor U2478 (N_2478,N_2397,N_2360);
nor U2479 (N_2479,N_2278,N_2348);
nor U2480 (N_2480,N_2254,N_2379);
or U2481 (N_2481,N_2263,N_2274);
and U2482 (N_2482,N_2331,N_2278);
and U2483 (N_2483,N_2390,N_2271);
nand U2484 (N_2484,N_2358,N_2253);
and U2485 (N_2485,N_2365,N_2336);
nand U2486 (N_2486,N_2322,N_2334);
xnor U2487 (N_2487,N_2321,N_2285);
xnor U2488 (N_2488,N_2294,N_2394);
nor U2489 (N_2489,N_2305,N_2329);
and U2490 (N_2490,N_2350,N_2297);
and U2491 (N_2491,N_2276,N_2257);
nor U2492 (N_2492,N_2261,N_2267);
nor U2493 (N_2493,N_2372,N_2304);
and U2494 (N_2494,N_2252,N_2372);
nor U2495 (N_2495,N_2294,N_2351);
nor U2496 (N_2496,N_2283,N_2341);
nand U2497 (N_2497,N_2358,N_2260);
nand U2498 (N_2498,N_2326,N_2259);
nor U2499 (N_2499,N_2297,N_2355);
or U2500 (N_2500,N_2266,N_2329);
nor U2501 (N_2501,N_2336,N_2322);
nand U2502 (N_2502,N_2284,N_2334);
and U2503 (N_2503,N_2322,N_2392);
nor U2504 (N_2504,N_2290,N_2308);
nand U2505 (N_2505,N_2288,N_2305);
nor U2506 (N_2506,N_2383,N_2325);
and U2507 (N_2507,N_2310,N_2350);
xnor U2508 (N_2508,N_2382,N_2293);
or U2509 (N_2509,N_2288,N_2376);
and U2510 (N_2510,N_2313,N_2372);
or U2511 (N_2511,N_2352,N_2313);
or U2512 (N_2512,N_2273,N_2306);
nand U2513 (N_2513,N_2383,N_2389);
nor U2514 (N_2514,N_2344,N_2302);
or U2515 (N_2515,N_2371,N_2301);
nand U2516 (N_2516,N_2270,N_2391);
xnor U2517 (N_2517,N_2321,N_2296);
or U2518 (N_2518,N_2261,N_2351);
and U2519 (N_2519,N_2304,N_2349);
and U2520 (N_2520,N_2256,N_2288);
and U2521 (N_2521,N_2289,N_2373);
nand U2522 (N_2522,N_2305,N_2373);
nor U2523 (N_2523,N_2377,N_2268);
nand U2524 (N_2524,N_2350,N_2278);
nand U2525 (N_2525,N_2273,N_2274);
or U2526 (N_2526,N_2336,N_2264);
xor U2527 (N_2527,N_2368,N_2390);
or U2528 (N_2528,N_2322,N_2398);
nor U2529 (N_2529,N_2289,N_2256);
xnor U2530 (N_2530,N_2326,N_2382);
nor U2531 (N_2531,N_2340,N_2260);
nor U2532 (N_2532,N_2361,N_2321);
xor U2533 (N_2533,N_2299,N_2355);
and U2534 (N_2534,N_2289,N_2281);
and U2535 (N_2535,N_2390,N_2258);
nor U2536 (N_2536,N_2368,N_2317);
nor U2537 (N_2537,N_2312,N_2350);
and U2538 (N_2538,N_2309,N_2264);
nand U2539 (N_2539,N_2299,N_2328);
nor U2540 (N_2540,N_2388,N_2267);
or U2541 (N_2541,N_2389,N_2265);
and U2542 (N_2542,N_2289,N_2359);
nor U2543 (N_2543,N_2372,N_2278);
nor U2544 (N_2544,N_2338,N_2356);
nand U2545 (N_2545,N_2302,N_2346);
nand U2546 (N_2546,N_2370,N_2337);
nor U2547 (N_2547,N_2311,N_2282);
nand U2548 (N_2548,N_2397,N_2271);
nand U2549 (N_2549,N_2309,N_2312);
nand U2550 (N_2550,N_2423,N_2453);
nand U2551 (N_2551,N_2432,N_2548);
or U2552 (N_2552,N_2431,N_2444);
and U2553 (N_2553,N_2443,N_2524);
xnor U2554 (N_2554,N_2469,N_2459);
nand U2555 (N_2555,N_2497,N_2414);
xnor U2556 (N_2556,N_2531,N_2514);
xor U2557 (N_2557,N_2536,N_2498);
nor U2558 (N_2558,N_2517,N_2437);
and U2559 (N_2559,N_2457,N_2480);
xor U2560 (N_2560,N_2513,N_2434);
nand U2561 (N_2561,N_2523,N_2521);
nor U2562 (N_2562,N_2403,N_2466);
nor U2563 (N_2563,N_2438,N_2463);
and U2564 (N_2564,N_2429,N_2458);
xnor U2565 (N_2565,N_2504,N_2418);
nand U2566 (N_2566,N_2533,N_2449);
and U2567 (N_2567,N_2472,N_2538);
nor U2568 (N_2568,N_2417,N_2507);
or U2569 (N_2569,N_2439,N_2527);
nor U2570 (N_2570,N_2430,N_2467);
nor U2571 (N_2571,N_2542,N_2499);
and U2572 (N_2572,N_2479,N_2428);
xor U2573 (N_2573,N_2446,N_2421);
nand U2574 (N_2574,N_2476,N_2516);
nor U2575 (N_2575,N_2400,N_2435);
nand U2576 (N_2576,N_2519,N_2478);
xnor U2577 (N_2577,N_2481,N_2475);
or U2578 (N_2578,N_2522,N_2473);
nand U2579 (N_2579,N_2515,N_2474);
nand U2580 (N_2580,N_2427,N_2455);
nor U2581 (N_2581,N_2452,N_2545);
and U2582 (N_2582,N_2506,N_2543);
and U2583 (N_2583,N_2407,N_2544);
nor U2584 (N_2584,N_2402,N_2483);
and U2585 (N_2585,N_2501,N_2505);
nor U2586 (N_2586,N_2450,N_2424);
and U2587 (N_2587,N_2535,N_2422);
and U2588 (N_2588,N_2492,N_2461);
or U2589 (N_2589,N_2488,N_2441);
nand U2590 (N_2590,N_2525,N_2528);
and U2591 (N_2591,N_2401,N_2408);
or U2592 (N_2592,N_2532,N_2487);
and U2593 (N_2593,N_2485,N_2433);
and U2594 (N_2594,N_2451,N_2425);
nor U2595 (N_2595,N_2420,N_2413);
and U2596 (N_2596,N_2460,N_2447);
nand U2597 (N_2597,N_2404,N_2415);
nor U2598 (N_2598,N_2489,N_2456);
and U2599 (N_2599,N_2416,N_2491);
or U2600 (N_2600,N_2436,N_2526);
and U2601 (N_2601,N_2454,N_2471);
xnor U2602 (N_2602,N_2529,N_2537);
or U2603 (N_2603,N_2442,N_2494);
nor U2604 (N_2604,N_2468,N_2534);
nand U2605 (N_2605,N_2470,N_2511);
or U2606 (N_2606,N_2465,N_2549);
nand U2607 (N_2607,N_2486,N_2547);
or U2608 (N_2608,N_2490,N_2512);
or U2609 (N_2609,N_2412,N_2409);
or U2610 (N_2610,N_2495,N_2508);
and U2611 (N_2611,N_2541,N_2405);
or U2612 (N_2612,N_2502,N_2509);
nand U2613 (N_2613,N_2445,N_2484);
nand U2614 (N_2614,N_2448,N_2510);
nor U2615 (N_2615,N_2540,N_2503);
or U2616 (N_2616,N_2482,N_2464);
or U2617 (N_2617,N_2419,N_2539);
nor U2618 (N_2618,N_2411,N_2493);
and U2619 (N_2619,N_2426,N_2546);
and U2620 (N_2620,N_2520,N_2410);
and U2621 (N_2621,N_2496,N_2406);
or U2622 (N_2622,N_2500,N_2462);
nor U2623 (N_2623,N_2477,N_2518);
or U2624 (N_2624,N_2440,N_2530);
xnor U2625 (N_2625,N_2527,N_2518);
or U2626 (N_2626,N_2461,N_2419);
and U2627 (N_2627,N_2421,N_2450);
nand U2628 (N_2628,N_2483,N_2420);
or U2629 (N_2629,N_2426,N_2543);
nand U2630 (N_2630,N_2401,N_2419);
nor U2631 (N_2631,N_2482,N_2516);
or U2632 (N_2632,N_2409,N_2400);
and U2633 (N_2633,N_2471,N_2404);
or U2634 (N_2634,N_2477,N_2449);
nor U2635 (N_2635,N_2410,N_2471);
nor U2636 (N_2636,N_2400,N_2426);
or U2637 (N_2637,N_2471,N_2431);
or U2638 (N_2638,N_2406,N_2432);
nand U2639 (N_2639,N_2505,N_2510);
nand U2640 (N_2640,N_2486,N_2499);
or U2641 (N_2641,N_2487,N_2540);
and U2642 (N_2642,N_2507,N_2472);
or U2643 (N_2643,N_2401,N_2534);
or U2644 (N_2644,N_2540,N_2510);
or U2645 (N_2645,N_2440,N_2507);
nor U2646 (N_2646,N_2405,N_2410);
nor U2647 (N_2647,N_2510,N_2423);
xor U2648 (N_2648,N_2509,N_2532);
nand U2649 (N_2649,N_2452,N_2499);
and U2650 (N_2650,N_2450,N_2447);
nor U2651 (N_2651,N_2428,N_2421);
nand U2652 (N_2652,N_2537,N_2426);
and U2653 (N_2653,N_2521,N_2502);
nand U2654 (N_2654,N_2444,N_2422);
nand U2655 (N_2655,N_2536,N_2402);
or U2656 (N_2656,N_2541,N_2526);
nand U2657 (N_2657,N_2524,N_2420);
xnor U2658 (N_2658,N_2547,N_2506);
or U2659 (N_2659,N_2462,N_2474);
nand U2660 (N_2660,N_2501,N_2425);
nand U2661 (N_2661,N_2452,N_2547);
nor U2662 (N_2662,N_2449,N_2404);
nor U2663 (N_2663,N_2474,N_2419);
or U2664 (N_2664,N_2402,N_2478);
or U2665 (N_2665,N_2488,N_2423);
xor U2666 (N_2666,N_2496,N_2499);
or U2667 (N_2667,N_2473,N_2513);
nand U2668 (N_2668,N_2485,N_2492);
or U2669 (N_2669,N_2422,N_2532);
nand U2670 (N_2670,N_2516,N_2541);
nand U2671 (N_2671,N_2424,N_2453);
nand U2672 (N_2672,N_2542,N_2543);
and U2673 (N_2673,N_2476,N_2534);
and U2674 (N_2674,N_2456,N_2499);
xor U2675 (N_2675,N_2441,N_2428);
nand U2676 (N_2676,N_2475,N_2536);
nand U2677 (N_2677,N_2519,N_2544);
nor U2678 (N_2678,N_2538,N_2440);
nor U2679 (N_2679,N_2523,N_2511);
nand U2680 (N_2680,N_2493,N_2517);
nand U2681 (N_2681,N_2438,N_2422);
or U2682 (N_2682,N_2446,N_2425);
nand U2683 (N_2683,N_2485,N_2474);
and U2684 (N_2684,N_2541,N_2533);
nor U2685 (N_2685,N_2494,N_2473);
xnor U2686 (N_2686,N_2489,N_2502);
xor U2687 (N_2687,N_2481,N_2510);
nor U2688 (N_2688,N_2548,N_2436);
nor U2689 (N_2689,N_2482,N_2422);
nor U2690 (N_2690,N_2502,N_2499);
or U2691 (N_2691,N_2509,N_2446);
xor U2692 (N_2692,N_2521,N_2470);
xnor U2693 (N_2693,N_2433,N_2494);
or U2694 (N_2694,N_2491,N_2502);
or U2695 (N_2695,N_2458,N_2460);
or U2696 (N_2696,N_2419,N_2488);
and U2697 (N_2697,N_2510,N_2517);
nand U2698 (N_2698,N_2452,N_2463);
and U2699 (N_2699,N_2469,N_2465);
xor U2700 (N_2700,N_2614,N_2688);
or U2701 (N_2701,N_2669,N_2588);
and U2702 (N_2702,N_2660,N_2643);
nor U2703 (N_2703,N_2573,N_2689);
nor U2704 (N_2704,N_2691,N_2628);
nand U2705 (N_2705,N_2570,N_2562);
nor U2706 (N_2706,N_2682,N_2574);
nand U2707 (N_2707,N_2676,N_2593);
xnor U2708 (N_2708,N_2563,N_2634);
nor U2709 (N_2709,N_2571,N_2678);
nor U2710 (N_2710,N_2603,N_2648);
nand U2711 (N_2711,N_2613,N_2637);
nand U2712 (N_2712,N_2619,N_2604);
xnor U2713 (N_2713,N_2679,N_2630);
or U2714 (N_2714,N_2599,N_2657);
nand U2715 (N_2715,N_2605,N_2572);
or U2716 (N_2716,N_2560,N_2677);
nand U2717 (N_2717,N_2653,N_2592);
or U2718 (N_2718,N_2683,N_2615);
and U2719 (N_2719,N_2641,N_2594);
nor U2720 (N_2720,N_2612,N_2597);
and U2721 (N_2721,N_2566,N_2576);
and U2722 (N_2722,N_2622,N_2556);
and U2723 (N_2723,N_2557,N_2674);
xnor U2724 (N_2724,N_2693,N_2681);
nand U2725 (N_2725,N_2649,N_2697);
and U2726 (N_2726,N_2647,N_2694);
xor U2727 (N_2727,N_2579,N_2554);
and U2728 (N_2728,N_2655,N_2591);
nor U2729 (N_2729,N_2640,N_2684);
and U2730 (N_2730,N_2661,N_2668);
or U2731 (N_2731,N_2629,N_2555);
or U2732 (N_2732,N_2602,N_2635);
nor U2733 (N_2733,N_2636,N_2652);
nand U2734 (N_2734,N_2582,N_2550);
nand U2735 (N_2735,N_2551,N_2624);
and U2736 (N_2736,N_2558,N_2561);
nand U2737 (N_2737,N_2598,N_2609);
nand U2738 (N_2738,N_2675,N_2610);
and U2739 (N_2739,N_2663,N_2618);
nor U2740 (N_2740,N_2621,N_2617);
and U2741 (N_2741,N_2656,N_2578);
or U2742 (N_2742,N_2627,N_2699);
or U2743 (N_2743,N_2631,N_2575);
nand U2744 (N_2744,N_2698,N_2671);
or U2745 (N_2745,N_2644,N_2586);
xnor U2746 (N_2746,N_2662,N_2685);
nor U2747 (N_2747,N_2639,N_2606);
nand U2748 (N_2748,N_2616,N_2658);
xor U2749 (N_2749,N_2585,N_2600);
xnor U2750 (N_2750,N_2553,N_2568);
or U2751 (N_2751,N_2589,N_2583);
nor U2752 (N_2752,N_2667,N_2611);
nand U2753 (N_2753,N_2587,N_2664);
nor U2754 (N_2754,N_2673,N_2577);
nand U2755 (N_2755,N_2650,N_2659);
nor U2756 (N_2756,N_2666,N_2638);
nor U2757 (N_2757,N_2665,N_2565);
nand U2758 (N_2758,N_2625,N_2695);
nand U2759 (N_2759,N_2646,N_2623);
xnor U2760 (N_2760,N_2651,N_2559);
nand U2761 (N_2761,N_2581,N_2552);
nand U2762 (N_2762,N_2670,N_2632);
or U2763 (N_2763,N_2626,N_2569);
and U2764 (N_2764,N_2672,N_2620);
nor U2765 (N_2765,N_2608,N_2580);
nand U2766 (N_2766,N_2690,N_2687);
and U2767 (N_2767,N_2654,N_2633);
nand U2768 (N_2768,N_2642,N_2696);
nand U2769 (N_2769,N_2567,N_2596);
nor U2770 (N_2770,N_2680,N_2607);
nand U2771 (N_2771,N_2601,N_2686);
or U2772 (N_2772,N_2584,N_2692);
nor U2773 (N_2773,N_2595,N_2590);
xor U2774 (N_2774,N_2564,N_2645);
and U2775 (N_2775,N_2606,N_2646);
nand U2776 (N_2776,N_2580,N_2689);
nor U2777 (N_2777,N_2639,N_2594);
and U2778 (N_2778,N_2635,N_2658);
and U2779 (N_2779,N_2621,N_2696);
nand U2780 (N_2780,N_2676,N_2658);
nor U2781 (N_2781,N_2568,N_2550);
nand U2782 (N_2782,N_2626,N_2688);
nor U2783 (N_2783,N_2606,N_2677);
or U2784 (N_2784,N_2630,N_2627);
nand U2785 (N_2785,N_2615,N_2600);
or U2786 (N_2786,N_2673,N_2686);
nand U2787 (N_2787,N_2683,N_2638);
xor U2788 (N_2788,N_2685,N_2668);
nand U2789 (N_2789,N_2685,N_2688);
or U2790 (N_2790,N_2601,N_2654);
and U2791 (N_2791,N_2695,N_2603);
or U2792 (N_2792,N_2571,N_2662);
or U2793 (N_2793,N_2656,N_2654);
and U2794 (N_2794,N_2679,N_2567);
and U2795 (N_2795,N_2681,N_2676);
or U2796 (N_2796,N_2612,N_2655);
or U2797 (N_2797,N_2642,N_2698);
and U2798 (N_2798,N_2643,N_2557);
or U2799 (N_2799,N_2605,N_2585);
or U2800 (N_2800,N_2607,N_2636);
nor U2801 (N_2801,N_2671,N_2584);
and U2802 (N_2802,N_2567,N_2658);
and U2803 (N_2803,N_2665,N_2606);
nor U2804 (N_2804,N_2674,N_2697);
or U2805 (N_2805,N_2650,N_2619);
xnor U2806 (N_2806,N_2590,N_2685);
nor U2807 (N_2807,N_2694,N_2646);
and U2808 (N_2808,N_2672,N_2556);
nand U2809 (N_2809,N_2560,N_2678);
or U2810 (N_2810,N_2669,N_2649);
nor U2811 (N_2811,N_2612,N_2660);
and U2812 (N_2812,N_2577,N_2638);
nand U2813 (N_2813,N_2563,N_2582);
nor U2814 (N_2814,N_2650,N_2697);
and U2815 (N_2815,N_2679,N_2688);
nand U2816 (N_2816,N_2695,N_2571);
and U2817 (N_2817,N_2628,N_2699);
nor U2818 (N_2818,N_2561,N_2582);
and U2819 (N_2819,N_2634,N_2617);
nor U2820 (N_2820,N_2570,N_2594);
or U2821 (N_2821,N_2601,N_2663);
or U2822 (N_2822,N_2583,N_2574);
and U2823 (N_2823,N_2576,N_2673);
xnor U2824 (N_2824,N_2556,N_2558);
and U2825 (N_2825,N_2606,N_2576);
nand U2826 (N_2826,N_2607,N_2679);
or U2827 (N_2827,N_2635,N_2687);
nor U2828 (N_2828,N_2593,N_2695);
nor U2829 (N_2829,N_2657,N_2681);
or U2830 (N_2830,N_2583,N_2564);
xor U2831 (N_2831,N_2551,N_2622);
or U2832 (N_2832,N_2691,N_2596);
nand U2833 (N_2833,N_2619,N_2661);
or U2834 (N_2834,N_2692,N_2695);
and U2835 (N_2835,N_2609,N_2697);
nor U2836 (N_2836,N_2571,N_2666);
or U2837 (N_2837,N_2598,N_2623);
and U2838 (N_2838,N_2663,N_2552);
or U2839 (N_2839,N_2676,N_2672);
xnor U2840 (N_2840,N_2631,N_2673);
and U2841 (N_2841,N_2682,N_2615);
or U2842 (N_2842,N_2691,N_2606);
or U2843 (N_2843,N_2555,N_2638);
or U2844 (N_2844,N_2576,N_2678);
or U2845 (N_2845,N_2592,N_2600);
nand U2846 (N_2846,N_2606,N_2694);
xnor U2847 (N_2847,N_2591,N_2667);
and U2848 (N_2848,N_2573,N_2583);
and U2849 (N_2849,N_2689,N_2664);
and U2850 (N_2850,N_2806,N_2711);
and U2851 (N_2851,N_2768,N_2762);
xor U2852 (N_2852,N_2810,N_2802);
and U2853 (N_2853,N_2775,N_2735);
xnor U2854 (N_2854,N_2812,N_2838);
and U2855 (N_2855,N_2710,N_2842);
nor U2856 (N_2856,N_2714,N_2736);
nand U2857 (N_2857,N_2748,N_2771);
or U2858 (N_2858,N_2799,N_2731);
and U2859 (N_2859,N_2786,N_2707);
nand U2860 (N_2860,N_2787,N_2840);
nand U2861 (N_2861,N_2738,N_2796);
and U2862 (N_2862,N_2844,N_2811);
and U2863 (N_2863,N_2713,N_2849);
nand U2864 (N_2864,N_2830,N_2766);
nor U2865 (N_2865,N_2832,N_2753);
or U2866 (N_2866,N_2730,N_2788);
xnor U2867 (N_2867,N_2760,N_2700);
nor U2868 (N_2868,N_2750,N_2761);
or U2869 (N_2869,N_2732,N_2848);
nand U2870 (N_2870,N_2729,N_2719);
xnor U2871 (N_2871,N_2767,N_2747);
nand U2872 (N_2872,N_2825,N_2827);
nand U2873 (N_2873,N_2764,N_2720);
nor U2874 (N_2874,N_2745,N_2826);
nor U2875 (N_2875,N_2726,N_2723);
and U2876 (N_2876,N_2807,N_2772);
nand U2877 (N_2877,N_2733,N_2743);
nor U2878 (N_2878,N_2789,N_2784);
and U2879 (N_2879,N_2763,N_2773);
nor U2880 (N_2880,N_2746,N_2722);
nand U2881 (N_2881,N_2847,N_2846);
or U2882 (N_2882,N_2823,N_2749);
nand U2883 (N_2883,N_2824,N_2765);
or U2884 (N_2884,N_2782,N_2790);
nor U2885 (N_2885,N_2769,N_2833);
nand U2886 (N_2886,N_2702,N_2803);
and U2887 (N_2887,N_2834,N_2754);
and U2888 (N_2888,N_2737,N_2839);
nand U2889 (N_2889,N_2739,N_2814);
nand U2890 (N_2890,N_2752,N_2703);
and U2891 (N_2891,N_2785,N_2800);
and U2892 (N_2892,N_2835,N_2706);
xnor U2893 (N_2893,N_2780,N_2818);
nor U2894 (N_2894,N_2819,N_2740);
and U2895 (N_2895,N_2721,N_2841);
nand U2896 (N_2896,N_2815,N_2717);
nor U2897 (N_2897,N_2822,N_2843);
and U2898 (N_2898,N_2777,N_2741);
or U2899 (N_2899,N_2783,N_2791);
or U2900 (N_2900,N_2774,N_2770);
and U2901 (N_2901,N_2758,N_2813);
nor U2902 (N_2902,N_2808,N_2701);
nand U2903 (N_2903,N_2781,N_2798);
and U2904 (N_2904,N_2794,N_2709);
xor U2905 (N_2905,N_2821,N_2718);
or U2906 (N_2906,N_2829,N_2797);
nand U2907 (N_2907,N_2805,N_2704);
and U2908 (N_2908,N_2836,N_2837);
or U2909 (N_2909,N_2820,N_2734);
and U2910 (N_2910,N_2757,N_2716);
nand U2911 (N_2911,N_2828,N_2816);
nand U2912 (N_2912,N_2792,N_2712);
and U2913 (N_2913,N_2708,N_2751);
and U2914 (N_2914,N_2804,N_2724);
nor U2915 (N_2915,N_2817,N_2756);
nor U2916 (N_2916,N_2744,N_2795);
nand U2917 (N_2917,N_2809,N_2755);
or U2918 (N_2918,N_2793,N_2759);
and U2919 (N_2919,N_2801,N_2779);
nand U2920 (N_2920,N_2725,N_2776);
or U2921 (N_2921,N_2728,N_2742);
and U2922 (N_2922,N_2727,N_2831);
nor U2923 (N_2923,N_2845,N_2705);
and U2924 (N_2924,N_2778,N_2715);
and U2925 (N_2925,N_2780,N_2762);
xor U2926 (N_2926,N_2736,N_2717);
nand U2927 (N_2927,N_2772,N_2784);
nor U2928 (N_2928,N_2837,N_2819);
nand U2929 (N_2929,N_2728,N_2706);
nor U2930 (N_2930,N_2718,N_2781);
or U2931 (N_2931,N_2732,N_2810);
and U2932 (N_2932,N_2751,N_2761);
or U2933 (N_2933,N_2835,N_2848);
or U2934 (N_2934,N_2839,N_2733);
and U2935 (N_2935,N_2713,N_2739);
nand U2936 (N_2936,N_2758,N_2721);
or U2937 (N_2937,N_2790,N_2703);
or U2938 (N_2938,N_2782,N_2774);
nor U2939 (N_2939,N_2758,N_2707);
xnor U2940 (N_2940,N_2811,N_2817);
nor U2941 (N_2941,N_2823,N_2814);
or U2942 (N_2942,N_2757,N_2736);
or U2943 (N_2943,N_2746,N_2797);
or U2944 (N_2944,N_2735,N_2817);
nand U2945 (N_2945,N_2721,N_2746);
xnor U2946 (N_2946,N_2772,N_2751);
nor U2947 (N_2947,N_2723,N_2802);
or U2948 (N_2948,N_2773,N_2841);
and U2949 (N_2949,N_2843,N_2764);
or U2950 (N_2950,N_2725,N_2782);
or U2951 (N_2951,N_2825,N_2766);
and U2952 (N_2952,N_2752,N_2730);
nor U2953 (N_2953,N_2752,N_2724);
nor U2954 (N_2954,N_2794,N_2745);
nor U2955 (N_2955,N_2813,N_2790);
nor U2956 (N_2956,N_2754,N_2707);
and U2957 (N_2957,N_2764,N_2802);
nor U2958 (N_2958,N_2779,N_2791);
and U2959 (N_2959,N_2730,N_2748);
nor U2960 (N_2960,N_2768,N_2764);
or U2961 (N_2961,N_2830,N_2761);
nor U2962 (N_2962,N_2791,N_2711);
nand U2963 (N_2963,N_2704,N_2785);
xnor U2964 (N_2964,N_2751,N_2713);
and U2965 (N_2965,N_2763,N_2805);
nand U2966 (N_2966,N_2767,N_2843);
xor U2967 (N_2967,N_2774,N_2742);
nor U2968 (N_2968,N_2827,N_2847);
nor U2969 (N_2969,N_2806,N_2836);
xnor U2970 (N_2970,N_2831,N_2715);
xnor U2971 (N_2971,N_2749,N_2707);
or U2972 (N_2972,N_2780,N_2727);
and U2973 (N_2973,N_2826,N_2842);
nand U2974 (N_2974,N_2760,N_2803);
nand U2975 (N_2975,N_2770,N_2818);
and U2976 (N_2976,N_2803,N_2801);
or U2977 (N_2977,N_2754,N_2820);
or U2978 (N_2978,N_2739,N_2784);
nor U2979 (N_2979,N_2720,N_2750);
nand U2980 (N_2980,N_2823,N_2825);
and U2981 (N_2981,N_2757,N_2715);
or U2982 (N_2982,N_2743,N_2804);
and U2983 (N_2983,N_2749,N_2783);
or U2984 (N_2984,N_2831,N_2846);
nor U2985 (N_2985,N_2737,N_2714);
nor U2986 (N_2986,N_2844,N_2720);
or U2987 (N_2987,N_2747,N_2824);
xor U2988 (N_2988,N_2819,N_2737);
xor U2989 (N_2989,N_2806,N_2725);
nor U2990 (N_2990,N_2848,N_2849);
xnor U2991 (N_2991,N_2791,N_2793);
and U2992 (N_2992,N_2727,N_2848);
xnor U2993 (N_2993,N_2763,N_2705);
or U2994 (N_2994,N_2740,N_2830);
and U2995 (N_2995,N_2780,N_2742);
or U2996 (N_2996,N_2717,N_2712);
nor U2997 (N_2997,N_2702,N_2795);
or U2998 (N_2998,N_2819,N_2795);
nor U2999 (N_2999,N_2732,N_2839);
or U3000 (N_3000,N_2854,N_2929);
nor U3001 (N_3001,N_2905,N_2993);
or U3002 (N_3002,N_2968,N_2872);
nor U3003 (N_3003,N_2878,N_2886);
xor U3004 (N_3004,N_2917,N_2920);
and U3005 (N_3005,N_2909,N_2856);
and U3006 (N_3006,N_2935,N_2932);
nor U3007 (N_3007,N_2904,N_2894);
nor U3008 (N_3008,N_2998,N_2992);
nor U3009 (N_3009,N_2960,N_2959);
and U3010 (N_3010,N_2943,N_2939);
or U3011 (N_3011,N_2956,N_2906);
nand U3012 (N_3012,N_2891,N_2850);
nand U3013 (N_3013,N_2977,N_2896);
and U3014 (N_3014,N_2936,N_2966);
or U3015 (N_3015,N_2903,N_2874);
nor U3016 (N_3016,N_2915,N_2884);
nor U3017 (N_3017,N_2898,N_2927);
or U3018 (N_3018,N_2853,N_2889);
or U3019 (N_3019,N_2969,N_2997);
nand U3020 (N_3020,N_2976,N_2875);
nand U3021 (N_3021,N_2924,N_2912);
nand U3022 (N_3022,N_2881,N_2910);
and U3023 (N_3023,N_2888,N_2944);
and U3024 (N_3024,N_2978,N_2855);
nor U3025 (N_3025,N_2858,N_2961);
nand U3026 (N_3026,N_2852,N_2964);
nor U3027 (N_3027,N_2907,N_2965);
or U3028 (N_3028,N_2922,N_2895);
nor U3029 (N_3029,N_2864,N_2983);
and U3030 (N_3030,N_2952,N_2989);
nor U3031 (N_3031,N_2911,N_2971);
or U3032 (N_3032,N_2974,N_2908);
or U3033 (N_3033,N_2879,N_2948);
nor U3034 (N_3034,N_2933,N_2876);
xnor U3035 (N_3035,N_2885,N_2962);
or U3036 (N_3036,N_2901,N_2902);
and U3037 (N_3037,N_2954,N_2914);
nand U3038 (N_3038,N_2860,N_2867);
and U3039 (N_3039,N_2893,N_2930);
or U3040 (N_3040,N_2980,N_2923);
nor U3041 (N_3041,N_2985,N_2851);
nor U3042 (N_3042,N_2925,N_2892);
and U3043 (N_3043,N_2987,N_2958);
nand U3044 (N_3044,N_2950,N_2940);
or U3045 (N_3045,N_2859,N_2880);
and U3046 (N_3046,N_2870,N_2866);
nor U3047 (N_3047,N_2955,N_2938);
and U3048 (N_3048,N_2890,N_2900);
or U3049 (N_3049,N_2986,N_2897);
or U3050 (N_3050,N_2995,N_2979);
or U3051 (N_3051,N_2973,N_2934);
and U3052 (N_3052,N_2899,N_2953);
nand U3053 (N_3053,N_2921,N_2967);
or U3054 (N_3054,N_2931,N_2941);
and U3055 (N_3055,N_2957,N_2877);
xor U3056 (N_3056,N_2942,N_2865);
or U3057 (N_3057,N_2975,N_2991);
or U3058 (N_3058,N_2926,N_2951);
nor U3059 (N_3059,N_2913,N_2869);
nor U3060 (N_3060,N_2883,N_2994);
nor U3061 (N_3061,N_2871,N_2947);
nor U3062 (N_3062,N_2862,N_2919);
nor U3063 (N_3063,N_2916,N_2972);
nand U3064 (N_3064,N_2857,N_2970);
or U3065 (N_3065,N_2861,N_2945);
xor U3066 (N_3066,N_2946,N_2882);
nor U3067 (N_3067,N_2990,N_2937);
and U3068 (N_3068,N_2963,N_2887);
nand U3069 (N_3069,N_2984,N_2873);
and U3070 (N_3070,N_2928,N_2868);
and U3071 (N_3071,N_2988,N_2982);
and U3072 (N_3072,N_2996,N_2999);
or U3073 (N_3073,N_2981,N_2918);
and U3074 (N_3074,N_2949,N_2863);
nor U3075 (N_3075,N_2909,N_2951);
and U3076 (N_3076,N_2945,N_2875);
and U3077 (N_3077,N_2922,N_2983);
or U3078 (N_3078,N_2896,N_2926);
xnor U3079 (N_3079,N_2969,N_2993);
nor U3080 (N_3080,N_2912,N_2914);
and U3081 (N_3081,N_2947,N_2948);
nor U3082 (N_3082,N_2929,N_2893);
and U3083 (N_3083,N_2889,N_2906);
nor U3084 (N_3084,N_2978,N_2860);
nand U3085 (N_3085,N_2852,N_2917);
or U3086 (N_3086,N_2853,N_2932);
and U3087 (N_3087,N_2984,N_2989);
and U3088 (N_3088,N_2892,N_2895);
or U3089 (N_3089,N_2951,N_2875);
nor U3090 (N_3090,N_2926,N_2996);
and U3091 (N_3091,N_2885,N_2949);
xnor U3092 (N_3092,N_2967,N_2942);
xnor U3093 (N_3093,N_2921,N_2857);
and U3094 (N_3094,N_2861,N_2994);
or U3095 (N_3095,N_2948,N_2916);
nand U3096 (N_3096,N_2931,N_2870);
nor U3097 (N_3097,N_2993,N_2936);
or U3098 (N_3098,N_2987,N_2946);
nand U3099 (N_3099,N_2985,N_2879);
or U3100 (N_3100,N_2936,N_2972);
nand U3101 (N_3101,N_2978,N_2929);
or U3102 (N_3102,N_2925,N_2854);
nor U3103 (N_3103,N_2957,N_2994);
nor U3104 (N_3104,N_2954,N_2970);
nand U3105 (N_3105,N_2972,N_2996);
and U3106 (N_3106,N_2979,N_2922);
and U3107 (N_3107,N_2872,N_2860);
nor U3108 (N_3108,N_2926,N_2978);
nand U3109 (N_3109,N_2940,N_2916);
and U3110 (N_3110,N_2948,N_2871);
or U3111 (N_3111,N_2868,N_2943);
and U3112 (N_3112,N_2970,N_2972);
nor U3113 (N_3113,N_2927,N_2855);
nor U3114 (N_3114,N_2954,N_2917);
or U3115 (N_3115,N_2994,N_2914);
or U3116 (N_3116,N_2963,N_2941);
nor U3117 (N_3117,N_2951,N_2945);
or U3118 (N_3118,N_2875,N_2957);
and U3119 (N_3119,N_2990,N_2974);
nor U3120 (N_3120,N_2894,N_2940);
nor U3121 (N_3121,N_2909,N_2924);
and U3122 (N_3122,N_2949,N_2998);
or U3123 (N_3123,N_2859,N_2933);
nor U3124 (N_3124,N_2926,N_2867);
nand U3125 (N_3125,N_2975,N_2967);
and U3126 (N_3126,N_2884,N_2901);
or U3127 (N_3127,N_2938,N_2890);
xnor U3128 (N_3128,N_2917,N_2906);
or U3129 (N_3129,N_2965,N_2924);
or U3130 (N_3130,N_2989,N_2853);
xnor U3131 (N_3131,N_2852,N_2923);
and U3132 (N_3132,N_2904,N_2874);
xnor U3133 (N_3133,N_2966,N_2916);
xnor U3134 (N_3134,N_2856,N_2985);
nand U3135 (N_3135,N_2955,N_2933);
and U3136 (N_3136,N_2904,N_2986);
and U3137 (N_3137,N_2941,N_2943);
or U3138 (N_3138,N_2923,N_2866);
or U3139 (N_3139,N_2912,N_2935);
xor U3140 (N_3140,N_2992,N_2890);
nand U3141 (N_3141,N_2902,N_2949);
or U3142 (N_3142,N_2995,N_2976);
or U3143 (N_3143,N_2982,N_2974);
nand U3144 (N_3144,N_2887,N_2961);
xnor U3145 (N_3145,N_2947,N_2889);
nor U3146 (N_3146,N_2852,N_2961);
nand U3147 (N_3147,N_2863,N_2884);
or U3148 (N_3148,N_2887,N_2983);
nand U3149 (N_3149,N_2889,N_2891);
or U3150 (N_3150,N_3124,N_3029);
nor U3151 (N_3151,N_3074,N_3054);
and U3152 (N_3152,N_3079,N_3114);
nor U3153 (N_3153,N_3131,N_3119);
nor U3154 (N_3154,N_3021,N_3042);
nor U3155 (N_3155,N_3082,N_3049);
and U3156 (N_3156,N_3084,N_3093);
nand U3157 (N_3157,N_3147,N_3098);
or U3158 (N_3158,N_3100,N_3135);
nand U3159 (N_3159,N_3089,N_3145);
nor U3160 (N_3160,N_3019,N_3081);
nor U3161 (N_3161,N_3051,N_3032);
or U3162 (N_3162,N_3066,N_3112);
nand U3163 (N_3163,N_3106,N_3103);
or U3164 (N_3164,N_3121,N_3075);
xor U3165 (N_3165,N_3039,N_3091);
nor U3166 (N_3166,N_3025,N_3101);
xor U3167 (N_3167,N_3016,N_3050);
nand U3168 (N_3168,N_3120,N_3006);
nor U3169 (N_3169,N_3001,N_3085);
and U3170 (N_3170,N_3064,N_3130);
nand U3171 (N_3171,N_3095,N_3113);
or U3172 (N_3172,N_3069,N_3127);
or U3173 (N_3173,N_3014,N_3140);
or U3174 (N_3174,N_3073,N_3088);
and U3175 (N_3175,N_3068,N_3026);
or U3176 (N_3176,N_3020,N_3031);
xnor U3177 (N_3177,N_3144,N_3022);
nor U3178 (N_3178,N_3062,N_3077);
and U3179 (N_3179,N_3004,N_3107);
nor U3180 (N_3180,N_3015,N_3109);
nor U3181 (N_3181,N_3046,N_3010);
or U3182 (N_3182,N_3133,N_3102);
and U3183 (N_3183,N_3137,N_3036);
and U3184 (N_3184,N_3094,N_3012);
or U3185 (N_3185,N_3055,N_3040);
and U3186 (N_3186,N_3017,N_3061);
nand U3187 (N_3187,N_3065,N_3000);
xnor U3188 (N_3188,N_3057,N_3033);
nand U3189 (N_3189,N_3059,N_3034);
or U3190 (N_3190,N_3018,N_3087);
and U3191 (N_3191,N_3125,N_3141);
nor U3192 (N_3192,N_3083,N_3013);
nor U3193 (N_3193,N_3071,N_3110);
xnor U3194 (N_3194,N_3070,N_3008);
or U3195 (N_3195,N_3105,N_3038);
nand U3196 (N_3196,N_3027,N_3134);
or U3197 (N_3197,N_3037,N_3148);
xnor U3198 (N_3198,N_3048,N_3090);
nand U3199 (N_3199,N_3096,N_3009);
nor U3200 (N_3200,N_3104,N_3142);
xor U3201 (N_3201,N_3005,N_3146);
or U3202 (N_3202,N_3007,N_3128);
and U3203 (N_3203,N_3086,N_3116);
nor U3204 (N_3204,N_3117,N_3002);
nand U3205 (N_3205,N_3011,N_3136);
and U3206 (N_3206,N_3149,N_3115);
or U3207 (N_3207,N_3139,N_3129);
nand U3208 (N_3208,N_3122,N_3044);
nor U3209 (N_3209,N_3092,N_3097);
or U3210 (N_3210,N_3052,N_3123);
nor U3211 (N_3211,N_3023,N_3080);
nor U3212 (N_3212,N_3067,N_3043);
nand U3213 (N_3213,N_3053,N_3045);
and U3214 (N_3214,N_3041,N_3058);
or U3215 (N_3215,N_3035,N_3047);
nand U3216 (N_3216,N_3078,N_3003);
and U3217 (N_3217,N_3118,N_3028);
nor U3218 (N_3218,N_3138,N_3063);
nor U3219 (N_3219,N_3111,N_3072);
nor U3220 (N_3220,N_3132,N_3076);
and U3221 (N_3221,N_3030,N_3143);
nand U3222 (N_3222,N_3024,N_3099);
and U3223 (N_3223,N_3108,N_3056);
or U3224 (N_3224,N_3060,N_3126);
nand U3225 (N_3225,N_3104,N_3078);
nor U3226 (N_3226,N_3092,N_3110);
nor U3227 (N_3227,N_3141,N_3134);
nand U3228 (N_3228,N_3127,N_3099);
and U3229 (N_3229,N_3054,N_3146);
nand U3230 (N_3230,N_3054,N_3143);
or U3231 (N_3231,N_3134,N_3051);
or U3232 (N_3232,N_3105,N_3141);
nand U3233 (N_3233,N_3061,N_3080);
or U3234 (N_3234,N_3033,N_3054);
or U3235 (N_3235,N_3101,N_3060);
nor U3236 (N_3236,N_3029,N_3051);
or U3237 (N_3237,N_3009,N_3007);
nor U3238 (N_3238,N_3142,N_3026);
nand U3239 (N_3239,N_3022,N_3018);
xnor U3240 (N_3240,N_3071,N_3100);
and U3241 (N_3241,N_3005,N_3039);
or U3242 (N_3242,N_3014,N_3141);
nor U3243 (N_3243,N_3130,N_3071);
nand U3244 (N_3244,N_3032,N_3083);
nand U3245 (N_3245,N_3105,N_3013);
nor U3246 (N_3246,N_3141,N_3122);
and U3247 (N_3247,N_3080,N_3143);
and U3248 (N_3248,N_3126,N_3008);
nor U3249 (N_3249,N_3117,N_3138);
nand U3250 (N_3250,N_3068,N_3144);
nor U3251 (N_3251,N_3015,N_3030);
and U3252 (N_3252,N_3037,N_3005);
xor U3253 (N_3253,N_3059,N_3145);
nand U3254 (N_3254,N_3064,N_3109);
nor U3255 (N_3255,N_3003,N_3048);
and U3256 (N_3256,N_3005,N_3093);
and U3257 (N_3257,N_3043,N_3006);
or U3258 (N_3258,N_3020,N_3137);
nand U3259 (N_3259,N_3147,N_3090);
and U3260 (N_3260,N_3070,N_3100);
xnor U3261 (N_3261,N_3010,N_3074);
nor U3262 (N_3262,N_3129,N_3038);
nand U3263 (N_3263,N_3122,N_3095);
and U3264 (N_3264,N_3049,N_3084);
nor U3265 (N_3265,N_3020,N_3110);
nand U3266 (N_3266,N_3011,N_3114);
and U3267 (N_3267,N_3145,N_3081);
nor U3268 (N_3268,N_3014,N_3076);
or U3269 (N_3269,N_3016,N_3004);
nand U3270 (N_3270,N_3122,N_3000);
nand U3271 (N_3271,N_3099,N_3043);
nand U3272 (N_3272,N_3080,N_3081);
nand U3273 (N_3273,N_3134,N_3052);
or U3274 (N_3274,N_3114,N_3095);
nand U3275 (N_3275,N_3136,N_3080);
and U3276 (N_3276,N_3146,N_3128);
nor U3277 (N_3277,N_3060,N_3080);
nand U3278 (N_3278,N_3110,N_3003);
or U3279 (N_3279,N_3074,N_3012);
or U3280 (N_3280,N_3003,N_3016);
nor U3281 (N_3281,N_3076,N_3022);
xnor U3282 (N_3282,N_3018,N_3057);
nand U3283 (N_3283,N_3013,N_3095);
nor U3284 (N_3284,N_3098,N_3135);
nand U3285 (N_3285,N_3042,N_3062);
nor U3286 (N_3286,N_3093,N_3081);
nand U3287 (N_3287,N_3005,N_3071);
and U3288 (N_3288,N_3122,N_3146);
nand U3289 (N_3289,N_3059,N_3013);
and U3290 (N_3290,N_3015,N_3142);
nand U3291 (N_3291,N_3108,N_3098);
and U3292 (N_3292,N_3117,N_3116);
and U3293 (N_3293,N_3124,N_3125);
xor U3294 (N_3294,N_3040,N_3014);
or U3295 (N_3295,N_3049,N_3107);
and U3296 (N_3296,N_3013,N_3010);
nand U3297 (N_3297,N_3056,N_3012);
and U3298 (N_3298,N_3036,N_3000);
and U3299 (N_3299,N_3077,N_3024);
and U3300 (N_3300,N_3165,N_3189);
or U3301 (N_3301,N_3282,N_3283);
xor U3302 (N_3302,N_3232,N_3218);
nand U3303 (N_3303,N_3276,N_3195);
or U3304 (N_3304,N_3216,N_3184);
and U3305 (N_3305,N_3272,N_3298);
nand U3306 (N_3306,N_3286,N_3220);
nor U3307 (N_3307,N_3243,N_3267);
xnor U3308 (N_3308,N_3200,N_3237);
nor U3309 (N_3309,N_3280,N_3211);
or U3310 (N_3310,N_3166,N_3169);
nor U3311 (N_3311,N_3222,N_3277);
nor U3312 (N_3312,N_3168,N_3201);
nor U3313 (N_3313,N_3246,N_3279);
xor U3314 (N_3314,N_3180,N_3265);
nor U3315 (N_3315,N_3238,N_3197);
or U3316 (N_3316,N_3186,N_3228);
nand U3317 (N_3317,N_3285,N_3212);
and U3318 (N_3318,N_3203,N_3198);
nand U3319 (N_3319,N_3163,N_3204);
nor U3320 (N_3320,N_3269,N_3288);
xor U3321 (N_3321,N_3260,N_3150);
and U3322 (N_3322,N_3161,N_3153);
xor U3323 (N_3323,N_3173,N_3236);
nor U3324 (N_3324,N_3241,N_3174);
xor U3325 (N_3325,N_3271,N_3281);
or U3326 (N_3326,N_3207,N_3188);
nand U3327 (N_3327,N_3217,N_3261);
or U3328 (N_3328,N_3176,N_3192);
nand U3329 (N_3329,N_3159,N_3299);
xnor U3330 (N_3330,N_3244,N_3291);
nor U3331 (N_3331,N_3177,N_3219);
nand U3332 (N_3332,N_3258,N_3160);
or U3333 (N_3333,N_3245,N_3182);
and U3334 (N_3334,N_3225,N_3259);
nand U3335 (N_3335,N_3294,N_3239);
nor U3336 (N_3336,N_3181,N_3226);
nor U3337 (N_3337,N_3205,N_3250);
nor U3338 (N_3338,N_3278,N_3234);
nor U3339 (N_3339,N_3156,N_3287);
nand U3340 (N_3340,N_3215,N_3202);
nand U3341 (N_3341,N_3268,N_3183);
nor U3342 (N_3342,N_3170,N_3297);
nand U3343 (N_3343,N_3175,N_3274);
xor U3344 (N_3344,N_3158,N_3249);
nand U3345 (N_3345,N_3263,N_3289);
xor U3346 (N_3346,N_3247,N_3157);
nor U3347 (N_3347,N_3206,N_3296);
or U3348 (N_3348,N_3185,N_3213);
and U3349 (N_3349,N_3248,N_3224);
or U3350 (N_3350,N_3209,N_3178);
nor U3351 (N_3351,N_3171,N_3151);
or U3352 (N_3352,N_3240,N_3164);
xnor U3353 (N_3353,N_3270,N_3293);
nor U3354 (N_3354,N_3242,N_3229);
nor U3355 (N_3355,N_3154,N_3167);
nand U3356 (N_3356,N_3155,N_3256);
xnor U3357 (N_3357,N_3196,N_3254);
nand U3358 (N_3358,N_3223,N_3266);
or U3359 (N_3359,N_3190,N_3199);
or U3360 (N_3360,N_3230,N_3253);
nand U3361 (N_3361,N_3193,N_3295);
and U3362 (N_3362,N_3252,N_3262);
or U3363 (N_3363,N_3257,N_3273);
or U3364 (N_3364,N_3264,N_3251);
or U3365 (N_3365,N_3194,N_3275);
and U3366 (N_3366,N_3191,N_3227);
or U3367 (N_3367,N_3233,N_3152);
and U3368 (N_3368,N_3221,N_3214);
nand U3369 (N_3369,N_3210,N_3284);
nand U3370 (N_3370,N_3162,N_3292);
or U3371 (N_3371,N_3208,N_3231);
xnor U3372 (N_3372,N_3235,N_3290);
nor U3373 (N_3373,N_3255,N_3179);
or U3374 (N_3374,N_3187,N_3172);
nor U3375 (N_3375,N_3266,N_3183);
nor U3376 (N_3376,N_3169,N_3202);
nor U3377 (N_3377,N_3204,N_3222);
xnor U3378 (N_3378,N_3296,N_3245);
nor U3379 (N_3379,N_3199,N_3257);
xnor U3380 (N_3380,N_3212,N_3190);
and U3381 (N_3381,N_3229,N_3174);
or U3382 (N_3382,N_3166,N_3175);
and U3383 (N_3383,N_3243,N_3265);
or U3384 (N_3384,N_3211,N_3162);
nor U3385 (N_3385,N_3233,N_3282);
nand U3386 (N_3386,N_3162,N_3204);
nor U3387 (N_3387,N_3261,N_3157);
nand U3388 (N_3388,N_3273,N_3253);
xnor U3389 (N_3389,N_3247,N_3238);
and U3390 (N_3390,N_3199,N_3181);
or U3391 (N_3391,N_3208,N_3182);
and U3392 (N_3392,N_3211,N_3242);
or U3393 (N_3393,N_3228,N_3174);
or U3394 (N_3394,N_3214,N_3275);
and U3395 (N_3395,N_3266,N_3257);
and U3396 (N_3396,N_3266,N_3249);
or U3397 (N_3397,N_3166,N_3230);
and U3398 (N_3398,N_3248,N_3263);
nor U3399 (N_3399,N_3233,N_3299);
nand U3400 (N_3400,N_3208,N_3256);
xnor U3401 (N_3401,N_3191,N_3152);
or U3402 (N_3402,N_3259,N_3294);
nor U3403 (N_3403,N_3150,N_3223);
and U3404 (N_3404,N_3253,N_3176);
nor U3405 (N_3405,N_3271,N_3221);
nor U3406 (N_3406,N_3254,N_3283);
and U3407 (N_3407,N_3282,N_3278);
or U3408 (N_3408,N_3191,N_3190);
nor U3409 (N_3409,N_3181,N_3197);
nand U3410 (N_3410,N_3269,N_3289);
or U3411 (N_3411,N_3173,N_3230);
nand U3412 (N_3412,N_3265,N_3257);
xor U3413 (N_3413,N_3159,N_3238);
and U3414 (N_3414,N_3212,N_3225);
and U3415 (N_3415,N_3243,N_3223);
nand U3416 (N_3416,N_3205,N_3200);
nor U3417 (N_3417,N_3168,N_3190);
nand U3418 (N_3418,N_3174,N_3219);
nand U3419 (N_3419,N_3257,N_3213);
and U3420 (N_3420,N_3189,N_3181);
nor U3421 (N_3421,N_3184,N_3235);
nor U3422 (N_3422,N_3231,N_3256);
nor U3423 (N_3423,N_3220,N_3245);
or U3424 (N_3424,N_3265,N_3198);
or U3425 (N_3425,N_3226,N_3252);
nand U3426 (N_3426,N_3248,N_3175);
nand U3427 (N_3427,N_3249,N_3160);
and U3428 (N_3428,N_3192,N_3239);
or U3429 (N_3429,N_3214,N_3285);
and U3430 (N_3430,N_3292,N_3179);
and U3431 (N_3431,N_3219,N_3216);
nand U3432 (N_3432,N_3210,N_3258);
nor U3433 (N_3433,N_3254,N_3217);
and U3434 (N_3434,N_3155,N_3203);
and U3435 (N_3435,N_3213,N_3276);
nor U3436 (N_3436,N_3267,N_3215);
nand U3437 (N_3437,N_3270,N_3273);
or U3438 (N_3438,N_3264,N_3172);
or U3439 (N_3439,N_3157,N_3297);
and U3440 (N_3440,N_3226,N_3228);
nand U3441 (N_3441,N_3171,N_3199);
and U3442 (N_3442,N_3225,N_3290);
nor U3443 (N_3443,N_3219,N_3180);
nand U3444 (N_3444,N_3234,N_3237);
and U3445 (N_3445,N_3219,N_3201);
nand U3446 (N_3446,N_3257,N_3264);
or U3447 (N_3447,N_3204,N_3259);
nor U3448 (N_3448,N_3253,N_3159);
nor U3449 (N_3449,N_3272,N_3167);
or U3450 (N_3450,N_3337,N_3325);
nor U3451 (N_3451,N_3367,N_3362);
nand U3452 (N_3452,N_3370,N_3369);
and U3453 (N_3453,N_3445,N_3322);
nand U3454 (N_3454,N_3351,N_3449);
or U3455 (N_3455,N_3341,N_3411);
nand U3456 (N_3456,N_3408,N_3430);
xor U3457 (N_3457,N_3318,N_3311);
nor U3458 (N_3458,N_3349,N_3344);
nand U3459 (N_3459,N_3397,N_3359);
nand U3460 (N_3460,N_3394,N_3429);
and U3461 (N_3461,N_3320,N_3372);
xnor U3462 (N_3462,N_3352,N_3390);
xor U3463 (N_3463,N_3376,N_3331);
or U3464 (N_3464,N_3401,N_3439);
nand U3465 (N_3465,N_3317,N_3353);
and U3466 (N_3466,N_3398,N_3332);
xnor U3467 (N_3467,N_3319,N_3307);
or U3468 (N_3468,N_3315,N_3312);
nand U3469 (N_3469,N_3304,N_3305);
xnor U3470 (N_3470,N_3327,N_3378);
and U3471 (N_3471,N_3436,N_3385);
and U3472 (N_3472,N_3358,N_3404);
and U3473 (N_3473,N_3392,N_3361);
or U3474 (N_3474,N_3314,N_3406);
nor U3475 (N_3475,N_3323,N_3448);
xnor U3476 (N_3476,N_3381,N_3432);
and U3477 (N_3477,N_3442,N_3321);
nand U3478 (N_3478,N_3384,N_3306);
or U3479 (N_3479,N_3380,N_3402);
or U3480 (N_3480,N_3389,N_3375);
nand U3481 (N_3481,N_3419,N_3386);
nor U3482 (N_3482,N_3328,N_3382);
nor U3483 (N_3483,N_3363,N_3330);
and U3484 (N_3484,N_3340,N_3405);
xnor U3485 (N_3485,N_3308,N_3422);
nor U3486 (N_3486,N_3447,N_3391);
xnor U3487 (N_3487,N_3440,N_3377);
or U3488 (N_3488,N_3357,N_3410);
nor U3489 (N_3489,N_3427,N_3425);
or U3490 (N_3490,N_3399,N_3443);
and U3491 (N_3491,N_3407,N_3444);
nor U3492 (N_3492,N_3409,N_3379);
and U3493 (N_3493,N_3438,N_3415);
or U3494 (N_3494,N_3336,N_3424);
xor U3495 (N_3495,N_3310,N_3413);
or U3496 (N_3496,N_3368,N_3302);
nor U3497 (N_3497,N_3396,N_3326);
or U3498 (N_3498,N_3416,N_3338);
or U3499 (N_3499,N_3324,N_3366);
xor U3500 (N_3500,N_3435,N_3346);
nor U3501 (N_3501,N_3423,N_3301);
or U3502 (N_3502,N_3309,N_3335);
and U3503 (N_3503,N_3329,N_3342);
or U3504 (N_3504,N_3371,N_3356);
and U3505 (N_3505,N_3365,N_3426);
nor U3506 (N_3506,N_3313,N_3428);
and U3507 (N_3507,N_3420,N_3339);
or U3508 (N_3508,N_3414,N_3350);
and U3509 (N_3509,N_3403,N_3374);
nand U3510 (N_3510,N_3418,N_3434);
and U3511 (N_3511,N_3383,N_3433);
and U3512 (N_3512,N_3421,N_3417);
and U3513 (N_3513,N_3347,N_3303);
or U3514 (N_3514,N_3373,N_3388);
nor U3515 (N_3515,N_3431,N_3300);
nor U3516 (N_3516,N_3441,N_3354);
nor U3517 (N_3517,N_3437,N_3393);
or U3518 (N_3518,N_3400,N_3343);
or U3519 (N_3519,N_3364,N_3334);
nand U3520 (N_3520,N_3345,N_3395);
or U3521 (N_3521,N_3355,N_3446);
or U3522 (N_3522,N_3360,N_3316);
nand U3523 (N_3523,N_3333,N_3387);
and U3524 (N_3524,N_3348,N_3412);
or U3525 (N_3525,N_3447,N_3326);
nor U3526 (N_3526,N_3335,N_3322);
and U3527 (N_3527,N_3443,N_3340);
nor U3528 (N_3528,N_3433,N_3359);
or U3529 (N_3529,N_3336,N_3318);
nor U3530 (N_3530,N_3313,N_3342);
and U3531 (N_3531,N_3438,N_3375);
or U3532 (N_3532,N_3368,N_3348);
nand U3533 (N_3533,N_3347,N_3389);
and U3534 (N_3534,N_3371,N_3398);
and U3535 (N_3535,N_3304,N_3361);
and U3536 (N_3536,N_3431,N_3390);
nor U3537 (N_3537,N_3385,N_3307);
or U3538 (N_3538,N_3403,N_3439);
nor U3539 (N_3539,N_3443,N_3314);
nor U3540 (N_3540,N_3323,N_3328);
and U3541 (N_3541,N_3319,N_3406);
nor U3542 (N_3542,N_3347,N_3349);
nand U3543 (N_3543,N_3435,N_3393);
or U3544 (N_3544,N_3315,N_3446);
nand U3545 (N_3545,N_3307,N_3369);
nand U3546 (N_3546,N_3320,N_3406);
or U3547 (N_3547,N_3364,N_3439);
or U3548 (N_3548,N_3449,N_3303);
nor U3549 (N_3549,N_3420,N_3436);
nand U3550 (N_3550,N_3349,N_3307);
or U3551 (N_3551,N_3405,N_3413);
and U3552 (N_3552,N_3396,N_3422);
and U3553 (N_3553,N_3367,N_3424);
nand U3554 (N_3554,N_3412,N_3408);
or U3555 (N_3555,N_3353,N_3432);
nand U3556 (N_3556,N_3393,N_3438);
nor U3557 (N_3557,N_3362,N_3438);
or U3558 (N_3558,N_3346,N_3320);
and U3559 (N_3559,N_3444,N_3441);
nor U3560 (N_3560,N_3376,N_3336);
or U3561 (N_3561,N_3397,N_3374);
nand U3562 (N_3562,N_3372,N_3352);
or U3563 (N_3563,N_3377,N_3411);
or U3564 (N_3564,N_3387,N_3348);
nand U3565 (N_3565,N_3340,N_3364);
nor U3566 (N_3566,N_3363,N_3382);
nand U3567 (N_3567,N_3433,N_3337);
xnor U3568 (N_3568,N_3376,N_3320);
and U3569 (N_3569,N_3374,N_3445);
and U3570 (N_3570,N_3381,N_3412);
or U3571 (N_3571,N_3337,N_3432);
or U3572 (N_3572,N_3448,N_3441);
nand U3573 (N_3573,N_3432,N_3358);
or U3574 (N_3574,N_3448,N_3449);
xor U3575 (N_3575,N_3366,N_3357);
xnor U3576 (N_3576,N_3352,N_3378);
nor U3577 (N_3577,N_3389,N_3349);
or U3578 (N_3578,N_3366,N_3423);
nor U3579 (N_3579,N_3378,N_3434);
nand U3580 (N_3580,N_3302,N_3421);
or U3581 (N_3581,N_3305,N_3365);
and U3582 (N_3582,N_3404,N_3375);
and U3583 (N_3583,N_3326,N_3370);
xnor U3584 (N_3584,N_3389,N_3340);
xnor U3585 (N_3585,N_3375,N_3434);
nor U3586 (N_3586,N_3302,N_3304);
nand U3587 (N_3587,N_3350,N_3371);
nand U3588 (N_3588,N_3323,N_3345);
or U3589 (N_3589,N_3368,N_3363);
or U3590 (N_3590,N_3338,N_3383);
or U3591 (N_3591,N_3321,N_3312);
nand U3592 (N_3592,N_3432,N_3433);
nor U3593 (N_3593,N_3303,N_3417);
and U3594 (N_3594,N_3435,N_3437);
nor U3595 (N_3595,N_3432,N_3386);
nor U3596 (N_3596,N_3440,N_3411);
nand U3597 (N_3597,N_3371,N_3347);
nor U3598 (N_3598,N_3313,N_3386);
or U3599 (N_3599,N_3388,N_3328);
nor U3600 (N_3600,N_3566,N_3461);
nor U3601 (N_3601,N_3578,N_3509);
xnor U3602 (N_3602,N_3507,N_3465);
or U3603 (N_3603,N_3551,N_3592);
xnor U3604 (N_3604,N_3453,N_3534);
nand U3605 (N_3605,N_3458,N_3575);
nand U3606 (N_3606,N_3524,N_3472);
nand U3607 (N_3607,N_3496,N_3519);
nor U3608 (N_3608,N_3469,N_3552);
or U3609 (N_3609,N_3466,N_3544);
or U3610 (N_3610,N_3591,N_3506);
nor U3611 (N_3611,N_3484,N_3573);
nor U3612 (N_3612,N_3590,N_3515);
and U3613 (N_3613,N_3473,N_3588);
or U3614 (N_3614,N_3530,N_3565);
nand U3615 (N_3615,N_3512,N_3491);
nor U3616 (N_3616,N_3475,N_3579);
or U3617 (N_3617,N_3486,N_3584);
nor U3618 (N_3618,N_3563,N_3554);
or U3619 (N_3619,N_3589,N_3535);
nor U3620 (N_3620,N_3489,N_3559);
xnor U3621 (N_3621,N_3558,N_3593);
or U3622 (N_3622,N_3479,N_3474);
and U3623 (N_3623,N_3570,N_3586);
and U3624 (N_3624,N_3462,N_3543);
and U3625 (N_3625,N_3504,N_3490);
xor U3626 (N_3626,N_3511,N_3582);
nor U3627 (N_3627,N_3599,N_3545);
nand U3628 (N_3628,N_3594,N_3540);
or U3629 (N_3629,N_3485,N_3457);
and U3630 (N_3630,N_3541,N_3546);
or U3631 (N_3631,N_3569,N_3539);
and U3632 (N_3632,N_3517,N_3567);
nor U3633 (N_3633,N_3527,N_3574);
and U3634 (N_3634,N_3580,N_3495);
nand U3635 (N_3635,N_3464,N_3556);
or U3636 (N_3636,N_3502,N_3467);
nor U3637 (N_3637,N_3459,N_3454);
nor U3638 (N_3638,N_3503,N_3493);
nand U3639 (N_3639,N_3487,N_3576);
and U3640 (N_3640,N_3568,N_3518);
nand U3641 (N_3641,N_3482,N_3450);
or U3642 (N_3642,N_3499,N_3585);
nand U3643 (N_3643,N_3596,N_3510);
nand U3644 (N_3644,N_3505,N_3581);
nand U3645 (N_3645,N_3494,N_3549);
and U3646 (N_3646,N_3597,N_3532);
nor U3647 (N_3647,N_3553,N_3480);
or U3648 (N_3648,N_3478,N_3555);
nand U3649 (N_3649,N_3587,N_3526);
xor U3650 (N_3650,N_3561,N_3477);
nand U3651 (N_3651,N_3521,N_3520);
nand U3652 (N_3652,N_3476,N_3531);
xnor U3653 (N_3653,N_3572,N_3488);
nor U3654 (N_3654,N_3548,N_3451);
nand U3655 (N_3655,N_3455,N_3481);
nand U3656 (N_3656,N_3571,N_3523);
nand U3657 (N_3657,N_3557,N_3468);
and U3658 (N_3658,N_3560,N_3497);
nor U3659 (N_3659,N_3528,N_3483);
nand U3660 (N_3660,N_3470,N_3547);
or U3661 (N_3661,N_3562,N_3529);
xor U3662 (N_3662,N_3564,N_3452);
nor U3663 (N_3663,N_3513,N_3522);
nand U3664 (N_3664,N_3460,N_3598);
or U3665 (N_3665,N_3583,N_3492);
and U3666 (N_3666,N_3536,N_3514);
or U3667 (N_3667,N_3508,N_3498);
nor U3668 (N_3668,N_3456,N_3471);
or U3669 (N_3669,N_3577,N_3500);
and U3670 (N_3670,N_3525,N_3550);
and U3671 (N_3671,N_3516,N_3538);
or U3672 (N_3672,N_3533,N_3537);
and U3673 (N_3673,N_3501,N_3595);
and U3674 (N_3674,N_3463,N_3542);
nand U3675 (N_3675,N_3466,N_3594);
nand U3676 (N_3676,N_3507,N_3514);
nor U3677 (N_3677,N_3454,N_3465);
nand U3678 (N_3678,N_3541,N_3518);
and U3679 (N_3679,N_3476,N_3545);
or U3680 (N_3680,N_3452,N_3517);
nand U3681 (N_3681,N_3544,N_3519);
and U3682 (N_3682,N_3501,N_3586);
or U3683 (N_3683,N_3464,N_3490);
nor U3684 (N_3684,N_3527,N_3504);
nand U3685 (N_3685,N_3467,N_3460);
or U3686 (N_3686,N_3465,N_3587);
and U3687 (N_3687,N_3545,N_3520);
nand U3688 (N_3688,N_3583,N_3455);
nor U3689 (N_3689,N_3563,N_3574);
or U3690 (N_3690,N_3533,N_3597);
nand U3691 (N_3691,N_3541,N_3462);
nor U3692 (N_3692,N_3531,N_3574);
or U3693 (N_3693,N_3581,N_3488);
nor U3694 (N_3694,N_3460,N_3457);
or U3695 (N_3695,N_3459,N_3554);
nand U3696 (N_3696,N_3465,N_3496);
and U3697 (N_3697,N_3550,N_3522);
nand U3698 (N_3698,N_3467,N_3515);
and U3699 (N_3699,N_3557,N_3550);
or U3700 (N_3700,N_3489,N_3517);
nand U3701 (N_3701,N_3486,N_3502);
or U3702 (N_3702,N_3452,N_3516);
and U3703 (N_3703,N_3461,N_3560);
nand U3704 (N_3704,N_3563,N_3551);
or U3705 (N_3705,N_3488,N_3525);
and U3706 (N_3706,N_3573,N_3558);
nor U3707 (N_3707,N_3534,N_3478);
and U3708 (N_3708,N_3594,N_3475);
xnor U3709 (N_3709,N_3537,N_3577);
or U3710 (N_3710,N_3576,N_3515);
nand U3711 (N_3711,N_3579,N_3479);
or U3712 (N_3712,N_3533,N_3455);
and U3713 (N_3713,N_3482,N_3580);
nand U3714 (N_3714,N_3588,N_3534);
or U3715 (N_3715,N_3516,N_3460);
nor U3716 (N_3716,N_3583,N_3472);
nand U3717 (N_3717,N_3467,N_3523);
or U3718 (N_3718,N_3577,N_3475);
or U3719 (N_3719,N_3531,N_3560);
nand U3720 (N_3720,N_3516,N_3553);
nand U3721 (N_3721,N_3495,N_3561);
nand U3722 (N_3722,N_3583,N_3550);
xor U3723 (N_3723,N_3477,N_3588);
or U3724 (N_3724,N_3450,N_3545);
xnor U3725 (N_3725,N_3595,N_3506);
nor U3726 (N_3726,N_3474,N_3524);
xnor U3727 (N_3727,N_3558,N_3565);
nand U3728 (N_3728,N_3491,N_3470);
or U3729 (N_3729,N_3505,N_3478);
and U3730 (N_3730,N_3558,N_3542);
nand U3731 (N_3731,N_3494,N_3513);
nor U3732 (N_3732,N_3471,N_3564);
xnor U3733 (N_3733,N_3570,N_3459);
nand U3734 (N_3734,N_3510,N_3563);
xor U3735 (N_3735,N_3599,N_3456);
or U3736 (N_3736,N_3595,N_3528);
or U3737 (N_3737,N_3514,N_3504);
nor U3738 (N_3738,N_3553,N_3483);
nor U3739 (N_3739,N_3516,N_3563);
nor U3740 (N_3740,N_3480,N_3556);
nor U3741 (N_3741,N_3507,N_3451);
nand U3742 (N_3742,N_3569,N_3574);
or U3743 (N_3743,N_3468,N_3550);
and U3744 (N_3744,N_3491,N_3481);
and U3745 (N_3745,N_3479,N_3569);
xor U3746 (N_3746,N_3587,N_3571);
nand U3747 (N_3747,N_3483,N_3456);
nand U3748 (N_3748,N_3561,N_3546);
or U3749 (N_3749,N_3588,N_3505);
or U3750 (N_3750,N_3664,N_3603);
and U3751 (N_3751,N_3711,N_3741);
and U3752 (N_3752,N_3702,N_3635);
or U3753 (N_3753,N_3642,N_3615);
or U3754 (N_3754,N_3637,N_3652);
or U3755 (N_3755,N_3728,N_3611);
and U3756 (N_3756,N_3659,N_3641);
and U3757 (N_3757,N_3684,N_3678);
nand U3758 (N_3758,N_3723,N_3616);
nor U3759 (N_3759,N_3651,N_3739);
and U3760 (N_3760,N_3688,N_3634);
and U3761 (N_3761,N_3705,N_3640);
nand U3762 (N_3762,N_3618,N_3690);
and U3763 (N_3763,N_3709,N_3719);
nand U3764 (N_3764,N_3696,N_3631);
nor U3765 (N_3765,N_3667,N_3692);
nand U3766 (N_3766,N_3710,N_3748);
nand U3767 (N_3767,N_3645,N_3636);
nand U3768 (N_3768,N_3715,N_3729);
or U3769 (N_3769,N_3689,N_3726);
nand U3770 (N_3770,N_3614,N_3621);
nand U3771 (N_3771,N_3721,N_3620);
or U3772 (N_3772,N_3745,N_3676);
or U3773 (N_3773,N_3720,N_3607);
or U3774 (N_3774,N_3675,N_3627);
or U3775 (N_3775,N_3732,N_3663);
and U3776 (N_3776,N_3612,N_3712);
or U3777 (N_3777,N_3630,N_3648);
and U3778 (N_3778,N_3738,N_3632);
or U3779 (N_3779,N_3646,N_3628);
or U3780 (N_3780,N_3613,N_3695);
or U3781 (N_3781,N_3622,N_3656);
and U3782 (N_3782,N_3691,N_3647);
and U3783 (N_3783,N_3682,N_3703);
nor U3784 (N_3784,N_3670,N_3734);
nor U3785 (N_3785,N_3725,N_3626);
nor U3786 (N_3786,N_3743,N_3742);
nor U3787 (N_3787,N_3669,N_3671);
xor U3788 (N_3788,N_3673,N_3713);
or U3789 (N_3789,N_3624,N_3658);
nand U3790 (N_3790,N_3707,N_3665);
nand U3791 (N_3791,N_3608,N_3714);
or U3792 (N_3792,N_3685,N_3638);
or U3793 (N_3793,N_3724,N_3700);
or U3794 (N_3794,N_3649,N_3683);
nor U3795 (N_3795,N_3679,N_3644);
xnor U3796 (N_3796,N_3746,N_3668);
xnor U3797 (N_3797,N_3602,N_3605);
nand U3798 (N_3798,N_3727,N_3699);
or U3799 (N_3799,N_3657,N_3701);
and U3800 (N_3800,N_3660,N_3693);
and U3801 (N_3801,N_3749,N_3672);
and U3802 (N_3802,N_3650,N_3731);
nand U3803 (N_3803,N_3604,N_3609);
nand U3804 (N_3804,N_3680,N_3600);
and U3805 (N_3805,N_3661,N_3643);
and U3806 (N_3806,N_3736,N_3718);
xor U3807 (N_3807,N_3735,N_3706);
nor U3808 (N_3808,N_3617,N_3677);
nand U3809 (N_3809,N_3606,N_3653);
nor U3810 (N_3810,N_3623,N_3740);
or U3811 (N_3811,N_3733,N_3674);
or U3812 (N_3812,N_3601,N_3629);
nand U3813 (N_3813,N_3654,N_3666);
nor U3814 (N_3814,N_3747,N_3730);
xnor U3815 (N_3815,N_3610,N_3697);
and U3816 (N_3816,N_3716,N_3708);
or U3817 (N_3817,N_3619,N_3704);
and U3818 (N_3818,N_3722,N_3744);
nand U3819 (N_3819,N_3639,N_3686);
or U3820 (N_3820,N_3694,N_3662);
or U3821 (N_3821,N_3717,N_3698);
nor U3822 (N_3822,N_3633,N_3655);
nand U3823 (N_3823,N_3681,N_3687);
and U3824 (N_3824,N_3737,N_3625);
and U3825 (N_3825,N_3710,N_3656);
nor U3826 (N_3826,N_3732,N_3643);
nor U3827 (N_3827,N_3732,N_3624);
and U3828 (N_3828,N_3646,N_3626);
and U3829 (N_3829,N_3693,N_3663);
or U3830 (N_3830,N_3685,N_3645);
or U3831 (N_3831,N_3743,N_3629);
nand U3832 (N_3832,N_3636,N_3648);
xnor U3833 (N_3833,N_3616,N_3649);
nand U3834 (N_3834,N_3615,N_3669);
nand U3835 (N_3835,N_3632,N_3605);
xnor U3836 (N_3836,N_3604,N_3710);
and U3837 (N_3837,N_3730,N_3709);
xnor U3838 (N_3838,N_3682,N_3653);
nand U3839 (N_3839,N_3602,N_3713);
or U3840 (N_3840,N_3617,N_3654);
or U3841 (N_3841,N_3610,N_3731);
and U3842 (N_3842,N_3690,N_3643);
nand U3843 (N_3843,N_3652,N_3635);
and U3844 (N_3844,N_3646,N_3742);
nor U3845 (N_3845,N_3694,N_3603);
and U3846 (N_3846,N_3677,N_3700);
nor U3847 (N_3847,N_3685,N_3615);
or U3848 (N_3848,N_3699,N_3673);
or U3849 (N_3849,N_3715,N_3634);
nand U3850 (N_3850,N_3713,N_3733);
or U3851 (N_3851,N_3615,N_3706);
or U3852 (N_3852,N_3653,N_3735);
nand U3853 (N_3853,N_3644,N_3621);
and U3854 (N_3854,N_3607,N_3672);
or U3855 (N_3855,N_3655,N_3682);
or U3856 (N_3856,N_3663,N_3679);
nand U3857 (N_3857,N_3624,N_3638);
or U3858 (N_3858,N_3743,N_3604);
nand U3859 (N_3859,N_3749,N_3698);
nor U3860 (N_3860,N_3630,N_3663);
nor U3861 (N_3861,N_3634,N_3723);
nor U3862 (N_3862,N_3666,N_3728);
nand U3863 (N_3863,N_3652,N_3684);
or U3864 (N_3864,N_3718,N_3623);
nand U3865 (N_3865,N_3703,N_3685);
and U3866 (N_3866,N_3737,N_3652);
or U3867 (N_3867,N_3685,N_3668);
or U3868 (N_3868,N_3748,N_3749);
xnor U3869 (N_3869,N_3636,N_3606);
nor U3870 (N_3870,N_3721,N_3686);
or U3871 (N_3871,N_3668,N_3712);
or U3872 (N_3872,N_3653,N_3691);
xnor U3873 (N_3873,N_3665,N_3734);
and U3874 (N_3874,N_3667,N_3725);
and U3875 (N_3875,N_3668,N_3682);
and U3876 (N_3876,N_3741,N_3729);
and U3877 (N_3877,N_3679,N_3658);
and U3878 (N_3878,N_3746,N_3661);
and U3879 (N_3879,N_3673,N_3730);
nor U3880 (N_3880,N_3642,N_3641);
nor U3881 (N_3881,N_3749,N_3652);
or U3882 (N_3882,N_3635,N_3726);
nor U3883 (N_3883,N_3634,N_3700);
nand U3884 (N_3884,N_3741,N_3665);
nor U3885 (N_3885,N_3696,N_3613);
or U3886 (N_3886,N_3704,N_3749);
and U3887 (N_3887,N_3649,N_3669);
and U3888 (N_3888,N_3644,N_3629);
nor U3889 (N_3889,N_3691,N_3655);
or U3890 (N_3890,N_3607,N_3719);
and U3891 (N_3891,N_3637,N_3671);
nor U3892 (N_3892,N_3727,N_3684);
nand U3893 (N_3893,N_3669,N_3628);
nor U3894 (N_3894,N_3657,N_3720);
nor U3895 (N_3895,N_3700,N_3664);
or U3896 (N_3896,N_3749,N_3709);
or U3897 (N_3897,N_3681,N_3677);
nor U3898 (N_3898,N_3671,N_3689);
nor U3899 (N_3899,N_3639,N_3625);
and U3900 (N_3900,N_3790,N_3769);
nor U3901 (N_3901,N_3801,N_3810);
nand U3902 (N_3902,N_3885,N_3827);
nor U3903 (N_3903,N_3891,N_3857);
nand U3904 (N_3904,N_3830,N_3869);
nand U3905 (N_3905,N_3836,N_3837);
and U3906 (N_3906,N_3792,N_3754);
nor U3907 (N_3907,N_3757,N_3751);
nand U3908 (N_3908,N_3785,N_3862);
or U3909 (N_3909,N_3794,N_3791);
xnor U3910 (N_3910,N_3882,N_3838);
nor U3911 (N_3911,N_3855,N_3848);
and U3912 (N_3912,N_3826,N_3783);
nor U3913 (N_3913,N_3880,N_3883);
or U3914 (N_3914,N_3818,N_3820);
nor U3915 (N_3915,N_3780,N_3898);
or U3916 (N_3916,N_3773,N_3888);
nand U3917 (N_3917,N_3872,N_3860);
nand U3918 (N_3918,N_3849,N_3805);
nand U3919 (N_3919,N_3853,N_3841);
nand U3920 (N_3920,N_3845,N_3859);
or U3921 (N_3921,N_3789,N_3798);
or U3922 (N_3922,N_3894,N_3868);
or U3923 (N_3923,N_3835,N_3847);
nand U3924 (N_3924,N_3759,N_3824);
nor U3925 (N_3925,N_3866,N_3800);
nand U3926 (N_3926,N_3776,N_3778);
or U3927 (N_3927,N_3832,N_3750);
or U3928 (N_3928,N_3877,N_3889);
or U3929 (N_3929,N_3875,N_3846);
or U3930 (N_3930,N_3899,N_3772);
or U3931 (N_3931,N_3895,N_3807);
or U3932 (N_3932,N_3756,N_3804);
and U3933 (N_3933,N_3850,N_3814);
nand U3934 (N_3934,N_3758,N_3799);
nand U3935 (N_3935,N_3768,N_3808);
nor U3936 (N_3936,N_3890,N_3876);
nand U3937 (N_3937,N_3802,N_3788);
nor U3938 (N_3938,N_3839,N_3755);
or U3939 (N_3939,N_3881,N_3787);
or U3940 (N_3940,N_3821,N_3886);
and U3941 (N_3941,N_3809,N_3828);
nor U3942 (N_3942,N_3873,N_3797);
nor U3943 (N_3943,N_3829,N_3834);
or U3944 (N_3944,N_3817,N_3842);
nor U3945 (N_3945,N_3867,N_3763);
or U3946 (N_3946,N_3812,N_3851);
nor U3947 (N_3947,N_3852,N_3833);
nor U3948 (N_3948,N_3753,N_3840);
or U3949 (N_3949,N_3878,N_3843);
and U3950 (N_3950,N_3854,N_3771);
nor U3951 (N_3951,N_3865,N_3892);
nand U3952 (N_3952,N_3779,N_3825);
nor U3953 (N_3953,N_3871,N_3806);
xnor U3954 (N_3954,N_3861,N_3765);
nor U3955 (N_3955,N_3796,N_3815);
or U3956 (N_3956,N_3856,N_3781);
nor U3957 (N_3957,N_3864,N_3884);
nand U3958 (N_3958,N_3803,N_3760);
and U3959 (N_3959,N_3887,N_3816);
and U3960 (N_3960,N_3897,N_3858);
nor U3961 (N_3961,N_3822,N_3764);
or U3962 (N_3962,N_3793,N_3766);
nand U3963 (N_3963,N_3896,N_3811);
nand U3964 (N_3964,N_3863,N_3870);
nand U3965 (N_3965,N_3844,N_3774);
or U3966 (N_3966,N_3752,N_3831);
xnor U3967 (N_3967,N_3770,N_3775);
nor U3968 (N_3968,N_3777,N_3795);
and U3969 (N_3969,N_3874,N_3819);
and U3970 (N_3970,N_3761,N_3879);
nand U3971 (N_3971,N_3767,N_3782);
nand U3972 (N_3972,N_3823,N_3813);
or U3973 (N_3973,N_3786,N_3784);
nand U3974 (N_3974,N_3893,N_3762);
nand U3975 (N_3975,N_3785,N_3884);
nand U3976 (N_3976,N_3770,N_3815);
xnor U3977 (N_3977,N_3859,N_3813);
or U3978 (N_3978,N_3754,N_3855);
or U3979 (N_3979,N_3866,N_3897);
nor U3980 (N_3980,N_3834,N_3789);
xor U3981 (N_3981,N_3831,N_3777);
nand U3982 (N_3982,N_3827,N_3779);
or U3983 (N_3983,N_3812,N_3784);
xor U3984 (N_3984,N_3869,N_3845);
nand U3985 (N_3985,N_3754,N_3883);
or U3986 (N_3986,N_3895,N_3894);
nand U3987 (N_3987,N_3778,N_3856);
nand U3988 (N_3988,N_3830,N_3813);
xor U3989 (N_3989,N_3792,N_3871);
and U3990 (N_3990,N_3850,N_3815);
nand U3991 (N_3991,N_3864,N_3856);
and U3992 (N_3992,N_3858,N_3809);
and U3993 (N_3993,N_3776,N_3768);
and U3994 (N_3994,N_3813,N_3795);
or U3995 (N_3995,N_3804,N_3878);
nor U3996 (N_3996,N_3884,N_3874);
or U3997 (N_3997,N_3795,N_3847);
and U3998 (N_3998,N_3882,N_3830);
or U3999 (N_3999,N_3873,N_3884);
and U4000 (N_4000,N_3844,N_3833);
and U4001 (N_4001,N_3875,N_3849);
or U4002 (N_4002,N_3752,N_3767);
nand U4003 (N_4003,N_3813,N_3774);
and U4004 (N_4004,N_3798,N_3863);
nand U4005 (N_4005,N_3759,N_3889);
or U4006 (N_4006,N_3848,N_3779);
nor U4007 (N_4007,N_3896,N_3822);
or U4008 (N_4008,N_3865,N_3773);
nor U4009 (N_4009,N_3785,N_3818);
xnor U4010 (N_4010,N_3792,N_3825);
and U4011 (N_4011,N_3826,N_3789);
xor U4012 (N_4012,N_3870,N_3796);
xor U4013 (N_4013,N_3860,N_3883);
or U4014 (N_4014,N_3773,N_3884);
or U4015 (N_4015,N_3854,N_3849);
and U4016 (N_4016,N_3776,N_3775);
nor U4017 (N_4017,N_3782,N_3779);
nor U4018 (N_4018,N_3885,N_3842);
xnor U4019 (N_4019,N_3875,N_3804);
nand U4020 (N_4020,N_3864,N_3783);
or U4021 (N_4021,N_3774,N_3885);
or U4022 (N_4022,N_3826,N_3780);
or U4023 (N_4023,N_3840,N_3770);
xnor U4024 (N_4024,N_3895,N_3827);
nand U4025 (N_4025,N_3773,N_3886);
nand U4026 (N_4026,N_3753,N_3791);
nor U4027 (N_4027,N_3813,N_3757);
and U4028 (N_4028,N_3851,N_3829);
or U4029 (N_4029,N_3785,N_3845);
nand U4030 (N_4030,N_3898,N_3865);
or U4031 (N_4031,N_3815,N_3804);
nor U4032 (N_4032,N_3871,N_3767);
or U4033 (N_4033,N_3802,N_3830);
nand U4034 (N_4034,N_3887,N_3790);
nor U4035 (N_4035,N_3889,N_3825);
nand U4036 (N_4036,N_3879,N_3790);
xor U4037 (N_4037,N_3854,N_3800);
nand U4038 (N_4038,N_3836,N_3786);
or U4039 (N_4039,N_3843,N_3867);
nand U4040 (N_4040,N_3883,N_3791);
nor U4041 (N_4041,N_3866,N_3810);
nor U4042 (N_4042,N_3765,N_3841);
nand U4043 (N_4043,N_3831,N_3820);
and U4044 (N_4044,N_3874,N_3826);
and U4045 (N_4045,N_3852,N_3786);
and U4046 (N_4046,N_3790,N_3811);
nor U4047 (N_4047,N_3778,N_3785);
nand U4048 (N_4048,N_3831,N_3880);
and U4049 (N_4049,N_3844,N_3836);
nand U4050 (N_4050,N_3988,N_4018);
nand U4051 (N_4051,N_3919,N_3991);
or U4052 (N_4052,N_3920,N_3926);
or U4053 (N_4053,N_3904,N_3948);
nor U4054 (N_4054,N_3933,N_3918);
or U4055 (N_4055,N_4032,N_3974);
xnor U4056 (N_4056,N_3987,N_3978);
or U4057 (N_4057,N_3911,N_3983);
nand U4058 (N_4058,N_4036,N_4038);
nand U4059 (N_4059,N_4002,N_3962);
and U4060 (N_4060,N_4049,N_3947);
or U4061 (N_4061,N_3992,N_3909);
nor U4062 (N_4062,N_3964,N_3939);
and U4063 (N_4063,N_3903,N_4016);
or U4064 (N_4064,N_4001,N_3938);
nand U4065 (N_4065,N_3967,N_3950);
and U4066 (N_4066,N_3996,N_3968);
nor U4067 (N_4067,N_4014,N_4029);
or U4068 (N_4068,N_4043,N_4004);
nand U4069 (N_4069,N_3913,N_3972);
nor U4070 (N_4070,N_3940,N_3901);
and U4071 (N_4071,N_3954,N_4047);
and U4072 (N_4072,N_4000,N_3998);
xor U4073 (N_4073,N_4012,N_4008);
nand U4074 (N_4074,N_4003,N_3980);
nand U4075 (N_4075,N_3923,N_3941);
nand U4076 (N_4076,N_3921,N_3994);
and U4077 (N_4077,N_3961,N_3986);
or U4078 (N_4078,N_3955,N_3984);
and U4079 (N_4079,N_3975,N_3970);
and U4080 (N_4080,N_3990,N_3957);
nor U4081 (N_4081,N_3971,N_3902);
nor U4082 (N_4082,N_3952,N_3932);
or U4083 (N_4083,N_4048,N_4041);
xnor U4084 (N_4084,N_3965,N_4044);
and U4085 (N_4085,N_3929,N_3956);
and U4086 (N_4086,N_3944,N_3949);
or U4087 (N_4087,N_3908,N_4034);
nor U4088 (N_4088,N_4030,N_4020);
nor U4089 (N_4089,N_3973,N_3900);
nand U4090 (N_4090,N_4007,N_4035);
xor U4091 (N_4091,N_4010,N_4006);
and U4092 (N_4092,N_3931,N_3942);
and U4093 (N_4093,N_4031,N_4037);
or U4094 (N_4094,N_3930,N_4022);
nor U4095 (N_4095,N_3985,N_3922);
and U4096 (N_4096,N_4040,N_3906);
xor U4097 (N_4097,N_4017,N_3916);
nor U4098 (N_4098,N_3979,N_4024);
nand U4099 (N_4099,N_3915,N_3914);
nand U4100 (N_4100,N_4028,N_3912);
and U4101 (N_4101,N_4027,N_3917);
and U4102 (N_4102,N_3927,N_4009);
nand U4103 (N_4103,N_3907,N_3905);
and U4104 (N_4104,N_4042,N_3959);
nand U4105 (N_4105,N_4045,N_3989);
and U4106 (N_4106,N_3936,N_3946);
nand U4107 (N_4107,N_3910,N_4013);
nor U4108 (N_4108,N_3945,N_4039);
and U4109 (N_4109,N_3963,N_3999);
and U4110 (N_4110,N_3997,N_4046);
or U4111 (N_4111,N_4023,N_4033);
nand U4112 (N_4112,N_4019,N_3935);
nor U4113 (N_4113,N_3976,N_3934);
nand U4114 (N_4114,N_4021,N_3928);
or U4115 (N_4115,N_4011,N_3960);
and U4116 (N_4116,N_3953,N_3995);
or U4117 (N_4117,N_3924,N_3966);
and U4118 (N_4118,N_3958,N_3937);
and U4119 (N_4119,N_3969,N_3982);
nor U4120 (N_4120,N_3925,N_4015);
nor U4121 (N_4121,N_4026,N_3981);
or U4122 (N_4122,N_4005,N_3977);
or U4123 (N_4123,N_3943,N_3951);
or U4124 (N_4124,N_4025,N_3993);
nor U4125 (N_4125,N_3926,N_3972);
nor U4126 (N_4126,N_3962,N_3991);
and U4127 (N_4127,N_3971,N_3955);
and U4128 (N_4128,N_3993,N_4041);
nor U4129 (N_4129,N_3982,N_3911);
nand U4130 (N_4130,N_3984,N_4004);
or U4131 (N_4131,N_3964,N_4022);
nand U4132 (N_4132,N_3941,N_3975);
or U4133 (N_4133,N_4041,N_4019);
or U4134 (N_4134,N_3967,N_3930);
or U4135 (N_4135,N_4030,N_4008);
nand U4136 (N_4136,N_3923,N_3950);
nand U4137 (N_4137,N_3977,N_4032);
nor U4138 (N_4138,N_3987,N_3928);
nand U4139 (N_4139,N_3995,N_3934);
nand U4140 (N_4140,N_4006,N_3950);
and U4141 (N_4141,N_3924,N_4027);
and U4142 (N_4142,N_4041,N_3939);
or U4143 (N_4143,N_4034,N_3931);
nand U4144 (N_4144,N_3977,N_3923);
or U4145 (N_4145,N_4028,N_3943);
nand U4146 (N_4146,N_4010,N_3965);
nor U4147 (N_4147,N_3934,N_3927);
or U4148 (N_4148,N_3971,N_4008);
nor U4149 (N_4149,N_3929,N_3972);
or U4150 (N_4150,N_3966,N_3951);
or U4151 (N_4151,N_3995,N_4026);
and U4152 (N_4152,N_4013,N_3940);
nand U4153 (N_4153,N_3910,N_3998);
nor U4154 (N_4154,N_3950,N_3985);
or U4155 (N_4155,N_4029,N_4000);
and U4156 (N_4156,N_4005,N_3964);
or U4157 (N_4157,N_4003,N_4019);
nand U4158 (N_4158,N_3942,N_3976);
nand U4159 (N_4159,N_3981,N_3977);
xnor U4160 (N_4160,N_4009,N_4024);
or U4161 (N_4161,N_3905,N_3915);
nor U4162 (N_4162,N_3944,N_3964);
nand U4163 (N_4163,N_3910,N_4006);
and U4164 (N_4164,N_4008,N_3976);
and U4165 (N_4165,N_4039,N_4014);
nand U4166 (N_4166,N_3969,N_4027);
nor U4167 (N_4167,N_4002,N_3914);
nor U4168 (N_4168,N_3982,N_3931);
nand U4169 (N_4169,N_3917,N_3934);
nor U4170 (N_4170,N_4030,N_3962);
nor U4171 (N_4171,N_3962,N_3980);
or U4172 (N_4172,N_3923,N_3990);
nor U4173 (N_4173,N_3930,N_3972);
and U4174 (N_4174,N_4002,N_4031);
nor U4175 (N_4175,N_4034,N_3907);
xor U4176 (N_4176,N_4042,N_3951);
and U4177 (N_4177,N_3971,N_3923);
or U4178 (N_4178,N_3900,N_4029);
nand U4179 (N_4179,N_3988,N_4032);
and U4180 (N_4180,N_4019,N_4028);
nand U4181 (N_4181,N_3990,N_3947);
xnor U4182 (N_4182,N_3929,N_4018);
nor U4183 (N_4183,N_4045,N_4004);
or U4184 (N_4184,N_3946,N_3928);
xor U4185 (N_4185,N_3968,N_3973);
or U4186 (N_4186,N_3904,N_3920);
nand U4187 (N_4187,N_4013,N_3950);
nor U4188 (N_4188,N_4015,N_4008);
or U4189 (N_4189,N_3979,N_4037);
and U4190 (N_4190,N_3942,N_3995);
nor U4191 (N_4191,N_3975,N_3926);
or U4192 (N_4192,N_3981,N_4006);
nand U4193 (N_4193,N_3991,N_4018);
nand U4194 (N_4194,N_3902,N_4025);
nor U4195 (N_4195,N_4004,N_3999);
nor U4196 (N_4196,N_3960,N_4013);
nor U4197 (N_4197,N_4023,N_3989);
xor U4198 (N_4198,N_3985,N_4021);
nand U4199 (N_4199,N_3998,N_4023);
nor U4200 (N_4200,N_4112,N_4083);
nand U4201 (N_4201,N_4185,N_4170);
nand U4202 (N_4202,N_4086,N_4127);
or U4203 (N_4203,N_4132,N_4070);
and U4204 (N_4204,N_4198,N_4152);
and U4205 (N_4205,N_4167,N_4129);
or U4206 (N_4206,N_4135,N_4187);
xor U4207 (N_4207,N_4105,N_4062);
nand U4208 (N_4208,N_4095,N_4162);
xor U4209 (N_4209,N_4145,N_4093);
or U4210 (N_4210,N_4121,N_4074);
xor U4211 (N_4211,N_4157,N_4098);
or U4212 (N_4212,N_4109,N_4190);
nor U4213 (N_4213,N_4097,N_4052);
nor U4214 (N_4214,N_4072,N_4182);
or U4215 (N_4215,N_4153,N_4136);
and U4216 (N_4216,N_4125,N_4173);
nand U4217 (N_4217,N_4056,N_4196);
and U4218 (N_4218,N_4067,N_4063);
and U4219 (N_4219,N_4068,N_4108);
nor U4220 (N_4220,N_4071,N_4172);
or U4221 (N_4221,N_4151,N_4106);
nor U4222 (N_4222,N_4119,N_4183);
and U4223 (N_4223,N_4138,N_4184);
and U4224 (N_4224,N_4165,N_4164);
nor U4225 (N_4225,N_4193,N_4148);
nor U4226 (N_4226,N_4124,N_4141);
nor U4227 (N_4227,N_4096,N_4117);
nor U4228 (N_4228,N_4100,N_4054);
nand U4229 (N_4229,N_4158,N_4065);
nand U4230 (N_4230,N_4103,N_4133);
and U4231 (N_4231,N_4059,N_4128);
nor U4232 (N_4232,N_4177,N_4080);
or U4233 (N_4233,N_4178,N_4149);
or U4234 (N_4234,N_4114,N_4050);
and U4235 (N_4235,N_4176,N_4092);
nand U4236 (N_4236,N_4102,N_4168);
nor U4237 (N_4237,N_4146,N_4180);
or U4238 (N_4238,N_4075,N_4191);
nand U4239 (N_4239,N_4150,N_4077);
xnor U4240 (N_4240,N_4104,N_4139);
and U4241 (N_4241,N_4197,N_4163);
nand U4242 (N_4242,N_4081,N_4194);
or U4243 (N_4243,N_4088,N_4144);
or U4244 (N_4244,N_4122,N_4174);
nor U4245 (N_4245,N_4130,N_4171);
nor U4246 (N_4246,N_4156,N_4115);
or U4247 (N_4247,N_4199,N_4142);
and U4248 (N_4248,N_4099,N_4084);
nand U4249 (N_4249,N_4131,N_4147);
nand U4250 (N_4250,N_4160,N_4123);
xor U4251 (N_4251,N_4087,N_4078);
nand U4252 (N_4252,N_4159,N_4101);
xnor U4253 (N_4253,N_4051,N_4094);
and U4254 (N_4254,N_4181,N_4189);
or U4255 (N_4255,N_4143,N_4069);
and U4256 (N_4256,N_4073,N_4188);
and U4257 (N_4257,N_4166,N_4154);
or U4258 (N_4258,N_4126,N_4082);
and U4259 (N_4259,N_4058,N_4085);
or U4260 (N_4260,N_4110,N_4076);
or U4261 (N_4261,N_4175,N_4118);
or U4262 (N_4262,N_4179,N_4192);
nor U4263 (N_4263,N_4091,N_4140);
and U4264 (N_4264,N_4079,N_4186);
and U4265 (N_4265,N_4120,N_4053);
or U4266 (N_4266,N_4137,N_4111);
xnor U4267 (N_4267,N_4055,N_4060);
and U4268 (N_4268,N_4155,N_4134);
nand U4269 (N_4269,N_4057,N_4161);
nand U4270 (N_4270,N_4116,N_4090);
nor U4271 (N_4271,N_4107,N_4061);
or U4272 (N_4272,N_4066,N_4064);
or U4273 (N_4273,N_4089,N_4113);
nand U4274 (N_4274,N_4195,N_4169);
or U4275 (N_4275,N_4106,N_4137);
nand U4276 (N_4276,N_4190,N_4114);
or U4277 (N_4277,N_4089,N_4064);
nand U4278 (N_4278,N_4137,N_4144);
and U4279 (N_4279,N_4162,N_4134);
nand U4280 (N_4280,N_4059,N_4187);
and U4281 (N_4281,N_4151,N_4146);
nor U4282 (N_4282,N_4198,N_4071);
nor U4283 (N_4283,N_4138,N_4158);
or U4284 (N_4284,N_4083,N_4147);
nand U4285 (N_4285,N_4107,N_4143);
and U4286 (N_4286,N_4142,N_4191);
or U4287 (N_4287,N_4071,N_4154);
nand U4288 (N_4288,N_4057,N_4124);
xnor U4289 (N_4289,N_4161,N_4103);
or U4290 (N_4290,N_4087,N_4093);
or U4291 (N_4291,N_4180,N_4074);
nand U4292 (N_4292,N_4061,N_4114);
nor U4293 (N_4293,N_4125,N_4087);
nor U4294 (N_4294,N_4089,N_4177);
or U4295 (N_4295,N_4112,N_4050);
or U4296 (N_4296,N_4093,N_4139);
nand U4297 (N_4297,N_4053,N_4094);
or U4298 (N_4298,N_4074,N_4197);
nor U4299 (N_4299,N_4115,N_4177);
or U4300 (N_4300,N_4199,N_4089);
or U4301 (N_4301,N_4075,N_4169);
or U4302 (N_4302,N_4056,N_4176);
nand U4303 (N_4303,N_4059,N_4155);
or U4304 (N_4304,N_4181,N_4145);
and U4305 (N_4305,N_4106,N_4089);
nand U4306 (N_4306,N_4146,N_4104);
nand U4307 (N_4307,N_4172,N_4120);
nor U4308 (N_4308,N_4186,N_4138);
nand U4309 (N_4309,N_4108,N_4081);
or U4310 (N_4310,N_4182,N_4064);
and U4311 (N_4311,N_4086,N_4108);
nand U4312 (N_4312,N_4183,N_4120);
and U4313 (N_4313,N_4181,N_4154);
or U4314 (N_4314,N_4121,N_4161);
and U4315 (N_4315,N_4101,N_4063);
nor U4316 (N_4316,N_4070,N_4053);
and U4317 (N_4317,N_4196,N_4189);
nand U4318 (N_4318,N_4094,N_4137);
and U4319 (N_4319,N_4093,N_4177);
xnor U4320 (N_4320,N_4164,N_4106);
nand U4321 (N_4321,N_4144,N_4071);
nand U4322 (N_4322,N_4189,N_4151);
xor U4323 (N_4323,N_4130,N_4187);
nand U4324 (N_4324,N_4153,N_4070);
and U4325 (N_4325,N_4115,N_4080);
nor U4326 (N_4326,N_4187,N_4172);
and U4327 (N_4327,N_4166,N_4100);
nand U4328 (N_4328,N_4056,N_4175);
nor U4329 (N_4329,N_4110,N_4078);
or U4330 (N_4330,N_4069,N_4128);
nand U4331 (N_4331,N_4066,N_4099);
nand U4332 (N_4332,N_4067,N_4130);
and U4333 (N_4333,N_4117,N_4073);
and U4334 (N_4334,N_4096,N_4154);
or U4335 (N_4335,N_4128,N_4169);
and U4336 (N_4336,N_4153,N_4141);
or U4337 (N_4337,N_4082,N_4197);
and U4338 (N_4338,N_4125,N_4073);
nor U4339 (N_4339,N_4122,N_4059);
nand U4340 (N_4340,N_4078,N_4195);
nand U4341 (N_4341,N_4192,N_4163);
or U4342 (N_4342,N_4100,N_4055);
nor U4343 (N_4343,N_4108,N_4153);
nand U4344 (N_4344,N_4185,N_4127);
nor U4345 (N_4345,N_4194,N_4103);
nand U4346 (N_4346,N_4151,N_4176);
or U4347 (N_4347,N_4069,N_4084);
nor U4348 (N_4348,N_4076,N_4174);
and U4349 (N_4349,N_4170,N_4106);
nand U4350 (N_4350,N_4316,N_4262);
nand U4351 (N_4351,N_4343,N_4223);
xnor U4352 (N_4352,N_4260,N_4339);
and U4353 (N_4353,N_4224,N_4243);
or U4354 (N_4354,N_4303,N_4221);
nand U4355 (N_4355,N_4225,N_4322);
or U4356 (N_4356,N_4329,N_4245);
and U4357 (N_4357,N_4204,N_4267);
or U4358 (N_4358,N_4206,N_4288);
nor U4359 (N_4359,N_4227,N_4349);
and U4360 (N_4360,N_4261,N_4340);
nand U4361 (N_4361,N_4337,N_4285);
nor U4362 (N_4362,N_4222,N_4219);
and U4363 (N_4363,N_4326,N_4323);
and U4364 (N_4364,N_4305,N_4237);
nand U4365 (N_4365,N_4319,N_4207);
nand U4366 (N_4366,N_4269,N_4286);
and U4367 (N_4367,N_4320,N_4300);
or U4368 (N_4368,N_4211,N_4255);
or U4369 (N_4369,N_4242,N_4279);
nor U4370 (N_4370,N_4331,N_4281);
or U4371 (N_4371,N_4330,N_4278);
and U4372 (N_4372,N_4333,N_4216);
nand U4373 (N_4373,N_4318,N_4209);
nand U4374 (N_4374,N_4200,N_4265);
and U4375 (N_4375,N_4250,N_4314);
and U4376 (N_4376,N_4298,N_4276);
nor U4377 (N_4377,N_4249,N_4271);
xnor U4378 (N_4378,N_4307,N_4263);
xnor U4379 (N_4379,N_4346,N_4234);
nor U4380 (N_4380,N_4345,N_4290);
and U4381 (N_4381,N_4247,N_4293);
nor U4382 (N_4382,N_4327,N_4254);
nor U4383 (N_4383,N_4287,N_4302);
and U4384 (N_4384,N_4310,N_4258);
nor U4385 (N_4385,N_4239,N_4308);
xor U4386 (N_4386,N_4273,N_4253);
xnor U4387 (N_4387,N_4232,N_4244);
nor U4388 (N_4388,N_4228,N_4274);
and U4389 (N_4389,N_4235,N_4335);
nor U4390 (N_4390,N_4205,N_4332);
or U4391 (N_4391,N_4313,N_4248);
xnor U4392 (N_4392,N_4272,N_4283);
or U4393 (N_4393,N_4240,N_4264);
and U4394 (N_4394,N_4309,N_4295);
and U4395 (N_4395,N_4210,N_4252);
and U4396 (N_4396,N_4321,N_4231);
nand U4397 (N_4397,N_4213,N_4238);
xor U4398 (N_4398,N_4292,N_4296);
nand U4399 (N_4399,N_4312,N_4325);
nor U4400 (N_4400,N_4217,N_4229);
or U4401 (N_4401,N_4241,N_4306);
xnor U4402 (N_4402,N_4214,N_4334);
nand U4403 (N_4403,N_4202,N_4338);
nor U4404 (N_4404,N_4291,N_4259);
xnor U4405 (N_4405,N_4233,N_4201);
nand U4406 (N_4406,N_4348,N_4251);
and U4407 (N_4407,N_4289,N_4215);
and U4408 (N_4408,N_4230,N_4344);
nor U4409 (N_4409,N_4304,N_4266);
nand U4410 (N_4410,N_4218,N_4317);
and U4411 (N_4411,N_4294,N_4256);
nand U4412 (N_4412,N_4270,N_4336);
nand U4413 (N_4413,N_4246,N_4257);
nor U4414 (N_4414,N_4324,N_4208);
nor U4415 (N_4415,N_4203,N_4341);
nand U4416 (N_4416,N_4280,N_4311);
nor U4417 (N_4417,N_4315,N_4226);
or U4418 (N_4418,N_4220,N_4347);
and U4419 (N_4419,N_4301,N_4284);
or U4420 (N_4420,N_4275,N_4236);
and U4421 (N_4421,N_4282,N_4268);
nand U4422 (N_4422,N_4212,N_4342);
nor U4423 (N_4423,N_4277,N_4299);
nand U4424 (N_4424,N_4297,N_4328);
xor U4425 (N_4425,N_4220,N_4313);
and U4426 (N_4426,N_4301,N_4229);
nor U4427 (N_4427,N_4291,N_4248);
nor U4428 (N_4428,N_4282,N_4213);
nor U4429 (N_4429,N_4249,N_4218);
xor U4430 (N_4430,N_4268,N_4312);
nor U4431 (N_4431,N_4333,N_4340);
and U4432 (N_4432,N_4337,N_4254);
xnor U4433 (N_4433,N_4342,N_4341);
or U4434 (N_4434,N_4305,N_4274);
nor U4435 (N_4435,N_4220,N_4321);
nor U4436 (N_4436,N_4310,N_4286);
nor U4437 (N_4437,N_4346,N_4337);
xnor U4438 (N_4438,N_4244,N_4220);
nand U4439 (N_4439,N_4277,N_4334);
nand U4440 (N_4440,N_4250,N_4255);
nand U4441 (N_4441,N_4241,N_4212);
or U4442 (N_4442,N_4307,N_4325);
and U4443 (N_4443,N_4257,N_4306);
and U4444 (N_4444,N_4259,N_4230);
or U4445 (N_4445,N_4260,N_4237);
nand U4446 (N_4446,N_4314,N_4338);
nand U4447 (N_4447,N_4274,N_4318);
and U4448 (N_4448,N_4285,N_4240);
and U4449 (N_4449,N_4293,N_4262);
or U4450 (N_4450,N_4302,N_4245);
xnor U4451 (N_4451,N_4242,N_4215);
nor U4452 (N_4452,N_4258,N_4205);
xnor U4453 (N_4453,N_4310,N_4267);
or U4454 (N_4454,N_4247,N_4246);
nor U4455 (N_4455,N_4205,N_4208);
and U4456 (N_4456,N_4285,N_4252);
and U4457 (N_4457,N_4242,N_4268);
and U4458 (N_4458,N_4333,N_4212);
nor U4459 (N_4459,N_4262,N_4284);
nor U4460 (N_4460,N_4339,N_4293);
and U4461 (N_4461,N_4299,N_4304);
nor U4462 (N_4462,N_4213,N_4316);
and U4463 (N_4463,N_4213,N_4277);
xor U4464 (N_4464,N_4206,N_4285);
nor U4465 (N_4465,N_4319,N_4234);
or U4466 (N_4466,N_4345,N_4242);
nor U4467 (N_4467,N_4265,N_4314);
xnor U4468 (N_4468,N_4224,N_4334);
or U4469 (N_4469,N_4317,N_4256);
or U4470 (N_4470,N_4227,N_4261);
or U4471 (N_4471,N_4233,N_4327);
and U4472 (N_4472,N_4214,N_4321);
xnor U4473 (N_4473,N_4284,N_4270);
nand U4474 (N_4474,N_4212,N_4213);
nand U4475 (N_4475,N_4228,N_4299);
and U4476 (N_4476,N_4233,N_4262);
nor U4477 (N_4477,N_4233,N_4342);
or U4478 (N_4478,N_4326,N_4335);
xnor U4479 (N_4479,N_4218,N_4346);
xor U4480 (N_4480,N_4324,N_4239);
and U4481 (N_4481,N_4256,N_4303);
or U4482 (N_4482,N_4216,N_4273);
and U4483 (N_4483,N_4325,N_4295);
xor U4484 (N_4484,N_4242,N_4260);
xnor U4485 (N_4485,N_4225,N_4232);
nor U4486 (N_4486,N_4292,N_4326);
nor U4487 (N_4487,N_4263,N_4272);
nor U4488 (N_4488,N_4258,N_4308);
and U4489 (N_4489,N_4247,N_4309);
nor U4490 (N_4490,N_4232,N_4301);
nor U4491 (N_4491,N_4224,N_4249);
nand U4492 (N_4492,N_4233,N_4255);
or U4493 (N_4493,N_4207,N_4206);
and U4494 (N_4494,N_4213,N_4328);
nand U4495 (N_4495,N_4346,N_4291);
nor U4496 (N_4496,N_4267,N_4258);
nor U4497 (N_4497,N_4275,N_4282);
or U4498 (N_4498,N_4267,N_4201);
nor U4499 (N_4499,N_4244,N_4291);
nand U4500 (N_4500,N_4492,N_4371);
and U4501 (N_4501,N_4375,N_4442);
nor U4502 (N_4502,N_4351,N_4489);
and U4503 (N_4503,N_4409,N_4397);
xnor U4504 (N_4504,N_4387,N_4389);
nand U4505 (N_4505,N_4367,N_4443);
or U4506 (N_4506,N_4459,N_4356);
or U4507 (N_4507,N_4476,N_4415);
nand U4508 (N_4508,N_4388,N_4416);
and U4509 (N_4509,N_4410,N_4378);
or U4510 (N_4510,N_4439,N_4484);
nor U4511 (N_4511,N_4462,N_4452);
and U4512 (N_4512,N_4391,N_4498);
nand U4513 (N_4513,N_4479,N_4486);
nand U4514 (N_4514,N_4419,N_4434);
nor U4515 (N_4515,N_4407,N_4399);
nor U4516 (N_4516,N_4418,N_4440);
nor U4517 (N_4517,N_4425,N_4398);
nand U4518 (N_4518,N_4355,N_4438);
nand U4519 (N_4519,N_4468,N_4413);
or U4520 (N_4520,N_4385,N_4475);
and U4521 (N_4521,N_4380,N_4386);
nor U4522 (N_4522,N_4376,N_4405);
nand U4523 (N_4523,N_4491,N_4404);
or U4524 (N_4524,N_4411,N_4495);
or U4525 (N_4525,N_4437,N_4396);
nor U4526 (N_4526,N_4402,N_4444);
nor U4527 (N_4527,N_4481,N_4382);
nor U4528 (N_4528,N_4456,N_4359);
and U4529 (N_4529,N_4364,N_4353);
nand U4530 (N_4530,N_4357,N_4424);
xnor U4531 (N_4531,N_4496,N_4370);
and U4532 (N_4532,N_4354,N_4360);
or U4533 (N_4533,N_4499,N_4395);
or U4534 (N_4534,N_4470,N_4473);
or U4535 (N_4535,N_4384,N_4478);
nor U4536 (N_4536,N_4430,N_4463);
and U4537 (N_4537,N_4494,N_4467);
xor U4538 (N_4538,N_4361,N_4460);
nand U4539 (N_4539,N_4432,N_4373);
nor U4540 (N_4540,N_4429,N_4426);
nand U4541 (N_4541,N_4403,N_4461);
or U4542 (N_4542,N_4406,N_4445);
nor U4543 (N_4543,N_4412,N_4472);
nor U4544 (N_4544,N_4451,N_4497);
and U4545 (N_4545,N_4457,N_4465);
nor U4546 (N_4546,N_4455,N_4377);
xor U4547 (N_4547,N_4352,N_4447);
and U4548 (N_4548,N_4358,N_4453);
and U4549 (N_4549,N_4420,N_4441);
nor U4550 (N_4550,N_4454,N_4368);
nor U4551 (N_4551,N_4390,N_4401);
or U4552 (N_4552,N_4400,N_4490);
and U4553 (N_4553,N_4435,N_4433);
nand U4554 (N_4554,N_4421,N_4362);
nor U4555 (N_4555,N_4383,N_4428);
nand U4556 (N_4556,N_4394,N_4469);
or U4557 (N_4557,N_4487,N_4392);
or U4558 (N_4558,N_4381,N_4417);
or U4559 (N_4559,N_4466,N_4449);
and U4560 (N_4560,N_4369,N_4488);
and U4561 (N_4561,N_4448,N_4483);
nand U4562 (N_4562,N_4423,N_4372);
nor U4563 (N_4563,N_4414,N_4493);
nor U4564 (N_4564,N_4363,N_4366);
and U4565 (N_4565,N_4350,N_4379);
or U4566 (N_4566,N_4427,N_4482);
nor U4567 (N_4567,N_4471,N_4485);
nand U4568 (N_4568,N_4408,N_4431);
nor U4569 (N_4569,N_4450,N_4446);
nor U4570 (N_4570,N_4374,N_4458);
or U4571 (N_4571,N_4393,N_4365);
or U4572 (N_4572,N_4464,N_4436);
xor U4573 (N_4573,N_4477,N_4480);
nand U4574 (N_4574,N_4422,N_4474);
or U4575 (N_4575,N_4454,N_4439);
and U4576 (N_4576,N_4478,N_4470);
nand U4577 (N_4577,N_4411,N_4447);
or U4578 (N_4578,N_4360,N_4392);
or U4579 (N_4579,N_4407,N_4457);
nor U4580 (N_4580,N_4364,N_4352);
nand U4581 (N_4581,N_4421,N_4400);
and U4582 (N_4582,N_4413,N_4356);
and U4583 (N_4583,N_4450,N_4454);
nor U4584 (N_4584,N_4363,N_4493);
or U4585 (N_4585,N_4486,N_4375);
xnor U4586 (N_4586,N_4440,N_4434);
nor U4587 (N_4587,N_4383,N_4392);
or U4588 (N_4588,N_4360,N_4462);
xor U4589 (N_4589,N_4416,N_4453);
nand U4590 (N_4590,N_4388,N_4355);
or U4591 (N_4591,N_4427,N_4478);
xnor U4592 (N_4592,N_4460,N_4441);
or U4593 (N_4593,N_4354,N_4383);
and U4594 (N_4594,N_4433,N_4406);
nand U4595 (N_4595,N_4447,N_4365);
or U4596 (N_4596,N_4477,N_4351);
nor U4597 (N_4597,N_4491,N_4449);
or U4598 (N_4598,N_4450,N_4423);
or U4599 (N_4599,N_4424,N_4398);
nor U4600 (N_4600,N_4351,N_4362);
nand U4601 (N_4601,N_4355,N_4456);
nand U4602 (N_4602,N_4418,N_4388);
xor U4603 (N_4603,N_4384,N_4455);
and U4604 (N_4604,N_4469,N_4479);
nand U4605 (N_4605,N_4397,N_4475);
or U4606 (N_4606,N_4455,N_4496);
nand U4607 (N_4607,N_4482,N_4363);
or U4608 (N_4608,N_4468,N_4436);
nand U4609 (N_4609,N_4364,N_4455);
nor U4610 (N_4610,N_4476,N_4429);
and U4611 (N_4611,N_4452,N_4405);
nor U4612 (N_4612,N_4463,N_4425);
and U4613 (N_4613,N_4453,N_4472);
xor U4614 (N_4614,N_4435,N_4368);
nor U4615 (N_4615,N_4453,N_4395);
and U4616 (N_4616,N_4357,N_4414);
or U4617 (N_4617,N_4456,N_4438);
or U4618 (N_4618,N_4465,N_4385);
and U4619 (N_4619,N_4397,N_4373);
or U4620 (N_4620,N_4483,N_4475);
and U4621 (N_4621,N_4458,N_4492);
nand U4622 (N_4622,N_4449,N_4388);
xnor U4623 (N_4623,N_4371,N_4481);
or U4624 (N_4624,N_4426,N_4479);
nand U4625 (N_4625,N_4383,N_4402);
xor U4626 (N_4626,N_4448,N_4437);
nand U4627 (N_4627,N_4461,N_4418);
nand U4628 (N_4628,N_4469,N_4461);
or U4629 (N_4629,N_4388,N_4352);
nand U4630 (N_4630,N_4486,N_4409);
xor U4631 (N_4631,N_4477,N_4449);
and U4632 (N_4632,N_4425,N_4400);
nand U4633 (N_4633,N_4402,N_4385);
nor U4634 (N_4634,N_4350,N_4492);
xnor U4635 (N_4635,N_4354,N_4363);
nand U4636 (N_4636,N_4430,N_4399);
and U4637 (N_4637,N_4492,N_4392);
and U4638 (N_4638,N_4484,N_4448);
nand U4639 (N_4639,N_4390,N_4425);
nand U4640 (N_4640,N_4398,N_4373);
and U4641 (N_4641,N_4494,N_4456);
nand U4642 (N_4642,N_4497,N_4452);
or U4643 (N_4643,N_4376,N_4373);
nand U4644 (N_4644,N_4401,N_4430);
nand U4645 (N_4645,N_4428,N_4493);
and U4646 (N_4646,N_4403,N_4433);
and U4647 (N_4647,N_4411,N_4476);
or U4648 (N_4648,N_4406,N_4375);
nor U4649 (N_4649,N_4432,N_4413);
or U4650 (N_4650,N_4610,N_4586);
xor U4651 (N_4651,N_4556,N_4632);
and U4652 (N_4652,N_4604,N_4574);
nand U4653 (N_4653,N_4522,N_4519);
or U4654 (N_4654,N_4527,N_4615);
or U4655 (N_4655,N_4543,N_4535);
nor U4656 (N_4656,N_4606,N_4517);
nor U4657 (N_4657,N_4501,N_4624);
and U4658 (N_4658,N_4513,N_4555);
nand U4659 (N_4659,N_4551,N_4608);
nand U4660 (N_4660,N_4622,N_4567);
nand U4661 (N_4661,N_4548,N_4540);
nor U4662 (N_4662,N_4623,N_4538);
and U4663 (N_4663,N_4628,N_4585);
nor U4664 (N_4664,N_4581,N_4573);
and U4665 (N_4665,N_4584,N_4518);
nand U4666 (N_4666,N_4642,N_4647);
and U4667 (N_4667,N_4635,N_4560);
and U4668 (N_4668,N_4524,N_4596);
nand U4669 (N_4669,N_4601,N_4578);
or U4670 (N_4670,N_4516,N_4599);
nor U4671 (N_4671,N_4609,N_4562);
xor U4672 (N_4672,N_4534,N_4568);
nor U4673 (N_4673,N_4515,N_4521);
and U4674 (N_4674,N_4545,N_4571);
nand U4675 (N_4675,N_4643,N_4607);
xor U4676 (N_4676,N_4554,N_4532);
nand U4677 (N_4677,N_4592,N_4621);
nand U4678 (N_4678,N_4637,N_4537);
nand U4679 (N_4679,N_4514,N_4593);
nand U4680 (N_4680,N_4566,N_4633);
or U4681 (N_4681,N_4549,N_4526);
or U4682 (N_4682,N_4544,N_4582);
nand U4683 (N_4683,N_4570,N_4631);
or U4684 (N_4684,N_4539,N_4546);
or U4685 (N_4685,N_4508,N_4505);
nand U4686 (N_4686,N_4618,N_4565);
nor U4687 (N_4687,N_4506,N_4591);
nor U4688 (N_4688,N_4520,N_4634);
nand U4689 (N_4689,N_4512,N_4588);
and U4690 (N_4690,N_4523,N_4504);
or U4691 (N_4691,N_4530,N_4583);
or U4692 (N_4692,N_4626,N_4620);
nand U4693 (N_4693,N_4595,N_4553);
nand U4694 (N_4694,N_4536,N_4507);
nand U4695 (N_4695,N_4630,N_4617);
nor U4696 (N_4696,N_4625,N_4603);
or U4697 (N_4697,N_4597,N_4531);
xnor U4698 (N_4698,N_4612,N_4528);
and U4699 (N_4699,N_4550,N_4525);
and U4700 (N_4700,N_4636,N_4502);
xnor U4701 (N_4701,N_4644,N_4638);
or U4702 (N_4702,N_4611,N_4598);
xnor U4703 (N_4703,N_4629,N_4589);
and U4704 (N_4704,N_4646,N_4529);
xor U4705 (N_4705,N_4641,N_4558);
and U4706 (N_4706,N_4600,N_4640);
nor U4707 (N_4707,N_4639,N_4572);
nor U4708 (N_4708,N_4561,N_4569);
nand U4709 (N_4709,N_4575,N_4509);
or U4710 (N_4710,N_4627,N_4511);
xnor U4711 (N_4711,N_4563,N_4541);
nor U4712 (N_4712,N_4576,N_4613);
xor U4713 (N_4713,N_4579,N_4645);
or U4714 (N_4714,N_4577,N_4559);
nor U4715 (N_4715,N_4533,N_4552);
xor U4716 (N_4716,N_4500,N_4547);
nand U4717 (N_4717,N_4649,N_4557);
nand U4718 (N_4718,N_4542,N_4602);
or U4719 (N_4719,N_4580,N_4605);
nor U4720 (N_4720,N_4510,N_4594);
nand U4721 (N_4721,N_4564,N_4590);
xnor U4722 (N_4722,N_4503,N_4614);
nor U4723 (N_4723,N_4619,N_4648);
nor U4724 (N_4724,N_4616,N_4587);
and U4725 (N_4725,N_4555,N_4503);
and U4726 (N_4726,N_4550,N_4627);
and U4727 (N_4727,N_4594,N_4577);
or U4728 (N_4728,N_4549,N_4586);
or U4729 (N_4729,N_4574,N_4600);
nand U4730 (N_4730,N_4523,N_4591);
nand U4731 (N_4731,N_4605,N_4550);
nor U4732 (N_4732,N_4626,N_4613);
nor U4733 (N_4733,N_4552,N_4554);
nor U4734 (N_4734,N_4553,N_4579);
and U4735 (N_4735,N_4590,N_4554);
or U4736 (N_4736,N_4625,N_4587);
or U4737 (N_4737,N_4526,N_4569);
and U4738 (N_4738,N_4534,N_4616);
or U4739 (N_4739,N_4555,N_4552);
nor U4740 (N_4740,N_4607,N_4503);
and U4741 (N_4741,N_4580,N_4506);
nand U4742 (N_4742,N_4605,N_4587);
nand U4743 (N_4743,N_4649,N_4577);
or U4744 (N_4744,N_4647,N_4573);
nand U4745 (N_4745,N_4600,N_4540);
nor U4746 (N_4746,N_4529,N_4511);
and U4747 (N_4747,N_4642,N_4608);
xor U4748 (N_4748,N_4502,N_4595);
or U4749 (N_4749,N_4623,N_4572);
nor U4750 (N_4750,N_4537,N_4549);
nand U4751 (N_4751,N_4519,N_4633);
xnor U4752 (N_4752,N_4513,N_4620);
nand U4753 (N_4753,N_4553,N_4645);
or U4754 (N_4754,N_4514,N_4616);
or U4755 (N_4755,N_4541,N_4588);
or U4756 (N_4756,N_4564,N_4613);
nor U4757 (N_4757,N_4641,N_4573);
xnor U4758 (N_4758,N_4513,N_4519);
and U4759 (N_4759,N_4607,N_4636);
and U4760 (N_4760,N_4635,N_4615);
nor U4761 (N_4761,N_4611,N_4533);
nand U4762 (N_4762,N_4567,N_4610);
or U4763 (N_4763,N_4575,N_4622);
nor U4764 (N_4764,N_4603,N_4518);
or U4765 (N_4765,N_4632,N_4639);
nor U4766 (N_4766,N_4639,N_4636);
nand U4767 (N_4767,N_4575,N_4538);
nor U4768 (N_4768,N_4580,N_4541);
xnor U4769 (N_4769,N_4508,N_4618);
or U4770 (N_4770,N_4543,N_4630);
nand U4771 (N_4771,N_4528,N_4581);
nor U4772 (N_4772,N_4502,N_4585);
and U4773 (N_4773,N_4561,N_4552);
or U4774 (N_4774,N_4628,N_4544);
nor U4775 (N_4775,N_4565,N_4598);
nor U4776 (N_4776,N_4600,N_4582);
nand U4777 (N_4777,N_4571,N_4625);
and U4778 (N_4778,N_4624,N_4527);
nor U4779 (N_4779,N_4569,N_4533);
nand U4780 (N_4780,N_4509,N_4592);
and U4781 (N_4781,N_4530,N_4566);
nand U4782 (N_4782,N_4586,N_4573);
and U4783 (N_4783,N_4622,N_4534);
xor U4784 (N_4784,N_4553,N_4525);
xor U4785 (N_4785,N_4606,N_4635);
or U4786 (N_4786,N_4576,N_4596);
or U4787 (N_4787,N_4533,N_4588);
and U4788 (N_4788,N_4605,N_4615);
nor U4789 (N_4789,N_4513,N_4526);
nor U4790 (N_4790,N_4642,N_4571);
nand U4791 (N_4791,N_4592,N_4598);
xnor U4792 (N_4792,N_4549,N_4564);
nor U4793 (N_4793,N_4588,N_4603);
nand U4794 (N_4794,N_4599,N_4571);
xor U4795 (N_4795,N_4644,N_4549);
or U4796 (N_4796,N_4528,N_4643);
nand U4797 (N_4797,N_4635,N_4546);
nor U4798 (N_4798,N_4544,N_4542);
xor U4799 (N_4799,N_4595,N_4566);
nand U4800 (N_4800,N_4718,N_4741);
nand U4801 (N_4801,N_4687,N_4708);
nor U4802 (N_4802,N_4724,N_4722);
nor U4803 (N_4803,N_4699,N_4666);
or U4804 (N_4804,N_4677,N_4705);
nand U4805 (N_4805,N_4692,N_4728);
or U4806 (N_4806,N_4753,N_4760);
and U4807 (N_4807,N_4788,N_4721);
and U4808 (N_4808,N_4653,N_4723);
nor U4809 (N_4809,N_4725,N_4787);
nand U4810 (N_4810,N_4650,N_4657);
and U4811 (N_4811,N_4763,N_4696);
or U4812 (N_4812,N_4765,N_4756);
xor U4813 (N_4813,N_4661,N_4748);
or U4814 (N_4814,N_4656,N_4668);
or U4815 (N_4815,N_4663,N_4738);
nor U4816 (N_4816,N_4700,N_4780);
nor U4817 (N_4817,N_4671,N_4710);
and U4818 (N_4818,N_4799,N_4676);
nor U4819 (N_4819,N_4703,N_4793);
and U4820 (N_4820,N_4698,N_4751);
nor U4821 (N_4821,N_4768,N_4706);
nor U4822 (N_4822,N_4680,N_4744);
nor U4823 (N_4823,N_4758,N_4777);
nor U4824 (N_4824,N_4735,N_4683);
and U4825 (N_4825,N_4673,N_4752);
nand U4826 (N_4826,N_4704,N_4659);
or U4827 (N_4827,N_4726,N_4757);
or U4828 (N_4828,N_4750,N_4767);
nor U4829 (N_4829,N_4747,N_4778);
and U4830 (N_4830,N_4690,N_4720);
and U4831 (N_4831,N_4679,N_4769);
nor U4832 (N_4832,N_4749,N_4798);
nand U4833 (N_4833,N_4740,N_4702);
nor U4834 (N_4834,N_4713,N_4717);
nand U4835 (N_4835,N_4662,N_4695);
or U4836 (N_4836,N_4784,N_4785);
nand U4837 (N_4837,N_4678,N_4754);
and U4838 (N_4838,N_4789,N_4736);
and U4839 (N_4839,N_4711,N_4783);
xnor U4840 (N_4840,N_4761,N_4693);
nand U4841 (N_4841,N_4770,N_4697);
and U4842 (N_4842,N_4782,N_4691);
and U4843 (N_4843,N_4727,N_4797);
and U4844 (N_4844,N_4762,N_4660);
xnor U4845 (N_4845,N_4779,N_4731);
and U4846 (N_4846,N_4701,N_4681);
nand U4847 (N_4847,N_4790,N_4688);
and U4848 (N_4848,N_4716,N_4792);
and U4849 (N_4849,N_4776,N_4652);
nor U4850 (N_4850,N_4732,N_4796);
nor U4851 (N_4851,N_4664,N_4774);
and U4852 (N_4852,N_4694,N_4743);
and U4853 (N_4853,N_4773,N_4794);
nand U4854 (N_4854,N_4654,N_4714);
nand U4855 (N_4855,N_4772,N_4675);
nand U4856 (N_4856,N_4759,N_4775);
nor U4857 (N_4857,N_4746,N_4665);
or U4858 (N_4858,N_4766,N_4669);
or U4859 (N_4859,N_4764,N_4771);
xor U4860 (N_4860,N_4730,N_4729);
and U4861 (N_4861,N_4682,N_4715);
or U4862 (N_4862,N_4674,N_4737);
nand U4863 (N_4863,N_4733,N_4719);
nand U4864 (N_4864,N_4670,N_4655);
or U4865 (N_4865,N_4739,N_4651);
and U4866 (N_4866,N_4684,N_4712);
and U4867 (N_4867,N_4742,N_4658);
nand U4868 (N_4868,N_4745,N_4755);
nor U4869 (N_4869,N_4709,N_4685);
and U4870 (N_4870,N_4686,N_4667);
nand U4871 (N_4871,N_4781,N_4734);
and U4872 (N_4872,N_4795,N_4786);
or U4873 (N_4873,N_4689,N_4791);
and U4874 (N_4874,N_4672,N_4707);
and U4875 (N_4875,N_4766,N_4777);
nor U4876 (N_4876,N_4688,N_4677);
or U4877 (N_4877,N_4680,N_4677);
or U4878 (N_4878,N_4721,N_4765);
nand U4879 (N_4879,N_4656,N_4650);
xor U4880 (N_4880,N_4720,N_4728);
nand U4881 (N_4881,N_4745,N_4660);
nand U4882 (N_4882,N_4718,N_4661);
nand U4883 (N_4883,N_4686,N_4669);
nor U4884 (N_4884,N_4692,N_4675);
nand U4885 (N_4885,N_4786,N_4778);
and U4886 (N_4886,N_4715,N_4795);
or U4887 (N_4887,N_4674,N_4698);
and U4888 (N_4888,N_4769,N_4759);
or U4889 (N_4889,N_4659,N_4748);
nand U4890 (N_4890,N_4737,N_4724);
nor U4891 (N_4891,N_4737,N_4706);
and U4892 (N_4892,N_4746,N_4724);
nor U4893 (N_4893,N_4780,N_4799);
and U4894 (N_4894,N_4694,N_4792);
and U4895 (N_4895,N_4681,N_4747);
and U4896 (N_4896,N_4746,N_4656);
and U4897 (N_4897,N_4746,N_4790);
nor U4898 (N_4898,N_4665,N_4772);
and U4899 (N_4899,N_4686,N_4725);
and U4900 (N_4900,N_4712,N_4737);
xor U4901 (N_4901,N_4739,N_4759);
or U4902 (N_4902,N_4721,N_4666);
nand U4903 (N_4903,N_4792,N_4665);
nor U4904 (N_4904,N_4654,N_4781);
nor U4905 (N_4905,N_4654,N_4739);
xor U4906 (N_4906,N_4753,N_4726);
and U4907 (N_4907,N_4767,N_4796);
nor U4908 (N_4908,N_4787,N_4741);
and U4909 (N_4909,N_4742,N_4724);
nand U4910 (N_4910,N_4650,N_4785);
xnor U4911 (N_4911,N_4716,N_4702);
nor U4912 (N_4912,N_4657,N_4786);
nand U4913 (N_4913,N_4782,N_4772);
and U4914 (N_4914,N_4793,N_4710);
and U4915 (N_4915,N_4718,N_4779);
and U4916 (N_4916,N_4710,N_4681);
nor U4917 (N_4917,N_4667,N_4705);
or U4918 (N_4918,N_4786,N_4762);
or U4919 (N_4919,N_4759,N_4698);
and U4920 (N_4920,N_4752,N_4769);
and U4921 (N_4921,N_4679,N_4719);
and U4922 (N_4922,N_4717,N_4731);
or U4923 (N_4923,N_4740,N_4695);
nand U4924 (N_4924,N_4732,N_4692);
or U4925 (N_4925,N_4683,N_4705);
nand U4926 (N_4926,N_4665,N_4768);
nor U4927 (N_4927,N_4741,N_4786);
and U4928 (N_4928,N_4672,N_4789);
nor U4929 (N_4929,N_4741,N_4799);
xor U4930 (N_4930,N_4727,N_4719);
nor U4931 (N_4931,N_4792,N_4687);
nand U4932 (N_4932,N_4698,N_4655);
xnor U4933 (N_4933,N_4722,N_4731);
or U4934 (N_4934,N_4764,N_4713);
nand U4935 (N_4935,N_4763,N_4796);
and U4936 (N_4936,N_4747,N_4667);
nor U4937 (N_4937,N_4793,N_4737);
nand U4938 (N_4938,N_4689,N_4666);
and U4939 (N_4939,N_4787,N_4747);
or U4940 (N_4940,N_4657,N_4700);
or U4941 (N_4941,N_4746,N_4714);
or U4942 (N_4942,N_4722,N_4655);
or U4943 (N_4943,N_4680,N_4746);
and U4944 (N_4944,N_4699,N_4753);
nor U4945 (N_4945,N_4763,N_4700);
or U4946 (N_4946,N_4710,N_4763);
nand U4947 (N_4947,N_4742,N_4783);
nor U4948 (N_4948,N_4767,N_4738);
nor U4949 (N_4949,N_4684,N_4762);
and U4950 (N_4950,N_4809,N_4931);
nand U4951 (N_4951,N_4932,N_4863);
xnor U4952 (N_4952,N_4850,N_4877);
nand U4953 (N_4953,N_4805,N_4858);
and U4954 (N_4954,N_4913,N_4866);
nor U4955 (N_4955,N_4845,N_4807);
nor U4956 (N_4956,N_4912,N_4859);
nor U4957 (N_4957,N_4928,N_4876);
or U4958 (N_4958,N_4848,N_4935);
or U4959 (N_4959,N_4884,N_4925);
nand U4960 (N_4960,N_4933,N_4904);
nand U4961 (N_4961,N_4829,N_4944);
nand U4962 (N_4962,N_4847,N_4869);
nor U4963 (N_4963,N_4834,N_4947);
nor U4964 (N_4964,N_4911,N_4801);
or U4965 (N_4965,N_4891,N_4810);
nor U4966 (N_4966,N_4818,N_4898);
and U4967 (N_4967,N_4846,N_4923);
and U4968 (N_4968,N_4890,N_4819);
and U4969 (N_4969,N_4835,N_4822);
or U4970 (N_4970,N_4856,N_4939);
nand U4971 (N_4971,N_4903,N_4815);
or U4972 (N_4972,N_4927,N_4878);
nand U4973 (N_4973,N_4907,N_4823);
nor U4974 (N_4974,N_4838,N_4942);
and U4975 (N_4975,N_4874,N_4906);
or U4976 (N_4976,N_4934,N_4905);
and U4977 (N_4977,N_4851,N_4888);
and U4978 (N_4978,N_4892,N_4832);
or U4979 (N_4979,N_4879,N_4864);
nor U4980 (N_4980,N_4826,N_4883);
or U4981 (N_4981,N_4875,N_4921);
and U4982 (N_4982,N_4841,N_4860);
nand U4983 (N_4983,N_4929,N_4893);
and U4984 (N_4984,N_4828,N_4861);
nand U4985 (N_4985,N_4889,N_4936);
and U4986 (N_4986,N_4894,N_4948);
nor U4987 (N_4987,N_4854,N_4836);
nor U4988 (N_4988,N_4867,N_4842);
or U4989 (N_4989,N_4817,N_4940);
nor U4990 (N_4990,N_4813,N_4821);
xnor U4991 (N_4991,N_4885,N_4849);
and U4992 (N_4992,N_4833,N_4831);
nand U4993 (N_4993,N_4872,N_4937);
or U4994 (N_4994,N_4895,N_4868);
nor U4995 (N_4995,N_4941,N_4824);
nor U4996 (N_4996,N_4945,N_4924);
xor U4997 (N_4997,N_4811,N_4896);
or U4998 (N_4998,N_4881,N_4816);
and U4999 (N_4999,N_4914,N_4910);
or U5000 (N_5000,N_4839,N_4837);
or U5001 (N_5001,N_4930,N_4800);
xor U5002 (N_5002,N_4915,N_4887);
or U5003 (N_5003,N_4926,N_4855);
nand U5004 (N_5004,N_4862,N_4871);
and U5005 (N_5005,N_4873,N_4844);
nor U5006 (N_5006,N_4857,N_4916);
or U5007 (N_5007,N_4840,N_4886);
nor U5008 (N_5008,N_4812,N_4899);
xnor U5009 (N_5009,N_4806,N_4946);
and U5010 (N_5010,N_4882,N_4897);
or U5011 (N_5011,N_4802,N_4922);
nor U5012 (N_5012,N_4804,N_4908);
nor U5013 (N_5013,N_4902,N_4909);
nor U5014 (N_5014,N_4917,N_4949);
nand U5015 (N_5015,N_4808,N_4827);
nand U5016 (N_5016,N_4938,N_4843);
nor U5017 (N_5017,N_4820,N_4920);
or U5018 (N_5018,N_4852,N_4814);
or U5019 (N_5019,N_4900,N_4830);
xnor U5020 (N_5020,N_4901,N_4943);
nor U5021 (N_5021,N_4918,N_4865);
and U5022 (N_5022,N_4803,N_4919);
or U5023 (N_5023,N_4880,N_4853);
and U5024 (N_5024,N_4870,N_4825);
and U5025 (N_5025,N_4938,N_4944);
and U5026 (N_5026,N_4941,N_4848);
and U5027 (N_5027,N_4922,N_4873);
and U5028 (N_5028,N_4871,N_4849);
nand U5029 (N_5029,N_4847,N_4820);
or U5030 (N_5030,N_4945,N_4824);
nor U5031 (N_5031,N_4814,N_4949);
or U5032 (N_5032,N_4863,N_4936);
nor U5033 (N_5033,N_4825,N_4883);
or U5034 (N_5034,N_4892,N_4814);
or U5035 (N_5035,N_4889,N_4919);
xnor U5036 (N_5036,N_4932,N_4856);
nor U5037 (N_5037,N_4887,N_4842);
nand U5038 (N_5038,N_4917,N_4831);
nand U5039 (N_5039,N_4824,N_4899);
nor U5040 (N_5040,N_4811,N_4849);
nand U5041 (N_5041,N_4932,N_4921);
nor U5042 (N_5042,N_4852,N_4881);
nor U5043 (N_5043,N_4891,N_4935);
and U5044 (N_5044,N_4913,N_4852);
and U5045 (N_5045,N_4870,N_4913);
or U5046 (N_5046,N_4923,N_4941);
and U5047 (N_5047,N_4882,N_4820);
nand U5048 (N_5048,N_4947,N_4943);
or U5049 (N_5049,N_4897,N_4817);
or U5050 (N_5050,N_4949,N_4810);
nor U5051 (N_5051,N_4939,N_4831);
and U5052 (N_5052,N_4937,N_4811);
and U5053 (N_5053,N_4892,N_4896);
nor U5054 (N_5054,N_4848,N_4910);
nor U5055 (N_5055,N_4869,N_4910);
or U5056 (N_5056,N_4892,N_4922);
xnor U5057 (N_5057,N_4882,N_4847);
nor U5058 (N_5058,N_4927,N_4817);
or U5059 (N_5059,N_4896,N_4940);
or U5060 (N_5060,N_4829,N_4925);
and U5061 (N_5061,N_4862,N_4948);
xnor U5062 (N_5062,N_4948,N_4856);
nor U5063 (N_5063,N_4843,N_4800);
nor U5064 (N_5064,N_4866,N_4923);
nand U5065 (N_5065,N_4858,N_4808);
or U5066 (N_5066,N_4915,N_4880);
and U5067 (N_5067,N_4939,N_4885);
nand U5068 (N_5068,N_4891,N_4880);
xnor U5069 (N_5069,N_4800,N_4832);
and U5070 (N_5070,N_4937,N_4916);
nor U5071 (N_5071,N_4943,N_4826);
nand U5072 (N_5072,N_4848,N_4922);
nand U5073 (N_5073,N_4810,N_4901);
and U5074 (N_5074,N_4850,N_4870);
nand U5075 (N_5075,N_4817,N_4830);
and U5076 (N_5076,N_4863,N_4923);
nor U5077 (N_5077,N_4887,N_4901);
nand U5078 (N_5078,N_4930,N_4922);
or U5079 (N_5079,N_4852,N_4900);
nor U5080 (N_5080,N_4875,N_4833);
or U5081 (N_5081,N_4830,N_4882);
nand U5082 (N_5082,N_4900,N_4940);
and U5083 (N_5083,N_4884,N_4816);
and U5084 (N_5084,N_4850,N_4911);
and U5085 (N_5085,N_4948,N_4857);
nand U5086 (N_5086,N_4874,N_4899);
xnor U5087 (N_5087,N_4810,N_4867);
or U5088 (N_5088,N_4938,N_4923);
or U5089 (N_5089,N_4933,N_4903);
nand U5090 (N_5090,N_4893,N_4874);
nor U5091 (N_5091,N_4860,N_4834);
xnor U5092 (N_5092,N_4882,N_4861);
or U5093 (N_5093,N_4851,N_4826);
and U5094 (N_5094,N_4948,N_4801);
or U5095 (N_5095,N_4814,N_4878);
nand U5096 (N_5096,N_4868,N_4839);
nor U5097 (N_5097,N_4806,N_4803);
nand U5098 (N_5098,N_4838,N_4802);
nand U5099 (N_5099,N_4841,N_4843);
nand U5100 (N_5100,N_5011,N_5063);
xnor U5101 (N_5101,N_5085,N_4974);
nand U5102 (N_5102,N_5049,N_5077);
and U5103 (N_5103,N_4970,N_5005);
or U5104 (N_5104,N_4957,N_4993);
and U5105 (N_5105,N_5089,N_4998);
and U5106 (N_5106,N_5054,N_5096);
and U5107 (N_5107,N_5012,N_5006);
or U5108 (N_5108,N_5080,N_5088);
nand U5109 (N_5109,N_5052,N_5059);
nor U5110 (N_5110,N_4973,N_5092);
or U5111 (N_5111,N_5032,N_5040);
and U5112 (N_5112,N_5016,N_4954);
nor U5113 (N_5113,N_5013,N_5081);
nand U5114 (N_5114,N_5015,N_5044);
and U5115 (N_5115,N_5064,N_5017);
nor U5116 (N_5116,N_5069,N_5036);
and U5117 (N_5117,N_4969,N_4985);
xor U5118 (N_5118,N_5055,N_5020);
nand U5119 (N_5119,N_5007,N_4962);
nand U5120 (N_5120,N_5002,N_4981);
xnor U5121 (N_5121,N_5071,N_5034);
or U5122 (N_5122,N_5062,N_5078);
nor U5123 (N_5123,N_4952,N_5030);
or U5124 (N_5124,N_4991,N_5082);
nor U5125 (N_5125,N_5065,N_4967);
nand U5126 (N_5126,N_4972,N_5087);
nand U5127 (N_5127,N_5084,N_5004);
and U5128 (N_5128,N_4990,N_4971);
or U5129 (N_5129,N_4995,N_5067);
or U5130 (N_5130,N_5043,N_4966);
nor U5131 (N_5131,N_5000,N_5097);
nand U5132 (N_5132,N_5056,N_5090);
xnor U5133 (N_5133,N_4997,N_5001);
xnor U5134 (N_5134,N_5031,N_5073);
nor U5135 (N_5135,N_4964,N_4983);
nor U5136 (N_5136,N_5099,N_5061);
nor U5137 (N_5137,N_4992,N_4977);
nand U5138 (N_5138,N_5074,N_4955);
nor U5139 (N_5139,N_5019,N_4975);
nor U5140 (N_5140,N_5083,N_5066);
nor U5141 (N_5141,N_4999,N_5094);
nor U5142 (N_5142,N_5039,N_5028);
nor U5143 (N_5143,N_4980,N_5047);
and U5144 (N_5144,N_5048,N_4953);
or U5145 (N_5145,N_5025,N_4956);
and U5146 (N_5146,N_5035,N_5042);
nor U5147 (N_5147,N_5023,N_5095);
nor U5148 (N_5148,N_5053,N_5051);
and U5149 (N_5149,N_4958,N_5070);
nand U5150 (N_5150,N_5046,N_4994);
nand U5151 (N_5151,N_5014,N_4982);
nand U5152 (N_5152,N_5050,N_5093);
nand U5153 (N_5153,N_4950,N_4976);
or U5154 (N_5154,N_5060,N_5038);
nand U5155 (N_5155,N_5029,N_4989);
nor U5156 (N_5156,N_4978,N_4960);
nand U5157 (N_5157,N_4986,N_4968);
or U5158 (N_5158,N_5041,N_5033);
nand U5159 (N_5159,N_4987,N_5072);
nand U5160 (N_5160,N_4965,N_5076);
or U5161 (N_5161,N_5068,N_5009);
or U5162 (N_5162,N_5018,N_5098);
nand U5163 (N_5163,N_5024,N_5021);
nand U5164 (N_5164,N_4959,N_5057);
nor U5165 (N_5165,N_5010,N_5086);
nand U5166 (N_5166,N_5027,N_5091);
or U5167 (N_5167,N_5075,N_4984);
nand U5168 (N_5168,N_4951,N_5022);
nand U5169 (N_5169,N_4996,N_5003);
and U5170 (N_5170,N_5058,N_4961);
and U5171 (N_5171,N_5008,N_5026);
nor U5172 (N_5172,N_5079,N_4979);
nor U5173 (N_5173,N_5045,N_4988);
or U5174 (N_5174,N_5037,N_4963);
or U5175 (N_5175,N_5092,N_5086);
xnor U5176 (N_5176,N_5095,N_5062);
and U5177 (N_5177,N_4995,N_5009);
nand U5178 (N_5178,N_5071,N_5082);
nor U5179 (N_5179,N_5029,N_4979);
nor U5180 (N_5180,N_4980,N_5010);
nand U5181 (N_5181,N_5011,N_5053);
or U5182 (N_5182,N_4966,N_5069);
nor U5183 (N_5183,N_5034,N_5002);
and U5184 (N_5184,N_5037,N_4961);
and U5185 (N_5185,N_5050,N_5095);
nand U5186 (N_5186,N_5055,N_5040);
nor U5187 (N_5187,N_5027,N_4974);
xor U5188 (N_5188,N_5050,N_5059);
nand U5189 (N_5189,N_5002,N_5062);
or U5190 (N_5190,N_4968,N_5070);
and U5191 (N_5191,N_4975,N_4984);
and U5192 (N_5192,N_4976,N_4975);
nand U5193 (N_5193,N_4961,N_5062);
and U5194 (N_5194,N_4954,N_5062);
and U5195 (N_5195,N_4982,N_5066);
and U5196 (N_5196,N_4986,N_4995);
and U5197 (N_5197,N_4955,N_4971);
nand U5198 (N_5198,N_5032,N_5024);
and U5199 (N_5199,N_5073,N_5000);
nor U5200 (N_5200,N_5028,N_5098);
nor U5201 (N_5201,N_4998,N_4984);
nand U5202 (N_5202,N_4955,N_5008);
and U5203 (N_5203,N_4972,N_5074);
or U5204 (N_5204,N_5009,N_4963);
xor U5205 (N_5205,N_5083,N_4982);
nand U5206 (N_5206,N_4956,N_4992);
or U5207 (N_5207,N_5004,N_4984);
and U5208 (N_5208,N_5016,N_4950);
or U5209 (N_5209,N_5024,N_4966);
or U5210 (N_5210,N_5036,N_4964);
and U5211 (N_5211,N_5014,N_5063);
or U5212 (N_5212,N_5012,N_5057);
nand U5213 (N_5213,N_5085,N_4962);
and U5214 (N_5214,N_5004,N_5056);
or U5215 (N_5215,N_5044,N_5068);
or U5216 (N_5216,N_5038,N_5007);
or U5217 (N_5217,N_4963,N_5089);
nor U5218 (N_5218,N_4996,N_4964);
xnor U5219 (N_5219,N_5015,N_5002);
nor U5220 (N_5220,N_5057,N_4985);
nor U5221 (N_5221,N_5054,N_5042);
nor U5222 (N_5222,N_5057,N_4991);
nand U5223 (N_5223,N_4989,N_5068);
and U5224 (N_5224,N_5003,N_4969);
nor U5225 (N_5225,N_5068,N_4961);
and U5226 (N_5226,N_5013,N_4959);
xor U5227 (N_5227,N_5066,N_5044);
nand U5228 (N_5228,N_4994,N_5061);
nor U5229 (N_5229,N_5061,N_4957);
nand U5230 (N_5230,N_4994,N_5066);
and U5231 (N_5231,N_4984,N_5030);
or U5232 (N_5232,N_5000,N_5061);
and U5233 (N_5233,N_5097,N_4972);
nand U5234 (N_5234,N_5011,N_4953);
nor U5235 (N_5235,N_5013,N_4989);
and U5236 (N_5236,N_4950,N_5023);
and U5237 (N_5237,N_4973,N_5072);
or U5238 (N_5238,N_4965,N_5008);
xnor U5239 (N_5239,N_4970,N_5086);
nand U5240 (N_5240,N_4979,N_4965);
nand U5241 (N_5241,N_4953,N_4992);
nor U5242 (N_5242,N_5008,N_5079);
or U5243 (N_5243,N_5023,N_5034);
or U5244 (N_5244,N_5018,N_5080);
or U5245 (N_5245,N_4952,N_5099);
or U5246 (N_5246,N_5029,N_4977);
or U5247 (N_5247,N_4972,N_5033);
nand U5248 (N_5248,N_5017,N_5021);
xnor U5249 (N_5249,N_5074,N_4960);
or U5250 (N_5250,N_5206,N_5138);
or U5251 (N_5251,N_5176,N_5132);
nor U5252 (N_5252,N_5187,N_5123);
nor U5253 (N_5253,N_5131,N_5189);
nand U5254 (N_5254,N_5129,N_5182);
or U5255 (N_5255,N_5185,N_5193);
or U5256 (N_5256,N_5183,N_5207);
nand U5257 (N_5257,N_5199,N_5103);
nor U5258 (N_5258,N_5155,N_5227);
or U5259 (N_5259,N_5229,N_5208);
xnor U5260 (N_5260,N_5109,N_5244);
nor U5261 (N_5261,N_5214,N_5130);
or U5262 (N_5262,N_5152,N_5234);
nor U5263 (N_5263,N_5168,N_5224);
or U5264 (N_5264,N_5160,N_5162);
nor U5265 (N_5265,N_5242,N_5197);
xor U5266 (N_5266,N_5105,N_5198);
or U5267 (N_5267,N_5125,N_5164);
nand U5268 (N_5268,N_5165,N_5108);
and U5269 (N_5269,N_5135,N_5142);
nand U5270 (N_5270,N_5205,N_5172);
nand U5271 (N_5271,N_5186,N_5213);
or U5272 (N_5272,N_5216,N_5243);
or U5273 (N_5273,N_5117,N_5167);
nand U5274 (N_5274,N_5128,N_5233);
nor U5275 (N_5275,N_5156,N_5111);
or U5276 (N_5276,N_5201,N_5173);
nand U5277 (N_5277,N_5226,N_5232);
nand U5278 (N_5278,N_5147,N_5113);
xnor U5279 (N_5279,N_5100,N_5222);
xor U5280 (N_5280,N_5166,N_5200);
or U5281 (N_5281,N_5220,N_5126);
xnor U5282 (N_5282,N_5212,N_5163);
or U5283 (N_5283,N_5110,N_5238);
nor U5284 (N_5284,N_5120,N_5121);
and U5285 (N_5285,N_5139,N_5116);
nor U5286 (N_5286,N_5159,N_5134);
nor U5287 (N_5287,N_5223,N_5191);
nor U5288 (N_5288,N_5118,N_5235);
nand U5289 (N_5289,N_5188,N_5115);
or U5290 (N_5290,N_5179,N_5248);
and U5291 (N_5291,N_5230,N_5127);
nand U5292 (N_5292,N_5209,N_5124);
xnor U5293 (N_5293,N_5175,N_5204);
and U5294 (N_5294,N_5211,N_5247);
nand U5295 (N_5295,N_5150,N_5202);
nor U5296 (N_5296,N_5239,N_5249);
or U5297 (N_5297,N_5145,N_5101);
and U5298 (N_5298,N_5144,N_5114);
nor U5299 (N_5299,N_5210,N_5236);
nor U5300 (N_5300,N_5104,N_5169);
and U5301 (N_5301,N_5148,N_5140);
nand U5302 (N_5302,N_5170,N_5180);
and U5303 (N_5303,N_5158,N_5141);
and U5304 (N_5304,N_5184,N_5107);
or U5305 (N_5305,N_5161,N_5143);
nand U5306 (N_5306,N_5225,N_5190);
and U5307 (N_5307,N_5157,N_5178);
or U5308 (N_5308,N_5219,N_5177);
xnor U5309 (N_5309,N_5106,N_5136);
and U5310 (N_5310,N_5203,N_5112);
nor U5311 (N_5311,N_5192,N_5194);
nor U5312 (N_5312,N_5149,N_5151);
or U5313 (N_5313,N_5196,N_5146);
nand U5314 (N_5314,N_5137,N_5174);
and U5315 (N_5315,N_5221,N_5246);
or U5316 (N_5316,N_5195,N_5133);
or U5317 (N_5317,N_5237,N_5215);
nand U5318 (N_5318,N_5241,N_5154);
nor U5319 (N_5319,N_5231,N_5218);
or U5320 (N_5320,N_5171,N_5102);
nand U5321 (N_5321,N_5217,N_5240);
and U5322 (N_5322,N_5119,N_5245);
and U5323 (N_5323,N_5122,N_5228);
nand U5324 (N_5324,N_5153,N_5181);
nand U5325 (N_5325,N_5129,N_5233);
or U5326 (N_5326,N_5161,N_5205);
nand U5327 (N_5327,N_5169,N_5232);
nand U5328 (N_5328,N_5161,N_5226);
nor U5329 (N_5329,N_5186,N_5229);
nor U5330 (N_5330,N_5212,N_5103);
and U5331 (N_5331,N_5196,N_5200);
or U5332 (N_5332,N_5196,N_5211);
and U5333 (N_5333,N_5178,N_5198);
and U5334 (N_5334,N_5167,N_5105);
nor U5335 (N_5335,N_5178,N_5118);
or U5336 (N_5336,N_5244,N_5121);
xor U5337 (N_5337,N_5134,N_5138);
and U5338 (N_5338,N_5157,N_5207);
and U5339 (N_5339,N_5224,N_5209);
nor U5340 (N_5340,N_5234,N_5188);
or U5341 (N_5341,N_5221,N_5125);
and U5342 (N_5342,N_5213,N_5247);
nor U5343 (N_5343,N_5226,N_5187);
nor U5344 (N_5344,N_5139,N_5123);
and U5345 (N_5345,N_5170,N_5246);
nor U5346 (N_5346,N_5185,N_5126);
and U5347 (N_5347,N_5133,N_5100);
or U5348 (N_5348,N_5115,N_5199);
nand U5349 (N_5349,N_5213,N_5128);
or U5350 (N_5350,N_5105,N_5130);
or U5351 (N_5351,N_5233,N_5155);
nor U5352 (N_5352,N_5183,N_5137);
nor U5353 (N_5353,N_5228,N_5189);
nand U5354 (N_5354,N_5167,N_5245);
nor U5355 (N_5355,N_5131,N_5136);
and U5356 (N_5356,N_5223,N_5113);
or U5357 (N_5357,N_5176,N_5216);
nor U5358 (N_5358,N_5177,N_5180);
xnor U5359 (N_5359,N_5127,N_5149);
and U5360 (N_5360,N_5201,N_5158);
and U5361 (N_5361,N_5107,N_5172);
or U5362 (N_5362,N_5203,N_5217);
nor U5363 (N_5363,N_5160,N_5114);
and U5364 (N_5364,N_5248,N_5227);
and U5365 (N_5365,N_5106,N_5134);
nor U5366 (N_5366,N_5106,N_5119);
nand U5367 (N_5367,N_5211,N_5110);
and U5368 (N_5368,N_5110,N_5154);
nand U5369 (N_5369,N_5199,N_5122);
nand U5370 (N_5370,N_5102,N_5188);
nor U5371 (N_5371,N_5141,N_5138);
xor U5372 (N_5372,N_5230,N_5163);
or U5373 (N_5373,N_5175,N_5242);
nor U5374 (N_5374,N_5238,N_5148);
or U5375 (N_5375,N_5183,N_5196);
or U5376 (N_5376,N_5201,N_5249);
and U5377 (N_5377,N_5108,N_5236);
or U5378 (N_5378,N_5140,N_5244);
or U5379 (N_5379,N_5138,N_5151);
nor U5380 (N_5380,N_5149,N_5161);
nor U5381 (N_5381,N_5164,N_5109);
or U5382 (N_5382,N_5104,N_5212);
or U5383 (N_5383,N_5189,N_5221);
and U5384 (N_5384,N_5187,N_5176);
and U5385 (N_5385,N_5220,N_5138);
nand U5386 (N_5386,N_5167,N_5101);
nand U5387 (N_5387,N_5203,N_5226);
or U5388 (N_5388,N_5248,N_5170);
nand U5389 (N_5389,N_5121,N_5162);
nand U5390 (N_5390,N_5130,N_5119);
nor U5391 (N_5391,N_5247,N_5186);
and U5392 (N_5392,N_5106,N_5139);
and U5393 (N_5393,N_5140,N_5152);
nor U5394 (N_5394,N_5210,N_5180);
or U5395 (N_5395,N_5135,N_5229);
and U5396 (N_5396,N_5138,N_5148);
nand U5397 (N_5397,N_5237,N_5100);
nor U5398 (N_5398,N_5122,N_5200);
nor U5399 (N_5399,N_5139,N_5144);
nand U5400 (N_5400,N_5387,N_5271);
or U5401 (N_5401,N_5377,N_5283);
xnor U5402 (N_5402,N_5267,N_5323);
nand U5403 (N_5403,N_5311,N_5365);
nor U5404 (N_5404,N_5253,N_5298);
nand U5405 (N_5405,N_5361,N_5368);
or U5406 (N_5406,N_5312,N_5362);
nand U5407 (N_5407,N_5356,N_5299);
nand U5408 (N_5408,N_5282,N_5303);
nor U5409 (N_5409,N_5364,N_5342);
or U5410 (N_5410,N_5250,N_5397);
nor U5411 (N_5411,N_5346,N_5383);
nor U5412 (N_5412,N_5294,N_5395);
or U5413 (N_5413,N_5334,N_5372);
nor U5414 (N_5414,N_5354,N_5319);
and U5415 (N_5415,N_5370,N_5369);
and U5416 (N_5416,N_5349,N_5313);
xor U5417 (N_5417,N_5310,N_5359);
or U5418 (N_5418,N_5269,N_5272);
nor U5419 (N_5419,N_5251,N_5281);
and U5420 (N_5420,N_5351,N_5285);
and U5421 (N_5421,N_5261,N_5392);
and U5422 (N_5422,N_5328,N_5270);
or U5423 (N_5423,N_5286,N_5389);
or U5424 (N_5424,N_5266,N_5398);
or U5425 (N_5425,N_5284,N_5339);
nor U5426 (N_5426,N_5264,N_5393);
nand U5427 (N_5427,N_5347,N_5260);
nand U5428 (N_5428,N_5278,N_5329);
or U5429 (N_5429,N_5341,N_5382);
and U5430 (N_5430,N_5338,N_5336);
or U5431 (N_5431,N_5288,N_5390);
and U5432 (N_5432,N_5366,N_5348);
or U5433 (N_5433,N_5296,N_5308);
or U5434 (N_5434,N_5274,N_5321);
xor U5435 (N_5435,N_5304,N_5381);
nor U5436 (N_5436,N_5316,N_5376);
nand U5437 (N_5437,N_5279,N_5344);
or U5438 (N_5438,N_5293,N_5324);
and U5439 (N_5439,N_5394,N_5378);
xnor U5440 (N_5440,N_5315,N_5326);
or U5441 (N_5441,N_5275,N_5391);
nand U5442 (N_5442,N_5340,N_5355);
nand U5443 (N_5443,N_5302,N_5384);
xnor U5444 (N_5444,N_5259,N_5314);
nand U5445 (N_5445,N_5327,N_5337);
nand U5446 (N_5446,N_5325,N_5371);
or U5447 (N_5447,N_5380,N_5295);
nand U5448 (N_5448,N_5345,N_5320);
nor U5449 (N_5449,N_5289,N_5396);
nor U5450 (N_5450,N_5335,N_5252);
or U5451 (N_5451,N_5258,N_5357);
nor U5452 (N_5452,N_5290,N_5276);
nand U5453 (N_5453,N_5363,N_5352);
and U5454 (N_5454,N_5385,N_5291);
nor U5455 (N_5455,N_5254,N_5255);
and U5456 (N_5456,N_5306,N_5263);
or U5457 (N_5457,N_5300,N_5386);
nor U5458 (N_5458,N_5265,N_5256);
or U5459 (N_5459,N_5367,N_5331);
and U5460 (N_5460,N_5353,N_5307);
or U5461 (N_5461,N_5374,N_5280);
nand U5462 (N_5462,N_5257,N_5297);
xnor U5463 (N_5463,N_5273,N_5375);
nor U5464 (N_5464,N_5309,N_5379);
nand U5465 (N_5465,N_5301,N_5292);
and U5466 (N_5466,N_5399,N_5322);
or U5467 (N_5467,N_5360,N_5332);
or U5468 (N_5468,N_5268,N_5343);
and U5469 (N_5469,N_5277,N_5388);
nand U5470 (N_5470,N_5318,N_5358);
nor U5471 (N_5471,N_5287,N_5373);
nor U5472 (N_5472,N_5317,N_5350);
nor U5473 (N_5473,N_5330,N_5305);
xor U5474 (N_5474,N_5262,N_5333);
and U5475 (N_5475,N_5269,N_5395);
or U5476 (N_5476,N_5393,N_5289);
nor U5477 (N_5477,N_5283,N_5321);
and U5478 (N_5478,N_5291,N_5311);
nor U5479 (N_5479,N_5367,N_5323);
and U5480 (N_5480,N_5322,N_5256);
nor U5481 (N_5481,N_5271,N_5372);
and U5482 (N_5482,N_5397,N_5399);
nor U5483 (N_5483,N_5361,N_5262);
or U5484 (N_5484,N_5371,N_5340);
nor U5485 (N_5485,N_5285,N_5303);
or U5486 (N_5486,N_5335,N_5373);
or U5487 (N_5487,N_5358,N_5377);
nor U5488 (N_5488,N_5363,N_5305);
or U5489 (N_5489,N_5396,N_5266);
nor U5490 (N_5490,N_5326,N_5298);
nand U5491 (N_5491,N_5325,N_5297);
nor U5492 (N_5492,N_5345,N_5318);
xnor U5493 (N_5493,N_5325,N_5295);
nand U5494 (N_5494,N_5291,N_5271);
or U5495 (N_5495,N_5356,N_5376);
or U5496 (N_5496,N_5265,N_5358);
xnor U5497 (N_5497,N_5287,N_5258);
xor U5498 (N_5498,N_5301,N_5382);
nand U5499 (N_5499,N_5254,N_5346);
and U5500 (N_5500,N_5384,N_5275);
and U5501 (N_5501,N_5279,N_5296);
nor U5502 (N_5502,N_5261,N_5292);
xor U5503 (N_5503,N_5363,N_5303);
or U5504 (N_5504,N_5260,N_5266);
nor U5505 (N_5505,N_5362,N_5364);
and U5506 (N_5506,N_5330,N_5361);
nor U5507 (N_5507,N_5350,N_5364);
xnor U5508 (N_5508,N_5393,N_5356);
or U5509 (N_5509,N_5311,N_5270);
nand U5510 (N_5510,N_5308,N_5305);
and U5511 (N_5511,N_5324,N_5365);
nand U5512 (N_5512,N_5292,N_5306);
and U5513 (N_5513,N_5397,N_5251);
nor U5514 (N_5514,N_5319,N_5350);
and U5515 (N_5515,N_5327,N_5280);
nand U5516 (N_5516,N_5276,N_5304);
nand U5517 (N_5517,N_5261,N_5255);
nand U5518 (N_5518,N_5285,N_5305);
and U5519 (N_5519,N_5367,N_5262);
nor U5520 (N_5520,N_5356,N_5276);
nor U5521 (N_5521,N_5372,N_5367);
nor U5522 (N_5522,N_5262,N_5353);
nor U5523 (N_5523,N_5321,N_5392);
or U5524 (N_5524,N_5328,N_5317);
nand U5525 (N_5525,N_5318,N_5301);
and U5526 (N_5526,N_5379,N_5347);
and U5527 (N_5527,N_5266,N_5355);
or U5528 (N_5528,N_5399,N_5293);
xnor U5529 (N_5529,N_5307,N_5334);
and U5530 (N_5530,N_5287,N_5363);
nor U5531 (N_5531,N_5389,N_5285);
nor U5532 (N_5532,N_5349,N_5336);
xor U5533 (N_5533,N_5349,N_5352);
or U5534 (N_5534,N_5312,N_5388);
nor U5535 (N_5535,N_5349,N_5396);
nand U5536 (N_5536,N_5287,N_5273);
and U5537 (N_5537,N_5260,N_5295);
and U5538 (N_5538,N_5295,N_5299);
or U5539 (N_5539,N_5272,N_5357);
and U5540 (N_5540,N_5264,N_5296);
nor U5541 (N_5541,N_5323,N_5329);
nor U5542 (N_5542,N_5326,N_5310);
nand U5543 (N_5543,N_5338,N_5335);
nor U5544 (N_5544,N_5272,N_5373);
and U5545 (N_5545,N_5358,N_5395);
or U5546 (N_5546,N_5370,N_5296);
xnor U5547 (N_5547,N_5319,N_5334);
nand U5548 (N_5548,N_5278,N_5385);
nand U5549 (N_5549,N_5258,N_5304);
and U5550 (N_5550,N_5534,N_5521);
xor U5551 (N_5551,N_5533,N_5491);
or U5552 (N_5552,N_5469,N_5514);
nor U5553 (N_5553,N_5421,N_5535);
and U5554 (N_5554,N_5466,N_5408);
xor U5555 (N_5555,N_5538,N_5516);
nand U5556 (N_5556,N_5510,N_5442);
and U5557 (N_5557,N_5423,N_5477);
nor U5558 (N_5558,N_5523,N_5415);
nand U5559 (N_5559,N_5494,N_5458);
or U5560 (N_5560,N_5409,N_5471);
or U5561 (N_5561,N_5508,N_5441);
or U5562 (N_5562,N_5498,N_5512);
or U5563 (N_5563,N_5457,N_5537);
or U5564 (N_5564,N_5492,N_5479);
and U5565 (N_5565,N_5518,N_5400);
nor U5566 (N_5566,N_5539,N_5414);
nand U5567 (N_5567,N_5517,N_5402);
or U5568 (N_5568,N_5502,N_5520);
or U5569 (N_5569,N_5434,N_5424);
nand U5570 (N_5570,N_5536,N_5447);
nand U5571 (N_5571,N_5459,N_5543);
nor U5572 (N_5572,N_5440,N_5485);
nor U5573 (N_5573,N_5481,N_5496);
nand U5574 (N_5574,N_5425,N_5401);
and U5575 (N_5575,N_5515,N_5405);
or U5576 (N_5576,N_5450,N_5433);
and U5577 (N_5577,N_5451,N_5422);
and U5578 (N_5578,N_5542,N_5439);
and U5579 (N_5579,N_5495,N_5449);
or U5580 (N_5580,N_5476,N_5429);
nor U5581 (N_5581,N_5541,N_5475);
nand U5582 (N_5582,N_5513,N_5482);
nor U5583 (N_5583,N_5407,N_5546);
or U5584 (N_5584,N_5505,N_5468);
nor U5585 (N_5585,N_5488,N_5437);
nor U5586 (N_5586,N_5493,N_5427);
and U5587 (N_5587,N_5460,N_5549);
nor U5588 (N_5588,N_5465,N_5464);
nand U5589 (N_5589,N_5443,N_5417);
nand U5590 (N_5590,N_5522,N_5462);
and U5591 (N_5591,N_5456,N_5487);
or U5592 (N_5592,N_5420,N_5410);
or U5593 (N_5593,N_5411,N_5444);
nand U5594 (N_5594,N_5431,N_5467);
nand U5595 (N_5595,N_5438,N_5470);
and U5596 (N_5596,N_5501,N_5540);
nand U5597 (N_5597,N_5529,N_5430);
nand U5598 (N_5598,N_5484,N_5473);
and U5599 (N_5599,N_5524,N_5412);
and U5600 (N_5600,N_5432,N_5454);
and U5601 (N_5601,N_5530,N_5499);
or U5602 (N_5602,N_5486,N_5503);
and U5603 (N_5603,N_5445,N_5506);
and U5604 (N_5604,N_5504,N_5497);
nand U5605 (N_5605,N_5419,N_5413);
nor U5606 (N_5606,N_5547,N_5448);
or U5607 (N_5607,N_5507,N_5483);
and U5608 (N_5608,N_5418,N_5472);
nor U5609 (N_5609,N_5463,N_5452);
nor U5610 (N_5610,N_5525,N_5490);
nor U5611 (N_5611,N_5480,N_5531);
xnor U5612 (N_5612,N_5404,N_5500);
nand U5613 (N_5613,N_5509,N_5527);
or U5614 (N_5614,N_5455,N_5416);
or U5615 (N_5615,N_5519,N_5478);
or U5616 (N_5616,N_5428,N_5453);
or U5617 (N_5617,N_5474,N_5435);
or U5618 (N_5618,N_5528,N_5544);
xor U5619 (N_5619,N_5489,N_5532);
nor U5620 (N_5620,N_5511,N_5406);
nand U5621 (N_5621,N_5446,N_5403);
nand U5622 (N_5622,N_5436,N_5426);
nand U5623 (N_5623,N_5548,N_5526);
xnor U5624 (N_5624,N_5461,N_5545);
nor U5625 (N_5625,N_5457,N_5425);
xor U5626 (N_5626,N_5476,N_5546);
nor U5627 (N_5627,N_5510,N_5502);
nor U5628 (N_5628,N_5454,N_5468);
and U5629 (N_5629,N_5501,N_5478);
nand U5630 (N_5630,N_5465,N_5423);
nand U5631 (N_5631,N_5404,N_5524);
nand U5632 (N_5632,N_5526,N_5497);
or U5633 (N_5633,N_5534,N_5465);
xor U5634 (N_5634,N_5463,N_5524);
nor U5635 (N_5635,N_5418,N_5519);
nand U5636 (N_5636,N_5412,N_5543);
or U5637 (N_5637,N_5467,N_5543);
nor U5638 (N_5638,N_5524,N_5425);
nor U5639 (N_5639,N_5520,N_5535);
and U5640 (N_5640,N_5494,N_5425);
nor U5641 (N_5641,N_5533,N_5440);
or U5642 (N_5642,N_5479,N_5429);
nor U5643 (N_5643,N_5472,N_5512);
nor U5644 (N_5644,N_5425,N_5441);
xnor U5645 (N_5645,N_5461,N_5482);
and U5646 (N_5646,N_5536,N_5517);
and U5647 (N_5647,N_5490,N_5518);
nand U5648 (N_5648,N_5530,N_5472);
nand U5649 (N_5649,N_5402,N_5539);
nor U5650 (N_5650,N_5497,N_5420);
and U5651 (N_5651,N_5544,N_5498);
or U5652 (N_5652,N_5493,N_5510);
nor U5653 (N_5653,N_5463,N_5475);
nor U5654 (N_5654,N_5434,N_5534);
or U5655 (N_5655,N_5459,N_5418);
nand U5656 (N_5656,N_5402,N_5442);
or U5657 (N_5657,N_5543,N_5507);
or U5658 (N_5658,N_5509,N_5534);
nand U5659 (N_5659,N_5517,N_5433);
nor U5660 (N_5660,N_5534,N_5482);
nand U5661 (N_5661,N_5547,N_5476);
nand U5662 (N_5662,N_5457,N_5449);
nor U5663 (N_5663,N_5408,N_5529);
nor U5664 (N_5664,N_5444,N_5463);
or U5665 (N_5665,N_5430,N_5471);
nor U5666 (N_5666,N_5429,N_5439);
and U5667 (N_5667,N_5435,N_5546);
nand U5668 (N_5668,N_5504,N_5549);
and U5669 (N_5669,N_5486,N_5430);
nand U5670 (N_5670,N_5499,N_5442);
and U5671 (N_5671,N_5463,N_5488);
xnor U5672 (N_5672,N_5461,N_5449);
and U5673 (N_5673,N_5547,N_5533);
and U5674 (N_5674,N_5534,N_5460);
nor U5675 (N_5675,N_5459,N_5426);
and U5676 (N_5676,N_5414,N_5522);
nand U5677 (N_5677,N_5526,N_5520);
nand U5678 (N_5678,N_5462,N_5489);
and U5679 (N_5679,N_5435,N_5493);
nor U5680 (N_5680,N_5402,N_5441);
nor U5681 (N_5681,N_5460,N_5418);
nand U5682 (N_5682,N_5496,N_5445);
and U5683 (N_5683,N_5439,N_5410);
or U5684 (N_5684,N_5540,N_5419);
or U5685 (N_5685,N_5453,N_5482);
nand U5686 (N_5686,N_5471,N_5470);
and U5687 (N_5687,N_5416,N_5447);
or U5688 (N_5688,N_5448,N_5490);
or U5689 (N_5689,N_5470,N_5528);
and U5690 (N_5690,N_5547,N_5434);
nand U5691 (N_5691,N_5537,N_5543);
nor U5692 (N_5692,N_5417,N_5493);
and U5693 (N_5693,N_5482,N_5492);
or U5694 (N_5694,N_5514,N_5526);
nand U5695 (N_5695,N_5452,N_5548);
or U5696 (N_5696,N_5539,N_5449);
nor U5697 (N_5697,N_5548,N_5519);
nand U5698 (N_5698,N_5480,N_5514);
nor U5699 (N_5699,N_5527,N_5492);
nor U5700 (N_5700,N_5683,N_5672);
nand U5701 (N_5701,N_5615,N_5613);
nand U5702 (N_5702,N_5693,N_5561);
xor U5703 (N_5703,N_5639,N_5697);
and U5704 (N_5704,N_5645,N_5653);
and U5705 (N_5705,N_5658,N_5643);
and U5706 (N_5706,N_5612,N_5650);
or U5707 (N_5707,N_5644,N_5629);
or U5708 (N_5708,N_5624,N_5573);
nor U5709 (N_5709,N_5553,N_5620);
xor U5710 (N_5710,N_5619,N_5638);
nand U5711 (N_5711,N_5649,N_5616);
or U5712 (N_5712,N_5609,N_5668);
and U5713 (N_5713,N_5567,N_5592);
nand U5714 (N_5714,N_5679,N_5669);
or U5715 (N_5715,N_5604,N_5694);
nand U5716 (N_5716,N_5552,N_5642);
and U5717 (N_5717,N_5593,N_5621);
or U5718 (N_5718,N_5654,N_5578);
nand U5719 (N_5719,N_5577,N_5602);
nor U5720 (N_5720,N_5594,N_5635);
and U5721 (N_5721,N_5684,N_5662);
nand U5722 (N_5722,N_5617,N_5631);
or U5723 (N_5723,N_5681,N_5647);
nand U5724 (N_5724,N_5574,N_5560);
nor U5725 (N_5725,N_5584,N_5640);
nor U5726 (N_5726,N_5607,N_5557);
nand U5727 (N_5727,N_5663,N_5588);
or U5728 (N_5728,N_5603,N_5698);
nor U5729 (N_5729,N_5575,N_5636);
xnor U5730 (N_5730,N_5692,N_5570);
and U5731 (N_5731,N_5565,N_5680);
nand U5732 (N_5732,N_5652,N_5656);
nor U5733 (N_5733,N_5589,N_5626);
and U5734 (N_5734,N_5558,N_5661);
nand U5735 (N_5735,N_5586,N_5676);
and U5736 (N_5736,N_5559,N_5597);
and U5737 (N_5737,N_5579,N_5699);
nand U5738 (N_5738,N_5600,N_5687);
nor U5739 (N_5739,N_5641,N_5655);
nor U5740 (N_5740,N_5566,N_5571);
and U5741 (N_5741,N_5611,N_5587);
nand U5742 (N_5742,N_5685,N_5550);
and U5743 (N_5743,N_5627,N_5666);
nor U5744 (N_5744,N_5595,N_5630);
and U5745 (N_5745,N_5606,N_5674);
nor U5746 (N_5746,N_5696,N_5551);
nand U5747 (N_5747,N_5665,N_5688);
nand U5748 (N_5748,N_5686,N_5648);
nand U5749 (N_5749,N_5610,N_5695);
xnor U5750 (N_5750,N_5625,N_5614);
nand U5751 (N_5751,N_5601,N_5618);
xnor U5752 (N_5752,N_5660,N_5596);
nor U5753 (N_5753,N_5576,N_5632);
nor U5754 (N_5754,N_5637,N_5634);
nor U5755 (N_5755,N_5556,N_5582);
or U5756 (N_5756,N_5568,N_5673);
xnor U5757 (N_5757,N_5623,N_5562);
or U5758 (N_5758,N_5691,N_5583);
xor U5759 (N_5759,N_5628,N_5690);
nand U5760 (N_5760,N_5678,N_5667);
and U5761 (N_5761,N_5555,N_5633);
nor U5762 (N_5762,N_5572,N_5599);
nand U5763 (N_5763,N_5569,N_5622);
nand U5764 (N_5764,N_5598,N_5659);
xor U5765 (N_5765,N_5651,N_5646);
or U5766 (N_5766,N_5677,N_5671);
nor U5767 (N_5767,N_5564,N_5590);
nor U5768 (N_5768,N_5664,N_5689);
nor U5769 (N_5769,N_5682,N_5675);
nor U5770 (N_5770,N_5554,N_5585);
nor U5771 (N_5771,N_5591,N_5670);
xor U5772 (N_5772,N_5581,N_5657);
and U5773 (N_5773,N_5605,N_5580);
nand U5774 (N_5774,N_5608,N_5563);
and U5775 (N_5775,N_5573,N_5668);
nand U5776 (N_5776,N_5674,N_5569);
or U5777 (N_5777,N_5685,N_5589);
and U5778 (N_5778,N_5667,N_5580);
nand U5779 (N_5779,N_5593,N_5658);
xnor U5780 (N_5780,N_5662,N_5590);
or U5781 (N_5781,N_5577,N_5668);
and U5782 (N_5782,N_5678,N_5672);
xnor U5783 (N_5783,N_5690,N_5580);
or U5784 (N_5784,N_5566,N_5599);
or U5785 (N_5785,N_5653,N_5678);
nor U5786 (N_5786,N_5556,N_5578);
nor U5787 (N_5787,N_5672,N_5594);
nor U5788 (N_5788,N_5683,N_5550);
and U5789 (N_5789,N_5678,N_5694);
or U5790 (N_5790,N_5576,N_5623);
or U5791 (N_5791,N_5582,N_5639);
and U5792 (N_5792,N_5654,N_5601);
and U5793 (N_5793,N_5647,N_5568);
nand U5794 (N_5794,N_5621,N_5635);
and U5795 (N_5795,N_5690,N_5574);
or U5796 (N_5796,N_5609,N_5696);
nor U5797 (N_5797,N_5668,N_5633);
or U5798 (N_5798,N_5634,N_5585);
xnor U5799 (N_5799,N_5668,N_5688);
or U5800 (N_5800,N_5578,N_5599);
or U5801 (N_5801,N_5579,N_5693);
or U5802 (N_5802,N_5565,N_5641);
nor U5803 (N_5803,N_5620,N_5673);
nor U5804 (N_5804,N_5642,N_5576);
xor U5805 (N_5805,N_5582,N_5619);
nor U5806 (N_5806,N_5606,N_5694);
and U5807 (N_5807,N_5573,N_5629);
nor U5808 (N_5808,N_5681,N_5636);
or U5809 (N_5809,N_5688,N_5552);
nor U5810 (N_5810,N_5580,N_5666);
and U5811 (N_5811,N_5602,N_5642);
nor U5812 (N_5812,N_5563,N_5561);
and U5813 (N_5813,N_5662,N_5682);
xnor U5814 (N_5814,N_5584,N_5683);
and U5815 (N_5815,N_5655,N_5627);
and U5816 (N_5816,N_5662,N_5699);
or U5817 (N_5817,N_5576,N_5635);
nand U5818 (N_5818,N_5684,N_5572);
nand U5819 (N_5819,N_5692,N_5664);
xnor U5820 (N_5820,N_5642,N_5659);
and U5821 (N_5821,N_5574,N_5646);
nand U5822 (N_5822,N_5550,N_5629);
nand U5823 (N_5823,N_5611,N_5616);
nand U5824 (N_5824,N_5592,N_5663);
and U5825 (N_5825,N_5645,N_5598);
nor U5826 (N_5826,N_5675,N_5570);
and U5827 (N_5827,N_5673,N_5572);
nand U5828 (N_5828,N_5681,N_5635);
and U5829 (N_5829,N_5583,N_5618);
nand U5830 (N_5830,N_5606,N_5568);
nor U5831 (N_5831,N_5567,N_5575);
nand U5832 (N_5832,N_5585,N_5572);
nor U5833 (N_5833,N_5652,N_5642);
or U5834 (N_5834,N_5572,N_5574);
and U5835 (N_5835,N_5585,N_5627);
and U5836 (N_5836,N_5579,N_5611);
or U5837 (N_5837,N_5683,N_5654);
or U5838 (N_5838,N_5611,N_5697);
nor U5839 (N_5839,N_5622,N_5631);
nand U5840 (N_5840,N_5627,N_5634);
nand U5841 (N_5841,N_5639,N_5657);
nor U5842 (N_5842,N_5607,N_5698);
xor U5843 (N_5843,N_5698,N_5658);
nor U5844 (N_5844,N_5668,N_5561);
and U5845 (N_5845,N_5693,N_5553);
nand U5846 (N_5846,N_5635,N_5578);
or U5847 (N_5847,N_5640,N_5682);
nor U5848 (N_5848,N_5561,N_5648);
nor U5849 (N_5849,N_5608,N_5615);
xor U5850 (N_5850,N_5708,N_5756);
and U5851 (N_5851,N_5822,N_5700);
nand U5852 (N_5852,N_5770,N_5796);
and U5853 (N_5853,N_5775,N_5765);
and U5854 (N_5854,N_5815,N_5758);
or U5855 (N_5855,N_5714,N_5736);
nor U5856 (N_5856,N_5723,N_5799);
or U5857 (N_5857,N_5771,N_5838);
nor U5858 (N_5858,N_5798,N_5840);
nor U5859 (N_5859,N_5819,N_5841);
and U5860 (N_5860,N_5707,N_5810);
nand U5861 (N_5861,N_5839,N_5788);
nor U5862 (N_5862,N_5833,N_5829);
xor U5863 (N_5863,N_5722,N_5844);
nand U5864 (N_5864,N_5849,N_5706);
nor U5865 (N_5865,N_5746,N_5814);
xnor U5866 (N_5866,N_5789,N_5848);
xnor U5867 (N_5867,N_5767,N_5701);
or U5868 (N_5868,N_5808,N_5741);
nor U5869 (N_5869,N_5715,N_5759);
nand U5870 (N_5870,N_5824,N_5845);
or U5871 (N_5871,N_5793,N_5740);
nor U5872 (N_5872,N_5735,N_5742);
or U5873 (N_5873,N_5817,N_5787);
and U5874 (N_5874,N_5768,N_5782);
xnor U5875 (N_5875,N_5769,N_5745);
or U5876 (N_5876,N_5725,N_5813);
xnor U5877 (N_5877,N_5794,N_5826);
nor U5878 (N_5878,N_5761,N_5842);
nand U5879 (N_5879,N_5760,N_5751);
nor U5880 (N_5880,N_5801,N_5785);
nor U5881 (N_5881,N_5713,N_5755);
and U5882 (N_5882,N_5710,N_5816);
or U5883 (N_5883,N_5802,N_5831);
and U5884 (N_5884,N_5795,N_5752);
nor U5885 (N_5885,N_5730,N_5704);
nand U5886 (N_5886,N_5772,N_5743);
nor U5887 (N_5887,N_5781,N_5712);
nand U5888 (N_5888,N_5747,N_5830);
and U5889 (N_5889,N_5820,N_5776);
nand U5890 (N_5890,N_5780,N_5719);
nor U5891 (N_5891,N_5800,N_5703);
and U5892 (N_5892,N_5702,N_5731);
and U5893 (N_5893,N_5727,N_5717);
nand U5894 (N_5894,N_5728,N_5726);
or U5895 (N_5895,N_5753,N_5846);
nand U5896 (N_5896,N_5748,N_5807);
nand U5897 (N_5897,N_5709,N_5729);
or U5898 (N_5898,N_5716,N_5737);
and U5899 (N_5899,N_5827,N_5818);
and U5900 (N_5900,N_5809,N_5754);
and U5901 (N_5901,N_5783,N_5744);
or U5902 (N_5902,N_5757,N_5811);
nand U5903 (N_5903,N_5773,N_5835);
or U5904 (N_5904,N_5721,N_5705);
nand U5905 (N_5905,N_5791,N_5790);
nand U5906 (N_5906,N_5738,N_5784);
xnor U5907 (N_5907,N_5832,N_5732);
and U5908 (N_5908,N_5797,N_5804);
and U5909 (N_5909,N_5779,N_5750);
nand U5910 (N_5910,N_5792,N_5764);
nor U5911 (N_5911,N_5763,N_5823);
nor U5912 (N_5912,N_5766,N_5720);
nand U5913 (N_5913,N_5825,N_5733);
nor U5914 (N_5914,N_5718,N_5828);
nand U5915 (N_5915,N_5762,N_5786);
or U5916 (N_5916,N_5777,N_5821);
nor U5917 (N_5917,N_5805,N_5803);
or U5918 (N_5918,N_5724,N_5834);
nor U5919 (N_5919,N_5734,N_5836);
nand U5920 (N_5920,N_5843,N_5711);
and U5921 (N_5921,N_5847,N_5778);
nor U5922 (N_5922,N_5739,N_5806);
nand U5923 (N_5923,N_5812,N_5774);
xor U5924 (N_5924,N_5837,N_5749);
nor U5925 (N_5925,N_5847,N_5720);
xnor U5926 (N_5926,N_5740,N_5739);
and U5927 (N_5927,N_5796,N_5785);
nand U5928 (N_5928,N_5837,N_5722);
or U5929 (N_5929,N_5802,N_5755);
nor U5930 (N_5930,N_5828,N_5762);
or U5931 (N_5931,N_5789,N_5773);
nand U5932 (N_5932,N_5848,N_5707);
and U5933 (N_5933,N_5786,N_5757);
or U5934 (N_5934,N_5784,N_5817);
or U5935 (N_5935,N_5823,N_5729);
or U5936 (N_5936,N_5717,N_5821);
or U5937 (N_5937,N_5793,N_5775);
and U5938 (N_5938,N_5847,N_5817);
and U5939 (N_5939,N_5781,N_5721);
nor U5940 (N_5940,N_5834,N_5787);
nand U5941 (N_5941,N_5735,N_5839);
xor U5942 (N_5942,N_5802,N_5709);
nand U5943 (N_5943,N_5814,N_5719);
or U5944 (N_5944,N_5808,N_5742);
or U5945 (N_5945,N_5820,N_5849);
nor U5946 (N_5946,N_5798,N_5721);
or U5947 (N_5947,N_5713,N_5813);
nand U5948 (N_5948,N_5769,N_5770);
nor U5949 (N_5949,N_5840,N_5770);
and U5950 (N_5950,N_5772,N_5776);
nand U5951 (N_5951,N_5800,N_5753);
and U5952 (N_5952,N_5826,N_5778);
and U5953 (N_5953,N_5781,N_5799);
or U5954 (N_5954,N_5756,N_5788);
xnor U5955 (N_5955,N_5749,N_5786);
nand U5956 (N_5956,N_5830,N_5751);
nor U5957 (N_5957,N_5831,N_5790);
nand U5958 (N_5958,N_5808,N_5809);
nand U5959 (N_5959,N_5723,N_5793);
nor U5960 (N_5960,N_5838,N_5764);
or U5961 (N_5961,N_5804,N_5815);
or U5962 (N_5962,N_5814,N_5709);
and U5963 (N_5963,N_5790,N_5752);
and U5964 (N_5964,N_5773,N_5733);
nand U5965 (N_5965,N_5782,N_5823);
nand U5966 (N_5966,N_5721,N_5767);
or U5967 (N_5967,N_5841,N_5758);
and U5968 (N_5968,N_5717,N_5723);
xnor U5969 (N_5969,N_5729,N_5716);
and U5970 (N_5970,N_5809,N_5748);
xnor U5971 (N_5971,N_5714,N_5742);
nor U5972 (N_5972,N_5796,N_5840);
nor U5973 (N_5973,N_5841,N_5721);
nor U5974 (N_5974,N_5766,N_5742);
xor U5975 (N_5975,N_5770,N_5764);
nand U5976 (N_5976,N_5746,N_5809);
xor U5977 (N_5977,N_5703,N_5839);
and U5978 (N_5978,N_5705,N_5725);
or U5979 (N_5979,N_5713,N_5848);
or U5980 (N_5980,N_5704,N_5802);
and U5981 (N_5981,N_5832,N_5745);
xnor U5982 (N_5982,N_5825,N_5739);
nand U5983 (N_5983,N_5841,N_5815);
or U5984 (N_5984,N_5835,N_5811);
nor U5985 (N_5985,N_5808,N_5714);
nor U5986 (N_5986,N_5775,N_5828);
nor U5987 (N_5987,N_5754,N_5813);
or U5988 (N_5988,N_5728,N_5720);
and U5989 (N_5989,N_5764,N_5760);
or U5990 (N_5990,N_5844,N_5784);
nand U5991 (N_5991,N_5729,N_5827);
nand U5992 (N_5992,N_5729,N_5708);
nor U5993 (N_5993,N_5787,N_5816);
and U5994 (N_5994,N_5816,N_5707);
xnor U5995 (N_5995,N_5703,N_5844);
and U5996 (N_5996,N_5803,N_5802);
or U5997 (N_5997,N_5736,N_5755);
nor U5998 (N_5998,N_5711,N_5785);
xor U5999 (N_5999,N_5727,N_5744);
nor U6000 (N_6000,N_5882,N_5992);
nor U6001 (N_6001,N_5908,N_5940);
and U6002 (N_6002,N_5968,N_5924);
nand U6003 (N_6003,N_5974,N_5887);
and U6004 (N_6004,N_5881,N_5872);
or U6005 (N_6005,N_5931,N_5930);
and U6006 (N_6006,N_5892,N_5921);
nor U6007 (N_6007,N_5987,N_5942);
nand U6008 (N_6008,N_5963,N_5912);
xnor U6009 (N_6009,N_5964,N_5855);
nor U6010 (N_6010,N_5856,N_5946);
or U6011 (N_6011,N_5989,N_5876);
nand U6012 (N_6012,N_5959,N_5917);
nand U6013 (N_6013,N_5919,N_5995);
and U6014 (N_6014,N_5975,N_5851);
nor U6015 (N_6015,N_5898,N_5877);
xor U6016 (N_6016,N_5867,N_5860);
xnor U6017 (N_6017,N_5865,N_5884);
nand U6018 (N_6018,N_5941,N_5988);
and U6019 (N_6019,N_5864,N_5936);
or U6020 (N_6020,N_5896,N_5944);
xnor U6021 (N_6021,N_5994,N_5868);
or U6022 (N_6022,N_5910,N_5949);
or U6023 (N_6023,N_5880,N_5971);
nand U6024 (N_6024,N_5926,N_5967);
nand U6025 (N_6025,N_5991,N_5945);
or U6026 (N_6026,N_5899,N_5960);
nor U6027 (N_6027,N_5857,N_5888);
nor U6028 (N_6028,N_5873,N_5979);
xnor U6029 (N_6029,N_5970,N_5958);
and U6030 (N_6030,N_5871,N_5937);
nand U6031 (N_6031,N_5999,N_5969);
nor U6032 (N_6032,N_5920,N_5886);
nand U6033 (N_6033,N_5966,N_5853);
or U6034 (N_6034,N_5905,N_5980);
or U6035 (N_6035,N_5933,N_5986);
nand U6036 (N_6036,N_5938,N_5874);
xnor U6037 (N_6037,N_5883,N_5918);
nor U6038 (N_6038,N_5914,N_5976);
xor U6039 (N_6039,N_5934,N_5906);
nor U6040 (N_6040,N_5947,N_5913);
nor U6041 (N_6041,N_5978,N_5925);
nor U6042 (N_6042,N_5911,N_5904);
xor U6043 (N_6043,N_5928,N_5901);
nand U6044 (N_6044,N_5990,N_5977);
or U6045 (N_6045,N_5954,N_5869);
and U6046 (N_6046,N_5951,N_5965);
xor U6047 (N_6047,N_5984,N_5927);
nand U6048 (N_6048,N_5915,N_5985);
nor U6049 (N_6049,N_5955,N_5962);
and U6050 (N_6050,N_5998,N_5997);
and U6051 (N_6051,N_5953,N_5993);
nand U6052 (N_6052,N_5854,N_5903);
or U6053 (N_6053,N_5923,N_5878);
and U6054 (N_6054,N_5932,N_5922);
or U6055 (N_6055,N_5973,N_5879);
or U6056 (N_6056,N_5950,N_5858);
xor U6057 (N_6057,N_5943,N_5863);
or U6058 (N_6058,N_5866,N_5916);
nand U6059 (N_6059,N_5900,N_5957);
and U6060 (N_6060,N_5961,N_5909);
xnor U6061 (N_6061,N_5893,N_5850);
or U6062 (N_6062,N_5890,N_5929);
and U6063 (N_6063,N_5972,N_5935);
nor U6064 (N_6064,N_5870,N_5956);
nand U6065 (N_6065,N_5895,N_5862);
or U6066 (N_6066,N_5861,N_5948);
or U6067 (N_6067,N_5894,N_5891);
nand U6068 (N_6068,N_5996,N_5902);
or U6069 (N_6069,N_5983,N_5982);
or U6070 (N_6070,N_5907,N_5859);
and U6071 (N_6071,N_5885,N_5981);
nor U6072 (N_6072,N_5939,N_5889);
and U6073 (N_6073,N_5952,N_5897);
nor U6074 (N_6074,N_5852,N_5875);
or U6075 (N_6075,N_5993,N_5998);
and U6076 (N_6076,N_5996,N_5904);
nor U6077 (N_6077,N_5895,N_5910);
nand U6078 (N_6078,N_5975,N_5852);
nor U6079 (N_6079,N_5974,N_5910);
nor U6080 (N_6080,N_5922,N_5929);
and U6081 (N_6081,N_5977,N_5864);
or U6082 (N_6082,N_5890,N_5972);
nor U6083 (N_6083,N_5990,N_5980);
nor U6084 (N_6084,N_5976,N_5974);
nor U6085 (N_6085,N_5982,N_5887);
xor U6086 (N_6086,N_5862,N_5944);
xnor U6087 (N_6087,N_5995,N_5981);
nor U6088 (N_6088,N_5999,N_5966);
or U6089 (N_6089,N_5971,N_5884);
or U6090 (N_6090,N_5963,N_5923);
xor U6091 (N_6091,N_5948,N_5879);
and U6092 (N_6092,N_5969,N_5864);
nand U6093 (N_6093,N_5957,N_5929);
or U6094 (N_6094,N_5978,N_5916);
nor U6095 (N_6095,N_5954,N_5905);
and U6096 (N_6096,N_5963,N_5979);
or U6097 (N_6097,N_5898,N_5986);
nor U6098 (N_6098,N_5938,N_5980);
nor U6099 (N_6099,N_5928,N_5925);
nor U6100 (N_6100,N_5994,N_5953);
or U6101 (N_6101,N_5904,N_5903);
nor U6102 (N_6102,N_5981,N_5991);
nand U6103 (N_6103,N_5983,N_5937);
or U6104 (N_6104,N_5850,N_5906);
nor U6105 (N_6105,N_5967,N_5949);
and U6106 (N_6106,N_5930,N_5875);
nand U6107 (N_6107,N_5945,N_5957);
or U6108 (N_6108,N_5933,N_5954);
and U6109 (N_6109,N_5861,N_5955);
and U6110 (N_6110,N_5947,N_5938);
nand U6111 (N_6111,N_5949,N_5955);
or U6112 (N_6112,N_5850,N_5889);
or U6113 (N_6113,N_5853,N_5933);
and U6114 (N_6114,N_5973,N_5959);
and U6115 (N_6115,N_5854,N_5901);
or U6116 (N_6116,N_5958,N_5922);
or U6117 (N_6117,N_5912,N_5977);
nor U6118 (N_6118,N_5932,N_5865);
nand U6119 (N_6119,N_5882,N_5928);
and U6120 (N_6120,N_5988,N_5867);
nand U6121 (N_6121,N_5993,N_5996);
and U6122 (N_6122,N_5879,N_5922);
and U6123 (N_6123,N_5989,N_5861);
nor U6124 (N_6124,N_5968,N_5961);
or U6125 (N_6125,N_5876,N_5967);
or U6126 (N_6126,N_5928,N_5978);
nand U6127 (N_6127,N_5871,N_5952);
nor U6128 (N_6128,N_5968,N_5879);
nor U6129 (N_6129,N_5984,N_5982);
and U6130 (N_6130,N_5953,N_5962);
and U6131 (N_6131,N_5895,N_5900);
xor U6132 (N_6132,N_5979,N_5880);
xor U6133 (N_6133,N_5882,N_5930);
and U6134 (N_6134,N_5994,N_5947);
and U6135 (N_6135,N_5940,N_5901);
nand U6136 (N_6136,N_5962,N_5950);
nor U6137 (N_6137,N_5887,N_5883);
and U6138 (N_6138,N_5975,N_5938);
nor U6139 (N_6139,N_5955,N_5856);
nor U6140 (N_6140,N_5999,N_5881);
nand U6141 (N_6141,N_5997,N_5923);
or U6142 (N_6142,N_5893,N_5940);
or U6143 (N_6143,N_5921,N_5891);
and U6144 (N_6144,N_5922,N_5886);
and U6145 (N_6145,N_5884,N_5952);
xor U6146 (N_6146,N_5891,N_5986);
nor U6147 (N_6147,N_5879,N_5931);
nand U6148 (N_6148,N_5881,N_5948);
nand U6149 (N_6149,N_5991,N_5977);
and U6150 (N_6150,N_6133,N_6126);
nor U6151 (N_6151,N_6109,N_6018);
nor U6152 (N_6152,N_6071,N_6130);
xnor U6153 (N_6153,N_6063,N_6125);
nor U6154 (N_6154,N_6138,N_6116);
nand U6155 (N_6155,N_6056,N_6127);
and U6156 (N_6156,N_6008,N_6146);
and U6157 (N_6157,N_6122,N_6048);
nor U6158 (N_6158,N_6084,N_6068);
nand U6159 (N_6159,N_6092,N_6110);
and U6160 (N_6160,N_6097,N_6064);
or U6161 (N_6161,N_6026,N_6055);
nand U6162 (N_6162,N_6010,N_6101);
nor U6163 (N_6163,N_6104,N_6080);
nand U6164 (N_6164,N_6076,N_6085);
xnor U6165 (N_6165,N_6052,N_6147);
or U6166 (N_6166,N_6087,N_6149);
and U6167 (N_6167,N_6066,N_6070);
or U6168 (N_6168,N_6030,N_6107);
nand U6169 (N_6169,N_6021,N_6136);
nand U6170 (N_6170,N_6096,N_6102);
nand U6171 (N_6171,N_6140,N_6073);
nand U6172 (N_6172,N_6108,N_6012);
nor U6173 (N_6173,N_6114,N_6049);
nor U6174 (N_6174,N_6115,N_6001);
nand U6175 (N_6175,N_6142,N_6094);
and U6176 (N_6176,N_6007,N_6131);
and U6177 (N_6177,N_6121,N_6047);
nand U6178 (N_6178,N_6119,N_6069);
or U6179 (N_6179,N_6144,N_6006);
nand U6180 (N_6180,N_6011,N_6015);
nor U6181 (N_6181,N_6041,N_6059);
or U6182 (N_6182,N_6062,N_6013);
xor U6183 (N_6183,N_6103,N_6123);
xor U6184 (N_6184,N_6105,N_6009);
nand U6185 (N_6185,N_6022,N_6091);
nand U6186 (N_6186,N_6016,N_6032);
nand U6187 (N_6187,N_6128,N_6028);
and U6188 (N_6188,N_6072,N_6118);
or U6189 (N_6189,N_6141,N_6139);
nand U6190 (N_6190,N_6098,N_6004);
or U6191 (N_6191,N_6029,N_6078);
nor U6192 (N_6192,N_6014,N_6113);
or U6193 (N_6193,N_6095,N_6086);
or U6194 (N_6194,N_6033,N_6077);
xor U6195 (N_6195,N_6044,N_6000);
nor U6196 (N_6196,N_6117,N_6017);
and U6197 (N_6197,N_6034,N_6089);
nor U6198 (N_6198,N_6020,N_6075);
or U6199 (N_6199,N_6023,N_6019);
nor U6200 (N_6200,N_6143,N_6065);
nor U6201 (N_6201,N_6099,N_6079);
or U6202 (N_6202,N_6039,N_6035);
and U6203 (N_6203,N_6050,N_6106);
xnor U6204 (N_6204,N_6124,N_6135);
and U6205 (N_6205,N_6081,N_6025);
or U6206 (N_6206,N_6067,N_6137);
and U6207 (N_6207,N_6037,N_6074);
and U6208 (N_6208,N_6054,N_6061);
and U6209 (N_6209,N_6024,N_6088);
or U6210 (N_6210,N_6046,N_6100);
nand U6211 (N_6211,N_6132,N_6003);
and U6212 (N_6212,N_6120,N_6090);
nor U6213 (N_6213,N_6051,N_6053);
nand U6214 (N_6214,N_6111,N_6005);
nand U6215 (N_6215,N_6058,N_6134);
or U6216 (N_6216,N_6027,N_6093);
xnor U6217 (N_6217,N_6040,N_6045);
nand U6218 (N_6218,N_6145,N_6082);
or U6219 (N_6219,N_6060,N_6031);
nor U6220 (N_6220,N_6083,N_6057);
nand U6221 (N_6221,N_6043,N_6038);
nor U6222 (N_6222,N_6112,N_6036);
nor U6223 (N_6223,N_6042,N_6002);
and U6224 (N_6224,N_6129,N_6148);
xor U6225 (N_6225,N_6069,N_6102);
nor U6226 (N_6226,N_6104,N_6039);
nand U6227 (N_6227,N_6096,N_6076);
or U6228 (N_6228,N_6097,N_6018);
or U6229 (N_6229,N_6052,N_6146);
nor U6230 (N_6230,N_6036,N_6064);
nor U6231 (N_6231,N_6018,N_6062);
nand U6232 (N_6232,N_6106,N_6005);
xnor U6233 (N_6233,N_6140,N_6033);
or U6234 (N_6234,N_6134,N_6096);
nand U6235 (N_6235,N_6048,N_6047);
nand U6236 (N_6236,N_6012,N_6056);
nor U6237 (N_6237,N_6137,N_6062);
or U6238 (N_6238,N_6021,N_6091);
nor U6239 (N_6239,N_6008,N_6031);
nand U6240 (N_6240,N_6045,N_6149);
xnor U6241 (N_6241,N_6124,N_6058);
xnor U6242 (N_6242,N_6115,N_6111);
nand U6243 (N_6243,N_6029,N_6025);
nand U6244 (N_6244,N_6005,N_6038);
nor U6245 (N_6245,N_6092,N_6143);
nor U6246 (N_6246,N_6121,N_6110);
and U6247 (N_6247,N_6062,N_6119);
or U6248 (N_6248,N_6087,N_6074);
and U6249 (N_6249,N_6062,N_6029);
nand U6250 (N_6250,N_6006,N_6044);
xnor U6251 (N_6251,N_6013,N_6118);
nand U6252 (N_6252,N_6079,N_6038);
and U6253 (N_6253,N_6040,N_6105);
and U6254 (N_6254,N_6140,N_6087);
nand U6255 (N_6255,N_6005,N_6056);
nor U6256 (N_6256,N_6100,N_6081);
or U6257 (N_6257,N_6129,N_6077);
nand U6258 (N_6258,N_6007,N_6022);
nor U6259 (N_6259,N_6065,N_6098);
nor U6260 (N_6260,N_6019,N_6013);
nor U6261 (N_6261,N_6106,N_6067);
nand U6262 (N_6262,N_6019,N_6017);
xor U6263 (N_6263,N_6076,N_6124);
and U6264 (N_6264,N_6129,N_6113);
or U6265 (N_6265,N_6024,N_6069);
or U6266 (N_6266,N_6014,N_6072);
or U6267 (N_6267,N_6066,N_6147);
xor U6268 (N_6268,N_6075,N_6129);
nand U6269 (N_6269,N_6111,N_6051);
nand U6270 (N_6270,N_6067,N_6136);
and U6271 (N_6271,N_6079,N_6002);
and U6272 (N_6272,N_6055,N_6054);
or U6273 (N_6273,N_6071,N_6058);
nor U6274 (N_6274,N_6087,N_6042);
nor U6275 (N_6275,N_6144,N_6139);
and U6276 (N_6276,N_6111,N_6136);
or U6277 (N_6277,N_6132,N_6059);
nand U6278 (N_6278,N_6120,N_6138);
and U6279 (N_6279,N_6127,N_6053);
or U6280 (N_6280,N_6092,N_6061);
nor U6281 (N_6281,N_6020,N_6104);
nand U6282 (N_6282,N_6144,N_6008);
nor U6283 (N_6283,N_6112,N_6009);
nor U6284 (N_6284,N_6143,N_6030);
nor U6285 (N_6285,N_6014,N_6137);
nand U6286 (N_6286,N_6101,N_6143);
and U6287 (N_6287,N_6128,N_6011);
xnor U6288 (N_6288,N_6146,N_6035);
and U6289 (N_6289,N_6026,N_6068);
or U6290 (N_6290,N_6083,N_6011);
nand U6291 (N_6291,N_6105,N_6052);
nand U6292 (N_6292,N_6022,N_6016);
nor U6293 (N_6293,N_6105,N_6034);
nand U6294 (N_6294,N_6067,N_6066);
nand U6295 (N_6295,N_6032,N_6009);
nor U6296 (N_6296,N_6138,N_6088);
or U6297 (N_6297,N_6031,N_6022);
nand U6298 (N_6298,N_6127,N_6003);
and U6299 (N_6299,N_6044,N_6104);
nand U6300 (N_6300,N_6211,N_6282);
nor U6301 (N_6301,N_6188,N_6232);
xor U6302 (N_6302,N_6244,N_6227);
xor U6303 (N_6303,N_6284,N_6201);
xor U6304 (N_6304,N_6174,N_6208);
nor U6305 (N_6305,N_6265,N_6212);
or U6306 (N_6306,N_6299,N_6296);
nand U6307 (N_6307,N_6195,N_6269);
nor U6308 (N_6308,N_6150,N_6190);
and U6309 (N_6309,N_6159,N_6266);
nand U6310 (N_6310,N_6181,N_6209);
nand U6311 (N_6311,N_6247,N_6226);
nand U6312 (N_6312,N_6224,N_6241);
nor U6313 (N_6313,N_6240,N_6267);
and U6314 (N_6314,N_6249,N_6218);
and U6315 (N_6315,N_6228,N_6191);
and U6316 (N_6316,N_6237,N_6170);
nor U6317 (N_6317,N_6245,N_6225);
nor U6318 (N_6318,N_6271,N_6261);
xor U6319 (N_6319,N_6289,N_6205);
and U6320 (N_6320,N_6210,N_6217);
and U6321 (N_6321,N_6256,N_6287);
xor U6322 (N_6322,N_6162,N_6221);
and U6323 (N_6323,N_6176,N_6273);
and U6324 (N_6324,N_6281,N_6157);
or U6325 (N_6325,N_6242,N_6297);
nand U6326 (N_6326,N_6153,N_6246);
or U6327 (N_6327,N_6268,N_6192);
xor U6328 (N_6328,N_6197,N_6152);
nand U6329 (N_6329,N_6216,N_6235);
nand U6330 (N_6330,N_6275,N_6290);
nand U6331 (N_6331,N_6236,N_6272);
nand U6332 (N_6332,N_6182,N_6166);
nand U6333 (N_6333,N_6215,N_6257);
or U6334 (N_6334,N_6204,N_6206);
and U6335 (N_6335,N_6203,N_6194);
nand U6336 (N_6336,N_6183,N_6156);
nor U6337 (N_6337,N_6283,N_6186);
or U6338 (N_6338,N_6270,N_6274);
or U6339 (N_6339,N_6151,N_6178);
or U6340 (N_6340,N_6260,N_6280);
xnor U6341 (N_6341,N_6158,N_6243);
nand U6342 (N_6342,N_6171,N_6251);
and U6343 (N_6343,N_6259,N_6179);
or U6344 (N_6344,N_6231,N_6161);
and U6345 (N_6345,N_6169,N_6165);
nand U6346 (N_6346,N_6276,N_6154);
nor U6347 (N_6347,N_6295,N_6175);
and U6348 (N_6348,N_6293,N_6248);
nor U6349 (N_6349,N_6279,N_6298);
and U6350 (N_6350,N_6263,N_6163);
or U6351 (N_6351,N_6254,N_6294);
nor U6352 (N_6352,N_6198,N_6250);
nor U6353 (N_6353,N_6189,N_6223);
and U6354 (N_6354,N_6264,N_6214);
nor U6355 (N_6355,N_6258,N_6173);
nor U6356 (N_6356,N_6213,N_6291);
nand U6357 (N_6357,N_6222,N_6239);
xnor U6358 (N_6358,N_6262,N_6207);
nor U6359 (N_6359,N_6200,N_6233);
xor U6360 (N_6360,N_6180,N_6196);
nand U6361 (N_6361,N_6187,N_6277);
nor U6362 (N_6362,N_6177,N_6238);
or U6363 (N_6363,N_6288,N_6286);
nand U6364 (N_6364,N_6255,N_6219);
and U6365 (N_6365,N_6285,N_6185);
or U6366 (N_6366,N_6193,N_6167);
or U6367 (N_6367,N_6234,N_6252);
xnor U6368 (N_6368,N_6184,N_6292);
nor U6369 (N_6369,N_6230,N_6253);
and U6370 (N_6370,N_6172,N_6278);
and U6371 (N_6371,N_6160,N_6199);
nand U6372 (N_6372,N_6202,N_6229);
or U6373 (N_6373,N_6164,N_6220);
or U6374 (N_6374,N_6168,N_6155);
nand U6375 (N_6375,N_6172,N_6258);
or U6376 (N_6376,N_6264,N_6197);
or U6377 (N_6377,N_6240,N_6211);
or U6378 (N_6378,N_6256,N_6203);
nand U6379 (N_6379,N_6275,N_6286);
or U6380 (N_6380,N_6278,N_6232);
nor U6381 (N_6381,N_6293,N_6272);
and U6382 (N_6382,N_6293,N_6253);
nand U6383 (N_6383,N_6233,N_6203);
nand U6384 (N_6384,N_6262,N_6252);
or U6385 (N_6385,N_6181,N_6196);
nand U6386 (N_6386,N_6152,N_6236);
xor U6387 (N_6387,N_6261,N_6228);
nor U6388 (N_6388,N_6198,N_6264);
or U6389 (N_6389,N_6224,N_6237);
and U6390 (N_6390,N_6249,N_6169);
and U6391 (N_6391,N_6167,N_6277);
nor U6392 (N_6392,N_6234,N_6281);
and U6393 (N_6393,N_6173,N_6154);
and U6394 (N_6394,N_6200,N_6162);
and U6395 (N_6395,N_6233,N_6268);
and U6396 (N_6396,N_6226,N_6221);
nand U6397 (N_6397,N_6176,N_6205);
or U6398 (N_6398,N_6267,N_6210);
nor U6399 (N_6399,N_6226,N_6263);
nor U6400 (N_6400,N_6195,N_6294);
nand U6401 (N_6401,N_6258,N_6155);
nand U6402 (N_6402,N_6186,N_6281);
nor U6403 (N_6403,N_6173,N_6227);
or U6404 (N_6404,N_6194,N_6167);
and U6405 (N_6405,N_6256,N_6189);
or U6406 (N_6406,N_6263,N_6297);
and U6407 (N_6407,N_6252,N_6177);
and U6408 (N_6408,N_6176,N_6295);
xor U6409 (N_6409,N_6258,N_6232);
xor U6410 (N_6410,N_6162,N_6192);
nand U6411 (N_6411,N_6196,N_6199);
and U6412 (N_6412,N_6271,N_6296);
or U6413 (N_6413,N_6172,N_6218);
nand U6414 (N_6414,N_6266,N_6269);
xnor U6415 (N_6415,N_6189,N_6247);
and U6416 (N_6416,N_6175,N_6150);
nor U6417 (N_6417,N_6181,N_6167);
and U6418 (N_6418,N_6276,N_6226);
nand U6419 (N_6419,N_6177,N_6170);
nand U6420 (N_6420,N_6252,N_6266);
xor U6421 (N_6421,N_6193,N_6180);
nand U6422 (N_6422,N_6192,N_6231);
and U6423 (N_6423,N_6166,N_6297);
nor U6424 (N_6424,N_6297,N_6170);
or U6425 (N_6425,N_6260,N_6226);
or U6426 (N_6426,N_6196,N_6233);
and U6427 (N_6427,N_6285,N_6157);
nand U6428 (N_6428,N_6184,N_6201);
and U6429 (N_6429,N_6296,N_6166);
or U6430 (N_6430,N_6168,N_6268);
and U6431 (N_6431,N_6175,N_6155);
xnor U6432 (N_6432,N_6238,N_6280);
or U6433 (N_6433,N_6266,N_6162);
or U6434 (N_6434,N_6251,N_6282);
nand U6435 (N_6435,N_6177,N_6183);
or U6436 (N_6436,N_6224,N_6280);
or U6437 (N_6437,N_6179,N_6286);
xnor U6438 (N_6438,N_6174,N_6168);
nand U6439 (N_6439,N_6242,N_6279);
or U6440 (N_6440,N_6171,N_6277);
nor U6441 (N_6441,N_6201,N_6167);
and U6442 (N_6442,N_6231,N_6181);
nor U6443 (N_6443,N_6250,N_6225);
nor U6444 (N_6444,N_6205,N_6288);
and U6445 (N_6445,N_6190,N_6276);
and U6446 (N_6446,N_6188,N_6221);
or U6447 (N_6447,N_6297,N_6249);
nor U6448 (N_6448,N_6188,N_6240);
nand U6449 (N_6449,N_6187,N_6184);
or U6450 (N_6450,N_6433,N_6392);
or U6451 (N_6451,N_6447,N_6401);
and U6452 (N_6452,N_6366,N_6420);
nor U6453 (N_6453,N_6425,N_6308);
or U6454 (N_6454,N_6375,N_6386);
or U6455 (N_6455,N_6443,N_6387);
nand U6456 (N_6456,N_6376,N_6396);
nand U6457 (N_6457,N_6402,N_6432);
nand U6458 (N_6458,N_6324,N_6332);
nand U6459 (N_6459,N_6361,N_6384);
and U6460 (N_6460,N_6318,N_6393);
and U6461 (N_6461,N_6403,N_6359);
and U6462 (N_6462,N_6441,N_6369);
nand U6463 (N_6463,N_6302,N_6426);
nand U6464 (N_6464,N_6325,N_6427);
or U6465 (N_6465,N_6343,N_6333);
or U6466 (N_6466,N_6335,N_6444);
nor U6467 (N_6467,N_6352,N_6394);
or U6468 (N_6468,N_6445,N_6310);
and U6469 (N_6469,N_6382,N_6309);
or U6470 (N_6470,N_6411,N_6312);
and U6471 (N_6471,N_6337,N_6364);
or U6472 (N_6472,N_6344,N_6347);
nand U6473 (N_6473,N_6349,N_6398);
nand U6474 (N_6474,N_6418,N_6415);
xor U6475 (N_6475,N_6301,N_6435);
or U6476 (N_6476,N_6336,N_6395);
and U6477 (N_6477,N_6306,N_6338);
or U6478 (N_6478,N_6400,N_6363);
and U6479 (N_6479,N_6404,N_6390);
nor U6480 (N_6480,N_6350,N_6331);
nand U6481 (N_6481,N_6323,N_6304);
nand U6482 (N_6482,N_6348,N_6383);
nand U6483 (N_6483,N_6367,N_6421);
nor U6484 (N_6484,N_6320,N_6365);
and U6485 (N_6485,N_6438,N_6431);
and U6486 (N_6486,N_6440,N_6407);
nand U6487 (N_6487,N_6428,N_6345);
nand U6488 (N_6488,N_6379,N_6409);
or U6489 (N_6489,N_6341,N_6340);
nand U6490 (N_6490,N_6448,N_6449);
and U6491 (N_6491,N_6354,N_6351);
and U6492 (N_6492,N_6436,N_6430);
and U6493 (N_6493,N_6300,N_6319);
and U6494 (N_6494,N_6374,N_6355);
and U6495 (N_6495,N_6327,N_6357);
or U6496 (N_6496,N_6362,N_6321);
or U6497 (N_6497,N_6405,N_6322);
xor U6498 (N_6498,N_6339,N_6391);
and U6499 (N_6499,N_6414,N_6388);
nor U6500 (N_6500,N_6358,N_6330);
or U6501 (N_6501,N_6397,N_6368);
xor U6502 (N_6502,N_6315,N_6303);
xnor U6503 (N_6503,N_6423,N_6371);
or U6504 (N_6504,N_6389,N_6378);
nor U6505 (N_6505,N_6417,N_6439);
nor U6506 (N_6506,N_6353,N_6437);
xor U6507 (N_6507,N_6377,N_6442);
nor U6508 (N_6508,N_6399,N_6381);
nand U6509 (N_6509,N_6316,N_6416);
or U6510 (N_6510,N_6360,N_6385);
nand U6511 (N_6511,N_6311,N_6356);
nor U6512 (N_6512,N_6408,N_6314);
nand U6513 (N_6513,N_6328,N_6424);
or U6514 (N_6514,N_6372,N_6346);
or U6515 (N_6515,N_6326,N_6406);
or U6516 (N_6516,N_6422,N_6434);
xnor U6517 (N_6517,N_6370,N_6413);
or U6518 (N_6518,N_6446,N_6334);
and U6519 (N_6519,N_6329,N_6313);
and U6520 (N_6520,N_6342,N_6305);
or U6521 (N_6521,N_6380,N_6419);
nor U6522 (N_6522,N_6410,N_6307);
nand U6523 (N_6523,N_6429,N_6373);
and U6524 (N_6524,N_6412,N_6317);
or U6525 (N_6525,N_6301,N_6380);
and U6526 (N_6526,N_6406,N_6325);
xor U6527 (N_6527,N_6315,N_6329);
or U6528 (N_6528,N_6435,N_6311);
nor U6529 (N_6529,N_6426,N_6412);
nor U6530 (N_6530,N_6301,N_6344);
nand U6531 (N_6531,N_6426,N_6344);
and U6532 (N_6532,N_6374,N_6402);
nor U6533 (N_6533,N_6355,N_6326);
or U6534 (N_6534,N_6403,N_6352);
and U6535 (N_6535,N_6423,N_6410);
or U6536 (N_6536,N_6327,N_6369);
xnor U6537 (N_6537,N_6366,N_6308);
and U6538 (N_6538,N_6396,N_6406);
xnor U6539 (N_6539,N_6423,N_6408);
nor U6540 (N_6540,N_6353,N_6407);
or U6541 (N_6541,N_6346,N_6327);
xnor U6542 (N_6542,N_6417,N_6369);
nand U6543 (N_6543,N_6408,N_6383);
or U6544 (N_6544,N_6422,N_6389);
nor U6545 (N_6545,N_6304,N_6379);
xnor U6546 (N_6546,N_6325,N_6309);
and U6547 (N_6547,N_6415,N_6304);
nand U6548 (N_6548,N_6330,N_6425);
nor U6549 (N_6549,N_6396,N_6311);
nand U6550 (N_6550,N_6349,N_6390);
and U6551 (N_6551,N_6369,N_6426);
or U6552 (N_6552,N_6326,N_6422);
nand U6553 (N_6553,N_6426,N_6416);
nor U6554 (N_6554,N_6328,N_6358);
and U6555 (N_6555,N_6303,N_6334);
nand U6556 (N_6556,N_6417,N_6364);
nor U6557 (N_6557,N_6326,N_6385);
xor U6558 (N_6558,N_6430,N_6415);
or U6559 (N_6559,N_6431,N_6430);
or U6560 (N_6560,N_6385,N_6333);
nor U6561 (N_6561,N_6398,N_6435);
or U6562 (N_6562,N_6420,N_6319);
or U6563 (N_6563,N_6365,N_6338);
nor U6564 (N_6564,N_6351,N_6385);
nor U6565 (N_6565,N_6330,N_6416);
or U6566 (N_6566,N_6411,N_6376);
nand U6567 (N_6567,N_6337,N_6349);
nand U6568 (N_6568,N_6324,N_6354);
or U6569 (N_6569,N_6379,N_6325);
xnor U6570 (N_6570,N_6378,N_6364);
nor U6571 (N_6571,N_6394,N_6330);
xnor U6572 (N_6572,N_6325,N_6307);
and U6573 (N_6573,N_6376,N_6324);
nand U6574 (N_6574,N_6424,N_6307);
xnor U6575 (N_6575,N_6363,N_6444);
or U6576 (N_6576,N_6306,N_6407);
or U6577 (N_6577,N_6312,N_6421);
nor U6578 (N_6578,N_6435,N_6416);
or U6579 (N_6579,N_6313,N_6354);
or U6580 (N_6580,N_6354,N_6339);
nor U6581 (N_6581,N_6444,N_6413);
and U6582 (N_6582,N_6434,N_6416);
nor U6583 (N_6583,N_6443,N_6350);
and U6584 (N_6584,N_6376,N_6418);
and U6585 (N_6585,N_6365,N_6307);
and U6586 (N_6586,N_6322,N_6385);
and U6587 (N_6587,N_6329,N_6405);
and U6588 (N_6588,N_6353,N_6375);
nand U6589 (N_6589,N_6379,N_6382);
and U6590 (N_6590,N_6374,N_6403);
and U6591 (N_6591,N_6398,N_6300);
and U6592 (N_6592,N_6398,N_6388);
or U6593 (N_6593,N_6355,N_6411);
or U6594 (N_6594,N_6386,N_6310);
nor U6595 (N_6595,N_6372,N_6384);
xor U6596 (N_6596,N_6309,N_6347);
nand U6597 (N_6597,N_6344,N_6328);
or U6598 (N_6598,N_6326,N_6374);
and U6599 (N_6599,N_6437,N_6444);
xor U6600 (N_6600,N_6464,N_6592);
xnor U6601 (N_6601,N_6453,N_6529);
nor U6602 (N_6602,N_6490,N_6575);
and U6603 (N_6603,N_6478,N_6546);
or U6604 (N_6604,N_6457,N_6485);
and U6605 (N_6605,N_6554,N_6562);
xor U6606 (N_6606,N_6527,N_6566);
and U6607 (N_6607,N_6551,N_6555);
nor U6608 (N_6608,N_6491,N_6567);
xnor U6609 (N_6609,N_6511,N_6458);
or U6610 (N_6610,N_6573,N_6514);
or U6611 (N_6611,N_6450,N_6472);
nand U6612 (N_6612,N_6599,N_6531);
nor U6613 (N_6613,N_6483,N_6545);
and U6614 (N_6614,N_6513,N_6556);
or U6615 (N_6615,N_6506,N_6536);
xnor U6616 (N_6616,N_6535,N_6508);
and U6617 (N_6617,N_6582,N_6578);
and U6618 (N_6618,N_6591,N_6540);
and U6619 (N_6619,N_6470,N_6523);
and U6620 (N_6620,N_6522,N_6524);
nand U6621 (N_6621,N_6565,N_6469);
or U6622 (N_6622,N_6560,N_6482);
nand U6623 (N_6623,N_6475,N_6509);
nand U6624 (N_6624,N_6494,N_6497);
xor U6625 (N_6625,N_6486,N_6585);
or U6626 (N_6626,N_6541,N_6595);
nand U6627 (N_6627,N_6452,N_6550);
and U6628 (N_6628,N_6539,N_6564);
or U6629 (N_6629,N_6476,N_6587);
xor U6630 (N_6630,N_6547,N_6576);
xor U6631 (N_6631,N_6520,N_6503);
nor U6632 (N_6632,N_6577,N_6574);
and U6633 (N_6633,N_6586,N_6559);
and U6634 (N_6634,N_6590,N_6583);
nor U6635 (N_6635,N_6563,N_6533);
nand U6636 (N_6636,N_6552,N_6537);
nand U6637 (N_6637,N_6543,N_6542);
nand U6638 (N_6638,N_6517,N_6515);
nor U6639 (N_6639,N_6549,N_6571);
xnor U6640 (N_6640,N_6459,N_6507);
xnor U6641 (N_6641,N_6568,N_6593);
or U6642 (N_6642,N_6468,N_6473);
and U6643 (N_6643,N_6488,N_6467);
xor U6644 (N_6644,N_6548,N_6597);
xnor U6645 (N_6645,N_6525,N_6489);
and U6646 (N_6646,N_6460,N_6579);
nand U6647 (N_6647,N_6484,N_6456);
nand U6648 (N_6648,N_6584,N_6501);
nand U6649 (N_6649,N_6500,N_6505);
nand U6650 (N_6650,N_6526,N_6471);
nand U6651 (N_6651,N_6461,N_6477);
and U6652 (N_6652,N_6479,N_6492);
nand U6653 (N_6653,N_6519,N_6496);
or U6654 (N_6654,N_6544,N_6454);
xnor U6655 (N_6655,N_6572,N_6495);
nor U6656 (N_6656,N_6451,N_6530);
or U6657 (N_6657,N_6588,N_6487);
nor U6658 (N_6658,N_6558,N_6518);
nor U6659 (N_6659,N_6480,N_6596);
nor U6660 (N_6660,N_6532,N_6557);
nor U6661 (N_6661,N_6516,N_6455);
or U6662 (N_6662,N_6553,N_6512);
and U6663 (N_6663,N_6493,N_6561);
nor U6664 (N_6664,N_6598,N_6581);
xnor U6665 (N_6665,N_6463,N_6462);
and U6666 (N_6666,N_6465,N_6504);
nor U6667 (N_6667,N_6570,N_6466);
or U6668 (N_6668,N_6589,N_6499);
or U6669 (N_6669,N_6498,N_6510);
nand U6670 (N_6670,N_6502,N_6528);
and U6671 (N_6671,N_6580,N_6474);
and U6672 (N_6672,N_6481,N_6569);
nand U6673 (N_6673,N_6594,N_6534);
and U6674 (N_6674,N_6521,N_6538);
or U6675 (N_6675,N_6455,N_6494);
or U6676 (N_6676,N_6458,N_6506);
or U6677 (N_6677,N_6530,N_6553);
or U6678 (N_6678,N_6453,N_6510);
and U6679 (N_6679,N_6487,N_6475);
nand U6680 (N_6680,N_6546,N_6498);
nor U6681 (N_6681,N_6491,N_6563);
and U6682 (N_6682,N_6563,N_6504);
nor U6683 (N_6683,N_6575,N_6530);
nor U6684 (N_6684,N_6502,N_6539);
xor U6685 (N_6685,N_6561,N_6576);
nor U6686 (N_6686,N_6524,N_6593);
or U6687 (N_6687,N_6593,N_6529);
and U6688 (N_6688,N_6502,N_6522);
nand U6689 (N_6689,N_6497,N_6524);
or U6690 (N_6690,N_6504,N_6487);
xor U6691 (N_6691,N_6529,N_6516);
or U6692 (N_6692,N_6548,N_6549);
or U6693 (N_6693,N_6508,N_6483);
nand U6694 (N_6694,N_6477,N_6493);
and U6695 (N_6695,N_6504,N_6598);
or U6696 (N_6696,N_6558,N_6463);
or U6697 (N_6697,N_6473,N_6499);
nand U6698 (N_6698,N_6557,N_6561);
nand U6699 (N_6699,N_6539,N_6463);
nor U6700 (N_6700,N_6548,N_6562);
nand U6701 (N_6701,N_6560,N_6474);
or U6702 (N_6702,N_6597,N_6450);
nor U6703 (N_6703,N_6471,N_6550);
or U6704 (N_6704,N_6508,N_6452);
or U6705 (N_6705,N_6480,N_6515);
nor U6706 (N_6706,N_6546,N_6545);
and U6707 (N_6707,N_6536,N_6563);
nor U6708 (N_6708,N_6567,N_6541);
or U6709 (N_6709,N_6509,N_6567);
xnor U6710 (N_6710,N_6584,N_6597);
nor U6711 (N_6711,N_6517,N_6587);
and U6712 (N_6712,N_6597,N_6555);
or U6713 (N_6713,N_6533,N_6459);
or U6714 (N_6714,N_6557,N_6555);
or U6715 (N_6715,N_6454,N_6497);
nor U6716 (N_6716,N_6525,N_6497);
nand U6717 (N_6717,N_6546,N_6457);
nand U6718 (N_6718,N_6552,N_6566);
or U6719 (N_6719,N_6540,N_6468);
nor U6720 (N_6720,N_6547,N_6584);
nor U6721 (N_6721,N_6471,N_6500);
and U6722 (N_6722,N_6508,N_6528);
or U6723 (N_6723,N_6473,N_6488);
and U6724 (N_6724,N_6480,N_6547);
nand U6725 (N_6725,N_6528,N_6583);
nand U6726 (N_6726,N_6553,N_6466);
or U6727 (N_6727,N_6527,N_6484);
or U6728 (N_6728,N_6598,N_6584);
nand U6729 (N_6729,N_6460,N_6550);
and U6730 (N_6730,N_6515,N_6589);
or U6731 (N_6731,N_6470,N_6478);
or U6732 (N_6732,N_6557,N_6593);
nand U6733 (N_6733,N_6513,N_6551);
and U6734 (N_6734,N_6463,N_6479);
and U6735 (N_6735,N_6493,N_6542);
or U6736 (N_6736,N_6559,N_6481);
and U6737 (N_6737,N_6509,N_6533);
nor U6738 (N_6738,N_6589,N_6580);
or U6739 (N_6739,N_6483,N_6590);
or U6740 (N_6740,N_6505,N_6548);
or U6741 (N_6741,N_6470,N_6491);
nand U6742 (N_6742,N_6498,N_6556);
or U6743 (N_6743,N_6534,N_6508);
nor U6744 (N_6744,N_6474,N_6594);
and U6745 (N_6745,N_6452,N_6460);
nand U6746 (N_6746,N_6502,N_6533);
nor U6747 (N_6747,N_6459,N_6598);
or U6748 (N_6748,N_6483,N_6596);
or U6749 (N_6749,N_6543,N_6495);
or U6750 (N_6750,N_6698,N_6608);
nor U6751 (N_6751,N_6748,N_6733);
nor U6752 (N_6752,N_6647,N_6614);
xor U6753 (N_6753,N_6669,N_6728);
nor U6754 (N_6754,N_6712,N_6702);
nor U6755 (N_6755,N_6622,N_6644);
and U6756 (N_6756,N_6711,N_6726);
or U6757 (N_6757,N_6679,N_6690);
nor U6758 (N_6758,N_6625,N_6600);
nand U6759 (N_6759,N_6727,N_6717);
and U6760 (N_6760,N_6675,N_6646);
nand U6761 (N_6761,N_6655,N_6616);
nor U6762 (N_6762,N_6657,N_6664);
nor U6763 (N_6763,N_6641,N_6709);
and U6764 (N_6764,N_6618,N_6610);
or U6765 (N_6765,N_6701,N_6639);
xor U6766 (N_6766,N_6694,N_6637);
nor U6767 (N_6767,N_6668,N_6674);
nor U6768 (N_6768,N_6615,N_6693);
or U6769 (N_6769,N_6627,N_6621);
and U6770 (N_6770,N_6628,N_6658);
and U6771 (N_6771,N_6603,N_6652);
nor U6772 (N_6772,N_6672,N_6602);
nand U6773 (N_6773,N_6700,N_6683);
nor U6774 (N_6774,N_6697,N_6643);
xor U6775 (N_6775,N_6740,N_6730);
or U6776 (N_6776,N_6629,N_6651);
and U6777 (N_6777,N_6634,N_6649);
xnor U6778 (N_6778,N_6689,N_6623);
nor U6779 (N_6779,N_6612,N_6656);
nor U6780 (N_6780,N_6636,N_6722);
or U6781 (N_6781,N_6613,N_6619);
nand U6782 (N_6782,N_6617,N_6737);
nor U6783 (N_6783,N_6666,N_6747);
and U6784 (N_6784,N_6638,N_6606);
xor U6785 (N_6785,N_6734,N_6654);
nor U6786 (N_6786,N_6601,N_6620);
xor U6787 (N_6787,N_6632,N_6681);
and U6788 (N_6788,N_6670,N_6745);
nand U6789 (N_6789,N_6631,N_6677);
nand U6790 (N_6790,N_6604,N_6626);
nand U6791 (N_6791,N_6715,N_6710);
nor U6792 (N_6792,N_6736,N_6741);
and U6793 (N_6793,N_6725,N_6744);
nor U6794 (N_6794,N_6721,N_6605);
and U6795 (N_6795,N_6706,N_6723);
or U6796 (N_6796,N_6718,N_6714);
or U6797 (N_6797,N_6716,N_6731);
or U6798 (N_6798,N_6673,N_6708);
nand U6799 (N_6799,N_6692,N_6633);
nand U6800 (N_6800,N_6635,N_6695);
xor U6801 (N_6801,N_6648,N_6720);
xnor U6802 (N_6802,N_6611,N_6703);
nor U6803 (N_6803,N_6665,N_6713);
nor U6804 (N_6804,N_6630,N_6724);
nor U6805 (N_6805,N_6686,N_6749);
or U6806 (N_6806,N_6688,N_6705);
or U6807 (N_6807,N_6660,N_6645);
or U6808 (N_6808,N_6739,N_6696);
nand U6809 (N_6809,N_6678,N_6653);
and U6810 (N_6810,N_6742,N_6704);
nor U6811 (N_6811,N_6661,N_6746);
or U6812 (N_6812,N_6691,N_6684);
or U6813 (N_6813,N_6687,N_6676);
and U6814 (N_6814,N_6659,N_6738);
nand U6815 (N_6815,N_6682,N_6667);
and U6816 (N_6816,N_6663,N_6743);
nand U6817 (N_6817,N_6685,N_6707);
nor U6818 (N_6818,N_6609,N_6650);
or U6819 (N_6819,N_6719,N_6662);
nand U6820 (N_6820,N_6699,N_6642);
and U6821 (N_6821,N_6624,N_6680);
nand U6822 (N_6822,N_6607,N_6732);
nand U6823 (N_6823,N_6671,N_6735);
and U6824 (N_6824,N_6640,N_6729);
or U6825 (N_6825,N_6727,N_6604);
and U6826 (N_6826,N_6701,N_6635);
or U6827 (N_6827,N_6672,N_6643);
nand U6828 (N_6828,N_6629,N_6690);
and U6829 (N_6829,N_6623,N_6705);
nand U6830 (N_6830,N_6689,N_6685);
and U6831 (N_6831,N_6705,N_6696);
nor U6832 (N_6832,N_6657,N_6644);
xnor U6833 (N_6833,N_6718,N_6635);
or U6834 (N_6834,N_6651,N_6648);
nand U6835 (N_6835,N_6663,N_6614);
or U6836 (N_6836,N_6628,N_6701);
and U6837 (N_6837,N_6641,N_6692);
nand U6838 (N_6838,N_6628,N_6632);
or U6839 (N_6839,N_6613,N_6728);
nor U6840 (N_6840,N_6601,N_6681);
nor U6841 (N_6841,N_6707,N_6684);
or U6842 (N_6842,N_6633,N_6668);
or U6843 (N_6843,N_6726,N_6721);
or U6844 (N_6844,N_6715,N_6730);
nor U6845 (N_6845,N_6636,N_6604);
or U6846 (N_6846,N_6600,N_6723);
nand U6847 (N_6847,N_6652,N_6671);
nor U6848 (N_6848,N_6616,N_6743);
nand U6849 (N_6849,N_6610,N_6600);
nand U6850 (N_6850,N_6674,N_6645);
nor U6851 (N_6851,N_6748,N_6724);
or U6852 (N_6852,N_6717,N_6631);
and U6853 (N_6853,N_6728,N_6693);
or U6854 (N_6854,N_6717,N_6744);
or U6855 (N_6855,N_6637,N_6622);
nor U6856 (N_6856,N_6717,N_6677);
or U6857 (N_6857,N_6732,N_6649);
nand U6858 (N_6858,N_6639,N_6610);
nor U6859 (N_6859,N_6730,N_6738);
nor U6860 (N_6860,N_6661,N_6640);
nor U6861 (N_6861,N_6658,N_6613);
nand U6862 (N_6862,N_6730,N_6660);
nand U6863 (N_6863,N_6682,N_6601);
nand U6864 (N_6864,N_6626,N_6685);
and U6865 (N_6865,N_6617,N_6632);
or U6866 (N_6866,N_6748,N_6610);
nor U6867 (N_6867,N_6715,N_6697);
nor U6868 (N_6868,N_6625,N_6658);
xor U6869 (N_6869,N_6607,N_6663);
nand U6870 (N_6870,N_6623,N_6633);
and U6871 (N_6871,N_6650,N_6645);
nor U6872 (N_6872,N_6666,N_6658);
nor U6873 (N_6873,N_6700,N_6746);
and U6874 (N_6874,N_6743,N_6747);
and U6875 (N_6875,N_6685,N_6632);
nand U6876 (N_6876,N_6633,N_6727);
nor U6877 (N_6877,N_6682,N_6744);
or U6878 (N_6878,N_6623,N_6620);
nand U6879 (N_6879,N_6668,N_6736);
nor U6880 (N_6880,N_6749,N_6625);
nor U6881 (N_6881,N_6600,N_6614);
nand U6882 (N_6882,N_6707,N_6725);
nand U6883 (N_6883,N_6680,N_6745);
or U6884 (N_6884,N_6720,N_6661);
or U6885 (N_6885,N_6663,N_6609);
and U6886 (N_6886,N_6719,N_6643);
xor U6887 (N_6887,N_6702,N_6678);
nand U6888 (N_6888,N_6679,N_6693);
nor U6889 (N_6889,N_6619,N_6685);
or U6890 (N_6890,N_6690,N_6606);
nor U6891 (N_6891,N_6682,N_6670);
nor U6892 (N_6892,N_6638,N_6653);
xnor U6893 (N_6893,N_6625,N_6660);
nor U6894 (N_6894,N_6641,N_6626);
and U6895 (N_6895,N_6606,N_6732);
nand U6896 (N_6896,N_6724,N_6703);
nor U6897 (N_6897,N_6646,N_6687);
nor U6898 (N_6898,N_6676,N_6724);
or U6899 (N_6899,N_6664,N_6667);
xnor U6900 (N_6900,N_6800,N_6772);
nand U6901 (N_6901,N_6805,N_6836);
nand U6902 (N_6902,N_6830,N_6886);
or U6903 (N_6903,N_6854,N_6813);
nor U6904 (N_6904,N_6823,N_6792);
xnor U6905 (N_6905,N_6751,N_6769);
nand U6906 (N_6906,N_6758,N_6812);
nand U6907 (N_6907,N_6819,N_6875);
and U6908 (N_6908,N_6787,N_6781);
nand U6909 (N_6909,N_6807,N_6871);
and U6910 (N_6910,N_6782,N_6859);
nand U6911 (N_6911,N_6778,N_6867);
nor U6912 (N_6912,N_6874,N_6788);
nor U6913 (N_6913,N_6882,N_6811);
and U6914 (N_6914,N_6761,N_6797);
or U6915 (N_6915,N_6780,N_6759);
or U6916 (N_6916,N_6771,N_6766);
and U6917 (N_6917,N_6833,N_6850);
nand U6918 (N_6918,N_6767,N_6808);
nor U6919 (N_6919,N_6831,N_6868);
or U6920 (N_6920,N_6869,N_6834);
xnor U6921 (N_6921,N_6757,N_6814);
nor U6922 (N_6922,N_6793,N_6750);
nand U6923 (N_6923,N_6784,N_6876);
nor U6924 (N_6924,N_6822,N_6764);
nor U6925 (N_6925,N_6885,N_6789);
nor U6926 (N_6926,N_6779,N_6775);
or U6927 (N_6927,N_6851,N_6818);
and U6928 (N_6928,N_6809,N_6873);
and U6929 (N_6929,N_6825,N_6796);
xor U6930 (N_6930,N_6752,N_6846);
nor U6931 (N_6931,N_6839,N_6877);
or U6932 (N_6932,N_6794,N_6849);
nor U6933 (N_6933,N_6858,N_6888);
or U6934 (N_6934,N_6754,N_6898);
nand U6935 (N_6935,N_6791,N_6817);
and U6936 (N_6936,N_6881,N_6860);
nand U6937 (N_6937,N_6899,N_6756);
and U6938 (N_6938,N_6861,N_6755);
and U6939 (N_6939,N_6820,N_6835);
nor U6940 (N_6940,N_6786,N_6847);
and U6941 (N_6941,N_6803,N_6856);
and U6942 (N_6942,N_6768,N_6765);
xnor U6943 (N_6943,N_6790,N_6845);
or U6944 (N_6944,N_6810,N_6855);
nor U6945 (N_6945,N_6897,N_6827);
nand U6946 (N_6946,N_6848,N_6777);
and U6947 (N_6947,N_6774,N_6798);
or U6948 (N_6948,N_6844,N_6872);
nand U6949 (N_6949,N_6773,N_6770);
and U6950 (N_6950,N_6870,N_6862);
nand U6951 (N_6951,N_6802,N_6890);
nor U6952 (N_6952,N_6864,N_6763);
nor U6953 (N_6953,N_6852,N_6795);
and U6954 (N_6954,N_6837,N_6896);
and U6955 (N_6955,N_6843,N_6762);
nand U6956 (N_6956,N_6884,N_6753);
or U6957 (N_6957,N_6783,N_6801);
and U6958 (N_6958,N_6829,N_6857);
nor U6959 (N_6959,N_6841,N_6895);
xnor U6960 (N_6960,N_6806,N_6826);
xnor U6961 (N_6961,N_6832,N_6799);
or U6962 (N_6962,N_6883,N_6866);
or U6963 (N_6963,N_6840,N_6894);
or U6964 (N_6964,N_6824,N_6815);
nor U6965 (N_6965,N_6887,N_6760);
nand U6966 (N_6966,N_6880,N_6892);
or U6967 (N_6967,N_6785,N_6879);
or U6968 (N_6968,N_6853,N_6893);
or U6969 (N_6969,N_6776,N_6838);
xor U6970 (N_6970,N_6816,N_6828);
xnor U6971 (N_6971,N_6821,N_6878);
or U6972 (N_6972,N_6804,N_6863);
nand U6973 (N_6973,N_6865,N_6842);
nor U6974 (N_6974,N_6889,N_6891);
and U6975 (N_6975,N_6856,N_6790);
xor U6976 (N_6976,N_6890,N_6898);
nor U6977 (N_6977,N_6798,N_6866);
and U6978 (N_6978,N_6752,N_6879);
nor U6979 (N_6979,N_6859,N_6848);
nor U6980 (N_6980,N_6887,N_6751);
nand U6981 (N_6981,N_6867,N_6765);
xnor U6982 (N_6982,N_6768,N_6870);
and U6983 (N_6983,N_6869,N_6831);
nand U6984 (N_6984,N_6850,N_6776);
and U6985 (N_6985,N_6828,N_6756);
nand U6986 (N_6986,N_6782,N_6886);
and U6987 (N_6987,N_6899,N_6896);
xnor U6988 (N_6988,N_6826,N_6779);
xor U6989 (N_6989,N_6867,N_6806);
nand U6990 (N_6990,N_6797,N_6795);
and U6991 (N_6991,N_6764,N_6867);
and U6992 (N_6992,N_6848,N_6802);
or U6993 (N_6993,N_6852,N_6817);
nor U6994 (N_6994,N_6855,N_6777);
xnor U6995 (N_6995,N_6858,N_6823);
nand U6996 (N_6996,N_6871,N_6768);
xnor U6997 (N_6997,N_6803,N_6771);
nand U6998 (N_6998,N_6764,N_6842);
nor U6999 (N_6999,N_6860,N_6830);
nor U7000 (N_7000,N_6791,N_6768);
nand U7001 (N_7001,N_6782,N_6800);
or U7002 (N_7002,N_6885,N_6836);
and U7003 (N_7003,N_6776,N_6899);
or U7004 (N_7004,N_6864,N_6808);
nor U7005 (N_7005,N_6831,N_6850);
and U7006 (N_7006,N_6771,N_6850);
nand U7007 (N_7007,N_6809,N_6885);
nor U7008 (N_7008,N_6890,N_6855);
nor U7009 (N_7009,N_6860,N_6868);
or U7010 (N_7010,N_6790,N_6781);
and U7011 (N_7011,N_6757,N_6889);
or U7012 (N_7012,N_6846,N_6859);
xnor U7013 (N_7013,N_6787,N_6798);
nor U7014 (N_7014,N_6855,N_6802);
and U7015 (N_7015,N_6847,N_6873);
and U7016 (N_7016,N_6866,N_6854);
and U7017 (N_7017,N_6889,N_6876);
xnor U7018 (N_7018,N_6877,N_6785);
nand U7019 (N_7019,N_6788,N_6803);
nor U7020 (N_7020,N_6888,N_6860);
nor U7021 (N_7021,N_6863,N_6801);
and U7022 (N_7022,N_6800,N_6864);
or U7023 (N_7023,N_6811,N_6763);
or U7024 (N_7024,N_6861,N_6882);
or U7025 (N_7025,N_6844,N_6791);
nand U7026 (N_7026,N_6804,N_6883);
xor U7027 (N_7027,N_6870,N_6802);
nor U7028 (N_7028,N_6884,N_6898);
and U7029 (N_7029,N_6758,N_6860);
and U7030 (N_7030,N_6820,N_6765);
or U7031 (N_7031,N_6897,N_6793);
xor U7032 (N_7032,N_6826,N_6805);
nor U7033 (N_7033,N_6898,N_6879);
or U7034 (N_7034,N_6872,N_6798);
and U7035 (N_7035,N_6757,N_6797);
nand U7036 (N_7036,N_6825,N_6821);
or U7037 (N_7037,N_6866,N_6806);
and U7038 (N_7038,N_6844,N_6893);
or U7039 (N_7039,N_6870,N_6899);
or U7040 (N_7040,N_6870,N_6769);
nor U7041 (N_7041,N_6838,N_6811);
xnor U7042 (N_7042,N_6843,N_6876);
nor U7043 (N_7043,N_6816,N_6757);
and U7044 (N_7044,N_6779,N_6791);
or U7045 (N_7045,N_6899,N_6857);
nor U7046 (N_7046,N_6797,N_6774);
and U7047 (N_7047,N_6823,N_6798);
nand U7048 (N_7048,N_6785,N_6795);
xor U7049 (N_7049,N_6787,N_6755);
and U7050 (N_7050,N_7001,N_7033);
nand U7051 (N_7051,N_6977,N_7000);
and U7052 (N_7052,N_6968,N_6934);
or U7053 (N_7053,N_6996,N_6950);
or U7054 (N_7054,N_6910,N_7012);
and U7055 (N_7055,N_6944,N_6901);
nand U7056 (N_7056,N_7035,N_6915);
and U7057 (N_7057,N_6923,N_6908);
xor U7058 (N_7058,N_7036,N_7037);
or U7059 (N_7059,N_7004,N_6964);
nand U7060 (N_7060,N_6993,N_6928);
and U7061 (N_7061,N_7046,N_6945);
and U7062 (N_7062,N_6920,N_7030);
nand U7063 (N_7063,N_6932,N_6998);
nor U7064 (N_7064,N_6965,N_7040);
nor U7065 (N_7065,N_6989,N_6984);
nand U7066 (N_7066,N_6999,N_6905);
or U7067 (N_7067,N_6921,N_6949);
nand U7068 (N_7068,N_7003,N_6995);
nand U7069 (N_7069,N_6971,N_7017);
or U7070 (N_7070,N_6969,N_6987);
or U7071 (N_7071,N_7042,N_6979);
nand U7072 (N_7072,N_6927,N_6967);
nor U7073 (N_7073,N_6904,N_7009);
or U7074 (N_7074,N_6930,N_6990);
nand U7075 (N_7075,N_6978,N_6980);
xnor U7076 (N_7076,N_6942,N_7026);
nor U7077 (N_7077,N_6939,N_7016);
or U7078 (N_7078,N_6983,N_6917);
nor U7079 (N_7079,N_7031,N_6992);
nor U7080 (N_7080,N_7002,N_6912);
xor U7081 (N_7081,N_7048,N_6955);
and U7082 (N_7082,N_6933,N_6937);
or U7083 (N_7083,N_7027,N_6974);
nand U7084 (N_7084,N_6960,N_7044);
nor U7085 (N_7085,N_7034,N_6941);
nor U7086 (N_7086,N_6936,N_7019);
and U7087 (N_7087,N_7006,N_7018);
nand U7088 (N_7088,N_7010,N_7014);
nand U7089 (N_7089,N_6966,N_6914);
nand U7090 (N_7090,N_7023,N_7025);
nor U7091 (N_7091,N_6970,N_6961);
xnor U7092 (N_7092,N_6900,N_6909);
nor U7093 (N_7093,N_7013,N_6952);
nand U7094 (N_7094,N_6976,N_6981);
nor U7095 (N_7095,N_7011,N_7029);
nor U7096 (N_7096,N_6958,N_6953);
xor U7097 (N_7097,N_6931,N_7032);
nand U7098 (N_7098,N_6906,N_6954);
nand U7099 (N_7099,N_6907,N_6988);
nand U7100 (N_7100,N_7015,N_7038);
nand U7101 (N_7101,N_6991,N_6922);
and U7102 (N_7102,N_6986,N_7043);
and U7103 (N_7103,N_6911,N_6929);
and U7104 (N_7104,N_6918,N_6924);
xor U7105 (N_7105,N_6940,N_7045);
xnor U7106 (N_7106,N_6994,N_6919);
nand U7107 (N_7107,N_6902,N_6946);
nand U7108 (N_7108,N_7047,N_6997);
and U7109 (N_7109,N_6903,N_6963);
and U7110 (N_7110,N_6938,N_6935);
and U7111 (N_7111,N_6948,N_7008);
xnor U7112 (N_7112,N_6916,N_6959);
and U7113 (N_7113,N_7039,N_6951);
nand U7114 (N_7114,N_6926,N_7028);
and U7115 (N_7115,N_7007,N_6947);
nand U7116 (N_7116,N_6962,N_7024);
nand U7117 (N_7117,N_6975,N_6982);
nand U7118 (N_7118,N_7049,N_7041);
or U7119 (N_7119,N_7021,N_6972);
or U7120 (N_7120,N_6956,N_6973);
xor U7121 (N_7121,N_6943,N_6985);
or U7122 (N_7122,N_7005,N_6925);
and U7123 (N_7123,N_6913,N_7022);
nand U7124 (N_7124,N_7020,N_6957);
or U7125 (N_7125,N_6994,N_6949);
or U7126 (N_7126,N_6970,N_7040);
or U7127 (N_7127,N_7011,N_7015);
nor U7128 (N_7128,N_6941,N_6997);
nor U7129 (N_7129,N_7039,N_6931);
nand U7130 (N_7130,N_6983,N_7036);
and U7131 (N_7131,N_6938,N_7001);
xor U7132 (N_7132,N_6968,N_6964);
nor U7133 (N_7133,N_6916,N_6995);
or U7134 (N_7134,N_7025,N_7046);
or U7135 (N_7135,N_6943,N_6969);
nand U7136 (N_7136,N_6997,N_7045);
and U7137 (N_7137,N_6927,N_6945);
nand U7138 (N_7138,N_6968,N_6910);
nor U7139 (N_7139,N_6948,N_7033);
or U7140 (N_7140,N_7045,N_6998);
nand U7141 (N_7141,N_7025,N_6931);
nor U7142 (N_7142,N_6964,N_6944);
or U7143 (N_7143,N_6993,N_6988);
nor U7144 (N_7144,N_7001,N_6912);
and U7145 (N_7145,N_6923,N_6926);
nor U7146 (N_7146,N_6902,N_6905);
or U7147 (N_7147,N_6996,N_7014);
nand U7148 (N_7148,N_6927,N_6938);
nor U7149 (N_7149,N_7024,N_6990);
nor U7150 (N_7150,N_7003,N_7025);
nand U7151 (N_7151,N_6990,N_7019);
and U7152 (N_7152,N_6910,N_7038);
and U7153 (N_7153,N_6963,N_6930);
and U7154 (N_7154,N_6901,N_6917);
or U7155 (N_7155,N_7022,N_7024);
nand U7156 (N_7156,N_6953,N_7037);
nor U7157 (N_7157,N_6991,N_7009);
or U7158 (N_7158,N_6905,N_6944);
xor U7159 (N_7159,N_6910,N_6991);
and U7160 (N_7160,N_6967,N_6902);
nand U7161 (N_7161,N_6950,N_7028);
nand U7162 (N_7162,N_6953,N_6999);
xor U7163 (N_7163,N_7020,N_7018);
and U7164 (N_7164,N_6941,N_6952);
nor U7165 (N_7165,N_7010,N_6949);
xor U7166 (N_7166,N_6924,N_6965);
xor U7167 (N_7167,N_6919,N_6959);
and U7168 (N_7168,N_6983,N_6999);
nor U7169 (N_7169,N_6979,N_6995);
and U7170 (N_7170,N_6990,N_6975);
or U7171 (N_7171,N_6918,N_6969);
and U7172 (N_7172,N_6923,N_6992);
and U7173 (N_7173,N_6965,N_7019);
and U7174 (N_7174,N_7039,N_6936);
or U7175 (N_7175,N_7003,N_6982);
xnor U7176 (N_7176,N_6954,N_6953);
xor U7177 (N_7177,N_6930,N_7026);
and U7178 (N_7178,N_6937,N_6913);
and U7179 (N_7179,N_7032,N_6995);
and U7180 (N_7180,N_7008,N_6904);
and U7181 (N_7181,N_6955,N_6904);
and U7182 (N_7182,N_7033,N_6929);
xor U7183 (N_7183,N_7007,N_6987);
or U7184 (N_7184,N_7000,N_6925);
nor U7185 (N_7185,N_6991,N_6964);
or U7186 (N_7186,N_7024,N_6910);
nand U7187 (N_7187,N_6978,N_7037);
and U7188 (N_7188,N_6994,N_6943);
xnor U7189 (N_7189,N_6952,N_7043);
and U7190 (N_7190,N_7001,N_6992);
xnor U7191 (N_7191,N_6955,N_7001);
and U7192 (N_7192,N_6913,N_7013);
and U7193 (N_7193,N_7030,N_6925);
and U7194 (N_7194,N_6947,N_6972);
and U7195 (N_7195,N_6952,N_6946);
nand U7196 (N_7196,N_6928,N_6939);
and U7197 (N_7197,N_6966,N_6974);
and U7198 (N_7198,N_6907,N_6908);
and U7199 (N_7199,N_6991,N_7048);
and U7200 (N_7200,N_7089,N_7167);
and U7201 (N_7201,N_7176,N_7172);
nor U7202 (N_7202,N_7066,N_7140);
and U7203 (N_7203,N_7179,N_7112);
nor U7204 (N_7204,N_7052,N_7150);
nand U7205 (N_7205,N_7165,N_7068);
nand U7206 (N_7206,N_7191,N_7080);
or U7207 (N_7207,N_7126,N_7163);
and U7208 (N_7208,N_7134,N_7155);
xnor U7209 (N_7209,N_7143,N_7103);
and U7210 (N_7210,N_7128,N_7161);
and U7211 (N_7211,N_7136,N_7056);
xor U7212 (N_7212,N_7147,N_7069);
nor U7213 (N_7213,N_7188,N_7197);
nor U7214 (N_7214,N_7109,N_7122);
nor U7215 (N_7215,N_7127,N_7100);
and U7216 (N_7216,N_7139,N_7146);
nor U7217 (N_7217,N_7116,N_7164);
or U7218 (N_7218,N_7120,N_7098);
nor U7219 (N_7219,N_7057,N_7123);
nor U7220 (N_7220,N_7158,N_7195);
and U7221 (N_7221,N_7105,N_7107);
and U7222 (N_7222,N_7153,N_7086);
nand U7223 (N_7223,N_7079,N_7177);
nor U7224 (N_7224,N_7131,N_7108);
nand U7225 (N_7225,N_7187,N_7111);
and U7226 (N_7226,N_7067,N_7106);
nor U7227 (N_7227,N_7169,N_7171);
or U7228 (N_7228,N_7117,N_7149);
nor U7229 (N_7229,N_7193,N_7118);
and U7230 (N_7230,N_7125,N_7144);
or U7231 (N_7231,N_7184,N_7054);
and U7232 (N_7232,N_7174,N_7119);
nand U7233 (N_7233,N_7115,N_7114);
nor U7234 (N_7234,N_7070,N_7138);
or U7235 (N_7235,N_7061,N_7186);
or U7236 (N_7236,N_7064,N_7137);
and U7237 (N_7237,N_7124,N_7190);
xnor U7238 (N_7238,N_7073,N_7074);
nand U7239 (N_7239,N_7183,N_7058);
nand U7240 (N_7240,N_7077,N_7053);
xnor U7241 (N_7241,N_7084,N_7078);
nand U7242 (N_7242,N_7159,N_7092);
xnor U7243 (N_7243,N_7059,N_7173);
and U7244 (N_7244,N_7083,N_7194);
and U7245 (N_7245,N_7180,N_7065);
nand U7246 (N_7246,N_7121,N_7170);
nor U7247 (N_7247,N_7091,N_7095);
nor U7248 (N_7248,N_7051,N_7063);
xnor U7249 (N_7249,N_7101,N_7182);
and U7250 (N_7250,N_7088,N_7130);
nand U7251 (N_7251,N_7189,N_7152);
nand U7252 (N_7252,N_7198,N_7175);
and U7253 (N_7253,N_7060,N_7132);
nor U7254 (N_7254,N_7097,N_7093);
and U7255 (N_7255,N_7090,N_7157);
nand U7256 (N_7256,N_7102,N_7062);
nand U7257 (N_7257,N_7178,N_7113);
nor U7258 (N_7258,N_7154,N_7055);
nand U7259 (N_7259,N_7142,N_7087);
nor U7260 (N_7260,N_7094,N_7168);
xnor U7261 (N_7261,N_7081,N_7082);
nand U7262 (N_7262,N_7076,N_7196);
xnor U7263 (N_7263,N_7085,N_7199);
nand U7264 (N_7264,N_7156,N_7104);
nand U7265 (N_7265,N_7071,N_7160);
xnor U7266 (N_7266,N_7141,N_7192);
xor U7267 (N_7267,N_7133,N_7151);
xnor U7268 (N_7268,N_7162,N_7166);
and U7269 (N_7269,N_7099,N_7145);
nand U7270 (N_7270,N_7185,N_7050);
or U7271 (N_7271,N_7110,N_7181);
and U7272 (N_7272,N_7135,N_7129);
xnor U7273 (N_7273,N_7072,N_7148);
nor U7274 (N_7274,N_7075,N_7096);
nor U7275 (N_7275,N_7076,N_7097);
or U7276 (N_7276,N_7179,N_7150);
and U7277 (N_7277,N_7075,N_7100);
and U7278 (N_7278,N_7107,N_7091);
xor U7279 (N_7279,N_7166,N_7195);
and U7280 (N_7280,N_7062,N_7169);
nor U7281 (N_7281,N_7176,N_7071);
nor U7282 (N_7282,N_7107,N_7128);
nand U7283 (N_7283,N_7127,N_7195);
xor U7284 (N_7284,N_7199,N_7105);
nand U7285 (N_7285,N_7152,N_7108);
nor U7286 (N_7286,N_7102,N_7192);
and U7287 (N_7287,N_7181,N_7136);
nand U7288 (N_7288,N_7114,N_7190);
nand U7289 (N_7289,N_7130,N_7059);
xnor U7290 (N_7290,N_7163,N_7140);
or U7291 (N_7291,N_7100,N_7162);
and U7292 (N_7292,N_7170,N_7171);
nand U7293 (N_7293,N_7071,N_7060);
nand U7294 (N_7294,N_7152,N_7053);
nor U7295 (N_7295,N_7083,N_7184);
or U7296 (N_7296,N_7060,N_7176);
or U7297 (N_7297,N_7094,N_7080);
nor U7298 (N_7298,N_7082,N_7117);
nor U7299 (N_7299,N_7052,N_7189);
and U7300 (N_7300,N_7131,N_7119);
nor U7301 (N_7301,N_7137,N_7173);
or U7302 (N_7302,N_7053,N_7093);
nand U7303 (N_7303,N_7191,N_7067);
and U7304 (N_7304,N_7122,N_7076);
and U7305 (N_7305,N_7074,N_7093);
nor U7306 (N_7306,N_7155,N_7147);
and U7307 (N_7307,N_7189,N_7127);
or U7308 (N_7308,N_7115,N_7150);
and U7309 (N_7309,N_7197,N_7170);
nand U7310 (N_7310,N_7087,N_7082);
and U7311 (N_7311,N_7113,N_7108);
nor U7312 (N_7312,N_7111,N_7105);
xor U7313 (N_7313,N_7064,N_7109);
xor U7314 (N_7314,N_7074,N_7137);
nor U7315 (N_7315,N_7078,N_7131);
and U7316 (N_7316,N_7198,N_7179);
or U7317 (N_7317,N_7175,N_7073);
nor U7318 (N_7318,N_7054,N_7168);
nand U7319 (N_7319,N_7135,N_7118);
and U7320 (N_7320,N_7075,N_7081);
or U7321 (N_7321,N_7103,N_7058);
and U7322 (N_7322,N_7162,N_7071);
xor U7323 (N_7323,N_7113,N_7072);
and U7324 (N_7324,N_7134,N_7061);
xor U7325 (N_7325,N_7102,N_7163);
nor U7326 (N_7326,N_7129,N_7077);
nand U7327 (N_7327,N_7115,N_7105);
nand U7328 (N_7328,N_7054,N_7176);
nor U7329 (N_7329,N_7127,N_7071);
and U7330 (N_7330,N_7094,N_7198);
nor U7331 (N_7331,N_7193,N_7191);
and U7332 (N_7332,N_7143,N_7064);
or U7333 (N_7333,N_7194,N_7139);
or U7334 (N_7334,N_7191,N_7185);
and U7335 (N_7335,N_7118,N_7055);
nor U7336 (N_7336,N_7153,N_7179);
or U7337 (N_7337,N_7119,N_7050);
xor U7338 (N_7338,N_7104,N_7134);
or U7339 (N_7339,N_7150,N_7169);
xnor U7340 (N_7340,N_7198,N_7071);
xnor U7341 (N_7341,N_7127,N_7056);
nor U7342 (N_7342,N_7114,N_7085);
nand U7343 (N_7343,N_7105,N_7123);
nand U7344 (N_7344,N_7072,N_7134);
and U7345 (N_7345,N_7173,N_7156);
xor U7346 (N_7346,N_7096,N_7154);
or U7347 (N_7347,N_7198,N_7166);
nor U7348 (N_7348,N_7061,N_7191);
and U7349 (N_7349,N_7092,N_7079);
nor U7350 (N_7350,N_7245,N_7277);
nand U7351 (N_7351,N_7230,N_7334);
nand U7352 (N_7352,N_7325,N_7235);
nor U7353 (N_7353,N_7328,N_7255);
nand U7354 (N_7354,N_7345,N_7201);
or U7355 (N_7355,N_7200,N_7215);
or U7356 (N_7356,N_7335,N_7257);
nand U7357 (N_7357,N_7224,N_7265);
nor U7358 (N_7358,N_7209,N_7264);
or U7359 (N_7359,N_7207,N_7319);
or U7360 (N_7360,N_7218,N_7300);
nor U7361 (N_7361,N_7336,N_7287);
nand U7362 (N_7362,N_7214,N_7327);
or U7363 (N_7363,N_7347,N_7253);
nor U7364 (N_7364,N_7221,N_7290);
or U7365 (N_7365,N_7315,N_7252);
nand U7366 (N_7366,N_7323,N_7313);
nor U7367 (N_7367,N_7250,N_7217);
nand U7368 (N_7368,N_7332,N_7339);
xor U7369 (N_7369,N_7274,N_7241);
nand U7370 (N_7370,N_7249,N_7340);
xnor U7371 (N_7371,N_7232,N_7322);
and U7372 (N_7372,N_7304,N_7329);
nor U7373 (N_7373,N_7278,N_7279);
or U7374 (N_7374,N_7211,N_7229);
nor U7375 (N_7375,N_7237,N_7247);
nand U7376 (N_7376,N_7318,N_7248);
nor U7377 (N_7377,N_7280,N_7321);
nor U7378 (N_7378,N_7288,N_7251);
nand U7379 (N_7379,N_7282,N_7244);
xnor U7380 (N_7380,N_7285,N_7305);
nor U7381 (N_7381,N_7291,N_7310);
nor U7382 (N_7382,N_7276,N_7337);
nand U7383 (N_7383,N_7240,N_7295);
nand U7384 (N_7384,N_7296,N_7260);
or U7385 (N_7385,N_7243,N_7317);
xor U7386 (N_7386,N_7349,N_7231);
nand U7387 (N_7387,N_7292,N_7326);
nand U7388 (N_7388,N_7269,N_7294);
nand U7389 (N_7389,N_7220,N_7271);
and U7390 (N_7390,N_7343,N_7342);
or U7391 (N_7391,N_7284,N_7289);
nand U7392 (N_7392,N_7216,N_7263);
and U7393 (N_7393,N_7307,N_7314);
nor U7394 (N_7394,N_7205,N_7286);
and U7395 (N_7395,N_7301,N_7259);
and U7396 (N_7396,N_7203,N_7258);
xnor U7397 (N_7397,N_7204,N_7303);
xor U7398 (N_7398,N_7306,N_7338);
and U7399 (N_7399,N_7256,N_7239);
nand U7400 (N_7400,N_7206,N_7312);
or U7401 (N_7401,N_7228,N_7297);
and U7402 (N_7402,N_7261,N_7299);
nand U7403 (N_7403,N_7270,N_7234);
and U7404 (N_7404,N_7330,N_7236);
xnor U7405 (N_7405,N_7272,N_7341);
and U7406 (N_7406,N_7281,N_7316);
nand U7407 (N_7407,N_7283,N_7309);
or U7408 (N_7408,N_7223,N_7275);
nand U7409 (N_7409,N_7308,N_7227);
and U7410 (N_7410,N_7333,N_7210);
nor U7411 (N_7411,N_7268,N_7346);
and U7412 (N_7412,N_7298,N_7202);
nor U7413 (N_7413,N_7302,N_7225);
xor U7414 (N_7414,N_7266,N_7324);
nand U7415 (N_7415,N_7219,N_7246);
or U7416 (N_7416,N_7208,N_7273);
nor U7417 (N_7417,N_7293,N_7348);
nor U7418 (N_7418,N_7262,N_7226);
nand U7419 (N_7419,N_7331,N_7254);
nor U7420 (N_7420,N_7212,N_7238);
and U7421 (N_7421,N_7233,N_7311);
or U7422 (N_7422,N_7267,N_7320);
nor U7423 (N_7423,N_7213,N_7242);
and U7424 (N_7424,N_7222,N_7344);
or U7425 (N_7425,N_7213,N_7343);
nand U7426 (N_7426,N_7329,N_7231);
or U7427 (N_7427,N_7268,N_7298);
or U7428 (N_7428,N_7349,N_7275);
nand U7429 (N_7429,N_7280,N_7217);
or U7430 (N_7430,N_7261,N_7203);
nand U7431 (N_7431,N_7245,N_7267);
nor U7432 (N_7432,N_7332,N_7289);
and U7433 (N_7433,N_7320,N_7200);
nand U7434 (N_7434,N_7233,N_7237);
xnor U7435 (N_7435,N_7270,N_7335);
nor U7436 (N_7436,N_7333,N_7242);
nor U7437 (N_7437,N_7249,N_7314);
xor U7438 (N_7438,N_7302,N_7324);
nor U7439 (N_7439,N_7252,N_7321);
nor U7440 (N_7440,N_7202,N_7253);
xnor U7441 (N_7441,N_7277,N_7255);
or U7442 (N_7442,N_7293,N_7318);
and U7443 (N_7443,N_7255,N_7204);
nor U7444 (N_7444,N_7338,N_7314);
nor U7445 (N_7445,N_7344,N_7217);
xnor U7446 (N_7446,N_7227,N_7255);
and U7447 (N_7447,N_7234,N_7266);
nand U7448 (N_7448,N_7272,N_7208);
xor U7449 (N_7449,N_7252,N_7337);
and U7450 (N_7450,N_7345,N_7269);
and U7451 (N_7451,N_7310,N_7325);
or U7452 (N_7452,N_7225,N_7210);
nor U7453 (N_7453,N_7298,N_7280);
or U7454 (N_7454,N_7347,N_7249);
nand U7455 (N_7455,N_7263,N_7306);
and U7456 (N_7456,N_7305,N_7317);
or U7457 (N_7457,N_7324,N_7205);
and U7458 (N_7458,N_7221,N_7311);
nor U7459 (N_7459,N_7203,N_7213);
nand U7460 (N_7460,N_7323,N_7200);
and U7461 (N_7461,N_7263,N_7331);
and U7462 (N_7462,N_7205,N_7201);
nand U7463 (N_7463,N_7280,N_7334);
nor U7464 (N_7464,N_7313,N_7279);
and U7465 (N_7465,N_7207,N_7253);
and U7466 (N_7466,N_7335,N_7225);
or U7467 (N_7467,N_7244,N_7223);
nand U7468 (N_7468,N_7227,N_7307);
or U7469 (N_7469,N_7261,N_7341);
and U7470 (N_7470,N_7303,N_7342);
nor U7471 (N_7471,N_7271,N_7327);
and U7472 (N_7472,N_7277,N_7243);
and U7473 (N_7473,N_7206,N_7320);
or U7474 (N_7474,N_7294,N_7246);
or U7475 (N_7475,N_7252,N_7261);
nand U7476 (N_7476,N_7337,N_7317);
nor U7477 (N_7477,N_7299,N_7204);
nor U7478 (N_7478,N_7301,N_7275);
xor U7479 (N_7479,N_7262,N_7326);
and U7480 (N_7480,N_7305,N_7219);
xnor U7481 (N_7481,N_7286,N_7214);
and U7482 (N_7482,N_7214,N_7244);
nand U7483 (N_7483,N_7283,N_7330);
xnor U7484 (N_7484,N_7345,N_7334);
and U7485 (N_7485,N_7297,N_7315);
and U7486 (N_7486,N_7216,N_7331);
xor U7487 (N_7487,N_7288,N_7250);
and U7488 (N_7488,N_7323,N_7234);
xor U7489 (N_7489,N_7212,N_7201);
or U7490 (N_7490,N_7305,N_7341);
and U7491 (N_7491,N_7201,N_7348);
or U7492 (N_7492,N_7324,N_7321);
or U7493 (N_7493,N_7312,N_7210);
and U7494 (N_7494,N_7250,N_7201);
nand U7495 (N_7495,N_7243,N_7348);
nor U7496 (N_7496,N_7229,N_7239);
or U7497 (N_7497,N_7295,N_7213);
or U7498 (N_7498,N_7215,N_7339);
nor U7499 (N_7499,N_7289,N_7298);
or U7500 (N_7500,N_7476,N_7429);
xnor U7501 (N_7501,N_7371,N_7498);
and U7502 (N_7502,N_7414,N_7456);
nor U7503 (N_7503,N_7353,N_7389);
and U7504 (N_7504,N_7404,N_7385);
and U7505 (N_7505,N_7352,N_7433);
nand U7506 (N_7506,N_7441,N_7478);
nand U7507 (N_7507,N_7426,N_7446);
and U7508 (N_7508,N_7401,N_7484);
and U7509 (N_7509,N_7378,N_7388);
xnor U7510 (N_7510,N_7440,N_7387);
nor U7511 (N_7511,N_7485,N_7483);
and U7512 (N_7512,N_7491,N_7434);
nand U7513 (N_7513,N_7412,N_7422);
xor U7514 (N_7514,N_7415,N_7374);
or U7515 (N_7515,N_7448,N_7355);
nor U7516 (N_7516,N_7410,N_7370);
nand U7517 (N_7517,N_7480,N_7470);
nand U7518 (N_7518,N_7396,N_7418);
nor U7519 (N_7519,N_7390,N_7377);
nor U7520 (N_7520,N_7425,N_7454);
nor U7521 (N_7521,N_7407,N_7488);
xnor U7522 (N_7522,N_7447,N_7361);
nand U7523 (N_7523,N_7357,N_7457);
nor U7524 (N_7524,N_7499,N_7375);
xor U7525 (N_7525,N_7413,N_7458);
nand U7526 (N_7526,N_7462,N_7427);
and U7527 (N_7527,N_7399,N_7445);
or U7528 (N_7528,N_7459,N_7438);
and U7529 (N_7529,N_7360,N_7432);
or U7530 (N_7530,N_7394,N_7487);
nor U7531 (N_7531,N_7467,N_7461);
nor U7532 (N_7532,N_7469,N_7479);
nand U7533 (N_7533,N_7493,N_7419);
nor U7534 (N_7534,N_7442,N_7383);
and U7535 (N_7535,N_7406,N_7443);
nand U7536 (N_7536,N_7372,N_7356);
nor U7537 (N_7537,N_7359,N_7451);
or U7538 (N_7538,N_7450,N_7421);
or U7539 (N_7539,N_7449,N_7382);
nand U7540 (N_7540,N_7452,N_7354);
nand U7541 (N_7541,N_7477,N_7475);
or U7542 (N_7542,N_7474,N_7397);
xor U7543 (N_7543,N_7492,N_7366);
nand U7544 (N_7544,N_7490,N_7365);
and U7545 (N_7545,N_7379,N_7496);
xor U7546 (N_7546,N_7391,N_7350);
and U7547 (N_7547,N_7453,N_7398);
and U7548 (N_7548,N_7369,N_7436);
nor U7549 (N_7549,N_7403,N_7494);
nor U7550 (N_7550,N_7393,N_7482);
nand U7551 (N_7551,N_7381,N_7455);
nand U7552 (N_7552,N_7380,N_7358);
nand U7553 (N_7553,N_7428,N_7463);
nor U7554 (N_7554,N_7435,N_7411);
nor U7555 (N_7555,N_7437,N_7468);
or U7556 (N_7556,N_7400,N_7416);
nor U7557 (N_7557,N_7431,N_7409);
and U7558 (N_7558,N_7423,N_7466);
nand U7559 (N_7559,N_7464,N_7489);
nand U7560 (N_7560,N_7486,N_7376);
xnor U7561 (N_7561,N_7497,N_7368);
and U7562 (N_7562,N_7471,N_7424);
and U7563 (N_7563,N_7408,N_7373);
nor U7564 (N_7564,N_7363,N_7367);
and U7565 (N_7565,N_7439,N_7402);
nand U7566 (N_7566,N_7444,N_7417);
or U7567 (N_7567,N_7473,N_7472);
nand U7568 (N_7568,N_7384,N_7351);
nand U7569 (N_7569,N_7460,N_7495);
nor U7570 (N_7570,N_7362,N_7395);
nor U7571 (N_7571,N_7481,N_7405);
or U7572 (N_7572,N_7392,N_7420);
and U7573 (N_7573,N_7465,N_7430);
and U7574 (N_7574,N_7364,N_7386);
and U7575 (N_7575,N_7429,N_7384);
nor U7576 (N_7576,N_7374,N_7351);
nand U7577 (N_7577,N_7380,N_7446);
xor U7578 (N_7578,N_7480,N_7368);
or U7579 (N_7579,N_7489,N_7468);
and U7580 (N_7580,N_7492,N_7469);
or U7581 (N_7581,N_7367,N_7492);
nor U7582 (N_7582,N_7359,N_7457);
or U7583 (N_7583,N_7462,N_7486);
nand U7584 (N_7584,N_7364,N_7409);
or U7585 (N_7585,N_7374,N_7378);
or U7586 (N_7586,N_7484,N_7422);
and U7587 (N_7587,N_7499,N_7478);
nor U7588 (N_7588,N_7449,N_7436);
nor U7589 (N_7589,N_7400,N_7496);
nand U7590 (N_7590,N_7440,N_7446);
nor U7591 (N_7591,N_7445,N_7384);
nor U7592 (N_7592,N_7472,N_7487);
nor U7593 (N_7593,N_7402,N_7495);
nand U7594 (N_7594,N_7397,N_7470);
nand U7595 (N_7595,N_7443,N_7488);
or U7596 (N_7596,N_7486,N_7444);
and U7597 (N_7597,N_7385,N_7398);
nor U7598 (N_7598,N_7467,N_7488);
and U7599 (N_7599,N_7389,N_7486);
nor U7600 (N_7600,N_7389,N_7387);
nor U7601 (N_7601,N_7371,N_7384);
nand U7602 (N_7602,N_7457,N_7454);
or U7603 (N_7603,N_7405,N_7439);
or U7604 (N_7604,N_7459,N_7414);
nor U7605 (N_7605,N_7479,N_7365);
xnor U7606 (N_7606,N_7443,N_7435);
nor U7607 (N_7607,N_7474,N_7415);
nor U7608 (N_7608,N_7484,N_7458);
or U7609 (N_7609,N_7489,N_7373);
and U7610 (N_7610,N_7392,N_7428);
or U7611 (N_7611,N_7366,N_7447);
nor U7612 (N_7612,N_7354,N_7400);
or U7613 (N_7613,N_7471,N_7413);
nor U7614 (N_7614,N_7375,N_7415);
nand U7615 (N_7615,N_7378,N_7442);
nand U7616 (N_7616,N_7357,N_7448);
nand U7617 (N_7617,N_7498,N_7355);
or U7618 (N_7618,N_7444,N_7453);
nor U7619 (N_7619,N_7390,N_7498);
nand U7620 (N_7620,N_7489,N_7463);
nand U7621 (N_7621,N_7383,N_7369);
or U7622 (N_7622,N_7383,N_7406);
and U7623 (N_7623,N_7428,N_7378);
nand U7624 (N_7624,N_7469,N_7436);
xnor U7625 (N_7625,N_7498,N_7478);
or U7626 (N_7626,N_7495,N_7421);
nor U7627 (N_7627,N_7426,N_7367);
nand U7628 (N_7628,N_7473,N_7424);
or U7629 (N_7629,N_7476,N_7390);
or U7630 (N_7630,N_7467,N_7415);
or U7631 (N_7631,N_7386,N_7350);
or U7632 (N_7632,N_7419,N_7494);
xor U7633 (N_7633,N_7495,N_7364);
nor U7634 (N_7634,N_7365,N_7389);
nor U7635 (N_7635,N_7455,N_7369);
xnor U7636 (N_7636,N_7438,N_7448);
nor U7637 (N_7637,N_7492,N_7459);
nor U7638 (N_7638,N_7437,N_7389);
nor U7639 (N_7639,N_7484,N_7408);
or U7640 (N_7640,N_7449,N_7423);
xor U7641 (N_7641,N_7392,N_7487);
xnor U7642 (N_7642,N_7406,N_7449);
and U7643 (N_7643,N_7358,N_7441);
or U7644 (N_7644,N_7483,N_7475);
or U7645 (N_7645,N_7428,N_7493);
or U7646 (N_7646,N_7354,N_7375);
nor U7647 (N_7647,N_7404,N_7397);
xor U7648 (N_7648,N_7393,N_7495);
nor U7649 (N_7649,N_7403,N_7401);
nand U7650 (N_7650,N_7560,N_7513);
and U7651 (N_7651,N_7540,N_7571);
nor U7652 (N_7652,N_7623,N_7503);
and U7653 (N_7653,N_7548,N_7567);
and U7654 (N_7654,N_7628,N_7642);
nor U7655 (N_7655,N_7529,N_7509);
or U7656 (N_7656,N_7616,N_7608);
and U7657 (N_7657,N_7520,N_7624);
and U7658 (N_7658,N_7576,N_7578);
or U7659 (N_7659,N_7588,N_7577);
nand U7660 (N_7660,N_7639,N_7641);
nand U7661 (N_7661,N_7627,N_7522);
nand U7662 (N_7662,N_7581,N_7603);
nor U7663 (N_7663,N_7533,N_7561);
nand U7664 (N_7664,N_7580,N_7619);
nand U7665 (N_7665,N_7600,N_7640);
nor U7666 (N_7666,N_7506,N_7618);
or U7667 (N_7667,N_7589,N_7620);
and U7668 (N_7668,N_7539,N_7644);
or U7669 (N_7669,N_7635,N_7518);
nand U7670 (N_7670,N_7617,N_7564);
nand U7671 (N_7671,N_7629,N_7528);
and U7672 (N_7672,N_7647,N_7634);
nor U7673 (N_7673,N_7582,N_7557);
xnor U7674 (N_7674,N_7625,N_7558);
and U7675 (N_7675,N_7643,N_7555);
or U7676 (N_7676,N_7607,N_7579);
or U7677 (N_7677,N_7559,N_7547);
and U7678 (N_7678,N_7584,N_7586);
and U7679 (N_7679,N_7645,N_7554);
nand U7680 (N_7680,N_7638,N_7596);
or U7681 (N_7681,N_7595,N_7510);
or U7682 (N_7682,N_7501,N_7553);
nor U7683 (N_7683,N_7572,N_7609);
nand U7684 (N_7684,N_7614,N_7562);
and U7685 (N_7685,N_7532,N_7519);
nor U7686 (N_7686,N_7621,N_7622);
xor U7687 (N_7687,N_7626,N_7505);
and U7688 (N_7688,N_7502,N_7597);
or U7689 (N_7689,N_7527,N_7605);
nand U7690 (N_7690,N_7537,N_7552);
nand U7691 (N_7691,N_7610,N_7538);
nand U7692 (N_7692,N_7546,N_7556);
nor U7693 (N_7693,N_7512,N_7568);
nor U7694 (N_7694,N_7525,N_7604);
xnor U7695 (N_7695,N_7631,N_7646);
nor U7696 (N_7696,N_7648,N_7599);
and U7697 (N_7697,N_7536,N_7602);
and U7698 (N_7698,N_7574,N_7598);
xor U7699 (N_7699,N_7535,N_7613);
nor U7700 (N_7700,N_7514,N_7592);
or U7701 (N_7701,N_7515,N_7585);
xnor U7702 (N_7702,N_7551,N_7570);
and U7703 (N_7703,N_7534,N_7508);
and U7704 (N_7704,N_7593,N_7611);
and U7705 (N_7705,N_7531,N_7507);
and U7706 (N_7706,N_7563,N_7517);
or U7707 (N_7707,N_7615,N_7612);
nor U7708 (N_7708,N_7569,N_7575);
nand U7709 (N_7709,N_7630,N_7583);
nand U7710 (N_7710,N_7542,N_7566);
and U7711 (N_7711,N_7565,N_7636);
nor U7712 (N_7712,N_7573,N_7587);
and U7713 (N_7713,N_7594,N_7526);
and U7714 (N_7714,N_7632,N_7541);
and U7715 (N_7715,N_7601,N_7523);
or U7716 (N_7716,N_7549,N_7524);
or U7717 (N_7717,N_7633,N_7606);
and U7718 (N_7718,N_7511,N_7550);
xor U7719 (N_7719,N_7521,N_7591);
nand U7720 (N_7720,N_7504,N_7543);
nand U7721 (N_7721,N_7590,N_7544);
xor U7722 (N_7722,N_7545,N_7637);
or U7723 (N_7723,N_7500,N_7530);
and U7724 (N_7724,N_7516,N_7649);
nor U7725 (N_7725,N_7536,N_7542);
or U7726 (N_7726,N_7633,N_7593);
or U7727 (N_7727,N_7594,N_7598);
and U7728 (N_7728,N_7582,N_7520);
nand U7729 (N_7729,N_7567,N_7536);
nand U7730 (N_7730,N_7649,N_7533);
nand U7731 (N_7731,N_7638,N_7558);
or U7732 (N_7732,N_7522,N_7595);
and U7733 (N_7733,N_7573,N_7584);
nor U7734 (N_7734,N_7516,N_7543);
nor U7735 (N_7735,N_7526,N_7570);
or U7736 (N_7736,N_7591,N_7585);
and U7737 (N_7737,N_7594,N_7601);
and U7738 (N_7738,N_7541,N_7567);
or U7739 (N_7739,N_7559,N_7635);
nand U7740 (N_7740,N_7535,N_7626);
xnor U7741 (N_7741,N_7587,N_7526);
and U7742 (N_7742,N_7530,N_7505);
xnor U7743 (N_7743,N_7519,N_7612);
nor U7744 (N_7744,N_7543,N_7614);
xnor U7745 (N_7745,N_7579,N_7523);
and U7746 (N_7746,N_7536,N_7582);
nand U7747 (N_7747,N_7576,N_7518);
nor U7748 (N_7748,N_7588,N_7513);
nand U7749 (N_7749,N_7591,N_7541);
and U7750 (N_7750,N_7553,N_7627);
or U7751 (N_7751,N_7605,N_7611);
nor U7752 (N_7752,N_7555,N_7517);
nor U7753 (N_7753,N_7545,N_7524);
xor U7754 (N_7754,N_7561,N_7598);
or U7755 (N_7755,N_7567,N_7633);
nand U7756 (N_7756,N_7567,N_7600);
or U7757 (N_7757,N_7603,N_7539);
and U7758 (N_7758,N_7640,N_7533);
nand U7759 (N_7759,N_7581,N_7604);
or U7760 (N_7760,N_7643,N_7621);
nor U7761 (N_7761,N_7629,N_7598);
or U7762 (N_7762,N_7613,N_7625);
or U7763 (N_7763,N_7617,N_7515);
and U7764 (N_7764,N_7588,N_7533);
and U7765 (N_7765,N_7626,N_7606);
nand U7766 (N_7766,N_7555,N_7607);
and U7767 (N_7767,N_7616,N_7518);
and U7768 (N_7768,N_7602,N_7531);
and U7769 (N_7769,N_7621,N_7593);
nor U7770 (N_7770,N_7649,N_7528);
nand U7771 (N_7771,N_7581,N_7628);
xnor U7772 (N_7772,N_7630,N_7584);
and U7773 (N_7773,N_7614,N_7566);
nand U7774 (N_7774,N_7620,N_7622);
nor U7775 (N_7775,N_7647,N_7500);
nand U7776 (N_7776,N_7536,N_7616);
and U7777 (N_7777,N_7639,N_7612);
or U7778 (N_7778,N_7521,N_7644);
xnor U7779 (N_7779,N_7570,N_7615);
or U7780 (N_7780,N_7624,N_7606);
nand U7781 (N_7781,N_7513,N_7583);
xnor U7782 (N_7782,N_7641,N_7518);
or U7783 (N_7783,N_7580,N_7608);
xor U7784 (N_7784,N_7549,N_7611);
and U7785 (N_7785,N_7594,N_7634);
or U7786 (N_7786,N_7552,N_7587);
nand U7787 (N_7787,N_7501,N_7621);
nor U7788 (N_7788,N_7517,N_7580);
nor U7789 (N_7789,N_7555,N_7576);
xnor U7790 (N_7790,N_7592,N_7601);
nand U7791 (N_7791,N_7637,N_7571);
nor U7792 (N_7792,N_7528,N_7512);
nand U7793 (N_7793,N_7515,N_7526);
and U7794 (N_7794,N_7590,N_7545);
or U7795 (N_7795,N_7606,N_7514);
nand U7796 (N_7796,N_7614,N_7542);
or U7797 (N_7797,N_7625,N_7572);
nand U7798 (N_7798,N_7611,N_7572);
nand U7799 (N_7799,N_7645,N_7542);
nand U7800 (N_7800,N_7757,N_7691);
or U7801 (N_7801,N_7708,N_7772);
and U7802 (N_7802,N_7786,N_7660);
and U7803 (N_7803,N_7732,N_7699);
or U7804 (N_7804,N_7693,N_7687);
nand U7805 (N_7805,N_7696,N_7725);
nor U7806 (N_7806,N_7743,N_7695);
nor U7807 (N_7807,N_7773,N_7728);
nor U7808 (N_7808,N_7763,N_7777);
or U7809 (N_7809,N_7726,N_7770);
nand U7810 (N_7810,N_7740,N_7710);
and U7811 (N_7811,N_7741,N_7657);
and U7812 (N_7812,N_7766,N_7672);
xor U7813 (N_7813,N_7659,N_7790);
nor U7814 (N_7814,N_7731,N_7735);
or U7815 (N_7815,N_7717,N_7679);
or U7816 (N_7816,N_7656,N_7650);
xnor U7817 (N_7817,N_7767,N_7780);
nand U7818 (N_7818,N_7667,N_7704);
and U7819 (N_7819,N_7745,N_7733);
xnor U7820 (N_7820,N_7689,N_7668);
or U7821 (N_7821,N_7700,N_7769);
nor U7822 (N_7822,N_7654,N_7782);
xor U7823 (N_7823,N_7738,N_7799);
or U7824 (N_7824,N_7758,N_7669);
nand U7825 (N_7825,N_7694,N_7755);
nand U7826 (N_7826,N_7764,N_7688);
nor U7827 (N_7827,N_7662,N_7722);
and U7828 (N_7828,N_7661,N_7734);
and U7829 (N_7829,N_7759,N_7666);
nand U7830 (N_7830,N_7751,N_7754);
and U7831 (N_7831,N_7697,N_7705);
or U7832 (N_7832,N_7765,N_7664);
nand U7833 (N_7833,N_7736,N_7761);
or U7834 (N_7834,N_7658,N_7762);
and U7835 (N_7835,N_7787,N_7748);
nand U7836 (N_7836,N_7682,N_7724);
nor U7837 (N_7837,N_7683,N_7715);
nand U7838 (N_7838,N_7709,N_7670);
nor U7839 (N_7839,N_7655,N_7652);
nand U7840 (N_7840,N_7680,N_7749);
and U7841 (N_7841,N_7727,N_7676);
nand U7842 (N_7842,N_7747,N_7685);
xnor U7843 (N_7843,N_7713,N_7692);
or U7844 (N_7844,N_7684,N_7718);
nand U7845 (N_7845,N_7796,N_7785);
nand U7846 (N_7846,N_7737,N_7720);
nand U7847 (N_7847,N_7703,N_7663);
and U7848 (N_7848,N_7714,N_7794);
or U7849 (N_7849,N_7702,N_7673);
and U7850 (N_7850,N_7678,N_7760);
and U7851 (N_7851,N_7776,N_7698);
xor U7852 (N_7852,N_7716,N_7779);
and U7853 (N_7853,N_7729,N_7753);
and U7854 (N_7854,N_7721,N_7771);
xnor U7855 (N_7855,N_7730,N_7723);
nor U7856 (N_7856,N_7671,N_7707);
and U7857 (N_7857,N_7752,N_7653);
nand U7858 (N_7858,N_7744,N_7719);
nand U7859 (N_7859,N_7778,N_7795);
nor U7860 (N_7860,N_7783,N_7768);
nand U7861 (N_7861,N_7797,N_7789);
and U7862 (N_7862,N_7665,N_7686);
or U7863 (N_7863,N_7791,N_7675);
nor U7864 (N_7864,N_7674,N_7701);
nor U7865 (N_7865,N_7681,N_7739);
nor U7866 (N_7866,N_7784,N_7788);
or U7867 (N_7867,N_7774,N_7651);
nand U7868 (N_7868,N_7706,N_7690);
and U7869 (N_7869,N_7711,N_7798);
nor U7870 (N_7870,N_7793,N_7781);
nor U7871 (N_7871,N_7792,N_7742);
nand U7872 (N_7872,N_7775,N_7756);
nor U7873 (N_7873,N_7746,N_7677);
nor U7874 (N_7874,N_7750,N_7712);
or U7875 (N_7875,N_7748,N_7798);
nor U7876 (N_7876,N_7658,N_7721);
or U7877 (N_7877,N_7665,N_7769);
nor U7878 (N_7878,N_7791,N_7747);
or U7879 (N_7879,N_7782,N_7679);
nor U7880 (N_7880,N_7787,N_7754);
xnor U7881 (N_7881,N_7756,N_7739);
and U7882 (N_7882,N_7774,N_7738);
nand U7883 (N_7883,N_7697,N_7776);
and U7884 (N_7884,N_7736,N_7728);
nor U7885 (N_7885,N_7781,N_7751);
xnor U7886 (N_7886,N_7661,N_7671);
nor U7887 (N_7887,N_7731,N_7714);
and U7888 (N_7888,N_7671,N_7734);
and U7889 (N_7889,N_7749,N_7716);
nor U7890 (N_7890,N_7650,N_7678);
nand U7891 (N_7891,N_7669,N_7695);
nor U7892 (N_7892,N_7662,N_7712);
and U7893 (N_7893,N_7742,N_7750);
and U7894 (N_7894,N_7678,N_7667);
nand U7895 (N_7895,N_7675,N_7704);
or U7896 (N_7896,N_7760,N_7751);
nand U7897 (N_7897,N_7747,N_7795);
nand U7898 (N_7898,N_7746,N_7760);
nand U7899 (N_7899,N_7668,N_7781);
nor U7900 (N_7900,N_7750,N_7753);
xnor U7901 (N_7901,N_7749,N_7671);
nor U7902 (N_7902,N_7667,N_7745);
and U7903 (N_7903,N_7701,N_7730);
or U7904 (N_7904,N_7655,N_7699);
and U7905 (N_7905,N_7696,N_7693);
nor U7906 (N_7906,N_7777,N_7666);
or U7907 (N_7907,N_7728,N_7755);
nand U7908 (N_7908,N_7687,N_7714);
or U7909 (N_7909,N_7693,N_7731);
nand U7910 (N_7910,N_7766,N_7789);
nand U7911 (N_7911,N_7665,N_7760);
nor U7912 (N_7912,N_7721,N_7753);
nand U7913 (N_7913,N_7788,N_7677);
or U7914 (N_7914,N_7799,N_7771);
or U7915 (N_7915,N_7703,N_7793);
or U7916 (N_7916,N_7673,N_7655);
and U7917 (N_7917,N_7776,N_7666);
and U7918 (N_7918,N_7789,N_7659);
and U7919 (N_7919,N_7723,N_7673);
nor U7920 (N_7920,N_7657,N_7778);
nand U7921 (N_7921,N_7730,N_7703);
nand U7922 (N_7922,N_7765,N_7772);
xnor U7923 (N_7923,N_7670,N_7712);
or U7924 (N_7924,N_7756,N_7697);
nor U7925 (N_7925,N_7788,N_7717);
or U7926 (N_7926,N_7745,N_7710);
nand U7927 (N_7927,N_7691,N_7733);
nand U7928 (N_7928,N_7712,N_7652);
and U7929 (N_7929,N_7783,N_7740);
or U7930 (N_7930,N_7785,N_7713);
or U7931 (N_7931,N_7667,N_7782);
nor U7932 (N_7932,N_7709,N_7711);
xor U7933 (N_7933,N_7689,N_7711);
and U7934 (N_7934,N_7754,N_7673);
or U7935 (N_7935,N_7701,N_7668);
xnor U7936 (N_7936,N_7713,N_7738);
nand U7937 (N_7937,N_7749,N_7715);
nand U7938 (N_7938,N_7741,N_7721);
nand U7939 (N_7939,N_7710,N_7705);
or U7940 (N_7940,N_7781,N_7725);
or U7941 (N_7941,N_7725,N_7788);
nor U7942 (N_7942,N_7736,N_7715);
nand U7943 (N_7943,N_7728,N_7720);
or U7944 (N_7944,N_7721,N_7698);
nand U7945 (N_7945,N_7724,N_7741);
and U7946 (N_7946,N_7777,N_7723);
or U7947 (N_7947,N_7664,N_7742);
or U7948 (N_7948,N_7709,N_7798);
nand U7949 (N_7949,N_7677,N_7741);
xnor U7950 (N_7950,N_7943,N_7938);
nand U7951 (N_7951,N_7827,N_7907);
xor U7952 (N_7952,N_7927,N_7912);
nand U7953 (N_7953,N_7930,N_7863);
nand U7954 (N_7954,N_7914,N_7920);
xnor U7955 (N_7955,N_7874,N_7910);
nor U7956 (N_7956,N_7859,N_7901);
xnor U7957 (N_7957,N_7828,N_7932);
nor U7958 (N_7958,N_7866,N_7842);
or U7959 (N_7959,N_7881,N_7856);
and U7960 (N_7960,N_7804,N_7861);
and U7961 (N_7961,N_7806,N_7857);
nand U7962 (N_7962,N_7825,N_7902);
or U7963 (N_7963,N_7811,N_7948);
and U7964 (N_7964,N_7869,N_7879);
nor U7965 (N_7965,N_7885,N_7872);
nand U7966 (N_7966,N_7936,N_7846);
nand U7967 (N_7967,N_7941,N_7864);
nand U7968 (N_7968,N_7934,N_7925);
or U7969 (N_7969,N_7841,N_7878);
and U7970 (N_7970,N_7911,N_7824);
nand U7971 (N_7971,N_7945,N_7826);
and U7972 (N_7972,N_7918,N_7875);
and U7973 (N_7973,N_7896,N_7838);
and U7974 (N_7974,N_7908,N_7916);
nor U7975 (N_7975,N_7933,N_7884);
and U7976 (N_7976,N_7801,N_7931);
nand U7977 (N_7977,N_7849,N_7873);
or U7978 (N_7978,N_7819,N_7891);
nor U7979 (N_7979,N_7928,N_7870);
nand U7980 (N_7980,N_7836,N_7882);
nand U7981 (N_7981,N_7820,N_7944);
nor U7982 (N_7982,N_7851,N_7913);
nand U7983 (N_7983,N_7844,N_7830);
nand U7984 (N_7984,N_7897,N_7829);
nand U7985 (N_7985,N_7823,N_7847);
nor U7986 (N_7986,N_7900,N_7853);
nor U7987 (N_7987,N_7837,N_7877);
xnor U7988 (N_7988,N_7890,N_7817);
and U7989 (N_7989,N_7803,N_7858);
or U7990 (N_7990,N_7888,N_7926);
or U7991 (N_7991,N_7894,N_7807);
or U7992 (N_7992,N_7946,N_7949);
and U7993 (N_7993,N_7818,N_7852);
nor U7994 (N_7994,N_7917,N_7924);
and U7995 (N_7995,N_7814,N_7923);
or U7996 (N_7996,N_7833,N_7909);
xor U7997 (N_7997,N_7889,N_7937);
nor U7998 (N_7998,N_7860,N_7843);
nand U7999 (N_7999,N_7903,N_7922);
or U8000 (N_8000,N_7809,N_7802);
nand U8001 (N_8001,N_7880,N_7831);
nor U8002 (N_8002,N_7834,N_7854);
nor U8003 (N_8003,N_7940,N_7832);
nor U8004 (N_8004,N_7871,N_7815);
or U8005 (N_8005,N_7821,N_7800);
nand U8006 (N_8006,N_7939,N_7906);
nor U8007 (N_8007,N_7904,N_7892);
nor U8008 (N_8008,N_7813,N_7898);
nand U8009 (N_8009,N_7899,N_7868);
nor U8010 (N_8010,N_7835,N_7812);
nand U8011 (N_8011,N_7808,N_7816);
and U8012 (N_8012,N_7919,N_7822);
nand U8013 (N_8013,N_7886,N_7905);
and U8014 (N_8014,N_7845,N_7855);
and U8015 (N_8015,N_7893,N_7887);
and U8016 (N_8016,N_7935,N_7805);
nor U8017 (N_8017,N_7883,N_7839);
nand U8018 (N_8018,N_7862,N_7867);
or U8019 (N_8019,N_7850,N_7942);
nand U8020 (N_8020,N_7947,N_7915);
or U8021 (N_8021,N_7810,N_7929);
or U8022 (N_8022,N_7840,N_7921);
and U8023 (N_8023,N_7876,N_7895);
and U8024 (N_8024,N_7848,N_7865);
nand U8025 (N_8025,N_7901,N_7800);
xor U8026 (N_8026,N_7885,N_7838);
nand U8027 (N_8027,N_7836,N_7896);
and U8028 (N_8028,N_7885,N_7897);
nand U8029 (N_8029,N_7802,N_7849);
nor U8030 (N_8030,N_7885,N_7917);
xor U8031 (N_8031,N_7805,N_7899);
or U8032 (N_8032,N_7919,N_7914);
or U8033 (N_8033,N_7942,N_7907);
and U8034 (N_8034,N_7853,N_7831);
nand U8035 (N_8035,N_7904,N_7936);
and U8036 (N_8036,N_7909,N_7920);
nor U8037 (N_8037,N_7934,N_7821);
nor U8038 (N_8038,N_7937,N_7941);
xnor U8039 (N_8039,N_7812,N_7806);
nor U8040 (N_8040,N_7858,N_7850);
nand U8041 (N_8041,N_7845,N_7899);
or U8042 (N_8042,N_7900,N_7909);
or U8043 (N_8043,N_7905,N_7917);
nor U8044 (N_8044,N_7914,N_7826);
and U8045 (N_8045,N_7808,N_7802);
nand U8046 (N_8046,N_7904,N_7813);
or U8047 (N_8047,N_7862,N_7869);
nand U8048 (N_8048,N_7893,N_7827);
nand U8049 (N_8049,N_7827,N_7850);
nand U8050 (N_8050,N_7825,N_7897);
and U8051 (N_8051,N_7822,N_7846);
or U8052 (N_8052,N_7925,N_7827);
nor U8053 (N_8053,N_7948,N_7823);
nor U8054 (N_8054,N_7922,N_7877);
and U8055 (N_8055,N_7934,N_7908);
nor U8056 (N_8056,N_7932,N_7846);
and U8057 (N_8057,N_7843,N_7866);
and U8058 (N_8058,N_7908,N_7910);
nor U8059 (N_8059,N_7861,N_7912);
and U8060 (N_8060,N_7807,N_7805);
nor U8061 (N_8061,N_7849,N_7915);
nand U8062 (N_8062,N_7860,N_7887);
xor U8063 (N_8063,N_7854,N_7879);
xnor U8064 (N_8064,N_7939,N_7924);
and U8065 (N_8065,N_7897,N_7808);
and U8066 (N_8066,N_7800,N_7917);
and U8067 (N_8067,N_7870,N_7824);
and U8068 (N_8068,N_7833,N_7832);
or U8069 (N_8069,N_7885,N_7870);
nor U8070 (N_8070,N_7936,N_7853);
and U8071 (N_8071,N_7842,N_7841);
nor U8072 (N_8072,N_7937,N_7857);
nand U8073 (N_8073,N_7944,N_7804);
and U8074 (N_8074,N_7898,N_7870);
and U8075 (N_8075,N_7907,N_7823);
and U8076 (N_8076,N_7806,N_7824);
nor U8077 (N_8077,N_7929,N_7864);
or U8078 (N_8078,N_7875,N_7898);
or U8079 (N_8079,N_7901,N_7894);
nand U8080 (N_8080,N_7874,N_7826);
or U8081 (N_8081,N_7820,N_7867);
and U8082 (N_8082,N_7941,N_7915);
or U8083 (N_8083,N_7807,N_7914);
and U8084 (N_8084,N_7910,N_7876);
nand U8085 (N_8085,N_7923,N_7844);
nand U8086 (N_8086,N_7844,N_7814);
or U8087 (N_8087,N_7840,N_7907);
nand U8088 (N_8088,N_7909,N_7843);
nor U8089 (N_8089,N_7936,N_7935);
xnor U8090 (N_8090,N_7925,N_7891);
xnor U8091 (N_8091,N_7901,N_7933);
nand U8092 (N_8092,N_7868,N_7919);
and U8093 (N_8093,N_7808,N_7852);
and U8094 (N_8094,N_7924,N_7821);
nand U8095 (N_8095,N_7843,N_7918);
and U8096 (N_8096,N_7933,N_7827);
and U8097 (N_8097,N_7949,N_7893);
nand U8098 (N_8098,N_7849,N_7913);
and U8099 (N_8099,N_7884,N_7813);
nand U8100 (N_8100,N_7963,N_8063);
nor U8101 (N_8101,N_7956,N_8023);
and U8102 (N_8102,N_7962,N_7973);
or U8103 (N_8103,N_7978,N_7992);
xnor U8104 (N_8104,N_8071,N_8084);
and U8105 (N_8105,N_8083,N_8027);
and U8106 (N_8106,N_7970,N_8093);
nand U8107 (N_8107,N_8098,N_8020);
and U8108 (N_8108,N_7960,N_7997);
or U8109 (N_8109,N_8058,N_8059);
and U8110 (N_8110,N_8051,N_8034);
or U8111 (N_8111,N_8017,N_7990);
nor U8112 (N_8112,N_7974,N_8039);
nand U8113 (N_8113,N_8054,N_8086);
xnor U8114 (N_8114,N_8036,N_8013);
or U8115 (N_8115,N_8021,N_8041);
and U8116 (N_8116,N_7981,N_8052);
xnor U8117 (N_8117,N_8061,N_7955);
xor U8118 (N_8118,N_8008,N_8022);
nor U8119 (N_8119,N_8043,N_8009);
nor U8120 (N_8120,N_8040,N_8010);
nor U8121 (N_8121,N_8028,N_8003);
and U8122 (N_8122,N_8062,N_8006);
and U8123 (N_8123,N_7994,N_8065);
nand U8124 (N_8124,N_7989,N_8091);
nand U8125 (N_8125,N_8056,N_8085);
or U8126 (N_8126,N_8069,N_8001);
nor U8127 (N_8127,N_8089,N_8088);
or U8128 (N_8128,N_8060,N_8070);
nor U8129 (N_8129,N_7988,N_7976);
nand U8130 (N_8130,N_8005,N_8057);
nand U8131 (N_8131,N_7985,N_8090);
nand U8132 (N_8132,N_8031,N_7959);
nor U8133 (N_8133,N_7980,N_7995);
or U8134 (N_8134,N_8004,N_7983);
or U8135 (N_8135,N_8045,N_7952);
or U8136 (N_8136,N_7954,N_7991);
nor U8137 (N_8137,N_7971,N_7975);
or U8138 (N_8138,N_7986,N_7999);
and U8139 (N_8139,N_8068,N_8077);
or U8140 (N_8140,N_7961,N_8015);
or U8141 (N_8141,N_7958,N_8047);
or U8142 (N_8142,N_7977,N_7979);
nand U8143 (N_8143,N_8035,N_8032);
xor U8144 (N_8144,N_8019,N_8064);
nor U8145 (N_8145,N_8029,N_8030);
or U8146 (N_8146,N_7993,N_8096);
and U8147 (N_8147,N_8072,N_8055);
nor U8148 (N_8148,N_7965,N_8038);
nor U8149 (N_8149,N_7984,N_7957);
nor U8150 (N_8150,N_8067,N_8037);
xnor U8151 (N_8151,N_8026,N_8079);
and U8152 (N_8152,N_8014,N_8073);
or U8153 (N_8153,N_8007,N_8053);
nand U8154 (N_8154,N_8012,N_7972);
nor U8155 (N_8155,N_8076,N_8092);
nand U8156 (N_8156,N_8042,N_8066);
or U8157 (N_8157,N_7967,N_8002);
and U8158 (N_8158,N_8099,N_8049);
and U8159 (N_8159,N_7996,N_7968);
nand U8160 (N_8160,N_8078,N_8025);
nor U8161 (N_8161,N_8080,N_7987);
and U8162 (N_8162,N_8050,N_8095);
and U8163 (N_8163,N_8018,N_7982);
nand U8164 (N_8164,N_7969,N_8097);
or U8165 (N_8165,N_8074,N_7998);
nor U8166 (N_8166,N_8011,N_8000);
nor U8167 (N_8167,N_8016,N_7951);
nand U8168 (N_8168,N_8087,N_7966);
nand U8169 (N_8169,N_8081,N_7950);
or U8170 (N_8170,N_8048,N_7964);
or U8171 (N_8171,N_8046,N_8033);
or U8172 (N_8172,N_8082,N_8024);
xnor U8173 (N_8173,N_7953,N_8075);
or U8174 (N_8174,N_8094,N_8044);
or U8175 (N_8175,N_8007,N_7958);
and U8176 (N_8176,N_8021,N_7983);
nor U8177 (N_8177,N_8067,N_7962);
nand U8178 (N_8178,N_8007,N_7969);
nor U8179 (N_8179,N_7961,N_7985);
or U8180 (N_8180,N_7978,N_7998);
nand U8181 (N_8181,N_7960,N_7973);
nor U8182 (N_8182,N_8016,N_8097);
xnor U8183 (N_8183,N_7954,N_8013);
nor U8184 (N_8184,N_8035,N_8003);
nand U8185 (N_8185,N_7993,N_8027);
or U8186 (N_8186,N_7996,N_8022);
or U8187 (N_8187,N_8058,N_8070);
and U8188 (N_8188,N_7971,N_8026);
nor U8189 (N_8189,N_8065,N_8078);
or U8190 (N_8190,N_7970,N_8095);
and U8191 (N_8191,N_7989,N_8046);
nand U8192 (N_8192,N_8066,N_8040);
nor U8193 (N_8193,N_7984,N_8050);
nor U8194 (N_8194,N_8057,N_8098);
or U8195 (N_8195,N_8036,N_8057);
nor U8196 (N_8196,N_7978,N_7986);
and U8197 (N_8197,N_7982,N_8046);
nor U8198 (N_8198,N_7961,N_8004);
nor U8199 (N_8199,N_8056,N_8000);
nor U8200 (N_8200,N_8070,N_8037);
nor U8201 (N_8201,N_7958,N_8067);
or U8202 (N_8202,N_8033,N_8047);
nor U8203 (N_8203,N_7972,N_8008);
nor U8204 (N_8204,N_8027,N_8008);
nand U8205 (N_8205,N_8099,N_8033);
nand U8206 (N_8206,N_8076,N_7990);
nor U8207 (N_8207,N_8082,N_8019);
nor U8208 (N_8208,N_7974,N_8052);
xnor U8209 (N_8209,N_8027,N_8043);
nor U8210 (N_8210,N_8079,N_8074);
nor U8211 (N_8211,N_8074,N_8054);
xor U8212 (N_8212,N_8084,N_7995);
nor U8213 (N_8213,N_8011,N_8012);
nor U8214 (N_8214,N_8077,N_8017);
or U8215 (N_8215,N_7988,N_8039);
xnor U8216 (N_8216,N_8075,N_7976);
nand U8217 (N_8217,N_7984,N_7988);
or U8218 (N_8218,N_8067,N_7984);
nor U8219 (N_8219,N_8089,N_7966);
or U8220 (N_8220,N_7987,N_8062);
nor U8221 (N_8221,N_8030,N_8048);
or U8222 (N_8222,N_8036,N_7984);
and U8223 (N_8223,N_7990,N_8044);
xnor U8224 (N_8224,N_8093,N_7972);
nand U8225 (N_8225,N_7996,N_8055);
nand U8226 (N_8226,N_7980,N_8028);
nand U8227 (N_8227,N_8018,N_8070);
nor U8228 (N_8228,N_8084,N_8022);
and U8229 (N_8229,N_8099,N_8042);
nor U8230 (N_8230,N_7980,N_8083);
nand U8231 (N_8231,N_8065,N_8019);
and U8232 (N_8232,N_8040,N_8076);
nor U8233 (N_8233,N_8018,N_7987);
and U8234 (N_8234,N_7979,N_8031);
nor U8235 (N_8235,N_7976,N_7959);
and U8236 (N_8236,N_8029,N_8051);
or U8237 (N_8237,N_8084,N_8046);
nor U8238 (N_8238,N_7969,N_7963);
nor U8239 (N_8239,N_7986,N_8044);
nand U8240 (N_8240,N_7985,N_7988);
xor U8241 (N_8241,N_8053,N_8015);
and U8242 (N_8242,N_8053,N_7967);
or U8243 (N_8243,N_8030,N_8065);
or U8244 (N_8244,N_8033,N_8045);
xor U8245 (N_8245,N_7995,N_8013);
or U8246 (N_8246,N_7995,N_7989);
or U8247 (N_8247,N_8082,N_7990);
xnor U8248 (N_8248,N_7956,N_8099);
nor U8249 (N_8249,N_7981,N_8087);
nand U8250 (N_8250,N_8117,N_8156);
xor U8251 (N_8251,N_8118,N_8146);
nor U8252 (N_8252,N_8245,N_8216);
and U8253 (N_8253,N_8176,N_8236);
nor U8254 (N_8254,N_8215,N_8208);
nor U8255 (N_8255,N_8140,N_8186);
and U8256 (N_8256,N_8242,N_8172);
nor U8257 (N_8257,N_8243,N_8100);
xor U8258 (N_8258,N_8161,N_8130);
xnor U8259 (N_8259,N_8137,N_8197);
and U8260 (N_8260,N_8225,N_8180);
or U8261 (N_8261,N_8145,N_8141);
or U8262 (N_8262,N_8151,N_8183);
xnor U8263 (N_8263,N_8219,N_8115);
or U8264 (N_8264,N_8101,N_8241);
nand U8265 (N_8265,N_8139,N_8160);
and U8266 (N_8266,N_8154,N_8249);
and U8267 (N_8267,N_8207,N_8111);
and U8268 (N_8268,N_8202,N_8175);
or U8269 (N_8269,N_8237,N_8187);
and U8270 (N_8270,N_8119,N_8201);
or U8271 (N_8271,N_8211,N_8158);
nor U8272 (N_8272,N_8195,N_8113);
nand U8273 (N_8273,N_8133,N_8179);
and U8274 (N_8274,N_8184,N_8230);
nor U8275 (N_8275,N_8238,N_8192);
nand U8276 (N_8276,N_8116,N_8205);
or U8277 (N_8277,N_8199,N_8165);
nor U8278 (N_8278,N_8200,N_8239);
and U8279 (N_8279,N_8226,N_8102);
nand U8280 (N_8280,N_8136,N_8214);
nor U8281 (N_8281,N_8108,N_8244);
and U8282 (N_8282,N_8203,N_8173);
nand U8283 (N_8283,N_8144,N_8220);
nand U8284 (N_8284,N_8232,N_8229);
nand U8285 (N_8285,N_8107,N_8122);
xnor U8286 (N_8286,N_8142,N_8174);
nor U8287 (N_8287,N_8128,N_8110);
nand U8288 (N_8288,N_8193,N_8114);
or U8289 (N_8289,N_8190,N_8228);
and U8290 (N_8290,N_8104,N_8170);
nand U8291 (N_8291,N_8152,N_8148);
or U8292 (N_8292,N_8134,N_8209);
nor U8293 (N_8293,N_8221,N_8204);
and U8294 (N_8294,N_8189,N_8248);
and U8295 (N_8295,N_8178,N_8135);
or U8296 (N_8296,N_8191,N_8149);
and U8297 (N_8297,N_8126,N_8233);
or U8298 (N_8298,N_8159,N_8227);
nand U8299 (N_8299,N_8121,N_8231);
and U8300 (N_8300,N_8109,N_8213);
nor U8301 (N_8301,N_8167,N_8123);
or U8302 (N_8302,N_8181,N_8166);
xor U8303 (N_8303,N_8235,N_8150);
nand U8304 (N_8304,N_8120,N_8105);
and U8305 (N_8305,N_8157,N_8171);
xnor U8306 (N_8306,N_8234,N_8196);
nor U8307 (N_8307,N_8132,N_8153);
xor U8308 (N_8308,N_8182,N_8106);
nor U8309 (N_8309,N_8131,N_8138);
nand U8310 (N_8310,N_8155,N_8223);
nand U8311 (N_8311,N_8188,N_8125);
or U8312 (N_8312,N_8162,N_8177);
and U8313 (N_8313,N_8217,N_8212);
nor U8314 (N_8314,N_8143,N_8222);
or U8315 (N_8315,N_8129,N_8124);
nand U8316 (N_8316,N_8147,N_8206);
nor U8317 (N_8317,N_8164,N_8224);
nor U8318 (N_8318,N_8168,N_8240);
nand U8319 (N_8319,N_8246,N_8198);
and U8320 (N_8320,N_8163,N_8103);
nand U8321 (N_8321,N_8127,N_8185);
nand U8322 (N_8322,N_8247,N_8194);
or U8323 (N_8323,N_8218,N_8210);
and U8324 (N_8324,N_8169,N_8112);
and U8325 (N_8325,N_8216,N_8243);
nor U8326 (N_8326,N_8228,N_8120);
nand U8327 (N_8327,N_8198,N_8108);
and U8328 (N_8328,N_8101,N_8152);
xor U8329 (N_8329,N_8201,N_8191);
or U8330 (N_8330,N_8212,N_8229);
nor U8331 (N_8331,N_8209,N_8240);
nor U8332 (N_8332,N_8175,N_8204);
nand U8333 (N_8333,N_8246,N_8170);
nand U8334 (N_8334,N_8114,N_8242);
nor U8335 (N_8335,N_8204,N_8121);
nor U8336 (N_8336,N_8142,N_8112);
nor U8337 (N_8337,N_8180,N_8138);
and U8338 (N_8338,N_8237,N_8146);
nor U8339 (N_8339,N_8183,N_8123);
or U8340 (N_8340,N_8206,N_8232);
and U8341 (N_8341,N_8200,N_8203);
nand U8342 (N_8342,N_8120,N_8217);
xnor U8343 (N_8343,N_8170,N_8159);
and U8344 (N_8344,N_8197,N_8173);
xnor U8345 (N_8345,N_8100,N_8187);
or U8346 (N_8346,N_8132,N_8129);
nor U8347 (N_8347,N_8132,N_8103);
and U8348 (N_8348,N_8104,N_8136);
or U8349 (N_8349,N_8246,N_8137);
nand U8350 (N_8350,N_8130,N_8182);
nand U8351 (N_8351,N_8122,N_8179);
nor U8352 (N_8352,N_8133,N_8218);
or U8353 (N_8353,N_8198,N_8209);
and U8354 (N_8354,N_8170,N_8102);
or U8355 (N_8355,N_8237,N_8148);
and U8356 (N_8356,N_8211,N_8136);
nor U8357 (N_8357,N_8136,N_8171);
and U8358 (N_8358,N_8235,N_8142);
nand U8359 (N_8359,N_8203,N_8216);
and U8360 (N_8360,N_8149,N_8171);
nand U8361 (N_8361,N_8240,N_8106);
or U8362 (N_8362,N_8142,N_8125);
nand U8363 (N_8363,N_8113,N_8118);
and U8364 (N_8364,N_8101,N_8157);
nand U8365 (N_8365,N_8213,N_8211);
and U8366 (N_8366,N_8117,N_8174);
nand U8367 (N_8367,N_8215,N_8132);
nand U8368 (N_8368,N_8124,N_8119);
or U8369 (N_8369,N_8114,N_8197);
xnor U8370 (N_8370,N_8167,N_8206);
and U8371 (N_8371,N_8236,N_8247);
or U8372 (N_8372,N_8218,N_8146);
nand U8373 (N_8373,N_8159,N_8173);
or U8374 (N_8374,N_8224,N_8128);
and U8375 (N_8375,N_8212,N_8152);
or U8376 (N_8376,N_8135,N_8159);
or U8377 (N_8377,N_8240,N_8222);
or U8378 (N_8378,N_8139,N_8198);
nand U8379 (N_8379,N_8219,N_8195);
and U8380 (N_8380,N_8134,N_8115);
nor U8381 (N_8381,N_8225,N_8175);
nor U8382 (N_8382,N_8162,N_8144);
and U8383 (N_8383,N_8147,N_8122);
or U8384 (N_8384,N_8133,N_8228);
nand U8385 (N_8385,N_8194,N_8231);
or U8386 (N_8386,N_8167,N_8218);
or U8387 (N_8387,N_8173,N_8132);
or U8388 (N_8388,N_8153,N_8140);
and U8389 (N_8389,N_8247,N_8171);
xnor U8390 (N_8390,N_8156,N_8249);
or U8391 (N_8391,N_8124,N_8208);
nand U8392 (N_8392,N_8248,N_8245);
or U8393 (N_8393,N_8195,N_8177);
or U8394 (N_8394,N_8156,N_8246);
nand U8395 (N_8395,N_8231,N_8232);
or U8396 (N_8396,N_8157,N_8190);
and U8397 (N_8397,N_8237,N_8215);
and U8398 (N_8398,N_8244,N_8169);
nor U8399 (N_8399,N_8168,N_8192);
xnor U8400 (N_8400,N_8299,N_8355);
xor U8401 (N_8401,N_8292,N_8290);
xor U8402 (N_8402,N_8351,N_8312);
and U8403 (N_8403,N_8372,N_8303);
nand U8404 (N_8404,N_8297,N_8311);
or U8405 (N_8405,N_8324,N_8395);
nor U8406 (N_8406,N_8268,N_8266);
xor U8407 (N_8407,N_8341,N_8285);
and U8408 (N_8408,N_8380,N_8274);
or U8409 (N_8409,N_8322,N_8252);
xnor U8410 (N_8410,N_8371,N_8353);
nor U8411 (N_8411,N_8314,N_8348);
nand U8412 (N_8412,N_8261,N_8317);
nor U8413 (N_8413,N_8326,N_8367);
nor U8414 (N_8414,N_8381,N_8366);
or U8415 (N_8415,N_8389,N_8387);
and U8416 (N_8416,N_8323,N_8272);
or U8417 (N_8417,N_8330,N_8345);
nand U8418 (N_8418,N_8358,N_8383);
and U8419 (N_8419,N_8321,N_8343);
nor U8420 (N_8420,N_8376,N_8319);
nand U8421 (N_8421,N_8393,N_8284);
nand U8422 (N_8422,N_8309,N_8397);
and U8423 (N_8423,N_8377,N_8291);
nand U8424 (N_8424,N_8255,N_8276);
or U8425 (N_8425,N_8265,N_8264);
nand U8426 (N_8426,N_8277,N_8335);
and U8427 (N_8427,N_8273,N_8289);
xnor U8428 (N_8428,N_8369,N_8315);
nand U8429 (N_8429,N_8281,N_8260);
or U8430 (N_8430,N_8263,N_8256);
nand U8431 (N_8431,N_8279,N_8270);
nand U8432 (N_8432,N_8275,N_8278);
and U8433 (N_8433,N_8384,N_8307);
nor U8434 (N_8434,N_8356,N_8357);
nor U8435 (N_8435,N_8251,N_8375);
nand U8436 (N_8436,N_8334,N_8313);
xor U8437 (N_8437,N_8385,N_8374);
nor U8438 (N_8438,N_8396,N_8294);
nor U8439 (N_8439,N_8368,N_8349);
and U8440 (N_8440,N_8286,N_8382);
nor U8441 (N_8441,N_8316,N_8362);
and U8442 (N_8442,N_8328,N_8300);
or U8443 (N_8443,N_8360,N_8388);
nor U8444 (N_8444,N_8331,N_8298);
and U8445 (N_8445,N_8399,N_8306);
or U8446 (N_8446,N_8390,N_8370);
or U8447 (N_8447,N_8386,N_8336);
nor U8448 (N_8448,N_8361,N_8259);
nand U8449 (N_8449,N_8347,N_8394);
nor U8450 (N_8450,N_8344,N_8359);
or U8451 (N_8451,N_8253,N_8379);
nand U8452 (N_8452,N_8391,N_8250);
nand U8453 (N_8453,N_8254,N_8282);
nand U8454 (N_8454,N_8304,N_8305);
or U8455 (N_8455,N_8337,N_8258);
nor U8456 (N_8456,N_8308,N_8378);
xor U8457 (N_8457,N_8364,N_8365);
nand U8458 (N_8458,N_8392,N_8296);
and U8459 (N_8459,N_8325,N_8267);
and U8460 (N_8460,N_8363,N_8302);
or U8461 (N_8461,N_8373,N_8333);
nand U8462 (N_8462,N_8293,N_8398);
nor U8463 (N_8463,N_8354,N_8310);
nor U8464 (N_8464,N_8332,N_8327);
or U8465 (N_8465,N_8346,N_8257);
nand U8466 (N_8466,N_8301,N_8342);
and U8467 (N_8467,N_8283,N_8338);
nand U8468 (N_8468,N_8339,N_8271);
xnor U8469 (N_8469,N_8340,N_8269);
or U8470 (N_8470,N_8288,N_8287);
and U8471 (N_8471,N_8318,N_8262);
xor U8472 (N_8472,N_8329,N_8295);
or U8473 (N_8473,N_8352,N_8280);
nand U8474 (N_8474,N_8320,N_8350);
nand U8475 (N_8475,N_8288,N_8276);
or U8476 (N_8476,N_8353,N_8389);
or U8477 (N_8477,N_8286,N_8354);
or U8478 (N_8478,N_8258,N_8347);
nand U8479 (N_8479,N_8309,N_8327);
and U8480 (N_8480,N_8361,N_8297);
nand U8481 (N_8481,N_8256,N_8283);
nand U8482 (N_8482,N_8359,N_8277);
nand U8483 (N_8483,N_8379,N_8340);
nor U8484 (N_8484,N_8327,N_8310);
nor U8485 (N_8485,N_8277,N_8383);
and U8486 (N_8486,N_8378,N_8318);
or U8487 (N_8487,N_8389,N_8319);
nor U8488 (N_8488,N_8251,N_8321);
nand U8489 (N_8489,N_8394,N_8305);
nand U8490 (N_8490,N_8377,N_8355);
nand U8491 (N_8491,N_8256,N_8251);
or U8492 (N_8492,N_8251,N_8276);
or U8493 (N_8493,N_8273,N_8320);
xnor U8494 (N_8494,N_8340,N_8258);
nand U8495 (N_8495,N_8271,N_8343);
or U8496 (N_8496,N_8320,N_8366);
nand U8497 (N_8497,N_8371,N_8263);
xnor U8498 (N_8498,N_8256,N_8250);
and U8499 (N_8499,N_8344,N_8317);
and U8500 (N_8500,N_8272,N_8280);
nand U8501 (N_8501,N_8330,N_8389);
and U8502 (N_8502,N_8364,N_8284);
or U8503 (N_8503,N_8352,N_8393);
and U8504 (N_8504,N_8342,N_8316);
nor U8505 (N_8505,N_8379,N_8322);
and U8506 (N_8506,N_8325,N_8315);
nand U8507 (N_8507,N_8323,N_8363);
or U8508 (N_8508,N_8323,N_8290);
or U8509 (N_8509,N_8326,N_8344);
nand U8510 (N_8510,N_8388,N_8274);
or U8511 (N_8511,N_8390,N_8316);
nand U8512 (N_8512,N_8314,N_8317);
xor U8513 (N_8513,N_8309,N_8359);
nor U8514 (N_8514,N_8396,N_8300);
and U8515 (N_8515,N_8288,N_8395);
nor U8516 (N_8516,N_8373,N_8331);
nor U8517 (N_8517,N_8364,N_8263);
nand U8518 (N_8518,N_8297,N_8257);
nor U8519 (N_8519,N_8393,N_8390);
and U8520 (N_8520,N_8367,N_8360);
xnor U8521 (N_8521,N_8347,N_8385);
and U8522 (N_8522,N_8395,N_8388);
and U8523 (N_8523,N_8359,N_8386);
nand U8524 (N_8524,N_8284,N_8375);
or U8525 (N_8525,N_8382,N_8295);
and U8526 (N_8526,N_8309,N_8332);
and U8527 (N_8527,N_8254,N_8318);
or U8528 (N_8528,N_8288,N_8282);
nand U8529 (N_8529,N_8289,N_8274);
or U8530 (N_8530,N_8372,N_8342);
and U8531 (N_8531,N_8340,N_8319);
nor U8532 (N_8532,N_8366,N_8279);
and U8533 (N_8533,N_8340,N_8327);
nand U8534 (N_8534,N_8362,N_8274);
or U8535 (N_8535,N_8336,N_8269);
nand U8536 (N_8536,N_8352,N_8365);
xor U8537 (N_8537,N_8337,N_8299);
nor U8538 (N_8538,N_8307,N_8398);
or U8539 (N_8539,N_8352,N_8270);
nor U8540 (N_8540,N_8289,N_8373);
xor U8541 (N_8541,N_8320,N_8267);
or U8542 (N_8542,N_8291,N_8268);
and U8543 (N_8543,N_8326,N_8280);
and U8544 (N_8544,N_8307,N_8279);
nand U8545 (N_8545,N_8263,N_8319);
and U8546 (N_8546,N_8346,N_8377);
and U8547 (N_8547,N_8341,N_8347);
nand U8548 (N_8548,N_8392,N_8281);
xor U8549 (N_8549,N_8394,N_8363);
nand U8550 (N_8550,N_8403,N_8473);
nand U8551 (N_8551,N_8540,N_8538);
and U8552 (N_8552,N_8543,N_8524);
xnor U8553 (N_8553,N_8466,N_8430);
nor U8554 (N_8554,N_8418,N_8433);
nand U8555 (N_8555,N_8472,N_8449);
and U8556 (N_8556,N_8499,N_8451);
xnor U8557 (N_8557,N_8535,N_8479);
and U8558 (N_8558,N_8445,N_8456);
xnor U8559 (N_8559,N_8471,N_8431);
xnor U8560 (N_8560,N_8469,N_8467);
nand U8561 (N_8561,N_8542,N_8498);
and U8562 (N_8562,N_8548,N_8484);
nand U8563 (N_8563,N_8470,N_8486);
and U8564 (N_8564,N_8432,N_8526);
and U8565 (N_8565,N_8491,N_8455);
and U8566 (N_8566,N_8406,N_8485);
nor U8567 (N_8567,N_8539,N_8423);
or U8568 (N_8568,N_8483,N_8530);
nand U8569 (N_8569,N_8411,N_8501);
xnor U8570 (N_8570,N_8459,N_8454);
nor U8571 (N_8571,N_8494,N_8520);
and U8572 (N_8572,N_8544,N_8518);
or U8573 (N_8573,N_8502,N_8489);
nand U8574 (N_8574,N_8514,N_8441);
and U8575 (N_8575,N_8528,N_8422);
xor U8576 (N_8576,N_8434,N_8405);
and U8577 (N_8577,N_8493,N_8437);
nor U8578 (N_8578,N_8508,N_8428);
nor U8579 (N_8579,N_8517,N_8410);
nor U8580 (N_8580,N_8481,N_8447);
xnor U8581 (N_8581,N_8438,N_8497);
and U8582 (N_8582,N_8490,N_8513);
nor U8583 (N_8583,N_8549,N_8420);
and U8584 (N_8584,N_8435,N_8407);
xor U8585 (N_8585,N_8427,N_8529);
or U8586 (N_8586,N_8426,N_8478);
and U8587 (N_8587,N_8442,N_8419);
xnor U8588 (N_8588,N_8461,N_8468);
or U8589 (N_8589,N_8452,N_8408);
and U8590 (N_8590,N_8487,N_8401);
nand U8591 (N_8591,N_8511,N_8450);
nor U8592 (N_8592,N_8474,N_8504);
and U8593 (N_8593,N_8523,N_8547);
nor U8594 (N_8594,N_8536,N_8436);
or U8595 (N_8595,N_8400,N_8477);
and U8596 (N_8596,N_8532,N_8534);
nor U8597 (N_8597,N_8492,N_8475);
or U8598 (N_8598,N_8421,N_8525);
and U8599 (N_8599,N_8521,N_8424);
xor U8600 (N_8600,N_8402,N_8488);
nand U8601 (N_8601,N_8537,N_8509);
nor U8602 (N_8602,N_8506,N_8500);
nor U8603 (N_8603,N_8516,N_8414);
or U8604 (N_8604,N_8448,N_8429);
and U8605 (N_8605,N_8503,N_8546);
xnor U8606 (N_8606,N_8413,N_8412);
nand U8607 (N_8607,N_8482,N_8443);
or U8608 (N_8608,N_8495,N_8496);
nand U8609 (N_8609,N_8505,N_8440);
and U8610 (N_8610,N_8507,N_8439);
nand U8611 (N_8611,N_8458,N_8545);
nand U8612 (N_8612,N_8417,N_8404);
and U8613 (N_8613,N_8444,N_8533);
nand U8614 (N_8614,N_8510,N_8465);
nand U8615 (N_8615,N_8457,N_8409);
xnor U8616 (N_8616,N_8515,N_8522);
or U8617 (N_8617,N_8460,N_8480);
and U8618 (N_8618,N_8446,N_8464);
xor U8619 (N_8619,N_8541,N_8463);
or U8620 (N_8620,N_8453,N_8415);
nor U8621 (N_8621,N_8527,N_8416);
nand U8622 (N_8622,N_8519,N_8512);
or U8623 (N_8623,N_8531,N_8462);
nand U8624 (N_8624,N_8476,N_8425);
nand U8625 (N_8625,N_8428,N_8515);
nand U8626 (N_8626,N_8423,N_8497);
nand U8627 (N_8627,N_8482,N_8534);
nand U8628 (N_8628,N_8483,N_8411);
or U8629 (N_8629,N_8478,N_8441);
nor U8630 (N_8630,N_8450,N_8423);
or U8631 (N_8631,N_8516,N_8437);
nand U8632 (N_8632,N_8401,N_8433);
or U8633 (N_8633,N_8508,N_8461);
nand U8634 (N_8634,N_8404,N_8548);
or U8635 (N_8635,N_8486,N_8422);
nor U8636 (N_8636,N_8457,N_8474);
and U8637 (N_8637,N_8451,N_8456);
or U8638 (N_8638,N_8444,N_8489);
nand U8639 (N_8639,N_8530,N_8527);
xnor U8640 (N_8640,N_8522,N_8544);
and U8641 (N_8641,N_8455,N_8525);
or U8642 (N_8642,N_8430,N_8424);
and U8643 (N_8643,N_8403,N_8412);
and U8644 (N_8644,N_8537,N_8542);
nand U8645 (N_8645,N_8547,N_8500);
nor U8646 (N_8646,N_8463,N_8506);
nor U8647 (N_8647,N_8538,N_8470);
nor U8648 (N_8648,N_8503,N_8411);
nor U8649 (N_8649,N_8405,N_8461);
or U8650 (N_8650,N_8533,N_8405);
nor U8651 (N_8651,N_8490,N_8408);
nor U8652 (N_8652,N_8453,N_8401);
nor U8653 (N_8653,N_8504,N_8518);
and U8654 (N_8654,N_8440,N_8489);
nor U8655 (N_8655,N_8448,N_8490);
nor U8656 (N_8656,N_8408,N_8549);
or U8657 (N_8657,N_8496,N_8440);
nor U8658 (N_8658,N_8477,N_8416);
xnor U8659 (N_8659,N_8460,N_8496);
nor U8660 (N_8660,N_8424,N_8509);
nor U8661 (N_8661,N_8521,N_8466);
nor U8662 (N_8662,N_8458,N_8449);
xor U8663 (N_8663,N_8470,N_8518);
nand U8664 (N_8664,N_8481,N_8503);
and U8665 (N_8665,N_8503,N_8500);
xnor U8666 (N_8666,N_8454,N_8464);
xor U8667 (N_8667,N_8441,N_8459);
nand U8668 (N_8668,N_8484,N_8421);
and U8669 (N_8669,N_8490,N_8512);
or U8670 (N_8670,N_8533,N_8478);
nand U8671 (N_8671,N_8426,N_8548);
nand U8672 (N_8672,N_8472,N_8505);
and U8673 (N_8673,N_8531,N_8473);
and U8674 (N_8674,N_8428,N_8402);
or U8675 (N_8675,N_8458,N_8453);
nor U8676 (N_8676,N_8548,N_8517);
nand U8677 (N_8677,N_8526,N_8465);
nor U8678 (N_8678,N_8453,N_8462);
and U8679 (N_8679,N_8427,N_8468);
nor U8680 (N_8680,N_8537,N_8508);
nor U8681 (N_8681,N_8424,N_8545);
nand U8682 (N_8682,N_8455,N_8450);
nand U8683 (N_8683,N_8421,N_8501);
and U8684 (N_8684,N_8540,N_8452);
nand U8685 (N_8685,N_8400,N_8401);
or U8686 (N_8686,N_8443,N_8547);
xnor U8687 (N_8687,N_8473,N_8422);
xnor U8688 (N_8688,N_8543,N_8505);
xnor U8689 (N_8689,N_8500,N_8499);
nand U8690 (N_8690,N_8504,N_8400);
and U8691 (N_8691,N_8450,N_8477);
or U8692 (N_8692,N_8414,N_8405);
nand U8693 (N_8693,N_8483,N_8456);
nor U8694 (N_8694,N_8427,N_8460);
or U8695 (N_8695,N_8546,N_8438);
nand U8696 (N_8696,N_8539,N_8427);
nor U8697 (N_8697,N_8527,N_8487);
nand U8698 (N_8698,N_8444,N_8432);
nor U8699 (N_8699,N_8527,N_8444);
nand U8700 (N_8700,N_8682,N_8579);
and U8701 (N_8701,N_8630,N_8645);
nand U8702 (N_8702,N_8672,N_8675);
nor U8703 (N_8703,N_8612,N_8596);
and U8704 (N_8704,N_8673,N_8623);
nand U8705 (N_8705,N_8565,N_8697);
nand U8706 (N_8706,N_8636,N_8571);
nand U8707 (N_8707,N_8691,N_8597);
nand U8708 (N_8708,N_8678,N_8559);
nor U8709 (N_8709,N_8670,N_8688);
or U8710 (N_8710,N_8555,N_8616);
nor U8711 (N_8711,N_8568,N_8581);
and U8712 (N_8712,N_8607,N_8569);
nand U8713 (N_8713,N_8633,N_8677);
nor U8714 (N_8714,N_8628,N_8694);
or U8715 (N_8715,N_8606,N_8564);
xnor U8716 (N_8716,N_8615,N_8562);
nand U8717 (N_8717,N_8580,N_8600);
nor U8718 (N_8718,N_8622,N_8593);
nand U8719 (N_8719,N_8576,N_8660);
nand U8720 (N_8720,N_8632,N_8595);
nor U8721 (N_8721,N_8646,N_8676);
or U8722 (N_8722,N_8649,N_8611);
nor U8723 (N_8723,N_8659,N_8619);
nand U8724 (N_8724,N_8693,N_8683);
and U8725 (N_8725,N_8613,N_8661);
nand U8726 (N_8726,N_8641,N_8586);
nand U8727 (N_8727,N_8644,N_8666);
nand U8728 (N_8728,N_8686,N_8639);
xnor U8729 (N_8729,N_8598,N_8654);
nand U8730 (N_8730,N_8668,N_8658);
nor U8731 (N_8731,N_8618,N_8674);
xor U8732 (N_8732,N_8588,N_8621);
and U8733 (N_8733,N_8584,N_8591);
and U8734 (N_8734,N_8601,N_8604);
nand U8735 (N_8735,N_8640,N_8656);
nor U8736 (N_8736,N_8599,N_8557);
nor U8737 (N_8737,N_8587,N_8589);
and U8738 (N_8738,N_8642,N_8651);
or U8739 (N_8739,N_8637,N_8608);
or U8740 (N_8740,N_8560,N_8681);
nor U8741 (N_8741,N_8647,N_8617);
nand U8742 (N_8742,N_8665,N_8610);
or U8743 (N_8743,N_8627,N_8638);
nor U8744 (N_8744,N_8648,N_8698);
and U8745 (N_8745,N_8662,N_8634);
xor U8746 (N_8746,N_8561,N_8663);
xor U8747 (N_8747,N_8554,N_8566);
nor U8748 (N_8748,N_8650,N_8563);
nand U8749 (N_8749,N_8655,N_8551);
or U8750 (N_8750,N_8590,N_8679);
nand U8751 (N_8751,N_8585,N_8609);
nand U8752 (N_8752,N_8553,N_8696);
nor U8753 (N_8753,N_8687,N_8690);
nor U8754 (N_8754,N_8652,N_8653);
and U8755 (N_8755,N_8552,N_8669);
nor U8756 (N_8756,N_8620,N_8624);
nor U8757 (N_8757,N_8684,N_8570);
nor U8758 (N_8758,N_8578,N_8657);
and U8759 (N_8759,N_8680,N_8574);
or U8760 (N_8760,N_8577,N_8699);
nand U8761 (N_8761,N_8592,N_8695);
xnor U8762 (N_8762,N_8556,N_8629);
nand U8763 (N_8763,N_8667,N_8692);
or U8764 (N_8764,N_8685,N_8643);
nand U8765 (N_8765,N_8625,N_8550);
and U8766 (N_8766,N_8664,N_8583);
xor U8767 (N_8767,N_8689,N_8603);
nand U8768 (N_8768,N_8635,N_8573);
or U8769 (N_8769,N_8582,N_8602);
and U8770 (N_8770,N_8567,N_8626);
xor U8771 (N_8771,N_8572,N_8671);
nand U8772 (N_8772,N_8594,N_8575);
nor U8773 (N_8773,N_8558,N_8614);
or U8774 (N_8774,N_8631,N_8605);
nand U8775 (N_8775,N_8628,N_8657);
and U8776 (N_8776,N_8687,N_8617);
nor U8777 (N_8777,N_8688,N_8572);
nor U8778 (N_8778,N_8647,N_8593);
or U8779 (N_8779,N_8692,N_8602);
nand U8780 (N_8780,N_8619,N_8594);
or U8781 (N_8781,N_8660,N_8674);
nand U8782 (N_8782,N_8600,N_8650);
nor U8783 (N_8783,N_8630,N_8602);
and U8784 (N_8784,N_8694,N_8560);
and U8785 (N_8785,N_8644,N_8684);
and U8786 (N_8786,N_8589,N_8606);
and U8787 (N_8787,N_8646,N_8585);
or U8788 (N_8788,N_8652,N_8691);
nand U8789 (N_8789,N_8595,N_8671);
and U8790 (N_8790,N_8588,N_8638);
nor U8791 (N_8791,N_8607,N_8683);
nor U8792 (N_8792,N_8585,N_8698);
xor U8793 (N_8793,N_8612,N_8690);
or U8794 (N_8794,N_8629,N_8604);
nand U8795 (N_8795,N_8663,N_8682);
or U8796 (N_8796,N_8644,N_8583);
nand U8797 (N_8797,N_8640,N_8555);
and U8798 (N_8798,N_8662,N_8659);
xnor U8799 (N_8799,N_8606,N_8649);
nor U8800 (N_8800,N_8616,N_8658);
nor U8801 (N_8801,N_8683,N_8670);
or U8802 (N_8802,N_8630,N_8665);
nor U8803 (N_8803,N_8609,N_8698);
nand U8804 (N_8804,N_8688,N_8618);
and U8805 (N_8805,N_8640,N_8631);
or U8806 (N_8806,N_8576,N_8629);
nor U8807 (N_8807,N_8628,N_8598);
and U8808 (N_8808,N_8636,N_8606);
or U8809 (N_8809,N_8681,N_8608);
nand U8810 (N_8810,N_8694,N_8678);
and U8811 (N_8811,N_8582,N_8578);
xnor U8812 (N_8812,N_8581,N_8579);
and U8813 (N_8813,N_8686,N_8633);
xnor U8814 (N_8814,N_8565,N_8609);
nor U8815 (N_8815,N_8642,N_8574);
and U8816 (N_8816,N_8673,N_8646);
and U8817 (N_8817,N_8582,N_8569);
nand U8818 (N_8818,N_8621,N_8635);
xnor U8819 (N_8819,N_8680,N_8634);
nor U8820 (N_8820,N_8621,N_8601);
or U8821 (N_8821,N_8672,N_8581);
and U8822 (N_8822,N_8578,N_8598);
and U8823 (N_8823,N_8677,N_8609);
xnor U8824 (N_8824,N_8561,N_8583);
and U8825 (N_8825,N_8686,N_8614);
xnor U8826 (N_8826,N_8590,N_8683);
nor U8827 (N_8827,N_8623,N_8584);
xnor U8828 (N_8828,N_8684,N_8688);
nand U8829 (N_8829,N_8602,N_8670);
nor U8830 (N_8830,N_8698,N_8633);
nor U8831 (N_8831,N_8637,N_8696);
nor U8832 (N_8832,N_8617,N_8628);
nor U8833 (N_8833,N_8694,N_8625);
or U8834 (N_8834,N_8552,N_8628);
nand U8835 (N_8835,N_8623,N_8698);
and U8836 (N_8836,N_8653,N_8590);
xnor U8837 (N_8837,N_8696,N_8617);
or U8838 (N_8838,N_8637,N_8580);
and U8839 (N_8839,N_8560,N_8664);
nor U8840 (N_8840,N_8567,N_8583);
or U8841 (N_8841,N_8622,N_8591);
nor U8842 (N_8842,N_8629,N_8692);
nor U8843 (N_8843,N_8659,N_8641);
and U8844 (N_8844,N_8627,N_8677);
nor U8845 (N_8845,N_8580,N_8613);
nor U8846 (N_8846,N_8675,N_8556);
nand U8847 (N_8847,N_8621,N_8677);
nor U8848 (N_8848,N_8580,N_8681);
or U8849 (N_8849,N_8571,N_8649);
and U8850 (N_8850,N_8847,N_8773);
and U8851 (N_8851,N_8794,N_8823);
nand U8852 (N_8852,N_8796,N_8762);
nand U8853 (N_8853,N_8706,N_8791);
or U8854 (N_8854,N_8744,N_8714);
nor U8855 (N_8855,N_8782,N_8781);
and U8856 (N_8856,N_8788,N_8831);
nand U8857 (N_8857,N_8735,N_8798);
xnor U8858 (N_8858,N_8777,N_8721);
nor U8859 (N_8859,N_8793,N_8713);
nor U8860 (N_8860,N_8790,N_8720);
or U8861 (N_8861,N_8797,N_8843);
or U8862 (N_8862,N_8813,N_8822);
nand U8863 (N_8863,N_8748,N_8743);
nand U8864 (N_8864,N_8703,N_8745);
nand U8865 (N_8865,N_8760,N_8836);
nor U8866 (N_8866,N_8815,N_8811);
nor U8867 (N_8867,N_8828,N_8768);
or U8868 (N_8868,N_8758,N_8741);
or U8869 (N_8869,N_8842,N_8759);
and U8870 (N_8870,N_8752,N_8807);
nand U8871 (N_8871,N_8709,N_8824);
nand U8872 (N_8872,N_8835,N_8783);
and U8873 (N_8873,N_8812,N_8784);
or U8874 (N_8874,N_8785,N_8751);
and U8875 (N_8875,N_8818,N_8849);
nor U8876 (N_8876,N_8731,N_8810);
nand U8877 (N_8877,N_8846,N_8786);
or U8878 (N_8878,N_8816,N_8707);
xnor U8879 (N_8879,N_8734,N_8806);
and U8880 (N_8880,N_8738,N_8761);
and U8881 (N_8881,N_8700,N_8756);
or U8882 (N_8882,N_8800,N_8844);
nand U8883 (N_8883,N_8817,N_8841);
and U8884 (N_8884,N_8737,N_8730);
or U8885 (N_8885,N_8755,N_8802);
or U8886 (N_8886,N_8845,N_8727);
xnor U8887 (N_8887,N_8719,N_8770);
xor U8888 (N_8888,N_8827,N_8778);
nor U8889 (N_8889,N_8747,N_8723);
or U8890 (N_8890,N_8712,N_8772);
or U8891 (N_8891,N_8739,N_8771);
nor U8892 (N_8892,N_8711,N_8763);
nand U8893 (N_8893,N_8808,N_8725);
nand U8894 (N_8894,N_8839,N_8814);
and U8895 (N_8895,N_8710,N_8795);
or U8896 (N_8896,N_8767,N_8833);
and U8897 (N_8897,N_8722,N_8825);
or U8898 (N_8898,N_8774,N_8779);
nand U8899 (N_8899,N_8840,N_8780);
nand U8900 (N_8900,N_8740,N_8749);
nand U8901 (N_8901,N_8757,N_8819);
nor U8902 (N_8902,N_8742,N_8718);
or U8903 (N_8903,N_8848,N_8805);
or U8904 (N_8904,N_8787,N_8769);
xor U8905 (N_8905,N_8821,N_8732);
or U8906 (N_8906,N_8789,N_8724);
or U8907 (N_8907,N_8804,N_8766);
nor U8908 (N_8908,N_8820,N_8705);
nand U8909 (N_8909,N_8826,N_8708);
and U8910 (N_8910,N_8834,N_8799);
xor U8911 (N_8911,N_8717,N_8701);
and U8912 (N_8912,N_8803,N_8832);
xor U8913 (N_8913,N_8809,N_8829);
and U8914 (N_8914,N_8837,N_8776);
nand U8915 (N_8915,N_8753,N_8750);
nand U8916 (N_8916,N_8729,N_8792);
nand U8917 (N_8917,N_8801,N_8736);
nand U8918 (N_8918,N_8830,N_8702);
and U8919 (N_8919,N_8726,N_8746);
nor U8920 (N_8920,N_8838,N_8716);
nand U8921 (N_8921,N_8733,N_8728);
or U8922 (N_8922,N_8704,N_8764);
nor U8923 (N_8923,N_8715,N_8765);
nor U8924 (N_8924,N_8775,N_8754);
nor U8925 (N_8925,N_8723,N_8835);
and U8926 (N_8926,N_8839,N_8821);
and U8927 (N_8927,N_8757,N_8720);
and U8928 (N_8928,N_8785,N_8810);
or U8929 (N_8929,N_8736,N_8841);
xnor U8930 (N_8930,N_8760,N_8753);
or U8931 (N_8931,N_8719,N_8756);
and U8932 (N_8932,N_8728,N_8798);
xnor U8933 (N_8933,N_8833,N_8804);
nand U8934 (N_8934,N_8823,N_8722);
xor U8935 (N_8935,N_8745,N_8738);
nand U8936 (N_8936,N_8827,N_8837);
nor U8937 (N_8937,N_8838,N_8818);
nand U8938 (N_8938,N_8828,N_8844);
nand U8939 (N_8939,N_8824,N_8790);
nor U8940 (N_8940,N_8842,N_8848);
nand U8941 (N_8941,N_8808,N_8707);
nand U8942 (N_8942,N_8813,N_8829);
xor U8943 (N_8943,N_8705,N_8734);
nand U8944 (N_8944,N_8713,N_8740);
and U8945 (N_8945,N_8783,N_8834);
and U8946 (N_8946,N_8770,N_8705);
xor U8947 (N_8947,N_8761,N_8787);
nor U8948 (N_8948,N_8841,N_8719);
or U8949 (N_8949,N_8771,N_8735);
or U8950 (N_8950,N_8754,N_8830);
nor U8951 (N_8951,N_8777,N_8768);
nor U8952 (N_8952,N_8716,N_8821);
and U8953 (N_8953,N_8814,N_8801);
nor U8954 (N_8954,N_8733,N_8758);
xnor U8955 (N_8955,N_8793,N_8787);
xor U8956 (N_8956,N_8847,N_8749);
nor U8957 (N_8957,N_8719,N_8711);
and U8958 (N_8958,N_8755,N_8777);
nor U8959 (N_8959,N_8724,N_8823);
or U8960 (N_8960,N_8733,N_8770);
xor U8961 (N_8961,N_8786,N_8779);
nand U8962 (N_8962,N_8758,N_8754);
nor U8963 (N_8963,N_8760,N_8737);
or U8964 (N_8964,N_8736,N_8717);
and U8965 (N_8965,N_8708,N_8745);
nand U8966 (N_8966,N_8732,N_8700);
nor U8967 (N_8967,N_8707,N_8817);
nor U8968 (N_8968,N_8770,N_8759);
nand U8969 (N_8969,N_8739,N_8737);
nand U8970 (N_8970,N_8737,N_8703);
and U8971 (N_8971,N_8808,N_8823);
nor U8972 (N_8972,N_8800,N_8833);
nor U8973 (N_8973,N_8847,N_8754);
and U8974 (N_8974,N_8817,N_8804);
nor U8975 (N_8975,N_8751,N_8790);
nor U8976 (N_8976,N_8720,N_8784);
and U8977 (N_8977,N_8750,N_8824);
and U8978 (N_8978,N_8725,N_8775);
and U8979 (N_8979,N_8760,N_8703);
nor U8980 (N_8980,N_8748,N_8740);
nand U8981 (N_8981,N_8833,N_8742);
nand U8982 (N_8982,N_8713,N_8722);
or U8983 (N_8983,N_8705,N_8738);
or U8984 (N_8984,N_8709,N_8830);
or U8985 (N_8985,N_8787,N_8792);
or U8986 (N_8986,N_8746,N_8816);
nor U8987 (N_8987,N_8722,N_8807);
or U8988 (N_8988,N_8797,N_8754);
and U8989 (N_8989,N_8799,N_8705);
and U8990 (N_8990,N_8823,N_8840);
and U8991 (N_8991,N_8752,N_8792);
or U8992 (N_8992,N_8786,N_8801);
or U8993 (N_8993,N_8764,N_8808);
nor U8994 (N_8994,N_8830,N_8802);
xnor U8995 (N_8995,N_8727,N_8752);
and U8996 (N_8996,N_8711,N_8734);
or U8997 (N_8997,N_8777,N_8833);
or U8998 (N_8998,N_8836,N_8763);
nor U8999 (N_8999,N_8803,N_8814);
and U9000 (N_9000,N_8920,N_8867);
or U9001 (N_9001,N_8885,N_8868);
xor U9002 (N_9002,N_8929,N_8884);
and U9003 (N_9003,N_8992,N_8932);
and U9004 (N_9004,N_8981,N_8854);
and U9005 (N_9005,N_8900,N_8955);
nand U9006 (N_9006,N_8873,N_8876);
and U9007 (N_9007,N_8972,N_8958);
xor U9008 (N_9008,N_8921,N_8925);
nor U9009 (N_9009,N_8903,N_8959);
xor U9010 (N_9010,N_8957,N_8927);
or U9011 (N_9011,N_8943,N_8917);
or U9012 (N_9012,N_8857,N_8978);
nor U9013 (N_9013,N_8971,N_8906);
nor U9014 (N_9014,N_8891,N_8950);
nor U9015 (N_9015,N_8938,N_8961);
or U9016 (N_9016,N_8912,N_8985);
or U9017 (N_9017,N_8913,N_8926);
and U9018 (N_9018,N_8969,N_8936);
nor U9019 (N_9019,N_8948,N_8907);
and U9020 (N_9020,N_8987,N_8939);
nor U9021 (N_9021,N_8979,N_8928);
xnor U9022 (N_9022,N_8931,N_8949);
and U9023 (N_9023,N_8942,N_8964);
and U9024 (N_9024,N_8894,N_8881);
nand U9025 (N_9025,N_8887,N_8982);
and U9026 (N_9026,N_8967,N_8883);
nand U9027 (N_9027,N_8863,N_8880);
nand U9028 (N_9028,N_8851,N_8915);
and U9029 (N_9029,N_8855,N_8997);
nand U9030 (N_9030,N_8898,N_8897);
nor U9031 (N_9031,N_8899,N_8944);
or U9032 (N_9032,N_8966,N_8914);
or U9033 (N_9033,N_8890,N_8924);
nand U9034 (N_9034,N_8945,N_8869);
nand U9035 (N_9035,N_8962,N_8879);
or U9036 (N_9036,N_8896,N_8940);
or U9037 (N_9037,N_8856,N_8953);
and U9038 (N_9038,N_8989,N_8963);
xnor U9039 (N_9039,N_8882,N_8996);
and U9040 (N_9040,N_8888,N_8970);
and U9041 (N_9041,N_8911,N_8946);
or U9042 (N_9042,N_8999,N_8954);
nor U9043 (N_9043,N_8935,N_8923);
nor U9044 (N_9044,N_8877,N_8995);
or U9045 (N_9045,N_8951,N_8991);
nand U9046 (N_9046,N_8910,N_8878);
or U9047 (N_9047,N_8968,N_8889);
nand U9048 (N_9048,N_8886,N_8993);
and U9049 (N_9049,N_8861,N_8941);
nor U9050 (N_9050,N_8918,N_8866);
or U9051 (N_9051,N_8956,N_8901);
nand U9052 (N_9052,N_8975,N_8974);
nor U9053 (N_9053,N_8976,N_8947);
or U9054 (N_9054,N_8870,N_8908);
nand U9055 (N_9055,N_8984,N_8850);
nand U9056 (N_9056,N_8960,N_8922);
xor U9057 (N_9057,N_8986,N_8916);
or U9058 (N_9058,N_8934,N_8871);
or U9059 (N_9059,N_8980,N_8998);
xnor U9060 (N_9060,N_8858,N_8973);
xnor U9061 (N_9061,N_8933,N_8983);
or U9062 (N_9062,N_8990,N_8875);
xnor U9063 (N_9063,N_8977,N_8862);
nand U9064 (N_9064,N_8965,N_8994);
nand U9065 (N_9065,N_8919,N_8904);
nor U9066 (N_9066,N_8893,N_8860);
and U9067 (N_9067,N_8853,N_8865);
nand U9068 (N_9068,N_8902,N_8892);
or U9069 (N_9069,N_8874,N_8930);
and U9070 (N_9070,N_8905,N_8909);
and U9071 (N_9071,N_8895,N_8872);
xnor U9072 (N_9072,N_8859,N_8864);
nor U9073 (N_9073,N_8852,N_8988);
xnor U9074 (N_9074,N_8937,N_8952);
nor U9075 (N_9075,N_8877,N_8952);
nor U9076 (N_9076,N_8895,N_8859);
nor U9077 (N_9077,N_8916,N_8985);
nand U9078 (N_9078,N_8941,N_8945);
or U9079 (N_9079,N_8869,N_8886);
and U9080 (N_9080,N_8920,N_8887);
or U9081 (N_9081,N_8993,N_8882);
or U9082 (N_9082,N_8893,N_8972);
or U9083 (N_9083,N_8920,N_8902);
nor U9084 (N_9084,N_8989,N_8962);
nor U9085 (N_9085,N_8981,N_8867);
and U9086 (N_9086,N_8973,N_8866);
or U9087 (N_9087,N_8997,N_8897);
nor U9088 (N_9088,N_8905,N_8925);
nor U9089 (N_9089,N_8935,N_8967);
and U9090 (N_9090,N_8880,N_8956);
and U9091 (N_9091,N_8924,N_8897);
and U9092 (N_9092,N_8963,N_8868);
and U9093 (N_9093,N_8876,N_8866);
and U9094 (N_9094,N_8998,N_8911);
or U9095 (N_9095,N_8924,N_8915);
and U9096 (N_9096,N_8961,N_8977);
nand U9097 (N_9097,N_8952,N_8936);
or U9098 (N_9098,N_8897,N_8941);
and U9099 (N_9099,N_8999,N_8965);
nor U9100 (N_9100,N_8875,N_8873);
and U9101 (N_9101,N_8883,N_8878);
xor U9102 (N_9102,N_8926,N_8995);
nand U9103 (N_9103,N_8971,N_8991);
nand U9104 (N_9104,N_8909,N_8900);
nand U9105 (N_9105,N_8981,N_8851);
nand U9106 (N_9106,N_8992,N_8867);
nor U9107 (N_9107,N_8897,N_8998);
and U9108 (N_9108,N_8973,N_8983);
nor U9109 (N_9109,N_8989,N_8863);
or U9110 (N_9110,N_8921,N_8973);
nor U9111 (N_9111,N_8954,N_8976);
and U9112 (N_9112,N_8899,N_8953);
nand U9113 (N_9113,N_8961,N_8864);
and U9114 (N_9114,N_8996,N_8997);
nand U9115 (N_9115,N_8992,N_8956);
and U9116 (N_9116,N_8898,N_8864);
or U9117 (N_9117,N_8879,N_8943);
or U9118 (N_9118,N_8989,N_8938);
nor U9119 (N_9119,N_8983,N_8981);
nand U9120 (N_9120,N_8953,N_8904);
nand U9121 (N_9121,N_8973,N_8954);
and U9122 (N_9122,N_8911,N_8901);
nand U9123 (N_9123,N_8972,N_8901);
xor U9124 (N_9124,N_8987,N_8920);
nor U9125 (N_9125,N_8926,N_8903);
and U9126 (N_9126,N_8891,N_8938);
nand U9127 (N_9127,N_8976,N_8918);
and U9128 (N_9128,N_8993,N_8984);
nor U9129 (N_9129,N_8940,N_8865);
xor U9130 (N_9130,N_8910,N_8951);
nand U9131 (N_9131,N_8964,N_8891);
and U9132 (N_9132,N_8929,N_8854);
nand U9133 (N_9133,N_8963,N_8946);
nand U9134 (N_9134,N_8981,N_8927);
nor U9135 (N_9135,N_8898,N_8986);
nor U9136 (N_9136,N_8875,N_8940);
and U9137 (N_9137,N_8894,N_8866);
nor U9138 (N_9138,N_8982,N_8905);
nor U9139 (N_9139,N_8928,N_8893);
and U9140 (N_9140,N_8947,N_8992);
nor U9141 (N_9141,N_8980,N_8887);
and U9142 (N_9142,N_8910,N_8892);
nor U9143 (N_9143,N_8967,N_8903);
and U9144 (N_9144,N_8993,N_8912);
xnor U9145 (N_9145,N_8910,N_8926);
or U9146 (N_9146,N_8916,N_8968);
xnor U9147 (N_9147,N_8965,N_8959);
nor U9148 (N_9148,N_8854,N_8868);
nor U9149 (N_9149,N_8898,N_8946);
nor U9150 (N_9150,N_9057,N_9003);
or U9151 (N_9151,N_9065,N_9109);
and U9152 (N_9152,N_9063,N_9002);
and U9153 (N_9153,N_9047,N_9056);
and U9154 (N_9154,N_9060,N_9114);
nor U9155 (N_9155,N_9007,N_9073);
or U9156 (N_9156,N_9134,N_9145);
and U9157 (N_9157,N_9126,N_9083);
nand U9158 (N_9158,N_9103,N_9029);
nor U9159 (N_9159,N_9024,N_9008);
or U9160 (N_9160,N_9064,N_9019);
and U9161 (N_9161,N_9107,N_9058);
nand U9162 (N_9162,N_9050,N_9105);
and U9163 (N_9163,N_9147,N_9072);
or U9164 (N_9164,N_9006,N_9089);
nor U9165 (N_9165,N_9099,N_9087);
nand U9166 (N_9166,N_9009,N_9020);
xor U9167 (N_9167,N_9055,N_9044);
nor U9168 (N_9168,N_9115,N_9113);
and U9169 (N_9169,N_9075,N_9022);
or U9170 (N_9170,N_9091,N_9021);
or U9171 (N_9171,N_9018,N_9026);
and U9172 (N_9172,N_9040,N_9149);
or U9173 (N_9173,N_9140,N_9052);
and U9174 (N_9174,N_9048,N_9117);
xor U9175 (N_9175,N_9144,N_9093);
nand U9176 (N_9176,N_9088,N_9137);
nor U9177 (N_9177,N_9118,N_9129);
or U9178 (N_9178,N_9030,N_9014);
nand U9179 (N_9179,N_9094,N_9053);
nor U9180 (N_9180,N_9121,N_9049);
or U9181 (N_9181,N_9069,N_9124);
nand U9182 (N_9182,N_9080,N_9092);
and U9183 (N_9183,N_9017,N_9120);
and U9184 (N_9184,N_9133,N_9098);
nand U9185 (N_9185,N_9025,N_9016);
or U9186 (N_9186,N_9061,N_9135);
and U9187 (N_9187,N_9082,N_9031);
nand U9188 (N_9188,N_9015,N_9136);
nor U9189 (N_9189,N_9138,N_9081);
and U9190 (N_9190,N_9085,N_9051);
or U9191 (N_9191,N_9000,N_9128);
xnor U9192 (N_9192,N_9059,N_9027);
nor U9193 (N_9193,N_9076,N_9038);
xnor U9194 (N_9194,N_9039,N_9013);
or U9195 (N_9195,N_9033,N_9077);
and U9196 (N_9196,N_9023,N_9012);
nor U9197 (N_9197,N_9102,N_9005);
or U9198 (N_9198,N_9148,N_9130);
nor U9199 (N_9199,N_9028,N_9146);
or U9200 (N_9200,N_9037,N_9042);
nand U9201 (N_9201,N_9035,N_9067);
nand U9202 (N_9202,N_9074,N_9101);
or U9203 (N_9203,N_9112,N_9086);
or U9204 (N_9204,N_9108,N_9070);
or U9205 (N_9205,N_9062,N_9111);
and U9206 (N_9206,N_9119,N_9127);
and U9207 (N_9207,N_9034,N_9054);
or U9208 (N_9208,N_9122,N_9097);
nor U9209 (N_9209,N_9011,N_9116);
xor U9210 (N_9210,N_9106,N_9090);
nor U9211 (N_9211,N_9142,N_9068);
nand U9212 (N_9212,N_9001,N_9139);
or U9213 (N_9213,N_9046,N_9110);
nand U9214 (N_9214,N_9036,N_9084);
and U9215 (N_9215,N_9096,N_9104);
nor U9216 (N_9216,N_9095,N_9131);
nor U9217 (N_9217,N_9045,N_9041);
nand U9218 (N_9218,N_9032,N_9132);
nor U9219 (N_9219,N_9141,N_9100);
and U9220 (N_9220,N_9010,N_9004);
nand U9221 (N_9221,N_9078,N_9125);
nor U9222 (N_9222,N_9071,N_9066);
and U9223 (N_9223,N_9079,N_9143);
nand U9224 (N_9224,N_9043,N_9123);
or U9225 (N_9225,N_9142,N_9004);
xnor U9226 (N_9226,N_9091,N_9011);
and U9227 (N_9227,N_9005,N_9096);
xor U9228 (N_9228,N_9094,N_9005);
or U9229 (N_9229,N_9063,N_9110);
nand U9230 (N_9230,N_9121,N_9070);
or U9231 (N_9231,N_9002,N_9091);
and U9232 (N_9232,N_9047,N_9089);
or U9233 (N_9233,N_9032,N_9142);
or U9234 (N_9234,N_9080,N_9034);
xor U9235 (N_9235,N_9126,N_9060);
nor U9236 (N_9236,N_9138,N_9014);
and U9237 (N_9237,N_9091,N_9081);
nor U9238 (N_9238,N_9015,N_9011);
and U9239 (N_9239,N_9143,N_9085);
or U9240 (N_9240,N_9088,N_9125);
or U9241 (N_9241,N_9118,N_9015);
and U9242 (N_9242,N_9002,N_9130);
nand U9243 (N_9243,N_9110,N_9061);
nor U9244 (N_9244,N_9128,N_9088);
xnor U9245 (N_9245,N_9125,N_9001);
nand U9246 (N_9246,N_9009,N_9115);
or U9247 (N_9247,N_9033,N_9141);
and U9248 (N_9248,N_9138,N_9061);
nand U9249 (N_9249,N_9059,N_9060);
nand U9250 (N_9250,N_9026,N_9144);
or U9251 (N_9251,N_9104,N_9080);
nand U9252 (N_9252,N_9133,N_9070);
nand U9253 (N_9253,N_9052,N_9005);
or U9254 (N_9254,N_9004,N_9136);
or U9255 (N_9255,N_9053,N_9061);
nor U9256 (N_9256,N_9146,N_9013);
nor U9257 (N_9257,N_9035,N_9033);
nand U9258 (N_9258,N_9104,N_9136);
nand U9259 (N_9259,N_9047,N_9038);
nor U9260 (N_9260,N_9110,N_9087);
nor U9261 (N_9261,N_9020,N_9133);
nor U9262 (N_9262,N_9126,N_9087);
nand U9263 (N_9263,N_9032,N_9031);
nand U9264 (N_9264,N_9075,N_9017);
or U9265 (N_9265,N_9099,N_9041);
or U9266 (N_9266,N_9070,N_9048);
or U9267 (N_9267,N_9100,N_9090);
or U9268 (N_9268,N_9004,N_9001);
xnor U9269 (N_9269,N_9082,N_9077);
nand U9270 (N_9270,N_9121,N_9002);
and U9271 (N_9271,N_9072,N_9146);
or U9272 (N_9272,N_9005,N_9047);
nor U9273 (N_9273,N_9042,N_9029);
nor U9274 (N_9274,N_9014,N_9108);
nand U9275 (N_9275,N_9077,N_9084);
and U9276 (N_9276,N_9122,N_9136);
nand U9277 (N_9277,N_9091,N_9100);
nand U9278 (N_9278,N_9112,N_9144);
nand U9279 (N_9279,N_9130,N_9061);
and U9280 (N_9280,N_9047,N_9077);
nand U9281 (N_9281,N_9018,N_9016);
and U9282 (N_9282,N_9144,N_9097);
and U9283 (N_9283,N_9013,N_9098);
nor U9284 (N_9284,N_9081,N_9112);
nor U9285 (N_9285,N_9016,N_9070);
nand U9286 (N_9286,N_9047,N_9081);
and U9287 (N_9287,N_9081,N_9128);
and U9288 (N_9288,N_9018,N_9146);
nor U9289 (N_9289,N_9109,N_9124);
nor U9290 (N_9290,N_9143,N_9107);
nor U9291 (N_9291,N_9061,N_9147);
nand U9292 (N_9292,N_9082,N_9064);
and U9293 (N_9293,N_9113,N_9048);
nand U9294 (N_9294,N_9086,N_9065);
or U9295 (N_9295,N_9078,N_9022);
nor U9296 (N_9296,N_9037,N_9133);
and U9297 (N_9297,N_9052,N_9013);
and U9298 (N_9298,N_9022,N_9137);
or U9299 (N_9299,N_9110,N_9070);
nor U9300 (N_9300,N_9227,N_9264);
nor U9301 (N_9301,N_9176,N_9289);
xor U9302 (N_9302,N_9153,N_9156);
nor U9303 (N_9303,N_9206,N_9291);
nor U9304 (N_9304,N_9271,N_9190);
nand U9305 (N_9305,N_9225,N_9188);
and U9306 (N_9306,N_9224,N_9258);
or U9307 (N_9307,N_9296,N_9164);
nor U9308 (N_9308,N_9237,N_9185);
or U9309 (N_9309,N_9154,N_9297);
nor U9310 (N_9310,N_9223,N_9247);
and U9311 (N_9311,N_9159,N_9282);
or U9312 (N_9312,N_9279,N_9201);
nand U9313 (N_9313,N_9276,N_9250);
and U9314 (N_9314,N_9230,N_9168);
xnor U9315 (N_9315,N_9261,N_9166);
nor U9316 (N_9316,N_9204,N_9212);
nor U9317 (N_9317,N_9244,N_9281);
nor U9318 (N_9318,N_9290,N_9200);
nor U9319 (N_9319,N_9266,N_9208);
nand U9320 (N_9320,N_9184,N_9293);
xnor U9321 (N_9321,N_9161,N_9202);
nor U9322 (N_9322,N_9243,N_9231);
and U9323 (N_9323,N_9182,N_9183);
nor U9324 (N_9324,N_9170,N_9292);
or U9325 (N_9325,N_9285,N_9259);
nor U9326 (N_9326,N_9226,N_9192);
xor U9327 (N_9327,N_9277,N_9254);
xnor U9328 (N_9328,N_9288,N_9160);
or U9329 (N_9329,N_9205,N_9255);
and U9330 (N_9330,N_9236,N_9217);
nor U9331 (N_9331,N_9169,N_9253);
nor U9332 (N_9332,N_9220,N_9171);
xnor U9333 (N_9333,N_9197,N_9219);
nor U9334 (N_9334,N_9260,N_9234);
nand U9335 (N_9335,N_9194,N_9249);
and U9336 (N_9336,N_9216,N_9270);
nor U9337 (N_9337,N_9193,N_9207);
nand U9338 (N_9338,N_9283,N_9240);
nor U9339 (N_9339,N_9242,N_9252);
and U9340 (N_9340,N_9211,N_9203);
and U9341 (N_9341,N_9175,N_9172);
and U9342 (N_9342,N_9246,N_9295);
and U9343 (N_9343,N_9165,N_9162);
nand U9344 (N_9344,N_9229,N_9241);
xnor U9345 (N_9345,N_9280,N_9245);
and U9346 (N_9346,N_9174,N_9178);
nand U9347 (N_9347,N_9209,N_9298);
or U9348 (N_9348,N_9198,N_9268);
or U9349 (N_9349,N_9235,N_9195);
nor U9350 (N_9350,N_9157,N_9187);
nand U9351 (N_9351,N_9181,N_9278);
xnor U9352 (N_9352,N_9155,N_9186);
nor U9353 (N_9353,N_9180,N_9218);
nor U9354 (N_9354,N_9228,N_9233);
or U9355 (N_9355,N_9191,N_9151);
or U9356 (N_9356,N_9167,N_9286);
nand U9357 (N_9357,N_9251,N_9196);
or U9358 (N_9358,N_9152,N_9274);
nand U9359 (N_9359,N_9265,N_9238);
nand U9360 (N_9360,N_9158,N_9232);
and U9361 (N_9361,N_9199,N_9163);
or U9362 (N_9362,N_9215,N_9189);
or U9363 (N_9363,N_9257,N_9173);
nor U9364 (N_9364,N_9262,N_9222);
and U9365 (N_9365,N_9239,N_9299);
xor U9366 (N_9366,N_9213,N_9177);
nor U9367 (N_9367,N_9269,N_9256);
nand U9368 (N_9368,N_9248,N_9179);
and U9369 (N_9369,N_9294,N_9267);
or U9370 (N_9370,N_9150,N_9284);
and U9371 (N_9371,N_9263,N_9272);
nand U9372 (N_9372,N_9273,N_9275);
or U9373 (N_9373,N_9287,N_9210);
or U9374 (N_9374,N_9221,N_9214);
nor U9375 (N_9375,N_9263,N_9211);
or U9376 (N_9376,N_9190,N_9254);
nor U9377 (N_9377,N_9272,N_9236);
or U9378 (N_9378,N_9161,N_9223);
nor U9379 (N_9379,N_9151,N_9270);
or U9380 (N_9380,N_9235,N_9292);
nor U9381 (N_9381,N_9211,N_9293);
nor U9382 (N_9382,N_9244,N_9162);
or U9383 (N_9383,N_9195,N_9243);
nor U9384 (N_9384,N_9224,N_9253);
and U9385 (N_9385,N_9164,N_9298);
or U9386 (N_9386,N_9222,N_9169);
and U9387 (N_9387,N_9291,N_9220);
nand U9388 (N_9388,N_9174,N_9258);
or U9389 (N_9389,N_9247,N_9267);
and U9390 (N_9390,N_9278,N_9219);
or U9391 (N_9391,N_9196,N_9261);
and U9392 (N_9392,N_9246,N_9198);
or U9393 (N_9393,N_9280,N_9201);
nor U9394 (N_9394,N_9168,N_9176);
or U9395 (N_9395,N_9239,N_9160);
nand U9396 (N_9396,N_9289,N_9225);
and U9397 (N_9397,N_9285,N_9299);
nor U9398 (N_9398,N_9289,N_9218);
or U9399 (N_9399,N_9179,N_9217);
or U9400 (N_9400,N_9224,N_9216);
or U9401 (N_9401,N_9270,N_9233);
or U9402 (N_9402,N_9245,N_9181);
or U9403 (N_9403,N_9246,N_9293);
nor U9404 (N_9404,N_9198,N_9260);
and U9405 (N_9405,N_9273,N_9194);
or U9406 (N_9406,N_9266,N_9192);
nand U9407 (N_9407,N_9254,N_9212);
nand U9408 (N_9408,N_9233,N_9238);
and U9409 (N_9409,N_9187,N_9209);
nor U9410 (N_9410,N_9189,N_9263);
or U9411 (N_9411,N_9225,N_9266);
or U9412 (N_9412,N_9171,N_9295);
nor U9413 (N_9413,N_9186,N_9160);
and U9414 (N_9414,N_9186,N_9234);
and U9415 (N_9415,N_9244,N_9285);
or U9416 (N_9416,N_9234,N_9294);
nor U9417 (N_9417,N_9205,N_9236);
or U9418 (N_9418,N_9285,N_9291);
and U9419 (N_9419,N_9255,N_9180);
and U9420 (N_9420,N_9203,N_9243);
nand U9421 (N_9421,N_9251,N_9192);
nor U9422 (N_9422,N_9205,N_9150);
nand U9423 (N_9423,N_9290,N_9193);
or U9424 (N_9424,N_9264,N_9191);
and U9425 (N_9425,N_9163,N_9206);
nand U9426 (N_9426,N_9215,N_9247);
and U9427 (N_9427,N_9183,N_9224);
nor U9428 (N_9428,N_9246,N_9248);
and U9429 (N_9429,N_9266,N_9294);
and U9430 (N_9430,N_9283,N_9192);
nand U9431 (N_9431,N_9250,N_9272);
or U9432 (N_9432,N_9227,N_9177);
or U9433 (N_9433,N_9180,N_9282);
nand U9434 (N_9434,N_9267,N_9254);
or U9435 (N_9435,N_9260,N_9263);
xnor U9436 (N_9436,N_9183,N_9256);
nor U9437 (N_9437,N_9270,N_9268);
xnor U9438 (N_9438,N_9205,N_9299);
or U9439 (N_9439,N_9189,N_9175);
nand U9440 (N_9440,N_9280,N_9184);
xnor U9441 (N_9441,N_9226,N_9196);
or U9442 (N_9442,N_9260,N_9267);
or U9443 (N_9443,N_9167,N_9216);
and U9444 (N_9444,N_9152,N_9168);
nand U9445 (N_9445,N_9239,N_9200);
nand U9446 (N_9446,N_9254,N_9214);
or U9447 (N_9447,N_9233,N_9153);
xnor U9448 (N_9448,N_9216,N_9269);
and U9449 (N_9449,N_9295,N_9161);
and U9450 (N_9450,N_9425,N_9370);
xor U9451 (N_9451,N_9392,N_9339);
or U9452 (N_9452,N_9366,N_9361);
or U9453 (N_9453,N_9341,N_9374);
nor U9454 (N_9454,N_9357,N_9420);
xor U9455 (N_9455,N_9421,N_9411);
or U9456 (N_9456,N_9423,N_9353);
or U9457 (N_9457,N_9356,N_9338);
nor U9458 (N_9458,N_9318,N_9383);
and U9459 (N_9459,N_9429,N_9372);
nor U9460 (N_9460,N_9319,N_9344);
or U9461 (N_9461,N_9363,N_9419);
and U9462 (N_9462,N_9393,N_9431);
nor U9463 (N_9463,N_9324,N_9352);
or U9464 (N_9464,N_9409,N_9444);
or U9465 (N_9465,N_9301,N_9428);
or U9466 (N_9466,N_9336,N_9384);
nor U9467 (N_9467,N_9448,N_9343);
nor U9468 (N_9468,N_9406,N_9333);
and U9469 (N_9469,N_9382,N_9377);
or U9470 (N_9470,N_9371,N_9325);
nor U9471 (N_9471,N_9368,N_9327);
nand U9472 (N_9472,N_9334,N_9446);
xor U9473 (N_9473,N_9426,N_9306);
nand U9474 (N_9474,N_9354,N_9331);
xor U9475 (N_9475,N_9346,N_9380);
nor U9476 (N_9476,N_9323,N_9410);
xnor U9477 (N_9477,N_9304,N_9391);
and U9478 (N_9478,N_9376,N_9389);
and U9479 (N_9479,N_9432,N_9300);
and U9480 (N_9480,N_9345,N_9385);
and U9481 (N_9481,N_9396,N_9309);
and U9482 (N_9482,N_9449,N_9332);
nor U9483 (N_9483,N_9404,N_9360);
or U9484 (N_9484,N_9315,N_9326);
and U9485 (N_9485,N_9388,N_9347);
or U9486 (N_9486,N_9413,N_9373);
nor U9487 (N_9487,N_9439,N_9310);
nor U9488 (N_9488,N_9364,N_9395);
nor U9489 (N_9489,N_9399,N_9422);
xor U9490 (N_9490,N_9375,N_9387);
and U9491 (N_9491,N_9302,N_9442);
nor U9492 (N_9492,N_9427,N_9416);
and U9493 (N_9493,N_9443,N_9348);
nor U9494 (N_9494,N_9414,N_9381);
nand U9495 (N_9495,N_9436,N_9328);
and U9496 (N_9496,N_9314,N_9320);
or U9497 (N_9497,N_9313,N_9312);
and U9498 (N_9498,N_9316,N_9350);
or U9499 (N_9499,N_9405,N_9397);
or U9500 (N_9500,N_9358,N_9330);
nand U9501 (N_9501,N_9433,N_9305);
xor U9502 (N_9502,N_9390,N_9438);
xnor U9503 (N_9503,N_9403,N_9430);
and U9504 (N_9504,N_9386,N_9340);
or U9505 (N_9505,N_9308,N_9398);
nand U9506 (N_9506,N_9317,N_9441);
nor U9507 (N_9507,N_9407,N_9367);
xnor U9508 (N_9508,N_9378,N_9342);
and U9509 (N_9509,N_9303,N_9447);
nand U9510 (N_9510,N_9307,N_9362);
or U9511 (N_9511,N_9412,N_9437);
or U9512 (N_9512,N_9418,N_9415);
and U9513 (N_9513,N_9337,N_9408);
or U9514 (N_9514,N_9401,N_9402);
or U9515 (N_9515,N_9394,N_9335);
or U9516 (N_9516,N_9435,N_9349);
nand U9517 (N_9517,N_9351,N_9311);
and U9518 (N_9518,N_9445,N_9434);
and U9519 (N_9519,N_9379,N_9369);
nand U9520 (N_9520,N_9321,N_9365);
nand U9521 (N_9521,N_9322,N_9440);
and U9522 (N_9522,N_9417,N_9400);
nor U9523 (N_9523,N_9359,N_9329);
or U9524 (N_9524,N_9424,N_9355);
or U9525 (N_9525,N_9375,N_9432);
nand U9526 (N_9526,N_9374,N_9309);
nor U9527 (N_9527,N_9428,N_9418);
or U9528 (N_9528,N_9426,N_9435);
and U9529 (N_9529,N_9385,N_9404);
nand U9530 (N_9530,N_9333,N_9398);
and U9531 (N_9531,N_9342,N_9307);
or U9532 (N_9532,N_9350,N_9429);
nor U9533 (N_9533,N_9386,N_9365);
nor U9534 (N_9534,N_9424,N_9438);
nand U9535 (N_9535,N_9362,N_9379);
and U9536 (N_9536,N_9428,N_9449);
or U9537 (N_9537,N_9341,N_9363);
and U9538 (N_9538,N_9380,N_9372);
nor U9539 (N_9539,N_9375,N_9391);
and U9540 (N_9540,N_9443,N_9430);
or U9541 (N_9541,N_9390,N_9380);
nand U9542 (N_9542,N_9324,N_9349);
and U9543 (N_9543,N_9418,N_9305);
nand U9544 (N_9544,N_9444,N_9436);
and U9545 (N_9545,N_9333,N_9340);
and U9546 (N_9546,N_9354,N_9305);
and U9547 (N_9547,N_9333,N_9321);
nor U9548 (N_9548,N_9412,N_9354);
and U9549 (N_9549,N_9402,N_9429);
xnor U9550 (N_9550,N_9313,N_9320);
nand U9551 (N_9551,N_9381,N_9304);
and U9552 (N_9552,N_9403,N_9393);
nor U9553 (N_9553,N_9413,N_9375);
or U9554 (N_9554,N_9331,N_9443);
xnor U9555 (N_9555,N_9371,N_9337);
and U9556 (N_9556,N_9388,N_9431);
nand U9557 (N_9557,N_9321,N_9407);
nor U9558 (N_9558,N_9322,N_9327);
nor U9559 (N_9559,N_9342,N_9356);
xnor U9560 (N_9560,N_9443,N_9339);
nor U9561 (N_9561,N_9305,N_9383);
or U9562 (N_9562,N_9301,N_9438);
nor U9563 (N_9563,N_9396,N_9409);
nand U9564 (N_9564,N_9443,N_9338);
xnor U9565 (N_9565,N_9442,N_9377);
nand U9566 (N_9566,N_9363,N_9449);
nand U9567 (N_9567,N_9442,N_9411);
or U9568 (N_9568,N_9328,N_9441);
xor U9569 (N_9569,N_9379,N_9319);
and U9570 (N_9570,N_9414,N_9384);
and U9571 (N_9571,N_9396,N_9395);
and U9572 (N_9572,N_9354,N_9323);
nand U9573 (N_9573,N_9428,N_9423);
or U9574 (N_9574,N_9428,N_9340);
nand U9575 (N_9575,N_9361,N_9448);
or U9576 (N_9576,N_9384,N_9300);
and U9577 (N_9577,N_9387,N_9442);
nor U9578 (N_9578,N_9383,N_9443);
or U9579 (N_9579,N_9391,N_9373);
and U9580 (N_9580,N_9380,N_9343);
nand U9581 (N_9581,N_9372,N_9365);
nand U9582 (N_9582,N_9363,N_9435);
and U9583 (N_9583,N_9343,N_9424);
nor U9584 (N_9584,N_9311,N_9336);
or U9585 (N_9585,N_9447,N_9382);
nand U9586 (N_9586,N_9313,N_9425);
and U9587 (N_9587,N_9389,N_9302);
or U9588 (N_9588,N_9391,N_9368);
nand U9589 (N_9589,N_9402,N_9390);
or U9590 (N_9590,N_9381,N_9398);
xnor U9591 (N_9591,N_9404,N_9436);
or U9592 (N_9592,N_9366,N_9358);
or U9593 (N_9593,N_9309,N_9425);
nand U9594 (N_9594,N_9410,N_9408);
xnor U9595 (N_9595,N_9420,N_9359);
nand U9596 (N_9596,N_9424,N_9366);
or U9597 (N_9597,N_9398,N_9402);
nor U9598 (N_9598,N_9328,N_9376);
or U9599 (N_9599,N_9313,N_9323);
nor U9600 (N_9600,N_9573,N_9495);
nand U9601 (N_9601,N_9542,N_9456);
nor U9602 (N_9602,N_9520,N_9560);
nand U9603 (N_9603,N_9535,N_9544);
nor U9604 (N_9604,N_9549,N_9530);
nor U9605 (N_9605,N_9484,N_9551);
nand U9606 (N_9606,N_9552,N_9509);
and U9607 (N_9607,N_9485,N_9585);
nand U9608 (N_9608,N_9505,N_9471);
and U9609 (N_9609,N_9525,N_9515);
or U9610 (N_9610,N_9540,N_9579);
nand U9611 (N_9611,N_9536,N_9528);
and U9612 (N_9612,N_9498,N_9455);
or U9613 (N_9613,N_9464,N_9458);
xor U9614 (N_9614,N_9516,N_9465);
and U9615 (N_9615,N_9514,N_9527);
or U9616 (N_9616,N_9594,N_9575);
nand U9617 (N_9617,N_9593,N_9591);
or U9618 (N_9618,N_9538,N_9453);
or U9619 (N_9619,N_9474,N_9497);
nand U9620 (N_9620,N_9496,N_9492);
nand U9621 (N_9621,N_9451,N_9524);
or U9622 (N_9622,N_9532,N_9486);
or U9623 (N_9623,N_9550,N_9555);
nand U9624 (N_9624,N_9523,N_9543);
xor U9625 (N_9625,N_9491,N_9480);
nor U9626 (N_9626,N_9577,N_9467);
nor U9627 (N_9627,N_9508,N_9469);
and U9628 (N_9628,N_9468,N_9513);
xor U9629 (N_9629,N_9569,N_9586);
or U9630 (N_9630,N_9481,N_9570);
xnor U9631 (N_9631,N_9587,N_9534);
xnor U9632 (N_9632,N_9592,N_9487);
nor U9633 (N_9633,N_9489,N_9501);
nor U9634 (N_9634,N_9598,N_9507);
xnor U9635 (N_9635,N_9460,N_9562);
nand U9636 (N_9636,N_9574,N_9559);
nor U9637 (N_9637,N_9561,N_9479);
or U9638 (N_9638,N_9596,N_9541);
and U9639 (N_9639,N_9580,N_9565);
or U9640 (N_9640,N_9472,N_9459);
nand U9641 (N_9641,N_9522,N_9450);
nor U9642 (N_9642,N_9556,N_9462);
or U9643 (N_9643,N_9548,N_9457);
nand U9644 (N_9644,N_9521,N_9564);
or U9645 (N_9645,N_9599,N_9510);
nand U9646 (N_9646,N_9519,N_9483);
nor U9647 (N_9647,N_9533,N_9539);
nand U9648 (N_9648,N_9563,N_9494);
and U9649 (N_9649,N_9576,N_9566);
or U9650 (N_9650,N_9557,N_9572);
or U9651 (N_9651,N_9503,N_9470);
and U9652 (N_9652,N_9517,N_9499);
nand U9653 (N_9653,N_9490,N_9506);
or U9654 (N_9654,N_9553,N_9578);
and U9655 (N_9655,N_9473,N_9526);
nor U9656 (N_9656,N_9581,N_9454);
nor U9657 (N_9657,N_9475,N_9582);
nor U9658 (N_9658,N_9545,N_9554);
nand U9659 (N_9659,N_9589,N_9511);
and U9660 (N_9660,N_9567,N_9482);
nand U9661 (N_9661,N_9537,N_9568);
and U9662 (N_9662,N_9583,N_9584);
xor U9663 (N_9663,N_9518,N_9531);
xnor U9664 (N_9664,N_9477,N_9512);
nor U9665 (N_9665,N_9461,N_9571);
nand U9666 (N_9666,N_9463,N_9500);
and U9667 (N_9667,N_9466,N_9597);
or U9668 (N_9668,N_9452,N_9476);
or U9669 (N_9669,N_9546,N_9529);
or U9670 (N_9670,N_9504,N_9558);
nand U9671 (N_9671,N_9478,N_9547);
or U9672 (N_9672,N_9502,N_9493);
nand U9673 (N_9673,N_9588,N_9590);
nor U9674 (N_9674,N_9595,N_9488);
nand U9675 (N_9675,N_9505,N_9543);
and U9676 (N_9676,N_9511,N_9487);
nor U9677 (N_9677,N_9578,N_9502);
nand U9678 (N_9678,N_9496,N_9555);
or U9679 (N_9679,N_9510,N_9514);
xor U9680 (N_9680,N_9480,N_9500);
and U9681 (N_9681,N_9570,N_9539);
xnor U9682 (N_9682,N_9582,N_9559);
nand U9683 (N_9683,N_9535,N_9477);
nor U9684 (N_9684,N_9453,N_9514);
nand U9685 (N_9685,N_9564,N_9559);
nor U9686 (N_9686,N_9537,N_9545);
nand U9687 (N_9687,N_9500,N_9550);
nand U9688 (N_9688,N_9523,N_9468);
nor U9689 (N_9689,N_9509,N_9540);
or U9690 (N_9690,N_9519,N_9454);
and U9691 (N_9691,N_9458,N_9551);
or U9692 (N_9692,N_9478,N_9483);
nor U9693 (N_9693,N_9552,N_9513);
or U9694 (N_9694,N_9496,N_9464);
or U9695 (N_9695,N_9468,N_9500);
and U9696 (N_9696,N_9542,N_9594);
and U9697 (N_9697,N_9535,N_9558);
nor U9698 (N_9698,N_9509,N_9516);
nand U9699 (N_9699,N_9467,N_9511);
and U9700 (N_9700,N_9561,N_9452);
or U9701 (N_9701,N_9493,N_9478);
nor U9702 (N_9702,N_9505,N_9465);
or U9703 (N_9703,N_9554,N_9581);
nor U9704 (N_9704,N_9488,N_9462);
nor U9705 (N_9705,N_9457,N_9563);
nor U9706 (N_9706,N_9509,N_9534);
nand U9707 (N_9707,N_9451,N_9589);
nor U9708 (N_9708,N_9596,N_9456);
and U9709 (N_9709,N_9472,N_9470);
and U9710 (N_9710,N_9594,N_9454);
and U9711 (N_9711,N_9515,N_9547);
nand U9712 (N_9712,N_9509,N_9522);
and U9713 (N_9713,N_9541,N_9527);
nand U9714 (N_9714,N_9541,N_9529);
nor U9715 (N_9715,N_9553,N_9505);
or U9716 (N_9716,N_9575,N_9533);
nand U9717 (N_9717,N_9498,N_9511);
or U9718 (N_9718,N_9560,N_9536);
nor U9719 (N_9719,N_9588,N_9472);
or U9720 (N_9720,N_9472,N_9573);
and U9721 (N_9721,N_9477,N_9581);
nand U9722 (N_9722,N_9515,N_9555);
nor U9723 (N_9723,N_9565,N_9509);
nor U9724 (N_9724,N_9592,N_9486);
or U9725 (N_9725,N_9500,N_9575);
and U9726 (N_9726,N_9479,N_9593);
or U9727 (N_9727,N_9469,N_9544);
and U9728 (N_9728,N_9516,N_9575);
nor U9729 (N_9729,N_9482,N_9450);
nand U9730 (N_9730,N_9573,N_9524);
xnor U9731 (N_9731,N_9491,N_9582);
nor U9732 (N_9732,N_9590,N_9520);
and U9733 (N_9733,N_9598,N_9465);
and U9734 (N_9734,N_9508,N_9470);
and U9735 (N_9735,N_9599,N_9452);
or U9736 (N_9736,N_9599,N_9513);
or U9737 (N_9737,N_9565,N_9583);
nand U9738 (N_9738,N_9588,N_9558);
or U9739 (N_9739,N_9503,N_9480);
nand U9740 (N_9740,N_9561,N_9469);
nand U9741 (N_9741,N_9583,N_9536);
and U9742 (N_9742,N_9482,N_9460);
or U9743 (N_9743,N_9491,N_9554);
and U9744 (N_9744,N_9599,N_9524);
nor U9745 (N_9745,N_9486,N_9454);
nand U9746 (N_9746,N_9476,N_9575);
nor U9747 (N_9747,N_9516,N_9550);
xnor U9748 (N_9748,N_9541,N_9458);
nor U9749 (N_9749,N_9554,N_9541);
and U9750 (N_9750,N_9662,N_9714);
nor U9751 (N_9751,N_9637,N_9740);
xnor U9752 (N_9752,N_9603,N_9649);
xor U9753 (N_9753,N_9707,N_9731);
nand U9754 (N_9754,N_9627,N_9695);
xnor U9755 (N_9755,N_9680,N_9720);
or U9756 (N_9756,N_9729,N_9696);
nor U9757 (N_9757,N_9744,N_9683);
or U9758 (N_9758,N_9640,N_9619);
and U9759 (N_9759,N_9721,N_9736);
and U9760 (N_9760,N_9608,N_9703);
xor U9761 (N_9761,N_9699,N_9725);
or U9762 (N_9762,N_9678,N_9743);
and U9763 (N_9763,N_9688,N_9613);
nor U9764 (N_9764,N_9705,N_9664);
or U9765 (N_9765,N_9681,N_9702);
or U9766 (N_9766,N_9738,N_9647);
nand U9767 (N_9767,N_9713,N_9636);
or U9768 (N_9768,N_9665,N_9739);
nor U9769 (N_9769,N_9661,N_9607);
nand U9770 (N_9770,N_9685,N_9717);
xnor U9771 (N_9771,N_9676,N_9642);
and U9772 (N_9772,N_9711,N_9633);
nand U9773 (N_9773,N_9639,N_9691);
nor U9774 (N_9774,N_9657,N_9614);
nor U9775 (N_9775,N_9622,N_9704);
xnor U9776 (N_9776,N_9667,N_9635);
or U9777 (N_9777,N_9710,N_9708);
and U9778 (N_9778,N_9656,N_9646);
and U9779 (N_9779,N_9727,N_9623);
nor U9780 (N_9780,N_9687,N_9610);
nand U9781 (N_9781,N_9722,N_9611);
or U9782 (N_9782,N_9605,N_9631);
nand U9783 (N_9783,N_9615,N_9666);
xnor U9784 (N_9784,N_9650,N_9748);
or U9785 (N_9785,N_9670,N_9658);
or U9786 (N_9786,N_9716,N_9625);
nor U9787 (N_9787,N_9629,N_9644);
nand U9788 (N_9788,N_9745,N_9674);
nand U9789 (N_9789,N_9728,N_9673);
xor U9790 (N_9790,N_9724,N_9634);
and U9791 (N_9791,N_9689,N_9630);
and U9792 (N_9792,N_9718,N_9672);
nand U9793 (N_9793,N_9715,N_9621);
nor U9794 (N_9794,N_9609,N_9620);
nor U9795 (N_9795,N_9660,N_9677);
or U9796 (N_9796,N_9632,N_9641);
and U9797 (N_9797,N_9675,N_9749);
nor U9798 (N_9798,N_9746,N_9730);
nor U9799 (N_9799,N_9700,N_9747);
nand U9800 (N_9800,N_9719,N_9638);
and U9801 (N_9801,N_9628,N_9697);
and U9802 (N_9802,N_9686,N_9617);
and U9803 (N_9803,N_9692,N_9669);
and U9804 (N_9804,N_9732,N_9653);
and U9805 (N_9805,N_9618,N_9709);
or U9806 (N_9806,N_9684,N_9624);
and U9807 (N_9807,N_9682,N_9741);
nand U9808 (N_9808,N_9742,N_9626);
nor U9809 (N_9809,N_9606,N_9712);
and U9810 (N_9810,N_9706,N_9690);
and U9811 (N_9811,N_9601,N_9663);
nand U9812 (N_9812,N_9726,N_9679);
or U9813 (N_9813,N_9659,N_9604);
nor U9814 (N_9814,N_9645,N_9648);
and U9815 (N_9815,N_9651,N_9735);
nor U9816 (N_9816,N_9643,N_9733);
nand U9817 (N_9817,N_9734,N_9616);
nor U9818 (N_9818,N_9723,N_9600);
nand U9819 (N_9819,N_9654,N_9602);
nor U9820 (N_9820,N_9671,N_9652);
and U9821 (N_9821,N_9737,N_9655);
and U9822 (N_9822,N_9612,N_9701);
or U9823 (N_9823,N_9694,N_9693);
nand U9824 (N_9824,N_9698,N_9668);
nor U9825 (N_9825,N_9612,N_9747);
nor U9826 (N_9826,N_9634,N_9625);
nor U9827 (N_9827,N_9651,N_9615);
xnor U9828 (N_9828,N_9662,N_9605);
nor U9829 (N_9829,N_9704,N_9652);
nand U9830 (N_9830,N_9600,N_9627);
or U9831 (N_9831,N_9706,N_9693);
nor U9832 (N_9832,N_9651,N_9662);
nand U9833 (N_9833,N_9708,N_9664);
nor U9834 (N_9834,N_9630,N_9701);
nand U9835 (N_9835,N_9602,N_9743);
or U9836 (N_9836,N_9696,N_9722);
and U9837 (N_9837,N_9654,N_9723);
nand U9838 (N_9838,N_9681,N_9667);
and U9839 (N_9839,N_9698,N_9643);
nor U9840 (N_9840,N_9605,N_9721);
or U9841 (N_9841,N_9626,N_9721);
xnor U9842 (N_9842,N_9673,N_9670);
and U9843 (N_9843,N_9645,N_9714);
nor U9844 (N_9844,N_9627,N_9746);
nand U9845 (N_9845,N_9726,N_9715);
or U9846 (N_9846,N_9740,N_9638);
and U9847 (N_9847,N_9663,N_9683);
xnor U9848 (N_9848,N_9687,N_9670);
nor U9849 (N_9849,N_9741,N_9729);
or U9850 (N_9850,N_9698,N_9619);
xnor U9851 (N_9851,N_9616,N_9651);
nor U9852 (N_9852,N_9640,N_9673);
and U9853 (N_9853,N_9708,N_9602);
nand U9854 (N_9854,N_9718,N_9686);
and U9855 (N_9855,N_9600,N_9705);
xor U9856 (N_9856,N_9695,N_9620);
nand U9857 (N_9857,N_9629,N_9736);
nor U9858 (N_9858,N_9686,N_9682);
and U9859 (N_9859,N_9666,N_9654);
and U9860 (N_9860,N_9671,N_9739);
xnor U9861 (N_9861,N_9663,N_9629);
xnor U9862 (N_9862,N_9665,N_9729);
xor U9863 (N_9863,N_9636,N_9708);
nand U9864 (N_9864,N_9648,N_9601);
or U9865 (N_9865,N_9615,N_9723);
nor U9866 (N_9866,N_9698,N_9709);
nor U9867 (N_9867,N_9684,N_9741);
and U9868 (N_9868,N_9695,N_9644);
and U9869 (N_9869,N_9689,N_9720);
nor U9870 (N_9870,N_9636,N_9679);
nor U9871 (N_9871,N_9684,N_9633);
or U9872 (N_9872,N_9715,N_9617);
nor U9873 (N_9873,N_9632,N_9665);
nor U9874 (N_9874,N_9630,N_9680);
or U9875 (N_9875,N_9649,N_9627);
nor U9876 (N_9876,N_9676,N_9699);
nand U9877 (N_9877,N_9649,N_9700);
or U9878 (N_9878,N_9712,N_9682);
xnor U9879 (N_9879,N_9740,N_9735);
nor U9880 (N_9880,N_9622,N_9626);
nor U9881 (N_9881,N_9693,N_9730);
and U9882 (N_9882,N_9660,N_9641);
nor U9883 (N_9883,N_9706,N_9625);
or U9884 (N_9884,N_9717,N_9658);
and U9885 (N_9885,N_9615,N_9658);
or U9886 (N_9886,N_9650,N_9729);
nand U9887 (N_9887,N_9643,N_9641);
nand U9888 (N_9888,N_9637,N_9689);
and U9889 (N_9889,N_9701,N_9728);
and U9890 (N_9890,N_9737,N_9651);
nand U9891 (N_9891,N_9722,N_9709);
and U9892 (N_9892,N_9705,N_9611);
or U9893 (N_9893,N_9732,N_9619);
nand U9894 (N_9894,N_9731,N_9679);
nor U9895 (N_9895,N_9676,N_9715);
nor U9896 (N_9896,N_9692,N_9618);
nand U9897 (N_9897,N_9616,N_9606);
and U9898 (N_9898,N_9672,N_9700);
or U9899 (N_9899,N_9690,N_9647);
or U9900 (N_9900,N_9773,N_9802);
xor U9901 (N_9901,N_9861,N_9766);
xor U9902 (N_9902,N_9870,N_9791);
nand U9903 (N_9903,N_9807,N_9768);
or U9904 (N_9904,N_9827,N_9760);
xor U9905 (N_9905,N_9793,N_9843);
nand U9906 (N_9906,N_9894,N_9761);
xnor U9907 (N_9907,N_9775,N_9830);
nand U9908 (N_9908,N_9875,N_9770);
xnor U9909 (N_9909,N_9840,N_9753);
xnor U9910 (N_9910,N_9757,N_9826);
or U9911 (N_9911,N_9790,N_9871);
nor U9912 (N_9912,N_9835,N_9891);
nand U9913 (N_9913,N_9774,N_9823);
nand U9914 (N_9914,N_9813,N_9805);
or U9915 (N_9915,N_9795,N_9881);
and U9916 (N_9916,N_9824,N_9752);
nand U9917 (N_9917,N_9819,N_9799);
and U9918 (N_9918,N_9817,N_9780);
nand U9919 (N_9919,N_9886,N_9837);
nor U9920 (N_9920,N_9816,N_9857);
nand U9921 (N_9921,N_9804,N_9789);
and U9922 (N_9922,N_9862,N_9765);
or U9923 (N_9923,N_9820,N_9899);
xnor U9924 (N_9924,N_9818,N_9821);
and U9925 (N_9925,N_9801,N_9879);
nor U9926 (N_9926,N_9772,N_9898);
xnor U9927 (N_9927,N_9853,N_9777);
xor U9928 (N_9928,N_9859,N_9841);
and U9929 (N_9929,N_9897,N_9781);
and U9930 (N_9930,N_9750,N_9833);
and U9931 (N_9931,N_9822,N_9872);
nand U9932 (N_9932,N_9842,N_9778);
and U9933 (N_9933,N_9769,N_9832);
and U9934 (N_9934,N_9812,N_9759);
or U9935 (N_9935,N_9852,N_9783);
or U9936 (N_9936,N_9851,N_9864);
nand U9937 (N_9937,N_9803,N_9885);
or U9938 (N_9938,N_9839,N_9877);
xnor U9939 (N_9939,N_9874,N_9856);
nand U9940 (N_9940,N_9882,N_9866);
nor U9941 (N_9941,N_9828,N_9779);
nor U9942 (N_9942,N_9858,N_9845);
and U9943 (N_9943,N_9836,N_9814);
nor U9944 (N_9944,N_9887,N_9834);
or U9945 (N_9945,N_9798,N_9878);
nor U9946 (N_9946,N_9800,N_9844);
or U9947 (N_9947,N_9896,N_9829);
nand U9948 (N_9948,N_9786,N_9763);
and U9949 (N_9949,N_9806,N_9854);
or U9950 (N_9950,N_9809,N_9811);
and U9951 (N_9951,N_9838,N_9855);
and U9952 (N_9952,N_9884,N_9767);
nand U9953 (N_9953,N_9762,N_9756);
nor U9954 (N_9954,N_9776,N_9847);
nor U9955 (N_9955,N_9880,N_9849);
nor U9956 (N_9956,N_9848,N_9888);
nand U9957 (N_9957,N_9782,N_9784);
nor U9958 (N_9958,N_9758,N_9846);
nand U9959 (N_9959,N_9764,N_9796);
or U9960 (N_9960,N_9825,N_9868);
nor U9961 (N_9961,N_9771,N_9869);
and U9962 (N_9962,N_9863,N_9873);
nor U9963 (N_9963,N_9895,N_9867);
nor U9964 (N_9964,N_9850,N_9876);
or U9965 (N_9965,N_9785,N_9794);
or U9966 (N_9966,N_9892,N_9810);
nand U9967 (N_9967,N_9755,N_9893);
nor U9968 (N_9968,N_9890,N_9751);
nor U9969 (N_9969,N_9883,N_9754);
xnor U9970 (N_9970,N_9792,N_9889);
nor U9971 (N_9971,N_9788,N_9860);
xnor U9972 (N_9972,N_9815,N_9797);
or U9973 (N_9973,N_9787,N_9865);
nand U9974 (N_9974,N_9808,N_9831);
nand U9975 (N_9975,N_9792,N_9859);
or U9976 (N_9976,N_9839,N_9838);
and U9977 (N_9977,N_9824,N_9803);
nand U9978 (N_9978,N_9802,N_9760);
nand U9979 (N_9979,N_9879,N_9831);
or U9980 (N_9980,N_9777,N_9851);
or U9981 (N_9981,N_9875,N_9873);
nand U9982 (N_9982,N_9789,N_9771);
nor U9983 (N_9983,N_9855,N_9861);
nand U9984 (N_9984,N_9756,N_9839);
or U9985 (N_9985,N_9778,N_9853);
or U9986 (N_9986,N_9778,N_9754);
or U9987 (N_9987,N_9841,N_9805);
and U9988 (N_9988,N_9854,N_9760);
nand U9989 (N_9989,N_9880,N_9878);
xor U9990 (N_9990,N_9865,N_9877);
xor U9991 (N_9991,N_9825,N_9835);
nor U9992 (N_9992,N_9822,N_9789);
or U9993 (N_9993,N_9860,N_9874);
and U9994 (N_9994,N_9830,N_9822);
nand U9995 (N_9995,N_9891,N_9811);
nand U9996 (N_9996,N_9806,N_9796);
nor U9997 (N_9997,N_9768,N_9816);
and U9998 (N_9998,N_9794,N_9872);
nor U9999 (N_9999,N_9849,N_9810);
xnor U10000 (N_10000,N_9849,N_9830);
and U10001 (N_10001,N_9806,N_9772);
or U10002 (N_10002,N_9779,N_9776);
nand U10003 (N_10003,N_9757,N_9885);
nand U10004 (N_10004,N_9860,N_9802);
nor U10005 (N_10005,N_9895,N_9794);
nor U10006 (N_10006,N_9893,N_9898);
and U10007 (N_10007,N_9884,N_9808);
nand U10008 (N_10008,N_9806,N_9859);
and U10009 (N_10009,N_9764,N_9832);
and U10010 (N_10010,N_9820,N_9781);
or U10011 (N_10011,N_9889,N_9843);
and U10012 (N_10012,N_9831,N_9886);
or U10013 (N_10013,N_9803,N_9871);
and U10014 (N_10014,N_9810,N_9896);
or U10015 (N_10015,N_9885,N_9752);
or U10016 (N_10016,N_9854,N_9778);
and U10017 (N_10017,N_9787,N_9829);
nand U10018 (N_10018,N_9843,N_9800);
nor U10019 (N_10019,N_9888,N_9875);
nand U10020 (N_10020,N_9821,N_9780);
and U10021 (N_10021,N_9772,N_9878);
nor U10022 (N_10022,N_9836,N_9769);
and U10023 (N_10023,N_9774,N_9778);
nor U10024 (N_10024,N_9777,N_9817);
nor U10025 (N_10025,N_9795,N_9875);
or U10026 (N_10026,N_9898,N_9792);
nand U10027 (N_10027,N_9898,N_9763);
nand U10028 (N_10028,N_9774,N_9842);
nor U10029 (N_10029,N_9751,N_9808);
or U10030 (N_10030,N_9792,N_9833);
or U10031 (N_10031,N_9789,N_9786);
and U10032 (N_10032,N_9822,N_9824);
or U10033 (N_10033,N_9890,N_9757);
nor U10034 (N_10034,N_9811,N_9822);
and U10035 (N_10035,N_9773,N_9768);
and U10036 (N_10036,N_9815,N_9786);
and U10037 (N_10037,N_9814,N_9857);
nor U10038 (N_10038,N_9751,N_9883);
or U10039 (N_10039,N_9757,N_9860);
and U10040 (N_10040,N_9862,N_9775);
or U10041 (N_10041,N_9758,N_9888);
or U10042 (N_10042,N_9862,N_9895);
nand U10043 (N_10043,N_9851,N_9784);
nand U10044 (N_10044,N_9846,N_9799);
nand U10045 (N_10045,N_9870,N_9865);
or U10046 (N_10046,N_9784,N_9887);
or U10047 (N_10047,N_9794,N_9811);
nor U10048 (N_10048,N_9786,N_9816);
xnor U10049 (N_10049,N_9809,N_9861);
or U10050 (N_10050,N_9981,N_9909);
nand U10051 (N_10051,N_10030,N_10016);
nor U10052 (N_10052,N_9949,N_10004);
nor U10053 (N_10053,N_9941,N_9910);
xnor U10054 (N_10054,N_9914,N_9960);
nand U10055 (N_10055,N_10021,N_10013);
nor U10056 (N_10056,N_10038,N_10035);
xor U10057 (N_10057,N_10031,N_9952);
nor U10058 (N_10058,N_9931,N_9978);
or U10059 (N_10059,N_9933,N_9943);
or U10060 (N_10060,N_9995,N_9936);
and U10061 (N_10061,N_9962,N_9983);
and U10062 (N_10062,N_9975,N_10010);
nand U10063 (N_10063,N_10009,N_9902);
and U10064 (N_10064,N_10014,N_10028);
or U10065 (N_10065,N_9958,N_9935);
nand U10066 (N_10066,N_10007,N_9993);
or U10067 (N_10067,N_9950,N_9944);
nor U10068 (N_10068,N_9930,N_9969);
xor U10069 (N_10069,N_10047,N_9955);
nand U10070 (N_10070,N_9903,N_9977);
nor U10071 (N_10071,N_10005,N_9912);
nor U10072 (N_10072,N_10034,N_9982);
and U10073 (N_10073,N_9932,N_10033);
or U10074 (N_10074,N_9907,N_10037);
and U10075 (N_10075,N_9940,N_9919);
nor U10076 (N_10076,N_10036,N_9948);
nand U10077 (N_10077,N_9963,N_9946);
or U10078 (N_10078,N_9991,N_9921);
nor U10079 (N_10079,N_9968,N_9924);
nand U10080 (N_10080,N_9984,N_10048);
or U10081 (N_10081,N_9938,N_10024);
and U10082 (N_10082,N_9913,N_10006);
nand U10083 (N_10083,N_9945,N_10027);
nand U10084 (N_10084,N_10000,N_10043);
nand U10085 (N_10085,N_9937,N_10017);
nor U10086 (N_10086,N_9906,N_10039);
nand U10087 (N_10087,N_9961,N_9934);
and U10088 (N_10088,N_9997,N_9972);
xnor U10089 (N_10089,N_9953,N_10002);
nand U10090 (N_10090,N_10008,N_9918);
nand U10091 (N_10091,N_9979,N_9900);
xnor U10092 (N_10092,N_9967,N_10026);
nor U10093 (N_10093,N_9917,N_9956);
nand U10094 (N_10094,N_9999,N_9920);
nand U10095 (N_10095,N_10018,N_10049);
and U10096 (N_10096,N_9916,N_9951);
xnor U10097 (N_10097,N_10044,N_10032);
or U10098 (N_10098,N_10012,N_9922);
xor U10099 (N_10099,N_9971,N_9908);
xor U10100 (N_10100,N_10001,N_10020);
and U10101 (N_10101,N_9974,N_9947);
nor U10102 (N_10102,N_9973,N_10040);
nor U10103 (N_10103,N_9966,N_9915);
xnor U10104 (N_10104,N_9926,N_10045);
or U10105 (N_10105,N_10011,N_9987);
xor U10106 (N_10106,N_9986,N_9965);
and U10107 (N_10107,N_9998,N_10003);
nand U10108 (N_10108,N_9989,N_9990);
xor U10109 (N_10109,N_10022,N_9970);
or U10110 (N_10110,N_9923,N_9901);
or U10111 (N_10111,N_9976,N_9925);
nand U10112 (N_10112,N_10019,N_10029);
and U10113 (N_10113,N_9904,N_9957);
xor U10114 (N_10114,N_9994,N_9980);
nand U10115 (N_10115,N_10015,N_9954);
and U10116 (N_10116,N_10025,N_9996);
or U10117 (N_10117,N_9964,N_9905);
nor U10118 (N_10118,N_9927,N_10042);
and U10119 (N_10119,N_9985,N_9988);
nand U10120 (N_10120,N_10023,N_9929);
xnor U10121 (N_10121,N_9942,N_10041);
nand U10122 (N_10122,N_10046,N_9992);
xnor U10123 (N_10123,N_9911,N_9959);
nand U10124 (N_10124,N_9928,N_9939);
and U10125 (N_10125,N_10039,N_9946);
and U10126 (N_10126,N_10049,N_9943);
and U10127 (N_10127,N_10048,N_10044);
nor U10128 (N_10128,N_9905,N_10020);
xor U10129 (N_10129,N_9952,N_10042);
and U10130 (N_10130,N_9948,N_9918);
or U10131 (N_10131,N_10027,N_9910);
xor U10132 (N_10132,N_9915,N_10010);
nor U10133 (N_10133,N_9948,N_10041);
nor U10134 (N_10134,N_10016,N_10029);
nand U10135 (N_10135,N_9919,N_10012);
nand U10136 (N_10136,N_9965,N_10046);
and U10137 (N_10137,N_10012,N_9911);
or U10138 (N_10138,N_9998,N_10045);
or U10139 (N_10139,N_9964,N_9931);
and U10140 (N_10140,N_10028,N_9914);
or U10141 (N_10141,N_9957,N_10027);
nand U10142 (N_10142,N_10035,N_9958);
nor U10143 (N_10143,N_9923,N_10038);
and U10144 (N_10144,N_10047,N_9944);
nand U10145 (N_10145,N_9922,N_9917);
nor U10146 (N_10146,N_9964,N_9965);
nor U10147 (N_10147,N_10014,N_9988);
and U10148 (N_10148,N_9946,N_9942);
nor U10149 (N_10149,N_9938,N_9947);
xor U10150 (N_10150,N_9906,N_9938);
xor U10151 (N_10151,N_9972,N_9936);
and U10152 (N_10152,N_10035,N_9988);
or U10153 (N_10153,N_9953,N_9905);
nor U10154 (N_10154,N_10043,N_10013);
nand U10155 (N_10155,N_9977,N_9908);
or U10156 (N_10156,N_10011,N_9954);
xnor U10157 (N_10157,N_10027,N_10016);
xor U10158 (N_10158,N_10028,N_10003);
and U10159 (N_10159,N_10046,N_9995);
nor U10160 (N_10160,N_9997,N_9918);
or U10161 (N_10161,N_10010,N_9941);
nor U10162 (N_10162,N_9937,N_9939);
and U10163 (N_10163,N_9957,N_9968);
nand U10164 (N_10164,N_9901,N_9939);
nand U10165 (N_10165,N_9926,N_9905);
or U10166 (N_10166,N_9992,N_9997);
nor U10167 (N_10167,N_10032,N_10037);
or U10168 (N_10168,N_9948,N_9909);
or U10169 (N_10169,N_10005,N_9999);
nor U10170 (N_10170,N_9999,N_9987);
nor U10171 (N_10171,N_10036,N_9952);
and U10172 (N_10172,N_9905,N_9916);
or U10173 (N_10173,N_9918,N_10046);
or U10174 (N_10174,N_9906,N_10025);
or U10175 (N_10175,N_9993,N_9907);
or U10176 (N_10176,N_9928,N_10034);
nor U10177 (N_10177,N_10023,N_9950);
nor U10178 (N_10178,N_10047,N_10003);
nand U10179 (N_10179,N_9937,N_9922);
xor U10180 (N_10180,N_9987,N_9988);
nor U10181 (N_10181,N_9956,N_9909);
nor U10182 (N_10182,N_9908,N_9962);
nand U10183 (N_10183,N_9964,N_9977);
nor U10184 (N_10184,N_10021,N_10004);
or U10185 (N_10185,N_10041,N_9983);
nor U10186 (N_10186,N_10029,N_9906);
nand U10187 (N_10187,N_10029,N_9914);
or U10188 (N_10188,N_9901,N_9942);
or U10189 (N_10189,N_10019,N_10021);
and U10190 (N_10190,N_9980,N_9971);
or U10191 (N_10191,N_9986,N_9974);
nor U10192 (N_10192,N_9996,N_9927);
or U10193 (N_10193,N_10027,N_10039);
nor U10194 (N_10194,N_10018,N_10045);
nand U10195 (N_10195,N_10048,N_9902);
and U10196 (N_10196,N_9985,N_9953);
or U10197 (N_10197,N_10004,N_9990);
and U10198 (N_10198,N_10009,N_9977);
and U10199 (N_10199,N_10002,N_10039);
nand U10200 (N_10200,N_10070,N_10083);
nand U10201 (N_10201,N_10073,N_10059);
nor U10202 (N_10202,N_10075,N_10187);
or U10203 (N_10203,N_10117,N_10142);
nand U10204 (N_10204,N_10094,N_10110);
xor U10205 (N_10205,N_10179,N_10111);
nor U10206 (N_10206,N_10149,N_10182);
or U10207 (N_10207,N_10162,N_10056);
and U10208 (N_10208,N_10119,N_10128);
nor U10209 (N_10209,N_10052,N_10164);
or U10210 (N_10210,N_10170,N_10064);
or U10211 (N_10211,N_10141,N_10125);
nand U10212 (N_10212,N_10077,N_10091);
nand U10213 (N_10213,N_10101,N_10103);
nand U10214 (N_10214,N_10107,N_10197);
and U10215 (N_10215,N_10175,N_10113);
nand U10216 (N_10216,N_10112,N_10050);
or U10217 (N_10217,N_10198,N_10134);
and U10218 (N_10218,N_10192,N_10074);
or U10219 (N_10219,N_10068,N_10086);
and U10220 (N_10220,N_10138,N_10136);
nor U10221 (N_10221,N_10131,N_10140);
nand U10222 (N_10222,N_10153,N_10060);
or U10223 (N_10223,N_10079,N_10161);
nand U10224 (N_10224,N_10171,N_10058);
or U10225 (N_10225,N_10055,N_10122);
or U10226 (N_10226,N_10051,N_10148);
and U10227 (N_10227,N_10053,N_10114);
nand U10228 (N_10228,N_10116,N_10144);
or U10229 (N_10229,N_10196,N_10145);
nand U10230 (N_10230,N_10098,N_10143);
and U10231 (N_10231,N_10106,N_10199);
or U10232 (N_10232,N_10066,N_10062);
nand U10233 (N_10233,N_10087,N_10186);
and U10234 (N_10234,N_10129,N_10155);
or U10235 (N_10235,N_10159,N_10193);
xnor U10236 (N_10236,N_10160,N_10067);
and U10237 (N_10237,N_10096,N_10154);
nand U10238 (N_10238,N_10105,N_10169);
xor U10239 (N_10239,N_10071,N_10081);
nand U10240 (N_10240,N_10057,N_10184);
nor U10241 (N_10241,N_10183,N_10178);
or U10242 (N_10242,N_10167,N_10089);
nand U10243 (N_10243,N_10185,N_10172);
nand U10244 (N_10244,N_10092,N_10102);
nor U10245 (N_10245,N_10133,N_10100);
and U10246 (N_10246,N_10189,N_10166);
xnor U10247 (N_10247,N_10115,N_10135);
and U10248 (N_10248,N_10176,N_10191);
xnor U10249 (N_10249,N_10181,N_10084);
nand U10250 (N_10250,N_10093,N_10146);
or U10251 (N_10251,N_10082,N_10099);
and U10252 (N_10252,N_10118,N_10151);
nor U10253 (N_10253,N_10127,N_10139);
nand U10254 (N_10254,N_10108,N_10095);
and U10255 (N_10255,N_10085,N_10180);
nand U10256 (N_10256,N_10150,N_10195);
xor U10257 (N_10257,N_10088,N_10120);
and U10258 (N_10258,N_10168,N_10076);
or U10259 (N_10259,N_10163,N_10156);
and U10260 (N_10260,N_10124,N_10104);
or U10261 (N_10261,N_10069,N_10061);
and U10262 (N_10262,N_10174,N_10188);
nand U10263 (N_10263,N_10063,N_10165);
or U10264 (N_10264,N_10097,N_10152);
or U10265 (N_10265,N_10137,N_10173);
and U10266 (N_10266,N_10121,N_10147);
nor U10267 (N_10267,N_10072,N_10190);
and U10268 (N_10268,N_10054,N_10109);
nand U10269 (N_10269,N_10177,N_10157);
nand U10270 (N_10270,N_10132,N_10078);
nor U10271 (N_10271,N_10130,N_10065);
and U10272 (N_10272,N_10090,N_10126);
nand U10273 (N_10273,N_10123,N_10080);
or U10274 (N_10274,N_10158,N_10194);
nand U10275 (N_10275,N_10167,N_10084);
or U10276 (N_10276,N_10098,N_10090);
nor U10277 (N_10277,N_10071,N_10104);
nand U10278 (N_10278,N_10076,N_10093);
or U10279 (N_10279,N_10090,N_10196);
nand U10280 (N_10280,N_10167,N_10118);
and U10281 (N_10281,N_10131,N_10168);
xor U10282 (N_10282,N_10109,N_10076);
nand U10283 (N_10283,N_10173,N_10135);
or U10284 (N_10284,N_10075,N_10157);
nor U10285 (N_10285,N_10191,N_10084);
and U10286 (N_10286,N_10166,N_10056);
or U10287 (N_10287,N_10141,N_10139);
and U10288 (N_10288,N_10102,N_10063);
nand U10289 (N_10289,N_10186,N_10136);
or U10290 (N_10290,N_10125,N_10198);
and U10291 (N_10291,N_10162,N_10132);
nand U10292 (N_10292,N_10108,N_10106);
nor U10293 (N_10293,N_10149,N_10191);
nand U10294 (N_10294,N_10163,N_10070);
nand U10295 (N_10295,N_10167,N_10105);
and U10296 (N_10296,N_10114,N_10156);
xnor U10297 (N_10297,N_10131,N_10155);
nor U10298 (N_10298,N_10183,N_10166);
nor U10299 (N_10299,N_10160,N_10091);
nand U10300 (N_10300,N_10056,N_10084);
nand U10301 (N_10301,N_10058,N_10090);
xor U10302 (N_10302,N_10169,N_10152);
or U10303 (N_10303,N_10194,N_10058);
and U10304 (N_10304,N_10126,N_10144);
xnor U10305 (N_10305,N_10158,N_10117);
and U10306 (N_10306,N_10085,N_10112);
nor U10307 (N_10307,N_10157,N_10102);
and U10308 (N_10308,N_10063,N_10179);
and U10309 (N_10309,N_10134,N_10072);
or U10310 (N_10310,N_10199,N_10051);
or U10311 (N_10311,N_10055,N_10058);
nor U10312 (N_10312,N_10095,N_10152);
xor U10313 (N_10313,N_10171,N_10130);
nand U10314 (N_10314,N_10101,N_10130);
and U10315 (N_10315,N_10060,N_10179);
nor U10316 (N_10316,N_10190,N_10182);
nand U10317 (N_10317,N_10050,N_10117);
and U10318 (N_10318,N_10116,N_10170);
nand U10319 (N_10319,N_10186,N_10091);
or U10320 (N_10320,N_10097,N_10158);
and U10321 (N_10321,N_10097,N_10127);
and U10322 (N_10322,N_10193,N_10186);
nand U10323 (N_10323,N_10054,N_10095);
nand U10324 (N_10324,N_10100,N_10128);
xnor U10325 (N_10325,N_10054,N_10057);
nor U10326 (N_10326,N_10099,N_10110);
nor U10327 (N_10327,N_10082,N_10108);
xnor U10328 (N_10328,N_10105,N_10082);
nor U10329 (N_10329,N_10105,N_10178);
or U10330 (N_10330,N_10066,N_10090);
nand U10331 (N_10331,N_10178,N_10134);
nand U10332 (N_10332,N_10081,N_10136);
nand U10333 (N_10333,N_10101,N_10153);
and U10334 (N_10334,N_10104,N_10093);
nor U10335 (N_10335,N_10078,N_10136);
and U10336 (N_10336,N_10163,N_10077);
nor U10337 (N_10337,N_10075,N_10104);
and U10338 (N_10338,N_10059,N_10136);
or U10339 (N_10339,N_10087,N_10170);
or U10340 (N_10340,N_10176,N_10172);
nor U10341 (N_10341,N_10117,N_10061);
nor U10342 (N_10342,N_10131,N_10072);
and U10343 (N_10343,N_10190,N_10152);
and U10344 (N_10344,N_10093,N_10169);
xnor U10345 (N_10345,N_10195,N_10123);
nand U10346 (N_10346,N_10136,N_10128);
or U10347 (N_10347,N_10182,N_10107);
nor U10348 (N_10348,N_10197,N_10137);
or U10349 (N_10349,N_10181,N_10138);
nor U10350 (N_10350,N_10234,N_10270);
and U10351 (N_10351,N_10317,N_10244);
and U10352 (N_10352,N_10273,N_10274);
or U10353 (N_10353,N_10211,N_10329);
and U10354 (N_10354,N_10291,N_10207);
and U10355 (N_10355,N_10213,N_10216);
nor U10356 (N_10356,N_10280,N_10328);
and U10357 (N_10357,N_10265,N_10271);
and U10358 (N_10358,N_10325,N_10278);
or U10359 (N_10359,N_10228,N_10302);
nor U10360 (N_10360,N_10266,N_10248);
and U10361 (N_10361,N_10263,N_10305);
nor U10362 (N_10362,N_10323,N_10322);
nor U10363 (N_10363,N_10343,N_10240);
nor U10364 (N_10364,N_10230,N_10320);
and U10365 (N_10365,N_10254,N_10201);
xnor U10366 (N_10366,N_10236,N_10324);
nand U10367 (N_10367,N_10326,N_10275);
nand U10368 (N_10368,N_10233,N_10268);
nand U10369 (N_10369,N_10225,N_10344);
nor U10370 (N_10370,N_10311,N_10220);
nand U10371 (N_10371,N_10241,N_10331);
and U10372 (N_10372,N_10229,N_10321);
xnor U10373 (N_10373,N_10204,N_10214);
or U10374 (N_10374,N_10261,N_10307);
or U10375 (N_10375,N_10330,N_10243);
nor U10376 (N_10376,N_10259,N_10277);
xnor U10377 (N_10377,N_10242,N_10289);
nand U10378 (N_10378,N_10205,N_10287);
and U10379 (N_10379,N_10202,N_10250);
nor U10380 (N_10380,N_10253,N_10313);
nor U10381 (N_10381,N_10338,N_10296);
xor U10382 (N_10382,N_10292,N_10286);
nor U10383 (N_10383,N_10224,N_10319);
or U10384 (N_10384,N_10279,N_10310);
and U10385 (N_10385,N_10297,N_10221);
and U10386 (N_10386,N_10298,N_10203);
nand U10387 (N_10387,N_10212,N_10312);
nor U10388 (N_10388,N_10249,N_10341);
and U10389 (N_10389,N_10335,N_10276);
nor U10390 (N_10390,N_10314,N_10300);
or U10391 (N_10391,N_10219,N_10245);
and U10392 (N_10392,N_10327,N_10258);
and U10393 (N_10393,N_10215,N_10227);
and U10394 (N_10394,N_10304,N_10255);
xor U10395 (N_10395,N_10235,N_10200);
or U10396 (N_10396,N_10299,N_10301);
nand U10397 (N_10397,N_10262,N_10348);
nand U10398 (N_10398,N_10308,N_10247);
nor U10399 (N_10399,N_10251,N_10246);
nand U10400 (N_10400,N_10285,N_10269);
and U10401 (N_10401,N_10282,N_10309);
nor U10402 (N_10402,N_10222,N_10206);
or U10403 (N_10403,N_10272,N_10303);
nor U10404 (N_10404,N_10256,N_10267);
or U10405 (N_10405,N_10232,N_10257);
xor U10406 (N_10406,N_10226,N_10264);
nor U10407 (N_10407,N_10333,N_10208);
xor U10408 (N_10408,N_10239,N_10345);
and U10409 (N_10409,N_10342,N_10293);
or U10410 (N_10410,N_10281,N_10209);
or U10411 (N_10411,N_10218,N_10290);
and U10412 (N_10412,N_10237,N_10223);
and U10413 (N_10413,N_10217,N_10315);
xor U10414 (N_10414,N_10346,N_10306);
or U10415 (N_10415,N_10336,N_10337);
nor U10416 (N_10416,N_10332,N_10340);
nand U10417 (N_10417,N_10339,N_10349);
xnor U10418 (N_10418,N_10252,N_10210);
xor U10419 (N_10419,N_10295,N_10283);
nor U10420 (N_10420,N_10260,N_10288);
nand U10421 (N_10421,N_10318,N_10316);
nand U10422 (N_10422,N_10294,N_10231);
and U10423 (N_10423,N_10238,N_10334);
and U10424 (N_10424,N_10284,N_10347);
nand U10425 (N_10425,N_10207,N_10223);
or U10426 (N_10426,N_10327,N_10308);
or U10427 (N_10427,N_10202,N_10333);
or U10428 (N_10428,N_10309,N_10319);
and U10429 (N_10429,N_10321,N_10314);
or U10430 (N_10430,N_10234,N_10315);
and U10431 (N_10431,N_10320,N_10308);
nor U10432 (N_10432,N_10337,N_10279);
nand U10433 (N_10433,N_10209,N_10274);
nand U10434 (N_10434,N_10214,N_10220);
nor U10435 (N_10435,N_10244,N_10230);
nand U10436 (N_10436,N_10201,N_10348);
and U10437 (N_10437,N_10290,N_10225);
nor U10438 (N_10438,N_10311,N_10309);
and U10439 (N_10439,N_10250,N_10305);
or U10440 (N_10440,N_10204,N_10318);
or U10441 (N_10441,N_10277,N_10256);
and U10442 (N_10442,N_10304,N_10336);
and U10443 (N_10443,N_10280,N_10254);
or U10444 (N_10444,N_10316,N_10275);
nand U10445 (N_10445,N_10254,N_10342);
nor U10446 (N_10446,N_10305,N_10346);
or U10447 (N_10447,N_10242,N_10237);
nand U10448 (N_10448,N_10324,N_10274);
nand U10449 (N_10449,N_10307,N_10252);
nand U10450 (N_10450,N_10295,N_10217);
and U10451 (N_10451,N_10277,N_10226);
nor U10452 (N_10452,N_10265,N_10316);
nand U10453 (N_10453,N_10311,N_10214);
nor U10454 (N_10454,N_10210,N_10218);
nor U10455 (N_10455,N_10211,N_10200);
nand U10456 (N_10456,N_10294,N_10206);
nand U10457 (N_10457,N_10266,N_10337);
or U10458 (N_10458,N_10226,N_10305);
nand U10459 (N_10459,N_10263,N_10294);
or U10460 (N_10460,N_10214,N_10211);
nand U10461 (N_10461,N_10204,N_10332);
nand U10462 (N_10462,N_10283,N_10241);
nor U10463 (N_10463,N_10234,N_10219);
xnor U10464 (N_10464,N_10260,N_10304);
xor U10465 (N_10465,N_10341,N_10280);
nor U10466 (N_10466,N_10272,N_10281);
or U10467 (N_10467,N_10267,N_10305);
nand U10468 (N_10468,N_10249,N_10331);
nor U10469 (N_10469,N_10280,N_10309);
or U10470 (N_10470,N_10312,N_10223);
xor U10471 (N_10471,N_10236,N_10334);
xor U10472 (N_10472,N_10212,N_10255);
xor U10473 (N_10473,N_10264,N_10330);
xnor U10474 (N_10474,N_10243,N_10308);
xor U10475 (N_10475,N_10318,N_10206);
and U10476 (N_10476,N_10236,N_10252);
and U10477 (N_10477,N_10296,N_10310);
or U10478 (N_10478,N_10329,N_10348);
or U10479 (N_10479,N_10208,N_10244);
nor U10480 (N_10480,N_10317,N_10201);
xnor U10481 (N_10481,N_10299,N_10326);
nand U10482 (N_10482,N_10349,N_10256);
or U10483 (N_10483,N_10281,N_10200);
nand U10484 (N_10484,N_10307,N_10227);
nand U10485 (N_10485,N_10297,N_10256);
or U10486 (N_10486,N_10313,N_10300);
nand U10487 (N_10487,N_10214,N_10317);
or U10488 (N_10488,N_10250,N_10336);
nor U10489 (N_10489,N_10345,N_10268);
and U10490 (N_10490,N_10296,N_10203);
nor U10491 (N_10491,N_10227,N_10318);
and U10492 (N_10492,N_10238,N_10317);
nor U10493 (N_10493,N_10306,N_10308);
xnor U10494 (N_10494,N_10290,N_10211);
xnor U10495 (N_10495,N_10239,N_10214);
or U10496 (N_10496,N_10313,N_10273);
nor U10497 (N_10497,N_10310,N_10328);
or U10498 (N_10498,N_10341,N_10235);
nor U10499 (N_10499,N_10329,N_10324);
nand U10500 (N_10500,N_10469,N_10384);
or U10501 (N_10501,N_10454,N_10370);
or U10502 (N_10502,N_10411,N_10453);
or U10503 (N_10503,N_10375,N_10423);
nor U10504 (N_10504,N_10353,N_10473);
or U10505 (N_10505,N_10461,N_10394);
or U10506 (N_10506,N_10464,N_10468);
xor U10507 (N_10507,N_10399,N_10412);
and U10508 (N_10508,N_10465,N_10404);
nor U10509 (N_10509,N_10463,N_10455);
nand U10510 (N_10510,N_10421,N_10418);
xor U10511 (N_10511,N_10407,N_10396);
and U10512 (N_10512,N_10400,N_10380);
nand U10513 (N_10513,N_10441,N_10382);
nor U10514 (N_10514,N_10378,N_10403);
nand U10515 (N_10515,N_10471,N_10478);
nor U10516 (N_10516,N_10429,N_10359);
nand U10517 (N_10517,N_10446,N_10477);
nand U10518 (N_10518,N_10430,N_10458);
and U10519 (N_10519,N_10467,N_10460);
nor U10520 (N_10520,N_10437,N_10493);
nand U10521 (N_10521,N_10443,N_10427);
or U10522 (N_10522,N_10413,N_10406);
nor U10523 (N_10523,N_10442,N_10414);
or U10524 (N_10524,N_10475,N_10439);
or U10525 (N_10525,N_10432,N_10474);
xor U10526 (N_10526,N_10386,N_10367);
nand U10527 (N_10527,N_10393,N_10425);
and U10528 (N_10528,N_10426,N_10420);
nand U10529 (N_10529,N_10488,N_10452);
or U10530 (N_10530,N_10436,N_10440);
nand U10531 (N_10531,N_10497,N_10369);
and U10532 (N_10532,N_10405,N_10409);
nor U10533 (N_10533,N_10438,N_10434);
or U10534 (N_10534,N_10444,N_10358);
and U10535 (N_10535,N_10388,N_10466);
or U10536 (N_10536,N_10355,N_10486);
and U10537 (N_10537,N_10435,N_10456);
or U10538 (N_10538,N_10374,N_10415);
nand U10539 (N_10539,N_10451,N_10470);
nand U10540 (N_10540,N_10422,N_10416);
or U10541 (N_10541,N_10499,N_10419);
xnor U10542 (N_10542,N_10480,N_10498);
nand U10543 (N_10543,N_10387,N_10401);
nand U10544 (N_10544,N_10372,N_10494);
and U10545 (N_10545,N_10483,N_10350);
xnor U10546 (N_10546,N_10364,N_10377);
xor U10547 (N_10547,N_10357,N_10495);
or U10548 (N_10548,N_10491,N_10365);
and U10549 (N_10549,N_10360,N_10356);
and U10550 (N_10550,N_10389,N_10424);
nor U10551 (N_10551,N_10433,N_10381);
nand U10552 (N_10552,N_10479,N_10361);
and U10553 (N_10553,N_10371,N_10410);
and U10554 (N_10554,N_10395,N_10391);
nor U10555 (N_10555,N_10481,N_10408);
nor U10556 (N_10556,N_10390,N_10448);
nor U10557 (N_10557,N_10449,N_10368);
nor U10558 (N_10558,N_10417,N_10431);
xor U10559 (N_10559,N_10476,N_10402);
nor U10560 (N_10560,N_10482,N_10459);
or U10561 (N_10561,N_10366,N_10445);
and U10562 (N_10562,N_10485,N_10379);
or U10563 (N_10563,N_10397,N_10484);
and U10564 (N_10564,N_10472,N_10487);
or U10565 (N_10565,N_10450,N_10354);
xor U10566 (N_10566,N_10383,N_10457);
nand U10567 (N_10567,N_10362,N_10492);
xnor U10568 (N_10568,N_10398,N_10376);
nand U10569 (N_10569,N_10490,N_10462);
or U10570 (N_10570,N_10373,N_10363);
or U10571 (N_10571,N_10352,N_10489);
and U10572 (N_10572,N_10496,N_10385);
nor U10573 (N_10573,N_10447,N_10428);
and U10574 (N_10574,N_10351,N_10392);
nor U10575 (N_10575,N_10442,N_10457);
and U10576 (N_10576,N_10354,N_10381);
nand U10577 (N_10577,N_10444,N_10357);
nand U10578 (N_10578,N_10459,N_10373);
and U10579 (N_10579,N_10488,N_10497);
and U10580 (N_10580,N_10481,N_10459);
nand U10581 (N_10581,N_10388,N_10389);
nor U10582 (N_10582,N_10397,N_10452);
nand U10583 (N_10583,N_10468,N_10498);
nand U10584 (N_10584,N_10386,N_10424);
xnor U10585 (N_10585,N_10390,N_10466);
or U10586 (N_10586,N_10485,N_10391);
nor U10587 (N_10587,N_10405,N_10374);
or U10588 (N_10588,N_10377,N_10389);
and U10589 (N_10589,N_10382,N_10358);
nand U10590 (N_10590,N_10382,N_10356);
or U10591 (N_10591,N_10412,N_10493);
nor U10592 (N_10592,N_10394,N_10400);
nor U10593 (N_10593,N_10476,N_10375);
or U10594 (N_10594,N_10473,N_10411);
nor U10595 (N_10595,N_10422,N_10426);
or U10596 (N_10596,N_10371,N_10489);
nand U10597 (N_10597,N_10401,N_10402);
nand U10598 (N_10598,N_10459,N_10375);
nand U10599 (N_10599,N_10460,N_10480);
and U10600 (N_10600,N_10476,N_10474);
or U10601 (N_10601,N_10353,N_10402);
nor U10602 (N_10602,N_10429,N_10449);
xor U10603 (N_10603,N_10379,N_10398);
and U10604 (N_10604,N_10451,N_10364);
nand U10605 (N_10605,N_10453,N_10437);
nor U10606 (N_10606,N_10388,N_10414);
and U10607 (N_10607,N_10351,N_10459);
xnor U10608 (N_10608,N_10377,N_10466);
and U10609 (N_10609,N_10360,N_10440);
and U10610 (N_10610,N_10499,N_10482);
or U10611 (N_10611,N_10481,N_10360);
and U10612 (N_10612,N_10488,N_10447);
nand U10613 (N_10613,N_10434,N_10427);
and U10614 (N_10614,N_10473,N_10426);
nand U10615 (N_10615,N_10414,N_10372);
xor U10616 (N_10616,N_10371,N_10480);
nand U10617 (N_10617,N_10350,N_10395);
and U10618 (N_10618,N_10398,N_10438);
xor U10619 (N_10619,N_10441,N_10384);
and U10620 (N_10620,N_10415,N_10409);
or U10621 (N_10621,N_10371,N_10458);
nand U10622 (N_10622,N_10490,N_10379);
and U10623 (N_10623,N_10379,N_10388);
xnor U10624 (N_10624,N_10413,N_10394);
or U10625 (N_10625,N_10391,N_10475);
nor U10626 (N_10626,N_10450,N_10463);
nor U10627 (N_10627,N_10460,N_10499);
and U10628 (N_10628,N_10472,N_10362);
nor U10629 (N_10629,N_10383,N_10432);
and U10630 (N_10630,N_10478,N_10418);
nand U10631 (N_10631,N_10391,N_10384);
and U10632 (N_10632,N_10355,N_10462);
or U10633 (N_10633,N_10476,N_10458);
and U10634 (N_10634,N_10422,N_10419);
nor U10635 (N_10635,N_10365,N_10441);
nor U10636 (N_10636,N_10380,N_10482);
nand U10637 (N_10637,N_10381,N_10439);
nor U10638 (N_10638,N_10371,N_10375);
nor U10639 (N_10639,N_10458,N_10422);
and U10640 (N_10640,N_10418,N_10432);
and U10641 (N_10641,N_10479,N_10358);
or U10642 (N_10642,N_10436,N_10361);
xor U10643 (N_10643,N_10376,N_10409);
nand U10644 (N_10644,N_10428,N_10408);
nand U10645 (N_10645,N_10351,N_10476);
or U10646 (N_10646,N_10444,N_10429);
nor U10647 (N_10647,N_10401,N_10366);
or U10648 (N_10648,N_10364,N_10471);
or U10649 (N_10649,N_10450,N_10446);
nand U10650 (N_10650,N_10596,N_10581);
and U10651 (N_10651,N_10521,N_10588);
nor U10652 (N_10652,N_10515,N_10540);
or U10653 (N_10653,N_10511,N_10523);
nand U10654 (N_10654,N_10535,N_10612);
or U10655 (N_10655,N_10551,N_10560);
nor U10656 (N_10656,N_10624,N_10520);
nor U10657 (N_10657,N_10580,N_10620);
and U10658 (N_10658,N_10538,N_10573);
nor U10659 (N_10659,N_10626,N_10501);
or U10660 (N_10660,N_10608,N_10539);
and U10661 (N_10661,N_10570,N_10512);
nor U10662 (N_10662,N_10563,N_10643);
nand U10663 (N_10663,N_10500,N_10553);
xor U10664 (N_10664,N_10633,N_10647);
or U10665 (N_10665,N_10627,N_10630);
or U10666 (N_10666,N_10556,N_10602);
or U10667 (N_10667,N_10531,N_10513);
nand U10668 (N_10668,N_10532,N_10536);
nand U10669 (N_10669,N_10530,N_10587);
or U10670 (N_10670,N_10564,N_10571);
nor U10671 (N_10671,N_10591,N_10507);
or U10672 (N_10672,N_10611,N_10613);
or U10673 (N_10673,N_10640,N_10557);
or U10674 (N_10674,N_10518,N_10522);
nor U10675 (N_10675,N_10648,N_10610);
nand U10676 (N_10676,N_10555,N_10582);
and U10677 (N_10677,N_10514,N_10525);
nand U10678 (N_10678,N_10604,N_10504);
or U10679 (N_10679,N_10508,N_10642);
or U10680 (N_10680,N_10519,N_10615);
or U10681 (N_10681,N_10609,N_10529);
nand U10682 (N_10682,N_10565,N_10569);
and U10683 (N_10683,N_10649,N_10509);
nand U10684 (N_10684,N_10619,N_10592);
or U10685 (N_10685,N_10506,N_10502);
and U10686 (N_10686,N_10550,N_10574);
and U10687 (N_10687,N_10632,N_10549);
and U10688 (N_10688,N_10637,N_10623);
xnor U10689 (N_10689,N_10526,N_10607);
or U10690 (N_10690,N_10566,N_10552);
nor U10691 (N_10691,N_10554,N_10543);
and U10692 (N_10692,N_10503,N_10598);
or U10693 (N_10693,N_10559,N_10562);
nor U10694 (N_10694,N_10614,N_10644);
xnor U10695 (N_10695,N_10597,N_10638);
nand U10696 (N_10696,N_10516,N_10586);
xnor U10697 (N_10697,N_10622,N_10544);
nor U10698 (N_10698,N_10528,N_10594);
or U10699 (N_10699,N_10629,N_10534);
and U10700 (N_10700,N_10567,N_10517);
nand U10701 (N_10701,N_10618,N_10524);
or U10702 (N_10702,N_10546,N_10616);
nand U10703 (N_10703,N_10601,N_10595);
or U10704 (N_10704,N_10641,N_10537);
or U10705 (N_10705,N_10636,N_10631);
and U10706 (N_10706,N_10645,N_10589);
or U10707 (N_10707,N_10576,N_10579);
and U10708 (N_10708,N_10599,N_10606);
nand U10709 (N_10709,N_10605,N_10600);
nor U10710 (N_10710,N_10583,N_10510);
nand U10711 (N_10711,N_10527,N_10561);
and U10712 (N_10712,N_10628,N_10646);
nand U10713 (N_10713,N_10568,N_10558);
nand U10714 (N_10714,N_10533,N_10578);
nor U10715 (N_10715,N_10541,N_10572);
nand U10716 (N_10716,N_10547,N_10545);
nand U10717 (N_10717,N_10639,N_10585);
or U10718 (N_10718,N_10577,N_10593);
and U10719 (N_10719,N_10548,N_10617);
nand U10720 (N_10720,N_10542,N_10603);
nor U10721 (N_10721,N_10621,N_10635);
and U10722 (N_10722,N_10575,N_10590);
nand U10723 (N_10723,N_10584,N_10634);
xnor U10724 (N_10724,N_10625,N_10505);
nor U10725 (N_10725,N_10512,N_10504);
nand U10726 (N_10726,N_10630,N_10529);
or U10727 (N_10727,N_10635,N_10574);
nand U10728 (N_10728,N_10590,N_10517);
nor U10729 (N_10729,N_10574,N_10554);
or U10730 (N_10730,N_10614,N_10508);
nand U10731 (N_10731,N_10561,N_10551);
and U10732 (N_10732,N_10603,N_10590);
nand U10733 (N_10733,N_10599,N_10580);
and U10734 (N_10734,N_10621,N_10586);
or U10735 (N_10735,N_10503,N_10560);
and U10736 (N_10736,N_10642,N_10529);
nor U10737 (N_10737,N_10646,N_10556);
nand U10738 (N_10738,N_10572,N_10620);
xnor U10739 (N_10739,N_10524,N_10582);
nor U10740 (N_10740,N_10549,N_10630);
and U10741 (N_10741,N_10626,N_10540);
and U10742 (N_10742,N_10563,N_10541);
nand U10743 (N_10743,N_10534,N_10539);
nor U10744 (N_10744,N_10596,N_10544);
nor U10745 (N_10745,N_10615,N_10530);
nand U10746 (N_10746,N_10555,N_10512);
nor U10747 (N_10747,N_10549,N_10589);
nand U10748 (N_10748,N_10638,N_10548);
or U10749 (N_10749,N_10505,N_10610);
and U10750 (N_10750,N_10601,N_10517);
nand U10751 (N_10751,N_10539,N_10573);
or U10752 (N_10752,N_10618,N_10511);
xnor U10753 (N_10753,N_10641,N_10560);
or U10754 (N_10754,N_10596,N_10585);
nand U10755 (N_10755,N_10630,N_10530);
xor U10756 (N_10756,N_10623,N_10507);
nor U10757 (N_10757,N_10519,N_10607);
and U10758 (N_10758,N_10612,N_10585);
and U10759 (N_10759,N_10607,N_10532);
nand U10760 (N_10760,N_10587,N_10580);
and U10761 (N_10761,N_10538,N_10608);
xor U10762 (N_10762,N_10568,N_10641);
nor U10763 (N_10763,N_10609,N_10518);
nand U10764 (N_10764,N_10508,N_10515);
xnor U10765 (N_10765,N_10563,N_10584);
nand U10766 (N_10766,N_10541,N_10624);
and U10767 (N_10767,N_10565,N_10514);
or U10768 (N_10768,N_10500,N_10635);
or U10769 (N_10769,N_10582,N_10588);
nor U10770 (N_10770,N_10646,N_10627);
xnor U10771 (N_10771,N_10575,N_10505);
nand U10772 (N_10772,N_10505,N_10595);
and U10773 (N_10773,N_10591,N_10598);
nand U10774 (N_10774,N_10545,N_10519);
xnor U10775 (N_10775,N_10598,N_10524);
and U10776 (N_10776,N_10556,N_10616);
or U10777 (N_10777,N_10635,N_10600);
and U10778 (N_10778,N_10545,N_10617);
nor U10779 (N_10779,N_10562,N_10584);
nand U10780 (N_10780,N_10582,N_10546);
nor U10781 (N_10781,N_10639,N_10597);
or U10782 (N_10782,N_10579,N_10563);
nand U10783 (N_10783,N_10585,N_10617);
and U10784 (N_10784,N_10508,N_10552);
and U10785 (N_10785,N_10587,N_10630);
or U10786 (N_10786,N_10589,N_10540);
nor U10787 (N_10787,N_10554,N_10562);
nand U10788 (N_10788,N_10541,N_10569);
and U10789 (N_10789,N_10646,N_10584);
and U10790 (N_10790,N_10506,N_10516);
and U10791 (N_10791,N_10616,N_10628);
nor U10792 (N_10792,N_10638,N_10620);
and U10793 (N_10793,N_10641,N_10592);
nor U10794 (N_10794,N_10622,N_10555);
nor U10795 (N_10795,N_10538,N_10588);
or U10796 (N_10796,N_10641,N_10580);
nand U10797 (N_10797,N_10534,N_10573);
or U10798 (N_10798,N_10572,N_10517);
and U10799 (N_10799,N_10521,N_10624);
nor U10800 (N_10800,N_10664,N_10759);
xnor U10801 (N_10801,N_10685,N_10711);
and U10802 (N_10802,N_10675,N_10706);
nand U10803 (N_10803,N_10704,N_10758);
nor U10804 (N_10804,N_10654,N_10714);
or U10805 (N_10805,N_10720,N_10795);
nand U10806 (N_10806,N_10674,N_10671);
or U10807 (N_10807,N_10652,N_10663);
and U10808 (N_10808,N_10776,N_10786);
nor U10809 (N_10809,N_10764,N_10673);
or U10810 (N_10810,N_10687,N_10682);
nand U10811 (N_10811,N_10698,N_10753);
xor U10812 (N_10812,N_10737,N_10740);
xnor U10813 (N_10813,N_10755,N_10686);
nand U10814 (N_10814,N_10728,N_10668);
nor U10815 (N_10815,N_10757,N_10703);
or U10816 (N_10816,N_10716,N_10696);
and U10817 (N_10817,N_10677,N_10700);
or U10818 (N_10818,N_10743,N_10708);
and U10819 (N_10819,N_10788,N_10688);
and U10820 (N_10820,N_10768,N_10713);
nand U10821 (N_10821,N_10779,N_10658);
or U10822 (N_10822,N_10705,N_10746);
or U10823 (N_10823,N_10756,N_10695);
nand U10824 (N_10824,N_10670,N_10791);
xor U10825 (N_10825,N_10747,N_10656);
nand U10826 (N_10826,N_10739,N_10683);
nand U10827 (N_10827,N_10702,N_10657);
and U10828 (N_10828,N_10774,N_10793);
nand U10829 (N_10829,N_10701,N_10731);
xor U10830 (N_10830,N_10699,N_10710);
nor U10831 (N_10831,N_10789,N_10717);
or U10832 (N_10832,N_10784,N_10722);
xor U10833 (N_10833,N_10678,N_10730);
nor U10834 (N_10834,N_10659,N_10761);
xor U10835 (N_10835,N_10715,N_10794);
nor U10836 (N_10836,N_10738,N_10787);
or U10837 (N_10837,N_10792,N_10766);
and U10838 (N_10838,N_10771,N_10735);
nor U10839 (N_10839,N_10729,N_10660);
nor U10840 (N_10840,N_10655,N_10751);
and U10841 (N_10841,N_10653,N_10726);
nor U10842 (N_10842,N_10721,N_10707);
or U10843 (N_10843,N_10797,N_10725);
nor U10844 (N_10844,N_10733,N_10681);
nor U10845 (N_10845,N_10773,N_10689);
nor U10846 (N_10846,N_10662,N_10679);
nor U10847 (N_10847,N_10763,N_10680);
nor U10848 (N_10848,N_10741,N_10749);
nand U10849 (N_10849,N_10667,N_10798);
nand U10850 (N_10850,N_10718,N_10790);
or U10851 (N_10851,N_10785,N_10781);
xnor U10852 (N_10852,N_10742,N_10734);
nand U10853 (N_10853,N_10650,N_10772);
or U10854 (N_10854,N_10752,N_10748);
and U10855 (N_10855,N_10672,N_10762);
and U10856 (N_10856,N_10691,N_10769);
nand U10857 (N_10857,N_10777,N_10727);
nand U10858 (N_10858,N_10669,N_10783);
and U10859 (N_10859,N_10778,N_10723);
xnor U10860 (N_10860,N_10676,N_10745);
and U10861 (N_10861,N_10661,N_10709);
nand U10862 (N_10862,N_10770,N_10775);
nor U10863 (N_10863,N_10719,N_10684);
nor U10864 (N_10864,N_10732,N_10693);
or U10865 (N_10865,N_10760,N_10750);
or U10866 (N_10866,N_10799,N_10744);
nand U10867 (N_10867,N_10690,N_10796);
or U10868 (N_10868,N_10736,N_10692);
nand U10869 (N_10869,N_10694,N_10665);
nand U10870 (N_10870,N_10780,N_10765);
nor U10871 (N_10871,N_10754,N_10651);
and U10872 (N_10872,N_10712,N_10724);
nor U10873 (N_10873,N_10666,N_10782);
and U10874 (N_10874,N_10697,N_10767);
or U10875 (N_10875,N_10717,N_10765);
nor U10876 (N_10876,N_10709,N_10721);
and U10877 (N_10877,N_10729,N_10730);
or U10878 (N_10878,N_10744,N_10696);
or U10879 (N_10879,N_10689,N_10734);
and U10880 (N_10880,N_10762,N_10660);
and U10881 (N_10881,N_10715,N_10664);
nor U10882 (N_10882,N_10691,N_10730);
and U10883 (N_10883,N_10751,N_10736);
xnor U10884 (N_10884,N_10750,N_10694);
and U10885 (N_10885,N_10756,N_10798);
nand U10886 (N_10886,N_10664,N_10766);
nand U10887 (N_10887,N_10690,N_10678);
or U10888 (N_10888,N_10748,N_10736);
nor U10889 (N_10889,N_10651,N_10665);
and U10890 (N_10890,N_10778,N_10682);
and U10891 (N_10891,N_10698,N_10736);
nand U10892 (N_10892,N_10697,N_10748);
nor U10893 (N_10893,N_10652,N_10674);
xor U10894 (N_10894,N_10686,N_10741);
or U10895 (N_10895,N_10755,N_10658);
and U10896 (N_10896,N_10731,N_10694);
nand U10897 (N_10897,N_10703,N_10709);
nand U10898 (N_10898,N_10736,N_10770);
and U10899 (N_10899,N_10741,N_10675);
xor U10900 (N_10900,N_10680,N_10789);
nor U10901 (N_10901,N_10685,N_10686);
or U10902 (N_10902,N_10662,N_10763);
or U10903 (N_10903,N_10799,N_10709);
nor U10904 (N_10904,N_10717,N_10666);
and U10905 (N_10905,N_10742,N_10656);
or U10906 (N_10906,N_10758,N_10710);
nand U10907 (N_10907,N_10739,N_10737);
or U10908 (N_10908,N_10668,N_10738);
xnor U10909 (N_10909,N_10753,N_10782);
or U10910 (N_10910,N_10697,N_10664);
nor U10911 (N_10911,N_10684,N_10657);
and U10912 (N_10912,N_10742,N_10759);
or U10913 (N_10913,N_10727,N_10743);
and U10914 (N_10914,N_10754,N_10700);
or U10915 (N_10915,N_10685,N_10767);
nand U10916 (N_10916,N_10765,N_10745);
xnor U10917 (N_10917,N_10775,N_10703);
nor U10918 (N_10918,N_10692,N_10729);
nor U10919 (N_10919,N_10682,N_10763);
nand U10920 (N_10920,N_10791,N_10676);
xnor U10921 (N_10921,N_10707,N_10703);
nand U10922 (N_10922,N_10780,N_10757);
and U10923 (N_10923,N_10688,N_10768);
nand U10924 (N_10924,N_10748,N_10666);
nand U10925 (N_10925,N_10760,N_10679);
or U10926 (N_10926,N_10748,N_10674);
nand U10927 (N_10927,N_10761,N_10790);
and U10928 (N_10928,N_10709,N_10771);
nand U10929 (N_10929,N_10723,N_10673);
nand U10930 (N_10930,N_10703,N_10745);
or U10931 (N_10931,N_10768,N_10666);
nand U10932 (N_10932,N_10661,N_10736);
xor U10933 (N_10933,N_10747,N_10736);
nor U10934 (N_10934,N_10758,N_10715);
and U10935 (N_10935,N_10784,N_10697);
nand U10936 (N_10936,N_10656,N_10774);
nor U10937 (N_10937,N_10720,N_10768);
or U10938 (N_10938,N_10671,N_10728);
or U10939 (N_10939,N_10799,N_10670);
nor U10940 (N_10940,N_10658,N_10743);
nand U10941 (N_10941,N_10769,N_10693);
nand U10942 (N_10942,N_10797,N_10653);
and U10943 (N_10943,N_10660,N_10750);
or U10944 (N_10944,N_10793,N_10722);
nand U10945 (N_10945,N_10705,N_10794);
and U10946 (N_10946,N_10660,N_10721);
xnor U10947 (N_10947,N_10726,N_10723);
nor U10948 (N_10948,N_10699,N_10716);
or U10949 (N_10949,N_10706,N_10685);
and U10950 (N_10950,N_10873,N_10827);
and U10951 (N_10951,N_10940,N_10942);
or U10952 (N_10952,N_10851,N_10880);
nor U10953 (N_10953,N_10914,N_10812);
or U10954 (N_10954,N_10815,N_10932);
nor U10955 (N_10955,N_10877,N_10903);
and U10956 (N_10956,N_10898,N_10947);
nor U10957 (N_10957,N_10829,N_10826);
or U10958 (N_10958,N_10806,N_10900);
nand U10959 (N_10959,N_10896,N_10853);
xnor U10960 (N_10960,N_10884,N_10869);
nor U10961 (N_10961,N_10852,N_10902);
nor U10962 (N_10962,N_10863,N_10872);
or U10963 (N_10963,N_10892,N_10839);
nand U10964 (N_10964,N_10838,N_10821);
and U10965 (N_10965,N_10890,N_10849);
nor U10966 (N_10966,N_10915,N_10921);
xnor U10967 (N_10967,N_10885,N_10943);
nand U10968 (N_10968,N_10830,N_10906);
and U10969 (N_10969,N_10866,N_10889);
nor U10970 (N_10970,N_10897,N_10822);
nand U10971 (N_10971,N_10928,N_10833);
and U10972 (N_10972,N_10917,N_10905);
or U10973 (N_10973,N_10816,N_10861);
nor U10974 (N_10974,N_10911,N_10819);
and U10975 (N_10975,N_10938,N_10842);
nor U10976 (N_10976,N_10926,N_10841);
nand U10977 (N_10977,N_10920,N_10811);
or U10978 (N_10978,N_10856,N_10931);
xor U10979 (N_10979,N_10860,N_10924);
xnor U10980 (N_10980,N_10882,N_10929);
nand U10981 (N_10981,N_10807,N_10946);
or U10982 (N_10982,N_10809,N_10803);
nor U10983 (N_10983,N_10824,N_10865);
or U10984 (N_10984,N_10840,N_10907);
nand U10985 (N_10985,N_10878,N_10944);
and U10986 (N_10986,N_10867,N_10904);
nor U10987 (N_10987,N_10883,N_10800);
or U10988 (N_10988,N_10808,N_10858);
nand U10989 (N_10989,N_10875,N_10941);
nand U10990 (N_10990,N_10848,N_10834);
nand U10991 (N_10991,N_10888,N_10870);
nand U10992 (N_10992,N_10881,N_10937);
nand U10993 (N_10993,N_10891,N_10876);
nor U10994 (N_10994,N_10908,N_10936);
or U10995 (N_10995,N_10930,N_10893);
nand U10996 (N_10996,N_10886,N_10933);
nor U10997 (N_10997,N_10948,N_10945);
nor U10998 (N_10998,N_10828,N_10817);
or U10999 (N_10999,N_10845,N_10820);
and U11000 (N_11000,N_10855,N_10802);
or U11001 (N_11001,N_10879,N_10887);
or U11002 (N_11002,N_10927,N_10805);
nand U11003 (N_11003,N_10949,N_10844);
nand U11004 (N_11004,N_10859,N_10899);
nand U11005 (N_11005,N_10854,N_10825);
nor U11006 (N_11006,N_10818,N_10874);
or U11007 (N_11007,N_10832,N_10801);
xor U11008 (N_11008,N_10895,N_10934);
nand U11009 (N_11009,N_10837,N_10918);
nor U11010 (N_11010,N_10909,N_10871);
nor U11011 (N_11011,N_10935,N_10846);
nand U11012 (N_11012,N_10850,N_10831);
xor U11013 (N_11013,N_10862,N_10814);
nand U11014 (N_11014,N_10910,N_10919);
and U11015 (N_11015,N_10894,N_10847);
xnor U11016 (N_11016,N_10836,N_10857);
and U11017 (N_11017,N_10939,N_10843);
and U11018 (N_11018,N_10868,N_10922);
nor U11019 (N_11019,N_10925,N_10864);
or U11020 (N_11020,N_10912,N_10835);
or U11021 (N_11021,N_10923,N_10901);
xor U11022 (N_11022,N_10804,N_10916);
xnor U11023 (N_11023,N_10810,N_10823);
or U11024 (N_11024,N_10813,N_10913);
xor U11025 (N_11025,N_10932,N_10865);
nand U11026 (N_11026,N_10878,N_10941);
or U11027 (N_11027,N_10938,N_10830);
nor U11028 (N_11028,N_10847,N_10860);
nand U11029 (N_11029,N_10906,N_10948);
and U11030 (N_11030,N_10942,N_10911);
nor U11031 (N_11031,N_10814,N_10929);
nand U11032 (N_11032,N_10867,N_10880);
or U11033 (N_11033,N_10906,N_10870);
nand U11034 (N_11034,N_10891,N_10921);
nor U11035 (N_11035,N_10807,N_10902);
and U11036 (N_11036,N_10893,N_10842);
nor U11037 (N_11037,N_10934,N_10941);
xor U11038 (N_11038,N_10896,N_10895);
xor U11039 (N_11039,N_10875,N_10800);
nand U11040 (N_11040,N_10840,N_10846);
or U11041 (N_11041,N_10814,N_10861);
nand U11042 (N_11042,N_10852,N_10938);
xnor U11043 (N_11043,N_10934,N_10944);
and U11044 (N_11044,N_10859,N_10872);
or U11045 (N_11045,N_10910,N_10936);
nand U11046 (N_11046,N_10879,N_10911);
nor U11047 (N_11047,N_10828,N_10853);
and U11048 (N_11048,N_10810,N_10948);
and U11049 (N_11049,N_10854,N_10842);
nor U11050 (N_11050,N_10862,N_10907);
or U11051 (N_11051,N_10916,N_10929);
and U11052 (N_11052,N_10828,N_10925);
nor U11053 (N_11053,N_10844,N_10825);
nor U11054 (N_11054,N_10842,N_10800);
nor U11055 (N_11055,N_10845,N_10948);
and U11056 (N_11056,N_10904,N_10918);
and U11057 (N_11057,N_10890,N_10932);
nor U11058 (N_11058,N_10859,N_10862);
nor U11059 (N_11059,N_10903,N_10926);
nor U11060 (N_11060,N_10825,N_10896);
nand U11061 (N_11061,N_10906,N_10935);
and U11062 (N_11062,N_10926,N_10891);
nor U11063 (N_11063,N_10941,N_10898);
xnor U11064 (N_11064,N_10914,N_10854);
and U11065 (N_11065,N_10862,N_10881);
nor U11066 (N_11066,N_10868,N_10813);
or U11067 (N_11067,N_10945,N_10847);
xnor U11068 (N_11068,N_10927,N_10835);
or U11069 (N_11069,N_10899,N_10817);
or U11070 (N_11070,N_10901,N_10832);
or U11071 (N_11071,N_10905,N_10808);
nand U11072 (N_11072,N_10816,N_10949);
nor U11073 (N_11073,N_10948,N_10904);
xor U11074 (N_11074,N_10941,N_10849);
or U11075 (N_11075,N_10900,N_10935);
or U11076 (N_11076,N_10919,N_10932);
nor U11077 (N_11077,N_10837,N_10817);
and U11078 (N_11078,N_10910,N_10844);
or U11079 (N_11079,N_10847,N_10879);
nor U11080 (N_11080,N_10926,N_10864);
xnor U11081 (N_11081,N_10898,N_10842);
xor U11082 (N_11082,N_10928,N_10838);
xor U11083 (N_11083,N_10873,N_10826);
or U11084 (N_11084,N_10852,N_10807);
or U11085 (N_11085,N_10924,N_10941);
xnor U11086 (N_11086,N_10848,N_10824);
nor U11087 (N_11087,N_10920,N_10938);
nand U11088 (N_11088,N_10870,N_10876);
nor U11089 (N_11089,N_10862,N_10852);
or U11090 (N_11090,N_10827,N_10922);
and U11091 (N_11091,N_10886,N_10830);
nand U11092 (N_11092,N_10806,N_10824);
nor U11093 (N_11093,N_10813,N_10935);
or U11094 (N_11094,N_10910,N_10862);
or U11095 (N_11095,N_10931,N_10875);
xor U11096 (N_11096,N_10947,N_10902);
xor U11097 (N_11097,N_10925,N_10907);
or U11098 (N_11098,N_10913,N_10886);
nor U11099 (N_11099,N_10891,N_10944);
xor U11100 (N_11100,N_10975,N_11017);
nand U11101 (N_11101,N_11072,N_11086);
and U11102 (N_11102,N_10996,N_11018);
xnor U11103 (N_11103,N_11024,N_11063);
nand U11104 (N_11104,N_11076,N_11020);
or U11105 (N_11105,N_11011,N_11037);
nand U11106 (N_11106,N_11029,N_11070);
nor U11107 (N_11107,N_11043,N_10990);
or U11108 (N_11108,N_11085,N_11016);
nand U11109 (N_11109,N_11044,N_11059);
nand U11110 (N_11110,N_11021,N_11040);
nor U11111 (N_11111,N_11054,N_11077);
xor U11112 (N_11112,N_11091,N_11071);
nor U11113 (N_11113,N_10976,N_10982);
nand U11114 (N_11114,N_11002,N_10994);
or U11115 (N_11115,N_11014,N_10952);
xor U11116 (N_11116,N_11045,N_10991);
and U11117 (N_11117,N_11039,N_11004);
and U11118 (N_11118,N_10983,N_10977);
xnor U11119 (N_11119,N_11060,N_11006);
and U11120 (N_11120,N_10987,N_10965);
xor U11121 (N_11121,N_11092,N_10953);
or U11122 (N_11122,N_10960,N_11010);
and U11123 (N_11123,N_11058,N_11097);
nand U11124 (N_11124,N_10968,N_10966);
and U11125 (N_11125,N_10951,N_11038);
and U11126 (N_11126,N_11025,N_10973);
nor U11127 (N_11127,N_11098,N_11003);
nand U11128 (N_11128,N_10964,N_11064);
and U11129 (N_11129,N_11046,N_10950);
or U11130 (N_11130,N_11000,N_10998);
and U11131 (N_11131,N_11047,N_10999);
nor U11132 (N_11132,N_10981,N_11087);
nor U11133 (N_11133,N_11026,N_10971);
and U11134 (N_11134,N_10961,N_11082);
nand U11135 (N_11135,N_11056,N_11096);
and U11136 (N_11136,N_11061,N_11093);
nand U11137 (N_11137,N_11009,N_11049);
and U11138 (N_11138,N_11074,N_11089);
or U11139 (N_11139,N_10985,N_11095);
xnor U11140 (N_11140,N_11055,N_11073);
nor U11141 (N_11141,N_11053,N_10954);
and U11142 (N_11142,N_11013,N_10988);
and U11143 (N_11143,N_10969,N_10967);
nor U11144 (N_11144,N_11062,N_11001);
and U11145 (N_11145,N_11050,N_10989);
or U11146 (N_11146,N_11041,N_11035);
nand U11147 (N_11147,N_11036,N_11084);
and U11148 (N_11148,N_10993,N_11042);
or U11149 (N_11149,N_11066,N_10958);
xor U11150 (N_11150,N_11080,N_10974);
nor U11151 (N_11151,N_10972,N_10970);
and U11152 (N_11152,N_10956,N_11081);
and U11153 (N_11153,N_11051,N_11012);
and U11154 (N_11154,N_10957,N_11094);
nand U11155 (N_11155,N_11083,N_11079);
nand U11156 (N_11156,N_10997,N_11057);
nand U11157 (N_11157,N_11068,N_10986);
and U11158 (N_11158,N_11015,N_10963);
or U11159 (N_11159,N_11075,N_10979);
nor U11160 (N_11160,N_11027,N_10955);
nor U11161 (N_11161,N_11005,N_11048);
or U11162 (N_11162,N_10978,N_10992);
and U11163 (N_11163,N_11030,N_11088);
or U11164 (N_11164,N_11034,N_10962);
or U11165 (N_11165,N_11032,N_11052);
and U11166 (N_11166,N_11019,N_10980);
or U11167 (N_11167,N_11067,N_11099);
xor U11168 (N_11168,N_10995,N_10959);
nand U11169 (N_11169,N_11090,N_10984);
nand U11170 (N_11170,N_11069,N_11007);
xor U11171 (N_11171,N_11022,N_11065);
nand U11172 (N_11172,N_11008,N_11078);
nand U11173 (N_11173,N_11028,N_11033);
xor U11174 (N_11174,N_11023,N_11031);
nand U11175 (N_11175,N_10976,N_11057);
nand U11176 (N_11176,N_11060,N_11077);
nand U11177 (N_11177,N_11012,N_10960);
xnor U11178 (N_11178,N_11031,N_10989);
nand U11179 (N_11179,N_11048,N_11039);
and U11180 (N_11180,N_11080,N_10960);
nor U11181 (N_11181,N_11073,N_11050);
xnor U11182 (N_11182,N_11071,N_10964);
and U11183 (N_11183,N_11091,N_10987);
nand U11184 (N_11184,N_11065,N_11080);
or U11185 (N_11185,N_11000,N_11021);
nand U11186 (N_11186,N_11001,N_10968);
nor U11187 (N_11187,N_10987,N_11096);
or U11188 (N_11188,N_10976,N_10968);
and U11189 (N_11189,N_10957,N_11077);
nand U11190 (N_11190,N_10970,N_11073);
xnor U11191 (N_11191,N_11069,N_10970);
xnor U11192 (N_11192,N_10985,N_11064);
or U11193 (N_11193,N_11083,N_11092);
or U11194 (N_11194,N_11081,N_11028);
nor U11195 (N_11195,N_10996,N_10992);
and U11196 (N_11196,N_11031,N_10986);
nor U11197 (N_11197,N_11009,N_11073);
or U11198 (N_11198,N_10988,N_11092);
nand U11199 (N_11199,N_11027,N_11080);
nand U11200 (N_11200,N_10983,N_10952);
nand U11201 (N_11201,N_11040,N_11069);
xor U11202 (N_11202,N_11064,N_11056);
and U11203 (N_11203,N_10970,N_11029);
xnor U11204 (N_11204,N_11004,N_11001);
nor U11205 (N_11205,N_11036,N_11038);
or U11206 (N_11206,N_10950,N_10963);
or U11207 (N_11207,N_10973,N_10969);
nand U11208 (N_11208,N_11001,N_11098);
nor U11209 (N_11209,N_10986,N_11095);
xnor U11210 (N_11210,N_11003,N_11099);
or U11211 (N_11211,N_10950,N_11099);
or U11212 (N_11212,N_11013,N_10968);
nand U11213 (N_11213,N_10956,N_11050);
or U11214 (N_11214,N_11016,N_10990);
or U11215 (N_11215,N_11088,N_11067);
nor U11216 (N_11216,N_11019,N_10950);
nor U11217 (N_11217,N_11087,N_11086);
nand U11218 (N_11218,N_11023,N_11059);
and U11219 (N_11219,N_10964,N_11085);
nor U11220 (N_11220,N_11083,N_11057);
nand U11221 (N_11221,N_11084,N_10984);
nor U11222 (N_11222,N_11081,N_11070);
or U11223 (N_11223,N_11080,N_11032);
and U11224 (N_11224,N_11001,N_11084);
nor U11225 (N_11225,N_10987,N_11068);
or U11226 (N_11226,N_11081,N_10959);
or U11227 (N_11227,N_11040,N_11097);
or U11228 (N_11228,N_11021,N_10958);
and U11229 (N_11229,N_11099,N_11056);
and U11230 (N_11230,N_11025,N_11026);
nand U11231 (N_11231,N_11016,N_11047);
xor U11232 (N_11232,N_11047,N_10992);
nand U11233 (N_11233,N_11087,N_11022);
nand U11234 (N_11234,N_11082,N_11068);
and U11235 (N_11235,N_10959,N_11008);
or U11236 (N_11236,N_11076,N_11091);
and U11237 (N_11237,N_11098,N_10986);
nor U11238 (N_11238,N_11017,N_10981);
nand U11239 (N_11239,N_11036,N_11088);
or U11240 (N_11240,N_11080,N_10966);
nor U11241 (N_11241,N_11049,N_10999);
xor U11242 (N_11242,N_10981,N_11005);
and U11243 (N_11243,N_10984,N_10979);
and U11244 (N_11244,N_11033,N_11052);
or U11245 (N_11245,N_11050,N_11060);
or U11246 (N_11246,N_11093,N_11065);
nand U11247 (N_11247,N_11034,N_10996);
nand U11248 (N_11248,N_11061,N_10979);
and U11249 (N_11249,N_11072,N_11037);
or U11250 (N_11250,N_11131,N_11245);
nand U11251 (N_11251,N_11236,N_11239);
xnor U11252 (N_11252,N_11249,N_11108);
nor U11253 (N_11253,N_11170,N_11198);
xor U11254 (N_11254,N_11174,N_11101);
nand U11255 (N_11255,N_11159,N_11242);
or U11256 (N_11256,N_11109,N_11221);
nor U11257 (N_11257,N_11199,N_11189);
nor U11258 (N_11258,N_11202,N_11179);
and U11259 (N_11259,N_11115,N_11120);
and U11260 (N_11260,N_11204,N_11243);
and U11261 (N_11261,N_11196,N_11223);
xnor U11262 (N_11262,N_11110,N_11100);
nor U11263 (N_11263,N_11232,N_11201);
nor U11264 (N_11264,N_11103,N_11205);
or U11265 (N_11265,N_11184,N_11144);
or U11266 (N_11266,N_11188,N_11134);
nor U11267 (N_11267,N_11225,N_11231);
nand U11268 (N_11268,N_11137,N_11146);
or U11269 (N_11269,N_11126,N_11162);
or U11270 (N_11270,N_11140,N_11186);
nor U11271 (N_11271,N_11234,N_11207);
or U11272 (N_11272,N_11136,N_11183);
and U11273 (N_11273,N_11133,N_11209);
or U11274 (N_11274,N_11244,N_11158);
or U11275 (N_11275,N_11116,N_11128);
or U11276 (N_11276,N_11104,N_11121);
or U11277 (N_11277,N_11138,N_11233);
or U11278 (N_11278,N_11241,N_11227);
nor U11279 (N_11279,N_11178,N_11155);
or U11280 (N_11280,N_11106,N_11210);
nor U11281 (N_11281,N_11102,N_11105);
or U11282 (N_11282,N_11139,N_11132);
xor U11283 (N_11283,N_11119,N_11224);
or U11284 (N_11284,N_11129,N_11226);
or U11285 (N_11285,N_11185,N_11117);
nor U11286 (N_11286,N_11157,N_11143);
nor U11287 (N_11287,N_11176,N_11194);
or U11288 (N_11288,N_11214,N_11216);
and U11289 (N_11289,N_11125,N_11169);
or U11290 (N_11290,N_11175,N_11180);
nor U11291 (N_11291,N_11152,N_11193);
or U11292 (N_11292,N_11248,N_11148);
and U11293 (N_11293,N_11177,N_11163);
nor U11294 (N_11294,N_11124,N_11111);
or U11295 (N_11295,N_11212,N_11215);
nor U11296 (N_11296,N_11208,N_11200);
or U11297 (N_11297,N_11171,N_11156);
nand U11298 (N_11298,N_11230,N_11166);
nand U11299 (N_11299,N_11122,N_11213);
or U11300 (N_11300,N_11167,N_11147);
nor U11301 (N_11301,N_11222,N_11246);
nor U11302 (N_11302,N_11150,N_11118);
nor U11303 (N_11303,N_11141,N_11135);
and U11304 (N_11304,N_11229,N_11191);
nand U11305 (N_11305,N_11203,N_11165);
and U11306 (N_11306,N_11219,N_11168);
or U11307 (N_11307,N_11187,N_11238);
nand U11308 (N_11308,N_11151,N_11114);
nor U11309 (N_11309,N_11211,N_11197);
and U11310 (N_11310,N_11195,N_11235);
and U11311 (N_11311,N_11123,N_11220);
xor U11312 (N_11312,N_11182,N_11142);
and U11313 (N_11313,N_11228,N_11247);
nor U11314 (N_11314,N_11160,N_11173);
or U11315 (N_11315,N_11164,N_11153);
or U11316 (N_11316,N_11145,N_11112);
nor U11317 (N_11317,N_11161,N_11240);
nor U11318 (N_11318,N_11237,N_11206);
nand U11319 (N_11319,N_11217,N_11127);
and U11320 (N_11320,N_11172,N_11218);
nor U11321 (N_11321,N_11181,N_11113);
or U11322 (N_11322,N_11190,N_11192);
or U11323 (N_11323,N_11130,N_11154);
or U11324 (N_11324,N_11107,N_11149);
or U11325 (N_11325,N_11194,N_11222);
nor U11326 (N_11326,N_11142,N_11238);
and U11327 (N_11327,N_11149,N_11109);
and U11328 (N_11328,N_11204,N_11129);
nand U11329 (N_11329,N_11184,N_11127);
or U11330 (N_11330,N_11137,N_11141);
or U11331 (N_11331,N_11105,N_11243);
nor U11332 (N_11332,N_11122,N_11148);
nand U11333 (N_11333,N_11191,N_11159);
nand U11334 (N_11334,N_11138,N_11202);
nor U11335 (N_11335,N_11102,N_11224);
and U11336 (N_11336,N_11180,N_11136);
and U11337 (N_11337,N_11236,N_11104);
nor U11338 (N_11338,N_11244,N_11120);
nand U11339 (N_11339,N_11235,N_11244);
nand U11340 (N_11340,N_11123,N_11180);
nand U11341 (N_11341,N_11128,N_11240);
or U11342 (N_11342,N_11189,N_11198);
or U11343 (N_11343,N_11183,N_11224);
nand U11344 (N_11344,N_11211,N_11165);
or U11345 (N_11345,N_11112,N_11109);
nor U11346 (N_11346,N_11171,N_11158);
nor U11347 (N_11347,N_11190,N_11127);
nor U11348 (N_11348,N_11163,N_11194);
xor U11349 (N_11349,N_11196,N_11183);
and U11350 (N_11350,N_11208,N_11131);
nand U11351 (N_11351,N_11243,N_11207);
or U11352 (N_11352,N_11196,N_11212);
nor U11353 (N_11353,N_11212,N_11121);
and U11354 (N_11354,N_11245,N_11234);
or U11355 (N_11355,N_11218,N_11249);
xor U11356 (N_11356,N_11137,N_11230);
nor U11357 (N_11357,N_11193,N_11122);
nand U11358 (N_11358,N_11226,N_11156);
nand U11359 (N_11359,N_11234,N_11109);
and U11360 (N_11360,N_11168,N_11147);
xnor U11361 (N_11361,N_11188,N_11174);
and U11362 (N_11362,N_11225,N_11139);
and U11363 (N_11363,N_11248,N_11190);
and U11364 (N_11364,N_11160,N_11207);
nor U11365 (N_11365,N_11180,N_11193);
nand U11366 (N_11366,N_11108,N_11106);
or U11367 (N_11367,N_11199,N_11177);
and U11368 (N_11368,N_11135,N_11148);
or U11369 (N_11369,N_11186,N_11183);
nor U11370 (N_11370,N_11231,N_11205);
and U11371 (N_11371,N_11222,N_11162);
nor U11372 (N_11372,N_11248,N_11157);
xor U11373 (N_11373,N_11245,N_11203);
and U11374 (N_11374,N_11211,N_11191);
or U11375 (N_11375,N_11157,N_11205);
or U11376 (N_11376,N_11102,N_11175);
and U11377 (N_11377,N_11113,N_11109);
nand U11378 (N_11378,N_11162,N_11246);
and U11379 (N_11379,N_11138,N_11211);
nor U11380 (N_11380,N_11246,N_11110);
xnor U11381 (N_11381,N_11240,N_11247);
xor U11382 (N_11382,N_11103,N_11197);
xnor U11383 (N_11383,N_11194,N_11228);
nor U11384 (N_11384,N_11248,N_11128);
or U11385 (N_11385,N_11237,N_11129);
nand U11386 (N_11386,N_11206,N_11193);
or U11387 (N_11387,N_11115,N_11160);
nor U11388 (N_11388,N_11248,N_11129);
nand U11389 (N_11389,N_11159,N_11139);
nand U11390 (N_11390,N_11236,N_11143);
nor U11391 (N_11391,N_11172,N_11103);
or U11392 (N_11392,N_11170,N_11103);
nor U11393 (N_11393,N_11107,N_11186);
and U11394 (N_11394,N_11247,N_11103);
or U11395 (N_11395,N_11210,N_11160);
nor U11396 (N_11396,N_11228,N_11173);
nand U11397 (N_11397,N_11187,N_11185);
nand U11398 (N_11398,N_11111,N_11150);
and U11399 (N_11399,N_11185,N_11180);
nand U11400 (N_11400,N_11395,N_11386);
and U11401 (N_11401,N_11353,N_11262);
nor U11402 (N_11402,N_11287,N_11374);
nor U11403 (N_11403,N_11277,N_11317);
or U11404 (N_11404,N_11267,N_11336);
nand U11405 (N_11405,N_11261,N_11278);
nand U11406 (N_11406,N_11371,N_11296);
nor U11407 (N_11407,N_11391,N_11310);
or U11408 (N_11408,N_11389,N_11297);
xor U11409 (N_11409,N_11368,N_11344);
and U11410 (N_11410,N_11376,N_11300);
nand U11411 (N_11411,N_11334,N_11303);
or U11412 (N_11412,N_11378,N_11316);
or U11413 (N_11413,N_11327,N_11359);
or U11414 (N_11414,N_11280,N_11363);
nor U11415 (N_11415,N_11319,N_11314);
and U11416 (N_11416,N_11292,N_11325);
xnor U11417 (N_11417,N_11388,N_11264);
or U11418 (N_11418,N_11383,N_11288);
nor U11419 (N_11419,N_11356,N_11259);
or U11420 (N_11420,N_11321,N_11322);
or U11421 (N_11421,N_11255,N_11384);
nand U11422 (N_11422,N_11290,N_11393);
or U11423 (N_11423,N_11329,N_11364);
and U11424 (N_11424,N_11279,N_11362);
and U11425 (N_11425,N_11373,N_11390);
or U11426 (N_11426,N_11294,N_11304);
or U11427 (N_11427,N_11355,N_11394);
nand U11428 (N_11428,N_11369,N_11380);
and U11429 (N_11429,N_11399,N_11252);
and U11430 (N_11430,N_11342,N_11269);
xor U11431 (N_11431,N_11349,N_11282);
nand U11432 (N_11432,N_11251,N_11268);
and U11433 (N_11433,N_11256,N_11347);
and U11434 (N_11434,N_11358,N_11375);
nor U11435 (N_11435,N_11324,N_11397);
and U11436 (N_11436,N_11345,N_11318);
nand U11437 (N_11437,N_11381,N_11293);
xnor U11438 (N_11438,N_11331,N_11270);
nor U11439 (N_11439,N_11265,N_11350);
nor U11440 (N_11440,N_11313,N_11257);
and U11441 (N_11441,N_11308,N_11352);
and U11442 (N_11442,N_11275,N_11366);
nand U11443 (N_11443,N_11299,N_11295);
and U11444 (N_11444,N_11340,N_11260);
or U11445 (N_11445,N_11354,N_11398);
or U11446 (N_11446,N_11289,N_11357);
or U11447 (N_11447,N_11272,N_11273);
nand U11448 (N_11448,N_11323,N_11337);
or U11449 (N_11449,N_11335,N_11339);
and U11450 (N_11450,N_11305,N_11320);
and U11451 (N_11451,N_11274,N_11254);
nand U11452 (N_11452,N_11382,N_11250);
nand U11453 (N_11453,N_11370,N_11286);
nor U11454 (N_11454,N_11379,N_11387);
nand U11455 (N_11455,N_11306,N_11253);
xor U11456 (N_11456,N_11309,N_11291);
nor U11457 (N_11457,N_11298,N_11281);
nand U11458 (N_11458,N_11258,N_11263);
nor U11459 (N_11459,N_11330,N_11307);
nor U11460 (N_11460,N_11348,N_11343);
and U11461 (N_11461,N_11301,N_11302);
and U11462 (N_11462,N_11328,N_11266);
nand U11463 (N_11463,N_11367,N_11341);
or U11464 (N_11464,N_11361,N_11315);
nor U11465 (N_11465,N_11326,N_11333);
and U11466 (N_11466,N_11284,N_11396);
and U11467 (N_11467,N_11392,N_11385);
nand U11468 (N_11468,N_11271,N_11365);
and U11469 (N_11469,N_11311,N_11338);
and U11470 (N_11470,N_11372,N_11276);
nor U11471 (N_11471,N_11377,N_11312);
or U11472 (N_11472,N_11351,N_11360);
nand U11473 (N_11473,N_11285,N_11346);
nand U11474 (N_11474,N_11332,N_11283);
and U11475 (N_11475,N_11290,N_11373);
nor U11476 (N_11476,N_11351,N_11268);
nor U11477 (N_11477,N_11344,N_11380);
nand U11478 (N_11478,N_11272,N_11380);
and U11479 (N_11479,N_11357,N_11288);
or U11480 (N_11480,N_11389,N_11285);
nor U11481 (N_11481,N_11354,N_11313);
nand U11482 (N_11482,N_11338,N_11372);
nand U11483 (N_11483,N_11393,N_11380);
and U11484 (N_11484,N_11301,N_11379);
and U11485 (N_11485,N_11367,N_11346);
xor U11486 (N_11486,N_11354,N_11295);
nand U11487 (N_11487,N_11295,N_11381);
nand U11488 (N_11488,N_11399,N_11322);
nand U11489 (N_11489,N_11285,N_11348);
or U11490 (N_11490,N_11366,N_11374);
nand U11491 (N_11491,N_11264,N_11297);
nor U11492 (N_11492,N_11318,N_11357);
nor U11493 (N_11493,N_11262,N_11327);
and U11494 (N_11494,N_11314,N_11253);
nand U11495 (N_11495,N_11354,N_11270);
and U11496 (N_11496,N_11373,N_11317);
nor U11497 (N_11497,N_11257,N_11310);
xor U11498 (N_11498,N_11271,N_11318);
and U11499 (N_11499,N_11315,N_11344);
xor U11500 (N_11500,N_11351,N_11329);
and U11501 (N_11501,N_11320,N_11273);
or U11502 (N_11502,N_11336,N_11261);
nand U11503 (N_11503,N_11354,N_11382);
and U11504 (N_11504,N_11280,N_11251);
nor U11505 (N_11505,N_11292,N_11268);
nor U11506 (N_11506,N_11288,N_11381);
or U11507 (N_11507,N_11363,N_11304);
or U11508 (N_11508,N_11353,N_11319);
and U11509 (N_11509,N_11274,N_11328);
nand U11510 (N_11510,N_11287,N_11286);
nor U11511 (N_11511,N_11370,N_11358);
nor U11512 (N_11512,N_11280,N_11257);
or U11513 (N_11513,N_11264,N_11308);
or U11514 (N_11514,N_11357,N_11262);
or U11515 (N_11515,N_11375,N_11251);
and U11516 (N_11516,N_11295,N_11259);
nor U11517 (N_11517,N_11392,N_11317);
nor U11518 (N_11518,N_11371,N_11322);
or U11519 (N_11519,N_11343,N_11271);
and U11520 (N_11520,N_11310,N_11367);
nand U11521 (N_11521,N_11305,N_11332);
and U11522 (N_11522,N_11337,N_11373);
and U11523 (N_11523,N_11347,N_11335);
nor U11524 (N_11524,N_11362,N_11319);
and U11525 (N_11525,N_11319,N_11253);
and U11526 (N_11526,N_11292,N_11274);
and U11527 (N_11527,N_11311,N_11289);
nand U11528 (N_11528,N_11376,N_11262);
nand U11529 (N_11529,N_11341,N_11312);
and U11530 (N_11530,N_11360,N_11304);
xor U11531 (N_11531,N_11300,N_11375);
or U11532 (N_11532,N_11324,N_11398);
nand U11533 (N_11533,N_11288,N_11368);
nand U11534 (N_11534,N_11279,N_11263);
nand U11535 (N_11535,N_11271,N_11257);
and U11536 (N_11536,N_11310,N_11327);
xor U11537 (N_11537,N_11369,N_11270);
nand U11538 (N_11538,N_11397,N_11358);
nor U11539 (N_11539,N_11283,N_11382);
nor U11540 (N_11540,N_11254,N_11387);
and U11541 (N_11541,N_11384,N_11324);
nand U11542 (N_11542,N_11251,N_11285);
or U11543 (N_11543,N_11390,N_11269);
nor U11544 (N_11544,N_11347,N_11368);
nor U11545 (N_11545,N_11261,N_11372);
and U11546 (N_11546,N_11312,N_11308);
nand U11547 (N_11547,N_11268,N_11278);
and U11548 (N_11548,N_11254,N_11372);
nand U11549 (N_11549,N_11349,N_11317);
xor U11550 (N_11550,N_11495,N_11474);
and U11551 (N_11551,N_11541,N_11419);
xor U11552 (N_11552,N_11532,N_11498);
or U11553 (N_11553,N_11483,N_11461);
xnor U11554 (N_11554,N_11432,N_11416);
nor U11555 (N_11555,N_11443,N_11452);
or U11556 (N_11556,N_11525,N_11517);
and U11557 (N_11557,N_11439,N_11431);
nor U11558 (N_11558,N_11481,N_11410);
xor U11559 (N_11559,N_11479,N_11464);
nor U11560 (N_11560,N_11454,N_11546);
or U11561 (N_11561,N_11408,N_11496);
xor U11562 (N_11562,N_11448,N_11426);
and U11563 (N_11563,N_11418,N_11515);
nor U11564 (N_11564,N_11476,N_11471);
nand U11565 (N_11565,N_11484,N_11433);
nand U11566 (N_11566,N_11421,N_11489);
nor U11567 (N_11567,N_11453,N_11523);
xor U11568 (N_11568,N_11466,N_11521);
xnor U11569 (N_11569,N_11405,N_11486);
and U11570 (N_11570,N_11442,N_11457);
nor U11571 (N_11571,N_11465,N_11492);
nor U11572 (N_11572,N_11530,N_11444);
nand U11573 (N_11573,N_11407,N_11445);
nand U11574 (N_11574,N_11460,N_11545);
nor U11575 (N_11575,N_11509,N_11503);
xor U11576 (N_11576,N_11406,N_11537);
nor U11577 (N_11577,N_11459,N_11548);
or U11578 (N_11578,N_11415,N_11516);
xor U11579 (N_11579,N_11539,N_11513);
nand U11580 (N_11580,N_11413,N_11529);
xnor U11581 (N_11581,N_11451,N_11424);
or U11582 (N_11582,N_11536,N_11543);
nand U11583 (N_11583,N_11508,N_11518);
xnor U11584 (N_11584,N_11535,N_11512);
nor U11585 (N_11585,N_11475,N_11469);
nand U11586 (N_11586,N_11429,N_11470);
nor U11587 (N_11587,N_11511,N_11531);
nand U11588 (N_11588,N_11506,N_11420);
and U11589 (N_11589,N_11544,N_11491);
xnor U11590 (N_11590,N_11458,N_11417);
nand U11591 (N_11591,N_11528,N_11425);
nand U11592 (N_11592,N_11542,N_11414);
nand U11593 (N_11593,N_11477,N_11501);
nor U11594 (N_11594,N_11463,N_11514);
nor U11595 (N_11595,N_11534,N_11409);
nor U11596 (N_11596,N_11480,N_11447);
nor U11597 (N_11597,N_11502,N_11423);
nor U11598 (N_11598,N_11450,N_11427);
nand U11599 (N_11599,N_11499,N_11526);
or U11600 (N_11600,N_11500,N_11504);
and U11601 (N_11601,N_11449,N_11497);
nand U11602 (N_11602,N_11527,N_11441);
xnor U11603 (N_11603,N_11403,N_11533);
nand U11604 (N_11604,N_11490,N_11422);
or U11605 (N_11605,N_11524,N_11507);
nor U11606 (N_11606,N_11434,N_11411);
and U11607 (N_11607,N_11485,N_11430);
and U11608 (N_11608,N_11473,N_11402);
and U11609 (N_11609,N_11437,N_11494);
and U11610 (N_11610,N_11467,N_11487);
nor U11611 (N_11611,N_11482,N_11478);
or U11612 (N_11612,N_11404,N_11401);
or U11613 (N_11613,N_11455,N_11538);
or U11614 (N_11614,N_11505,N_11519);
or U11615 (N_11615,N_11440,N_11446);
or U11616 (N_11616,N_11438,N_11522);
and U11617 (N_11617,N_11549,N_11547);
nand U11618 (N_11618,N_11493,N_11472);
nor U11619 (N_11619,N_11400,N_11468);
and U11620 (N_11620,N_11428,N_11540);
or U11621 (N_11621,N_11456,N_11488);
and U11622 (N_11622,N_11435,N_11412);
and U11623 (N_11623,N_11520,N_11510);
nand U11624 (N_11624,N_11462,N_11436);
or U11625 (N_11625,N_11412,N_11443);
or U11626 (N_11626,N_11531,N_11480);
or U11627 (N_11627,N_11549,N_11431);
nand U11628 (N_11628,N_11460,N_11471);
nor U11629 (N_11629,N_11407,N_11538);
and U11630 (N_11630,N_11506,N_11446);
or U11631 (N_11631,N_11525,N_11484);
nor U11632 (N_11632,N_11482,N_11509);
and U11633 (N_11633,N_11403,N_11477);
or U11634 (N_11634,N_11415,N_11494);
xnor U11635 (N_11635,N_11454,N_11526);
nand U11636 (N_11636,N_11482,N_11485);
or U11637 (N_11637,N_11448,N_11511);
and U11638 (N_11638,N_11547,N_11431);
nor U11639 (N_11639,N_11401,N_11530);
and U11640 (N_11640,N_11418,N_11529);
nand U11641 (N_11641,N_11444,N_11450);
xnor U11642 (N_11642,N_11436,N_11458);
nor U11643 (N_11643,N_11449,N_11471);
or U11644 (N_11644,N_11445,N_11467);
xor U11645 (N_11645,N_11453,N_11434);
xor U11646 (N_11646,N_11403,N_11501);
nand U11647 (N_11647,N_11537,N_11444);
xnor U11648 (N_11648,N_11534,N_11491);
nor U11649 (N_11649,N_11410,N_11409);
or U11650 (N_11650,N_11464,N_11424);
or U11651 (N_11651,N_11513,N_11453);
xor U11652 (N_11652,N_11492,N_11523);
or U11653 (N_11653,N_11407,N_11457);
or U11654 (N_11654,N_11425,N_11518);
nor U11655 (N_11655,N_11471,N_11507);
or U11656 (N_11656,N_11544,N_11549);
nor U11657 (N_11657,N_11533,N_11433);
nand U11658 (N_11658,N_11506,N_11445);
xor U11659 (N_11659,N_11487,N_11544);
and U11660 (N_11660,N_11549,N_11546);
nor U11661 (N_11661,N_11493,N_11525);
and U11662 (N_11662,N_11458,N_11524);
and U11663 (N_11663,N_11510,N_11493);
nor U11664 (N_11664,N_11513,N_11401);
and U11665 (N_11665,N_11483,N_11455);
and U11666 (N_11666,N_11483,N_11499);
nor U11667 (N_11667,N_11470,N_11418);
or U11668 (N_11668,N_11493,N_11543);
nor U11669 (N_11669,N_11409,N_11427);
nor U11670 (N_11670,N_11419,N_11490);
nand U11671 (N_11671,N_11454,N_11446);
xor U11672 (N_11672,N_11502,N_11429);
nand U11673 (N_11673,N_11490,N_11446);
nand U11674 (N_11674,N_11487,N_11409);
nor U11675 (N_11675,N_11524,N_11476);
nand U11676 (N_11676,N_11408,N_11502);
xnor U11677 (N_11677,N_11430,N_11415);
nor U11678 (N_11678,N_11437,N_11422);
or U11679 (N_11679,N_11421,N_11542);
and U11680 (N_11680,N_11509,N_11496);
and U11681 (N_11681,N_11451,N_11509);
nand U11682 (N_11682,N_11452,N_11524);
or U11683 (N_11683,N_11435,N_11513);
nand U11684 (N_11684,N_11452,N_11466);
and U11685 (N_11685,N_11538,N_11541);
xnor U11686 (N_11686,N_11424,N_11433);
or U11687 (N_11687,N_11532,N_11410);
nor U11688 (N_11688,N_11447,N_11543);
nand U11689 (N_11689,N_11450,N_11489);
nor U11690 (N_11690,N_11496,N_11514);
nor U11691 (N_11691,N_11477,N_11506);
or U11692 (N_11692,N_11480,N_11472);
nand U11693 (N_11693,N_11521,N_11504);
or U11694 (N_11694,N_11440,N_11466);
nand U11695 (N_11695,N_11533,N_11490);
xor U11696 (N_11696,N_11545,N_11530);
nor U11697 (N_11697,N_11419,N_11448);
or U11698 (N_11698,N_11459,N_11425);
nor U11699 (N_11699,N_11521,N_11487);
xnor U11700 (N_11700,N_11628,N_11626);
nor U11701 (N_11701,N_11666,N_11682);
nand U11702 (N_11702,N_11603,N_11675);
and U11703 (N_11703,N_11601,N_11575);
nand U11704 (N_11704,N_11595,N_11661);
nor U11705 (N_11705,N_11642,N_11645);
nand U11706 (N_11706,N_11663,N_11664);
nor U11707 (N_11707,N_11632,N_11689);
nor U11708 (N_11708,N_11611,N_11670);
nor U11709 (N_11709,N_11580,N_11563);
nand U11710 (N_11710,N_11690,N_11568);
and U11711 (N_11711,N_11684,N_11556);
or U11712 (N_11712,N_11625,N_11636);
nor U11713 (N_11713,N_11671,N_11565);
or U11714 (N_11714,N_11630,N_11660);
or U11715 (N_11715,N_11559,N_11685);
xor U11716 (N_11716,N_11620,N_11695);
and U11717 (N_11717,N_11607,N_11589);
or U11718 (N_11718,N_11644,N_11581);
or U11719 (N_11719,N_11653,N_11584);
nand U11720 (N_11720,N_11631,N_11696);
or U11721 (N_11721,N_11615,N_11606);
nor U11722 (N_11722,N_11564,N_11640);
or U11723 (N_11723,N_11635,N_11567);
nor U11724 (N_11724,N_11588,N_11698);
or U11725 (N_11725,N_11592,N_11597);
nor U11726 (N_11726,N_11674,N_11639);
nor U11727 (N_11727,N_11649,N_11554);
or U11728 (N_11728,N_11622,N_11599);
nor U11729 (N_11729,N_11629,N_11657);
and U11730 (N_11730,N_11551,N_11694);
xnor U11731 (N_11731,N_11573,N_11619);
nand U11732 (N_11732,N_11687,N_11633);
nand U11733 (N_11733,N_11656,N_11553);
nand U11734 (N_11734,N_11693,N_11651);
or U11735 (N_11735,N_11550,N_11621);
and U11736 (N_11736,N_11624,N_11688);
nand U11737 (N_11737,N_11578,N_11579);
nand U11738 (N_11738,N_11654,N_11591);
nand U11739 (N_11739,N_11600,N_11561);
xnor U11740 (N_11740,N_11623,N_11634);
and U11741 (N_11741,N_11638,N_11614);
nor U11742 (N_11742,N_11678,N_11557);
nor U11743 (N_11743,N_11604,N_11667);
nand U11744 (N_11744,N_11570,N_11583);
xor U11745 (N_11745,N_11683,N_11594);
nand U11746 (N_11746,N_11655,N_11598);
and U11747 (N_11747,N_11691,N_11648);
or U11748 (N_11748,N_11608,N_11569);
or U11749 (N_11749,N_11587,N_11571);
nand U11750 (N_11750,N_11646,N_11586);
or U11751 (N_11751,N_11665,N_11617);
or U11752 (N_11752,N_11555,N_11652);
nand U11753 (N_11753,N_11676,N_11643);
and U11754 (N_11754,N_11596,N_11552);
and U11755 (N_11755,N_11610,N_11616);
nand U11756 (N_11756,N_11612,N_11647);
and U11757 (N_11757,N_11699,N_11593);
nand U11758 (N_11758,N_11577,N_11613);
nor U11759 (N_11759,N_11641,N_11680);
nor U11760 (N_11760,N_11692,N_11672);
nand U11761 (N_11761,N_11560,N_11627);
nor U11762 (N_11762,N_11677,N_11576);
or U11763 (N_11763,N_11668,N_11679);
nor U11764 (N_11764,N_11686,N_11609);
xnor U11765 (N_11765,N_11659,N_11650);
nand U11766 (N_11766,N_11562,N_11697);
and U11767 (N_11767,N_11572,N_11681);
nand U11768 (N_11768,N_11618,N_11637);
and U11769 (N_11769,N_11574,N_11582);
and U11770 (N_11770,N_11673,N_11590);
nand U11771 (N_11771,N_11658,N_11602);
nand U11772 (N_11772,N_11585,N_11566);
nor U11773 (N_11773,N_11558,N_11669);
nor U11774 (N_11774,N_11662,N_11605);
and U11775 (N_11775,N_11565,N_11584);
nand U11776 (N_11776,N_11550,N_11695);
and U11777 (N_11777,N_11562,N_11690);
nor U11778 (N_11778,N_11640,N_11587);
nor U11779 (N_11779,N_11669,N_11673);
xor U11780 (N_11780,N_11667,N_11568);
xnor U11781 (N_11781,N_11616,N_11633);
and U11782 (N_11782,N_11667,N_11576);
or U11783 (N_11783,N_11622,N_11619);
or U11784 (N_11784,N_11691,N_11644);
nand U11785 (N_11785,N_11631,N_11560);
nand U11786 (N_11786,N_11681,N_11551);
nand U11787 (N_11787,N_11643,N_11639);
nand U11788 (N_11788,N_11622,N_11573);
nor U11789 (N_11789,N_11612,N_11689);
or U11790 (N_11790,N_11608,N_11582);
or U11791 (N_11791,N_11576,N_11554);
nand U11792 (N_11792,N_11685,N_11626);
or U11793 (N_11793,N_11617,N_11673);
and U11794 (N_11794,N_11670,N_11675);
or U11795 (N_11795,N_11593,N_11605);
nand U11796 (N_11796,N_11593,N_11567);
or U11797 (N_11797,N_11695,N_11555);
xor U11798 (N_11798,N_11601,N_11627);
or U11799 (N_11799,N_11683,N_11682);
and U11800 (N_11800,N_11576,N_11599);
xnor U11801 (N_11801,N_11559,N_11646);
nand U11802 (N_11802,N_11655,N_11592);
nor U11803 (N_11803,N_11643,N_11615);
or U11804 (N_11804,N_11591,N_11565);
nand U11805 (N_11805,N_11653,N_11669);
nor U11806 (N_11806,N_11672,N_11571);
nor U11807 (N_11807,N_11607,N_11602);
nor U11808 (N_11808,N_11670,N_11639);
or U11809 (N_11809,N_11653,N_11576);
and U11810 (N_11810,N_11594,N_11668);
and U11811 (N_11811,N_11642,N_11652);
and U11812 (N_11812,N_11627,N_11564);
xor U11813 (N_11813,N_11618,N_11644);
nand U11814 (N_11814,N_11570,N_11625);
and U11815 (N_11815,N_11662,N_11612);
nand U11816 (N_11816,N_11582,N_11664);
xnor U11817 (N_11817,N_11592,N_11699);
and U11818 (N_11818,N_11567,N_11550);
and U11819 (N_11819,N_11599,N_11616);
or U11820 (N_11820,N_11615,N_11695);
nor U11821 (N_11821,N_11695,N_11688);
or U11822 (N_11822,N_11584,N_11647);
xor U11823 (N_11823,N_11648,N_11631);
nand U11824 (N_11824,N_11679,N_11587);
nand U11825 (N_11825,N_11689,N_11664);
nand U11826 (N_11826,N_11607,N_11658);
nand U11827 (N_11827,N_11678,N_11683);
nand U11828 (N_11828,N_11569,N_11566);
and U11829 (N_11829,N_11560,N_11592);
and U11830 (N_11830,N_11622,N_11698);
nand U11831 (N_11831,N_11589,N_11643);
or U11832 (N_11832,N_11574,N_11683);
nand U11833 (N_11833,N_11654,N_11652);
or U11834 (N_11834,N_11663,N_11566);
or U11835 (N_11835,N_11563,N_11647);
or U11836 (N_11836,N_11618,N_11690);
and U11837 (N_11837,N_11645,N_11683);
and U11838 (N_11838,N_11645,N_11599);
and U11839 (N_11839,N_11654,N_11658);
nor U11840 (N_11840,N_11579,N_11619);
nor U11841 (N_11841,N_11605,N_11555);
nor U11842 (N_11842,N_11648,N_11693);
or U11843 (N_11843,N_11636,N_11696);
nor U11844 (N_11844,N_11679,N_11691);
xor U11845 (N_11845,N_11619,N_11657);
nand U11846 (N_11846,N_11616,N_11576);
or U11847 (N_11847,N_11564,N_11674);
nand U11848 (N_11848,N_11593,N_11659);
and U11849 (N_11849,N_11580,N_11626);
nor U11850 (N_11850,N_11813,N_11715);
and U11851 (N_11851,N_11777,N_11759);
xor U11852 (N_11852,N_11797,N_11744);
nor U11853 (N_11853,N_11749,N_11748);
nor U11854 (N_11854,N_11703,N_11712);
and U11855 (N_11855,N_11783,N_11757);
nor U11856 (N_11856,N_11820,N_11816);
and U11857 (N_11857,N_11745,N_11761);
or U11858 (N_11858,N_11836,N_11730);
nand U11859 (N_11859,N_11723,N_11787);
or U11860 (N_11860,N_11778,N_11746);
or U11861 (N_11861,N_11701,N_11741);
xor U11862 (N_11862,N_11734,N_11831);
nor U11863 (N_11863,N_11768,N_11829);
and U11864 (N_11864,N_11817,N_11824);
nor U11865 (N_11865,N_11789,N_11728);
or U11866 (N_11866,N_11747,N_11733);
and U11867 (N_11867,N_11830,N_11843);
nand U11868 (N_11868,N_11832,N_11835);
nor U11869 (N_11869,N_11839,N_11731);
nor U11870 (N_11870,N_11738,N_11841);
or U11871 (N_11871,N_11785,N_11807);
xor U11872 (N_11872,N_11826,N_11848);
or U11873 (N_11873,N_11794,N_11706);
and U11874 (N_11874,N_11849,N_11709);
nor U11875 (N_11875,N_11795,N_11707);
nor U11876 (N_11876,N_11773,N_11827);
nand U11877 (N_11877,N_11722,N_11729);
or U11878 (N_11878,N_11786,N_11798);
or U11879 (N_11879,N_11705,N_11711);
nand U11880 (N_11880,N_11751,N_11825);
and U11881 (N_11881,N_11803,N_11811);
and U11882 (N_11882,N_11823,N_11846);
and U11883 (N_11883,N_11737,N_11735);
and U11884 (N_11884,N_11790,N_11765);
nand U11885 (N_11885,N_11812,N_11834);
and U11886 (N_11886,N_11847,N_11821);
nor U11887 (N_11887,N_11784,N_11800);
nor U11888 (N_11888,N_11822,N_11718);
and U11889 (N_11889,N_11838,N_11717);
and U11890 (N_11890,N_11774,N_11770);
or U11891 (N_11891,N_11719,N_11810);
or U11892 (N_11892,N_11805,N_11743);
and U11893 (N_11893,N_11842,N_11726);
nor U11894 (N_11894,N_11764,N_11809);
nor U11895 (N_11895,N_11776,N_11742);
and U11896 (N_11896,N_11767,N_11708);
and U11897 (N_11897,N_11775,N_11725);
xnor U11898 (N_11898,N_11771,N_11755);
nor U11899 (N_11899,N_11716,N_11754);
nor U11900 (N_11900,N_11844,N_11721);
nor U11901 (N_11901,N_11801,N_11702);
nand U11902 (N_11902,N_11806,N_11819);
nand U11903 (N_11903,N_11762,N_11796);
nor U11904 (N_11904,N_11840,N_11766);
or U11905 (N_11905,N_11791,N_11780);
nand U11906 (N_11906,N_11740,N_11700);
nand U11907 (N_11907,N_11802,N_11752);
or U11908 (N_11908,N_11753,N_11769);
and U11909 (N_11909,N_11814,N_11837);
xnor U11910 (N_11910,N_11724,N_11760);
nand U11911 (N_11911,N_11845,N_11782);
and U11912 (N_11912,N_11727,N_11714);
xnor U11913 (N_11913,N_11736,N_11704);
nand U11914 (N_11914,N_11710,N_11815);
or U11915 (N_11915,N_11788,N_11756);
and U11916 (N_11916,N_11799,N_11732);
nor U11917 (N_11917,N_11739,N_11720);
nand U11918 (N_11918,N_11750,N_11808);
and U11919 (N_11919,N_11804,N_11772);
xor U11920 (N_11920,N_11763,N_11758);
xnor U11921 (N_11921,N_11781,N_11713);
nand U11922 (N_11922,N_11793,N_11779);
nand U11923 (N_11923,N_11792,N_11833);
nand U11924 (N_11924,N_11828,N_11818);
xor U11925 (N_11925,N_11735,N_11722);
and U11926 (N_11926,N_11802,N_11705);
nand U11927 (N_11927,N_11703,N_11805);
or U11928 (N_11928,N_11762,N_11708);
or U11929 (N_11929,N_11731,N_11767);
nor U11930 (N_11930,N_11713,N_11715);
nor U11931 (N_11931,N_11843,N_11817);
nand U11932 (N_11932,N_11767,N_11733);
xnor U11933 (N_11933,N_11705,N_11728);
and U11934 (N_11934,N_11768,N_11717);
nand U11935 (N_11935,N_11738,N_11703);
nor U11936 (N_11936,N_11818,N_11732);
and U11937 (N_11937,N_11741,N_11803);
nor U11938 (N_11938,N_11794,N_11826);
nor U11939 (N_11939,N_11846,N_11797);
or U11940 (N_11940,N_11817,N_11840);
nor U11941 (N_11941,N_11704,N_11775);
or U11942 (N_11942,N_11745,N_11787);
nor U11943 (N_11943,N_11803,N_11740);
nand U11944 (N_11944,N_11809,N_11771);
nor U11945 (N_11945,N_11758,N_11735);
nor U11946 (N_11946,N_11824,N_11828);
nor U11947 (N_11947,N_11791,N_11823);
or U11948 (N_11948,N_11770,N_11847);
and U11949 (N_11949,N_11753,N_11782);
nand U11950 (N_11950,N_11847,N_11749);
nor U11951 (N_11951,N_11827,N_11803);
and U11952 (N_11952,N_11755,N_11700);
nor U11953 (N_11953,N_11825,N_11842);
nand U11954 (N_11954,N_11755,N_11820);
xnor U11955 (N_11955,N_11768,N_11718);
xnor U11956 (N_11956,N_11725,N_11791);
nand U11957 (N_11957,N_11754,N_11773);
and U11958 (N_11958,N_11731,N_11813);
or U11959 (N_11959,N_11815,N_11706);
and U11960 (N_11960,N_11790,N_11744);
nor U11961 (N_11961,N_11811,N_11703);
or U11962 (N_11962,N_11789,N_11829);
nor U11963 (N_11963,N_11832,N_11768);
nand U11964 (N_11964,N_11820,N_11718);
and U11965 (N_11965,N_11756,N_11737);
xnor U11966 (N_11966,N_11808,N_11805);
nand U11967 (N_11967,N_11723,N_11733);
or U11968 (N_11968,N_11812,N_11824);
nor U11969 (N_11969,N_11742,N_11814);
or U11970 (N_11970,N_11753,N_11813);
nor U11971 (N_11971,N_11772,N_11757);
and U11972 (N_11972,N_11828,N_11735);
and U11973 (N_11973,N_11774,N_11808);
and U11974 (N_11974,N_11829,N_11760);
xor U11975 (N_11975,N_11794,N_11792);
and U11976 (N_11976,N_11836,N_11837);
and U11977 (N_11977,N_11726,N_11767);
or U11978 (N_11978,N_11714,N_11706);
nand U11979 (N_11979,N_11830,N_11815);
xnor U11980 (N_11980,N_11785,N_11702);
nand U11981 (N_11981,N_11753,N_11787);
and U11982 (N_11982,N_11709,N_11741);
nor U11983 (N_11983,N_11751,N_11813);
nand U11984 (N_11984,N_11841,N_11832);
nor U11985 (N_11985,N_11716,N_11791);
and U11986 (N_11986,N_11813,N_11704);
nand U11987 (N_11987,N_11820,N_11722);
or U11988 (N_11988,N_11790,N_11734);
and U11989 (N_11989,N_11806,N_11720);
xnor U11990 (N_11990,N_11796,N_11706);
nand U11991 (N_11991,N_11824,N_11728);
or U11992 (N_11992,N_11778,N_11743);
nand U11993 (N_11993,N_11801,N_11779);
or U11994 (N_11994,N_11738,N_11727);
nor U11995 (N_11995,N_11803,N_11822);
or U11996 (N_11996,N_11735,N_11745);
or U11997 (N_11997,N_11700,N_11769);
nand U11998 (N_11998,N_11776,N_11753);
nand U11999 (N_11999,N_11846,N_11781);
or U12000 (N_12000,N_11860,N_11975);
or U12001 (N_12001,N_11919,N_11897);
nor U12002 (N_12002,N_11889,N_11993);
nand U12003 (N_12003,N_11969,N_11998);
and U12004 (N_12004,N_11927,N_11955);
and U12005 (N_12005,N_11922,N_11950);
xor U12006 (N_12006,N_11946,N_11866);
nand U12007 (N_12007,N_11994,N_11882);
nor U12008 (N_12008,N_11964,N_11872);
nand U12009 (N_12009,N_11990,N_11989);
nand U12010 (N_12010,N_11867,N_11907);
nand U12011 (N_12011,N_11985,N_11931);
and U12012 (N_12012,N_11963,N_11874);
and U12013 (N_12013,N_11906,N_11914);
or U12014 (N_12014,N_11978,N_11908);
and U12015 (N_12015,N_11999,N_11968);
and U12016 (N_12016,N_11971,N_11984);
xor U12017 (N_12017,N_11869,N_11979);
xor U12018 (N_12018,N_11970,N_11851);
or U12019 (N_12019,N_11965,N_11988);
or U12020 (N_12020,N_11932,N_11953);
nor U12021 (N_12021,N_11992,N_11973);
nand U12022 (N_12022,N_11996,N_11977);
nand U12023 (N_12023,N_11859,N_11972);
or U12024 (N_12024,N_11890,N_11921);
and U12025 (N_12025,N_11938,N_11850);
nand U12026 (N_12026,N_11949,N_11870);
and U12027 (N_12027,N_11960,N_11920);
and U12028 (N_12028,N_11959,N_11934);
nor U12029 (N_12029,N_11944,N_11913);
or U12030 (N_12030,N_11967,N_11982);
or U12031 (N_12031,N_11986,N_11974);
or U12032 (N_12032,N_11943,N_11864);
or U12033 (N_12033,N_11935,N_11905);
and U12034 (N_12034,N_11853,N_11954);
xor U12035 (N_12035,N_11856,N_11880);
nor U12036 (N_12036,N_11981,N_11892);
and U12037 (N_12037,N_11879,N_11854);
nand U12038 (N_12038,N_11912,N_11951);
or U12039 (N_12039,N_11862,N_11858);
or U12040 (N_12040,N_11885,N_11895);
nor U12041 (N_12041,N_11875,N_11857);
nand U12042 (N_12042,N_11861,N_11909);
nand U12043 (N_12043,N_11942,N_11936);
nand U12044 (N_12044,N_11940,N_11991);
xor U12045 (N_12045,N_11997,N_11980);
nand U12046 (N_12046,N_11983,N_11995);
or U12047 (N_12047,N_11899,N_11900);
nand U12048 (N_12048,N_11947,N_11952);
and U12049 (N_12049,N_11930,N_11976);
and U12050 (N_12050,N_11877,N_11911);
and U12051 (N_12051,N_11956,N_11902);
and U12052 (N_12052,N_11966,N_11884);
and U12053 (N_12053,N_11893,N_11987);
nor U12054 (N_12054,N_11915,N_11852);
nand U12055 (N_12055,N_11863,N_11876);
and U12056 (N_12056,N_11894,N_11888);
xor U12057 (N_12057,N_11939,N_11945);
nor U12058 (N_12058,N_11933,N_11962);
nor U12059 (N_12059,N_11957,N_11941);
nor U12060 (N_12060,N_11898,N_11948);
nand U12061 (N_12061,N_11928,N_11958);
or U12062 (N_12062,N_11926,N_11917);
nor U12063 (N_12063,N_11881,N_11887);
and U12064 (N_12064,N_11855,N_11865);
or U12065 (N_12065,N_11871,N_11937);
nor U12066 (N_12066,N_11923,N_11886);
and U12067 (N_12067,N_11873,N_11901);
and U12068 (N_12068,N_11878,N_11891);
nand U12069 (N_12069,N_11961,N_11903);
nor U12070 (N_12070,N_11924,N_11916);
or U12071 (N_12071,N_11883,N_11929);
nor U12072 (N_12072,N_11904,N_11896);
nand U12073 (N_12073,N_11925,N_11868);
nor U12074 (N_12074,N_11918,N_11910);
xnor U12075 (N_12075,N_11995,N_11888);
nor U12076 (N_12076,N_11935,N_11917);
or U12077 (N_12077,N_11944,N_11992);
and U12078 (N_12078,N_11910,N_11928);
nor U12079 (N_12079,N_11972,N_11994);
nand U12080 (N_12080,N_11977,N_11895);
or U12081 (N_12081,N_11925,N_11890);
nand U12082 (N_12082,N_11919,N_11978);
and U12083 (N_12083,N_11930,N_11967);
xor U12084 (N_12084,N_11867,N_11992);
and U12085 (N_12085,N_11945,N_11904);
and U12086 (N_12086,N_11998,N_11924);
xor U12087 (N_12087,N_11979,N_11937);
nand U12088 (N_12088,N_11947,N_11945);
or U12089 (N_12089,N_11944,N_11901);
nor U12090 (N_12090,N_11852,N_11880);
nand U12091 (N_12091,N_11961,N_11922);
nand U12092 (N_12092,N_11939,N_11919);
nand U12093 (N_12093,N_11955,N_11922);
xor U12094 (N_12094,N_11996,N_11919);
xnor U12095 (N_12095,N_11984,N_11906);
and U12096 (N_12096,N_11977,N_11984);
nor U12097 (N_12097,N_11868,N_11934);
nor U12098 (N_12098,N_11983,N_11963);
xnor U12099 (N_12099,N_11890,N_11983);
nor U12100 (N_12100,N_11852,N_11868);
xnor U12101 (N_12101,N_11852,N_11924);
nand U12102 (N_12102,N_11998,N_11915);
nor U12103 (N_12103,N_11999,N_11904);
or U12104 (N_12104,N_11931,N_11944);
xnor U12105 (N_12105,N_11934,N_11914);
or U12106 (N_12106,N_11986,N_11914);
nor U12107 (N_12107,N_11896,N_11997);
and U12108 (N_12108,N_11890,N_11871);
nor U12109 (N_12109,N_11914,N_11963);
nand U12110 (N_12110,N_11952,N_11983);
nand U12111 (N_12111,N_11869,N_11946);
nand U12112 (N_12112,N_11850,N_11992);
nand U12113 (N_12113,N_11899,N_11999);
nand U12114 (N_12114,N_11947,N_11961);
nand U12115 (N_12115,N_11933,N_11939);
nand U12116 (N_12116,N_11871,N_11944);
nor U12117 (N_12117,N_11921,N_11919);
nand U12118 (N_12118,N_11981,N_11883);
xor U12119 (N_12119,N_11920,N_11953);
nand U12120 (N_12120,N_11880,N_11858);
nor U12121 (N_12121,N_11970,N_11927);
or U12122 (N_12122,N_11934,N_11875);
and U12123 (N_12123,N_11901,N_11864);
xnor U12124 (N_12124,N_11979,N_11885);
nand U12125 (N_12125,N_11969,N_11999);
nand U12126 (N_12126,N_11850,N_11961);
and U12127 (N_12127,N_11926,N_11937);
nor U12128 (N_12128,N_11890,N_11956);
or U12129 (N_12129,N_11890,N_11987);
or U12130 (N_12130,N_11881,N_11985);
nor U12131 (N_12131,N_11956,N_11979);
or U12132 (N_12132,N_11945,N_11899);
nand U12133 (N_12133,N_11921,N_11988);
and U12134 (N_12134,N_11976,N_11911);
or U12135 (N_12135,N_11947,N_11873);
xnor U12136 (N_12136,N_11901,N_11921);
or U12137 (N_12137,N_11891,N_11885);
nor U12138 (N_12138,N_11875,N_11886);
and U12139 (N_12139,N_11918,N_11892);
nand U12140 (N_12140,N_11927,N_11999);
xor U12141 (N_12141,N_11938,N_11996);
xnor U12142 (N_12142,N_11851,N_11999);
and U12143 (N_12143,N_11943,N_11859);
or U12144 (N_12144,N_11947,N_11915);
nand U12145 (N_12145,N_11996,N_11969);
nor U12146 (N_12146,N_11904,N_11880);
xor U12147 (N_12147,N_11853,N_11964);
nor U12148 (N_12148,N_11889,N_11945);
or U12149 (N_12149,N_11936,N_11993);
nand U12150 (N_12150,N_12047,N_12124);
or U12151 (N_12151,N_12028,N_12078);
nor U12152 (N_12152,N_12116,N_12013);
xnor U12153 (N_12153,N_12121,N_12147);
xor U12154 (N_12154,N_12072,N_12042);
xor U12155 (N_12155,N_12085,N_12045);
nand U12156 (N_12156,N_12083,N_12105);
xor U12157 (N_12157,N_12025,N_12104);
and U12158 (N_12158,N_12034,N_12031);
nand U12159 (N_12159,N_12090,N_12016);
and U12160 (N_12160,N_12117,N_12055);
nor U12161 (N_12161,N_12046,N_12009);
nand U12162 (N_12162,N_12026,N_12063);
and U12163 (N_12163,N_12077,N_12087);
and U12164 (N_12164,N_12021,N_12107);
and U12165 (N_12165,N_12128,N_12136);
nand U12166 (N_12166,N_12129,N_12109);
nor U12167 (N_12167,N_12007,N_12041);
or U12168 (N_12168,N_12050,N_12066);
xnor U12169 (N_12169,N_12131,N_12029);
nand U12170 (N_12170,N_12056,N_12126);
nand U12171 (N_12171,N_12108,N_12100);
xor U12172 (N_12172,N_12118,N_12122);
xor U12173 (N_12173,N_12082,N_12096);
and U12174 (N_12174,N_12140,N_12127);
and U12175 (N_12175,N_12142,N_12064);
nand U12176 (N_12176,N_12114,N_12018);
xnor U12177 (N_12177,N_12032,N_12070);
or U12178 (N_12178,N_12051,N_12098);
nor U12179 (N_12179,N_12125,N_12111);
and U12180 (N_12180,N_12065,N_12054);
nor U12181 (N_12181,N_12020,N_12033);
xor U12182 (N_12182,N_12091,N_12001);
or U12183 (N_12183,N_12086,N_12134);
nor U12184 (N_12184,N_12141,N_12052);
and U12185 (N_12185,N_12068,N_12004);
xor U12186 (N_12186,N_12071,N_12089);
nor U12187 (N_12187,N_12076,N_12097);
and U12188 (N_12188,N_12137,N_12144);
nand U12189 (N_12189,N_12138,N_12080);
xor U12190 (N_12190,N_12048,N_12035);
and U12191 (N_12191,N_12123,N_12120);
xor U12192 (N_12192,N_12103,N_12084);
and U12193 (N_12193,N_12060,N_12119);
nand U12194 (N_12194,N_12106,N_12081);
or U12195 (N_12195,N_12073,N_12102);
xor U12196 (N_12196,N_12133,N_12139);
and U12197 (N_12197,N_12015,N_12115);
and U12198 (N_12198,N_12059,N_12075);
and U12199 (N_12199,N_12130,N_12093);
nor U12200 (N_12200,N_12095,N_12146);
nor U12201 (N_12201,N_12074,N_12010);
nand U12202 (N_12202,N_12053,N_12069);
nand U12203 (N_12203,N_12002,N_12088);
nor U12204 (N_12204,N_12043,N_12143);
and U12205 (N_12205,N_12017,N_12058);
nor U12206 (N_12206,N_12145,N_12148);
nand U12207 (N_12207,N_12039,N_12019);
or U12208 (N_12208,N_12044,N_12040);
nand U12209 (N_12209,N_12110,N_12000);
nand U12210 (N_12210,N_12049,N_12024);
and U12211 (N_12211,N_12062,N_12061);
and U12212 (N_12212,N_12135,N_12038);
or U12213 (N_12213,N_12112,N_12057);
nand U12214 (N_12214,N_12030,N_12036);
and U12215 (N_12215,N_12094,N_12037);
and U12216 (N_12216,N_12132,N_12003);
nand U12217 (N_12217,N_12022,N_12005);
nor U12218 (N_12218,N_12012,N_12113);
nand U12219 (N_12219,N_12023,N_12101);
nand U12220 (N_12220,N_12099,N_12092);
nand U12221 (N_12221,N_12011,N_12006);
and U12222 (N_12222,N_12079,N_12067);
and U12223 (N_12223,N_12027,N_12149);
nand U12224 (N_12224,N_12014,N_12008);
nor U12225 (N_12225,N_12068,N_12031);
nand U12226 (N_12226,N_12076,N_12012);
and U12227 (N_12227,N_12029,N_12053);
and U12228 (N_12228,N_12132,N_12022);
xor U12229 (N_12229,N_12095,N_12106);
nor U12230 (N_12230,N_12045,N_12080);
and U12231 (N_12231,N_12127,N_12021);
nor U12232 (N_12232,N_12110,N_12133);
and U12233 (N_12233,N_12143,N_12010);
nand U12234 (N_12234,N_12046,N_12059);
nand U12235 (N_12235,N_12066,N_12004);
and U12236 (N_12236,N_12014,N_12145);
nand U12237 (N_12237,N_12057,N_12140);
or U12238 (N_12238,N_12101,N_12140);
or U12239 (N_12239,N_12038,N_12007);
nor U12240 (N_12240,N_12147,N_12118);
nand U12241 (N_12241,N_12138,N_12145);
and U12242 (N_12242,N_12133,N_12042);
nor U12243 (N_12243,N_12090,N_12080);
xor U12244 (N_12244,N_12060,N_12088);
or U12245 (N_12245,N_12115,N_12008);
nand U12246 (N_12246,N_12037,N_12033);
nand U12247 (N_12247,N_12128,N_12001);
nand U12248 (N_12248,N_12075,N_12083);
and U12249 (N_12249,N_12023,N_12088);
nor U12250 (N_12250,N_12142,N_12117);
nor U12251 (N_12251,N_12113,N_12064);
xnor U12252 (N_12252,N_12019,N_12043);
and U12253 (N_12253,N_12082,N_12103);
nor U12254 (N_12254,N_12035,N_12096);
or U12255 (N_12255,N_12096,N_12097);
nor U12256 (N_12256,N_12067,N_12062);
nor U12257 (N_12257,N_12138,N_12101);
xnor U12258 (N_12258,N_12022,N_12122);
and U12259 (N_12259,N_12147,N_12081);
or U12260 (N_12260,N_12147,N_12073);
nand U12261 (N_12261,N_12115,N_12093);
or U12262 (N_12262,N_12063,N_12028);
nor U12263 (N_12263,N_12097,N_12112);
and U12264 (N_12264,N_12014,N_12051);
xor U12265 (N_12265,N_12057,N_12050);
nand U12266 (N_12266,N_12064,N_12128);
nand U12267 (N_12267,N_12068,N_12067);
nand U12268 (N_12268,N_12056,N_12038);
nor U12269 (N_12269,N_12025,N_12034);
and U12270 (N_12270,N_12138,N_12016);
nor U12271 (N_12271,N_12080,N_12141);
nand U12272 (N_12272,N_12047,N_12114);
and U12273 (N_12273,N_12007,N_12141);
or U12274 (N_12274,N_12110,N_12091);
and U12275 (N_12275,N_12149,N_12077);
or U12276 (N_12276,N_12113,N_12051);
nand U12277 (N_12277,N_12006,N_12143);
nor U12278 (N_12278,N_12040,N_12120);
nor U12279 (N_12279,N_12138,N_12123);
nand U12280 (N_12280,N_12137,N_12028);
and U12281 (N_12281,N_12057,N_12105);
xnor U12282 (N_12282,N_12065,N_12001);
and U12283 (N_12283,N_12087,N_12144);
nor U12284 (N_12284,N_12132,N_12130);
or U12285 (N_12285,N_12031,N_12088);
nand U12286 (N_12286,N_12136,N_12026);
nand U12287 (N_12287,N_12112,N_12134);
or U12288 (N_12288,N_12107,N_12058);
and U12289 (N_12289,N_12064,N_12141);
nand U12290 (N_12290,N_12090,N_12038);
or U12291 (N_12291,N_12029,N_12115);
nand U12292 (N_12292,N_12013,N_12117);
or U12293 (N_12293,N_12084,N_12028);
or U12294 (N_12294,N_12119,N_12090);
xnor U12295 (N_12295,N_12096,N_12022);
or U12296 (N_12296,N_12016,N_12142);
and U12297 (N_12297,N_12083,N_12057);
and U12298 (N_12298,N_12067,N_12119);
nand U12299 (N_12299,N_12092,N_12012);
and U12300 (N_12300,N_12171,N_12293);
nand U12301 (N_12301,N_12284,N_12223);
nand U12302 (N_12302,N_12162,N_12181);
and U12303 (N_12303,N_12286,N_12177);
nor U12304 (N_12304,N_12267,N_12192);
nor U12305 (N_12305,N_12174,N_12282);
nand U12306 (N_12306,N_12152,N_12239);
nand U12307 (N_12307,N_12250,N_12194);
or U12308 (N_12308,N_12243,N_12206);
nor U12309 (N_12309,N_12288,N_12165);
and U12310 (N_12310,N_12270,N_12185);
nor U12311 (N_12311,N_12246,N_12207);
or U12312 (N_12312,N_12274,N_12178);
and U12313 (N_12313,N_12179,N_12285);
nand U12314 (N_12314,N_12297,N_12222);
xor U12315 (N_12315,N_12220,N_12264);
nand U12316 (N_12316,N_12216,N_12299);
and U12317 (N_12317,N_12217,N_12227);
nor U12318 (N_12318,N_12164,N_12235);
nor U12319 (N_12319,N_12200,N_12189);
and U12320 (N_12320,N_12266,N_12191);
and U12321 (N_12321,N_12158,N_12218);
nor U12322 (N_12322,N_12213,N_12225);
nand U12323 (N_12323,N_12224,N_12298);
and U12324 (N_12324,N_12255,N_12170);
nand U12325 (N_12325,N_12219,N_12184);
and U12326 (N_12326,N_12245,N_12168);
nand U12327 (N_12327,N_12161,N_12252);
nand U12328 (N_12328,N_12268,N_12287);
or U12329 (N_12329,N_12229,N_12249);
or U12330 (N_12330,N_12291,N_12237);
and U12331 (N_12331,N_12160,N_12241);
or U12332 (N_12332,N_12190,N_12151);
and U12333 (N_12333,N_12197,N_12154);
nand U12334 (N_12334,N_12281,N_12155);
nand U12335 (N_12335,N_12230,N_12240);
xor U12336 (N_12336,N_12188,N_12159);
nor U12337 (N_12337,N_12166,N_12261);
or U12338 (N_12338,N_12257,N_12163);
or U12339 (N_12339,N_12279,N_12262);
nor U12340 (N_12340,N_12292,N_12153);
nand U12341 (N_12341,N_12272,N_12269);
nor U12342 (N_12342,N_12254,N_12228);
nand U12343 (N_12343,N_12290,N_12209);
nand U12344 (N_12344,N_12199,N_12195);
or U12345 (N_12345,N_12294,N_12221);
or U12346 (N_12346,N_12212,N_12280);
xor U12347 (N_12347,N_12242,N_12296);
nand U12348 (N_12348,N_12258,N_12289);
nor U12349 (N_12349,N_12182,N_12201);
or U12350 (N_12350,N_12278,N_12295);
nor U12351 (N_12351,N_12202,N_12283);
or U12352 (N_12352,N_12208,N_12231);
nand U12353 (N_12353,N_12205,N_12210);
nand U12354 (N_12354,N_12172,N_12193);
xnor U12355 (N_12355,N_12175,N_12263);
and U12356 (N_12356,N_12183,N_12180);
nand U12357 (N_12357,N_12238,N_12157);
or U12358 (N_12358,N_12214,N_12253);
or U12359 (N_12359,N_12271,N_12204);
xor U12360 (N_12360,N_12232,N_12156);
and U12361 (N_12361,N_12276,N_12215);
nand U12362 (N_12362,N_12196,N_12167);
or U12363 (N_12363,N_12256,N_12173);
or U12364 (N_12364,N_12273,N_12150);
nand U12365 (N_12365,N_12248,N_12169);
nand U12366 (N_12366,N_12247,N_12203);
nor U12367 (N_12367,N_12176,N_12275);
nand U12368 (N_12368,N_12277,N_12236);
or U12369 (N_12369,N_12251,N_12211);
nor U12370 (N_12370,N_12234,N_12226);
nand U12371 (N_12371,N_12244,N_12265);
nor U12372 (N_12372,N_12186,N_12198);
nor U12373 (N_12373,N_12187,N_12260);
or U12374 (N_12374,N_12259,N_12233);
nor U12375 (N_12375,N_12219,N_12251);
and U12376 (N_12376,N_12249,N_12272);
xnor U12377 (N_12377,N_12233,N_12290);
and U12378 (N_12378,N_12284,N_12214);
or U12379 (N_12379,N_12165,N_12245);
or U12380 (N_12380,N_12245,N_12196);
nand U12381 (N_12381,N_12248,N_12178);
or U12382 (N_12382,N_12162,N_12211);
xnor U12383 (N_12383,N_12211,N_12180);
nor U12384 (N_12384,N_12163,N_12282);
nand U12385 (N_12385,N_12207,N_12270);
nand U12386 (N_12386,N_12227,N_12160);
nor U12387 (N_12387,N_12291,N_12153);
or U12388 (N_12388,N_12165,N_12218);
nor U12389 (N_12389,N_12186,N_12285);
and U12390 (N_12390,N_12294,N_12199);
nand U12391 (N_12391,N_12263,N_12226);
nand U12392 (N_12392,N_12182,N_12203);
and U12393 (N_12393,N_12177,N_12163);
and U12394 (N_12394,N_12286,N_12160);
nor U12395 (N_12395,N_12162,N_12270);
nand U12396 (N_12396,N_12193,N_12205);
and U12397 (N_12397,N_12179,N_12222);
nand U12398 (N_12398,N_12222,N_12159);
nor U12399 (N_12399,N_12284,N_12183);
nand U12400 (N_12400,N_12295,N_12150);
xor U12401 (N_12401,N_12248,N_12162);
nor U12402 (N_12402,N_12230,N_12223);
or U12403 (N_12403,N_12198,N_12253);
nor U12404 (N_12404,N_12215,N_12177);
nor U12405 (N_12405,N_12194,N_12174);
or U12406 (N_12406,N_12173,N_12198);
nor U12407 (N_12407,N_12187,N_12172);
or U12408 (N_12408,N_12279,N_12201);
and U12409 (N_12409,N_12153,N_12195);
nor U12410 (N_12410,N_12230,N_12201);
and U12411 (N_12411,N_12271,N_12287);
nor U12412 (N_12412,N_12164,N_12236);
nand U12413 (N_12413,N_12264,N_12246);
nor U12414 (N_12414,N_12212,N_12285);
xnor U12415 (N_12415,N_12267,N_12295);
nand U12416 (N_12416,N_12254,N_12173);
or U12417 (N_12417,N_12241,N_12196);
nor U12418 (N_12418,N_12238,N_12231);
or U12419 (N_12419,N_12208,N_12243);
or U12420 (N_12420,N_12241,N_12207);
nand U12421 (N_12421,N_12176,N_12193);
and U12422 (N_12422,N_12182,N_12246);
and U12423 (N_12423,N_12280,N_12221);
nor U12424 (N_12424,N_12258,N_12167);
nor U12425 (N_12425,N_12180,N_12258);
nand U12426 (N_12426,N_12267,N_12166);
and U12427 (N_12427,N_12279,N_12230);
xnor U12428 (N_12428,N_12204,N_12226);
xnor U12429 (N_12429,N_12175,N_12286);
and U12430 (N_12430,N_12254,N_12225);
nor U12431 (N_12431,N_12185,N_12239);
nand U12432 (N_12432,N_12237,N_12156);
or U12433 (N_12433,N_12211,N_12288);
nor U12434 (N_12434,N_12211,N_12274);
xnor U12435 (N_12435,N_12273,N_12215);
and U12436 (N_12436,N_12275,N_12209);
nor U12437 (N_12437,N_12201,N_12274);
and U12438 (N_12438,N_12232,N_12234);
or U12439 (N_12439,N_12271,N_12189);
nor U12440 (N_12440,N_12254,N_12274);
nand U12441 (N_12441,N_12291,N_12198);
nand U12442 (N_12442,N_12169,N_12244);
or U12443 (N_12443,N_12207,N_12279);
and U12444 (N_12444,N_12208,N_12278);
nor U12445 (N_12445,N_12227,N_12274);
nand U12446 (N_12446,N_12263,N_12156);
and U12447 (N_12447,N_12190,N_12223);
nand U12448 (N_12448,N_12164,N_12279);
and U12449 (N_12449,N_12221,N_12283);
nor U12450 (N_12450,N_12350,N_12442);
nor U12451 (N_12451,N_12354,N_12334);
or U12452 (N_12452,N_12411,N_12312);
nor U12453 (N_12453,N_12348,N_12340);
nor U12454 (N_12454,N_12316,N_12445);
xnor U12455 (N_12455,N_12349,N_12372);
or U12456 (N_12456,N_12380,N_12434);
or U12457 (N_12457,N_12359,N_12381);
nor U12458 (N_12458,N_12443,N_12362);
nor U12459 (N_12459,N_12426,N_12429);
nand U12460 (N_12460,N_12424,N_12325);
nand U12461 (N_12461,N_12422,N_12369);
and U12462 (N_12462,N_12378,N_12310);
or U12463 (N_12463,N_12315,N_12421);
nor U12464 (N_12464,N_12430,N_12416);
or U12465 (N_12465,N_12387,N_12368);
nand U12466 (N_12466,N_12399,N_12337);
nor U12467 (N_12467,N_12413,N_12400);
and U12468 (N_12468,N_12360,N_12447);
or U12469 (N_12469,N_12420,N_12365);
or U12470 (N_12470,N_12355,N_12393);
and U12471 (N_12471,N_12409,N_12407);
nand U12472 (N_12472,N_12376,N_12335);
nor U12473 (N_12473,N_12302,N_12389);
and U12474 (N_12474,N_12308,N_12404);
nor U12475 (N_12475,N_12383,N_12345);
nand U12476 (N_12476,N_12336,N_12436);
or U12477 (N_12477,N_12382,N_12344);
nor U12478 (N_12478,N_12401,N_12437);
nor U12479 (N_12479,N_12391,N_12419);
nor U12480 (N_12480,N_12343,N_12415);
nand U12481 (N_12481,N_12448,N_12338);
nand U12482 (N_12482,N_12300,N_12398);
or U12483 (N_12483,N_12418,N_12386);
and U12484 (N_12484,N_12402,N_12446);
and U12485 (N_12485,N_12331,N_12326);
nand U12486 (N_12486,N_12414,N_12439);
or U12487 (N_12487,N_12395,N_12431);
nand U12488 (N_12488,N_12396,N_12384);
and U12489 (N_12489,N_12352,N_12367);
xor U12490 (N_12490,N_12324,N_12363);
nand U12491 (N_12491,N_12394,N_12390);
nor U12492 (N_12492,N_12423,N_12449);
nor U12493 (N_12493,N_12427,N_12327);
nor U12494 (N_12494,N_12317,N_12309);
nor U12495 (N_12495,N_12403,N_12332);
or U12496 (N_12496,N_12371,N_12373);
nand U12497 (N_12497,N_12346,N_12375);
nand U12498 (N_12498,N_12441,N_12339);
nand U12499 (N_12499,N_12412,N_12307);
or U12500 (N_12500,N_12330,N_12320);
nor U12501 (N_12501,N_12356,N_12314);
xnor U12502 (N_12502,N_12374,N_12385);
nand U12503 (N_12503,N_12318,N_12392);
nor U12504 (N_12504,N_12342,N_12388);
nor U12505 (N_12505,N_12329,N_12311);
xor U12506 (N_12506,N_12432,N_12319);
and U12507 (N_12507,N_12306,N_12438);
nor U12508 (N_12508,N_12333,N_12444);
nand U12509 (N_12509,N_12433,N_12364);
and U12510 (N_12510,N_12397,N_12305);
or U12511 (N_12511,N_12301,N_12353);
xnor U12512 (N_12512,N_12357,N_12366);
nor U12513 (N_12513,N_12428,N_12370);
nand U12514 (N_12514,N_12321,N_12410);
and U12515 (N_12515,N_12303,N_12408);
and U12516 (N_12516,N_12440,N_12406);
and U12517 (N_12517,N_12341,N_12435);
or U12518 (N_12518,N_12405,N_12361);
xor U12519 (N_12519,N_12358,N_12304);
or U12520 (N_12520,N_12351,N_12323);
or U12521 (N_12521,N_12417,N_12347);
or U12522 (N_12522,N_12425,N_12328);
nor U12523 (N_12523,N_12377,N_12313);
nand U12524 (N_12524,N_12322,N_12379);
and U12525 (N_12525,N_12313,N_12366);
and U12526 (N_12526,N_12345,N_12350);
nand U12527 (N_12527,N_12319,N_12429);
nand U12528 (N_12528,N_12426,N_12380);
nand U12529 (N_12529,N_12378,N_12305);
nor U12530 (N_12530,N_12361,N_12364);
or U12531 (N_12531,N_12354,N_12387);
nand U12532 (N_12532,N_12415,N_12352);
or U12533 (N_12533,N_12425,N_12448);
nand U12534 (N_12534,N_12427,N_12384);
or U12535 (N_12535,N_12404,N_12414);
or U12536 (N_12536,N_12432,N_12436);
and U12537 (N_12537,N_12361,N_12339);
or U12538 (N_12538,N_12340,N_12362);
nand U12539 (N_12539,N_12384,N_12319);
and U12540 (N_12540,N_12422,N_12364);
nand U12541 (N_12541,N_12346,N_12391);
nand U12542 (N_12542,N_12365,N_12350);
nand U12543 (N_12543,N_12446,N_12393);
or U12544 (N_12544,N_12397,N_12387);
xor U12545 (N_12545,N_12308,N_12439);
nor U12546 (N_12546,N_12387,N_12303);
or U12547 (N_12547,N_12431,N_12416);
and U12548 (N_12548,N_12364,N_12395);
xnor U12549 (N_12549,N_12357,N_12303);
and U12550 (N_12550,N_12426,N_12306);
or U12551 (N_12551,N_12312,N_12394);
and U12552 (N_12552,N_12365,N_12339);
nor U12553 (N_12553,N_12419,N_12351);
nor U12554 (N_12554,N_12317,N_12327);
nor U12555 (N_12555,N_12426,N_12349);
nand U12556 (N_12556,N_12394,N_12435);
xnor U12557 (N_12557,N_12422,N_12372);
or U12558 (N_12558,N_12309,N_12400);
or U12559 (N_12559,N_12445,N_12350);
or U12560 (N_12560,N_12438,N_12414);
nand U12561 (N_12561,N_12401,N_12342);
nand U12562 (N_12562,N_12417,N_12415);
or U12563 (N_12563,N_12406,N_12340);
or U12564 (N_12564,N_12442,N_12420);
or U12565 (N_12565,N_12330,N_12369);
or U12566 (N_12566,N_12399,N_12448);
nand U12567 (N_12567,N_12318,N_12442);
and U12568 (N_12568,N_12446,N_12335);
nor U12569 (N_12569,N_12309,N_12416);
nor U12570 (N_12570,N_12443,N_12407);
nand U12571 (N_12571,N_12374,N_12333);
nand U12572 (N_12572,N_12396,N_12445);
or U12573 (N_12573,N_12322,N_12366);
nand U12574 (N_12574,N_12420,N_12385);
nor U12575 (N_12575,N_12357,N_12365);
xor U12576 (N_12576,N_12324,N_12360);
and U12577 (N_12577,N_12399,N_12394);
nor U12578 (N_12578,N_12375,N_12404);
and U12579 (N_12579,N_12346,N_12395);
and U12580 (N_12580,N_12392,N_12343);
nand U12581 (N_12581,N_12314,N_12403);
or U12582 (N_12582,N_12386,N_12416);
or U12583 (N_12583,N_12387,N_12312);
nor U12584 (N_12584,N_12321,N_12324);
and U12585 (N_12585,N_12341,N_12306);
nor U12586 (N_12586,N_12428,N_12433);
or U12587 (N_12587,N_12330,N_12371);
and U12588 (N_12588,N_12307,N_12431);
nand U12589 (N_12589,N_12345,N_12369);
nand U12590 (N_12590,N_12317,N_12389);
or U12591 (N_12591,N_12405,N_12403);
and U12592 (N_12592,N_12395,N_12415);
nand U12593 (N_12593,N_12301,N_12418);
nor U12594 (N_12594,N_12353,N_12388);
nand U12595 (N_12595,N_12319,N_12404);
nand U12596 (N_12596,N_12350,N_12300);
or U12597 (N_12597,N_12331,N_12384);
xnor U12598 (N_12598,N_12307,N_12340);
xor U12599 (N_12599,N_12404,N_12311);
nor U12600 (N_12600,N_12476,N_12511);
xor U12601 (N_12601,N_12564,N_12531);
and U12602 (N_12602,N_12575,N_12493);
nand U12603 (N_12603,N_12462,N_12507);
or U12604 (N_12604,N_12577,N_12563);
xor U12605 (N_12605,N_12571,N_12463);
and U12606 (N_12606,N_12516,N_12514);
nor U12607 (N_12607,N_12509,N_12555);
or U12608 (N_12608,N_12484,N_12473);
nor U12609 (N_12609,N_12537,N_12482);
or U12610 (N_12610,N_12512,N_12536);
nor U12611 (N_12611,N_12456,N_12502);
and U12612 (N_12612,N_12595,N_12508);
nor U12613 (N_12613,N_12561,N_12539);
nor U12614 (N_12614,N_12573,N_12542);
and U12615 (N_12615,N_12551,N_12547);
nor U12616 (N_12616,N_12568,N_12597);
or U12617 (N_12617,N_12584,N_12469);
nor U12618 (N_12618,N_12591,N_12501);
nor U12619 (N_12619,N_12588,N_12500);
nand U12620 (N_12620,N_12593,N_12479);
nor U12621 (N_12621,N_12465,N_12589);
nor U12622 (N_12622,N_12454,N_12585);
xnor U12623 (N_12623,N_12517,N_12590);
and U12624 (N_12624,N_12552,N_12594);
or U12625 (N_12625,N_12540,N_12504);
nand U12626 (N_12626,N_12578,N_12560);
or U12627 (N_12627,N_12579,N_12467);
and U12628 (N_12628,N_12523,N_12475);
nand U12629 (N_12629,N_12529,N_12474);
nor U12630 (N_12630,N_12544,N_12567);
xor U12631 (N_12631,N_12470,N_12553);
or U12632 (N_12632,N_12535,N_12580);
nand U12633 (N_12633,N_12581,N_12489);
nor U12634 (N_12634,N_12554,N_12486);
nor U12635 (N_12635,N_12520,N_12570);
nor U12636 (N_12636,N_12488,N_12513);
or U12637 (N_12637,N_12521,N_12527);
or U12638 (N_12638,N_12598,N_12546);
nand U12639 (N_12639,N_12559,N_12528);
nor U12640 (N_12640,N_12556,N_12483);
nor U12641 (N_12641,N_12480,N_12518);
nor U12642 (N_12642,N_12565,N_12450);
or U12643 (N_12643,N_12499,N_12582);
or U12644 (N_12644,N_12481,N_12453);
nand U12645 (N_12645,N_12583,N_12461);
and U12646 (N_12646,N_12457,N_12505);
or U12647 (N_12647,N_12534,N_12558);
nand U12648 (N_12648,N_12587,N_12452);
nand U12649 (N_12649,N_12468,N_12472);
and U12650 (N_12650,N_12503,N_12557);
nand U12651 (N_12651,N_12574,N_12522);
or U12652 (N_12652,N_12569,N_12494);
nor U12653 (N_12653,N_12485,N_12530);
or U12654 (N_12654,N_12596,N_12533);
or U12655 (N_12655,N_12592,N_12532);
xor U12656 (N_12656,N_12543,N_12599);
nor U12657 (N_12657,N_12478,N_12458);
and U12658 (N_12658,N_12576,N_12586);
nor U12659 (N_12659,N_12510,N_12538);
nand U12660 (N_12660,N_12566,N_12460);
or U12661 (N_12661,N_12572,N_12459);
or U12662 (N_12662,N_12506,N_12487);
or U12663 (N_12663,N_12451,N_12515);
and U12664 (N_12664,N_12524,N_12545);
and U12665 (N_12665,N_12477,N_12548);
and U12666 (N_12666,N_12497,N_12496);
or U12667 (N_12667,N_12498,N_12491);
nor U12668 (N_12668,N_12549,N_12526);
nand U12669 (N_12669,N_12525,N_12464);
or U12670 (N_12670,N_12471,N_12519);
nor U12671 (N_12671,N_12495,N_12492);
and U12672 (N_12672,N_12490,N_12562);
or U12673 (N_12673,N_12541,N_12550);
nor U12674 (N_12674,N_12455,N_12466);
and U12675 (N_12675,N_12596,N_12507);
or U12676 (N_12676,N_12540,N_12465);
nand U12677 (N_12677,N_12460,N_12495);
and U12678 (N_12678,N_12472,N_12594);
nand U12679 (N_12679,N_12580,N_12527);
or U12680 (N_12680,N_12539,N_12523);
nand U12681 (N_12681,N_12496,N_12571);
nand U12682 (N_12682,N_12546,N_12480);
xnor U12683 (N_12683,N_12511,N_12516);
nand U12684 (N_12684,N_12464,N_12451);
and U12685 (N_12685,N_12565,N_12585);
nor U12686 (N_12686,N_12564,N_12578);
and U12687 (N_12687,N_12530,N_12479);
and U12688 (N_12688,N_12491,N_12567);
nor U12689 (N_12689,N_12546,N_12552);
and U12690 (N_12690,N_12473,N_12573);
and U12691 (N_12691,N_12512,N_12561);
and U12692 (N_12692,N_12569,N_12464);
nand U12693 (N_12693,N_12538,N_12451);
nand U12694 (N_12694,N_12518,N_12527);
nor U12695 (N_12695,N_12456,N_12452);
nor U12696 (N_12696,N_12501,N_12461);
nand U12697 (N_12697,N_12595,N_12524);
or U12698 (N_12698,N_12485,N_12573);
or U12699 (N_12699,N_12505,N_12592);
nand U12700 (N_12700,N_12535,N_12488);
nand U12701 (N_12701,N_12543,N_12467);
or U12702 (N_12702,N_12461,N_12527);
or U12703 (N_12703,N_12475,N_12559);
xnor U12704 (N_12704,N_12562,N_12492);
nor U12705 (N_12705,N_12573,N_12502);
and U12706 (N_12706,N_12491,N_12559);
xnor U12707 (N_12707,N_12536,N_12478);
nand U12708 (N_12708,N_12484,N_12583);
nor U12709 (N_12709,N_12535,N_12536);
nor U12710 (N_12710,N_12564,N_12582);
nand U12711 (N_12711,N_12529,N_12497);
xnor U12712 (N_12712,N_12549,N_12592);
nor U12713 (N_12713,N_12480,N_12456);
nor U12714 (N_12714,N_12536,N_12534);
nor U12715 (N_12715,N_12548,N_12456);
or U12716 (N_12716,N_12530,N_12577);
nand U12717 (N_12717,N_12514,N_12511);
nor U12718 (N_12718,N_12566,N_12534);
xnor U12719 (N_12719,N_12565,N_12513);
and U12720 (N_12720,N_12511,N_12452);
nand U12721 (N_12721,N_12541,N_12529);
or U12722 (N_12722,N_12551,N_12569);
and U12723 (N_12723,N_12501,N_12454);
nor U12724 (N_12724,N_12506,N_12551);
and U12725 (N_12725,N_12457,N_12473);
and U12726 (N_12726,N_12575,N_12582);
and U12727 (N_12727,N_12495,N_12571);
nand U12728 (N_12728,N_12479,N_12543);
nor U12729 (N_12729,N_12496,N_12589);
or U12730 (N_12730,N_12456,N_12561);
or U12731 (N_12731,N_12471,N_12515);
nand U12732 (N_12732,N_12573,N_12595);
nor U12733 (N_12733,N_12499,N_12518);
or U12734 (N_12734,N_12462,N_12466);
nand U12735 (N_12735,N_12597,N_12561);
xor U12736 (N_12736,N_12558,N_12595);
nand U12737 (N_12737,N_12457,N_12584);
nor U12738 (N_12738,N_12527,N_12483);
and U12739 (N_12739,N_12554,N_12501);
nor U12740 (N_12740,N_12528,N_12564);
or U12741 (N_12741,N_12574,N_12491);
or U12742 (N_12742,N_12565,N_12596);
or U12743 (N_12743,N_12539,N_12518);
and U12744 (N_12744,N_12493,N_12587);
and U12745 (N_12745,N_12543,N_12544);
nor U12746 (N_12746,N_12533,N_12550);
and U12747 (N_12747,N_12453,N_12492);
nor U12748 (N_12748,N_12523,N_12554);
nor U12749 (N_12749,N_12588,N_12489);
and U12750 (N_12750,N_12747,N_12688);
and U12751 (N_12751,N_12644,N_12735);
and U12752 (N_12752,N_12720,N_12667);
nor U12753 (N_12753,N_12689,N_12725);
or U12754 (N_12754,N_12648,N_12623);
xor U12755 (N_12755,N_12712,N_12716);
xnor U12756 (N_12756,N_12603,N_12741);
xor U12757 (N_12757,N_12730,N_12654);
nand U12758 (N_12758,N_12671,N_12633);
or U12759 (N_12759,N_12727,N_12622);
nand U12760 (N_12760,N_12736,N_12637);
nor U12761 (N_12761,N_12641,N_12699);
nor U12762 (N_12762,N_12728,N_12615);
or U12763 (N_12763,N_12690,N_12605);
nor U12764 (N_12764,N_12620,N_12652);
xnor U12765 (N_12765,N_12729,N_12706);
or U12766 (N_12766,N_12744,N_12634);
or U12767 (N_12767,N_12681,N_12610);
nor U12768 (N_12768,N_12711,N_12626);
nand U12769 (N_12769,N_12650,N_12701);
nand U12770 (N_12770,N_12670,N_12635);
or U12771 (N_12771,N_12638,N_12657);
nor U12772 (N_12772,N_12694,N_12703);
or U12773 (N_12773,N_12674,N_12684);
nand U12774 (N_12774,N_12613,N_12697);
nor U12775 (N_12775,N_12672,N_12614);
or U12776 (N_12776,N_12616,N_12748);
or U12777 (N_12777,N_12708,N_12721);
nand U12778 (N_12778,N_12602,N_12642);
or U12779 (N_12779,N_12737,N_12609);
or U12780 (N_12780,N_12612,N_12619);
nand U12781 (N_12781,N_12719,N_12700);
xnor U12782 (N_12782,N_12643,N_12669);
nand U12783 (N_12783,N_12646,N_12679);
and U12784 (N_12784,N_12621,N_12702);
nor U12785 (N_12785,N_12718,N_12695);
nand U12786 (N_12786,N_12601,N_12691);
nor U12787 (N_12787,N_12743,N_12604);
nand U12788 (N_12788,N_12606,N_12661);
or U12789 (N_12789,N_12723,N_12731);
or U12790 (N_12790,N_12707,N_12739);
and U12791 (N_12791,N_12732,N_12649);
xnor U12792 (N_12792,N_12715,N_12660);
nand U12793 (N_12793,N_12713,N_12636);
nor U12794 (N_12794,N_12631,N_12710);
and U12795 (N_12795,N_12709,N_12717);
nor U12796 (N_12796,N_12668,N_12617);
and U12797 (N_12797,N_12632,N_12628);
or U12798 (N_12798,N_12675,N_12704);
nand U12799 (N_12799,N_12663,N_12733);
and U12800 (N_12800,N_12625,N_12607);
and U12801 (N_12801,N_12692,N_12693);
nor U12802 (N_12802,N_12659,N_12705);
nor U12803 (N_12803,N_12742,N_12611);
or U12804 (N_12804,N_12624,N_12738);
xor U12805 (N_12805,N_12724,N_12745);
nor U12806 (N_12806,N_12656,N_12645);
nand U12807 (N_12807,N_12714,N_12665);
or U12808 (N_12808,N_12629,N_12627);
or U12809 (N_12809,N_12618,N_12658);
nor U12810 (N_12810,N_12640,N_12746);
nand U12811 (N_12811,N_12662,N_12653);
or U12812 (N_12812,N_12651,N_12683);
and U12813 (N_12813,N_12676,N_12687);
nor U12814 (N_12814,N_12677,N_12734);
and U12815 (N_12815,N_12682,N_12655);
nand U12816 (N_12816,N_12673,N_12630);
nor U12817 (N_12817,N_12698,N_12664);
nor U12818 (N_12818,N_12680,N_12678);
xnor U12819 (N_12819,N_12726,N_12666);
or U12820 (N_12820,N_12722,N_12686);
or U12821 (N_12821,N_12647,N_12685);
and U12822 (N_12822,N_12749,N_12608);
or U12823 (N_12823,N_12696,N_12600);
nor U12824 (N_12824,N_12740,N_12639);
nand U12825 (N_12825,N_12692,N_12724);
nand U12826 (N_12826,N_12687,N_12609);
xor U12827 (N_12827,N_12729,N_12638);
nand U12828 (N_12828,N_12704,N_12737);
nand U12829 (N_12829,N_12698,N_12686);
nand U12830 (N_12830,N_12600,N_12708);
and U12831 (N_12831,N_12684,N_12697);
nor U12832 (N_12832,N_12604,N_12626);
xnor U12833 (N_12833,N_12738,N_12608);
nor U12834 (N_12834,N_12604,N_12671);
and U12835 (N_12835,N_12718,N_12666);
nand U12836 (N_12836,N_12626,N_12732);
nand U12837 (N_12837,N_12697,N_12628);
and U12838 (N_12838,N_12736,N_12633);
nor U12839 (N_12839,N_12671,N_12628);
or U12840 (N_12840,N_12681,N_12636);
nor U12841 (N_12841,N_12660,N_12601);
or U12842 (N_12842,N_12600,N_12711);
or U12843 (N_12843,N_12602,N_12669);
and U12844 (N_12844,N_12677,N_12671);
nor U12845 (N_12845,N_12702,N_12694);
nand U12846 (N_12846,N_12625,N_12626);
or U12847 (N_12847,N_12710,N_12650);
nand U12848 (N_12848,N_12633,N_12620);
nand U12849 (N_12849,N_12749,N_12701);
nand U12850 (N_12850,N_12685,N_12725);
and U12851 (N_12851,N_12703,N_12670);
nor U12852 (N_12852,N_12718,N_12603);
and U12853 (N_12853,N_12645,N_12693);
nor U12854 (N_12854,N_12613,N_12609);
xor U12855 (N_12855,N_12622,N_12606);
nand U12856 (N_12856,N_12685,N_12681);
nor U12857 (N_12857,N_12674,N_12646);
and U12858 (N_12858,N_12664,N_12691);
nand U12859 (N_12859,N_12713,N_12726);
nand U12860 (N_12860,N_12694,N_12679);
xnor U12861 (N_12861,N_12722,N_12680);
or U12862 (N_12862,N_12676,N_12725);
or U12863 (N_12863,N_12692,N_12613);
and U12864 (N_12864,N_12624,N_12605);
or U12865 (N_12865,N_12690,N_12643);
nor U12866 (N_12866,N_12697,N_12603);
xnor U12867 (N_12867,N_12627,N_12674);
and U12868 (N_12868,N_12716,N_12631);
and U12869 (N_12869,N_12694,N_12640);
xnor U12870 (N_12870,N_12636,N_12746);
nand U12871 (N_12871,N_12684,N_12660);
and U12872 (N_12872,N_12613,N_12735);
nor U12873 (N_12873,N_12607,N_12614);
and U12874 (N_12874,N_12746,N_12606);
nor U12875 (N_12875,N_12626,N_12601);
and U12876 (N_12876,N_12689,N_12614);
nand U12877 (N_12877,N_12707,N_12654);
xor U12878 (N_12878,N_12635,N_12668);
nor U12879 (N_12879,N_12640,N_12685);
nand U12880 (N_12880,N_12661,N_12699);
and U12881 (N_12881,N_12636,N_12626);
or U12882 (N_12882,N_12652,N_12640);
nor U12883 (N_12883,N_12656,N_12742);
and U12884 (N_12884,N_12708,N_12695);
and U12885 (N_12885,N_12608,N_12723);
nand U12886 (N_12886,N_12638,N_12669);
nand U12887 (N_12887,N_12726,N_12643);
and U12888 (N_12888,N_12693,N_12653);
nand U12889 (N_12889,N_12685,N_12691);
nor U12890 (N_12890,N_12730,N_12723);
nor U12891 (N_12891,N_12697,N_12630);
and U12892 (N_12892,N_12641,N_12688);
and U12893 (N_12893,N_12619,N_12701);
nand U12894 (N_12894,N_12720,N_12613);
and U12895 (N_12895,N_12603,N_12723);
or U12896 (N_12896,N_12670,N_12610);
or U12897 (N_12897,N_12617,N_12711);
nor U12898 (N_12898,N_12620,N_12712);
and U12899 (N_12899,N_12613,N_12628);
or U12900 (N_12900,N_12852,N_12872);
nor U12901 (N_12901,N_12858,N_12860);
and U12902 (N_12902,N_12897,N_12878);
nor U12903 (N_12903,N_12841,N_12887);
nand U12904 (N_12904,N_12877,N_12757);
and U12905 (N_12905,N_12770,N_12783);
or U12906 (N_12906,N_12828,N_12755);
nor U12907 (N_12907,N_12801,N_12827);
and U12908 (N_12908,N_12809,N_12888);
nand U12909 (N_12909,N_12787,N_12855);
nor U12910 (N_12910,N_12797,N_12843);
nand U12911 (N_12911,N_12867,N_12895);
nor U12912 (N_12912,N_12874,N_12778);
nor U12913 (N_12913,N_12847,N_12898);
and U12914 (N_12914,N_12825,N_12870);
nor U12915 (N_12915,N_12826,N_12844);
and U12916 (N_12916,N_12873,N_12869);
or U12917 (N_12917,N_12823,N_12790);
nor U12918 (N_12918,N_12818,N_12892);
or U12919 (N_12919,N_12875,N_12880);
nand U12920 (N_12920,N_12794,N_12891);
nand U12921 (N_12921,N_12798,N_12863);
or U12922 (N_12922,N_12767,N_12805);
nand U12923 (N_12923,N_12859,N_12806);
nand U12924 (N_12924,N_12807,N_12829);
and U12925 (N_12925,N_12853,N_12845);
and U12926 (N_12926,N_12754,N_12899);
xor U12927 (N_12927,N_12791,N_12766);
or U12928 (N_12928,N_12882,N_12784);
and U12929 (N_12929,N_12884,N_12820);
xor U12930 (N_12930,N_12832,N_12883);
nand U12931 (N_12931,N_12851,N_12840);
nand U12932 (N_12932,N_12751,N_12865);
xnor U12933 (N_12933,N_12868,N_12881);
nand U12934 (N_12934,N_12804,N_12765);
nor U12935 (N_12935,N_12803,N_12792);
xnor U12936 (N_12936,N_12812,N_12822);
nand U12937 (N_12937,N_12854,N_12759);
nor U12938 (N_12938,N_12779,N_12810);
nor U12939 (N_12939,N_12835,N_12893);
nand U12940 (N_12940,N_12890,N_12876);
and U12941 (N_12941,N_12814,N_12824);
nor U12942 (N_12942,N_12813,N_12815);
and U12943 (N_12943,N_12793,N_12802);
nand U12944 (N_12944,N_12830,N_12795);
nand U12945 (N_12945,N_12842,N_12856);
xor U12946 (N_12946,N_12771,N_12821);
nand U12947 (N_12947,N_12864,N_12889);
nand U12948 (N_12948,N_12789,N_12816);
or U12949 (N_12949,N_12837,N_12773);
and U12950 (N_12950,N_12811,N_12800);
or U12951 (N_12951,N_12808,N_12871);
and U12952 (N_12952,N_12846,N_12750);
and U12953 (N_12953,N_12760,N_12799);
nand U12954 (N_12954,N_12761,N_12831);
and U12955 (N_12955,N_12753,N_12777);
or U12956 (N_12956,N_12862,N_12817);
xnor U12957 (N_12957,N_12879,N_12763);
nor U12958 (N_12958,N_12886,N_12833);
nand U12959 (N_12959,N_12752,N_12861);
or U12960 (N_12960,N_12781,N_12850);
or U12961 (N_12961,N_12849,N_12896);
and U12962 (N_12962,N_12756,N_12836);
and U12963 (N_12963,N_12782,N_12819);
and U12964 (N_12964,N_12762,N_12776);
nor U12965 (N_12965,N_12780,N_12796);
nand U12966 (N_12966,N_12769,N_12834);
and U12967 (N_12967,N_12839,N_12885);
or U12968 (N_12968,N_12785,N_12775);
and U12969 (N_12969,N_12772,N_12866);
or U12970 (N_12970,N_12838,N_12764);
and U12971 (N_12971,N_12758,N_12786);
nor U12972 (N_12972,N_12848,N_12774);
and U12973 (N_12973,N_12857,N_12894);
or U12974 (N_12974,N_12788,N_12768);
nor U12975 (N_12975,N_12848,N_12881);
or U12976 (N_12976,N_12781,N_12796);
nor U12977 (N_12977,N_12778,N_12872);
xnor U12978 (N_12978,N_12778,N_12826);
nor U12979 (N_12979,N_12764,N_12858);
nand U12980 (N_12980,N_12832,N_12826);
and U12981 (N_12981,N_12799,N_12883);
and U12982 (N_12982,N_12788,N_12885);
nor U12983 (N_12983,N_12791,N_12823);
nand U12984 (N_12984,N_12760,N_12871);
and U12985 (N_12985,N_12870,N_12828);
and U12986 (N_12986,N_12803,N_12770);
nand U12987 (N_12987,N_12836,N_12863);
nor U12988 (N_12988,N_12799,N_12814);
nor U12989 (N_12989,N_12870,N_12763);
and U12990 (N_12990,N_12799,N_12865);
and U12991 (N_12991,N_12898,N_12884);
nand U12992 (N_12992,N_12801,N_12803);
or U12993 (N_12993,N_12844,N_12786);
or U12994 (N_12994,N_12899,N_12826);
nor U12995 (N_12995,N_12761,N_12848);
or U12996 (N_12996,N_12868,N_12753);
nand U12997 (N_12997,N_12837,N_12755);
and U12998 (N_12998,N_12837,N_12809);
nor U12999 (N_12999,N_12887,N_12867);
and U13000 (N_13000,N_12806,N_12787);
nand U13001 (N_13001,N_12850,N_12807);
nand U13002 (N_13002,N_12854,N_12864);
xnor U13003 (N_13003,N_12866,N_12814);
or U13004 (N_13004,N_12826,N_12891);
or U13005 (N_13005,N_12801,N_12879);
nor U13006 (N_13006,N_12899,N_12820);
or U13007 (N_13007,N_12849,N_12869);
or U13008 (N_13008,N_12776,N_12789);
and U13009 (N_13009,N_12756,N_12897);
xnor U13010 (N_13010,N_12892,N_12774);
xor U13011 (N_13011,N_12794,N_12882);
or U13012 (N_13012,N_12813,N_12847);
xor U13013 (N_13013,N_12867,N_12846);
xnor U13014 (N_13014,N_12893,N_12795);
or U13015 (N_13015,N_12851,N_12815);
and U13016 (N_13016,N_12814,N_12879);
nand U13017 (N_13017,N_12754,N_12803);
or U13018 (N_13018,N_12800,N_12873);
and U13019 (N_13019,N_12868,N_12892);
xnor U13020 (N_13020,N_12810,N_12879);
nand U13021 (N_13021,N_12806,N_12825);
and U13022 (N_13022,N_12897,N_12849);
nor U13023 (N_13023,N_12818,N_12868);
nand U13024 (N_13024,N_12808,N_12753);
and U13025 (N_13025,N_12810,N_12892);
nand U13026 (N_13026,N_12791,N_12878);
nand U13027 (N_13027,N_12864,N_12832);
nor U13028 (N_13028,N_12783,N_12752);
and U13029 (N_13029,N_12750,N_12865);
or U13030 (N_13030,N_12782,N_12800);
or U13031 (N_13031,N_12893,N_12782);
and U13032 (N_13032,N_12783,N_12862);
nor U13033 (N_13033,N_12786,N_12755);
nor U13034 (N_13034,N_12809,N_12751);
nand U13035 (N_13035,N_12828,N_12832);
nor U13036 (N_13036,N_12819,N_12781);
and U13037 (N_13037,N_12870,N_12779);
and U13038 (N_13038,N_12781,N_12831);
and U13039 (N_13039,N_12775,N_12784);
nand U13040 (N_13040,N_12823,N_12858);
or U13041 (N_13041,N_12811,N_12847);
nor U13042 (N_13042,N_12764,N_12895);
nand U13043 (N_13043,N_12769,N_12850);
nand U13044 (N_13044,N_12866,N_12840);
nor U13045 (N_13045,N_12798,N_12894);
nand U13046 (N_13046,N_12854,N_12890);
nor U13047 (N_13047,N_12879,N_12796);
or U13048 (N_13048,N_12859,N_12876);
or U13049 (N_13049,N_12857,N_12860);
nand U13050 (N_13050,N_12908,N_13026);
nor U13051 (N_13051,N_12985,N_13020);
and U13052 (N_13052,N_13048,N_13033);
nand U13053 (N_13053,N_12914,N_13029);
xnor U13054 (N_13054,N_12978,N_13010);
or U13055 (N_13055,N_12915,N_12929);
nor U13056 (N_13056,N_12995,N_13047);
and U13057 (N_13057,N_12917,N_12948);
xor U13058 (N_13058,N_12916,N_12909);
nand U13059 (N_13059,N_12990,N_12949);
nor U13060 (N_13060,N_12927,N_13014);
nand U13061 (N_13061,N_13038,N_12960);
and U13062 (N_13062,N_12986,N_12998);
xor U13063 (N_13063,N_13021,N_12934);
nor U13064 (N_13064,N_13018,N_12944);
nor U13065 (N_13065,N_13005,N_13031);
nand U13066 (N_13066,N_13017,N_12906);
xnor U13067 (N_13067,N_12994,N_12970);
or U13068 (N_13068,N_12968,N_13028);
and U13069 (N_13069,N_13036,N_13012);
xnor U13070 (N_13070,N_12937,N_12969);
nor U13071 (N_13071,N_12953,N_12936);
nand U13072 (N_13072,N_13039,N_13003);
nand U13073 (N_13073,N_12935,N_12910);
and U13074 (N_13074,N_13007,N_12976);
nor U13075 (N_13075,N_12942,N_12923);
nand U13076 (N_13076,N_13037,N_12973);
nand U13077 (N_13077,N_12901,N_13049);
nand U13078 (N_13078,N_13001,N_12967);
or U13079 (N_13079,N_12919,N_13024);
nand U13080 (N_13080,N_12931,N_12912);
nand U13081 (N_13081,N_12954,N_12974);
or U13082 (N_13082,N_13015,N_12925);
nand U13083 (N_13083,N_12932,N_13004);
nand U13084 (N_13084,N_12913,N_12947);
nor U13085 (N_13085,N_13011,N_12930);
nor U13086 (N_13086,N_12982,N_13006);
nand U13087 (N_13087,N_12965,N_12922);
and U13088 (N_13088,N_12996,N_12950);
xnor U13089 (N_13089,N_12933,N_13045);
nor U13090 (N_13090,N_12962,N_12971);
and U13091 (N_13091,N_12964,N_12905);
nor U13092 (N_13092,N_12946,N_12939);
nand U13093 (N_13093,N_12924,N_12981);
nor U13094 (N_13094,N_12918,N_13000);
or U13095 (N_13095,N_13019,N_12988);
and U13096 (N_13096,N_12993,N_13044);
nand U13097 (N_13097,N_13030,N_12980);
nand U13098 (N_13098,N_12997,N_13013);
nand U13099 (N_13099,N_12921,N_12940);
or U13100 (N_13100,N_12999,N_12963);
and U13101 (N_13101,N_12987,N_12957);
nand U13102 (N_13102,N_12938,N_12975);
nor U13103 (N_13103,N_13002,N_13040);
xnor U13104 (N_13104,N_12951,N_12958);
or U13105 (N_13105,N_12928,N_12903);
and U13106 (N_13106,N_13042,N_13023);
nand U13107 (N_13107,N_12977,N_13046);
nor U13108 (N_13108,N_13043,N_13032);
xor U13109 (N_13109,N_12941,N_12900);
or U13110 (N_13110,N_13035,N_12943);
nor U13111 (N_13111,N_13025,N_12945);
nor U13112 (N_13112,N_12952,N_12989);
or U13113 (N_13113,N_12983,N_13022);
or U13114 (N_13114,N_12992,N_12979);
or U13115 (N_13115,N_13034,N_13009);
and U13116 (N_13116,N_12984,N_12959);
nand U13117 (N_13117,N_12920,N_12911);
or U13118 (N_13118,N_12926,N_12956);
xnor U13119 (N_13119,N_13008,N_13027);
xor U13120 (N_13120,N_12991,N_12907);
and U13121 (N_13121,N_12902,N_12955);
or U13122 (N_13122,N_13016,N_12972);
or U13123 (N_13123,N_12961,N_12966);
and U13124 (N_13124,N_13041,N_12904);
and U13125 (N_13125,N_12947,N_12904);
nor U13126 (N_13126,N_13040,N_12961);
nor U13127 (N_13127,N_13006,N_12992);
and U13128 (N_13128,N_12909,N_12968);
nand U13129 (N_13129,N_13029,N_12969);
xor U13130 (N_13130,N_12998,N_13007);
nand U13131 (N_13131,N_12991,N_12927);
nor U13132 (N_13132,N_12990,N_12904);
nand U13133 (N_13133,N_12949,N_12977);
nand U13134 (N_13134,N_12947,N_13040);
xor U13135 (N_13135,N_13025,N_12922);
xor U13136 (N_13136,N_12969,N_12947);
xnor U13137 (N_13137,N_12978,N_12974);
and U13138 (N_13138,N_12974,N_12903);
and U13139 (N_13139,N_13033,N_12913);
or U13140 (N_13140,N_12948,N_12983);
and U13141 (N_13141,N_12985,N_12972);
nor U13142 (N_13142,N_13018,N_13043);
nand U13143 (N_13143,N_12909,N_13020);
and U13144 (N_13144,N_12966,N_12910);
or U13145 (N_13145,N_12955,N_13022);
xnor U13146 (N_13146,N_13011,N_13014);
and U13147 (N_13147,N_13022,N_13009);
or U13148 (N_13148,N_12922,N_12985);
nand U13149 (N_13149,N_13009,N_12940);
nand U13150 (N_13150,N_13043,N_13033);
or U13151 (N_13151,N_12903,N_13047);
and U13152 (N_13152,N_13048,N_12930);
nand U13153 (N_13153,N_13000,N_13035);
and U13154 (N_13154,N_13003,N_13036);
nand U13155 (N_13155,N_13003,N_13008);
xor U13156 (N_13156,N_12979,N_12976);
and U13157 (N_13157,N_12948,N_13048);
nor U13158 (N_13158,N_13043,N_12971);
and U13159 (N_13159,N_13043,N_12995);
xnor U13160 (N_13160,N_12973,N_12922);
and U13161 (N_13161,N_12996,N_13013);
nand U13162 (N_13162,N_12912,N_13006);
or U13163 (N_13163,N_12999,N_13024);
nand U13164 (N_13164,N_13020,N_12900);
or U13165 (N_13165,N_12975,N_13035);
xnor U13166 (N_13166,N_13016,N_12945);
nand U13167 (N_13167,N_12996,N_12943);
nand U13168 (N_13168,N_12991,N_12947);
nor U13169 (N_13169,N_13028,N_12921);
nand U13170 (N_13170,N_12945,N_13047);
or U13171 (N_13171,N_13049,N_12993);
xnor U13172 (N_13172,N_13010,N_12925);
nor U13173 (N_13173,N_12972,N_12970);
nor U13174 (N_13174,N_13040,N_12945);
or U13175 (N_13175,N_13011,N_12909);
and U13176 (N_13176,N_12999,N_13044);
nand U13177 (N_13177,N_13009,N_13023);
xor U13178 (N_13178,N_12962,N_12978);
nand U13179 (N_13179,N_13016,N_12996);
or U13180 (N_13180,N_12908,N_12978);
nor U13181 (N_13181,N_13010,N_13032);
nand U13182 (N_13182,N_12922,N_12913);
or U13183 (N_13183,N_12961,N_12975);
and U13184 (N_13184,N_13042,N_13049);
nor U13185 (N_13185,N_13017,N_13016);
nand U13186 (N_13186,N_12988,N_12918);
nand U13187 (N_13187,N_12923,N_12924);
nand U13188 (N_13188,N_12979,N_12940);
and U13189 (N_13189,N_12914,N_12962);
or U13190 (N_13190,N_13010,N_12956);
nand U13191 (N_13191,N_13013,N_12907);
and U13192 (N_13192,N_12908,N_13039);
nor U13193 (N_13193,N_12958,N_12950);
xnor U13194 (N_13194,N_12993,N_13010);
and U13195 (N_13195,N_12965,N_12946);
or U13196 (N_13196,N_12960,N_12901);
or U13197 (N_13197,N_12902,N_12920);
and U13198 (N_13198,N_12919,N_12940);
or U13199 (N_13199,N_12968,N_12954);
nand U13200 (N_13200,N_13085,N_13070);
nand U13201 (N_13201,N_13186,N_13082);
or U13202 (N_13202,N_13062,N_13162);
and U13203 (N_13203,N_13163,N_13118);
nor U13204 (N_13204,N_13127,N_13172);
or U13205 (N_13205,N_13181,N_13164);
nor U13206 (N_13206,N_13170,N_13199);
and U13207 (N_13207,N_13138,N_13130);
nor U13208 (N_13208,N_13132,N_13159);
and U13209 (N_13209,N_13120,N_13153);
and U13210 (N_13210,N_13165,N_13072);
and U13211 (N_13211,N_13089,N_13140);
and U13212 (N_13212,N_13080,N_13068);
nor U13213 (N_13213,N_13125,N_13103);
nand U13214 (N_13214,N_13106,N_13101);
nor U13215 (N_13215,N_13099,N_13161);
or U13216 (N_13216,N_13098,N_13086);
and U13217 (N_13217,N_13056,N_13176);
nand U13218 (N_13218,N_13150,N_13185);
and U13219 (N_13219,N_13087,N_13108);
or U13220 (N_13220,N_13105,N_13104);
nand U13221 (N_13221,N_13054,N_13193);
and U13222 (N_13222,N_13197,N_13050);
nand U13223 (N_13223,N_13183,N_13173);
and U13224 (N_13224,N_13175,N_13198);
and U13225 (N_13225,N_13188,N_13077);
or U13226 (N_13226,N_13128,N_13195);
nor U13227 (N_13227,N_13121,N_13133);
and U13228 (N_13228,N_13079,N_13191);
nand U13229 (N_13229,N_13129,N_13112);
nor U13230 (N_13230,N_13078,N_13053);
and U13231 (N_13231,N_13083,N_13126);
xnor U13232 (N_13232,N_13136,N_13100);
and U13233 (N_13233,N_13114,N_13180);
and U13234 (N_13234,N_13184,N_13156);
nor U13235 (N_13235,N_13073,N_13143);
or U13236 (N_13236,N_13051,N_13182);
xnor U13237 (N_13237,N_13142,N_13057);
nand U13238 (N_13238,N_13190,N_13096);
nand U13239 (N_13239,N_13144,N_13061);
and U13240 (N_13240,N_13154,N_13075);
xor U13241 (N_13241,N_13052,N_13091);
or U13242 (N_13242,N_13139,N_13064);
or U13243 (N_13243,N_13157,N_13145);
or U13244 (N_13244,N_13187,N_13189);
and U13245 (N_13245,N_13093,N_13076);
and U13246 (N_13246,N_13192,N_13092);
xnor U13247 (N_13247,N_13117,N_13081);
xor U13248 (N_13248,N_13137,N_13074);
nor U13249 (N_13249,N_13169,N_13178);
or U13250 (N_13250,N_13090,N_13088);
nand U13251 (N_13251,N_13059,N_13148);
or U13252 (N_13252,N_13151,N_13119);
nor U13253 (N_13253,N_13167,N_13131);
or U13254 (N_13254,N_13152,N_13113);
nor U13255 (N_13255,N_13060,N_13058);
or U13256 (N_13256,N_13147,N_13067);
and U13257 (N_13257,N_13122,N_13123);
or U13258 (N_13258,N_13102,N_13110);
or U13259 (N_13259,N_13069,N_13174);
and U13260 (N_13260,N_13071,N_13177);
or U13261 (N_13261,N_13109,N_13155);
or U13262 (N_13262,N_13097,N_13111);
xnor U13263 (N_13263,N_13134,N_13194);
nand U13264 (N_13264,N_13146,N_13107);
or U13265 (N_13265,N_13171,N_13066);
nor U13266 (N_13266,N_13095,N_13055);
nand U13267 (N_13267,N_13084,N_13166);
xor U13268 (N_13268,N_13115,N_13160);
nor U13269 (N_13269,N_13124,N_13196);
or U13270 (N_13270,N_13116,N_13135);
nand U13271 (N_13271,N_13065,N_13168);
nand U13272 (N_13272,N_13094,N_13158);
nor U13273 (N_13273,N_13063,N_13179);
nand U13274 (N_13274,N_13149,N_13141);
nand U13275 (N_13275,N_13138,N_13117);
or U13276 (N_13276,N_13131,N_13115);
or U13277 (N_13277,N_13096,N_13092);
or U13278 (N_13278,N_13082,N_13119);
xor U13279 (N_13279,N_13117,N_13112);
or U13280 (N_13280,N_13141,N_13076);
and U13281 (N_13281,N_13106,N_13118);
and U13282 (N_13282,N_13165,N_13175);
nor U13283 (N_13283,N_13183,N_13057);
nand U13284 (N_13284,N_13102,N_13082);
xor U13285 (N_13285,N_13172,N_13072);
or U13286 (N_13286,N_13158,N_13115);
and U13287 (N_13287,N_13157,N_13055);
nand U13288 (N_13288,N_13128,N_13089);
nor U13289 (N_13289,N_13050,N_13193);
nor U13290 (N_13290,N_13143,N_13192);
and U13291 (N_13291,N_13065,N_13115);
and U13292 (N_13292,N_13069,N_13074);
and U13293 (N_13293,N_13058,N_13153);
nor U13294 (N_13294,N_13151,N_13070);
nor U13295 (N_13295,N_13176,N_13134);
nor U13296 (N_13296,N_13062,N_13125);
nand U13297 (N_13297,N_13150,N_13071);
and U13298 (N_13298,N_13106,N_13144);
xor U13299 (N_13299,N_13056,N_13196);
nor U13300 (N_13300,N_13150,N_13135);
or U13301 (N_13301,N_13152,N_13158);
and U13302 (N_13302,N_13086,N_13129);
and U13303 (N_13303,N_13108,N_13127);
nand U13304 (N_13304,N_13077,N_13052);
nor U13305 (N_13305,N_13181,N_13152);
or U13306 (N_13306,N_13071,N_13060);
nand U13307 (N_13307,N_13150,N_13139);
and U13308 (N_13308,N_13150,N_13137);
and U13309 (N_13309,N_13184,N_13132);
nand U13310 (N_13310,N_13163,N_13170);
nand U13311 (N_13311,N_13084,N_13196);
nand U13312 (N_13312,N_13138,N_13114);
nand U13313 (N_13313,N_13096,N_13191);
nand U13314 (N_13314,N_13072,N_13146);
or U13315 (N_13315,N_13061,N_13198);
or U13316 (N_13316,N_13108,N_13100);
and U13317 (N_13317,N_13092,N_13050);
nand U13318 (N_13318,N_13059,N_13093);
and U13319 (N_13319,N_13096,N_13091);
and U13320 (N_13320,N_13115,N_13143);
and U13321 (N_13321,N_13177,N_13152);
nand U13322 (N_13322,N_13087,N_13179);
nor U13323 (N_13323,N_13065,N_13093);
nor U13324 (N_13324,N_13188,N_13112);
and U13325 (N_13325,N_13103,N_13153);
nand U13326 (N_13326,N_13159,N_13137);
and U13327 (N_13327,N_13154,N_13146);
and U13328 (N_13328,N_13084,N_13104);
nor U13329 (N_13329,N_13164,N_13107);
nand U13330 (N_13330,N_13090,N_13141);
and U13331 (N_13331,N_13152,N_13084);
or U13332 (N_13332,N_13107,N_13197);
or U13333 (N_13333,N_13110,N_13116);
nor U13334 (N_13334,N_13142,N_13099);
nor U13335 (N_13335,N_13118,N_13117);
and U13336 (N_13336,N_13162,N_13091);
nand U13337 (N_13337,N_13069,N_13194);
nand U13338 (N_13338,N_13131,N_13158);
or U13339 (N_13339,N_13055,N_13174);
or U13340 (N_13340,N_13133,N_13059);
nand U13341 (N_13341,N_13129,N_13172);
nor U13342 (N_13342,N_13172,N_13073);
nor U13343 (N_13343,N_13051,N_13132);
and U13344 (N_13344,N_13115,N_13050);
and U13345 (N_13345,N_13079,N_13193);
nand U13346 (N_13346,N_13082,N_13060);
xnor U13347 (N_13347,N_13133,N_13149);
nand U13348 (N_13348,N_13063,N_13187);
nand U13349 (N_13349,N_13086,N_13063);
nand U13350 (N_13350,N_13218,N_13296);
or U13351 (N_13351,N_13318,N_13252);
nor U13352 (N_13352,N_13311,N_13214);
nand U13353 (N_13353,N_13337,N_13270);
nor U13354 (N_13354,N_13259,N_13266);
nand U13355 (N_13355,N_13275,N_13328);
nor U13356 (N_13356,N_13297,N_13329);
xor U13357 (N_13357,N_13344,N_13294);
nor U13358 (N_13358,N_13308,N_13211);
nand U13359 (N_13359,N_13342,N_13242);
and U13360 (N_13360,N_13249,N_13298);
and U13361 (N_13361,N_13343,N_13234);
nand U13362 (N_13362,N_13248,N_13282);
xor U13363 (N_13363,N_13295,N_13307);
and U13364 (N_13364,N_13280,N_13274);
and U13365 (N_13365,N_13209,N_13217);
or U13366 (N_13366,N_13320,N_13278);
or U13367 (N_13367,N_13306,N_13335);
and U13368 (N_13368,N_13221,N_13247);
and U13369 (N_13369,N_13310,N_13265);
or U13370 (N_13370,N_13314,N_13333);
and U13371 (N_13371,N_13207,N_13228);
nor U13372 (N_13372,N_13345,N_13271);
nor U13373 (N_13373,N_13347,N_13288);
and U13374 (N_13374,N_13290,N_13230);
or U13375 (N_13375,N_13201,N_13348);
nand U13376 (N_13376,N_13276,N_13309);
or U13377 (N_13377,N_13303,N_13219);
or U13378 (N_13378,N_13220,N_13237);
and U13379 (N_13379,N_13240,N_13215);
and U13380 (N_13380,N_13272,N_13317);
xor U13381 (N_13381,N_13305,N_13299);
nor U13382 (N_13382,N_13269,N_13331);
xor U13383 (N_13383,N_13202,N_13263);
nor U13384 (N_13384,N_13206,N_13289);
nor U13385 (N_13385,N_13256,N_13205);
or U13386 (N_13386,N_13339,N_13319);
nand U13387 (N_13387,N_13284,N_13203);
nand U13388 (N_13388,N_13236,N_13225);
nor U13389 (N_13389,N_13224,N_13268);
nand U13390 (N_13390,N_13302,N_13233);
or U13391 (N_13391,N_13281,N_13255);
nand U13392 (N_13392,N_13216,N_13287);
nor U13393 (N_13393,N_13283,N_13291);
and U13394 (N_13394,N_13251,N_13332);
nor U13395 (N_13395,N_13300,N_13244);
nand U13396 (N_13396,N_13349,N_13315);
nand U13397 (N_13397,N_13235,N_13267);
and U13398 (N_13398,N_13254,N_13323);
nand U13399 (N_13399,N_13273,N_13212);
nor U13400 (N_13400,N_13312,N_13250);
or U13401 (N_13401,N_13338,N_13210);
nand U13402 (N_13402,N_13293,N_13346);
nand U13403 (N_13403,N_13301,N_13223);
or U13404 (N_13404,N_13279,N_13246);
nand U13405 (N_13405,N_13286,N_13226);
nor U13406 (N_13406,N_13261,N_13243);
and U13407 (N_13407,N_13325,N_13257);
and U13408 (N_13408,N_13262,N_13260);
nand U13409 (N_13409,N_13330,N_13322);
xnor U13410 (N_13410,N_13258,N_13341);
nand U13411 (N_13411,N_13208,N_13292);
xnor U13412 (N_13412,N_13204,N_13231);
nand U13413 (N_13413,N_13253,N_13327);
nand U13414 (N_13414,N_13340,N_13285);
nor U13415 (N_13415,N_13245,N_13304);
nor U13416 (N_13416,N_13213,N_13232);
and U13417 (N_13417,N_13264,N_13326);
nand U13418 (N_13418,N_13227,N_13222);
nor U13419 (N_13419,N_13239,N_13316);
nor U13420 (N_13420,N_13324,N_13313);
or U13421 (N_13421,N_13241,N_13321);
or U13422 (N_13422,N_13277,N_13229);
and U13423 (N_13423,N_13334,N_13200);
nand U13424 (N_13424,N_13238,N_13336);
nor U13425 (N_13425,N_13226,N_13258);
and U13426 (N_13426,N_13299,N_13240);
and U13427 (N_13427,N_13210,N_13308);
or U13428 (N_13428,N_13233,N_13346);
nand U13429 (N_13429,N_13240,N_13234);
nand U13430 (N_13430,N_13236,N_13213);
nor U13431 (N_13431,N_13215,N_13245);
or U13432 (N_13432,N_13311,N_13289);
nor U13433 (N_13433,N_13285,N_13335);
nor U13434 (N_13434,N_13204,N_13283);
nor U13435 (N_13435,N_13343,N_13299);
or U13436 (N_13436,N_13333,N_13229);
nand U13437 (N_13437,N_13223,N_13271);
nor U13438 (N_13438,N_13327,N_13237);
nand U13439 (N_13439,N_13270,N_13348);
and U13440 (N_13440,N_13336,N_13214);
or U13441 (N_13441,N_13267,N_13261);
nand U13442 (N_13442,N_13209,N_13202);
and U13443 (N_13443,N_13291,N_13280);
nor U13444 (N_13444,N_13307,N_13277);
or U13445 (N_13445,N_13204,N_13280);
nand U13446 (N_13446,N_13310,N_13231);
nand U13447 (N_13447,N_13230,N_13298);
nor U13448 (N_13448,N_13306,N_13329);
nor U13449 (N_13449,N_13234,N_13292);
nor U13450 (N_13450,N_13331,N_13292);
and U13451 (N_13451,N_13265,N_13281);
and U13452 (N_13452,N_13261,N_13215);
nand U13453 (N_13453,N_13279,N_13267);
xor U13454 (N_13454,N_13260,N_13247);
nand U13455 (N_13455,N_13339,N_13213);
and U13456 (N_13456,N_13320,N_13249);
nand U13457 (N_13457,N_13290,N_13208);
nand U13458 (N_13458,N_13268,N_13270);
nor U13459 (N_13459,N_13249,N_13210);
and U13460 (N_13460,N_13257,N_13273);
nor U13461 (N_13461,N_13291,N_13286);
nor U13462 (N_13462,N_13259,N_13268);
or U13463 (N_13463,N_13267,N_13237);
or U13464 (N_13464,N_13225,N_13306);
or U13465 (N_13465,N_13305,N_13204);
or U13466 (N_13466,N_13317,N_13263);
and U13467 (N_13467,N_13283,N_13206);
and U13468 (N_13468,N_13225,N_13289);
or U13469 (N_13469,N_13278,N_13231);
or U13470 (N_13470,N_13228,N_13261);
nand U13471 (N_13471,N_13323,N_13279);
nand U13472 (N_13472,N_13213,N_13334);
and U13473 (N_13473,N_13261,N_13303);
nand U13474 (N_13474,N_13283,N_13231);
and U13475 (N_13475,N_13347,N_13316);
or U13476 (N_13476,N_13254,N_13212);
nand U13477 (N_13477,N_13240,N_13322);
and U13478 (N_13478,N_13325,N_13295);
xnor U13479 (N_13479,N_13211,N_13291);
or U13480 (N_13480,N_13297,N_13226);
nor U13481 (N_13481,N_13312,N_13295);
nand U13482 (N_13482,N_13238,N_13202);
or U13483 (N_13483,N_13341,N_13347);
or U13484 (N_13484,N_13298,N_13315);
xor U13485 (N_13485,N_13229,N_13251);
and U13486 (N_13486,N_13329,N_13282);
and U13487 (N_13487,N_13251,N_13240);
or U13488 (N_13488,N_13323,N_13225);
and U13489 (N_13489,N_13239,N_13262);
xor U13490 (N_13490,N_13331,N_13333);
and U13491 (N_13491,N_13313,N_13346);
and U13492 (N_13492,N_13226,N_13288);
nor U13493 (N_13493,N_13321,N_13232);
or U13494 (N_13494,N_13223,N_13250);
xor U13495 (N_13495,N_13239,N_13319);
or U13496 (N_13496,N_13301,N_13345);
nand U13497 (N_13497,N_13212,N_13255);
nand U13498 (N_13498,N_13327,N_13225);
nor U13499 (N_13499,N_13220,N_13332);
or U13500 (N_13500,N_13386,N_13480);
xor U13501 (N_13501,N_13395,N_13441);
and U13502 (N_13502,N_13471,N_13406);
and U13503 (N_13503,N_13353,N_13485);
or U13504 (N_13504,N_13352,N_13379);
nor U13505 (N_13505,N_13392,N_13458);
and U13506 (N_13506,N_13482,N_13421);
or U13507 (N_13507,N_13368,N_13469);
nand U13508 (N_13508,N_13449,N_13437);
and U13509 (N_13509,N_13397,N_13398);
xnor U13510 (N_13510,N_13410,N_13427);
and U13511 (N_13511,N_13390,N_13381);
nand U13512 (N_13512,N_13380,N_13457);
and U13513 (N_13513,N_13370,N_13434);
and U13514 (N_13514,N_13383,N_13402);
nor U13515 (N_13515,N_13375,N_13371);
or U13516 (N_13516,N_13497,N_13451);
nor U13517 (N_13517,N_13444,N_13414);
xnor U13518 (N_13518,N_13445,N_13465);
nor U13519 (N_13519,N_13473,N_13376);
nand U13520 (N_13520,N_13424,N_13422);
or U13521 (N_13521,N_13431,N_13420);
xnor U13522 (N_13522,N_13474,N_13439);
nor U13523 (N_13523,N_13433,N_13401);
nor U13524 (N_13524,N_13430,N_13400);
and U13525 (N_13525,N_13394,N_13389);
xnor U13526 (N_13526,N_13483,N_13452);
or U13527 (N_13527,N_13355,N_13432);
or U13528 (N_13528,N_13388,N_13374);
or U13529 (N_13529,N_13476,N_13396);
or U13530 (N_13530,N_13470,N_13372);
and U13531 (N_13531,N_13387,N_13498);
or U13532 (N_13532,N_13450,N_13484);
and U13533 (N_13533,N_13418,N_13463);
nor U13534 (N_13534,N_13479,N_13385);
nand U13535 (N_13535,N_13373,N_13436);
xnor U13536 (N_13536,N_13453,N_13423);
or U13537 (N_13537,N_13351,N_13364);
nand U13538 (N_13538,N_13363,N_13384);
and U13539 (N_13539,N_13362,N_13489);
and U13540 (N_13540,N_13358,N_13350);
nor U13541 (N_13541,N_13412,N_13496);
and U13542 (N_13542,N_13366,N_13499);
xnor U13543 (N_13543,N_13417,N_13391);
nand U13544 (N_13544,N_13454,N_13487);
and U13545 (N_13545,N_13378,N_13475);
and U13546 (N_13546,N_13357,N_13440);
or U13547 (N_13547,N_13495,N_13354);
nand U13548 (N_13548,N_13442,N_13472);
xnor U13549 (N_13549,N_13478,N_13425);
nand U13550 (N_13550,N_13435,N_13466);
nor U13551 (N_13551,N_13367,N_13443);
or U13552 (N_13552,N_13456,N_13369);
nand U13553 (N_13553,N_13356,N_13464);
and U13554 (N_13554,N_13403,N_13447);
or U13555 (N_13555,N_13404,N_13393);
and U13556 (N_13556,N_13407,N_13494);
xor U13557 (N_13557,N_13409,N_13377);
nand U13558 (N_13558,N_13408,N_13491);
and U13559 (N_13559,N_13359,N_13492);
or U13560 (N_13560,N_13477,N_13461);
nor U13561 (N_13561,N_13493,N_13488);
and U13562 (N_13562,N_13365,N_13360);
nor U13563 (N_13563,N_13467,N_13428);
nand U13564 (N_13564,N_13468,N_13462);
or U13565 (N_13565,N_13455,N_13399);
nand U13566 (N_13566,N_13448,N_13361);
or U13567 (N_13567,N_13446,N_13413);
and U13568 (N_13568,N_13416,N_13411);
or U13569 (N_13569,N_13405,N_13429);
nand U13570 (N_13570,N_13481,N_13426);
or U13571 (N_13571,N_13438,N_13460);
nand U13572 (N_13572,N_13419,N_13415);
or U13573 (N_13573,N_13382,N_13490);
nand U13574 (N_13574,N_13459,N_13486);
nand U13575 (N_13575,N_13390,N_13460);
nand U13576 (N_13576,N_13393,N_13454);
or U13577 (N_13577,N_13396,N_13446);
and U13578 (N_13578,N_13454,N_13391);
or U13579 (N_13579,N_13448,N_13375);
and U13580 (N_13580,N_13380,N_13448);
nor U13581 (N_13581,N_13442,N_13410);
or U13582 (N_13582,N_13385,N_13362);
xor U13583 (N_13583,N_13380,N_13441);
xor U13584 (N_13584,N_13424,N_13409);
and U13585 (N_13585,N_13379,N_13355);
and U13586 (N_13586,N_13496,N_13422);
or U13587 (N_13587,N_13465,N_13460);
nor U13588 (N_13588,N_13354,N_13397);
nand U13589 (N_13589,N_13459,N_13440);
and U13590 (N_13590,N_13428,N_13423);
nand U13591 (N_13591,N_13358,N_13471);
nor U13592 (N_13592,N_13356,N_13364);
nand U13593 (N_13593,N_13430,N_13483);
and U13594 (N_13594,N_13489,N_13407);
and U13595 (N_13595,N_13409,N_13456);
nand U13596 (N_13596,N_13444,N_13438);
nand U13597 (N_13597,N_13404,N_13462);
and U13598 (N_13598,N_13423,N_13410);
xnor U13599 (N_13599,N_13457,N_13379);
nand U13600 (N_13600,N_13428,N_13395);
and U13601 (N_13601,N_13426,N_13495);
and U13602 (N_13602,N_13365,N_13372);
xor U13603 (N_13603,N_13365,N_13481);
nand U13604 (N_13604,N_13385,N_13465);
and U13605 (N_13605,N_13456,N_13355);
nor U13606 (N_13606,N_13409,N_13497);
and U13607 (N_13607,N_13470,N_13407);
or U13608 (N_13608,N_13372,N_13461);
xnor U13609 (N_13609,N_13430,N_13485);
nand U13610 (N_13610,N_13443,N_13499);
nor U13611 (N_13611,N_13353,N_13416);
nor U13612 (N_13612,N_13406,N_13381);
or U13613 (N_13613,N_13428,N_13411);
nand U13614 (N_13614,N_13398,N_13370);
nor U13615 (N_13615,N_13376,N_13402);
nor U13616 (N_13616,N_13491,N_13477);
and U13617 (N_13617,N_13378,N_13412);
nand U13618 (N_13618,N_13491,N_13470);
nor U13619 (N_13619,N_13457,N_13368);
nor U13620 (N_13620,N_13499,N_13444);
nor U13621 (N_13621,N_13401,N_13475);
and U13622 (N_13622,N_13499,N_13422);
nand U13623 (N_13623,N_13399,N_13430);
and U13624 (N_13624,N_13462,N_13489);
nand U13625 (N_13625,N_13478,N_13398);
nor U13626 (N_13626,N_13450,N_13351);
nand U13627 (N_13627,N_13467,N_13486);
and U13628 (N_13628,N_13471,N_13498);
and U13629 (N_13629,N_13361,N_13419);
nand U13630 (N_13630,N_13477,N_13394);
and U13631 (N_13631,N_13407,N_13413);
xnor U13632 (N_13632,N_13353,N_13356);
nor U13633 (N_13633,N_13390,N_13425);
nor U13634 (N_13634,N_13428,N_13451);
xor U13635 (N_13635,N_13437,N_13469);
nor U13636 (N_13636,N_13361,N_13477);
or U13637 (N_13637,N_13421,N_13409);
and U13638 (N_13638,N_13474,N_13485);
nand U13639 (N_13639,N_13437,N_13459);
xnor U13640 (N_13640,N_13448,N_13381);
or U13641 (N_13641,N_13385,N_13493);
or U13642 (N_13642,N_13496,N_13481);
and U13643 (N_13643,N_13413,N_13396);
and U13644 (N_13644,N_13371,N_13469);
nor U13645 (N_13645,N_13369,N_13429);
nor U13646 (N_13646,N_13499,N_13417);
nor U13647 (N_13647,N_13410,N_13450);
or U13648 (N_13648,N_13463,N_13407);
or U13649 (N_13649,N_13362,N_13484);
and U13650 (N_13650,N_13525,N_13508);
and U13651 (N_13651,N_13535,N_13582);
nand U13652 (N_13652,N_13576,N_13533);
nor U13653 (N_13653,N_13560,N_13596);
nand U13654 (N_13654,N_13631,N_13648);
nand U13655 (N_13655,N_13540,N_13557);
and U13656 (N_13656,N_13520,N_13617);
nand U13657 (N_13657,N_13556,N_13623);
nand U13658 (N_13658,N_13615,N_13643);
or U13659 (N_13659,N_13517,N_13539);
nand U13660 (N_13660,N_13641,N_13592);
nand U13661 (N_13661,N_13604,N_13545);
and U13662 (N_13662,N_13642,N_13633);
nor U13663 (N_13663,N_13521,N_13632);
and U13664 (N_13664,N_13571,N_13563);
nand U13665 (N_13665,N_13630,N_13566);
nand U13666 (N_13666,N_13606,N_13528);
xnor U13667 (N_13667,N_13628,N_13640);
or U13668 (N_13668,N_13608,N_13534);
and U13669 (N_13669,N_13583,N_13523);
or U13670 (N_13670,N_13589,N_13618);
nand U13671 (N_13671,N_13512,N_13531);
or U13672 (N_13672,N_13624,N_13616);
nor U13673 (N_13673,N_13518,N_13603);
and U13674 (N_13674,N_13522,N_13547);
nor U13675 (N_13675,N_13567,N_13532);
or U13676 (N_13676,N_13519,N_13502);
nor U13677 (N_13677,N_13639,N_13568);
nand U13678 (N_13678,N_13538,N_13587);
xnor U13679 (N_13679,N_13501,N_13597);
nor U13680 (N_13680,N_13645,N_13551);
nand U13681 (N_13681,N_13605,N_13621);
and U13682 (N_13682,N_13637,N_13586);
nor U13683 (N_13683,N_13644,N_13613);
and U13684 (N_13684,N_13509,N_13504);
nand U13685 (N_13685,N_13553,N_13541);
nand U13686 (N_13686,N_13585,N_13578);
or U13687 (N_13687,N_13552,N_13544);
nor U13688 (N_13688,N_13626,N_13530);
nand U13689 (N_13689,N_13505,N_13607);
nand U13690 (N_13690,N_13565,N_13572);
nand U13691 (N_13691,N_13584,N_13562);
or U13692 (N_13692,N_13590,N_13647);
and U13693 (N_13693,N_13515,N_13574);
nor U13694 (N_13694,N_13638,N_13500);
and U13695 (N_13695,N_13620,N_13646);
or U13696 (N_13696,N_13510,N_13542);
and U13697 (N_13697,N_13595,N_13614);
xnor U13698 (N_13698,N_13543,N_13507);
and U13699 (N_13699,N_13526,N_13610);
nand U13700 (N_13700,N_13629,N_13527);
nand U13701 (N_13701,N_13602,N_13588);
nand U13702 (N_13702,N_13564,N_13577);
nor U13703 (N_13703,N_13549,N_13514);
and U13704 (N_13704,N_13649,N_13622);
nand U13705 (N_13705,N_13612,N_13516);
or U13706 (N_13706,N_13579,N_13581);
nand U13707 (N_13707,N_13573,N_13511);
nand U13708 (N_13708,N_13570,N_13524);
or U13709 (N_13709,N_13599,N_13634);
or U13710 (N_13710,N_13548,N_13636);
nand U13711 (N_13711,N_13627,N_13506);
xor U13712 (N_13712,N_13611,N_13550);
xnor U13713 (N_13713,N_13554,N_13575);
nand U13714 (N_13714,N_13619,N_13591);
or U13715 (N_13715,N_13601,N_13546);
and U13716 (N_13716,N_13529,N_13598);
and U13717 (N_13717,N_13537,N_13513);
or U13718 (N_13718,N_13635,N_13580);
nor U13719 (N_13719,N_13569,N_13561);
or U13720 (N_13720,N_13609,N_13559);
xnor U13721 (N_13721,N_13558,N_13593);
nor U13722 (N_13722,N_13503,N_13536);
nand U13723 (N_13723,N_13594,N_13625);
nand U13724 (N_13724,N_13555,N_13600);
or U13725 (N_13725,N_13500,N_13627);
nor U13726 (N_13726,N_13626,N_13644);
nor U13727 (N_13727,N_13585,N_13515);
nand U13728 (N_13728,N_13628,N_13546);
nor U13729 (N_13729,N_13616,N_13509);
and U13730 (N_13730,N_13638,N_13572);
nor U13731 (N_13731,N_13524,N_13509);
and U13732 (N_13732,N_13522,N_13553);
nand U13733 (N_13733,N_13562,N_13612);
nand U13734 (N_13734,N_13569,N_13536);
and U13735 (N_13735,N_13600,N_13612);
or U13736 (N_13736,N_13548,N_13531);
xnor U13737 (N_13737,N_13525,N_13569);
nor U13738 (N_13738,N_13501,N_13586);
or U13739 (N_13739,N_13635,N_13630);
or U13740 (N_13740,N_13574,N_13524);
and U13741 (N_13741,N_13638,N_13564);
and U13742 (N_13742,N_13526,N_13585);
nand U13743 (N_13743,N_13619,N_13516);
nor U13744 (N_13744,N_13640,N_13554);
nand U13745 (N_13745,N_13577,N_13503);
or U13746 (N_13746,N_13524,N_13567);
nor U13747 (N_13747,N_13605,N_13532);
or U13748 (N_13748,N_13564,N_13562);
or U13749 (N_13749,N_13520,N_13589);
nor U13750 (N_13750,N_13579,N_13586);
nor U13751 (N_13751,N_13608,N_13645);
and U13752 (N_13752,N_13518,N_13581);
nand U13753 (N_13753,N_13604,N_13591);
nor U13754 (N_13754,N_13646,N_13525);
and U13755 (N_13755,N_13620,N_13606);
or U13756 (N_13756,N_13610,N_13623);
or U13757 (N_13757,N_13514,N_13609);
or U13758 (N_13758,N_13511,N_13614);
nand U13759 (N_13759,N_13632,N_13589);
xnor U13760 (N_13760,N_13552,N_13617);
nand U13761 (N_13761,N_13566,N_13509);
nand U13762 (N_13762,N_13567,N_13517);
or U13763 (N_13763,N_13524,N_13604);
nand U13764 (N_13764,N_13648,N_13503);
and U13765 (N_13765,N_13534,N_13579);
or U13766 (N_13766,N_13633,N_13520);
nor U13767 (N_13767,N_13586,N_13578);
and U13768 (N_13768,N_13588,N_13540);
and U13769 (N_13769,N_13576,N_13537);
nand U13770 (N_13770,N_13553,N_13626);
nor U13771 (N_13771,N_13567,N_13564);
nor U13772 (N_13772,N_13550,N_13532);
nand U13773 (N_13773,N_13573,N_13646);
or U13774 (N_13774,N_13590,N_13593);
or U13775 (N_13775,N_13617,N_13641);
nand U13776 (N_13776,N_13501,N_13609);
or U13777 (N_13777,N_13566,N_13532);
nor U13778 (N_13778,N_13522,N_13622);
or U13779 (N_13779,N_13639,N_13574);
and U13780 (N_13780,N_13537,N_13567);
nor U13781 (N_13781,N_13606,N_13502);
nand U13782 (N_13782,N_13601,N_13505);
nor U13783 (N_13783,N_13593,N_13641);
xor U13784 (N_13784,N_13538,N_13575);
nand U13785 (N_13785,N_13607,N_13640);
nand U13786 (N_13786,N_13621,N_13566);
and U13787 (N_13787,N_13539,N_13617);
and U13788 (N_13788,N_13609,N_13581);
nand U13789 (N_13789,N_13528,N_13504);
nand U13790 (N_13790,N_13611,N_13601);
or U13791 (N_13791,N_13609,N_13611);
and U13792 (N_13792,N_13595,N_13624);
and U13793 (N_13793,N_13640,N_13519);
nor U13794 (N_13794,N_13618,N_13518);
nand U13795 (N_13795,N_13506,N_13572);
nor U13796 (N_13796,N_13523,N_13507);
xor U13797 (N_13797,N_13554,N_13514);
nand U13798 (N_13798,N_13572,N_13581);
nand U13799 (N_13799,N_13572,N_13556);
or U13800 (N_13800,N_13777,N_13749);
or U13801 (N_13801,N_13711,N_13781);
nor U13802 (N_13802,N_13699,N_13723);
and U13803 (N_13803,N_13785,N_13752);
or U13804 (N_13804,N_13758,N_13669);
xnor U13805 (N_13805,N_13718,N_13698);
and U13806 (N_13806,N_13693,N_13690);
nor U13807 (N_13807,N_13717,N_13757);
or U13808 (N_13808,N_13755,N_13675);
xor U13809 (N_13809,N_13786,N_13797);
or U13810 (N_13810,N_13673,N_13790);
or U13811 (N_13811,N_13651,N_13659);
nand U13812 (N_13812,N_13671,N_13665);
xor U13813 (N_13813,N_13776,N_13658);
and U13814 (N_13814,N_13736,N_13733);
nor U13815 (N_13815,N_13778,N_13714);
nand U13816 (N_13816,N_13783,N_13697);
and U13817 (N_13817,N_13687,N_13799);
and U13818 (N_13818,N_13760,N_13789);
or U13819 (N_13819,N_13731,N_13674);
or U13820 (N_13820,N_13771,N_13684);
and U13821 (N_13821,N_13670,N_13650);
nand U13822 (N_13822,N_13732,N_13796);
nand U13823 (N_13823,N_13729,N_13748);
xnor U13824 (N_13824,N_13681,N_13740);
xor U13825 (N_13825,N_13759,N_13677);
nand U13826 (N_13826,N_13739,N_13792);
nand U13827 (N_13827,N_13712,N_13662);
nor U13828 (N_13828,N_13657,N_13691);
or U13829 (N_13829,N_13705,N_13680);
or U13830 (N_13830,N_13751,N_13703);
nand U13831 (N_13831,N_13767,N_13768);
or U13832 (N_13832,N_13769,N_13761);
nor U13833 (N_13833,N_13772,N_13694);
nand U13834 (N_13834,N_13721,N_13728);
or U13835 (N_13835,N_13676,N_13747);
and U13836 (N_13836,N_13734,N_13793);
xor U13837 (N_13837,N_13730,N_13738);
nor U13838 (N_13838,N_13754,N_13794);
or U13839 (N_13839,N_13689,N_13745);
nand U13840 (N_13840,N_13780,N_13656);
nor U13841 (N_13841,N_13688,N_13765);
or U13842 (N_13842,N_13775,N_13716);
xnor U13843 (N_13843,N_13737,N_13666);
nor U13844 (N_13844,N_13795,N_13722);
nand U13845 (N_13845,N_13741,N_13696);
nand U13846 (N_13846,N_13764,N_13713);
nor U13847 (N_13847,N_13720,N_13791);
or U13848 (N_13848,N_13726,N_13743);
xor U13849 (N_13849,N_13685,N_13679);
nand U13850 (N_13850,N_13709,N_13766);
or U13851 (N_13851,N_13655,N_13700);
nand U13852 (N_13852,N_13742,N_13710);
and U13853 (N_13853,N_13750,N_13653);
or U13854 (N_13854,N_13784,N_13708);
or U13855 (N_13855,N_13763,N_13664);
or U13856 (N_13856,N_13692,N_13756);
nor U13857 (N_13857,N_13744,N_13678);
xor U13858 (N_13858,N_13683,N_13701);
nand U13859 (N_13859,N_13773,N_13682);
and U13860 (N_13860,N_13753,N_13667);
nand U13861 (N_13861,N_13654,N_13706);
xnor U13862 (N_13862,N_13663,N_13727);
nor U13863 (N_13863,N_13660,N_13652);
and U13864 (N_13864,N_13715,N_13762);
and U13865 (N_13865,N_13788,N_13724);
or U13866 (N_13866,N_13704,N_13782);
or U13867 (N_13867,N_13787,N_13661);
nand U13868 (N_13868,N_13725,N_13779);
nor U13869 (N_13869,N_13746,N_13672);
nand U13870 (N_13870,N_13702,N_13668);
or U13871 (N_13871,N_13774,N_13798);
nand U13872 (N_13872,N_13695,N_13735);
nand U13873 (N_13873,N_13770,N_13719);
xor U13874 (N_13874,N_13707,N_13686);
and U13875 (N_13875,N_13784,N_13731);
and U13876 (N_13876,N_13738,N_13712);
xnor U13877 (N_13877,N_13653,N_13767);
nand U13878 (N_13878,N_13709,N_13679);
xnor U13879 (N_13879,N_13697,N_13711);
xor U13880 (N_13880,N_13781,N_13750);
xnor U13881 (N_13881,N_13662,N_13700);
nand U13882 (N_13882,N_13684,N_13731);
or U13883 (N_13883,N_13735,N_13668);
nor U13884 (N_13884,N_13782,N_13752);
nand U13885 (N_13885,N_13715,N_13768);
nor U13886 (N_13886,N_13799,N_13763);
nand U13887 (N_13887,N_13690,N_13651);
and U13888 (N_13888,N_13772,N_13734);
xnor U13889 (N_13889,N_13693,N_13755);
nor U13890 (N_13890,N_13794,N_13650);
nor U13891 (N_13891,N_13660,N_13736);
or U13892 (N_13892,N_13695,N_13716);
and U13893 (N_13893,N_13668,N_13673);
nor U13894 (N_13894,N_13730,N_13719);
nor U13895 (N_13895,N_13657,N_13738);
and U13896 (N_13896,N_13766,N_13694);
nor U13897 (N_13897,N_13750,N_13771);
and U13898 (N_13898,N_13782,N_13699);
nand U13899 (N_13899,N_13663,N_13684);
and U13900 (N_13900,N_13660,N_13654);
and U13901 (N_13901,N_13732,N_13714);
and U13902 (N_13902,N_13760,N_13681);
nand U13903 (N_13903,N_13737,N_13774);
or U13904 (N_13904,N_13724,N_13743);
nor U13905 (N_13905,N_13797,N_13783);
nor U13906 (N_13906,N_13709,N_13660);
and U13907 (N_13907,N_13698,N_13710);
nor U13908 (N_13908,N_13786,N_13728);
and U13909 (N_13909,N_13683,N_13659);
and U13910 (N_13910,N_13740,N_13799);
nand U13911 (N_13911,N_13679,N_13768);
nor U13912 (N_13912,N_13732,N_13742);
nor U13913 (N_13913,N_13753,N_13650);
nand U13914 (N_13914,N_13705,N_13757);
nor U13915 (N_13915,N_13716,N_13785);
nand U13916 (N_13916,N_13689,N_13681);
and U13917 (N_13917,N_13698,N_13766);
or U13918 (N_13918,N_13738,N_13748);
or U13919 (N_13919,N_13706,N_13792);
nand U13920 (N_13920,N_13718,N_13705);
and U13921 (N_13921,N_13734,N_13668);
xor U13922 (N_13922,N_13678,N_13771);
nor U13923 (N_13923,N_13652,N_13755);
nor U13924 (N_13924,N_13755,N_13670);
or U13925 (N_13925,N_13740,N_13668);
nand U13926 (N_13926,N_13790,N_13757);
nand U13927 (N_13927,N_13755,N_13737);
nor U13928 (N_13928,N_13663,N_13694);
and U13929 (N_13929,N_13752,N_13766);
and U13930 (N_13930,N_13689,N_13712);
nor U13931 (N_13931,N_13704,N_13710);
nand U13932 (N_13932,N_13796,N_13775);
nand U13933 (N_13933,N_13681,N_13693);
nand U13934 (N_13934,N_13780,N_13793);
nand U13935 (N_13935,N_13775,N_13693);
nand U13936 (N_13936,N_13725,N_13694);
nor U13937 (N_13937,N_13719,N_13696);
nand U13938 (N_13938,N_13667,N_13709);
xor U13939 (N_13939,N_13752,N_13661);
nand U13940 (N_13940,N_13741,N_13655);
xnor U13941 (N_13941,N_13739,N_13674);
nand U13942 (N_13942,N_13747,N_13731);
or U13943 (N_13943,N_13769,N_13745);
nand U13944 (N_13944,N_13788,N_13722);
and U13945 (N_13945,N_13659,N_13712);
nand U13946 (N_13946,N_13762,N_13787);
and U13947 (N_13947,N_13674,N_13753);
nand U13948 (N_13948,N_13740,N_13651);
and U13949 (N_13949,N_13669,N_13782);
nor U13950 (N_13950,N_13863,N_13800);
nor U13951 (N_13951,N_13865,N_13849);
and U13952 (N_13952,N_13929,N_13934);
nand U13953 (N_13953,N_13896,N_13831);
or U13954 (N_13954,N_13893,N_13888);
nor U13955 (N_13955,N_13946,N_13851);
or U13956 (N_13956,N_13919,N_13869);
nand U13957 (N_13957,N_13852,N_13921);
and U13958 (N_13958,N_13949,N_13948);
nand U13959 (N_13959,N_13828,N_13804);
nor U13960 (N_13960,N_13819,N_13872);
nand U13961 (N_13961,N_13813,N_13871);
xor U13962 (N_13962,N_13923,N_13853);
nor U13963 (N_13963,N_13801,N_13862);
nand U13964 (N_13964,N_13864,N_13944);
nor U13965 (N_13965,N_13889,N_13916);
nor U13966 (N_13966,N_13850,N_13860);
and U13967 (N_13967,N_13809,N_13902);
or U13968 (N_13968,N_13811,N_13906);
nand U13969 (N_13969,N_13841,N_13947);
and U13970 (N_13970,N_13917,N_13897);
and U13971 (N_13971,N_13867,N_13821);
or U13972 (N_13972,N_13855,N_13918);
and U13973 (N_13973,N_13832,N_13942);
nor U13974 (N_13974,N_13812,N_13901);
nand U13975 (N_13975,N_13880,N_13909);
and U13976 (N_13976,N_13892,N_13905);
and U13977 (N_13977,N_13899,N_13915);
or U13978 (N_13978,N_13943,N_13903);
nand U13979 (N_13979,N_13907,N_13856);
or U13980 (N_13980,N_13936,N_13882);
or U13981 (N_13981,N_13830,N_13818);
nand U13982 (N_13982,N_13808,N_13807);
and U13983 (N_13983,N_13913,N_13866);
nand U13984 (N_13984,N_13920,N_13922);
and U13985 (N_13985,N_13904,N_13834);
or U13986 (N_13986,N_13854,N_13900);
nand U13987 (N_13987,N_13824,N_13817);
and U13988 (N_13988,N_13927,N_13885);
nor U13989 (N_13989,N_13816,N_13875);
and U13990 (N_13990,N_13910,N_13810);
nand U13991 (N_13991,N_13928,N_13829);
nand U13992 (N_13992,N_13937,N_13868);
or U13993 (N_13993,N_13814,N_13802);
nand U13994 (N_13994,N_13940,N_13826);
and U13995 (N_13995,N_13881,N_13840);
nand U13996 (N_13996,N_13931,N_13835);
and U13997 (N_13997,N_13898,N_13861);
nand U13998 (N_13998,N_13877,N_13823);
and U13999 (N_13999,N_13805,N_13939);
and U14000 (N_14000,N_13932,N_13891);
or U14001 (N_14001,N_13878,N_13879);
nor U14002 (N_14002,N_13858,N_13925);
nor U14003 (N_14003,N_13836,N_13838);
and U14004 (N_14004,N_13874,N_13803);
or U14005 (N_14005,N_13933,N_13837);
nor U14006 (N_14006,N_13822,N_13833);
nor U14007 (N_14007,N_13876,N_13859);
and U14008 (N_14008,N_13884,N_13908);
nor U14009 (N_14009,N_13844,N_13895);
xnor U14010 (N_14010,N_13843,N_13941);
and U14011 (N_14011,N_13894,N_13870);
nor U14012 (N_14012,N_13886,N_13846);
nor U14013 (N_14013,N_13926,N_13945);
and U14014 (N_14014,N_13873,N_13890);
nor U14015 (N_14015,N_13842,N_13924);
and U14016 (N_14016,N_13815,N_13839);
nand U14017 (N_14017,N_13912,N_13887);
nor U14018 (N_14018,N_13848,N_13847);
nor U14019 (N_14019,N_13938,N_13825);
and U14020 (N_14020,N_13806,N_13827);
nand U14021 (N_14021,N_13857,N_13930);
xnor U14022 (N_14022,N_13845,N_13883);
xnor U14023 (N_14023,N_13935,N_13820);
nand U14024 (N_14024,N_13911,N_13914);
or U14025 (N_14025,N_13810,N_13826);
xnor U14026 (N_14026,N_13896,N_13848);
nor U14027 (N_14027,N_13875,N_13895);
or U14028 (N_14028,N_13945,N_13914);
xnor U14029 (N_14029,N_13891,N_13947);
nor U14030 (N_14030,N_13819,N_13833);
and U14031 (N_14031,N_13826,N_13914);
nor U14032 (N_14032,N_13925,N_13800);
xor U14033 (N_14033,N_13888,N_13923);
or U14034 (N_14034,N_13941,N_13855);
nand U14035 (N_14035,N_13844,N_13801);
or U14036 (N_14036,N_13939,N_13942);
or U14037 (N_14037,N_13910,N_13908);
nand U14038 (N_14038,N_13939,N_13858);
nor U14039 (N_14039,N_13880,N_13847);
and U14040 (N_14040,N_13852,N_13919);
nor U14041 (N_14041,N_13812,N_13928);
nor U14042 (N_14042,N_13844,N_13865);
nor U14043 (N_14043,N_13925,N_13905);
nor U14044 (N_14044,N_13929,N_13836);
and U14045 (N_14045,N_13930,N_13937);
xnor U14046 (N_14046,N_13811,N_13858);
nor U14047 (N_14047,N_13822,N_13935);
nand U14048 (N_14048,N_13824,N_13910);
and U14049 (N_14049,N_13881,N_13943);
and U14050 (N_14050,N_13935,N_13864);
and U14051 (N_14051,N_13931,N_13949);
and U14052 (N_14052,N_13891,N_13882);
and U14053 (N_14053,N_13874,N_13804);
and U14054 (N_14054,N_13912,N_13805);
and U14055 (N_14055,N_13909,N_13924);
or U14056 (N_14056,N_13825,N_13829);
xnor U14057 (N_14057,N_13940,N_13815);
nand U14058 (N_14058,N_13837,N_13911);
and U14059 (N_14059,N_13927,N_13850);
and U14060 (N_14060,N_13834,N_13887);
nor U14061 (N_14061,N_13893,N_13903);
or U14062 (N_14062,N_13895,N_13945);
xor U14063 (N_14063,N_13941,N_13811);
and U14064 (N_14064,N_13823,N_13822);
or U14065 (N_14065,N_13823,N_13811);
nand U14066 (N_14066,N_13937,N_13898);
and U14067 (N_14067,N_13835,N_13855);
and U14068 (N_14068,N_13837,N_13851);
nor U14069 (N_14069,N_13925,N_13840);
nor U14070 (N_14070,N_13828,N_13882);
nor U14071 (N_14071,N_13882,N_13821);
nand U14072 (N_14072,N_13896,N_13890);
or U14073 (N_14073,N_13808,N_13865);
nor U14074 (N_14074,N_13894,N_13852);
and U14075 (N_14075,N_13855,N_13809);
or U14076 (N_14076,N_13860,N_13830);
nor U14077 (N_14077,N_13801,N_13942);
and U14078 (N_14078,N_13875,N_13910);
nand U14079 (N_14079,N_13936,N_13914);
or U14080 (N_14080,N_13904,N_13852);
or U14081 (N_14081,N_13814,N_13860);
nor U14082 (N_14082,N_13855,N_13881);
nand U14083 (N_14083,N_13910,N_13912);
and U14084 (N_14084,N_13893,N_13855);
or U14085 (N_14085,N_13934,N_13866);
and U14086 (N_14086,N_13883,N_13825);
or U14087 (N_14087,N_13874,N_13839);
or U14088 (N_14088,N_13932,N_13842);
nor U14089 (N_14089,N_13911,N_13820);
or U14090 (N_14090,N_13811,N_13853);
and U14091 (N_14091,N_13864,N_13819);
and U14092 (N_14092,N_13939,N_13911);
xnor U14093 (N_14093,N_13930,N_13881);
or U14094 (N_14094,N_13918,N_13842);
nand U14095 (N_14095,N_13855,N_13859);
nor U14096 (N_14096,N_13879,N_13829);
or U14097 (N_14097,N_13874,N_13901);
and U14098 (N_14098,N_13893,N_13837);
or U14099 (N_14099,N_13927,N_13886);
and U14100 (N_14100,N_14003,N_14065);
or U14101 (N_14101,N_14018,N_14032);
nand U14102 (N_14102,N_13969,N_14012);
xnor U14103 (N_14103,N_14078,N_14082);
or U14104 (N_14104,N_14056,N_14016);
and U14105 (N_14105,N_14044,N_14052);
xor U14106 (N_14106,N_13997,N_13955);
or U14107 (N_14107,N_14015,N_14086);
nand U14108 (N_14108,N_14030,N_14099);
nor U14109 (N_14109,N_14061,N_14046);
and U14110 (N_14110,N_13987,N_14013);
and U14111 (N_14111,N_14010,N_13960);
nor U14112 (N_14112,N_13982,N_13976);
and U14113 (N_14113,N_14024,N_14088);
nor U14114 (N_14114,N_14017,N_14026);
or U14115 (N_14115,N_13978,N_14069);
and U14116 (N_14116,N_14001,N_13986);
nor U14117 (N_14117,N_13983,N_14094);
nand U14118 (N_14118,N_14090,N_14093);
and U14119 (N_14119,N_13972,N_14058);
and U14120 (N_14120,N_13981,N_13963);
or U14121 (N_14121,N_13995,N_13991);
nand U14122 (N_14122,N_14051,N_13998);
nand U14123 (N_14123,N_14047,N_13968);
and U14124 (N_14124,N_14073,N_13965);
nor U14125 (N_14125,N_14079,N_14048);
xnor U14126 (N_14126,N_14080,N_14040);
nor U14127 (N_14127,N_14083,N_14011);
nor U14128 (N_14128,N_14004,N_14055);
nand U14129 (N_14129,N_14045,N_14054);
xnor U14130 (N_14130,N_14041,N_13993);
or U14131 (N_14131,N_14008,N_14059);
nor U14132 (N_14132,N_13989,N_14025);
nor U14133 (N_14133,N_14060,N_14087);
xnor U14134 (N_14134,N_14057,N_13980);
nand U14135 (N_14135,N_14072,N_14029);
nand U14136 (N_14136,N_13977,N_14089);
nand U14137 (N_14137,N_13954,N_14019);
or U14138 (N_14138,N_14053,N_13975);
and U14139 (N_14139,N_14035,N_14020);
nand U14140 (N_14140,N_13952,N_13967);
xor U14141 (N_14141,N_14021,N_13970);
nand U14142 (N_14142,N_13957,N_14014);
or U14143 (N_14143,N_14076,N_14007);
nor U14144 (N_14144,N_14098,N_13992);
nor U14145 (N_14145,N_13999,N_14006);
nor U14146 (N_14146,N_14074,N_14034);
nand U14147 (N_14147,N_14023,N_13984);
nand U14148 (N_14148,N_14042,N_14064);
or U14149 (N_14149,N_14049,N_14027);
nand U14150 (N_14150,N_13964,N_13959);
or U14151 (N_14151,N_13994,N_14081);
and U14152 (N_14152,N_14075,N_14009);
or U14153 (N_14153,N_14066,N_14033);
xor U14154 (N_14154,N_13988,N_14095);
nor U14155 (N_14155,N_14070,N_14031);
xor U14156 (N_14156,N_13966,N_13961);
nand U14157 (N_14157,N_14071,N_14005);
nor U14158 (N_14158,N_13958,N_14002);
and U14159 (N_14159,N_13996,N_13985);
nor U14160 (N_14160,N_14037,N_13956);
nor U14161 (N_14161,N_14068,N_14039);
or U14162 (N_14162,N_14067,N_14043);
nor U14163 (N_14163,N_13962,N_14038);
nor U14164 (N_14164,N_14050,N_14022);
and U14165 (N_14165,N_14091,N_14097);
nor U14166 (N_14166,N_13950,N_13990);
and U14167 (N_14167,N_13951,N_13953);
nand U14168 (N_14168,N_13973,N_14085);
or U14169 (N_14169,N_14036,N_13979);
nand U14170 (N_14170,N_14096,N_14028);
or U14171 (N_14171,N_14077,N_14084);
or U14172 (N_14172,N_13974,N_14000);
and U14173 (N_14173,N_14062,N_14063);
nor U14174 (N_14174,N_13971,N_14092);
nand U14175 (N_14175,N_14006,N_14026);
xnor U14176 (N_14176,N_13991,N_14054);
xor U14177 (N_14177,N_14084,N_14091);
nor U14178 (N_14178,N_14040,N_13955);
xnor U14179 (N_14179,N_14022,N_14029);
nor U14180 (N_14180,N_13950,N_14066);
nand U14181 (N_14181,N_14049,N_14052);
and U14182 (N_14182,N_14082,N_14005);
nand U14183 (N_14183,N_13956,N_13993);
xor U14184 (N_14184,N_14010,N_14035);
and U14185 (N_14185,N_14098,N_14095);
or U14186 (N_14186,N_13951,N_14042);
or U14187 (N_14187,N_14094,N_14086);
xnor U14188 (N_14188,N_14015,N_14016);
or U14189 (N_14189,N_14039,N_14088);
nand U14190 (N_14190,N_13959,N_13990);
or U14191 (N_14191,N_14029,N_14001);
or U14192 (N_14192,N_13985,N_13973);
and U14193 (N_14193,N_14022,N_13978);
and U14194 (N_14194,N_14089,N_13953);
nor U14195 (N_14195,N_14077,N_13956);
nor U14196 (N_14196,N_14068,N_14093);
or U14197 (N_14197,N_13985,N_14064);
nor U14198 (N_14198,N_14072,N_14098);
nand U14199 (N_14199,N_14049,N_14006);
nand U14200 (N_14200,N_14067,N_14078);
or U14201 (N_14201,N_14065,N_13998);
nor U14202 (N_14202,N_14035,N_13992);
or U14203 (N_14203,N_14068,N_14099);
nor U14204 (N_14204,N_14064,N_14004);
nor U14205 (N_14205,N_14002,N_13950);
or U14206 (N_14206,N_14008,N_14043);
and U14207 (N_14207,N_14006,N_14031);
nand U14208 (N_14208,N_14006,N_14042);
nor U14209 (N_14209,N_13966,N_14023);
nand U14210 (N_14210,N_14014,N_14065);
and U14211 (N_14211,N_13962,N_14090);
nand U14212 (N_14212,N_14071,N_14060);
nor U14213 (N_14213,N_14088,N_14097);
xnor U14214 (N_14214,N_14002,N_14098);
nand U14215 (N_14215,N_13974,N_13998);
or U14216 (N_14216,N_14086,N_14098);
nand U14217 (N_14217,N_13981,N_14005);
nor U14218 (N_14218,N_13994,N_14088);
and U14219 (N_14219,N_14079,N_13987);
and U14220 (N_14220,N_14063,N_14060);
or U14221 (N_14221,N_14021,N_14071);
nand U14222 (N_14222,N_14083,N_13997);
nor U14223 (N_14223,N_13990,N_14028);
or U14224 (N_14224,N_14035,N_14060);
nand U14225 (N_14225,N_14022,N_13965);
nand U14226 (N_14226,N_14040,N_14013);
or U14227 (N_14227,N_14098,N_14001);
and U14228 (N_14228,N_13958,N_13965);
or U14229 (N_14229,N_13958,N_14075);
nor U14230 (N_14230,N_14033,N_14029);
or U14231 (N_14231,N_14040,N_13973);
and U14232 (N_14232,N_14045,N_13963);
and U14233 (N_14233,N_14046,N_14018);
nor U14234 (N_14234,N_14022,N_13982);
nand U14235 (N_14235,N_13983,N_13950);
nor U14236 (N_14236,N_14081,N_14075);
nor U14237 (N_14237,N_14016,N_13977);
and U14238 (N_14238,N_14045,N_14096);
xor U14239 (N_14239,N_13952,N_14022);
or U14240 (N_14240,N_13982,N_14047);
nor U14241 (N_14241,N_14012,N_14028);
nand U14242 (N_14242,N_13974,N_13960);
xnor U14243 (N_14243,N_13984,N_14045);
or U14244 (N_14244,N_14043,N_14090);
and U14245 (N_14245,N_14000,N_13979);
nor U14246 (N_14246,N_14015,N_14034);
nand U14247 (N_14247,N_14039,N_13993);
nand U14248 (N_14248,N_13989,N_14094);
nand U14249 (N_14249,N_14055,N_13976);
or U14250 (N_14250,N_14134,N_14193);
nor U14251 (N_14251,N_14203,N_14244);
nand U14252 (N_14252,N_14122,N_14131);
or U14253 (N_14253,N_14169,N_14218);
or U14254 (N_14254,N_14128,N_14160);
or U14255 (N_14255,N_14240,N_14100);
nand U14256 (N_14256,N_14147,N_14148);
and U14257 (N_14257,N_14127,N_14198);
nor U14258 (N_14258,N_14199,N_14186);
and U14259 (N_14259,N_14145,N_14138);
and U14260 (N_14260,N_14158,N_14235);
nor U14261 (N_14261,N_14130,N_14227);
nand U14262 (N_14262,N_14179,N_14137);
nor U14263 (N_14263,N_14230,N_14216);
and U14264 (N_14264,N_14117,N_14205);
and U14265 (N_14265,N_14183,N_14237);
nand U14266 (N_14266,N_14223,N_14239);
xnor U14267 (N_14267,N_14207,N_14221);
nand U14268 (N_14268,N_14104,N_14157);
nand U14269 (N_14269,N_14125,N_14204);
and U14270 (N_14270,N_14119,N_14167);
and U14271 (N_14271,N_14110,N_14202);
nand U14272 (N_14272,N_14133,N_14180);
xor U14273 (N_14273,N_14236,N_14114);
xnor U14274 (N_14274,N_14209,N_14220);
or U14275 (N_14275,N_14124,N_14222);
nand U14276 (N_14276,N_14159,N_14109);
nand U14277 (N_14277,N_14155,N_14185);
and U14278 (N_14278,N_14108,N_14211);
nand U14279 (N_14279,N_14201,N_14247);
and U14280 (N_14280,N_14233,N_14187);
and U14281 (N_14281,N_14245,N_14243);
and U14282 (N_14282,N_14139,N_14214);
xnor U14283 (N_14283,N_14142,N_14162);
or U14284 (N_14284,N_14234,N_14150);
nand U14285 (N_14285,N_14215,N_14118);
nand U14286 (N_14286,N_14144,N_14165);
nand U14287 (N_14287,N_14192,N_14136);
nor U14288 (N_14288,N_14101,N_14241);
xor U14289 (N_14289,N_14174,N_14184);
and U14290 (N_14290,N_14103,N_14248);
or U14291 (N_14291,N_14102,N_14189);
and U14292 (N_14292,N_14229,N_14123);
and U14293 (N_14293,N_14213,N_14140);
nor U14294 (N_14294,N_14152,N_14132);
xor U14295 (N_14295,N_14176,N_14194);
xor U14296 (N_14296,N_14195,N_14197);
or U14297 (N_14297,N_14170,N_14238);
nor U14298 (N_14298,N_14166,N_14224);
nand U14299 (N_14299,N_14190,N_14141);
or U14300 (N_14300,N_14212,N_14210);
and U14301 (N_14301,N_14126,N_14219);
or U14302 (N_14302,N_14107,N_14168);
nand U14303 (N_14303,N_14161,N_14129);
nand U14304 (N_14304,N_14106,N_14151);
or U14305 (N_14305,N_14177,N_14156);
and U14306 (N_14306,N_14112,N_14172);
nand U14307 (N_14307,N_14171,N_14188);
or U14308 (N_14308,N_14178,N_14249);
xor U14309 (N_14309,N_14191,N_14121);
and U14310 (N_14310,N_14232,N_14182);
nor U14311 (N_14311,N_14164,N_14196);
nor U14312 (N_14312,N_14163,N_14225);
and U14313 (N_14313,N_14173,N_14146);
nand U14314 (N_14314,N_14231,N_14115);
nor U14315 (N_14315,N_14208,N_14154);
nand U14316 (N_14316,N_14246,N_14116);
or U14317 (N_14317,N_14200,N_14111);
and U14318 (N_14318,N_14242,N_14135);
and U14319 (N_14319,N_14228,N_14149);
nor U14320 (N_14320,N_14217,N_14153);
nand U14321 (N_14321,N_14143,N_14226);
or U14322 (N_14322,N_14181,N_14120);
xor U14323 (N_14323,N_14105,N_14206);
or U14324 (N_14324,N_14113,N_14175);
nand U14325 (N_14325,N_14246,N_14134);
or U14326 (N_14326,N_14234,N_14126);
or U14327 (N_14327,N_14240,N_14133);
or U14328 (N_14328,N_14215,N_14155);
xor U14329 (N_14329,N_14104,N_14224);
nand U14330 (N_14330,N_14131,N_14218);
xnor U14331 (N_14331,N_14113,N_14156);
nand U14332 (N_14332,N_14216,N_14109);
nor U14333 (N_14333,N_14230,N_14210);
nand U14334 (N_14334,N_14129,N_14112);
and U14335 (N_14335,N_14183,N_14109);
or U14336 (N_14336,N_14122,N_14218);
nand U14337 (N_14337,N_14170,N_14225);
xor U14338 (N_14338,N_14184,N_14142);
nor U14339 (N_14339,N_14129,N_14245);
and U14340 (N_14340,N_14150,N_14166);
nor U14341 (N_14341,N_14234,N_14141);
nand U14342 (N_14342,N_14214,N_14229);
nand U14343 (N_14343,N_14245,N_14162);
and U14344 (N_14344,N_14219,N_14215);
nand U14345 (N_14345,N_14130,N_14155);
xnor U14346 (N_14346,N_14129,N_14108);
xnor U14347 (N_14347,N_14195,N_14184);
nand U14348 (N_14348,N_14233,N_14203);
nand U14349 (N_14349,N_14164,N_14142);
or U14350 (N_14350,N_14195,N_14175);
nor U14351 (N_14351,N_14106,N_14208);
and U14352 (N_14352,N_14245,N_14130);
or U14353 (N_14353,N_14175,N_14200);
nand U14354 (N_14354,N_14209,N_14111);
nor U14355 (N_14355,N_14103,N_14107);
and U14356 (N_14356,N_14117,N_14187);
nand U14357 (N_14357,N_14121,N_14216);
or U14358 (N_14358,N_14221,N_14235);
or U14359 (N_14359,N_14108,N_14133);
or U14360 (N_14360,N_14203,N_14221);
nand U14361 (N_14361,N_14208,N_14186);
and U14362 (N_14362,N_14121,N_14156);
nand U14363 (N_14363,N_14188,N_14202);
nand U14364 (N_14364,N_14209,N_14186);
and U14365 (N_14365,N_14191,N_14159);
nand U14366 (N_14366,N_14249,N_14203);
nand U14367 (N_14367,N_14244,N_14147);
nor U14368 (N_14368,N_14205,N_14224);
or U14369 (N_14369,N_14111,N_14225);
nand U14370 (N_14370,N_14248,N_14142);
or U14371 (N_14371,N_14216,N_14141);
and U14372 (N_14372,N_14207,N_14170);
nand U14373 (N_14373,N_14145,N_14118);
or U14374 (N_14374,N_14143,N_14169);
nor U14375 (N_14375,N_14220,N_14217);
and U14376 (N_14376,N_14183,N_14166);
xnor U14377 (N_14377,N_14245,N_14158);
or U14378 (N_14378,N_14231,N_14142);
nand U14379 (N_14379,N_14169,N_14175);
and U14380 (N_14380,N_14137,N_14200);
nor U14381 (N_14381,N_14191,N_14218);
nor U14382 (N_14382,N_14103,N_14177);
nand U14383 (N_14383,N_14113,N_14234);
nor U14384 (N_14384,N_14156,N_14115);
nand U14385 (N_14385,N_14120,N_14153);
and U14386 (N_14386,N_14204,N_14140);
nor U14387 (N_14387,N_14176,N_14204);
or U14388 (N_14388,N_14170,N_14158);
nor U14389 (N_14389,N_14124,N_14123);
xnor U14390 (N_14390,N_14246,N_14224);
nor U14391 (N_14391,N_14187,N_14196);
and U14392 (N_14392,N_14175,N_14114);
nor U14393 (N_14393,N_14179,N_14222);
nor U14394 (N_14394,N_14233,N_14241);
and U14395 (N_14395,N_14131,N_14249);
or U14396 (N_14396,N_14190,N_14152);
xor U14397 (N_14397,N_14144,N_14124);
nand U14398 (N_14398,N_14148,N_14209);
and U14399 (N_14399,N_14140,N_14136);
and U14400 (N_14400,N_14330,N_14358);
nor U14401 (N_14401,N_14399,N_14308);
nor U14402 (N_14402,N_14262,N_14251);
xor U14403 (N_14403,N_14398,N_14278);
xnor U14404 (N_14404,N_14311,N_14359);
nor U14405 (N_14405,N_14356,N_14272);
nor U14406 (N_14406,N_14310,N_14287);
nand U14407 (N_14407,N_14261,N_14275);
xor U14408 (N_14408,N_14294,N_14268);
and U14409 (N_14409,N_14352,N_14302);
and U14410 (N_14410,N_14291,N_14269);
nand U14411 (N_14411,N_14381,N_14342);
or U14412 (N_14412,N_14367,N_14260);
and U14413 (N_14413,N_14364,N_14267);
nand U14414 (N_14414,N_14341,N_14327);
nor U14415 (N_14415,N_14321,N_14313);
and U14416 (N_14416,N_14351,N_14375);
nor U14417 (N_14417,N_14271,N_14304);
nand U14418 (N_14418,N_14376,N_14334);
nand U14419 (N_14419,N_14284,N_14357);
nand U14420 (N_14420,N_14360,N_14259);
and U14421 (N_14421,N_14368,N_14333);
and U14422 (N_14422,N_14331,N_14325);
nand U14423 (N_14423,N_14343,N_14288);
nor U14424 (N_14424,N_14329,N_14257);
or U14425 (N_14425,N_14350,N_14253);
and U14426 (N_14426,N_14309,N_14322);
xnor U14427 (N_14427,N_14361,N_14396);
and U14428 (N_14428,N_14323,N_14346);
nor U14429 (N_14429,N_14389,N_14395);
or U14430 (N_14430,N_14254,N_14377);
nor U14431 (N_14431,N_14374,N_14289);
nor U14432 (N_14432,N_14305,N_14281);
nand U14433 (N_14433,N_14348,N_14392);
and U14434 (N_14434,N_14298,N_14336);
and U14435 (N_14435,N_14293,N_14332);
and U14436 (N_14436,N_14378,N_14372);
nor U14437 (N_14437,N_14353,N_14382);
and U14438 (N_14438,N_14383,N_14393);
and U14439 (N_14439,N_14264,N_14379);
nand U14440 (N_14440,N_14397,N_14344);
nor U14441 (N_14441,N_14285,N_14337);
and U14442 (N_14442,N_14290,N_14282);
or U14443 (N_14443,N_14283,N_14354);
or U14444 (N_14444,N_14306,N_14369);
or U14445 (N_14445,N_14265,N_14320);
and U14446 (N_14446,N_14385,N_14324);
nor U14447 (N_14447,N_14340,N_14373);
and U14448 (N_14448,N_14349,N_14316);
nand U14449 (N_14449,N_14391,N_14386);
or U14450 (N_14450,N_14263,N_14345);
nand U14451 (N_14451,N_14280,N_14266);
nor U14452 (N_14452,N_14328,N_14273);
or U14453 (N_14453,N_14303,N_14371);
nand U14454 (N_14454,N_14318,N_14286);
or U14455 (N_14455,N_14295,N_14380);
nand U14456 (N_14456,N_14388,N_14312);
xor U14457 (N_14457,N_14362,N_14317);
or U14458 (N_14458,N_14252,N_14363);
or U14459 (N_14459,N_14296,N_14319);
nand U14460 (N_14460,N_14299,N_14274);
xor U14461 (N_14461,N_14366,N_14258);
and U14462 (N_14462,N_14390,N_14326);
nand U14463 (N_14463,N_14314,N_14255);
nand U14464 (N_14464,N_14339,N_14394);
nand U14465 (N_14465,N_14250,N_14300);
nand U14466 (N_14466,N_14370,N_14270);
nand U14467 (N_14467,N_14276,N_14384);
xnor U14468 (N_14468,N_14297,N_14307);
nand U14469 (N_14469,N_14315,N_14387);
nand U14470 (N_14470,N_14355,N_14365);
nand U14471 (N_14471,N_14338,N_14292);
nand U14472 (N_14472,N_14277,N_14301);
nand U14473 (N_14473,N_14335,N_14279);
nand U14474 (N_14474,N_14347,N_14256);
and U14475 (N_14475,N_14342,N_14388);
nand U14476 (N_14476,N_14396,N_14324);
xor U14477 (N_14477,N_14383,N_14281);
nand U14478 (N_14478,N_14351,N_14343);
and U14479 (N_14479,N_14255,N_14265);
and U14480 (N_14480,N_14306,N_14382);
nand U14481 (N_14481,N_14337,N_14381);
nor U14482 (N_14482,N_14349,N_14262);
or U14483 (N_14483,N_14337,N_14308);
nor U14484 (N_14484,N_14346,N_14351);
or U14485 (N_14485,N_14296,N_14259);
nor U14486 (N_14486,N_14309,N_14327);
xnor U14487 (N_14487,N_14306,N_14314);
or U14488 (N_14488,N_14391,N_14344);
or U14489 (N_14489,N_14290,N_14289);
or U14490 (N_14490,N_14256,N_14375);
nor U14491 (N_14491,N_14317,N_14370);
nand U14492 (N_14492,N_14318,N_14280);
or U14493 (N_14493,N_14369,N_14390);
nor U14494 (N_14494,N_14345,N_14271);
nand U14495 (N_14495,N_14375,N_14282);
or U14496 (N_14496,N_14281,N_14374);
nand U14497 (N_14497,N_14277,N_14330);
and U14498 (N_14498,N_14353,N_14311);
or U14499 (N_14499,N_14350,N_14307);
nand U14500 (N_14500,N_14256,N_14329);
or U14501 (N_14501,N_14346,N_14389);
nand U14502 (N_14502,N_14349,N_14397);
or U14503 (N_14503,N_14319,N_14368);
xnor U14504 (N_14504,N_14251,N_14339);
nor U14505 (N_14505,N_14357,N_14270);
nand U14506 (N_14506,N_14264,N_14316);
and U14507 (N_14507,N_14318,N_14335);
and U14508 (N_14508,N_14363,N_14328);
nand U14509 (N_14509,N_14389,N_14317);
nor U14510 (N_14510,N_14316,N_14330);
nor U14511 (N_14511,N_14305,N_14386);
and U14512 (N_14512,N_14340,N_14298);
and U14513 (N_14513,N_14281,N_14345);
nand U14514 (N_14514,N_14359,N_14390);
nor U14515 (N_14515,N_14339,N_14286);
and U14516 (N_14516,N_14264,N_14361);
and U14517 (N_14517,N_14269,N_14330);
and U14518 (N_14518,N_14366,N_14371);
nor U14519 (N_14519,N_14280,N_14327);
nand U14520 (N_14520,N_14287,N_14311);
nand U14521 (N_14521,N_14354,N_14371);
nor U14522 (N_14522,N_14350,N_14397);
xnor U14523 (N_14523,N_14323,N_14287);
nor U14524 (N_14524,N_14350,N_14368);
nand U14525 (N_14525,N_14353,N_14293);
or U14526 (N_14526,N_14309,N_14371);
and U14527 (N_14527,N_14345,N_14332);
or U14528 (N_14528,N_14375,N_14310);
xor U14529 (N_14529,N_14331,N_14293);
nand U14530 (N_14530,N_14340,N_14348);
nand U14531 (N_14531,N_14317,N_14387);
nand U14532 (N_14532,N_14318,N_14294);
nand U14533 (N_14533,N_14381,N_14324);
and U14534 (N_14534,N_14256,N_14359);
nand U14535 (N_14535,N_14381,N_14361);
and U14536 (N_14536,N_14325,N_14393);
and U14537 (N_14537,N_14323,N_14349);
or U14538 (N_14538,N_14392,N_14351);
nand U14539 (N_14539,N_14368,N_14329);
nor U14540 (N_14540,N_14329,N_14327);
nand U14541 (N_14541,N_14289,N_14254);
and U14542 (N_14542,N_14372,N_14270);
nand U14543 (N_14543,N_14287,N_14280);
and U14544 (N_14544,N_14318,N_14288);
or U14545 (N_14545,N_14331,N_14258);
or U14546 (N_14546,N_14323,N_14252);
nand U14547 (N_14547,N_14326,N_14361);
nand U14548 (N_14548,N_14353,N_14396);
and U14549 (N_14549,N_14270,N_14310);
nand U14550 (N_14550,N_14490,N_14412);
nand U14551 (N_14551,N_14456,N_14463);
or U14552 (N_14552,N_14421,N_14440);
or U14553 (N_14553,N_14454,N_14447);
or U14554 (N_14554,N_14507,N_14503);
nand U14555 (N_14555,N_14538,N_14488);
nand U14556 (N_14556,N_14427,N_14438);
and U14557 (N_14557,N_14466,N_14467);
nor U14558 (N_14558,N_14497,N_14529);
nand U14559 (N_14559,N_14434,N_14506);
and U14560 (N_14560,N_14522,N_14544);
nand U14561 (N_14561,N_14465,N_14549);
and U14562 (N_14562,N_14539,N_14432);
and U14563 (N_14563,N_14448,N_14401);
nand U14564 (N_14564,N_14457,N_14410);
nand U14565 (N_14565,N_14513,N_14474);
or U14566 (N_14566,N_14403,N_14535);
nand U14567 (N_14567,N_14523,N_14437);
or U14568 (N_14568,N_14458,N_14512);
or U14569 (N_14569,N_14479,N_14422);
nor U14570 (N_14570,N_14477,N_14408);
nand U14571 (N_14571,N_14473,N_14429);
or U14572 (N_14572,N_14433,N_14493);
nand U14573 (N_14573,N_14514,N_14540);
and U14574 (N_14574,N_14472,N_14496);
or U14575 (N_14575,N_14519,N_14436);
and U14576 (N_14576,N_14545,N_14431);
nor U14577 (N_14577,N_14521,N_14486);
or U14578 (N_14578,N_14464,N_14543);
nor U14579 (N_14579,N_14409,N_14527);
nor U14580 (N_14580,N_14536,N_14475);
or U14581 (N_14581,N_14418,N_14469);
and U14582 (N_14582,N_14520,N_14495);
nor U14583 (N_14583,N_14498,N_14483);
or U14584 (N_14584,N_14532,N_14413);
or U14585 (N_14585,N_14443,N_14500);
xor U14586 (N_14586,N_14482,N_14402);
and U14587 (N_14587,N_14445,N_14492);
and U14588 (N_14588,N_14491,N_14450);
or U14589 (N_14589,N_14439,N_14476);
and U14590 (N_14590,N_14547,N_14404);
and U14591 (N_14591,N_14487,N_14459);
nor U14592 (N_14592,N_14419,N_14415);
or U14593 (N_14593,N_14517,N_14504);
or U14594 (N_14594,N_14426,N_14411);
and U14595 (N_14595,N_14533,N_14537);
nand U14596 (N_14596,N_14405,N_14470);
nand U14597 (N_14597,N_14478,N_14518);
or U14598 (N_14598,N_14453,N_14424);
nor U14599 (N_14599,N_14508,N_14420);
nand U14600 (N_14600,N_14510,N_14416);
nand U14601 (N_14601,N_14499,N_14428);
nand U14602 (N_14602,N_14528,N_14541);
or U14603 (N_14603,N_14468,N_14516);
and U14604 (N_14604,N_14423,N_14441);
or U14605 (N_14605,N_14524,N_14501);
or U14606 (N_14606,N_14531,N_14455);
nor U14607 (N_14607,N_14542,N_14484);
or U14608 (N_14608,N_14494,N_14525);
nor U14609 (N_14609,N_14451,N_14471);
and U14610 (N_14610,N_14406,N_14407);
and U14611 (N_14611,N_14509,N_14449);
or U14612 (N_14612,N_14446,N_14430);
nand U14613 (N_14613,N_14452,N_14460);
and U14614 (N_14614,N_14485,N_14546);
nand U14615 (N_14615,N_14435,N_14442);
or U14616 (N_14616,N_14489,N_14526);
nor U14617 (N_14617,N_14400,N_14511);
nand U14618 (N_14618,N_14414,N_14444);
or U14619 (N_14619,N_14480,N_14534);
nor U14620 (N_14620,N_14505,N_14502);
nor U14621 (N_14621,N_14548,N_14417);
or U14622 (N_14622,N_14530,N_14481);
xor U14623 (N_14623,N_14462,N_14425);
or U14624 (N_14624,N_14461,N_14515);
nor U14625 (N_14625,N_14517,N_14425);
or U14626 (N_14626,N_14459,N_14450);
and U14627 (N_14627,N_14460,N_14480);
nor U14628 (N_14628,N_14525,N_14422);
or U14629 (N_14629,N_14431,N_14484);
nor U14630 (N_14630,N_14457,N_14513);
nand U14631 (N_14631,N_14488,N_14537);
nor U14632 (N_14632,N_14484,N_14547);
nand U14633 (N_14633,N_14451,N_14441);
nand U14634 (N_14634,N_14475,N_14505);
and U14635 (N_14635,N_14509,N_14452);
or U14636 (N_14636,N_14438,N_14494);
and U14637 (N_14637,N_14446,N_14467);
and U14638 (N_14638,N_14473,N_14463);
or U14639 (N_14639,N_14505,N_14420);
nand U14640 (N_14640,N_14466,N_14418);
nor U14641 (N_14641,N_14532,N_14418);
xor U14642 (N_14642,N_14465,N_14546);
nand U14643 (N_14643,N_14510,N_14417);
or U14644 (N_14644,N_14491,N_14533);
nor U14645 (N_14645,N_14531,N_14433);
or U14646 (N_14646,N_14497,N_14452);
nand U14647 (N_14647,N_14482,N_14454);
or U14648 (N_14648,N_14465,N_14438);
or U14649 (N_14649,N_14470,N_14484);
nor U14650 (N_14650,N_14446,N_14488);
xor U14651 (N_14651,N_14428,N_14482);
or U14652 (N_14652,N_14427,N_14497);
nor U14653 (N_14653,N_14508,N_14495);
nand U14654 (N_14654,N_14469,N_14482);
nand U14655 (N_14655,N_14455,N_14476);
xnor U14656 (N_14656,N_14540,N_14408);
nor U14657 (N_14657,N_14489,N_14487);
and U14658 (N_14658,N_14511,N_14467);
xor U14659 (N_14659,N_14407,N_14410);
or U14660 (N_14660,N_14518,N_14440);
nand U14661 (N_14661,N_14445,N_14488);
nor U14662 (N_14662,N_14443,N_14477);
xnor U14663 (N_14663,N_14532,N_14498);
nor U14664 (N_14664,N_14459,N_14529);
and U14665 (N_14665,N_14440,N_14413);
nand U14666 (N_14666,N_14426,N_14480);
and U14667 (N_14667,N_14484,N_14452);
nand U14668 (N_14668,N_14413,N_14400);
or U14669 (N_14669,N_14519,N_14478);
or U14670 (N_14670,N_14431,N_14542);
or U14671 (N_14671,N_14426,N_14420);
or U14672 (N_14672,N_14468,N_14486);
and U14673 (N_14673,N_14526,N_14464);
nand U14674 (N_14674,N_14478,N_14411);
nand U14675 (N_14675,N_14505,N_14426);
or U14676 (N_14676,N_14416,N_14525);
or U14677 (N_14677,N_14479,N_14432);
nor U14678 (N_14678,N_14537,N_14412);
and U14679 (N_14679,N_14539,N_14423);
nand U14680 (N_14680,N_14500,N_14525);
nand U14681 (N_14681,N_14525,N_14435);
or U14682 (N_14682,N_14426,N_14463);
and U14683 (N_14683,N_14534,N_14467);
and U14684 (N_14684,N_14548,N_14475);
and U14685 (N_14685,N_14548,N_14479);
and U14686 (N_14686,N_14480,N_14542);
nor U14687 (N_14687,N_14402,N_14423);
nand U14688 (N_14688,N_14404,N_14521);
or U14689 (N_14689,N_14499,N_14522);
or U14690 (N_14690,N_14537,N_14417);
and U14691 (N_14691,N_14546,N_14436);
and U14692 (N_14692,N_14513,N_14530);
nor U14693 (N_14693,N_14425,N_14451);
nand U14694 (N_14694,N_14455,N_14480);
or U14695 (N_14695,N_14480,N_14519);
nand U14696 (N_14696,N_14547,N_14511);
nand U14697 (N_14697,N_14438,N_14514);
nand U14698 (N_14698,N_14469,N_14475);
xor U14699 (N_14699,N_14547,N_14442);
nor U14700 (N_14700,N_14588,N_14687);
xnor U14701 (N_14701,N_14586,N_14660);
xor U14702 (N_14702,N_14632,N_14637);
or U14703 (N_14703,N_14675,N_14620);
nand U14704 (N_14704,N_14564,N_14651);
nor U14705 (N_14705,N_14593,N_14611);
nor U14706 (N_14706,N_14655,N_14619);
nor U14707 (N_14707,N_14666,N_14551);
xor U14708 (N_14708,N_14571,N_14584);
xor U14709 (N_14709,N_14669,N_14635);
nor U14710 (N_14710,N_14668,N_14598);
or U14711 (N_14711,N_14640,N_14605);
nand U14712 (N_14712,N_14657,N_14566);
xor U14713 (N_14713,N_14689,N_14608);
and U14714 (N_14714,N_14656,N_14633);
nor U14715 (N_14715,N_14610,N_14587);
and U14716 (N_14716,N_14557,N_14628);
and U14717 (N_14717,N_14692,N_14562);
nand U14718 (N_14718,N_14648,N_14638);
nor U14719 (N_14719,N_14606,N_14677);
xor U14720 (N_14720,N_14603,N_14630);
and U14721 (N_14721,N_14568,N_14665);
nor U14722 (N_14722,N_14672,N_14686);
nor U14723 (N_14723,N_14644,N_14622);
nor U14724 (N_14724,N_14618,N_14574);
xnor U14725 (N_14725,N_14678,N_14581);
nor U14726 (N_14726,N_14636,N_14600);
or U14727 (N_14727,N_14639,N_14573);
nand U14728 (N_14728,N_14558,N_14662);
nor U14729 (N_14729,N_14627,N_14621);
nor U14730 (N_14730,N_14589,N_14645);
or U14731 (N_14731,N_14694,N_14682);
nor U14732 (N_14732,N_14681,N_14591);
nor U14733 (N_14733,N_14592,N_14577);
nor U14734 (N_14734,N_14623,N_14609);
and U14735 (N_14735,N_14691,N_14646);
nor U14736 (N_14736,N_14601,N_14642);
or U14737 (N_14737,N_14699,N_14583);
or U14738 (N_14738,N_14579,N_14670);
and U14739 (N_14739,N_14597,N_14652);
nand U14740 (N_14740,N_14659,N_14576);
and U14741 (N_14741,N_14679,N_14614);
and U14742 (N_14742,N_14688,N_14553);
nor U14743 (N_14743,N_14599,N_14680);
nand U14744 (N_14744,N_14570,N_14676);
and U14745 (N_14745,N_14596,N_14664);
or U14746 (N_14746,N_14556,N_14634);
nand U14747 (N_14747,N_14561,N_14667);
nand U14748 (N_14748,N_14616,N_14554);
or U14749 (N_14749,N_14590,N_14555);
nor U14750 (N_14750,N_14612,N_14565);
and U14751 (N_14751,N_14641,N_14683);
and U14752 (N_14752,N_14673,N_14684);
nor U14753 (N_14753,N_14582,N_14643);
xor U14754 (N_14754,N_14578,N_14647);
and U14755 (N_14755,N_14580,N_14626);
nand U14756 (N_14756,N_14602,N_14625);
and U14757 (N_14757,N_14697,N_14663);
nand U14758 (N_14758,N_14671,N_14604);
and U14759 (N_14759,N_14615,N_14613);
nand U14760 (N_14760,N_14653,N_14595);
and U14761 (N_14761,N_14654,N_14661);
xnor U14762 (N_14762,N_14696,N_14631);
and U14763 (N_14763,N_14567,N_14693);
and U14764 (N_14764,N_14560,N_14685);
nor U14765 (N_14765,N_14563,N_14695);
nor U14766 (N_14766,N_14585,N_14569);
nand U14767 (N_14767,N_14607,N_14698);
or U14768 (N_14768,N_14572,N_14650);
xor U14769 (N_14769,N_14624,N_14552);
nand U14770 (N_14770,N_14617,N_14594);
or U14771 (N_14771,N_14690,N_14674);
or U14772 (N_14772,N_14649,N_14559);
nor U14773 (N_14773,N_14575,N_14629);
or U14774 (N_14774,N_14658,N_14550);
xnor U14775 (N_14775,N_14658,N_14642);
nor U14776 (N_14776,N_14689,N_14694);
and U14777 (N_14777,N_14557,N_14602);
nor U14778 (N_14778,N_14559,N_14561);
nand U14779 (N_14779,N_14593,N_14614);
and U14780 (N_14780,N_14602,N_14655);
nand U14781 (N_14781,N_14635,N_14693);
nand U14782 (N_14782,N_14650,N_14661);
nor U14783 (N_14783,N_14556,N_14598);
nor U14784 (N_14784,N_14568,N_14699);
nand U14785 (N_14785,N_14647,N_14572);
nand U14786 (N_14786,N_14626,N_14569);
and U14787 (N_14787,N_14570,N_14626);
nor U14788 (N_14788,N_14613,N_14640);
xor U14789 (N_14789,N_14646,N_14650);
nand U14790 (N_14790,N_14642,N_14628);
xnor U14791 (N_14791,N_14648,N_14579);
and U14792 (N_14792,N_14578,N_14639);
nand U14793 (N_14793,N_14592,N_14641);
or U14794 (N_14794,N_14616,N_14644);
and U14795 (N_14795,N_14593,N_14694);
or U14796 (N_14796,N_14626,N_14575);
and U14797 (N_14797,N_14569,N_14587);
xnor U14798 (N_14798,N_14572,N_14590);
and U14799 (N_14799,N_14643,N_14688);
and U14800 (N_14800,N_14563,N_14688);
xor U14801 (N_14801,N_14551,N_14616);
and U14802 (N_14802,N_14694,N_14586);
or U14803 (N_14803,N_14671,N_14615);
nor U14804 (N_14804,N_14654,N_14602);
and U14805 (N_14805,N_14607,N_14631);
nand U14806 (N_14806,N_14672,N_14688);
nor U14807 (N_14807,N_14589,N_14695);
xor U14808 (N_14808,N_14684,N_14557);
nand U14809 (N_14809,N_14617,N_14561);
nor U14810 (N_14810,N_14611,N_14618);
nand U14811 (N_14811,N_14658,N_14647);
or U14812 (N_14812,N_14660,N_14569);
nand U14813 (N_14813,N_14693,N_14654);
nor U14814 (N_14814,N_14676,N_14581);
nand U14815 (N_14815,N_14686,N_14581);
or U14816 (N_14816,N_14591,N_14653);
nand U14817 (N_14817,N_14585,N_14676);
or U14818 (N_14818,N_14643,N_14598);
nand U14819 (N_14819,N_14573,N_14622);
and U14820 (N_14820,N_14591,N_14627);
nand U14821 (N_14821,N_14591,N_14675);
or U14822 (N_14822,N_14662,N_14675);
and U14823 (N_14823,N_14650,N_14612);
nand U14824 (N_14824,N_14645,N_14613);
nor U14825 (N_14825,N_14582,N_14634);
nand U14826 (N_14826,N_14576,N_14630);
xor U14827 (N_14827,N_14683,N_14678);
and U14828 (N_14828,N_14675,N_14598);
nand U14829 (N_14829,N_14653,N_14630);
or U14830 (N_14830,N_14673,N_14693);
nand U14831 (N_14831,N_14678,N_14660);
and U14832 (N_14832,N_14558,N_14643);
nand U14833 (N_14833,N_14578,N_14658);
or U14834 (N_14834,N_14576,N_14638);
xor U14835 (N_14835,N_14626,N_14669);
and U14836 (N_14836,N_14668,N_14599);
or U14837 (N_14837,N_14604,N_14635);
nor U14838 (N_14838,N_14590,N_14681);
nor U14839 (N_14839,N_14628,N_14665);
nand U14840 (N_14840,N_14637,N_14668);
nor U14841 (N_14841,N_14653,N_14570);
and U14842 (N_14842,N_14604,N_14695);
and U14843 (N_14843,N_14604,N_14603);
xor U14844 (N_14844,N_14671,N_14579);
and U14845 (N_14845,N_14625,N_14588);
or U14846 (N_14846,N_14590,N_14689);
or U14847 (N_14847,N_14641,N_14585);
nor U14848 (N_14848,N_14550,N_14614);
nor U14849 (N_14849,N_14553,N_14651);
or U14850 (N_14850,N_14820,N_14833);
nand U14851 (N_14851,N_14705,N_14713);
and U14852 (N_14852,N_14789,N_14840);
and U14853 (N_14853,N_14721,N_14745);
nor U14854 (N_14854,N_14826,N_14783);
nor U14855 (N_14855,N_14706,N_14709);
and U14856 (N_14856,N_14780,N_14844);
nor U14857 (N_14857,N_14843,N_14792);
nor U14858 (N_14858,N_14726,N_14708);
and U14859 (N_14859,N_14725,N_14822);
nand U14860 (N_14860,N_14757,N_14740);
xnor U14861 (N_14861,N_14775,N_14765);
or U14862 (N_14862,N_14785,N_14774);
nor U14863 (N_14863,N_14782,N_14763);
nand U14864 (N_14864,N_14715,N_14716);
and U14865 (N_14865,N_14787,N_14804);
nand U14866 (N_14866,N_14809,N_14735);
nand U14867 (N_14867,N_14835,N_14823);
nand U14868 (N_14868,N_14802,N_14811);
and U14869 (N_14869,N_14751,N_14733);
nand U14870 (N_14870,N_14712,N_14827);
nand U14871 (N_14871,N_14773,N_14825);
nor U14872 (N_14872,N_14776,N_14788);
xnor U14873 (N_14873,N_14846,N_14753);
or U14874 (N_14874,N_14727,N_14808);
xor U14875 (N_14875,N_14800,N_14761);
or U14876 (N_14876,N_14842,N_14828);
and U14877 (N_14877,N_14832,N_14806);
and U14878 (N_14878,N_14817,N_14710);
nor U14879 (N_14879,N_14766,N_14805);
or U14880 (N_14880,N_14724,N_14801);
nor U14881 (N_14881,N_14719,N_14769);
and U14882 (N_14882,N_14836,N_14730);
or U14883 (N_14883,N_14847,N_14772);
nand U14884 (N_14884,N_14704,N_14759);
or U14885 (N_14885,N_14781,N_14750);
nor U14886 (N_14886,N_14746,N_14810);
or U14887 (N_14887,N_14824,N_14830);
or U14888 (N_14888,N_14729,N_14762);
nand U14889 (N_14889,N_14819,N_14786);
xnor U14890 (N_14890,N_14779,N_14731);
and U14891 (N_14891,N_14758,N_14791);
xor U14892 (N_14892,N_14734,N_14702);
nor U14893 (N_14893,N_14807,N_14790);
xnor U14894 (N_14894,N_14818,N_14723);
or U14895 (N_14895,N_14849,N_14738);
xnor U14896 (N_14896,N_14777,N_14747);
and U14897 (N_14897,N_14815,N_14837);
or U14898 (N_14898,N_14794,N_14839);
nand U14899 (N_14899,N_14797,N_14718);
xor U14900 (N_14900,N_14829,N_14814);
and U14901 (N_14901,N_14764,N_14760);
and U14902 (N_14902,N_14793,N_14799);
and U14903 (N_14903,N_14831,N_14771);
or U14904 (N_14904,N_14767,N_14796);
xnor U14905 (N_14905,N_14841,N_14778);
nand U14906 (N_14906,N_14752,N_14845);
or U14907 (N_14907,N_14834,N_14739);
nor U14908 (N_14908,N_14742,N_14728);
and U14909 (N_14909,N_14722,N_14720);
nand U14910 (N_14910,N_14812,N_14754);
xor U14911 (N_14911,N_14816,N_14700);
and U14912 (N_14912,N_14717,N_14703);
or U14913 (N_14913,N_14798,N_14821);
or U14914 (N_14914,N_14756,N_14737);
and U14915 (N_14915,N_14744,N_14701);
and U14916 (N_14916,N_14838,N_14770);
nor U14917 (N_14917,N_14748,N_14755);
xor U14918 (N_14918,N_14741,N_14743);
nor U14919 (N_14919,N_14714,N_14711);
and U14920 (N_14920,N_14784,N_14749);
and U14921 (N_14921,N_14707,N_14803);
nor U14922 (N_14922,N_14795,N_14848);
or U14923 (N_14923,N_14768,N_14732);
nor U14924 (N_14924,N_14813,N_14736);
nand U14925 (N_14925,N_14806,N_14721);
nor U14926 (N_14926,N_14837,N_14772);
xor U14927 (N_14927,N_14753,N_14737);
or U14928 (N_14928,N_14763,N_14807);
or U14929 (N_14929,N_14781,N_14807);
and U14930 (N_14930,N_14718,N_14834);
or U14931 (N_14931,N_14747,N_14754);
or U14932 (N_14932,N_14798,N_14833);
nand U14933 (N_14933,N_14753,N_14769);
nand U14934 (N_14934,N_14786,N_14710);
and U14935 (N_14935,N_14708,N_14753);
nor U14936 (N_14936,N_14837,N_14807);
and U14937 (N_14937,N_14806,N_14742);
nor U14938 (N_14938,N_14786,N_14765);
nor U14939 (N_14939,N_14737,N_14735);
nand U14940 (N_14940,N_14730,N_14722);
or U14941 (N_14941,N_14829,N_14786);
nand U14942 (N_14942,N_14803,N_14701);
and U14943 (N_14943,N_14763,N_14824);
and U14944 (N_14944,N_14847,N_14803);
and U14945 (N_14945,N_14782,N_14762);
nand U14946 (N_14946,N_14793,N_14837);
and U14947 (N_14947,N_14788,N_14792);
and U14948 (N_14948,N_14808,N_14744);
or U14949 (N_14949,N_14801,N_14777);
and U14950 (N_14950,N_14845,N_14806);
nor U14951 (N_14951,N_14771,N_14762);
nand U14952 (N_14952,N_14733,N_14724);
or U14953 (N_14953,N_14753,N_14823);
or U14954 (N_14954,N_14793,N_14786);
nor U14955 (N_14955,N_14777,N_14744);
or U14956 (N_14956,N_14705,N_14848);
nor U14957 (N_14957,N_14775,N_14847);
and U14958 (N_14958,N_14747,N_14706);
nor U14959 (N_14959,N_14817,N_14780);
and U14960 (N_14960,N_14740,N_14739);
nor U14961 (N_14961,N_14739,N_14738);
xor U14962 (N_14962,N_14749,N_14742);
nor U14963 (N_14963,N_14762,N_14827);
nand U14964 (N_14964,N_14800,N_14840);
nor U14965 (N_14965,N_14755,N_14728);
and U14966 (N_14966,N_14770,N_14735);
and U14967 (N_14967,N_14742,N_14714);
and U14968 (N_14968,N_14849,N_14823);
and U14969 (N_14969,N_14762,N_14712);
or U14970 (N_14970,N_14827,N_14768);
nand U14971 (N_14971,N_14818,N_14713);
and U14972 (N_14972,N_14817,N_14830);
nor U14973 (N_14973,N_14756,N_14805);
xnor U14974 (N_14974,N_14732,N_14835);
nand U14975 (N_14975,N_14735,N_14829);
or U14976 (N_14976,N_14765,N_14780);
and U14977 (N_14977,N_14703,N_14770);
and U14978 (N_14978,N_14839,N_14828);
xor U14979 (N_14979,N_14747,N_14712);
nand U14980 (N_14980,N_14712,N_14763);
and U14981 (N_14981,N_14732,N_14713);
and U14982 (N_14982,N_14787,N_14846);
nand U14983 (N_14983,N_14825,N_14720);
and U14984 (N_14984,N_14781,N_14819);
and U14985 (N_14985,N_14833,N_14710);
or U14986 (N_14986,N_14763,N_14836);
or U14987 (N_14987,N_14811,N_14701);
nor U14988 (N_14988,N_14834,N_14806);
nor U14989 (N_14989,N_14845,N_14788);
nand U14990 (N_14990,N_14714,N_14789);
nand U14991 (N_14991,N_14764,N_14814);
or U14992 (N_14992,N_14721,N_14760);
nand U14993 (N_14993,N_14766,N_14748);
nor U14994 (N_14994,N_14765,N_14846);
and U14995 (N_14995,N_14799,N_14741);
xor U14996 (N_14996,N_14707,N_14732);
and U14997 (N_14997,N_14836,N_14806);
nand U14998 (N_14998,N_14849,N_14734);
or U14999 (N_14999,N_14771,N_14758);
nand UO_0 (O_0,N_14852,N_14949);
nand UO_1 (O_1,N_14882,N_14998);
xor UO_2 (O_2,N_14918,N_14991);
and UO_3 (O_3,N_14967,N_14945);
nand UO_4 (O_4,N_14870,N_14965);
or UO_5 (O_5,N_14922,N_14934);
or UO_6 (O_6,N_14974,N_14981);
nor UO_7 (O_7,N_14952,N_14961);
nor UO_8 (O_8,N_14940,N_14871);
nand UO_9 (O_9,N_14976,N_14951);
nand UO_10 (O_10,N_14873,N_14862);
and UO_11 (O_11,N_14968,N_14957);
nor UO_12 (O_12,N_14985,N_14878);
nand UO_13 (O_13,N_14860,N_14912);
nand UO_14 (O_14,N_14863,N_14916);
nor UO_15 (O_15,N_14901,N_14928);
nand UO_16 (O_16,N_14921,N_14902);
nand UO_17 (O_17,N_14954,N_14980);
nor UO_18 (O_18,N_14992,N_14869);
or UO_19 (O_19,N_14899,N_14960);
or UO_20 (O_20,N_14897,N_14861);
or UO_21 (O_21,N_14910,N_14859);
nor UO_22 (O_22,N_14973,N_14854);
nor UO_23 (O_23,N_14975,N_14911);
nand UO_24 (O_24,N_14875,N_14950);
and UO_25 (O_25,N_14903,N_14850);
and UO_26 (O_26,N_14933,N_14892);
or UO_27 (O_27,N_14906,N_14932);
and UO_28 (O_28,N_14956,N_14881);
nand UO_29 (O_29,N_14872,N_14986);
or UO_30 (O_30,N_14885,N_14994);
or UO_31 (O_31,N_14925,N_14941);
and UO_32 (O_32,N_14983,N_14888);
nor UO_33 (O_33,N_14936,N_14977);
or UO_34 (O_34,N_14930,N_14913);
xnor UO_35 (O_35,N_14879,N_14939);
nor UO_36 (O_36,N_14895,N_14864);
nor UO_37 (O_37,N_14890,N_14935);
and UO_38 (O_38,N_14964,N_14953);
nor UO_39 (O_39,N_14943,N_14924);
or UO_40 (O_40,N_14905,N_14857);
xor UO_41 (O_41,N_14937,N_14867);
nor UO_42 (O_42,N_14927,N_14993);
xor UO_43 (O_43,N_14987,N_14963);
nand UO_44 (O_44,N_14900,N_14978);
or UO_45 (O_45,N_14990,N_14989);
and UO_46 (O_46,N_14995,N_14942);
nor UO_47 (O_47,N_14884,N_14877);
nand UO_48 (O_48,N_14887,N_14926);
nand UO_49 (O_49,N_14891,N_14946);
or UO_50 (O_50,N_14979,N_14896);
nand UO_51 (O_51,N_14868,N_14988);
nand UO_52 (O_52,N_14908,N_14889);
nand UO_53 (O_53,N_14904,N_14919);
nor UO_54 (O_54,N_14947,N_14856);
or UO_55 (O_55,N_14959,N_14898);
nand UO_56 (O_56,N_14958,N_14893);
nor UO_57 (O_57,N_14907,N_14915);
nand UO_58 (O_58,N_14909,N_14999);
nand UO_59 (O_59,N_14876,N_14920);
or UO_60 (O_60,N_14883,N_14955);
or UO_61 (O_61,N_14880,N_14948);
or UO_62 (O_62,N_14997,N_14853);
and UO_63 (O_63,N_14866,N_14982);
nand UO_64 (O_64,N_14938,N_14886);
or UO_65 (O_65,N_14962,N_14894);
xor UO_66 (O_66,N_14855,N_14874);
nor UO_67 (O_67,N_14931,N_14996);
or UO_68 (O_68,N_14929,N_14966);
and UO_69 (O_69,N_14984,N_14865);
nand UO_70 (O_70,N_14944,N_14858);
xnor UO_71 (O_71,N_14971,N_14969);
nand UO_72 (O_72,N_14923,N_14914);
or UO_73 (O_73,N_14972,N_14917);
and UO_74 (O_74,N_14851,N_14970);
nand UO_75 (O_75,N_14908,N_14919);
and UO_76 (O_76,N_14978,N_14950);
and UO_77 (O_77,N_14913,N_14872);
and UO_78 (O_78,N_14931,N_14972);
xor UO_79 (O_79,N_14890,N_14865);
nor UO_80 (O_80,N_14917,N_14979);
nor UO_81 (O_81,N_14971,N_14943);
or UO_82 (O_82,N_14976,N_14989);
nand UO_83 (O_83,N_14939,N_14884);
nand UO_84 (O_84,N_14870,N_14900);
or UO_85 (O_85,N_14934,N_14936);
nor UO_86 (O_86,N_14972,N_14907);
or UO_87 (O_87,N_14920,N_14959);
and UO_88 (O_88,N_14894,N_14885);
or UO_89 (O_89,N_14947,N_14930);
and UO_90 (O_90,N_14961,N_14904);
nand UO_91 (O_91,N_14895,N_14887);
or UO_92 (O_92,N_14931,N_14995);
nor UO_93 (O_93,N_14905,N_14895);
and UO_94 (O_94,N_14995,N_14948);
and UO_95 (O_95,N_14950,N_14905);
nand UO_96 (O_96,N_14901,N_14866);
or UO_97 (O_97,N_14891,N_14930);
nand UO_98 (O_98,N_14887,N_14951);
or UO_99 (O_99,N_14874,N_14945);
and UO_100 (O_100,N_14878,N_14993);
xor UO_101 (O_101,N_14924,N_14886);
xor UO_102 (O_102,N_14917,N_14986);
nand UO_103 (O_103,N_14977,N_14909);
xnor UO_104 (O_104,N_14858,N_14984);
and UO_105 (O_105,N_14999,N_14953);
nor UO_106 (O_106,N_14978,N_14870);
nor UO_107 (O_107,N_14892,N_14982);
nand UO_108 (O_108,N_14997,N_14954);
nor UO_109 (O_109,N_14958,N_14948);
nand UO_110 (O_110,N_14852,N_14888);
or UO_111 (O_111,N_14956,N_14867);
and UO_112 (O_112,N_14947,N_14977);
nor UO_113 (O_113,N_14874,N_14956);
and UO_114 (O_114,N_14852,N_14867);
nand UO_115 (O_115,N_14900,N_14926);
and UO_116 (O_116,N_14984,N_14937);
or UO_117 (O_117,N_14892,N_14997);
nor UO_118 (O_118,N_14921,N_14944);
nand UO_119 (O_119,N_14923,N_14983);
and UO_120 (O_120,N_14935,N_14942);
and UO_121 (O_121,N_14852,N_14957);
and UO_122 (O_122,N_14929,N_14932);
and UO_123 (O_123,N_14998,N_14938);
nand UO_124 (O_124,N_14894,N_14953);
nor UO_125 (O_125,N_14935,N_14857);
and UO_126 (O_126,N_14869,N_14870);
nand UO_127 (O_127,N_14859,N_14971);
nand UO_128 (O_128,N_14898,N_14885);
and UO_129 (O_129,N_14856,N_14852);
or UO_130 (O_130,N_14990,N_14916);
nor UO_131 (O_131,N_14855,N_14939);
xnor UO_132 (O_132,N_14975,N_14946);
or UO_133 (O_133,N_14924,N_14986);
and UO_134 (O_134,N_14902,N_14890);
nor UO_135 (O_135,N_14855,N_14978);
xor UO_136 (O_136,N_14902,N_14893);
and UO_137 (O_137,N_14854,N_14974);
nand UO_138 (O_138,N_14948,N_14857);
and UO_139 (O_139,N_14933,N_14891);
xor UO_140 (O_140,N_14887,N_14855);
and UO_141 (O_141,N_14857,N_14934);
or UO_142 (O_142,N_14859,N_14915);
nand UO_143 (O_143,N_14906,N_14985);
nand UO_144 (O_144,N_14896,N_14864);
or UO_145 (O_145,N_14961,N_14986);
and UO_146 (O_146,N_14961,N_14855);
nor UO_147 (O_147,N_14978,N_14909);
and UO_148 (O_148,N_14878,N_14976);
or UO_149 (O_149,N_14933,N_14858);
nor UO_150 (O_150,N_14865,N_14933);
xnor UO_151 (O_151,N_14879,N_14980);
and UO_152 (O_152,N_14855,N_14977);
or UO_153 (O_153,N_14953,N_14998);
xor UO_154 (O_154,N_14888,N_14967);
nor UO_155 (O_155,N_14937,N_14952);
and UO_156 (O_156,N_14905,N_14894);
nor UO_157 (O_157,N_14890,N_14968);
and UO_158 (O_158,N_14947,N_14900);
nor UO_159 (O_159,N_14854,N_14905);
xnor UO_160 (O_160,N_14952,N_14869);
xnor UO_161 (O_161,N_14906,N_14894);
nor UO_162 (O_162,N_14939,N_14853);
xnor UO_163 (O_163,N_14937,N_14916);
nor UO_164 (O_164,N_14994,N_14854);
or UO_165 (O_165,N_14876,N_14974);
xor UO_166 (O_166,N_14852,N_14953);
nor UO_167 (O_167,N_14996,N_14908);
nand UO_168 (O_168,N_14947,N_14986);
nor UO_169 (O_169,N_14898,N_14991);
xor UO_170 (O_170,N_14961,N_14910);
nand UO_171 (O_171,N_14956,N_14924);
or UO_172 (O_172,N_14923,N_14868);
nor UO_173 (O_173,N_14858,N_14917);
and UO_174 (O_174,N_14998,N_14929);
and UO_175 (O_175,N_14853,N_14952);
nor UO_176 (O_176,N_14942,N_14949);
nand UO_177 (O_177,N_14856,N_14921);
nand UO_178 (O_178,N_14887,N_14954);
or UO_179 (O_179,N_14890,N_14864);
xnor UO_180 (O_180,N_14946,N_14854);
nand UO_181 (O_181,N_14906,N_14988);
and UO_182 (O_182,N_14964,N_14892);
and UO_183 (O_183,N_14922,N_14953);
and UO_184 (O_184,N_14882,N_14960);
nor UO_185 (O_185,N_14957,N_14894);
nor UO_186 (O_186,N_14877,N_14931);
xnor UO_187 (O_187,N_14982,N_14934);
nand UO_188 (O_188,N_14852,N_14919);
nand UO_189 (O_189,N_14873,N_14981);
or UO_190 (O_190,N_14953,N_14952);
nand UO_191 (O_191,N_14907,N_14952);
and UO_192 (O_192,N_14904,N_14941);
nor UO_193 (O_193,N_14976,N_14900);
nand UO_194 (O_194,N_14944,N_14857);
and UO_195 (O_195,N_14965,N_14864);
or UO_196 (O_196,N_14950,N_14900);
nand UO_197 (O_197,N_14858,N_14865);
nor UO_198 (O_198,N_14951,N_14921);
nand UO_199 (O_199,N_14988,N_14991);
or UO_200 (O_200,N_14970,N_14874);
nor UO_201 (O_201,N_14995,N_14936);
and UO_202 (O_202,N_14922,N_14899);
xnor UO_203 (O_203,N_14949,N_14962);
or UO_204 (O_204,N_14979,N_14892);
nor UO_205 (O_205,N_14851,N_14934);
or UO_206 (O_206,N_14956,N_14993);
nor UO_207 (O_207,N_14895,N_14857);
nor UO_208 (O_208,N_14859,N_14939);
nand UO_209 (O_209,N_14953,N_14909);
nand UO_210 (O_210,N_14877,N_14948);
or UO_211 (O_211,N_14976,N_14975);
nor UO_212 (O_212,N_14854,N_14995);
nor UO_213 (O_213,N_14958,N_14981);
or UO_214 (O_214,N_14880,N_14919);
and UO_215 (O_215,N_14953,N_14945);
or UO_216 (O_216,N_14961,N_14918);
nor UO_217 (O_217,N_14885,N_14902);
and UO_218 (O_218,N_14936,N_14903);
or UO_219 (O_219,N_14952,N_14920);
nor UO_220 (O_220,N_14858,N_14934);
nor UO_221 (O_221,N_14869,N_14996);
nor UO_222 (O_222,N_14897,N_14877);
xnor UO_223 (O_223,N_14914,N_14984);
and UO_224 (O_224,N_14880,N_14861);
or UO_225 (O_225,N_14904,N_14983);
nand UO_226 (O_226,N_14860,N_14890);
nor UO_227 (O_227,N_14882,N_14984);
nor UO_228 (O_228,N_14999,N_14924);
or UO_229 (O_229,N_14912,N_14872);
and UO_230 (O_230,N_14982,N_14917);
and UO_231 (O_231,N_14874,N_14998);
nand UO_232 (O_232,N_14936,N_14887);
or UO_233 (O_233,N_14932,N_14854);
xnor UO_234 (O_234,N_14942,N_14903);
nor UO_235 (O_235,N_14920,N_14917);
nand UO_236 (O_236,N_14879,N_14928);
or UO_237 (O_237,N_14946,N_14895);
and UO_238 (O_238,N_14962,N_14898);
or UO_239 (O_239,N_14911,N_14989);
xor UO_240 (O_240,N_14932,N_14899);
nor UO_241 (O_241,N_14865,N_14962);
nor UO_242 (O_242,N_14981,N_14895);
and UO_243 (O_243,N_14901,N_14937);
nand UO_244 (O_244,N_14993,N_14991);
nor UO_245 (O_245,N_14877,N_14894);
nor UO_246 (O_246,N_14994,N_14961);
or UO_247 (O_247,N_14959,N_14886);
and UO_248 (O_248,N_14884,N_14861);
nor UO_249 (O_249,N_14868,N_14922);
nor UO_250 (O_250,N_14855,N_14924);
xnor UO_251 (O_251,N_14977,N_14854);
nor UO_252 (O_252,N_14971,N_14938);
nand UO_253 (O_253,N_14871,N_14967);
nand UO_254 (O_254,N_14869,N_14884);
and UO_255 (O_255,N_14995,N_14972);
and UO_256 (O_256,N_14996,N_14917);
or UO_257 (O_257,N_14999,N_14926);
xnor UO_258 (O_258,N_14916,N_14899);
or UO_259 (O_259,N_14887,N_14878);
nor UO_260 (O_260,N_14933,N_14951);
and UO_261 (O_261,N_14855,N_14952);
nor UO_262 (O_262,N_14959,N_14961);
and UO_263 (O_263,N_14889,N_14915);
nand UO_264 (O_264,N_14965,N_14904);
nor UO_265 (O_265,N_14850,N_14899);
nand UO_266 (O_266,N_14876,N_14904);
xor UO_267 (O_267,N_14987,N_14943);
nand UO_268 (O_268,N_14876,N_14968);
and UO_269 (O_269,N_14879,N_14874);
nor UO_270 (O_270,N_14995,N_14879);
or UO_271 (O_271,N_14975,N_14864);
xor UO_272 (O_272,N_14875,N_14904);
or UO_273 (O_273,N_14984,N_14972);
or UO_274 (O_274,N_14924,N_14946);
nor UO_275 (O_275,N_14989,N_14908);
xor UO_276 (O_276,N_14876,N_14941);
nand UO_277 (O_277,N_14905,N_14911);
nand UO_278 (O_278,N_14851,N_14964);
nor UO_279 (O_279,N_14856,N_14977);
nand UO_280 (O_280,N_14988,N_14931);
nor UO_281 (O_281,N_14896,N_14986);
or UO_282 (O_282,N_14872,N_14877);
and UO_283 (O_283,N_14850,N_14951);
or UO_284 (O_284,N_14955,N_14890);
or UO_285 (O_285,N_14867,N_14915);
and UO_286 (O_286,N_14938,N_14974);
nor UO_287 (O_287,N_14868,N_14867);
and UO_288 (O_288,N_14997,N_14943);
or UO_289 (O_289,N_14913,N_14949);
nand UO_290 (O_290,N_14910,N_14982);
and UO_291 (O_291,N_14923,N_14977);
or UO_292 (O_292,N_14956,N_14940);
xnor UO_293 (O_293,N_14873,N_14966);
nand UO_294 (O_294,N_14963,N_14986);
xor UO_295 (O_295,N_14893,N_14956);
nor UO_296 (O_296,N_14850,N_14925);
or UO_297 (O_297,N_14866,N_14932);
and UO_298 (O_298,N_14918,N_14915);
nand UO_299 (O_299,N_14851,N_14901);
nand UO_300 (O_300,N_14875,N_14905);
nor UO_301 (O_301,N_14957,N_14925);
nand UO_302 (O_302,N_14880,N_14960);
and UO_303 (O_303,N_14940,N_14883);
and UO_304 (O_304,N_14895,N_14908);
and UO_305 (O_305,N_14914,N_14924);
nor UO_306 (O_306,N_14982,N_14873);
or UO_307 (O_307,N_14908,N_14944);
or UO_308 (O_308,N_14991,N_14879);
nor UO_309 (O_309,N_14878,N_14948);
xnor UO_310 (O_310,N_14943,N_14854);
or UO_311 (O_311,N_14886,N_14995);
or UO_312 (O_312,N_14912,N_14924);
xnor UO_313 (O_313,N_14967,N_14905);
nor UO_314 (O_314,N_14983,N_14886);
nand UO_315 (O_315,N_14933,N_14996);
or UO_316 (O_316,N_14888,N_14997);
and UO_317 (O_317,N_14972,N_14898);
nand UO_318 (O_318,N_14860,N_14879);
nor UO_319 (O_319,N_14888,N_14901);
nand UO_320 (O_320,N_14931,N_14919);
nor UO_321 (O_321,N_14914,N_14968);
nand UO_322 (O_322,N_14890,N_14967);
or UO_323 (O_323,N_14912,N_14931);
and UO_324 (O_324,N_14860,N_14985);
nand UO_325 (O_325,N_14999,N_14958);
and UO_326 (O_326,N_14938,N_14959);
nand UO_327 (O_327,N_14868,N_14967);
or UO_328 (O_328,N_14892,N_14978);
nor UO_329 (O_329,N_14945,N_14991);
or UO_330 (O_330,N_14904,N_14988);
nor UO_331 (O_331,N_14938,N_14888);
nand UO_332 (O_332,N_14870,N_14896);
or UO_333 (O_333,N_14988,N_14941);
or UO_334 (O_334,N_14853,N_14983);
and UO_335 (O_335,N_14957,N_14934);
or UO_336 (O_336,N_14949,N_14911);
and UO_337 (O_337,N_14886,N_14858);
xor UO_338 (O_338,N_14993,N_14988);
nand UO_339 (O_339,N_14859,N_14927);
or UO_340 (O_340,N_14922,N_14965);
or UO_341 (O_341,N_14916,N_14947);
xnor UO_342 (O_342,N_14892,N_14994);
nand UO_343 (O_343,N_14912,N_14975);
and UO_344 (O_344,N_14902,N_14899);
nand UO_345 (O_345,N_14972,N_14874);
or UO_346 (O_346,N_14882,N_14985);
and UO_347 (O_347,N_14893,N_14915);
nor UO_348 (O_348,N_14935,N_14859);
nand UO_349 (O_349,N_14967,N_14960);
nor UO_350 (O_350,N_14932,N_14961);
nand UO_351 (O_351,N_14979,N_14887);
and UO_352 (O_352,N_14935,N_14946);
and UO_353 (O_353,N_14957,N_14905);
and UO_354 (O_354,N_14912,N_14922);
nand UO_355 (O_355,N_14855,N_14963);
or UO_356 (O_356,N_14984,N_14857);
and UO_357 (O_357,N_14945,N_14889);
and UO_358 (O_358,N_14879,N_14967);
nand UO_359 (O_359,N_14903,N_14966);
and UO_360 (O_360,N_14919,N_14991);
and UO_361 (O_361,N_14890,N_14986);
or UO_362 (O_362,N_14907,N_14905);
xor UO_363 (O_363,N_14887,N_14924);
or UO_364 (O_364,N_14937,N_14985);
nand UO_365 (O_365,N_14893,N_14910);
xnor UO_366 (O_366,N_14936,N_14991);
nand UO_367 (O_367,N_14906,N_14853);
or UO_368 (O_368,N_14874,N_14927);
nor UO_369 (O_369,N_14858,N_14891);
nand UO_370 (O_370,N_14908,N_14938);
or UO_371 (O_371,N_14940,N_14855);
and UO_372 (O_372,N_14876,N_14961);
and UO_373 (O_373,N_14997,N_14872);
or UO_374 (O_374,N_14853,N_14996);
or UO_375 (O_375,N_14914,N_14932);
nor UO_376 (O_376,N_14967,N_14907);
nand UO_377 (O_377,N_14915,N_14939);
or UO_378 (O_378,N_14994,N_14933);
and UO_379 (O_379,N_14889,N_14881);
nor UO_380 (O_380,N_14927,N_14853);
or UO_381 (O_381,N_14962,N_14915);
nand UO_382 (O_382,N_14988,N_14888);
xor UO_383 (O_383,N_14894,N_14978);
and UO_384 (O_384,N_14965,N_14962);
or UO_385 (O_385,N_14944,N_14886);
or UO_386 (O_386,N_14898,N_14889);
and UO_387 (O_387,N_14986,N_14974);
or UO_388 (O_388,N_14997,N_14908);
nor UO_389 (O_389,N_14969,N_14892);
or UO_390 (O_390,N_14877,N_14981);
or UO_391 (O_391,N_14876,N_14871);
or UO_392 (O_392,N_14874,N_14933);
nor UO_393 (O_393,N_14917,N_14933);
xnor UO_394 (O_394,N_14850,N_14937);
nand UO_395 (O_395,N_14970,N_14920);
nor UO_396 (O_396,N_14964,N_14893);
or UO_397 (O_397,N_14989,N_14995);
and UO_398 (O_398,N_14959,N_14933);
or UO_399 (O_399,N_14950,N_14932);
nor UO_400 (O_400,N_14937,N_14933);
nand UO_401 (O_401,N_14946,N_14979);
or UO_402 (O_402,N_14924,N_14991);
and UO_403 (O_403,N_14893,N_14967);
nor UO_404 (O_404,N_14969,N_14995);
or UO_405 (O_405,N_14921,N_14949);
nand UO_406 (O_406,N_14851,N_14875);
nor UO_407 (O_407,N_14870,N_14862);
or UO_408 (O_408,N_14889,N_14959);
nor UO_409 (O_409,N_14947,N_14896);
nor UO_410 (O_410,N_14969,N_14964);
or UO_411 (O_411,N_14993,N_14926);
nor UO_412 (O_412,N_14907,N_14948);
and UO_413 (O_413,N_14955,N_14895);
and UO_414 (O_414,N_14853,N_14951);
or UO_415 (O_415,N_14997,N_14940);
or UO_416 (O_416,N_14921,N_14930);
or UO_417 (O_417,N_14958,N_14856);
and UO_418 (O_418,N_14992,N_14881);
nor UO_419 (O_419,N_14924,N_14958);
and UO_420 (O_420,N_14898,N_14967);
or UO_421 (O_421,N_14868,N_14951);
nand UO_422 (O_422,N_14949,N_14891);
and UO_423 (O_423,N_14857,N_14876);
nand UO_424 (O_424,N_14944,N_14979);
or UO_425 (O_425,N_14853,N_14880);
nand UO_426 (O_426,N_14869,N_14998);
and UO_427 (O_427,N_14888,N_14900);
or UO_428 (O_428,N_14971,N_14982);
or UO_429 (O_429,N_14909,N_14989);
nand UO_430 (O_430,N_14960,N_14996);
and UO_431 (O_431,N_14985,N_14934);
and UO_432 (O_432,N_14886,N_14927);
nand UO_433 (O_433,N_14925,N_14912);
nor UO_434 (O_434,N_14973,N_14956);
nand UO_435 (O_435,N_14902,N_14956);
and UO_436 (O_436,N_14989,N_14879);
nand UO_437 (O_437,N_14880,N_14867);
nand UO_438 (O_438,N_14935,N_14909);
xor UO_439 (O_439,N_14877,N_14970);
nor UO_440 (O_440,N_14856,N_14880);
and UO_441 (O_441,N_14922,N_14850);
nand UO_442 (O_442,N_14869,N_14936);
and UO_443 (O_443,N_14913,N_14943);
nor UO_444 (O_444,N_14957,N_14959);
and UO_445 (O_445,N_14906,N_14915);
or UO_446 (O_446,N_14989,N_14897);
xor UO_447 (O_447,N_14962,N_14863);
nand UO_448 (O_448,N_14930,N_14881);
or UO_449 (O_449,N_14981,N_14851);
and UO_450 (O_450,N_14971,N_14890);
nand UO_451 (O_451,N_14882,N_14919);
and UO_452 (O_452,N_14943,N_14970);
or UO_453 (O_453,N_14957,N_14975);
nand UO_454 (O_454,N_14850,N_14890);
nand UO_455 (O_455,N_14909,N_14911);
nand UO_456 (O_456,N_14950,N_14941);
nor UO_457 (O_457,N_14926,N_14948);
nor UO_458 (O_458,N_14909,N_14991);
nor UO_459 (O_459,N_14905,N_14985);
or UO_460 (O_460,N_14942,N_14897);
or UO_461 (O_461,N_14934,N_14927);
and UO_462 (O_462,N_14886,N_14948);
nor UO_463 (O_463,N_14997,N_14972);
nand UO_464 (O_464,N_14852,N_14864);
nand UO_465 (O_465,N_14912,N_14883);
or UO_466 (O_466,N_14937,N_14965);
and UO_467 (O_467,N_14891,N_14920);
and UO_468 (O_468,N_14957,N_14891);
nor UO_469 (O_469,N_14917,N_14869);
and UO_470 (O_470,N_14871,N_14966);
nor UO_471 (O_471,N_14902,N_14995);
nor UO_472 (O_472,N_14903,N_14917);
and UO_473 (O_473,N_14871,N_14948);
or UO_474 (O_474,N_14960,N_14874);
and UO_475 (O_475,N_14863,N_14946);
nand UO_476 (O_476,N_14925,N_14996);
nor UO_477 (O_477,N_14966,N_14959);
and UO_478 (O_478,N_14951,N_14989);
nor UO_479 (O_479,N_14911,N_14902);
and UO_480 (O_480,N_14926,N_14860);
and UO_481 (O_481,N_14943,N_14894);
or UO_482 (O_482,N_14875,N_14966);
and UO_483 (O_483,N_14905,N_14984);
and UO_484 (O_484,N_14955,N_14945);
or UO_485 (O_485,N_14901,N_14968);
nand UO_486 (O_486,N_14870,N_14945);
nand UO_487 (O_487,N_14931,N_14973);
nand UO_488 (O_488,N_14858,N_14971);
and UO_489 (O_489,N_14962,N_14861);
and UO_490 (O_490,N_14966,N_14904);
xor UO_491 (O_491,N_14892,N_14869);
and UO_492 (O_492,N_14895,N_14880);
or UO_493 (O_493,N_14915,N_14942);
and UO_494 (O_494,N_14908,N_14973);
and UO_495 (O_495,N_14989,N_14997);
nand UO_496 (O_496,N_14881,N_14897);
nand UO_497 (O_497,N_14869,N_14851);
nor UO_498 (O_498,N_14856,N_14937);
or UO_499 (O_499,N_14887,N_14891);
nor UO_500 (O_500,N_14878,N_14940);
or UO_501 (O_501,N_14861,N_14899);
and UO_502 (O_502,N_14909,N_14925);
or UO_503 (O_503,N_14968,N_14904);
and UO_504 (O_504,N_14948,N_14859);
xor UO_505 (O_505,N_14970,N_14936);
nor UO_506 (O_506,N_14899,N_14896);
nand UO_507 (O_507,N_14921,N_14966);
nor UO_508 (O_508,N_14878,N_14990);
and UO_509 (O_509,N_14950,N_14893);
and UO_510 (O_510,N_14868,N_14870);
and UO_511 (O_511,N_14870,N_14908);
nor UO_512 (O_512,N_14945,N_14993);
nand UO_513 (O_513,N_14851,N_14908);
nor UO_514 (O_514,N_14976,N_14856);
or UO_515 (O_515,N_14866,N_14963);
nor UO_516 (O_516,N_14929,N_14983);
nor UO_517 (O_517,N_14993,N_14946);
nor UO_518 (O_518,N_14882,N_14886);
nor UO_519 (O_519,N_14920,N_14854);
or UO_520 (O_520,N_14968,N_14958);
nand UO_521 (O_521,N_14972,N_14926);
nand UO_522 (O_522,N_14977,N_14919);
nor UO_523 (O_523,N_14975,N_14879);
or UO_524 (O_524,N_14918,N_14883);
nor UO_525 (O_525,N_14927,N_14899);
and UO_526 (O_526,N_14892,N_14906);
and UO_527 (O_527,N_14854,N_14965);
or UO_528 (O_528,N_14864,N_14901);
or UO_529 (O_529,N_14894,N_14875);
and UO_530 (O_530,N_14876,N_14981);
and UO_531 (O_531,N_14995,N_14896);
nand UO_532 (O_532,N_14981,N_14867);
and UO_533 (O_533,N_14992,N_14850);
nand UO_534 (O_534,N_14872,N_14964);
nand UO_535 (O_535,N_14883,N_14986);
nor UO_536 (O_536,N_14879,N_14861);
or UO_537 (O_537,N_14862,N_14946);
nand UO_538 (O_538,N_14877,N_14882);
nor UO_539 (O_539,N_14915,N_14979);
nand UO_540 (O_540,N_14898,N_14968);
nor UO_541 (O_541,N_14902,N_14977);
nand UO_542 (O_542,N_14996,N_14954);
and UO_543 (O_543,N_14856,N_14961);
and UO_544 (O_544,N_14987,N_14893);
nor UO_545 (O_545,N_14951,N_14914);
xor UO_546 (O_546,N_14975,N_14973);
nand UO_547 (O_547,N_14980,N_14973);
or UO_548 (O_548,N_14919,N_14900);
and UO_549 (O_549,N_14962,N_14933);
or UO_550 (O_550,N_14858,N_14893);
or UO_551 (O_551,N_14889,N_14866);
xor UO_552 (O_552,N_14947,N_14883);
and UO_553 (O_553,N_14959,N_14998);
nor UO_554 (O_554,N_14898,N_14892);
or UO_555 (O_555,N_14928,N_14981);
nand UO_556 (O_556,N_14939,N_14975);
and UO_557 (O_557,N_14865,N_14949);
or UO_558 (O_558,N_14852,N_14924);
or UO_559 (O_559,N_14904,N_14905);
or UO_560 (O_560,N_14927,N_14880);
nand UO_561 (O_561,N_14930,N_14861);
nor UO_562 (O_562,N_14894,N_14916);
xor UO_563 (O_563,N_14987,N_14863);
nor UO_564 (O_564,N_14857,N_14931);
nor UO_565 (O_565,N_14863,N_14974);
nor UO_566 (O_566,N_14948,N_14999);
nor UO_567 (O_567,N_14968,N_14926);
and UO_568 (O_568,N_14863,N_14937);
or UO_569 (O_569,N_14998,N_14927);
or UO_570 (O_570,N_14904,N_14962);
and UO_571 (O_571,N_14897,N_14966);
nor UO_572 (O_572,N_14999,N_14861);
nor UO_573 (O_573,N_14921,N_14863);
nor UO_574 (O_574,N_14981,N_14947);
or UO_575 (O_575,N_14887,N_14989);
and UO_576 (O_576,N_14992,N_14914);
nor UO_577 (O_577,N_14949,N_14879);
nor UO_578 (O_578,N_14970,N_14933);
or UO_579 (O_579,N_14885,N_14853);
nor UO_580 (O_580,N_14919,N_14916);
nor UO_581 (O_581,N_14858,N_14967);
nor UO_582 (O_582,N_14997,N_14966);
or UO_583 (O_583,N_14881,N_14971);
nand UO_584 (O_584,N_14932,N_14934);
and UO_585 (O_585,N_14999,N_14963);
nand UO_586 (O_586,N_14889,N_14904);
nand UO_587 (O_587,N_14993,N_14955);
and UO_588 (O_588,N_14850,N_14990);
nor UO_589 (O_589,N_14978,N_14982);
xnor UO_590 (O_590,N_14954,N_14871);
and UO_591 (O_591,N_14960,N_14890);
or UO_592 (O_592,N_14963,N_14906);
xnor UO_593 (O_593,N_14917,N_14954);
and UO_594 (O_594,N_14993,N_14867);
xnor UO_595 (O_595,N_14920,N_14937);
nand UO_596 (O_596,N_14922,N_14854);
or UO_597 (O_597,N_14931,N_14874);
nand UO_598 (O_598,N_14970,N_14982);
and UO_599 (O_599,N_14994,N_14950);
nor UO_600 (O_600,N_14964,N_14879);
or UO_601 (O_601,N_14979,N_14964);
nand UO_602 (O_602,N_14974,N_14935);
xnor UO_603 (O_603,N_14935,N_14854);
or UO_604 (O_604,N_14901,N_14890);
nand UO_605 (O_605,N_14884,N_14859);
and UO_606 (O_606,N_14923,N_14958);
nand UO_607 (O_607,N_14993,N_14924);
nand UO_608 (O_608,N_14965,N_14982);
or UO_609 (O_609,N_14943,N_14944);
xor UO_610 (O_610,N_14890,N_14978);
or UO_611 (O_611,N_14908,N_14854);
xnor UO_612 (O_612,N_14899,N_14874);
nor UO_613 (O_613,N_14871,N_14925);
nand UO_614 (O_614,N_14905,N_14891);
nand UO_615 (O_615,N_14967,N_14927);
or UO_616 (O_616,N_14866,N_14938);
nor UO_617 (O_617,N_14955,N_14858);
and UO_618 (O_618,N_14952,N_14976);
nand UO_619 (O_619,N_14954,N_14870);
nor UO_620 (O_620,N_14994,N_14902);
or UO_621 (O_621,N_14992,N_14898);
or UO_622 (O_622,N_14959,N_14905);
or UO_623 (O_623,N_14933,N_14902);
nor UO_624 (O_624,N_14891,N_14959);
and UO_625 (O_625,N_14875,N_14886);
nor UO_626 (O_626,N_14877,N_14957);
or UO_627 (O_627,N_14954,N_14867);
nand UO_628 (O_628,N_14877,N_14965);
nand UO_629 (O_629,N_14961,N_14861);
nor UO_630 (O_630,N_14948,N_14977);
and UO_631 (O_631,N_14995,N_14949);
and UO_632 (O_632,N_14917,N_14885);
and UO_633 (O_633,N_14926,N_14852);
nor UO_634 (O_634,N_14875,N_14867);
xor UO_635 (O_635,N_14935,N_14892);
and UO_636 (O_636,N_14980,N_14870);
nand UO_637 (O_637,N_14899,N_14900);
and UO_638 (O_638,N_14942,N_14945);
and UO_639 (O_639,N_14909,N_14855);
nand UO_640 (O_640,N_14908,N_14855);
nand UO_641 (O_641,N_14981,N_14880);
and UO_642 (O_642,N_14874,N_14882);
nand UO_643 (O_643,N_14890,N_14930);
or UO_644 (O_644,N_14940,N_14907);
or UO_645 (O_645,N_14948,N_14998);
nand UO_646 (O_646,N_14928,N_14953);
nor UO_647 (O_647,N_14860,N_14852);
and UO_648 (O_648,N_14862,N_14951);
xnor UO_649 (O_649,N_14932,N_14978);
nand UO_650 (O_650,N_14918,N_14872);
nor UO_651 (O_651,N_14874,N_14958);
and UO_652 (O_652,N_14866,N_14919);
nand UO_653 (O_653,N_14954,N_14912);
or UO_654 (O_654,N_14901,N_14885);
and UO_655 (O_655,N_14958,N_14997);
nand UO_656 (O_656,N_14859,N_14894);
or UO_657 (O_657,N_14871,N_14979);
nor UO_658 (O_658,N_14913,N_14889);
nand UO_659 (O_659,N_14968,N_14918);
nand UO_660 (O_660,N_14917,N_14969);
and UO_661 (O_661,N_14900,N_14853);
nor UO_662 (O_662,N_14980,N_14907);
or UO_663 (O_663,N_14982,N_14913);
or UO_664 (O_664,N_14864,N_14886);
or UO_665 (O_665,N_14888,N_14998);
or UO_666 (O_666,N_14942,N_14999);
or UO_667 (O_667,N_14948,N_14904);
nand UO_668 (O_668,N_14990,N_14903);
and UO_669 (O_669,N_14920,N_14914);
or UO_670 (O_670,N_14955,N_14959);
nand UO_671 (O_671,N_14933,N_14978);
and UO_672 (O_672,N_14949,N_14970);
xor UO_673 (O_673,N_14974,N_14963);
nand UO_674 (O_674,N_14901,N_14954);
and UO_675 (O_675,N_14859,N_14887);
or UO_676 (O_676,N_14989,N_14953);
nor UO_677 (O_677,N_14947,N_14956);
nand UO_678 (O_678,N_14984,N_14871);
xor UO_679 (O_679,N_14985,N_14893);
or UO_680 (O_680,N_14897,N_14885);
xnor UO_681 (O_681,N_14959,N_14942);
and UO_682 (O_682,N_14997,N_14921);
or UO_683 (O_683,N_14880,N_14890);
and UO_684 (O_684,N_14988,N_14902);
nor UO_685 (O_685,N_14961,N_14966);
xor UO_686 (O_686,N_14861,N_14985);
and UO_687 (O_687,N_14885,N_14864);
nor UO_688 (O_688,N_14879,N_14899);
or UO_689 (O_689,N_14886,N_14910);
nand UO_690 (O_690,N_14967,N_14959);
nand UO_691 (O_691,N_14879,N_14960);
nand UO_692 (O_692,N_14917,N_14937);
nand UO_693 (O_693,N_14866,N_14914);
or UO_694 (O_694,N_14873,N_14874);
or UO_695 (O_695,N_14940,N_14980);
nand UO_696 (O_696,N_14929,N_14908);
or UO_697 (O_697,N_14916,N_14978);
xor UO_698 (O_698,N_14903,N_14863);
nand UO_699 (O_699,N_14922,N_14851);
or UO_700 (O_700,N_14923,N_14942);
and UO_701 (O_701,N_14855,N_14984);
or UO_702 (O_702,N_14945,N_14863);
nand UO_703 (O_703,N_14887,N_14912);
nand UO_704 (O_704,N_14889,N_14990);
nand UO_705 (O_705,N_14921,N_14999);
nor UO_706 (O_706,N_14973,N_14963);
nor UO_707 (O_707,N_14966,N_14910);
nor UO_708 (O_708,N_14926,N_14920);
nor UO_709 (O_709,N_14856,N_14866);
or UO_710 (O_710,N_14864,N_14883);
nand UO_711 (O_711,N_14927,N_14909);
and UO_712 (O_712,N_14987,N_14990);
nor UO_713 (O_713,N_14934,N_14993);
nand UO_714 (O_714,N_14882,N_14989);
nor UO_715 (O_715,N_14960,N_14974);
or UO_716 (O_716,N_14920,N_14954);
or UO_717 (O_717,N_14883,N_14919);
or UO_718 (O_718,N_14913,N_14855);
xnor UO_719 (O_719,N_14902,N_14851);
nor UO_720 (O_720,N_14879,N_14880);
nand UO_721 (O_721,N_14898,N_14939);
nor UO_722 (O_722,N_14983,N_14988);
and UO_723 (O_723,N_14936,N_14920);
or UO_724 (O_724,N_14912,N_14904);
and UO_725 (O_725,N_14928,N_14949);
or UO_726 (O_726,N_14920,N_14933);
and UO_727 (O_727,N_14996,N_14945);
nor UO_728 (O_728,N_14995,N_14895);
nor UO_729 (O_729,N_14947,N_14871);
and UO_730 (O_730,N_14929,N_14879);
or UO_731 (O_731,N_14889,N_14909);
or UO_732 (O_732,N_14892,N_14887);
nor UO_733 (O_733,N_14853,N_14955);
nand UO_734 (O_734,N_14894,N_14944);
nor UO_735 (O_735,N_14986,N_14909);
or UO_736 (O_736,N_14983,N_14885);
or UO_737 (O_737,N_14923,N_14995);
and UO_738 (O_738,N_14992,N_14853);
nor UO_739 (O_739,N_14904,N_14959);
and UO_740 (O_740,N_14958,N_14995);
xor UO_741 (O_741,N_14920,N_14948);
nand UO_742 (O_742,N_14867,N_14974);
and UO_743 (O_743,N_14947,N_14879);
nor UO_744 (O_744,N_14954,N_14907);
or UO_745 (O_745,N_14964,N_14963);
or UO_746 (O_746,N_14887,N_14860);
xor UO_747 (O_747,N_14902,N_14975);
and UO_748 (O_748,N_14938,N_14953);
nand UO_749 (O_749,N_14884,N_14883);
nor UO_750 (O_750,N_14957,N_14950);
or UO_751 (O_751,N_14960,N_14997);
nor UO_752 (O_752,N_14866,N_14927);
and UO_753 (O_753,N_14917,N_14892);
nor UO_754 (O_754,N_14993,N_14915);
nand UO_755 (O_755,N_14887,N_14983);
or UO_756 (O_756,N_14964,N_14921);
nor UO_757 (O_757,N_14943,N_14917);
and UO_758 (O_758,N_14921,N_14936);
nor UO_759 (O_759,N_14975,N_14930);
nor UO_760 (O_760,N_14923,N_14992);
nand UO_761 (O_761,N_14963,N_14948);
xor UO_762 (O_762,N_14898,N_14978);
or UO_763 (O_763,N_14881,N_14980);
nand UO_764 (O_764,N_14870,N_14976);
and UO_765 (O_765,N_14984,N_14851);
or UO_766 (O_766,N_14940,N_14919);
or UO_767 (O_767,N_14988,N_14932);
nor UO_768 (O_768,N_14914,N_14856);
or UO_769 (O_769,N_14960,N_14961);
nand UO_770 (O_770,N_14869,N_14972);
and UO_771 (O_771,N_14926,N_14882);
or UO_772 (O_772,N_14982,N_14963);
or UO_773 (O_773,N_14886,N_14876);
nor UO_774 (O_774,N_14898,N_14900);
and UO_775 (O_775,N_14893,N_14901);
and UO_776 (O_776,N_14869,N_14888);
nand UO_777 (O_777,N_14962,N_14916);
nor UO_778 (O_778,N_14862,N_14937);
xor UO_779 (O_779,N_14869,N_14909);
nor UO_780 (O_780,N_14852,N_14982);
or UO_781 (O_781,N_14935,N_14969);
or UO_782 (O_782,N_14936,N_14918);
nand UO_783 (O_783,N_14944,N_14973);
xor UO_784 (O_784,N_14926,N_14976);
or UO_785 (O_785,N_14990,N_14917);
or UO_786 (O_786,N_14951,N_14946);
nor UO_787 (O_787,N_14911,N_14924);
and UO_788 (O_788,N_14974,N_14900);
nor UO_789 (O_789,N_14878,N_14979);
or UO_790 (O_790,N_14919,N_14917);
xnor UO_791 (O_791,N_14935,N_14875);
nand UO_792 (O_792,N_14990,N_14961);
xnor UO_793 (O_793,N_14873,N_14913);
or UO_794 (O_794,N_14998,N_14910);
nand UO_795 (O_795,N_14887,N_14873);
or UO_796 (O_796,N_14943,N_14957);
and UO_797 (O_797,N_14859,N_14922);
and UO_798 (O_798,N_14850,N_14929);
and UO_799 (O_799,N_14914,N_14939);
and UO_800 (O_800,N_14950,N_14851);
nand UO_801 (O_801,N_14858,N_14964);
nand UO_802 (O_802,N_14977,N_14910);
or UO_803 (O_803,N_14865,N_14972);
nand UO_804 (O_804,N_14918,N_14854);
or UO_805 (O_805,N_14989,N_14933);
nor UO_806 (O_806,N_14929,N_14990);
nand UO_807 (O_807,N_14973,N_14885);
nor UO_808 (O_808,N_14968,N_14944);
xnor UO_809 (O_809,N_14932,N_14917);
or UO_810 (O_810,N_14877,N_14928);
and UO_811 (O_811,N_14902,N_14852);
nor UO_812 (O_812,N_14933,N_14888);
and UO_813 (O_813,N_14982,N_14920);
nand UO_814 (O_814,N_14887,N_14874);
nand UO_815 (O_815,N_14883,N_14949);
and UO_816 (O_816,N_14926,N_14957);
and UO_817 (O_817,N_14871,N_14919);
nand UO_818 (O_818,N_14966,N_14982);
and UO_819 (O_819,N_14982,N_14974);
nand UO_820 (O_820,N_14955,N_14893);
and UO_821 (O_821,N_14904,N_14939);
nor UO_822 (O_822,N_14891,N_14854);
xnor UO_823 (O_823,N_14858,N_14906);
nor UO_824 (O_824,N_14970,N_14926);
and UO_825 (O_825,N_14878,N_14875);
and UO_826 (O_826,N_14985,N_14998);
or UO_827 (O_827,N_14964,N_14952);
and UO_828 (O_828,N_14991,N_14927);
or UO_829 (O_829,N_14877,N_14952);
or UO_830 (O_830,N_14998,N_14930);
and UO_831 (O_831,N_14986,N_14983);
nand UO_832 (O_832,N_14922,N_14872);
or UO_833 (O_833,N_14859,N_14983);
nand UO_834 (O_834,N_14973,N_14946);
nor UO_835 (O_835,N_14867,N_14893);
or UO_836 (O_836,N_14951,N_14902);
or UO_837 (O_837,N_14930,N_14872);
nand UO_838 (O_838,N_14992,N_14908);
nor UO_839 (O_839,N_14942,N_14924);
and UO_840 (O_840,N_14888,N_14894);
xor UO_841 (O_841,N_14964,N_14850);
and UO_842 (O_842,N_14989,N_14968);
and UO_843 (O_843,N_14882,N_14864);
and UO_844 (O_844,N_14892,N_14857);
or UO_845 (O_845,N_14896,N_14872);
xor UO_846 (O_846,N_14946,N_14914);
or UO_847 (O_847,N_14987,N_14854);
xor UO_848 (O_848,N_14892,N_14907);
nor UO_849 (O_849,N_14937,N_14970);
and UO_850 (O_850,N_14850,N_14895);
or UO_851 (O_851,N_14988,N_14898);
or UO_852 (O_852,N_14931,N_14855);
nor UO_853 (O_853,N_14906,N_14854);
and UO_854 (O_854,N_14971,N_14952);
or UO_855 (O_855,N_14890,N_14918);
nor UO_856 (O_856,N_14864,N_14909);
nor UO_857 (O_857,N_14955,N_14901);
nor UO_858 (O_858,N_14931,N_14864);
nor UO_859 (O_859,N_14912,N_14929);
and UO_860 (O_860,N_14917,N_14866);
nand UO_861 (O_861,N_14937,N_14955);
and UO_862 (O_862,N_14956,N_14877);
or UO_863 (O_863,N_14996,N_14975);
and UO_864 (O_864,N_14914,N_14978);
and UO_865 (O_865,N_14912,N_14867);
nor UO_866 (O_866,N_14942,N_14938);
nor UO_867 (O_867,N_14938,N_14853);
or UO_868 (O_868,N_14991,N_14897);
or UO_869 (O_869,N_14987,N_14853);
nor UO_870 (O_870,N_14931,N_14939);
nand UO_871 (O_871,N_14914,N_14960);
and UO_872 (O_872,N_14907,N_14921);
nor UO_873 (O_873,N_14974,N_14920);
nor UO_874 (O_874,N_14955,N_14914);
nand UO_875 (O_875,N_14947,N_14997);
or UO_876 (O_876,N_14884,N_14994);
nor UO_877 (O_877,N_14996,N_14929);
xor UO_878 (O_878,N_14851,N_14926);
and UO_879 (O_879,N_14961,N_14871);
or UO_880 (O_880,N_14924,N_14907);
and UO_881 (O_881,N_14908,N_14977);
or UO_882 (O_882,N_14858,N_14953);
nand UO_883 (O_883,N_14934,N_14929);
nor UO_884 (O_884,N_14886,N_14891);
or UO_885 (O_885,N_14997,N_14877);
nand UO_886 (O_886,N_14895,N_14941);
or UO_887 (O_887,N_14919,N_14983);
xnor UO_888 (O_888,N_14954,N_14860);
nand UO_889 (O_889,N_14877,N_14986);
and UO_890 (O_890,N_14867,N_14904);
or UO_891 (O_891,N_14996,N_14974);
and UO_892 (O_892,N_14880,N_14866);
and UO_893 (O_893,N_14865,N_14964);
and UO_894 (O_894,N_14886,N_14917);
and UO_895 (O_895,N_14911,N_14947);
and UO_896 (O_896,N_14930,N_14853);
nor UO_897 (O_897,N_14890,N_14910);
xor UO_898 (O_898,N_14897,N_14992);
and UO_899 (O_899,N_14941,N_14916);
xor UO_900 (O_900,N_14983,N_14858);
or UO_901 (O_901,N_14851,N_14986);
nand UO_902 (O_902,N_14880,N_14978);
nor UO_903 (O_903,N_14939,N_14857);
nand UO_904 (O_904,N_14877,N_14857);
nor UO_905 (O_905,N_14907,N_14893);
or UO_906 (O_906,N_14913,N_14964);
nor UO_907 (O_907,N_14859,N_14987);
and UO_908 (O_908,N_14926,N_14916);
or UO_909 (O_909,N_14957,N_14910);
or UO_910 (O_910,N_14948,N_14942);
nand UO_911 (O_911,N_14956,N_14883);
nand UO_912 (O_912,N_14981,N_14936);
nor UO_913 (O_913,N_14968,N_14999);
nor UO_914 (O_914,N_14963,N_14939);
nor UO_915 (O_915,N_14925,N_14863);
xor UO_916 (O_916,N_14850,N_14919);
or UO_917 (O_917,N_14855,N_14879);
or UO_918 (O_918,N_14932,N_14879);
and UO_919 (O_919,N_14913,N_14884);
or UO_920 (O_920,N_14896,N_14990);
nand UO_921 (O_921,N_14910,N_14917);
nor UO_922 (O_922,N_14880,N_14992);
or UO_923 (O_923,N_14977,N_14953);
nand UO_924 (O_924,N_14950,N_14852);
nor UO_925 (O_925,N_14927,N_14936);
nor UO_926 (O_926,N_14879,N_14873);
xor UO_927 (O_927,N_14934,N_14859);
and UO_928 (O_928,N_14889,N_14863);
nor UO_929 (O_929,N_14908,N_14850);
and UO_930 (O_930,N_14921,N_14879);
nor UO_931 (O_931,N_14936,N_14952);
nand UO_932 (O_932,N_14920,N_14938);
nand UO_933 (O_933,N_14970,N_14918);
and UO_934 (O_934,N_14894,N_14919);
xnor UO_935 (O_935,N_14884,N_14929);
nor UO_936 (O_936,N_14876,N_14946);
xnor UO_937 (O_937,N_14896,N_14853);
nand UO_938 (O_938,N_14947,N_14862);
nand UO_939 (O_939,N_14956,N_14988);
or UO_940 (O_940,N_14949,N_14931);
or UO_941 (O_941,N_14933,N_14885);
and UO_942 (O_942,N_14990,N_14870);
and UO_943 (O_943,N_14997,N_14876);
nor UO_944 (O_944,N_14931,N_14892);
or UO_945 (O_945,N_14998,N_14873);
nor UO_946 (O_946,N_14868,N_14955);
and UO_947 (O_947,N_14936,N_14915);
and UO_948 (O_948,N_14915,N_14995);
nor UO_949 (O_949,N_14974,N_14921);
or UO_950 (O_950,N_14985,N_14981);
nor UO_951 (O_951,N_14864,N_14972);
or UO_952 (O_952,N_14938,N_14930);
nor UO_953 (O_953,N_14995,N_14976);
and UO_954 (O_954,N_14902,N_14878);
nor UO_955 (O_955,N_14982,N_14958);
and UO_956 (O_956,N_14882,N_14855);
or UO_957 (O_957,N_14965,N_14973);
nand UO_958 (O_958,N_14953,N_14969);
nor UO_959 (O_959,N_14929,N_14977);
or UO_960 (O_960,N_14952,N_14859);
nor UO_961 (O_961,N_14896,N_14925);
nand UO_962 (O_962,N_14944,N_14936);
or UO_963 (O_963,N_14865,N_14994);
xor UO_964 (O_964,N_14981,N_14952);
xnor UO_965 (O_965,N_14913,N_14944);
and UO_966 (O_966,N_14949,N_14899);
nand UO_967 (O_967,N_14883,N_14908);
nand UO_968 (O_968,N_14967,N_14990);
xnor UO_969 (O_969,N_14928,N_14998);
or UO_970 (O_970,N_14872,N_14990);
or UO_971 (O_971,N_14875,N_14960);
nand UO_972 (O_972,N_14894,N_14970);
xnor UO_973 (O_973,N_14893,N_14895);
and UO_974 (O_974,N_14853,N_14907);
nand UO_975 (O_975,N_14878,N_14929);
nor UO_976 (O_976,N_14875,N_14996);
and UO_977 (O_977,N_14905,N_14866);
nand UO_978 (O_978,N_14951,N_14880);
and UO_979 (O_979,N_14970,N_14997);
and UO_980 (O_980,N_14918,N_14895);
nand UO_981 (O_981,N_14892,N_14988);
and UO_982 (O_982,N_14994,N_14999);
nor UO_983 (O_983,N_14852,N_14904);
and UO_984 (O_984,N_14971,N_14954);
nand UO_985 (O_985,N_14891,N_14955);
and UO_986 (O_986,N_14957,N_14945);
nand UO_987 (O_987,N_14911,N_14879);
nor UO_988 (O_988,N_14878,N_14874);
and UO_989 (O_989,N_14876,N_14935);
xor UO_990 (O_990,N_14890,N_14866);
and UO_991 (O_991,N_14933,N_14856);
nor UO_992 (O_992,N_14880,N_14876);
and UO_993 (O_993,N_14944,N_14872);
or UO_994 (O_994,N_14970,N_14884);
nor UO_995 (O_995,N_14905,N_14943);
nor UO_996 (O_996,N_14988,N_14916);
nor UO_997 (O_997,N_14947,N_14899);
or UO_998 (O_998,N_14904,N_14882);
and UO_999 (O_999,N_14873,N_14960);
or UO_1000 (O_1000,N_14923,N_14991);
nand UO_1001 (O_1001,N_14871,N_14962);
nor UO_1002 (O_1002,N_14902,N_14889);
nand UO_1003 (O_1003,N_14912,N_14859);
nor UO_1004 (O_1004,N_14866,N_14996);
or UO_1005 (O_1005,N_14877,N_14863);
nand UO_1006 (O_1006,N_14888,N_14962);
and UO_1007 (O_1007,N_14987,N_14918);
nor UO_1008 (O_1008,N_14924,N_14920);
nand UO_1009 (O_1009,N_14986,N_14998);
nor UO_1010 (O_1010,N_14932,N_14936);
and UO_1011 (O_1011,N_14886,N_14872);
and UO_1012 (O_1012,N_14883,N_14889);
nand UO_1013 (O_1013,N_14912,N_14882);
and UO_1014 (O_1014,N_14925,N_14880);
or UO_1015 (O_1015,N_14920,N_14873);
and UO_1016 (O_1016,N_14868,N_14855);
nor UO_1017 (O_1017,N_14930,N_14884);
and UO_1018 (O_1018,N_14876,N_14873);
and UO_1019 (O_1019,N_14986,N_14921);
xnor UO_1020 (O_1020,N_14930,N_14863);
nor UO_1021 (O_1021,N_14921,N_14991);
nor UO_1022 (O_1022,N_14909,N_14993);
xnor UO_1023 (O_1023,N_14868,N_14872);
xnor UO_1024 (O_1024,N_14921,N_14855);
nand UO_1025 (O_1025,N_14901,N_14982);
nand UO_1026 (O_1026,N_14931,N_14928);
nand UO_1027 (O_1027,N_14895,N_14855);
and UO_1028 (O_1028,N_14993,N_14900);
nand UO_1029 (O_1029,N_14852,N_14975);
nand UO_1030 (O_1030,N_14865,N_14968);
xnor UO_1031 (O_1031,N_14860,N_14948);
nand UO_1032 (O_1032,N_14984,N_14958);
nand UO_1033 (O_1033,N_14932,N_14975);
and UO_1034 (O_1034,N_14932,N_14955);
and UO_1035 (O_1035,N_14938,N_14964);
nand UO_1036 (O_1036,N_14928,N_14957);
nand UO_1037 (O_1037,N_14924,N_14889);
or UO_1038 (O_1038,N_14906,N_14987);
and UO_1039 (O_1039,N_14874,N_14928);
nand UO_1040 (O_1040,N_14923,N_14990);
and UO_1041 (O_1041,N_14933,N_14867);
xor UO_1042 (O_1042,N_14920,N_14987);
and UO_1043 (O_1043,N_14899,N_14872);
nand UO_1044 (O_1044,N_14907,N_14861);
and UO_1045 (O_1045,N_14916,N_14851);
and UO_1046 (O_1046,N_14967,N_14903);
or UO_1047 (O_1047,N_14982,N_14872);
nand UO_1048 (O_1048,N_14858,N_14880);
or UO_1049 (O_1049,N_14887,N_14890);
or UO_1050 (O_1050,N_14903,N_14937);
or UO_1051 (O_1051,N_14942,N_14868);
and UO_1052 (O_1052,N_14904,N_14975);
or UO_1053 (O_1053,N_14961,N_14975);
nor UO_1054 (O_1054,N_14907,N_14887);
and UO_1055 (O_1055,N_14912,N_14952);
nor UO_1056 (O_1056,N_14853,N_14905);
nor UO_1057 (O_1057,N_14869,N_14949);
and UO_1058 (O_1058,N_14935,N_14920);
or UO_1059 (O_1059,N_14963,N_14977);
or UO_1060 (O_1060,N_14968,N_14933);
nand UO_1061 (O_1061,N_14862,N_14897);
and UO_1062 (O_1062,N_14997,N_14992);
or UO_1063 (O_1063,N_14891,N_14999);
and UO_1064 (O_1064,N_14993,N_14930);
nor UO_1065 (O_1065,N_14988,N_14877);
xnor UO_1066 (O_1066,N_14858,N_14999);
nor UO_1067 (O_1067,N_14952,N_14906);
or UO_1068 (O_1068,N_14917,N_14912);
or UO_1069 (O_1069,N_14965,N_14915);
nor UO_1070 (O_1070,N_14913,N_14955);
nor UO_1071 (O_1071,N_14850,N_14943);
or UO_1072 (O_1072,N_14863,N_14990);
nand UO_1073 (O_1073,N_14954,N_14861);
and UO_1074 (O_1074,N_14913,N_14934);
xor UO_1075 (O_1075,N_14866,N_14896);
nand UO_1076 (O_1076,N_14929,N_14904);
nand UO_1077 (O_1077,N_14974,N_14882);
and UO_1078 (O_1078,N_14982,N_14977);
nand UO_1079 (O_1079,N_14900,N_14901);
or UO_1080 (O_1080,N_14996,N_14884);
nor UO_1081 (O_1081,N_14979,N_14914);
nand UO_1082 (O_1082,N_14892,N_14876);
and UO_1083 (O_1083,N_14941,N_14924);
nand UO_1084 (O_1084,N_14865,N_14874);
nand UO_1085 (O_1085,N_14905,N_14999);
nor UO_1086 (O_1086,N_14939,N_14987);
nand UO_1087 (O_1087,N_14907,N_14883);
and UO_1088 (O_1088,N_14867,N_14864);
or UO_1089 (O_1089,N_14888,N_14931);
and UO_1090 (O_1090,N_14918,N_14982);
nand UO_1091 (O_1091,N_14891,N_14873);
nand UO_1092 (O_1092,N_14922,N_14925);
and UO_1093 (O_1093,N_14947,N_14912);
or UO_1094 (O_1094,N_14983,N_14962);
or UO_1095 (O_1095,N_14988,N_14975);
or UO_1096 (O_1096,N_14896,N_14996);
nand UO_1097 (O_1097,N_14938,N_14994);
and UO_1098 (O_1098,N_14873,N_14938);
nand UO_1099 (O_1099,N_14882,N_14899);
nand UO_1100 (O_1100,N_14872,N_14960);
xnor UO_1101 (O_1101,N_14924,N_14864);
nand UO_1102 (O_1102,N_14857,N_14888);
xor UO_1103 (O_1103,N_14998,N_14937);
nor UO_1104 (O_1104,N_14949,N_14920);
nor UO_1105 (O_1105,N_14931,N_14967);
or UO_1106 (O_1106,N_14874,N_14904);
nor UO_1107 (O_1107,N_14981,N_14993);
or UO_1108 (O_1108,N_14865,N_14915);
nand UO_1109 (O_1109,N_14914,N_14956);
nor UO_1110 (O_1110,N_14851,N_14858);
xnor UO_1111 (O_1111,N_14982,N_14904);
and UO_1112 (O_1112,N_14928,N_14873);
and UO_1113 (O_1113,N_14956,N_14938);
nand UO_1114 (O_1114,N_14911,N_14872);
and UO_1115 (O_1115,N_14867,N_14962);
and UO_1116 (O_1116,N_14994,N_14970);
xor UO_1117 (O_1117,N_14852,N_14877);
nor UO_1118 (O_1118,N_14887,N_14987);
and UO_1119 (O_1119,N_14888,N_14957);
xor UO_1120 (O_1120,N_14924,N_14850);
nor UO_1121 (O_1121,N_14984,N_14944);
nand UO_1122 (O_1122,N_14935,N_14908);
xor UO_1123 (O_1123,N_14938,N_14931);
or UO_1124 (O_1124,N_14925,N_14948);
nand UO_1125 (O_1125,N_14984,N_14856);
or UO_1126 (O_1126,N_14894,N_14990);
or UO_1127 (O_1127,N_14906,N_14925);
nand UO_1128 (O_1128,N_14880,N_14924);
nand UO_1129 (O_1129,N_14895,N_14875);
or UO_1130 (O_1130,N_14855,N_14979);
nand UO_1131 (O_1131,N_14924,N_14978);
or UO_1132 (O_1132,N_14919,N_14973);
nand UO_1133 (O_1133,N_14929,N_14875);
nor UO_1134 (O_1134,N_14919,N_14952);
nand UO_1135 (O_1135,N_14981,N_14863);
xnor UO_1136 (O_1136,N_14874,N_14922);
and UO_1137 (O_1137,N_14911,N_14938);
and UO_1138 (O_1138,N_14861,N_14876);
or UO_1139 (O_1139,N_14854,N_14899);
and UO_1140 (O_1140,N_14863,N_14942);
and UO_1141 (O_1141,N_14978,N_14948);
nand UO_1142 (O_1142,N_14941,N_14901);
and UO_1143 (O_1143,N_14877,N_14881);
nor UO_1144 (O_1144,N_14906,N_14895);
and UO_1145 (O_1145,N_14917,N_14904);
or UO_1146 (O_1146,N_14887,N_14990);
xor UO_1147 (O_1147,N_14887,N_14997);
or UO_1148 (O_1148,N_14996,N_14898);
nand UO_1149 (O_1149,N_14935,N_14915);
nand UO_1150 (O_1150,N_14945,N_14857);
nand UO_1151 (O_1151,N_14940,N_14979);
nand UO_1152 (O_1152,N_14945,N_14892);
nor UO_1153 (O_1153,N_14952,N_14934);
and UO_1154 (O_1154,N_14988,N_14963);
nand UO_1155 (O_1155,N_14911,N_14887);
xnor UO_1156 (O_1156,N_14971,N_14991);
nor UO_1157 (O_1157,N_14885,N_14980);
and UO_1158 (O_1158,N_14944,N_14867);
or UO_1159 (O_1159,N_14913,N_14891);
or UO_1160 (O_1160,N_14928,N_14992);
or UO_1161 (O_1161,N_14894,N_14902);
nand UO_1162 (O_1162,N_14901,N_14991);
and UO_1163 (O_1163,N_14982,N_14862);
and UO_1164 (O_1164,N_14927,N_14988);
and UO_1165 (O_1165,N_14964,N_14978);
or UO_1166 (O_1166,N_14930,N_14914);
and UO_1167 (O_1167,N_14879,N_14913);
nor UO_1168 (O_1168,N_14976,N_14884);
and UO_1169 (O_1169,N_14975,N_14920);
nand UO_1170 (O_1170,N_14854,N_14927);
xor UO_1171 (O_1171,N_14961,N_14905);
xor UO_1172 (O_1172,N_14894,N_14873);
nor UO_1173 (O_1173,N_14906,N_14953);
nor UO_1174 (O_1174,N_14954,N_14977);
and UO_1175 (O_1175,N_14901,N_14952);
nand UO_1176 (O_1176,N_14864,N_14880);
nand UO_1177 (O_1177,N_14986,N_14996);
or UO_1178 (O_1178,N_14879,N_14968);
and UO_1179 (O_1179,N_14868,N_14873);
and UO_1180 (O_1180,N_14936,N_14922);
or UO_1181 (O_1181,N_14920,N_14969);
xnor UO_1182 (O_1182,N_14894,N_14887);
nand UO_1183 (O_1183,N_14914,N_14958);
or UO_1184 (O_1184,N_14881,N_14973);
or UO_1185 (O_1185,N_14925,N_14930);
nor UO_1186 (O_1186,N_14880,N_14934);
nor UO_1187 (O_1187,N_14962,N_14990);
or UO_1188 (O_1188,N_14862,N_14975);
and UO_1189 (O_1189,N_14882,N_14858);
and UO_1190 (O_1190,N_14869,N_14970);
or UO_1191 (O_1191,N_14942,N_14851);
nand UO_1192 (O_1192,N_14851,N_14879);
nor UO_1193 (O_1193,N_14909,N_14901);
xor UO_1194 (O_1194,N_14879,N_14850);
xnor UO_1195 (O_1195,N_14932,N_14963);
or UO_1196 (O_1196,N_14892,N_14851);
or UO_1197 (O_1197,N_14996,N_14957);
nand UO_1198 (O_1198,N_14935,N_14896);
or UO_1199 (O_1199,N_14956,N_14941);
or UO_1200 (O_1200,N_14980,N_14916);
nor UO_1201 (O_1201,N_14982,N_14994);
or UO_1202 (O_1202,N_14859,N_14895);
xnor UO_1203 (O_1203,N_14967,N_14892);
nand UO_1204 (O_1204,N_14908,N_14999);
nor UO_1205 (O_1205,N_14916,N_14861);
nand UO_1206 (O_1206,N_14885,N_14899);
and UO_1207 (O_1207,N_14855,N_14973);
nor UO_1208 (O_1208,N_14877,N_14914);
nor UO_1209 (O_1209,N_14955,N_14920);
nand UO_1210 (O_1210,N_14890,N_14951);
and UO_1211 (O_1211,N_14996,N_14999);
nand UO_1212 (O_1212,N_14870,N_14905);
nor UO_1213 (O_1213,N_14859,N_14861);
nand UO_1214 (O_1214,N_14864,N_14905);
or UO_1215 (O_1215,N_14969,N_14945);
nor UO_1216 (O_1216,N_14955,N_14855);
and UO_1217 (O_1217,N_14954,N_14923);
and UO_1218 (O_1218,N_14995,N_14883);
or UO_1219 (O_1219,N_14931,N_14876);
nand UO_1220 (O_1220,N_14954,N_14962);
nor UO_1221 (O_1221,N_14911,N_14925);
xor UO_1222 (O_1222,N_14979,N_14869);
xor UO_1223 (O_1223,N_14963,N_14934);
nand UO_1224 (O_1224,N_14983,N_14976);
and UO_1225 (O_1225,N_14879,N_14999);
or UO_1226 (O_1226,N_14896,N_14955);
nand UO_1227 (O_1227,N_14856,N_14951);
nand UO_1228 (O_1228,N_14933,N_14990);
and UO_1229 (O_1229,N_14870,N_14926);
and UO_1230 (O_1230,N_14915,N_14908);
nand UO_1231 (O_1231,N_14948,N_14921);
nor UO_1232 (O_1232,N_14987,N_14969);
or UO_1233 (O_1233,N_14928,N_14967);
nor UO_1234 (O_1234,N_14869,N_14878);
nor UO_1235 (O_1235,N_14853,N_14862);
nand UO_1236 (O_1236,N_14969,N_14983);
or UO_1237 (O_1237,N_14887,N_14938);
and UO_1238 (O_1238,N_14983,N_14905);
or UO_1239 (O_1239,N_14912,N_14903);
and UO_1240 (O_1240,N_14944,N_14948);
nand UO_1241 (O_1241,N_14954,N_14976);
nor UO_1242 (O_1242,N_14900,N_14889);
and UO_1243 (O_1243,N_14883,N_14869);
nand UO_1244 (O_1244,N_14987,N_14970);
and UO_1245 (O_1245,N_14919,N_14942);
nand UO_1246 (O_1246,N_14886,N_14912);
and UO_1247 (O_1247,N_14912,N_14868);
nor UO_1248 (O_1248,N_14908,N_14911);
and UO_1249 (O_1249,N_14924,N_14951);
and UO_1250 (O_1250,N_14993,N_14963);
nor UO_1251 (O_1251,N_14939,N_14900);
xor UO_1252 (O_1252,N_14921,N_14885);
nand UO_1253 (O_1253,N_14923,N_14913);
nand UO_1254 (O_1254,N_14923,N_14907);
and UO_1255 (O_1255,N_14991,N_14970);
or UO_1256 (O_1256,N_14993,N_14880);
and UO_1257 (O_1257,N_14900,N_14911);
and UO_1258 (O_1258,N_14873,N_14929);
nor UO_1259 (O_1259,N_14926,N_14989);
or UO_1260 (O_1260,N_14978,N_14919);
nand UO_1261 (O_1261,N_14887,N_14942);
and UO_1262 (O_1262,N_14949,N_14906);
nor UO_1263 (O_1263,N_14933,N_14859);
and UO_1264 (O_1264,N_14907,N_14877);
and UO_1265 (O_1265,N_14988,N_14976);
or UO_1266 (O_1266,N_14899,N_14983);
and UO_1267 (O_1267,N_14987,N_14953);
or UO_1268 (O_1268,N_14873,N_14940);
or UO_1269 (O_1269,N_14961,N_14950);
nor UO_1270 (O_1270,N_14936,N_14872);
nand UO_1271 (O_1271,N_14937,N_14876);
and UO_1272 (O_1272,N_14907,N_14933);
nor UO_1273 (O_1273,N_14976,N_14896);
nor UO_1274 (O_1274,N_14905,N_14975);
xor UO_1275 (O_1275,N_14877,N_14992);
nor UO_1276 (O_1276,N_14873,N_14907);
nor UO_1277 (O_1277,N_14878,N_14923);
or UO_1278 (O_1278,N_14876,N_14960);
xor UO_1279 (O_1279,N_14935,N_14941);
and UO_1280 (O_1280,N_14912,N_14992);
xor UO_1281 (O_1281,N_14889,N_14992);
and UO_1282 (O_1282,N_14892,N_14924);
xor UO_1283 (O_1283,N_14865,N_14935);
nand UO_1284 (O_1284,N_14946,N_14910);
or UO_1285 (O_1285,N_14882,N_14990);
nor UO_1286 (O_1286,N_14882,N_14944);
and UO_1287 (O_1287,N_14934,N_14866);
nor UO_1288 (O_1288,N_14880,N_14886);
and UO_1289 (O_1289,N_14867,N_14911);
or UO_1290 (O_1290,N_14912,N_14852);
or UO_1291 (O_1291,N_14906,N_14979);
nand UO_1292 (O_1292,N_14870,N_14963);
and UO_1293 (O_1293,N_14867,N_14957);
nand UO_1294 (O_1294,N_14868,N_14970);
nor UO_1295 (O_1295,N_14921,N_14861);
and UO_1296 (O_1296,N_14850,N_14979);
xor UO_1297 (O_1297,N_14952,N_14987);
nor UO_1298 (O_1298,N_14922,N_14956);
or UO_1299 (O_1299,N_14875,N_14988);
nand UO_1300 (O_1300,N_14963,N_14953);
and UO_1301 (O_1301,N_14968,N_14996);
nor UO_1302 (O_1302,N_14938,N_14936);
and UO_1303 (O_1303,N_14914,N_14898);
or UO_1304 (O_1304,N_14947,N_14975);
xnor UO_1305 (O_1305,N_14974,N_14926);
or UO_1306 (O_1306,N_14870,N_14982);
or UO_1307 (O_1307,N_14977,N_14998);
nand UO_1308 (O_1308,N_14938,N_14914);
xor UO_1309 (O_1309,N_14902,N_14958);
nand UO_1310 (O_1310,N_14894,N_14954);
xnor UO_1311 (O_1311,N_14980,N_14892);
nor UO_1312 (O_1312,N_14861,N_14936);
and UO_1313 (O_1313,N_14899,N_14857);
and UO_1314 (O_1314,N_14964,N_14983);
nor UO_1315 (O_1315,N_14898,N_14936);
nor UO_1316 (O_1316,N_14966,N_14924);
or UO_1317 (O_1317,N_14870,N_14890);
xor UO_1318 (O_1318,N_14877,N_14984);
nor UO_1319 (O_1319,N_14876,N_14983);
and UO_1320 (O_1320,N_14943,N_14955);
and UO_1321 (O_1321,N_14897,N_14882);
and UO_1322 (O_1322,N_14875,N_14869);
xor UO_1323 (O_1323,N_14851,N_14853);
nand UO_1324 (O_1324,N_14913,N_14937);
xnor UO_1325 (O_1325,N_14993,N_14976);
nor UO_1326 (O_1326,N_14881,N_14998);
or UO_1327 (O_1327,N_14991,N_14992);
and UO_1328 (O_1328,N_14961,N_14878);
and UO_1329 (O_1329,N_14868,N_14954);
nor UO_1330 (O_1330,N_14908,N_14878);
xnor UO_1331 (O_1331,N_14916,N_14939);
nor UO_1332 (O_1332,N_14850,N_14935);
nor UO_1333 (O_1333,N_14903,N_14904);
nor UO_1334 (O_1334,N_14935,N_14950);
and UO_1335 (O_1335,N_14978,N_14955);
or UO_1336 (O_1336,N_14915,N_14948);
nand UO_1337 (O_1337,N_14920,N_14905);
nor UO_1338 (O_1338,N_14876,N_14980);
nor UO_1339 (O_1339,N_14884,N_14952);
and UO_1340 (O_1340,N_14914,N_14999);
nand UO_1341 (O_1341,N_14998,N_14983);
nand UO_1342 (O_1342,N_14891,N_14943);
or UO_1343 (O_1343,N_14960,N_14962);
nor UO_1344 (O_1344,N_14955,N_14944);
or UO_1345 (O_1345,N_14908,N_14867);
nor UO_1346 (O_1346,N_14938,N_14966);
nor UO_1347 (O_1347,N_14936,N_14888);
xor UO_1348 (O_1348,N_14882,N_14898);
or UO_1349 (O_1349,N_14962,N_14899);
nor UO_1350 (O_1350,N_14947,N_14952);
nor UO_1351 (O_1351,N_14853,N_14899);
and UO_1352 (O_1352,N_14911,N_14855);
nand UO_1353 (O_1353,N_14854,N_14997);
and UO_1354 (O_1354,N_14903,N_14892);
and UO_1355 (O_1355,N_14960,N_14881);
and UO_1356 (O_1356,N_14901,N_14951);
and UO_1357 (O_1357,N_14900,N_14882);
or UO_1358 (O_1358,N_14956,N_14870);
nor UO_1359 (O_1359,N_14961,N_14973);
or UO_1360 (O_1360,N_14867,N_14869);
or UO_1361 (O_1361,N_14930,N_14911);
or UO_1362 (O_1362,N_14853,N_14924);
nor UO_1363 (O_1363,N_14903,N_14971);
nor UO_1364 (O_1364,N_14854,N_14962);
xor UO_1365 (O_1365,N_14867,N_14959);
or UO_1366 (O_1366,N_14972,N_14861);
and UO_1367 (O_1367,N_14860,N_14923);
and UO_1368 (O_1368,N_14966,N_14905);
nor UO_1369 (O_1369,N_14898,N_14943);
and UO_1370 (O_1370,N_14949,N_14856);
nor UO_1371 (O_1371,N_14875,N_14893);
nand UO_1372 (O_1372,N_14976,N_14876);
and UO_1373 (O_1373,N_14851,N_14854);
and UO_1374 (O_1374,N_14962,N_14924);
xnor UO_1375 (O_1375,N_14915,N_14988);
nor UO_1376 (O_1376,N_14928,N_14902);
and UO_1377 (O_1377,N_14873,N_14866);
nand UO_1378 (O_1378,N_14987,N_14864);
and UO_1379 (O_1379,N_14930,N_14970);
nor UO_1380 (O_1380,N_14994,N_14991);
and UO_1381 (O_1381,N_14866,N_14850);
nor UO_1382 (O_1382,N_14987,N_14986);
and UO_1383 (O_1383,N_14911,N_14852);
or UO_1384 (O_1384,N_14897,N_14949);
and UO_1385 (O_1385,N_14860,N_14924);
xnor UO_1386 (O_1386,N_14878,N_14989);
and UO_1387 (O_1387,N_14965,N_14929);
and UO_1388 (O_1388,N_14907,N_14968);
nand UO_1389 (O_1389,N_14879,N_14910);
nand UO_1390 (O_1390,N_14928,N_14979);
and UO_1391 (O_1391,N_14906,N_14930);
and UO_1392 (O_1392,N_14975,N_14944);
nand UO_1393 (O_1393,N_14866,N_14857);
xor UO_1394 (O_1394,N_14873,N_14896);
and UO_1395 (O_1395,N_14966,N_14950);
and UO_1396 (O_1396,N_14958,N_14895);
nor UO_1397 (O_1397,N_14978,N_14954);
xor UO_1398 (O_1398,N_14989,N_14871);
nor UO_1399 (O_1399,N_14904,N_14998);
nand UO_1400 (O_1400,N_14920,N_14963);
and UO_1401 (O_1401,N_14956,N_14971);
and UO_1402 (O_1402,N_14977,N_14866);
nor UO_1403 (O_1403,N_14871,N_14908);
or UO_1404 (O_1404,N_14952,N_14984);
or UO_1405 (O_1405,N_14993,N_14967);
nand UO_1406 (O_1406,N_14953,N_14918);
nor UO_1407 (O_1407,N_14881,N_14924);
nor UO_1408 (O_1408,N_14904,N_14886);
or UO_1409 (O_1409,N_14941,N_14938);
nor UO_1410 (O_1410,N_14938,N_14876);
nand UO_1411 (O_1411,N_14977,N_14872);
nand UO_1412 (O_1412,N_14866,N_14949);
nor UO_1413 (O_1413,N_14852,N_14862);
or UO_1414 (O_1414,N_14906,N_14878);
or UO_1415 (O_1415,N_14981,N_14973);
or UO_1416 (O_1416,N_14948,N_14867);
xnor UO_1417 (O_1417,N_14930,N_14981);
and UO_1418 (O_1418,N_14945,N_14915);
nand UO_1419 (O_1419,N_14901,N_14945);
nand UO_1420 (O_1420,N_14984,N_14870);
nand UO_1421 (O_1421,N_14878,N_14914);
or UO_1422 (O_1422,N_14898,N_14903);
nor UO_1423 (O_1423,N_14861,N_14947);
xor UO_1424 (O_1424,N_14858,N_14985);
xnor UO_1425 (O_1425,N_14880,N_14976);
xnor UO_1426 (O_1426,N_14911,N_14853);
nand UO_1427 (O_1427,N_14892,N_14954);
nor UO_1428 (O_1428,N_14970,N_14992);
xnor UO_1429 (O_1429,N_14942,N_14958);
nor UO_1430 (O_1430,N_14983,N_14922);
xor UO_1431 (O_1431,N_14875,N_14957);
nor UO_1432 (O_1432,N_14953,N_14980);
nor UO_1433 (O_1433,N_14931,N_14890);
nor UO_1434 (O_1434,N_14922,N_14972);
and UO_1435 (O_1435,N_14906,N_14888);
or UO_1436 (O_1436,N_14970,N_14909);
or UO_1437 (O_1437,N_14868,N_14956);
nor UO_1438 (O_1438,N_14884,N_14870);
and UO_1439 (O_1439,N_14949,N_14987);
nand UO_1440 (O_1440,N_14912,N_14981);
or UO_1441 (O_1441,N_14882,N_14941);
nand UO_1442 (O_1442,N_14961,N_14963);
nand UO_1443 (O_1443,N_14970,N_14863);
nand UO_1444 (O_1444,N_14955,N_14957);
and UO_1445 (O_1445,N_14938,N_14897);
nor UO_1446 (O_1446,N_14977,N_14979);
or UO_1447 (O_1447,N_14933,N_14953);
nor UO_1448 (O_1448,N_14867,N_14900);
nor UO_1449 (O_1449,N_14948,N_14951);
and UO_1450 (O_1450,N_14874,N_14901);
nand UO_1451 (O_1451,N_14948,N_14893);
or UO_1452 (O_1452,N_14925,N_14956);
nand UO_1453 (O_1453,N_14928,N_14959);
and UO_1454 (O_1454,N_14943,N_14969);
and UO_1455 (O_1455,N_14906,N_14900);
and UO_1456 (O_1456,N_14900,N_14994);
and UO_1457 (O_1457,N_14894,N_14855);
or UO_1458 (O_1458,N_14985,N_14948);
and UO_1459 (O_1459,N_14901,N_14976);
nor UO_1460 (O_1460,N_14979,N_14971);
and UO_1461 (O_1461,N_14987,N_14937);
and UO_1462 (O_1462,N_14998,N_14892);
and UO_1463 (O_1463,N_14964,N_14884);
nor UO_1464 (O_1464,N_14922,N_14898);
nor UO_1465 (O_1465,N_14911,N_14976);
nor UO_1466 (O_1466,N_14939,N_14885);
nand UO_1467 (O_1467,N_14927,N_14989);
nand UO_1468 (O_1468,N_14880,N_14901);
nor UO_1469 (O_1469,N_14908,N_14897);
xnor UO_1470 (O_1470,N_14887,N_14966);
nor UO_1471 (O_1471,N_14988,N_14910);
xor UO_1472 (O_1472,N_14940,N_14866);
nand UO_1473 (O_1473,N_14908,N_14906);
and UO_1474 (O_1474,N_14908,N_14863);
xnor UO_1475 (O_1475,N_14883,N_14880);
nor UO_1476 (O_1476,N_14856,N_14967);
nand UO_1477 (O_1477,N_14892,N_14908);
and UO_1478 (O_1478,N_14911,N_14873);
and UO_1479 (O_1479,N_14966,N_14896);
nand UO_1480 (O_1480,N_14913,N_14876);
nand UO_1481 (O_1481,N_14860,N_14909);
or UO_1482 (O_1482,N_14980,N_14948);
or UO_1483 (O_1483,N_14875,N_14857);
and UO_1484 (O_1484,N_14913,N_14995);
nand UO_1485 (O_1485,N_14884,N_14945);
nor UO_1486 (O_1486,N_14890,N_14873);
and UO_1487 (O_1487,N_14972,N_14876);
xor UO_1488 (O_1488,N_14855,N_14970);
or UO_1489 (O_1489,N_14888,N_14961);
nand UO_1490 (O_1490,N_14894,N_14939);
and UO_1491 (O_1491,N_14989,N_14861);
nor UO_1492 (O_1492,N_14892,N_14993);
or UO_1493 (O_1493,N_14881,N_14884);
nor UO_1494 (O_1494,N_14914,N_14977);
nand UO_1495 (O_1495,N_14969,N_14886);
and UO_1496 (O_1496,N_14894,N_14879);
nand UO_1497 (O_1497,N_14980,N_14942);
or UO_1498 (O_1498,N_14869,N_14855);
nand UO_1499 (O_1499,N_14886,N_14884);
nor UO_1500 (O_1500,N_14862,N_14878);
and UO_1501 (O_1501,N_14986,N_14902);
nand UO_1502 (O_1502,N_14998,N_14856);
nor UO_1503 (O_1503,N_14859,N_14972);
nor UO_1504 (O_1504,N_14885,N_14943);
or UO_1505 (O_1505,N_14981,N_14879);
and UO_1506 (O_1506,N_14967,N_14996);
and UO_1507 (O_1507,N_14850,N_14855);
nand UO_1508 (O_1508,N_14934,N_14975);
nor UO_1509 (O_1509,N_14963,N_14869);
or UO_1510 (O_1510,N_14852,N_14931);
or UO_1511 (O_1511,N_14870,N_14960);
and UO_1512 (O_1512,N_14965,N_14907);
nor UO_1513 (O_1513,N_14893,N_14908);
nor UO_1514 (O_1514,N_14988,N_14858);
xnor UO_1515 (O_1515,N_14987,N_14956);
nand UO_1516 (O_1516,N_14907,N_14876);
nor UO_1517 (O_1517,N_14859,N_14994);
or UO_1518 (O_1518,N_14862,N_14879);
or UO_1519 (O_1519,N_14937,N_14966);
or UO_1520 (O_1520,N_14996,N_14981);
and UO_1521 (O_1521,N_14869,N_14879);
or UO_1522 (O_1522,N_14910,N_14873);
or UO_1523 (O_1523,N_14869,N_14922);
nor UO_1524 (O_1524,N_14882,N_14887);
xnor UO_1525 (O_1525,N_14903,N_14910);
xor UO_1526 (O_1526,N_14871,N_14892);
nor UO_1527 (O_1527,N_14997,N_14965);
xnor UO_1528 (O_1528,N_14897,N_14909);
or UO_1529 (O_1529,N_14962,N_14943);
nor UO_1530 (O_1530,N_14978,N_14946);
nand UO_1531 (O_1531,N_14865,N_14898);
nor UO_1532 (O_1532,N_14936,N_14873);
nor UO_1533 (O_1533,N_14917,N_14941);
nand UO_1534 (O_1534,N_14894,N_14856);
or UO_1535 (O_1535,N_14895,N_14884);
and UO_1536 (O_1536,N_14936,N_14945);
nor UO_1537 (O_1537,N_14864,N_14897);
or UO_1538 (O_1538,N_14869,N_14889);
or UO_1539 (O_1539,N_14855,N_14953);
nand UO_1540 (O_1540,N_14850,N_14884);
and UO_1541 (O_1541,N_14905,N_14953);
nor UO_1542 (O_1542,N_14972,N_14928);
and UO_1543 (O_1543,N_14922,N_14966);
nor UO_1544 (O_1544,N_14962,N_14911);
or UO_1545 (O_1545,N_14899,N_14966);
or UO_1546 (O_1546,N_14899,N_14969);
nand UO_1547 (O_1547,N_14967,N_14942);
nor UO_1548 (O_1548,N_14917,N_14901);
nor UO_1549 (O_1549,N_14981,N_14883);
and UO_1550 (O_1550,N_14879,N_14866);
nand UO_1551 (O_1551,N_14916,N_14896);
nor UO_1552 (O_1552,N_14905,N_14936);
xnor UO_1553 (O_1553,N_14950,N_14992);
nor UO_1554 (O_1554,N_14928,N_14914);
or UO_1555 (O_1555,N_14960,N_14930);
xor UO_1556 (O_1556,N_14921,N_14891);
or UO_1557 (O_1557,N_14885,N_14862);
nor UO_1558 (O_1558,N_14980,N_14853);
nand UO_1559 (O_1559,N_14913,N_14887);
and UO_1560 (O_1560,N_14918,N_14905);
xnor UO_1561 (O_1561,N_14877,N_14949);
nand UO_1562 (O_1562,N_14934,N_14911);
and UO_1563 (O_1563,N_14856,N_14926);
or UO_1564 (O_1564,N_14898,N_14879);
and UO_1565 (O_1565,N_14982,N_14895);
or UO_1566 (O_1566,N_14954,N_14936);
or UO_1567 (O_1567,N_14991,N_14890);
xnor UO_1568 (O_1568,N_14989,N_14998);
or UO_1569 (O_1569,N_14855,N_14950);
or UO_1570 (O_1570,N_14862,N_14894);
nand UO_1571 (O_1571,N_14939,N_14877);
or UO_1572 (O_1572,N_14901,N_14942);
nor UO_1573 (O_1573,N_14895,N_14992);
and UO_1574 (O_1574,N_14994,N_14920);
or UO_1575 (O_1575,N_14963,N_14896);
nor UO_1576 (O_1576,N_14934,N_14942);
or UO_1577 (O_1577,N_14929,N_14942);
xor UO_1578 (O_1578,N_14882,N_14940);
or UO_1579 (O_1579,N_14935,N_14887);
nor UO_1580 (O_1580,N_14970,N_14886);
and UO_1581 (O_1581,N_14974,N_14977);
nand UO_1582 (O_1582,N_14989,N_14851);
or UO_1583 (O_1583,N_14878,N_14957);
nor UO_1584 (O_1584,N_14878,N_14996);
or UO_1585 (O_1585,N_14869,N_14950);
or UO_1586 (O_1586,N_14914,N_14896);
nor UO_1587 (O_1587,N_14897,N_14906);
nand UO_1588 (O_1588,N_14949,N_14975);
nor UO_1589 (O_1589,N_14975,N_14972);
or UO_1590 (O_1590,N_14921,N_14985);
or UO_1591 (O_1591,N_14884,N_14896);
nor UO_1592 (O_1592,N_14990,N_14921);
nand UO_1593 (O_1593,N_14907,N_14973);
and UO_1594 (O_1594,N_14989,N_14934);
and UO_1595 (O_1595,N_14866,N_14913);
and UO_1596 (O_1596,N_14891,N_14958);
nand UO_1597 (O_1597,N_14909,N_14881);
nand UO_1598 (O_1598,N_14991,N_14958);
or UO_1599 (O_1599,N_14903,N_14916);
and UO_1600 (O_1600,N_14881,N_14874);
and UO_1601 (O_1601,N_14886,N_14976);
nand UO_1602 (O_1602,N_14869,N_14931);
nand UO_1603 (O_1603,N_14992,N_14989);
nor UO_1604 (O_1604,N_14873,N_14851);
or UO_1605 (O_1605,N_14900,N_14875);
nand UO_1606 (O_1606,N_14885,N_14990);
and UO_1607 (O_1607,N_14876,N_14999);
nor UO_1608 (O_1608,N_14989,N_14940);
xor UO_1609 (O_1609,N_14950,N_14973);
or UO_1610 (O_1610,N_14922,N_14889);
nor UO_1611 (O_1611,N_14978,N_14956);
and UO_1612 (O_1612,N_14876,N_14902);
nor UO_1613 (O_1613,N_14917,N_14899);
nor UO_1614 (O_1614,N_14882,N_14909);
or UO_1615 (O_1615,N_14886,N_14907);
or UO_1616 (O_1616,N_14912,N_14945);
nand UO_1617 (O_1617,N_14988,N_14855);
and UO_1618 (O_1618,N_14879,N_14888);
nand UO_1619 (O_1619,N_14927,N_14879);
nor UO_1620 (O_1620,N_14859,N_14953);
nand UO_1621 (O_1621,N_14962,N_14981);
or UO_1622 (O_1622,N_14866,N_14935);
nand UO_1623 (O_1623,N_14949,N_14885);
and UO_1624 (O_1624,N_14967,N_14963);
or UO_1625 (O_1625,N_14953,N_14973);
or UO_1626 (O_1626,N_14967,N_14997);
nand UO_1627 (O_1627,N_14982,N_14987);
or UO_1628 (O_1628,N_14993,N_14996);
or UO_1629 (O_1629,N_14907,N_14851);
nand UO_1630 (O_1630,N_14876,N_14956);
or UO_1631 (O_1631,N_14901,N_14972);
xnor UO_1632 (O_1632,N_14931,N_14930);
or UO_1633 (O_1633,N_14914,N_14862);
or UO_1634 (O_1634,N_14966,N_14935);
nand UO_1635 (O_1635,N_14934,N_14940);
nor UO_1636 (O_1636,N_14882,N_14977);
nor UO_1637 (O_1637,N_14900,N_14998);
nand UO_1638 (O_1638,N_14939,N_14911);
or UO_1639 (O_1639,N_14869,N_14914);
xnor UO_1640 (O_1640,N_14865,N_14916);
nor UO_1641 (O_1641,N_14923,N_14852);
nor UO_1642 (O_1642,N_14896,N_14927);
nor UO_1643 (O_1643,N_14982,N_14928);
nor UO_1644 (O_1644,N_14872,N_14866);
and UO_1645 (O_1645,N_14994,N_14989);
and UO_1646 (O_1646,N_14864,N_14944);
and UO_1647 (O_1647,N_14864,N_14977);
xor UO_1648 (O_1648,N_14930,N_14949);
or UO_1649 (O_1649,N_14926,N_14862);
or UO_1650 (O_1650,N_14921,N_14955);
or UO_1651 (O_1651,N_14851,N_14924);
and UO_1652 (O_1652,N_14866,N_14962);
nand UO_1653 (O_1653,N_14851,N_14918);
nor UO_1654 (O_1654,N_14970,N_14983);
or UO_1655 (O_1655,N_14946,N_14857);
xnor UO_1656 (O_1656,N_14958,N_14971);
or UO_1657 (O_1657,N_14924,N_14895);
xnor UO_1658 (O_1658,N_14957,N_14906);
and UO_1659 (O_1659,N_14857,N_14996);
or UO_1660 (O_1660,N_14926,N_14956);
and UO_1661 (O_1661,N_14994,N_14861);
or UO_1662 (O_1662,N_14856,N_14863);
or UO_1663 (O_1663,N_14886,N_14937);
nor UO_1664 (O_1664,N_14869,N_14852);
or UO_1665 (O_1665,N_14887,N_14958);
nor UO_1666 (O_1666,N_14968,N_14920);
or UO_1667 (O_1667,N_14964,N_14982);
or UO_1668 (O_1668,N_14918,N_14884);
or UO_1669 (O_1669,N_14879,N_14985);
nand UO_1670 (O_1670,N_14863,N_14909);
and UO_1671 (O_1671,N_14976,N_14924);
nor UO_1672 (O_1672,N_14942,N_14983);
nor UO_1673 (O_1673,N_14881,N_14929);
or UO_1674 (O_1674,N_14945,N_14903);
nor UO_1675 (O_1675,N_14983,N_14984);
nand UO_1676 (O_1676,N_14960,N_14965);
or UO_1677 (O_1677,N_14962,N_14937);
or UO_1678 (O_1678,N_14929,N_14888);
or UO_1679 (O_1679,N_14891,N_14877);
and UO_1680 (O_1680,N_14923,N_14917);
and UO_1681 (O_1681,N_14896,N_14888);
xnor UO_1682 (O_1682,N_14971,N_14919);
nand UO_1683 (O_1683,N_14866,N_14947);
and UO_1684 (O_1684,N_14934,N_14967);
nor UO_1685 (O_1685,N_14965,N_14896);
xnor UO_1686 (O_1686,N_14969,N_14906);
and UO_1687 (O_1687,N_14973,N_14894);
and UO_1688 (O_1688,N_14938,N_14937);
or UO_1689 (O_1689,N_14980,N_14998);
and UO_1690 (O_1690,N_14947,N_14885);
nand UO_1691 (O_1691,N_14862,N_14996);
nand UO_1692 (O_1692,N_14879,N_14990);
nand UO_1693 (O_1693,N_14925,N_14953);
nand UO_1694 (O_1694,N_14971,N_14989);
nor UO_1695 (O_1695,N_14979,N_14967);
nor UO_1696 (O_1696,N_14965,N_14956);
or UO_1697 (O_1697,N_14907,N_14904);
and UO_1698 (O_1698,N_14986,N_14879);
and UO_1699 (O_1699,N_14985,N_14958);
and UO_1700 (O_1700,N_14963,N_14962);
or UO_1701 (O_1701,N_14891,N_14876);
or UO_1702 (O_1702,N_14978,N_14980);
and UO_1703 (O_1703,N_14940,N_14944);
nor UO_1704 (O_1704,N_14920,N_14985);
and UO_1705 (O_1705,N_14884,N_14890);
nand UO_1706 (O_1706,N_14999,N_14873);
nor UO_1707 (O_1707,N_14891,N_14872);
nand UO_1708 (O_1708,N_14998,N_14941);
nand UO_1709 (O_1709,N_14921,N_14993);
or UO_1710 (O_1710,N_14878,N_14917);
and UO_1711 (O_1711,N_14928,N_14929);
nor UO_1712 (O_1712,N_14963,N_14942);
and UO_1713 (O_1713,N_14929,N_14985);
nand UO_1714 (O_1714,N_14926,N_14949);
and UO_1715 (O_1715,N_14935,N_14864);
nand UO_1716 (O_1716,N_14892,N_14948);
nor UO_1717 (O_1717,N_14988,N_14918);
or UO_1718 (O_1718,N_14946,N_14868);
or UO_1719 (O_1719,N_14959,N_14963);
xnor UO_1720 (O_1720,N_14880,N_14857);
or UO_1721 (O_1721,N_14878,N_14858);
nor UO_1722 (O_1722,N_14856,N_14888);
or UO_1723 (O_1723,N_14966,N_14973);
and UO_1724 (O_1724,N_14931,N_14887);
or UO_1725 (O_1725,N_14885,N_14908);
or UO_1726 (O_1726,N_14854,N_14948);
xnor UO_1727 (O_1727,N_14948,N_14991);
nor UO_1728 (O_1728,N_14992,N_14879);
nand UO_1729 (O_1729,N_14884,N_14891);
or UO_1730 (O_1730,N_14886,N_14851);
nand UO_1731 (O_1731,N_14900,N_14918);
and UO_1732 (O_1732,N_14927,N_14855);
nand UO_1733 (O_1733,N_14890,N_14851);
nand UO_1734 (O_1734,N_14984,N_14872);
or UO_1735 (O_1735,N_14859,N_14924);
or UO_1736 (O_1736,N_14921,N_14945);
nand UO_1737 (O_1737,N_14891,N_14923);
nand UO_1738 (O_1738,N_14924,N_14876);
nor UO_1739 (O_1739,N_14922,N_14911);
nor UO_1740 (O_1740,N_14920,N_14925);
or UO_1741 (O_1741,N_14973,N_14913);
nor UO_1742 (O_1742,N_14996,N_14873);
nand UO_1743 (O_1743,N_14961,N_14944);
nor UO_1744 (O_1744,N_14863,N_14896);
or UO_1745 (O_1745,N_14962,N_14908);
nor UO_1746 (O_1746,N_14930,N_14862);
and UO_1747 (O_1747,N_14850,N_14995);
and UO_1748 (O_1748,N_14994,N_14952);
or UO_1749 (O_1749,N_14870,N_14860);
nand UO_1750 (O_1750,N_14985,N_14960);
xor UO_1751 (O_1751,N_14904,N_14883);
nor UO_1752 (O_1752,N_14859,N_14899);
nand UO_1753 (O_1753,N_14892,N_14990);
nand UO_1754 (O_1754,N_14913,N_14905);
and UO_1755 (O_1755,N_14909,N_14933);
nand UO_1756 (O_1756,N_14953,N_14936);
and UO_1757 (O_1757,N_14994,N_14969);
nor UO_1758 (O_1758,N_14990,N_14898);
nand UO_1759 (O_1759,N_14941,N_14959);
and UO_1760 (O_1760,N_14945,N_14898);
and UO_1761 (O_1761,N_14921,N_14871);
nor UO_1762 (O_1762,N_14871,N_14978);
nor UO_1763 (O_1763,N_14857,N_14989);
and UO_1764 (O_1764,N_14932,N_14949);
or UO_1765 (O_1765,N_14870,N_14930);
nor UO_1766 (O_1766,N_14877,N_14851);
nor UO_1767 (O_1767,N_14884,N_14910);
and UO_1768 (O_1768,N_14951,N_14983);
or UO_1769 (O_1769,N_14885,N_14946);
nand UO_1770 (O_1770,N_14964,N_14962);
and UO_1771 (O_1771,N_14933,N_14991);
or UO_1772 (O_1772,N_14871,N_14981);
nand UO_1773 (O_1773,N_14949,N_14853);
or UO_1774 (O_1774,N_14994,N_14997);
nand UO_1775 (O_1775,N_14857,N_14911);
xor UO_1776 (O_1776,N_14946,N_14941);
nand UO_1777 (O_1777,N_14932,N_14926);
nor UO_1778 (O_1778,N_14943,N_14983);
nand UO_1779 (O_1779,N_14879,N_14941);
and UO_1780 (O_1780,N_14921,N_14872);
nand UO_1781 (O_1781,N_14890,N_14888);
nand UO_1782 (O_1782,N_14859,N_14973);
nand UO_1783 (O_1783,N_14929,N_14986);
nor UO_1784 (O_1784,N_14991,N_14872);
nand UO_1785 (O_1785,N_14854,N_14999);
nand UO_1786 (O_1786,N_14895,N_14856);
xnor UO_1787 (O_1787,N_14871,N_14972);
xnor UO_1788 (O_1788,N_14947,N_14978);
nor UO_1789 (O_1789,N_14930,N_14875);
nand UO_1790 (O_1790,N_14963,N_14996);
or UO_1791 (O_1791,N_14913,N_14882);
and UO_1792 (O_1792,N_14991,N_14930);
xor UO_1793 (O_1793,N_14928,N_14909);
nor UO_1794 (O_1794,N_14951,N_14896);
or UO_1795 (O_1795,N_14993,N_14994);
nor UO_1796 (O_1796,N_14865,N_14861);
xnor UO_1797 (O_1797,N_14942,N_14890);
nor UO_1798 (O_1798,N_14984,N_14899);
nand UO_1799 (O_1799,N_14873,N_14884);
and UO_1800 (O_1800,N_14871,N_14982);
and UO_1801 (O_1801,N_14854,N_14870);
nand UO_1802 (O_1802,N_14877,N_14895);
or UO_1803 (O_1803,N_14890,N_14981);
or UO_1804 (O_1804,N_14988,N_14900);
and UO_1805 (O_1805,N_14886,N_14968);
xnor UO_1806 (O_1806,N_14974,N_14869);
or UO_1807 (O_1807,N_14877,N_14868);
and UO_1808 (O_1808,N_14905,N_14910);
nor UO_1809 (O_1809,N_14913,N_14910);
or UO_1810 (O_1810,N_14880,N_14852);
and UO_1811 (O_1811,N_14917,N_14864);
xnor UO_1812 (O_1812,N_14952,N_14959);
and UO_1813 (O_1813,N_14872,N_14893);
nand UO_1814 (O_1814,N_14951,N_14963);
nand UO_1815 (O_1815,N_14852,N_14976);
nor UO_1816 (O_1816,N_14981,N_14910);
nor UO_1817 (O_1817,N_14912,N_14909);
nor UO_1818 (O_1818,N_14969,N_14924);
nand UO_1819 (O_1819,N_14853,N_14861);
nand UO_1820 (O_1820,N_14891,N_14995);
xor UO_1821 (O_1821,N_14898,N_14854);
or UO_1822 (O_1822,N_14950,N_14857);
and UO_1823 (O_1823,N_14981,N_14866);
nand UO_1824 (O_1824,N_14909,N_14985);
or UO_1825 (O_1825,N_14969,N_14908);
nand UO_1826 (O_1826,N_14930,N_14868);
nor UO_1827 (O_1827,N_14988,N_14899);
nor UO_1828 (O_1828,N_14883,N_14961);
and UO_1829 (O_1829,N_14941,N_14942);
and UO_1830 (O_1830,N_14984,N_14961);
xor UO_1831 (O_1831,N_14977,N_14964);
nand UO_1832 (O_1832,N_14866,N_14871);
or UO_1833 (O_1833,N_14973,N_14958);
and UO_1834 (O_1834,N_14879,N_14982);
and UO_1835 (O_1835,N_14971,N_14874);
nand UO_1836 (O_1836,N_14959,N_14975);
or UO_1837 (O_1837,N_14926,N_14895);
and UO_1838 (O_1838,N_14881,N_14950);
or UO_1839 (O_1839,N_14982,N_14943);
nor UO_1840 (O_1840,N_14906,N_14850);
nand UO_1841 (O_1841,N_14910,N_14883);
and UO_1842 (O_1842,N_14941,N_14974);
or UO_1843 (O_1843,N_14936,N_14923);
and UO_1844 (O_1844,N_14933,N_14930);
and UO_1845 (O_1845,N_14978,N_14850);
and UO_1846 (O_1846,N_14924,N_14869);
nand UO_1847 (O_1847,N_14918,N_14958);
or UO_1848 (O_1848,N_14985,N_14980);
or UO_1849 (O_1849,N_14991,N_14911);
nand UO_1850 (O_1850,N_14897,N_14940);
nor UO_1851 (O_1851,N_14933,N_14914);
and UO_1852 (O_1852,N_14907,N_14961);
nor UO_1853 (O_1853,N_14861,N_14862);
or UO_1854 (O_1854,N_14860,N_14945);
nand UO_1855 (O_1855,N_14853,N_14909);
and UO_1856 (O_1856,N_14931,N_14945);
nor UO_1857 (O_1857,N_14914,N_14855);
xor UO_1858 (O_1858,N_14997,N_14891);
and UO_1859 (O_1859,N_14915,N_14854);
or UO_1860 (O_1860,N_14931,N_14985);
or UO_1861 (O_1861,N_14953,N_14956);
or UO_1862 (O_1862,N_14920,N_14862);
nor UO_1863 (O_1863,N_14941,N_14857);
or UO_1864 (O_1864,N_14879,N_14961);
nor UO_1865 (O_1865,N_14955,N_14876);
nor UO_1866 (O_1866,N_14929,N_14980);
and UO_1867 (O_1867,N_14966,N_14946);
nand UO_1868 (O_1868,N_14993,N_14908);
nor UO_1869 (O_1869,N_14969,N_14970);
nor UO_1870 (O_1870,N_14900,N_14979);
or UO_1871 (O_1871,N_14903,N_14981);
nor UO_1872 (O_1872,N_14933,N_14866);
and UO_1873 (O_1873,N_14950,N_14926);
nand UO_1874 (O_1874,N_14961,N_14926);
or UO_1875 (O_1875,N_14855,N_14901);
nor UO_1876 (O_1876,N_14878,N_14885);
nor UO_1877 (O_1877,N_14972,N_14971);
xnor UO_1878 (O_1878,N_14933,N_14887);
nor UO_1879 (O_1879,N_14976,N_14929);
nand UO_1880 (O_1880,N_14885,N_14935);
or UO_1881 (O_1881,N_14870,N_14983);
and UO_1882 (O_1882,N_14874,N_14967);
nor UO_1883 (O_1883,N_14868,N_14878);
nand UO_1884 (O_1884,N_14906,N_14922);
or UO_1885 (O_1885,N_14859,N_14879);
and UO_1886 (O_1886,N_14885,N_14883);
or UO_1887 (O_1887,N_14880,N_14916);
and UO_1888 (O_1888,N_14865,N_14892);
or UO_1889 (O_1889,N_14945,N_14893);
nand UO_1890 (O_1890,N_14909,N_14919);
xor UO_1891 (O_1891,N_14963,N_14860);
or UO_1892 (O_1892,N_14950,N_14975);
xor UO_1893 (O_1893,N_14878,N_14980);
nor UO_1894 (O_1894,N_14923,N_14964);
nor UO_1895 (O_1895,N_14971,N_14902);
nand UO_1896 (O_1896,N_14866,N_14874);
nor UO_1897 (O_1897,N_14948,N_14889);
or UO_1898 (O_1898,N_14969,N_14893);
xnor UO_1899 (O_1899,N_14977,N_14945);
and UO_1900 (O_1900,N_14943,N_14993);
nand UO_1901 (O_1901,N_14916,N_14888);
nand UO_1902 (O_1902,N_14895,N_14913);
or UO_1903 (O_1903,N_14994,N_14882);
and UO_1904 (O_1904,N_14942,N_14882);
nand UO_1905 (O_1905,N_14894,N_14918);
xnor UO_1906 (O_1906,N_14873,N_14921);
or UO_1907 (O_1907,N_14918,N_14889);
nor UO_1908 (O_1908,N_14858,N_14942);
or UO_1909 (O_1909,N_14978,N_14908);
nand UO_1910 (O_1910,N_14882,N_14988);
nor UO_1911 (O_1911,N_14986,N_14907);
and UO_1912 (O_1912,N_14962,N_14882);
or UO_1913 (O_1913,N_14939,N_14977);
xnor UO_1914 (O_1914,N_14944,N_14998);
or UO_1915 (O_1915,N_14893,N_14903);
xnor UO_1916 (O_1916,N_14861,N_14909);
nand UO_1917 (O_1917,N_14946,N_14850);
nor UO_1918 (O_1918,N_14910,N_14994);
or UO_1919 (O_1919,N_14968,N_14994);
or UO_1920 (O_1920,N_14923,N_14981);
nand UO_1921 (O_1921,N_14877,N_14861);
or UO_1922 (O_1922,N_14919,N_14939);
nand UO_1923 (O_1923,N_14954,N_14890);
and UO_1924 (O_1924,N_14885,N_14940);
or UO_1925 (O_1925,N_14984,N_14879);
or UO_1926 (O_1926,N_14998,N_14911);
or UO_1927 (O_1927,N_14954,N_14979);
nand UO_1928 (O_1928,N_14891,N_14941);
nor UO_1929 (O_1929,N_14922,N_14862);
nand UO_1930 (O_1930,N_14941,N_14963);
and UO_1931 (O_1931,N_14984,N_14907);
nor UO_1932 (O_1932,N_14932,N_14909);
or UO_1933 (O_1933,N_14954,N_14914);
nor UO_1934 (O_1934,N_14941,N_14947);
nor UO_1935 (O_1935,N_14872,N_14998);
nand UO_1936 (O_1936,N_14948,N_14946);
or UO_1937 (O_1937,N_14994,N_14894);
nand UO_1938 (O_1938,N_14996,N_14992);
xor UO_1939 (O_1939,N_14956,N_14910);
or UO_1940 (O_1940,N_14965,N_14874);
xor UO_1941 (O_1941,N_14962,N_14971);
nor UO_1942 (O_1942,N_14976,N_14996);
nand UO_1943 (O_1943,N_14954,N_14989);
or UO_1944 (O_1944,N_14947,N_14915);
nor UO_1945 (O_1945,N_14966,N_14865);
nand UO_1946 (O_1946,N_14885,N_14911);
nand UO_1947 (O_1947,N_14927,N_14891);
and UO_1948 (O_1948,N_14909,N_14957);
nand UO_1949 (O_1949,N_14922,N_14873);
and UO_1950 (O_1950,N_14860,N_14988);
and UO_1951 (O_1951,N_14989,N_14853);
nand UO_1952 (O_1952,N_14917,N_14942);
or UO_1953 (O_1953,N_14969,N_14859);
or UO_1954 (O_1954,N_14959,N_14940);
or UO_1955 (O_1955,N_14963,N_14865);
and UO_1956 (O_1956,N_14874,N_14943);
nand UO_1957 (O_1957,N_14978,N_14857);
nand UO_1958 (O_1958,N_14900,N_14960);
nand UO_1959 (O_1959,N_14880,N_14973);
and UO_1960 (O_1960,N_14980,N_14858);
nor UO_1961 (O_1961,N_14934,N_14883);
xor UO_1962 (O_1962,N_14943,N_14961);
xor UO_1963 (O_1963,N_14896,N_14892);
nor UO_1964 (O_1964,N_14906,N_14872);
or UO_1965 (O_1965,N_14885,N_14907);
nand UO_1966 (O_1966,N_14851,N_14914);
nand UO_1967 (O_1967,N_14856,N_14957);
nor UO_1968 (O_1968,N_14860,N_14940);
or UO_1969 (O_1969,N_14911,N_14903);
or UO_1970 (O_1970,N_14867,N_14949);
nand UO_1971 (O_1971,N_14865,N_14925);
nand UO_1972 (O_1972,N_14934,N_14877);
nand UO_1973 (O_1973,N_14948,N_14934);
xor UO_1974 (O_1974,N_14989,N_14969);
nor UO_1975 (O_1975,N_14898,N_14860);
nand UO_1976 (O_1976,N_14950,N_14879);
and UO_1977 (O_1977,N_14927,N_14968);
xnor UO_1978 (O_1978,N_14913,N_14865);
and UO_1979 (O_1979,N_14911,N_14915);
and UO_1980 (O_1980,N_14860,N_14987);
nor UO_1981 (O_1981,N_14865,N_14917);
nor UO_1982 (O_1982,N_14852,N_14907);
xnor UO_1983 (O_1983,N_14918,N_14997);
and UO_1984 (O_1984,N_14963,N_14908);
nand UO_1985 (O_1985,N_14927,N_14897);
or UO_1986 (O_1986,N_14865,N_14883);
nand UO_1987 (O_1987,N_14908,N_14918);
or UO_1988 (O_1988,N_14852,N_14925);
xnor UO_1989 (O_1989,N_14887,N_14899);
and UO_1990 (O_1990,N_14928,N_14911);
or UO_1991 (O_1991,N_14977,N_14980);
or UO_1992 (O_1992,N_14915,N_14982);
xor UO_1993 (O_1993,N_14967,N_14910);
nor UO_1994 (O_1994,N_14967,N_14906);
nor UO_1995 (O_1995,N_14960,N_14856);
nand UO_1996 (O_1996,N_14891,N_14994);
and UO_1997 (O_1997,N_14909,N_14871);
or UO_1998 (O_1998,N_14855,N_14859);
nand UO_1999 (O_1999,N_14923,N_14905);
endmodule