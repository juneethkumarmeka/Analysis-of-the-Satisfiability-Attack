module basic_750_5000_1000_5_levels_1xor_9(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
or U0 (N_0,In_323,In_417);
and U1 (N_1,In_521,In_454);
and U2 (N_2,In_382,In_407);
and U3 (N_3,In_44,In_485);
xor U4 (N_4,In_303,In_476);
or U5 (N_5,In_171,In_673);
nor U6 (N_6,In_462,In_448);
and U7 (N_7,In_88,In_249);
or U8 (N_8,In_165,In_368);
and U9 (N_9,In_461,In_341);
or U10 (N_10,In_99,In_439);
and U11 (N_11,In_525,In_39);
nand U12 (N_12,In_213,In_666);
and U13 (N_13,In_0,In_327);
nand U14 (N_14,In_189,In_505);
and U15 (N_15,In_349,In_107);
nor U16 (N_16,In_43,In_489);
and U17 (N_17,In_124,In_490);
or U18 (N_18,In_64,In_394);
nor U19 (N_19,In_142,In_616);
nor U20 (N_20,In_528,In_231);
or U21 (N_21,In_289,In_545);
and U22 (N_22,In_531,In_533);
or U23 (N_23,In_274,In_593);
or U24 (N_24,In_672,In_187);
and U25 (N_25,In_66,In_60);
nor U26 (N_26,In_559,In_728);
or U27 (N_27,In_63,In_282);
nand U28 (N_28,In_603,In_431);
nand U29 (N_29,In_591,In_413);
nor U30 (N_30,In_714,In_319);
nor U31 (N_31,In_281,In_152);
and U32 (N_32,In_4,In_625);
and U33 (N_33,In_600,In_446);
nand U34 (N_34,In_713,In_638);
or U35 (N_35,In_538,In_79);
nor U36 (N_36,In_566,In_710);
or U37 (N_37,In_55,In_73);
nor U38 (N_38,In_720,In_364);
or U39 (N_39,In_381,In_23);
nand U40 (N_40,In_61,In_272);
nor U41 (N_41,In_84,In_645);
or U42 (N_42,In_547,In_300);
nand U43 (N_43,In_299,In_238);
nor U44 (N_44,In_614,In_258);
nor U45 (N_45,In_575,In_749);
nand U46 (N_46,In_199,In_702);
nor U47 (N_47,In_352,In_144);
nor U48 (N_48,In_599,In_111);
nand U49 (N_49,In_255,In_346);
nor U50 (N_50,In_733,In_378);
or U51 (N_51,In_71,In_83);
or U52 (N_52,In_594,In_340);
nand U53 (N_53,In_100,In_621);
nand U54 (N_54,In_206,In_504);
nor U55 (N_55,In_17,In_421);
xnor U56 (N_56,In_304,In_511);
and U57 (N_57,In_656,In_706);
nor U58 (N_58,In_363,In_522);
nor U59 (N_59,In_445,In_471);
nand U60 (N_60,In_130,In_606);
nor U61 (N_61,In_338,In_390);
or U62 (N_62,In_653,In_428);
nor U63 (N_63,In_290,In_184);
and U64 (N_64,In_21,In_316);
or U65 (N_65,In_365,In_174);
nand U66 (N_66,In_337,In_440);
nor U67 (N_67,In_432,In_496);
nor U68 (N_68,In_226,In_333);
nor U69 (N_69,In_186,In_604);
and U70 (N_70,In_267,In_134);
or U71 (N_71,In_208,In_123);
or U72 (N_72,In_644,In_302);
and U73 (N_73,In_449,In_564);
nand U74 (N_74,In_580,In_483);
and U75 (N_75,In_217,In_177);
and U76 (N_76,In_307,In_135);
nor U77 (N_77,In_204,In_326);
and U78 (N_78,In_414,In_59);
and U79 (N_79,In_450,In_48);
nor U80 (N_80,In_585,In_509);
nor U81 (N_81,In_242,In_336);
or U82 (N_82,In_607,In_699);
nand U83 (N_83,In_278,In_424);
nor U84 (N_84,In_704,In_369);
or U85 (N_85,In_532,In_136);
nor U86 (N_86,In_370,In_596);
nand U87 (N_87,In_551,In_542);
or U88 (N_88,In_172,In_16);
xor U89 (N_89,In_402,In_259);
and U90 (N_90,In_403,In_510);
nand U91 (N_91,In_423,In_126);
nand U92 (N_92,In_694,In_253);
nor U93 (N_93,In_711,In_161);
nand U94 (N_94,In_7,In_548);
nor U95 (N_95,In_32,In_194);
nor U96 (N_96,In_419,In_313);
and U97 (N_97,In_487,In_434);
or U98 (N_98,In_641,In_516);
nor U99 (N_99,In_457,In_701);
or U100 (N_100,In_555,In_214);
and U101 (N_101,In_425,In_650);
or U102 (N_102,In_75,In_149);
nor U103 (N_103,In_26,In_264);
nor U104 (N_104,In_193,In_718);
nand U105 (N_105,In_544,In_72);
or U106 (N_106,In_148,In_245);
nand U107 (N_107,In_597,In_467);
or U108 (N_108,In_668,In_230);
nand U109 (N_109,In_624,In_375);
and U110 (N_110,In_464,In_309);
or U111 (N_111,In_380,In_203);
nor U112 (N_112,In_328,In_637);
or U113 (N_113,In_164,In_477);
or U114 (N_114,In_721,In_411);
or U115 (N_115,In_9,In_583);
and U116 (N_116,In_279,In_590);
nor U117 (N_117,In_97,In_92);
nand U118 (N_118,In_655,In_615);
or U119 (N_119,In_125,In_629);
or U120 (N_120,In_141,In_652);
nor U121 (N_121,In_717,In_58);
nand U122 (N_122,In_235,In_420);
nor U123 (N_123,In_85,In_488);
nor U124 (N_124,In_497,In_169);
nand U125 (N_125,In_246,In_686);
and U126 (N_126,In_353,In_628);
nand U127 (N_127,In_620,In_513);
or U128 (N_128,In_395,In_315);
nand U129 (N_129,In_318,In_680);
nor U130 (N_130,In_133,In_601);
nand U131 (N_131,In_35,In_158);
nand U132 (N_132,In_503,In_38);
nor U133 (N_133,In_581,In_687);
nor U134 (N_134,In_173,In_605);
nor U135 (N_135,In_740,In_140);
and U136 (N_136,In_563,In_371);
nand U137 (N_137,In_348,In_106);
nand U138 (N_138,In_103,In_465);
and U139 (N_139,In_62,In_356);
or U140 (N_140,In_659,In_286);
nand U141 (N_141,In_660,In_216);
or U142 (N_142,In_639,In_310);
and U143 (N_143,In_81,In_466);
or U144 (N_144,In_37,In_735);
nand U145 (N_145,In_667,In_202);
and U146 (N_146,In_447,In_13);
or U147 (N_147,In_225,In_138);
and U148 (N_148,In_479,In_578);
nand U149 (N_149,In_143,In_3);
nor U150 (N_150,In_192,In_478);
nand U151 (N_151,In_69,In_287);
or U152 (N_152,In_263,In_53);
nor U153 (N_153,In_561,In_619);
nand U154 (N_154,In_308,In_345);
nor U155 (N_155,In_635,In_670);
nor U156 (N_156,In_507,In_705);
nand U157 (N_157,In_543,In_367);
and U158 (N_158,In_347,In_209);
nand U159 (N_159,In_181,In_18);
nor U160 (N_160,In_95,In_685);
nand U161 (N_161,In_211,In_669);
nor U162 (N_162,In_212,In_384);
or U163 (N_163,In_87,In_683);
xnor U164 (N_164,In_643,In_730);
nand U165 (N_165,In_10,In_560);
or U166 (N_166,In_709,In_738);
or U167 (N_167,In_396,In_233);
nor U168 (N_168,In_321,In_374);
and U169 (N_169,In_684,In_529);
nor U170 (N_170,In_314,In_692);
nor U171 (N_171,In_618,In_159);
and U172 (N_172,In_351,In_15);
nand U173 (N_173,In_400,In_250);
nand U174 (N_174,In_359,In_435);
nand U175 (N_175,In_523,In_636);
nand U176 (N_176,In_535,In_220);
and U177 (N_177,In_160,In_569);
nand U178 (N_178,In_179,In_554);
and U179 (N_179,In_28,In_549);
nand U180 (N_180,In_571,In_248);
nand U181 (N_181,In_546,In_630);
or U182 (N_182,In_147,In_501);
nor U183 (N_183,In_305,In_582);
nand U184 (N_184,In_320,In_361);
or U185 (N_185,In_224,In_33);
nor U186 (N_186,In_726,In_584);
and U187 (N_187,In_362,In_12);
nor U188 (N_188,In_240,In_86);
or U189 (N_189,In_681,In_283);
nand U190 (N_190,In_422,In_167);
and U191 (N_191,In_222,In_696);
nand U192 (N_192,In_661,In_139);
and U193 (N_193,In_470,In_617);
or U194 (N_194,In_241,In_312);
nand U195 (N_195,In_25,In_688);
and U196 (N_196,In_389,In_627);
nand U197 (N_197,In_116,In_530);
nor U198 (N_198,In_708,In_634);
nor U199 (N_199,In_266,In_460);
nor U200 (N_200,In_19,In_405);
nand U201 (N_201,In_611,In_243);
nand U202 (N_202,In_553,In_577);
nand U203 (N_203,In_24,In_132);
or U204 (N_204,In_385,In_1);
nand U205 (N_205,In_188,In_256);
or U206 (N_206,In_56,In_589);
or U207 (N_207,In_11,In_739);
nand U208 (N_208,In_301,In_647);
and U209 (N_209,In_429,In_244);
and U210 (N_210,In_120,In_335);
or U211 (N_211,In_418,In_502);
nand U212 (N_212,In_49,In_68);
xnor U213 (N_213,In_157,In_292);
nand U214 (N_214,In_689,In_745);
nor U215 (N_215,In_398,In_379);
nor U216 (N_216,In_52,In_74);
xnor U217 (N_217,In_567,In_646);
nand U218 (N_218,In_27,In_703);
nand U219 (N_219,In_732,In_67);
and U220 (N_220,In_237,In_122);
nor U221 (N_221,In_500,In_664);
and U222 (N_222,In_288,In_119);
or U223 (N_223,In_261,In_196);
nor U224 (N_224,In_269,In_262);
and U225 (N_225,In_239,In_118);
and U226 (N_226,In_633,In_127);
nand U227 (N_227,In_154,In_695);
nor U228 (N_228,In_610,In_234);
nand U229 (N_229,In_552,In_153);
and U230 (N_230,In_30,In_499);
nand U231 (N_231,In_608,In_273);
nand U232 (N_232,In_441,In_558);
nor U233 (N_233,In_46,In_406);
nand U234 (N_234,In_155,In_562);
nand U235 (N_235,In_185,In_678);
nand U236 (N_236,In_393,In_207);
and U237 (N_237,In_276,In_227);
nor U238 (N_238,In_190,In_388);
and U239 (N_239,In_50,In_724);
or U240 (N_240,In_463,In_156);
nand U241 (N_241,In_570,In_451);
and U242 (N_242,In_453,In_372);
nand U243 (N_243,In_108,In_498);
nor U244 (N_244,In_40,In_251);
or U245 (N_245,In_275,In_105);
nand U246 (N_246,In_195,In_293);
or U247 (N_247,In_342,In_14);
nand U248 (N_248,In_679,In_725);
or U249 (N_249,In_729,In_70);
nand U250 (N_250,In_2,In_587);
nand U251 (N_251,In_183,In_537);
nand U252 (N_252,In_662,In_257);
xor U253 (N_253,In_182,In_254);
nor U254 (N_254,In_205,In_722);
nand U255 (N_255,In_663,In_514);
or U256 (N_256,In_332,In_524);
or U257 (N_257,In_376,In_416);
or U258 (N_258,In_145,In_576);
nand U259 (N_259,In_109,In_518);
and U260 (N_260,In_329,In_744);
and U261 (N_261,In_715,In_442);
nand U262 (N_262,In_383,In_612);
or U263 (N_263,In_459,In_215);
or U264 (N_264,In_102,In_654);
or U265 (N_265,In_210,In_350);
or U266 (N_266,In_331,In_175);
or U267 (N_267,In_539,In_178);
nand U268 (N_268,In_41,In_343);
and U269 (N_269,In_42,In_77);
or U270 (N_270,In_360,In_676);
nand U271 (N_271,In_65,In_712);
nor U272 (N_272,In_236,In_291);
nand U273 (N_273,In_520,In_201);
nor U274 (N_274,In_592,In_622);
or U275 (N_275,In_412,In_298);
and U276 (N_276,In_354,In_579);
and U277 (N_277,In_426,In_723);
nor U278 (N_278,In_166,In_677);
nand U279 (N_279,In_748,In_115);
nor U280 (N_280,In_430,In_716);
and U281 (N_281,In_146,In_737);
nand U282 (N_282,In_339,In_306);
or U283 (N_283,In_180,In_588);
nand U284 (N_284,In_556,In_613);
nor U285 (N_285,In_191,In_91);
or U286 (N_286,In_437,In_640);
nor U287 (N_287,In_280,In_736);
nor U288 (N_288,In_508,In_741);
nand U289 (N_289,In_117,In_492);
and U290 (N_290,In_129,In_334);
and U291 (N_291,In_47,In_691);
nand U292 (N_292,In_493,In_151);
or U293 (N_293,In_480,In_330);
nor U294 (N_294,In_527,In_541);
nand U295 (N_295,In_260,In_410);
nand U296 (N_296,In_658,In_131);
or U297 (N_297,In_82,In_540);
nand U298 (N_298,In_344,In_631);
nand U299 (N_299,In_693,In_358);
nor U300 (N_300,In_742,In_671);
nand U301 (N_301,In_475,In_626);
or U302 (N_302,In_455,In_357);
nand U303 (N_303,In_6,In_574);
nor U304 (N_304,In_268,In_697);
and U305 (N_305,In_651,In_317);
or U306 (N_306,In_114,In_150);
or U307 (N_307,In_557,In_648);
and U308 (N_308,In_98,In_8);
nor U309 (N_309,In_270,In_128);
or U310 (N_310,In_22,In_265);
nor U311 (N_311,In_387,In_29);
or U312 (N_312,In_104,In_391);
or U313 (N_313,In_200,In_284);
nand U314 (N_314,In_93,In_386);
or U315 (N_315,In_609,In_5);
or U316 (N_316,In_57,In_573);
or U317 (N_317,In_456,In_586);
and U318 (N_318,In_649,In_452);
nor U319 (N_319,In_436,In_366);
and U320 (N_320,In_443,In_473);
nor U321 (N_321,In_285,In_271);
and U322 (N_322,In_698,In_743);
and U323 (N_323,In_565,In_45);
and U324 (N_324,In_322,In_469);
and U325 (N_325,In_484,In_198);
and U326 (N_326,In_294,In_137);
nor U327 (N_327,In_163,In_598);
nand U328 (N_328,In_168,In_197);
nor U329 (N_329,In_427,In_34);
nor U330 (N_330,In_415,In_229);
and U331 (N_331,In_221,In_623);
and U332 (N_332,In_731,In_700);
or U333 (N_333,In_632,In_550);
or U334 (N_334,In_665,In_162);
nor U335 (N_335,In_657,In_719);
nor U336 (N_336,In_727,In_232);
and U337 (N_337,In_392,In_80);
or U338 (N_338,In_486,In_495);
or U339 (N_339,In_31,In_247);
and U340 (N_340,In_474,In_94);
and U341 (N_341,In_519,In_517);
or U342 (N_342,In_494,In_90);
xor U343 (N_343,In_399,In_295);
or U344 (N_344,In_96,In_20);
nand U345 (N_345,In_482,In_112);
nor U346 (N_346,In_682,In_277);
and U347 (N_347,In_642,In_444);
or U348 (N_348,In_409,In_572);
or U349 (N_349,In_76,In_404);
and U350 (N_350,In_401,In_223);
nor U351 (N_351,In_481,In_675);
nand U352 (N_352,In_674,In_707);
or U353 (N_353,In_113,In_170);
and U354 (N_354,In_408,In_311);
or U355 (N_355,In_472,In_89);
nor U356 (N_356,In_252,In_506);
nand U357 (N_357,In_433,In_54);
and U358 (N_358,In_568,In_110);
or U359 (N_359,In_746,In_36);
and U360 (N_360,In_602,In_296);
nor U361 (N_361,In_595,In_78);
or U362 (N_362,In_219,In_526);
and U363 (N_363,In_101,In_373);
nor U364 (N_364,In_536,In_734);
or U365 (N_365,In_534,In_468);
nor U366 (N_366,In_228,In_325);
nor U367 (N_367,In_355,In_297);
nor U368 (N_368,In_747,In_512);
and U369 (N_369,In_377,In_121);
and U370 (N_370,In_324,In_515);
nand U371 (N_371,In_176,In_218);
and U372 (N_372,In_458,In_690);
or U373 (N_373,In_491,In_438);
nand U374 (N_374,In_51,In_397);
nor U375 (N_375,In_442,In_478);
or U376 (N_376,In_505,In_548);
nor U377 (N_377,In_1,In_334);
or U378 (N_378,In_446,In_68);
or U379 (N_379,In_432,In_35);
nor U380 (N_380,In_624,In_491);
nor U381 (N_381,In_483,In_378);
and U382 (N_382,In_220,In_12);
and U383 (N_383,In_236,In_437);
or U384 (N_384,In_466,In_676);
nand U385 (N_385,In_32,In_284);
or U386 (N_386,In_698,In_565);
nand U387 (N_387,In_688,In_110);
nand U388 (N_388,In_498,In_471);
nand U389 (N_389,In_507,In_537);
and U390 (N_390,In_190,In_154);
and U391 (N_391,In_278,In_454);
and U392 (N_392,In_507,In_249);
or U393 (N_393,In_394,In_13);
and U394 (N_394,In_65,In_708);
or U395 (N_395,In_646,In_31);
nor U396 (N_396,In_459,In_48);
nand U397 (N_397,In_504,In_325);
nand U398 (N_398,In_42,In_449);
and U399 (N_399,In_688,In_383);
or U400 (N_400,In_232,In_138);
nor U401 (N_401,In_171,In_276);
nand U402 (N_402,In_217,In_725);
and U403 (N_403,In_555,In_106);
or U404 (N_404,In_6,In_235);
and U405 (N_405,In_701,In_372);
nor U406 (N_406,In_204,In_397);
and U407 (N_407,In_362,In_463);
and U408 (N_408,In_3,In_408);
and U409 (N_409,In_135,In_231);
nor U410 (N_410,In_138,In_312);
and U411 (N_411,In_233,In_34);
nor U412 (N_412,In_720,In_199);
or U413 (N_413,In_51,In_523);
nand U414 (N_414,In_738,In_453);
xor U415 (N_415,In_136,In_448);
and U416 (N_416,In_521,In_308);
and U417 (N_417,In_7,In_509);
and U418 (N_418,In_466,In_730);
and U419 (N_419,In_208,In_232);
nor U420 (N_420,In_419,In_571);
nor U421 (N_421,In_238,In_711);
nor U422 (N_422,In_297,In_111);
or U423 (N_423,In_743,In_614);
nand U424 (N_424,In_12,In_400);
and U425 (N_425,In_486,In_666);
and U426 (N_426,In_0,In_129);
and U427 (N_427,In_167,In_281);
or U428 (N_428,In_282,In_208);
nand U429 (N_429,In_604,In_598);
and U430 (N_430,In_584,In_499);
nand U431 (N_431,In_709,In_146);
or U432 (N_432,In_17,In_135);
and U433 (N_433,In_40,In_7);
nand U434 (N_434,In_584,In_520);
or U435 (N_435,In_141,In_54);
nand U436 (N_436,In_547,In_150);
nor U437 (N_437,In_55,In_517);
nor U438 (N_438,In_149,In_552);
or U439 (N_439,In_526,In_594);
and U440 (N_440,In_233,In_539);
nand U441 (N_441,In_257,In_407);
nand U442 (N_442,In_353,In_120);
nor U443 (N_443,In_183,In_261);
nor U444 (N_444,In_129,In_1);
or U445 (N_445,In_628,In_166);
nand U446 (N_446,In_278,In_204);
nand U447 (N_447,In_551,In_616);
nor U448 (N_448,In_643,In_542);
and U449 (N_449,In_443,In_209);
and U450 (N_450,In_483,In_283);
nor U451 (N_451,In_363,In_679);
or U452 (N_452,In_262,In_16);
nand U453 (N_453,In_300,In_150);
nand U454 (N_454,In_124,In_82);
nand U455 (N_455,In_330,In_580);
or U456 (N_456,In_463,In_123);
nand U457 (N_457,In_429,In_632);
or U458 (N_458,In_123,In_568);
or U459 (N_459,In_177,In_144);
nor U460 (N_460,In_472,In_491);
nand U461 (N_461,In_671,In_538);
nand U462 (N_462,In_32,In_103);
nor U463 (N_463,In_371,In_67);
nand U464 (N_464,In_653,In_108);
nor U465 (N_465,In_568,In_84);
and U466 (N_466,In_732,In_347);
or U467 (N_467,In_550,In_700);
and U468 (N_468,In_369,In_59);
nand U469 (N_469,In_54,In_635);
and U470 (N_470,In_18,In_440);
nand U471 (N_471,In_78,In_161);
or U472 (N_472,In_551,In_273);
nand U473 (N_473,In_186,In_237);
nand U474 (N_474,In_307,In_291);
and U475 (N_475,In_104,In_586);
nand U476 (N_476,In_683,In_436);
and U477 (N_477,In_592,In_189);
nand U478 (N_478,In_548,In_22);
and U479 (N_479,In_272,In_237);
nor U480 (N_480,In_53,In_508);
or U481 (N_481,In_391,In_52);
nand U482 (N_482,In_112,In_480);
nor U483 (N_483,In_405,In_20);
or U484 (N_484,In_86,In_142);
or U485 (N_485,In_412,In_273);
nand U486 (N_486,In_597,In_87);
and U487 (N_487,In_352,In_242);
and U488 (N_488,In_42,In_673);
or U489 (N_489,In_382,In_432);
nor U490 (N_490,In_112,In_140);
or U491 (N_491,In_729,In_56);
nand U492 (N_492,In_561,In_364);
nor U493 (N_493,In_326,In_580);
nand U494 (N_494,In_435,In_176);
and U495 (N_495,In_572,In_469);
nor U496 (N_496,In_582,In_178);
or U497 (N_497,In_388,In_637);
or U498 (N_498,In_252,In_439);
nand U499 (N_499,In_472,In_389);
nand U500 (N_500,In_54,In_729);
nand U501 (N_501,In_154,In_3);
or U502 (N_502,In_106,In_33);
or U503 (N_503,In_456,In_541);
nor U504 (N_504,In_304,In_721);
or U505 (N_505,In_668,In_599);
and U506 (N_506,In_599,In_312);
nor U507 (N_507,In_581,In_43);
nand U508 (N_508,In_703,In_88);
and U509 (N_509,In_126,In_653);
and U510 (N_510,In_502,In_426);
or U511 (N_511,In_437,In_581);
nor U512 (N_512,In_460,In_551);
and U513 (N_513,In_379,In_0);
and U514 (N_514,In_275,In_527);
nor U515 (N_515,In_267,In_268);
or U516 (N_516,In_545,In_451);
and U517 (N_517,In_565,In_450);
xor U518 (N_518,In_741,In_57);
and U519 (N_519,In_239,In_553);
nor U520 (N_520,In_609,In_529);
nor U521 (N_521,In_211,In_355);
xnor U522 (N_522,In_284,In_199);
nand U523 (N_523,In_48,In_540);
nand U524 (N_524,In_535,In_122);
nand U525 (N_525,In_48,In_743);
nor U526 (N_526,In_148,In_465);
and U527 (N_527,In_619,In_75);
nand U528 (N_528,In_8,In_562);
or U529 (N_529,In_274,In_14);
nand U530 (N_530,In_156,In_280);
or U531 (N_531,In_170,In_580);
or U532 (N_532,In_577,In_107);
and U533 (N_533,In_482,In_383);
nand U534 (N_534,In_492,In_292);
nor U535 (N_535,In_362,In_636);
or U536 (N_536,In_8,In_740);
nand U537 (N_537,In_411,In_551);
nor U538 (N_538,In_104,In_347);
nand U539 (N_539,In_722,In_322);
and U540 (N_540,In_378,In_647);
and U541 (N_541,In_55,In_345);
nand U542 (N_542,In_514,In_192);
or U543 (N_543,In_648,In_278);
nand U544 (N_544,In_632,In_174);
or U545 (N_545,In_270,In_582);
nand U546 (N_546,In_59,In_31);
or U547 (N_547,In_635,In_92);
nand U548 (N_548,In_87,In_142);
or U549 (N_549,In_407,In_18);
or U550 (N_550,In_70,In_736);
and U551 (N_551,In_287,In_449);
nand U552 (N_552,In_746,In_383);
nor U553 (N_553,In_535,In_51);
nor U554 (N_554,In_107,In_56);
and U555 (N_555,In_559,In_684);
nor U556 (N_556,In_406,In_635);
and U557 (N_557,In_294,In_95);
or U558 (N_558,In_152,In_17);
nand U559 (N_559,In_244,In_350);
nand U560 (N_560,In_475,In_99);
nand U561 (N_561,In_153,In_67);
nor U562 (N_562,In_282,In_731);
or U563 (N_563,In_326,In_245);
and U564 (N_564,In_542,In_461);
and U565 (N_565,In_115,In_228);
or U566 (N_566,In_383,In_606);
xor U567 (N_567,In_569,In_96);
and U568 (N_568,In_40,In_155);
or U569 (N_569,In_116,In_547);
nor U570 (N_570,In_607,In_153);
nor U571 (N_571,In_64,In_68);
nand U572 (N_572,In_621,In_282);
nand U573 (N_573,In_529,In_291);
or U574 (N_574,In_678,In_137);
nor U575 (N_575,In_721,In_621);
or U576 (N_576,In_493,In_290);
and U577 (N_577,In_537,In_157);
nand U578 (N_578,In_150,In_468);
nor U579 (N_579,In_256,In_675);
or U580 (N_580,In_274,In_306);
nor U581 (N_581,In_456,In_699);
nor U582 (N_582,In_375,In_410);
nand U583 (N_583,In_413,In_739);
nor U584 (N_584,In_205,In_671);
and U585 (N_585,In_519,In_311);
and U586 (N_586,In_603,In_707);
and U587 (N_587,In_685,In_362);
nor U588 (N_588,In_73,In_56);
and U589 (N_589,In_463,In_739);
or U590 (N_590,In_682,In_717);
and U591 (N_591,In_37,In_273);
nand U592 (N_592,In_141,In_174);
or U593 (N_593,In_410,In_101);
nor U594 (N_594,In_393,In_645);
and U595 (N_595,In_449,In_120);
nand U596 (N_596,In_195,In_218);
nor U597 (N_597,In_128,In_716);
and U598 (N_598,In_301,In_271);
and U599 (N_599,In_213,In_577);
nand U600 (N_600,In_341,In_17);
nor U601 (N_601,In_484,In_725);
or U602 (N_602,In_662,In_74);
or U603 (N_603,In_396,In_99);
nand U604 (N_604,In_669,In_115);
nor U605 (N_605,In_725,In_25);
nand U606 (N_606,In_545,In_86);
nor U607 (N_607,In_75,In_596);
and U608 (N_608,In_36,In_167);
nand U609 (N_609,In_392,In_305);
or U610 (N_610,In_377,In_592);
and U611 (N_611,In_248,In_738);
nand U612 (N_612,In_510,In_710);
nand U613 (N_613,In_216,In_465);
nand U614 (N_614,In_715,In_315);
or U615 (N_615,In_572,In_670);
and U616 (N_616,In_474,In_113);
nor U617 (N_617,In_425,In_195);
nor U618 (N_618,In_461,In_610);
or U619 (N_619,In_567,In_370);
nor U620 (N_620,In_48,In_94);
nand U621 (N_621,In_238,In_119);
nand U622 (N_622,In_17,In_547);
or U623 (N_623,In_735,In_730);
nor U624 (N_624,In_160,In_724);
or U625 (N_625,In_508,In_490);
and U626 (N_626,In_319,In_527);
or U627 (N_627,In_253,In_214);
nor U628 (N_628,In_120,In_398);
or U629 (N_629,In_650,In_642);
and U630 (N_630,In_716,In_110);
or U631 (N_631,In_593,In_121);
nand U632 (N_632,In_351,In_499);
or U633 (N_633,In_379,In_697);
and U634 (N_634,In_510,In_601);
nand U635 (N_635,In_573,In_136);
nand U636 (N_636,In_98,In_396);
nand U637 (N_637,In_299,In_53);
and U638 (N_638,In_95,In_195);
and U639 (N_639,In_664,In_302);
nor U640 (N_640,In_643,In_81);
or U641 (N_641,In_731,In_399);
or U642 (N_642,In_291,In_371);
nor U643 (N_643,In_627,In_275);
nor U644 (N_644,In_282,In_555);
and U645 (N_645,In_629,In_585);
nor U646 (N_646,In_532,In_359);
nor U647 (N_647,In_249,In_717);
nor U648 (N_648,In_153,In_628);
nand U649 (N_649,In_554,In_528);
nand U650 (N_650,In_371,In_581);
nand U651 (N_651,In_103,In_237);
nor U652 (N_652,In_76,In_341);
and U653 (N_653,In_333,In_707);
or U654 (N_654,In_417,In_479);
nand U655 (N_655,In_466,In_481);
nor U656 (N_656,In_467,In_247);
and U657 (N_657,In_552,In_94);
and U658 (N_658,In_588,In_734);
nor U659 (N_659,In_380,In_45);
nand U660 (N_660,In_505,In_255);
nand U661 (N_661,In_383,In_117);
and U662 (N_662,In_506,In_25);
nor U663 (N_663,In_596,In_212);
or U664 (N_664,In_182,In_600);
nor U665 (N_665,In_528,In_570);
nand U666 (N_666,In_658,In_558);
and U667 (N_667,In_185,In_501);
nor U668 (N_668,In_60,In_147);
nor U669 (N_669,In_308,In_257);
or U670 (N_670,In_354,In_713);
or U671 (N_671,In_444,In_363);
or U672 (N_672,In_6,In_605);
nand U673 (N_673,In_703,In_335);
nor U674 (N_674,In_420,In_126);
nand U675 (N_675,In_114,In_292);
nand U676 (N_676,In_108,In_514);
nand U677 (N_677,In_621,In_647);
nor U678 (N_678,In_435,In_368);
and U679 (N_679,In_116,In_558);
or U680 (N_680,In_115,In_80);
or U681 (N_681,In_468,In_121);
or U682 (N_682,In_7,In_279);
nor U683 (N_683,In_54,In_529);
and U684 (N_684,In_5,In_622);
nand U685 (N_685,In_391,In_322);
and U686 (N_686,In_245,In_353);
and U687 (N_687,In_186,In_106);
nor U688 (N_688,In_141,In_417);
nand U689 (N_689,In_187,In_725);
and U690 (N_690,In_94,In_710);
and U691 (N_691,In_346,In_294);
nand U692 (N_692,In_144,In_165);
or U693 (N_693,In_370,In_582);
nor U694 (N_694,In_476,In_453);
and U695 (N_695,In_415,In_358);
nor U696 (N_696,In_237,In_605);
or U697 (N_697,In_302,In_330);
or U698 (N_698,In_542,In_529);
or U699 (N_699,In_335,In_414);
or U700 (N_700,In_575,In_397);
nor U701 (N_701,In_104,In_57);
or U702 (N_702,In_14,In_733);
nor U703 (N_703,In_424,In_175);
xnor U704 (N_704,In_583,In_286);
nand U705 (N_705,In_305,In_402);
nor U706 (N_706,In_404,In_200);
nor U707 (N_707,In_288,In_329);
or U708 (N_708,In_431,In_607);
nor U709 (N_709,In_676,In_206);
and U710 (N_710,In_724,In_567);
or U711 (N_711,In_375,In_379);
nand U712 (N_712,In_141,In_188);
or U713 (N_713,In_203,In_510);
and U714 (N_714,In_358,In_120);
nand U715 (N_715,In_629,In_430);
or U716 (N_716,In_731,In_631);
nor U717 (N_717,In_562,In_611);
or U718 (N_718,In_675,In_57);
and U719 (N_719,In_471,In_143);
nand U720 (N_720,In_496,In_167);
and U721 (N_721,In_501,In_152);
nand U722 (N_722,In_437,In_721);
or U723 (N_723,In_439,In_12);
or U724 (N_724,In_288,In_430);
or U725 (N_725,In_441,In_411);
nor U726 (N_726,In_299,In_487);
and U727 (N_727,In_716,In_372);
nor U728 (N_728,In_209,In_358);
or U729 (N_729,In_331,In_111);
or U730 (N_730,In_550,In_664);
nand U731 (N_731,In_220,In_14);
or U732 (N_732,In_176,In_167);
nand U733 (N_733,In_348,In_238);
nand U734 (N_734,In_471,In_621);
nand U735 (N_735,In_645,In_463);
and U736 (N_736,In_244,In_293);
nor U737 (N_737,In_483,In_596);
and U738 (N_738,In_117,In_286);
nor U739 (N_739,In_527,In_713);
or U740 (N_740,In_240,In_245);
or U741 (N_741,In_233,In_251);
and U742 (N_742,In_190,In_287);
or U743 (N_743,In_271,In_142);
or U744 (N_744,In_568,In_223);
and U745 (N_745,In_710,In_360);
nand U746 (N_746,In_693,In_45);
or U747 (N_747,In_300,In_31);
nand U748 (N_748,In_418,In_123);
nor U749 (N_749,In_124,In_17);
and U750 (N_750,In_356,In_454);
nand U751 (N_751,In_555,In_179);
nor U752 (N_752,In_126,In_330);
or U753 (N_753,In_329,In_466);
or U754 (N_754,In_502,In_31);
nand U755 (N_755,In_197,In_402);
nor U756 (N_756,In_640,In_67);
nand U757 (N_757,In_22,In_172);
and U758 (N_758,In_451,In_521);
or U759 (N_759,In_294,In_482);
or U760 (N_760,In_191,In_428);
and U761 (N_761,In_380,In_117);
or U762 (N_762,In_308,In_58);
or U763 (N_763,In_290,In_491);
and U764 (N_764,In_690,In_120);
or U765 (N_765,In_523,In_683);
xnor U766 (N_766,In_203,In_456);
nor U767 (N_767,In_412,In_480);
nor U768 (N_768,In_651,In_275);
or U769 (N_769,In_19,In_15);
nor U770 (N_770,In_681,In_114);
and U771 (N_771,In_291,In_211);
and U772 (N_772,In_603,In_667);
or U773 (N_773,In_461,In_671);
or U774 (N_774,In_599,In_130);
xor U775 (N_775,In_96,In_394);
nand U776 (N_776,In_119,In_628);
nand U777 (N_777,In_159,In_337);
nor U778 (N_778,In_51,In_490);
and U779 (N_779,In_51,In_314);
nor U780 (N_780,In_26,In_126);
or U781 (N_781,In_714,In_289);
or U782 (N_782,In_720,In_188);
or U783 (N_783,In_740,In_569);
nand U784 (N_784,In_262,In_631);
nor U785 (N_785,In_708,In_223);
and U786 (N_786,In_362,In_662);
and U787 (N_787,In_539,In_125);
nand U788 (N_788,In_590,In_159);
and U789 (N_789,In_489,In_368);
nand U790 (N_790,In_398,In_234);
or U791 (N_791,In_361,In_337);
nor U792 (N_792,In_539,In_186);
nand U793 (N_793,In_116,In_58);
and U794 (N_794,In_26,In_715);
or U795 (N_795,In_370,In_533);
xor U796 (N_796,In_241,In_629);
nand U797 (N_797,In_176,In_94);
nor U798 (N_798,In_737,In_642);
nand U799 (N_799,In_658,In_512);
or U800 (N_800,In_639,In_603);
nor U801 (N_801,In_527,In_288);
or U802 (N_802,In_319,In_9);
or U803 (N_803,In_162,In_463);
nor U804 (N_804,In_726,In_683);
nor U805 (N_805,In_641,In_522);
and U806 (N_806,In_419,In_637);
and U807 (N_807,In_543,In_630);
nor U808 (N_808,In_610,In_691);
xnor U809 (N_809,In_162,In_565);
nand U810 (N_810,In_251,In_707);
nand U811 (N_811,In_107,In_680);
nand U812 (N_812,In_163,In_245);
nor U813 (N_813,In_292,In_347);
nand U814 (N_814,In_449,In_180);
or U815 (N_815,In_347,In_477);
and U816 (N_816,In_78,In_659);
nand U817 (N_817,In_644,In_716);
or U818 (N_818,In_409,In_45);
or U819 (N_819,In_121,In_127);
nand U820 (N_820,In_291,In_420);
nand U821 (N_821,In_740,In_602);
and U822 (N_822,In_273,In_602);
or U823 (N_823,In_674,In_289);
or U824 (N_824,In_480,In_61);
and U825 (N_825,In_383,In_561);
nor U826 (N_826,In_459,In_255);
nor U827 (N_827,In_51,In_704);
or U828 (N_828,In_155,In_187);
nand U829 (N_829,In_455,In_628);
nand U830 (N_830,In_45,In_581);
and U831 (N_831,In_165,In_503);
nand U832 (N_832,In_535,In_251);
and U833 (N_833,In_475,In_86);
or U834 (N_834,In_131,In_129);
nand U835 (N_835,In_442,In_430);
nand U836 (N_836,In_273,In_539);
nor U837 (N_837,In_449,In_408);
or U838 (N_838,In_310,In_745);
and U839 (N_839,In_421,In_425);
or U840 (N_840,In_47,In_356);
nand U841 (N_841,In_745,In_718);
nand U842 (N_842,In_691,In_703);
and U843 (N_843,In_111,In_742);
nor U844 (N_844,In_140,In_306);
nor U845 (N_845,In_274,In_588);
nand U846 (N_846,In_56,In_97);
and U847 (N_847,In_379,In_481);
nor U848 (N_848,In_575,In_43);
nand U849 (N_849,In_310,In_114);
and U850 (N_850,In_69,In_672);
nand U851 (N_851,In_587,In_62);
and U852 (N_852,In_260,In_393);
nand U853 (N_853,In_546,In_663);
or U854 (N_854,In_536,In_302);
and U855 (N_855,In_512,In_345);
nor U856 (N_856,In_359,In_746);
nor U857 (N_857,In_411,In_594);
or U858 (N_858,In_385,In_690);
nand U859 (N_859,In_725,In_435);
or U860 (N_860,In_455,In_655);
and U861 (N_861,In_584,In_507);
or U862 (N_862,In_426,In_39);
nand U863 (N_863,In_14,In_301);
nor U864 (N_864,In_573,In_190);
nor U865 (N_865,In_199,In_335);
and U866 (N_866,In_438,In_346);
or U867 (N_867,In_735,In_486);
nor U868 (N_868,In_93,In_422);
or U869 (N_869,In_488,In_130);
nand U870 (N_870,In_188,In_482);
and U871 (N_871,In_720,In_78);
or U872 (N_872,In_28,In_274);
and U873 (N_873,In_250,In_438);
and U874 (N_874,In_120,In_271);
nor U875 (N_875,In_217,In_738);
nand U876 (N_876,In_320,In_675);
and U877 (N_877,In_30,In_468);
or U878 (N_878,In_444,In_551);
or U879 (N_879,In_87,In_187);
nand U880 (N_880,In_633,In_659);
or U881 (N_881,In_173,In_742);
and U882 (N_882,In_401,In_121);
nand U883 (N_883,In_214,In_364);
and U884 (N_884,In_249,In_335);
nor U885 (N_885,In_587,In_100);
or U886 (N_886,In_193,In_81);
and U887 (N_887,In_630,In_244);
and U888 (N_888,In_428,In_692);
nand U889 (N_889,In_612,In_0);
nor U890 (N_890,In_568,In_246);
and U891 (N_891,In_446,In_164);
nand U892 (N_892,In_375,In_507);
or U893 (N_893,In_525,In_18);
xor U894 (N_894,In_349,In_516);
nor U895 (N_895,In_319,In_225);
and U896 (N_896,In_531,In_453);
nand U897 (N_897,In_99,In_368);
nor U898 (N_898,In_143,In_435);
and U899 (N_899,In_344,In_153);
nand U900 (N_900,In_669,In_439);
nand U901 (N_901,In_441,In_412);
and U902 (N_902,In_537,In_246);
or U903 (N_903,In_159,In_287);
or U904 (N_904,In_249,In_674);
nor U905 (N_905,In_75,In_420);
or U906 (N_906,In_203,In_576);
nand U907 (N_907,In_601,In_63);
and U908 (N_908,In_131,In_62);
nand U909 (N_909,In_595,In_456);
nand U910 (N_910,In_54,In_294);
and U911 (N_911,In_238,In_566);
and U912 (N_912,In_153,In_704);
nor U913 (N_913,In_142,In_174);
nand U914 (N_914,In_177,In_470);
and U915 (N_915,In_162,In_613);
or U916 (N_916,In_297,In_294);
nor U917 (N_917,In_552,In_86);
nor U918 (N_918,In_510,In_619);
nor U919 (N_919,In_236,In_239);
or U920 (N_920,In_244,In_655);
and U921 (N_921,In_377,In_717);
and U922 (N_922,In_428,In_267);
nor U923 (N_923,In_457,In_230);
nand U924 (N_924,In_745,In_546);
nand U925 (N_925,In_136,In_15);
nor U926 (N_926,In_420,In_255);
nor U927 (N_927,In_80,In_665);
or U928 (N_928,In_220,In_68);
or U929 (N_929,In_68,In_635);
nor U930 (N_930,In_545,In_547);
nand U931 (N_931,In_581,In_10);
and U932 (N_932,In_130,In_172);
or U933 (N_933,In_229,In_277);
or U934 (N_934,In_569,In_646);
xnor U935 (N_935,In_373,In_661);
nor U936 (N_936,In_633,In_707);
nand U937 (N_937,In_275,In_455);
or U938 (N_938,In_564,In_600);
xnor U939 (N_939,In_509,In_678);
nor U940 (N_940,In_238,In_188);
nor U941 (N_941,In_50,In_620);
and U942 (N_942,In_539,In_378);
nor U943 (N_943,In_728,In_325);
nor U944 (N_944,In_180,In_579);
and U945 (N_945,In_218,In_527);
nor U946 (N_946,In_71,In_521);
nand U947 (N_947,In_163,In_150);
nand U948 (N_948,In_738,In_257);
nor U949 (N_949,In_569,In_351);
or U950 (N_950,In_621,In_713);
nand U951 (N_951,In_9,In_161);
and U952 (N_952,In_21,In_475);
nor U953 (N_953,In_634,In_277);
and U954 (N_954,In_140,In_741);
or U955 (N_955,In_236,In_195);
or U956 (N_956,In_134,In_573);
nand U957 (N_957,In_735,In_169);
or U958 (N_958,In_481,In_212);
nand U959 (N_959,In_227,In_218);
nand U960 (N_960,In_198,In_503);
or U961 (N_961,In_209,In_404);
nand U962 (N_962,In_618,In_236);
and U963 (N_963,In_384,In_297);
and U964 (N_964,In_479,In_39);
and U965 (N_965,In_389,In_467);
nand U966 (N_966,In_161,In_284);
and U967 (N_967,In_4,In_716);
nand U968 (N_968,In_115,In_43);
xnor U969 (N_969,In_16,In_494);
or U970 (N_970,In_579,In_523);
nor U971 (N_971,In_310,In_278);
nor U972 (N_972,In_86,In_639);
or U973 (N_973,In_479,In_34);
and U974 (N_974,In_651,In_244);
nor U975 (N_975,In_168,In_436);
nand U976 (N_976,In_20,In_729);
or U977 (N_977,In_177,In_437);
nand U978 (N_978,In_644,In_282);
or U979 (N_979,In_243,In_318);
nand U980 (N_980,In_689,In_539);
or U981 (N_981,In_192,In_159);
nand U982 (N_982,In_290,In_304);
and U983 (N_983,In_525,In_1);
nand U984 (N_984,In_744,In_132);
nor U985 (N_985,In_539,In_341);
nor U986 (N_986,In_581,In_267);
or U987 (N_987,In_235,In_437);
nor U988 (N_988,In_122,In_556);
and U989 (N_989,In_132,In_701);
and U990 (N_990,In_214,In_156);
or U991 (N_991,In_322,In_98);
nor U992 (N_992,In_617,In_462);
and U993 (N_993,In_106,In_627);
nor U994 (N_994,In_430,In_551);
or U995 (N_995,In_130,In_350);
nand U996 (N_996,In_731,In_429);
or U997 (N_997,In_380,In_582);
nor U998 (N_998,In_32,In_338);
or U999 (N_999,In_415,In_88);
nor U1000 (N_1000,N_383,N_773);
and U1001 (N_1001,N_24,N_781);
nor U1002 (N_1002,N_3,N_654);
nor U1003 (N_1003,N_254,N_125);
nor U1004 (N_1004,N_339,N_474);
and U1005 (N_1005,N_257,N_958);
and U1006 (N_1006,N_107,N_671);
and U1007 (N_1007,N_798,N_522);
or U1008 (N_1008,N_42,N_811);
or U1009 (N_1009,N_963,N_21);
nand U1010 (N_1010,N_552,N_808);
nand U1011 (N_1011,N_580,N_959);
or U1012 (N_1012,N_572,N_47);
nand U1013 (N_1013,N_241,N_78);
nor U1014 (N_1014,N_236,N_22);
nor U1015 (N_1015,N_68,N_11);
and U1016 (N_1016,N_907,N_222);
nor U1017 (N_1017,N_15,N_690);
nand U1018 (N_1018,N_727,N_33);
or U1019 (N_1019,N_457,N_848);
nand U1020 (N_1020,N_469,N_716);
nor U1021 (N_1021,N_590,N_37);
and U1022 (N_1022,N_458,N_7);
or U1023 (N_1023,N_938,N_59);
or U1024 (N_1024,N_542,N_696);
or U1025 (N_1025,N_6,N_679);
and U1026 (N_1026,N_672,N_620);
nor U1027 (N_1027,N_543,N_331);
nor U1028 (N_1028,N_110,N_105);
nand U1029 (N_1029,N_280,N_817);
nor U1030 (N_1030,N_746,N_9);
nand U1031 (N_1031,N_205,N_568);
and U1032 (N_1032,N_533,N_253);
and U1033 (N_1033,N_738,N_956);
nor U1034 (N_1034,N_686,N_816);
or U1035 (N_1035,N_667,N_987);
or U1036 (N_1036,N_459,N_585);
or U1037 (N_1037,N_197,N_677);
nor U1038 (N_1038,N_61,N_111);
nor U1039 (N_1039,N_234,N_424);
nor U1040 (N_1040,N_176,N_614);
and U1041 (N_1041,N_683,N_661);
nor U1042 (N_1042,N_190,N_181);
xnor U1043 (N_1043,N_507,N_855);
and U1044 (N_1044,N_351,N_944);
nor U1045 (N_1045,N_137,N_906);
nand U1046 (N_1046,N_829,N_199);
nand U1047 (N_1047,N_18,N_289);
or U1048 (N_1048,N_266,N_264);
and U1049 (N_1049,N_597,N_286);
and U1050 (N_1050,N_516,N_536);
nand U1051 (N_1051,N_307,N_853);
or U1052 (N_1052,N_731,N_297);
nand U1053 (N_1053,N_885,N_739);
nand U1054 (N_1054,N_612,N_931);
and U1055 (N_1055,N_640,N_606);
nand U1056 (N_1056,N_185,N_36);
xnor U1057 (N_1057,N_503,N_326);
nand U1058 (N_1058,N_991,N_518);
nor U1059 (N_1059,N_616,N_563);
and U1060 (N_1060,N_418,N_615);
nand U1061 (N_1061,N_64,N_208);
nor U1062 (N_1062,N_407,N_428);
or U1063 (N_1063,N_20,N_796);
and U1064 (N_1064,N_415,N_335);
nor U1065 (N_1065,N_734,N_506);
or U1066 (N_1066,N_475,N_421);
nand U1067 (N_1067,N_873,N_934);
and U1068 (N_1068,N_665,N_823);
nand U1069 (N_1069,N_594,N_336);
or U1070 (N_1070,N_344,N_687);
nand U1071 (N_1071,N_652,N_30);
and U1072 (N_1072,N_399,N_322);
nand U1073 (N_1073,N_79,N_557);
nor U1074 (N_1074,N_630,N_911);
nand U1075 (N_1075,N_814,N_549);
or U1076 (N_1076,N_939,N_998);
nand U1077 (N_1077,N_485,N_251);
nand U1078 (N_1078,N_699,N_901);
or U1079 (N_1079,N_281,N_218);
or U1080 (N_1080,N_454,N_278);
or U1081 (N_1081,N_584,N_363);
or U1082 (N_1082,N_747,N_760);
and U1083 (N_1083,N_519,N_427);
or U1084 (N_1084,N_362,N_138);
and U1085 (N_1085,N_910,N_919);
or U1086 (N_1086,N_131,N_388);
and U1087 (N_1087,N_139,N_573);
nor U1088 (N_1088,N_41,N_882);
or U1089 (N_1089,N_118,N_969);
and U1090 (N_1090,N_327,N_170);
nand U1091 (N_1091,N_980,N_409);
or U1092 (N_1092,N_722,N_957);
or U1093 (N_1093,N_318,N_724);
nor U1094 (N_1094,N_601,N_488);
nor U1095 (N_1095,N_210,N_420);
nor U1096 (N_1096,N_26,N_358);
or U1097 (N_1097,N_124,N_688);
and U1098 (N_1098,N_451,N_613);
or U1099 (N_1099,N_864,N_52);
xor U1100 (N_1100,N_617,N_341);
or U1101 (N_1101,N_247,N_789);
xnor U1102 (N_1102,N_35,N_513);
and U1103 (N_1103,N_345,N_762);
or U1104 (N_1104,N_444,N_115);
and U1105 (N_1105,N_728,N_733);
and U1106 (N_1106,N_847,N_877);
or U1107 (N_1107,N_741,N_482);
and U1108 (N_1108,N_876,N_730);
or U1109 (N_1109,N_135,N_430);
nand U1110 (N_1110,N_132,N_763);
or U1111 (N_1111,N_926,N_631);
nand U1112 (N_1112,N_530,N_397);
nand U1113 (N_1113,N_870,N_863);
and U1114 (N_1114,N_250,N_865);
nor U1115 (N_1115,N_279,N_100);
nor U1116 (N_1116,N_647,N_788);
and U1117 (N_1117,N_492,N_570);
nor U1118 (N_1118,N_224,N_213);
nand U1119 (N_1119,N_604,N_403);
nor U1120 (N_1120,N_66,N_146);
nor U1121 (N_1121,N_866,N_802);
and U1122 (N_1122,N_971,N_942);
and U1123 (N_1123,N_676,N_499);
nor U1124 (N_1124,N_94,N_13);
nand U1125 (N_1125,N_862,N_954);
and U1126 (N_1126,N_774,N_902);
or U1127 (N_1127,N_869,N_650);
nand U1128 (N_1128,N_439,N_152);
or U1129 (N_1129,N_517,N_160);
and U1130 (N_1130,N_150,N_525);
nand U1131 (N_1131,N_221,N_288);
or U1132 (N_1132,N_861,N_607);
or U1133 (N_1133,N_524,N_719);
and U1134 (N_1134,N_410,N_621);
nand U1135 (N_1135,N_95,N_768);
and U1136 (N_1136,N_382,N_897);
nand U1137 (N_1137,N_765,N_841);
nand U1138 (N_1138,N_225,N_933);
and U1139 (N_1139,N_282,N_813);
or U1140 (N_1140,N_365,N_843);
and U1141 (N_1141,N_504,N_28);
and U1142 (N_1142,N_592,N_596);
nand U1143 (N_1143,N_541,N_134);
and U1144 (N_1144,N_92,N_554);
nor U1145 (N_1145,N_249,N_858);
and U1146 (N_1146,N_978,N_332);
and U1147 (N_1147,N_779,N_836);
nand U1148 (N_1148,N_638,N_361);
or U1149 (N_1149,N_311,N_308);
and U1150 (N_1150,N_149,N_967);
or U1151 (N_1151,N_357,N_31);
nand U1152 (N_1152,N_992,N_772);
nor U1153 (N_1153,N_745,N_545);
nand U1154 (N_1154,N_29,N_743);
nand U1155 (N_1155,N_86,N_408);
nor U1156 (N_1156,N_759,N_913);
or U1157 (N_1157,N_697,N_941);
and U1158 (N_1158,N_639,N_182);
nor U1159 (N_1159,N_501,N_396);
and U1160 (N_1160,N_562,N_764);
and U1161 (N_1161,N_313,N_411);
and U1162 (N_1162,N_995,N_751);
and U1163 (N_1163,N_434,N_949);
nor U1164 (N_1164,N_229,N_867);
nor U1165 (N_1165,N_72,N_782);
and U1166 (N_1166,N_443,N_809);
nor U1167 (N_1167,N_588,N_512);
and U1168 (N_1168,N_16,N_359);
nand U1169 (N_1169,N_40,N_771);
nand U1170 (N_1170,N_223,N_790);
nor U1171 (N_1171,N_883,N_438);
nand U1172 (N_1172,N_548,N_900);
and U1173 (N_1173,N_46,N_818);
and U1174 (N_1174,N_918,N_255);
nand U1175 (N_1175,N_478,N_104);
and U1176 (N_1176,N_398,N_356);
and U1177 (N_1177,N_414,N_186);
and U1178 (N_1178,N_975,N_277);
or U1179 (N_1179,N_915,N_171);
nor U1180 (N_1180,N_385,N_908);
and U1181 (N_1181,N_239,N_209);
and U1182 (N_1182,N_710,N_845);
or U1183 (N_1183,N_660,N_994);
nand U1184 (N_1184,N_348,N_940);
or U1185 (N_1185,N_756,N_200);
and U1186 (N_1186,N_39,N_860);
nor U1187 (N_1187,N_752,N_532);
nor U1188 (N_1188,N_950,N_304);
nor U1189 (N_1189,N_894,N_214);
nand U1190 (N_1190,N_819,N_168);
and U1191 (N_1191,N_82,N_714);
or U1192 (N_1192,N_58,N_153);
nand U1193 (N_1193,N_502,N_188);
nand U1194 (N_1194,N_232,N_384);
and U1195 (N_1195,N_425,N_825);
nor U1196 (N_1196,N_314,N_509);
or U1197 (N_1197,N_821,N_44);
nor U1198 (N_1198,N_903,N_446);
xor U1199 (N_1199,N_744,N_17);
nor U1200 (N_1200,N_535,N_62);
and U1201 (N_1201,N_970,N_912);
or U1202 (N_1202,N_923,N_932);
nand U1203 (N_1203,N_642,N_355);
nand U1204 (N_1204,N_986,N_67);
nand U1205 (N_1205,N_441,N_997);
nand U1206 (N_1206,N_142,N_662);
nor U1207 (N_1207,N_787,N_284);
or U1208 (N_1208,N_979,N_328);
nor U1209 (N_1209,N_498,N_784);
nor U1210 (N_1210,N_128,N_511);
or U1211 (N_1211,N_936,N_742);
nor U1212 (N_1212,N_569,N_989);
or U1213 (N_1213,N_786,N_755);
xor U1214 (N_1214,N_175,N_810);
or U1215 (N_1215,N_163,N_377);
or U1216 (N_1216,N_822,N_644);
nand U1217 (N_1217,N_292,N_849);
nor U1218 (N_1218,N_27,N_436);
nor U1219 (N_1219,N_837,N_364);
or U1220 (N_1220,N_211,N_645);
or U1221 (N_1221,N_974,N_114);
nand U1222 (N_1222,N_462,N_404);
nor U1223 (N_1223,N_96,N_216);
nand U1224 (N_1224,N_57,N_448);
or U1225 (N_1225,N_129,N_723);
nor U1226 (N_1226,N_528,N_447);
xnor U1227 (N_1227,N_682,N_347);
or U1228 (N_1228,N_627,N_832);
nand U1229 (N_1229,N_663,N_538);
nor U1230 (N_1230,N_985,N_405);
xnor U1231 (N_1231,N_120,N_141);
nor U1232 (N_1232,N_19,N_892);
nand U1233 (N_1233,N_93,N_801);
nand U1234 (N_1234,N_648,N_178);
nor U1235 (N_1235,N_729,N_343);
and U1236 (N_1236,N_38,N_898);
nand U1237 (N_1237,N_889,N_196);
or U1238 (N_1238,N_375,N_487);
nor U1239 (N_1239,N_922,N_283);
nor U1240 (N_1240,N_206,N_905);
nor U1241 (N_1241,N_466,N_157);
or U1242 (N_1242,N_852,N_372);
and U1243 (N_1243,N_928,N_965);
or U1244 (N_1244,N_432,N_393);
or U1245 (N_1245,N_147,N_704);
nand U1246 (N_1246,N_574,N_180);
nand U1247 (N_1247,N_184,N_674);
and U1248 (N_1248,N_490,N_8);
nor U1249 (N_1249,N_593,N_419);
nand U1250 (N_1250,N_203,N_761);
and U1251 (N_1251,N_953,N_287);
and U1252 (N_1252,N_556,N_472);
nor U1253 (N_1253,N_700,N_632);
nor U1254 (N_1254,N_201,N_962);
and U1255 (N_1255,N_60,N_207);
nor U1256 (N_1256,N_269,N_945);
or U1257 (N_1257,N_136,N_740);
nand U1258 (N_1258,N_527,N_769);
nand U1259 (N_1259,N_749,N_732);
and U1260 (N_1260,N_303,N_896);
nor U1261 (N_1261,N_169,N_565);
nor U1262 (N_1262,N_489,N_123);
nor U1263 (N_1263,N_324,N_387);
and U1264 (N_1264,N_685,N_566);
nand U1265 (N_1265,N_582,N_243);
and U1266 (N_1266,N_815,N_140);
and U1267 (N_1267,N_193,N_794);
and U1268 (N_1268,N_930,N_678);
or U1269 (N_1269,N_245,N_56);
or U1270 (N_1270,N_329,N_248);
and U1271 (N_1271,N_812,N_851);
and U1272 (N_1272,N_204,N_274);
or U1273 (N_1273,N_634,N_844);
nor U1274 (N_1274,N_0,N_785);
and U1275 (N_1275,N_982,N_258);
or U1276 (N_1276,N_702,N_996);
nand U1277 (N_1277,N_505,N_468);
and U1278 (N_1278,N_651,N_888);
nor U1279 (N_1279,N_878,N_453);
nand U1280 (N_1280,N_887,N_879);
nor U1281 (N_1281,N_999,N_579);
and U1282 (N_1282,N_256,N_74);
and U1283 (N_1283,N_390,N_680);
and U1284 (N_1284,N_968,N_49);
nor U1285 (N_1285,N_103,N_917);
or U1286 (N_1286,N_725,N_833);
and U1287 (N_1287,N_551,N_155);
nor U1288 (N_1288,N_435,N_976);
nor U1289 (N_1289,N_943,N_412);
nor U1290 (N_1290,N_754,N_797);
xnor U1291 (N_1291,N_602,N_895);
and U1292 (N_1292,N_497,N_559);
or U1293 (N_1293,N_85,N_461);
nor U1294 (N_1294,N_846,N_477);
or U1295 (N_1295,N_291,N_984);
nor U1296 (N_1296,N_575,N_805);
nor U1297 (N_1297,N_881,N_440);
nand U1298 (N_1298,N_544,N_927);
or U1299 (N_1299,N_736,N_159);
and U1300 (N_1300,N_493,N_600);
and U1301 (N_1301,N_70,N_133);
or U1302 (N_1302,N_857,N_87);
and U1303 (N_1303,N_369,N_212);
and U1304 (N_1304,N_55,N_367);
nor U1305 (N_1305,N_293,N_422);
or U1306 (N_1306,N_633,N_433);
nor U1307 (N_1307,N_350,N_770);
and U1308 (N_1308,N_546,N_81);
and U1309 (N_1309,N_299,N_309);
nor U1310 (N_1310,N_321,N_479);
nor U1311 (N_1311,N_301,N_381);
or U1312 (N_1312,N_413,N_323);
and U1313 (N_1313,N_715,N_748);
and U1314 (N_1314,N_317,N_791);
or U1315 (N_1315,N_521,N_981);
and U1316 (N_1316,N_450,N_273);
or U1317 (N_1317,N_792,N_402);
nor U1318 (N_1318,N_767,N_628);
or U1319 (N_1319,N_776,N_5);
and U1320 (N_1320,N_4,N_442);
and U1321 (N_1321,N_587,N_330);
or U1322 (N_1322,N_609,N_240);
nor U1323 (N_1323,N_583,N_990);
or U1324 (N_1324,N_757,N_400);
or U1325 (N_1325,N_655,N_373);
nand U1326 (N_1326,N_455,N_290);
and U1327 (N_1327,N_76,N_603);
nor U1328 (N_1328,N_98,N_198);
nand U1329 (N_1329,N_717,N_599);
or U1330 (N_1330,N_539,N_244);
nand U1331 (N_1331,N_668,N_859);
nand U1332 (N_1332,N_401,N_558);
or U1333 (N_1333,N_578,N_102);
nor U1334 (N_1334,N_871,N_354);
or U1335 (N_1335,N_227,N_820);
or U1336 (N_1336,N_302,N_611);
or U1337 (N_1337,N_673,N_179);
and U1338 (N_1338,N_705,N_483);
nor U1339 (N_1339,N_220,N_342);
nor U1340 (N_1340,N_707,N_54);
and U1341 (N_1341,N_948,N_629);
or U1342 (N_1342,N_955,N_34);
and U1343 (N_1343,N_694,N_276);
and U1344 (N_1344,N_156,N_481);
nand U1345 (N_1345,N_161,N_973);
nand U1346 (N_1346,N_777,N_653);
nand U1347 (N_1347,N_766,N_649);
or U1348 (N_1348,N_25,N_709);
or U1349 (N_1349,N_778,N_718);
nor U1350 (N_1350,N_53,N_657);
and U1351 (N_1351,N_296,N_426);
and U1352 (N_1352,N_352,N_465);
or U1353 (N_1353,N_899,N_547);
nor U1354 (N_1354,N_840,N_228);
nand U1355 (N_1355,N_495,N_456);
and U1356 (N_1356,N_144,N_158);
nor U1357 (N_1357,N_116,N_534);
nor U1358 (N_1358,N_389,N_340);
and U1359 (N_1359,N_90,N_262);
nand U1360 (N_1360,N_564,N_856);
or U1361 (N_1361,N_692,N_924);
and U1362 (N_1362,N_374,N_32);
or U1363 (N_1363,N_550,N_643);
or U1364 (N_1364,N_242,N_246);
nand U1365 (N_1365,N_300,N_476);
or U1366 (N_1366,N_315,N_263);
nor U1367 (N_1367,N_235,N_540);
and U1368 (N_1368,N_467,N_589);
nand U1369 (N_1369,N_50,N_154);
nor U1370 (N_1370,N_946,N_964);
and U1371 (N_1371,N_464,N_577);
and U1372 (N_1372,N_127,N_929);
nand U1373 (N_1373,N_626,N_445);
nor U1374 (N_1374,N_567,N_43);
and U1375 (N_1375,N_598,N_108);
or U1376 (N_1376,N_97,N_463);
nand U1377 (N_1377,N_830,N_394);
and U1378 (N_1378,N_925,N_219);
nand U1379 (N_1379,N_803,N_122);
or U1380 (N_1380,N_799,N_298);
xor U1381 (N_1381,N_555,N_595);
or U1382 (N_1382,N_272,N_75);
or U1383 (N_1383,N_780,N_712);
nand U1384 (N_1384,N_1,N_109);
and U1385 (N_1385,N_491,N_698);
or U1386 (N_1386,N_65,N_71);
or U1387 (N_1387,N_960,N_84);
nor U1388 (N_1388,N_2,N_921);
and U1389 (N_1389,N_916,N_961);
or U1390 (N_1390,N_353,N_429);
or U1391 (N_1391,N_909,N_312);
and U1392 (N_1392,N_252,N_368);
nor U1393 (N_1393,N_431,N_553);
and U1394 (N_1394,N_735,N_187);
nand U1395 (N_1395,N_473,N_51);
nand U1396 (N_1396,N_783,N_316);
and U1397 (N_1397,N_689,N_265);
and U1398 (N_1398,N_711,N_386);
or U1399 (N_1399,N_151,N_376);
nor U1400 (N_1400,N_423,N_636);
or U1401 (N_1401,N_720,N_623);
or U1402 (N_1402,N_793,N_192);
and U1403 (N_1403,N_77,N_360);
or U1404 (N_1404,N_531,N_183);
or U1405 (N_1405,N_189,N_130);
nand U1406 (N_1406,N_664,N_260);
and U1407 (N_1407,N_666,N_804);
or U1408 (N_1408,N_839,N_486);
nor U1409 (N_1409,N_306,N_23);
and U1410 (N_1410,N_172,N_775);
and U1411 (N_1411,N_480,N_177);
or U1412 (N_1412,N_195,N_379);
or U1413 (N_1413,N_691,N_835);
or U1414 (N_1414,N_993,N_148);
nor U1415 (N_1415,N_145,N_523);
nor U1416 (N_1416,N_449,N_670);
or U1417 (N_1417,N_850,N_635);
nor U1418 (N_1418,N_226,N_370);
nor U1419 (N_1419,N_935,N_726);
and U1420 (N_1420,N_294,N_952);
nand U1421 (N_1421,N_618,N_378);
or U1422 (N_1422,N_101,N_333);
or U1423 (N_1423,N_675,N_63);
nand U1424 (N_1424,N_701,N_591);
nand U1425 (N_1425,N_893,N_831);
nor U1426 (N_1426,N_167,N_366);
and U1427 (N_1427,N_417,N_658);
nor U1428 (N_1428,N_261,N_460);
or U1429 (N_1429,N_194,N_121);
nand U1430 (N_1430,N_162,N_69);
and U1431 (N_1431,N_113,N_656);
or U1432 (N_1432,N_164,N_721);
and U1433 (N_1433,N_325,N_703);
and U1434 (N_1434,N_510,N_106);
nor U1435 (N_1435,N_807,N_983);
nor U1436 (N_1436,N_904,N_537);
or U1437 (N_1437,N_624,N_337);
nor U1438 (N_1438,N_320,N_231);
and U1439 (N_1439,N_920,N_143);
nand U1440 (N_1440,N_576,N_619);
or U1441 (N_1441,N_795,N_295);
nor U1442 (N_1442,N_706,N_496);
nor U1443 (N_1443,N_238,N_827);
nand U1444 (N_1444,N_89,N_800);
or U1445 (N_1445,N_268,N_659);
nand U1446 (N_1446,N_608,N_515);
nand U1447 (N_1447,N_868,N_684);
and U1448 (N_1448,N_605,N_230);
and U1449 (N_1449,N_622,N_237);
nand U1450 (N_1450,N_112,N_470);
or U1451 (N_1451,N_452,N_750);
and U1452 (N_1452,N_753,N_437);
xor U1453 (N_1453,N_319,N_951);
nand U1454 (N_1454,N_275,N_334);
and U1455 (N_1455,N_826,N_202);
nand U1456 (N_1456,N_625,N_884);
and U1457 (N_1457,N_416,N_271);
nand U1458 (N_1458,N_270,N_83);
and U1459 (N_1459,N_681,N_708);
nor U1460 (N_1460,N_669,N_126);
nor U1461 (N_1461,N_637,N_641);
and U1462 (N_1462,N_834,N_215);
nand U1463 (N_1463,N_484,N_526);
nor U1464 (N_1464,N_561,N_14);
xnor U1465 (N_1465,N_117,N_174);
nand U1466 (N_1466,N_838,N_166);
nand U1467 (N_1467,N_806,N_842);
nor U1468 (N_1468,N_494,N_285);
or U1469 (N_1469,N_346,N_854);
and U1470 (N_1470,N_165,N_571);
and U1471 (N_1471,N_824,N_12);
or U1472 (N_1472,N_45,N_529);
nor U1473 (N_1473,N_508,N_890);
and U1474 (N_1474,N_310,N_695);
nand U1475 (N_1475,N_217,N_966);
and U1476 (N_1476,N_886,N_874);
or U1477 (N_1477,N_73,N_392);
or U1478 (N_1478,N_80,N_371);
nor U1479 (N_1479,N_99,N_977);
nor U1480 (N_1480,N_520,N_380);
nor U1481 (N_1481,N_471,N_267);
and U1482 (N_1482,N_988,N_581);
nor U1483 (N_1483,N_349,N_500);
nor U1484 (N_1484,N_758,N_88);
and U1485 (N_1485,N_173,N_191);
nor U1486 (N_1486,N_233,N_972);
nor U1487 (N_1487,N_305,N_737);
or U1488 (N_1488,N_338,N_891);
nor U1489 (N_1489,N_914,N_119);
nor U1490 (N_1490,N_872,N_91);
and U1491 (N_1491,N_406,N_395);
nand U1492 (N_1492,N_875,N_828);
or U1493 (N_1493,N_646,N_48);
or U1494 (N_1494,N_259,N_514);
nand U1495 (N_1495,N_586,N_610);
nand U1496 (N_1496,N_10,N_560);
or U1497 (N_1497,N_391,N_947);
and U1498 (N_1498,N_713,N_693);
or U1499 (N_1499,N_880,N_937);
nor U1500 (N_1500,N_201,N_758);
nor U1501 (N_1501,N_927,N_173);
and U1502 (N_1502,N_351,N_787);
or U1503 (N_1503,N_981,N_472);
nand U1504 (N_1504,N_150,N_341);
or U1505 (N_1505,N_211,N_605);
and U1506 (N_1506,N_363,N_637);
nand U1507 (N_1507,N_310,N_433);
or U1508 (N_1508,N_491,N_207);
nand U1509 (N_1509,N_337,N_53);
nand U1510 (N_1510,N_76,N_99);
or U1511 (N_1511,N_857,N_821);
nor U1512 (N_1512,N_676,N_982);
or U1513 (N_1513,N_856,N_58);
nor U1514 (N_1514,N_113,N_819);
nand U1515 (N_1515,N_159,N_187);
nand U1516 (N_1516,N_857,N_212);
and U1517 (N_1517,N_754,N_95);
or U1518 (N_1518,N_153,N_714);
or U1519 (N_1519,N_262,N_933);
or U1520 (N_1520,N_74,N_721);
and U1521 (N_1521,N_415,N_99);
and U1522 (N_1522,N_989,N_638);
or U1523 (N_1523,N_918,N_224);
and U1524 (N_1524,N_908,N_161);
nor U1525 (N_1525,N_144,N_793);
and U1526 (N_1526,N_944,N_179);
and U1527 (N_1527,N_380,N_191);
nand U1528 (N_1528,N_691,N_285);
and U1529 (N_1529,N_608,N_849);
nor U1530 (N_1530,N_36,N_702);
and U1531 (N_1531,N_867,N_323);
or U1532 (N_1532,N_183,N_338);
and U1533 (N_1533,N_476,N_532);
and U1534 (N_1534,N_757,N_911);
and U1535 (N_1535,N_328,N_46);
nand U1536 (N_1536,N_862,N_534);
or U1537 (N_1537,N_558,N_692);
nand U1538 (N_1538,N_673,N_161);
nor U1539 (N_1539,N_887,N_361);
and U1540 (N_1540,N_603,N_903);
or U1541 (N_1541,N_377,N_455);
and U1542 (N_1542,N_183,N_622);
or U1543 (N_1543,N_703,N_714);
or U1544 (N_1544,N_525,N_940);
or U1545 (N_1545,N_882,N_168);
or U1546 (N_1546,N_240,N_378);
or U1547 (N_1547,N_207,N_361);
and U1548 (N_1548,N_112,N_581);
nand U1549 (N_1549,N_20,N_370);
and U1550 (N_1550,N_588,N_131);
and U1551 (N_1551,N_436,N_156);
nand U1552 (N_1552,N_853,N_801);
nand U1553 (N_1553,N_836,N_85);
and U1554 (N_1554,N_583,N_671);
nand U1555 (N_1555,N_49,N_892);
and U1556 (N_1556,N_726,N_813);
nand U1557 (N_1557,N_794,N_110);
or U1558 (N_1558,N_12,N_559);
and U1559 (N_1559,N_722,N_136);
or U1560 (N_1560,N_128,N_468);
nand U1561 (N_1561,N_426,N_777);
nor U1562 (N_1562,N_292,N_271);
nand U1563 (N_1563,N_210,N_292);
nand U1564 (N_1564,N_464,N_274);
and U1565 (N_1565,N_707,N_922);
and U1566 (N_1566,N_674,N_785);
nor U1567 (N_1567,N_491,N_556);
xor U1568 (N_1568,N_230,N_468);
nand U1569 (N_1569,N_277,N_404);
nand U1570 (N_1570,N_553,N_784);
nor U1571 (N_1571,N_211,N_539);
and U1572 (N_1572,N_691,N_728);
nand U1573 (N_1573,N_638,N_350);
nand U1574 (N_1574,N_484,N_602);
nor U1575 (N_1575,N_101,N_600);
nor U1576 (N_1576,N_552,N_891);
and U1577 (N_1577,N_496,N_604);
and U1578 (N_1578,N_336,N_337);
nand U1579 (N_1579,N_170,N_567);
nor U1580 (N_1580,N_302,N_508);
and U1581 (N_1581,N_297,N_641);
or U1582 (N_1582,N_603,N_4);
nor U1583 (N_1583,N_945,N_552);
and U1584 (N_1584,N_846,N_84);
and U1585 (N_1585,N_24,N_147);
and U1586 (N_1586,N_894,N_742);
nor U1587 (N_1587,N_745,N_949);
nor U1588 (N_1588,N_139,N_868);
or U1589 (N_1589,N_834,N_988);
nand U1590 (N_1590,N_763,N_660);
and U1591 (N_1591,N_90,N_957);
or U1592 (N_1592,N_413,N_548);
nor U1593 (N_1593,N_666,N_640);
and U1594 (N_1594,N_592,N_259);
or U1595 (N_1595,N_104,N_562);
or U1596 (N_1596,N_768,N_366);
nand U1597 (N_1597,N_253,N_51);
and U1598 (N_1598,N_328,N_18);
or U1599 (N_1599,N_807,N_804);
nor U1600 (N_1600,N_229,N_923);
or U1601 (N_1601,N_921,N_463);
nor U1602 (N_1602,N_386,N_595);
nand U1603 (N_1603,N_658,N_921);
nor U1604 (N_1604,N_820,N_43);
or U1605 (N_1605,N_467,N_656);
and U1606 (N_1606,N_207,N_521);
and U1607 (N_1607,N_822,N_195);
or U1608 (N_1608,N_312,N_853);
nand U1609 (N_1609,N_531,N_255);
nand U1610 (N_1610,N_181,N_314);
and U1611 (N_1611,N_542,N_258);
nand U1612 (N_1612,N_890,N_847);
or U1613 (N_1613,N_118,N_976);
nor U1614 (N_1614,N_235,N_659);
nor U1615 (N_1615,N_966,N_850);
or U1616 (N_1616,N_991,N_507);
and U1617 (N_1617,N_694,N_523);
nand U1618 (N_1618,N_380,N_409);
nand U1619 (N_1619,N_484,N_597);
nand U1620 (N_1620,N_756,N_875);
nand U1621 (N_1621,N_461,N_609);
nand U1622 (N_1622,N_17,N_594);
and U1623 (N_1623,N_953,N_644);
nor U1624 (N_1624,N_144,N_981);
and U1625 (N_1625,N_840,N_884);
or U1626 (N_1626,N_531,N_916);
nand U1627 (N_1627,N_361,N_565);
and U1628 (N_1628,N_670,N_327);
xnor U1629 (N_1629,N_69,N_120);
nand U1630 (N_1630,N_827,N_764);
and U1631 (N_1631,N_297,N_314);
or U1632 (N_1632,N_522,N_193);
and U1633 (N_1633,N_486,N_235);
nor U1634 (N_1634,N_813,N_380);
nor U1635 (N_1635,N_861,N_243);
nand U1636 (N_1636,N_26,N_61);
nor U1637 (N_1637,N_932,N_236);
and U1638 (N_1638,N_581,N_330);
nor U1639 (N_1639,N_706,N_982);
or U1640 (N_1640,N_353,N_714);
or U1641 (N_1641,N_275,N_955);
nand U1642 (N_1642,N_341,N_69);
nor U1643 (N_1643,N_978,N_368);
nand U1644 (N_1644,N_157,N_357);
or U1645 (N_1645,N_759,N_701);
and U1646 (N_1646,N_708,N_933);
nor U1647 (N_1647,N_332,N_575);
nor U1648 (N_1648,N_985,N_404);
nand U1649 (N_1649,N_151,N_71);
nand U1650 (N_1650,N_227,N_786);
nor U1651 (N_1651,N_433,N_966);
and U1652 (N_1652,N_979,N_467);
and U1653 (N_1653,N_299,N_294);
or U1654 (N_1654,N_145,N_293);
nor U1655 (N_1655,N_122,N_222);
nor U1656 (N_1656,N_131,N_85);
or U1657 (N_1657,N_744,N_313);
and U1658 (N_1658,N_131,N_631);
or U1659 (N_1659,N_743,N_151);
and U1660 (N_1660,N_508,N_836);
nand U1661 (N_1661,N_983,N_339);
nor U1662 (N_1662,N_493,N_145);
or U1663 (N_1663,N_669,N_623);
nand U1664 (N_1664,N_25,N_795);
and U1665 (N_1665,N_527,N_714);
nor U1666 (N_1666,N_87,N_832);
nand U1667 (N_1667,N_185,N_965);
or U1668 (N_1668,N_36,N_321);
or U1669 (N_1669,N_742,N_73);
nand U1670 (N_1670,N_840,N_20);
nand U1671 (N_1671,N_460,N_34);
xor U1672 (N_1672,N_305,N_23);
xnor U1673 (N_1673,N_239,N_68);
or U1674 (N_1674,N_983,N_291);
nor U1675 (N_1675,N_46,N_35);
nand U1676 (N_1676,N_705,N_896);
or U1677 (N_1677,N_713,N_729);
or U1678 (N_1678,N_41,N_664);
and U1679 (N_1679,N_456,N_357);
nor U1680 (N_1680,N_240,N_574);
or U1681 (N_1681,N_355,N_208);
and U1682 (N_1682,N_699,N_442);
nand U1683 (N_1683,N_784,N_12);
and U1684 (N_1684,N_133,N_572);
and U1685 (N_1685,N_293,N_0);
or U1686 (N_1686,N_854,N_751);
nand U1687 (N_1687,N_794,N_236);
or U1688 (N_1688,N_712,N_820);
nand U1689 (N_1689,N_300,N_877);
nand U1690 (N_1690,N_961,N_946);
nor U1691 (N_1691,N_174,N_871);
nor U1692 (N_1692,N_320,N_348);
and U1693 (N_1693,N_506,N_216);
or U1694 (N_1694,N_544,N_773);
and U1695 (N_1695,N_306,N_169);
or U1696 (N_1696,N_494,N_800);
nor U1697 (N_1697,N_96,N_356);
or U1698 (N_1698,N_834,N_198);
or U1699 (N_1699,N_949,N_510);
and U1700 (N_1700,N_992,N_271);
or U1701 (N_1701,N_181,N_676);
or U1702 (N_1702,N_867,N_745);
and U1703 (N_1703,N_143,N_777);
nand U1704 (N_1704,N_640,N_277);
or U1705 (N_1705,N_430,N_14);
nand U1706 (N_1706,N_615,N_362);
and U1707 (N_1707,N_972,N_729);
and U1708 (N_1708,N_296,N_97);
and U1709 (N_1709,N_538,N_551);
nand U1710 (N_1710,N_589,N_136);
and U1711 (N_1711,N_183,N_86);
or U1712 (N_1712,N_24,N_778);
nor U1713 (N_1713,N_787,N_822);
and U1714 (N_1714,N_159,N_687);
nor U1715 (N_1715,N_305,N_456);
and U1716 (N_1716,N_245,N_147);
and U1717 (N_1717,N_518,N_280);
or U1718 (N_1718,N_718,N_607);
and U1719 (N_1719,N_188,N_160);
or U1720 (N_1720,N_269,N_762);
nand U1721 (N_1721,N_433,N_715);
nor U1722 (N_1722,N_374,N_865);
nor U1723 (N_1723,N_386,N_415);
nor U1724 (N_1724,N_270,N_449);
nand U1725 (N_1725,N_780,N_669);
xnor U1726 (N_1726,N_581,N_873);
nor U1727 (N_1727,N_235,N_533);
nand U1728 (N_1728,N_840,N_640);
and U1729 (N_1729,N_684,N_186);
xnor U1730 (N_1730,N_681,N_873);
and U1731 (N_1731,N_188,N_204);
or U1732 (N_1732,N_865,N_300);
and U1733 (N_1733,N_54,N_23);
or U1734 (N_1734,N_165,N_80);
and U1735 (N_1735,N_957,N_964);
and U1736 (N_1736,N_392,N_576);
and U1737 (N_1737,N_825,N_228);
and U1738 (N_1738,N_208,N_724);
nand U1739 (N_1739,N_15,N_541);
nor U1740 (N_1740,N_832,N_421);
nor U1741 (N_1741,N_711,N_323);
nand U1742 (N_1742,N_85,N_444);
nor U1743 (N_1743,N_64,N_651);
nor U1744 (N_1744,N_548,N_777);
nand U1745 (N_1745,N_203,N_439);
or U1746 (N_1746,N_961,N_370);
and U1747 (N_1747,N_836,N_255);
nor U1748 (N_1748,N_209,N_509);
and U1749 (N_1749,N_223,N_759);
and U1750 (N_1750,N_168,N_811);
nor U1751 (N_1751,N_72,N_804);
and U1752 (N_1752,N_253,N_480);
nor U1753 (N_1753,N_808,N_114);
nand U1754 (N_1754,N_291,N_160);
nand U1755 (N_1755,N_325,N_13);
or U1756 (N_1756,N_853,N_547);
nand U1757 (N_1757,N_312,N_193);
nor U1758 (N_1758,N_101,N_908);
nor U1759 (N_1759,N_374,N_574);
nor U1760 (N_1760,N_412,N_75);
nand U1761 (N_1761,N_410,N_9);
or U1762 (N_1762,N_960,N_980);
and U1763 (N_1763,N_860,N_161);
nor U1764 (N_1764,N_468,N_284);
or U1765 (N_1765,N_895,N_986);
nand U1766 (N_1766,N_199,N_759);
nor U1767 (N_1767,N_770,N_390);
or U1768 (N_1768,N_803,N_906);
and U1769 (N_1769,N_299,N_6);
nand U1770 (N_1770,N_776,N_652);
nand U1771 (N_1771,N_58,N_977);
and U1772 (N_1772,N_787,N_778);
nor U1773 (N_1773,N_47,N_984);
and U1774 (N_1774,N_350,N_448);
nand U1775 (N_1775,N_785,N_373);
nand U1776 (N_1776,N_30,N_905);
nor U1777 (N_1777,N_128,N_879);
or U1778 (N_1778,N_552,N_259);
nor U1779 (N_1779,N_453,N_656);
nand U1780 (N_1780,N_120,N_489);
nand U1781 (N_1781,N_622,N_13);
or U1782 (N_1782,N_602,N_985);
nor U1783 (N_1783,N_542,N_487);
nand U1784 (N_1784,N_456,N_145);
nor U1785 (N_1785,N_545,N_926);
nand U1786 (N_1786,N_549,N_111);
nor U1787 (N_1787,N_826,N_78);
and U1788 (N_1788,N_190,N_236);
or U1789 (N_1789,N_392,N_561);
or U1790 (N_1790,N_634,N_735);
nand U1791 (N_1791,N_651,N_368);
nor U1792 (N_1792,N_318,N_424);
or U1793 (N_1793,N_628,N_153);
nand U1794 (N_1794,N_464,N_318);
nor U1795 (N_1795,N_90,N_270);
nand U1796 (N_1796,N_487,N_529);
nand U1797 (N_1797,N_788,N_274);
and U1798 (N_1798,N_867,N_619);
nand U1799 (N_1799,N_454,N_728);
or U1800 (N_1800,N_851,N_871);
or U1801 (N_1801,N_709,N_747);
or U1802 (N_1802,N_444,N_742);
or U1803 (N_1803,N_6,N_960);
and U1804 (N_1804,N_603,N_105);
or U1805 (N_1805,N_799,N_211);
and U1806 (N_1806,N_576,N_202);
or U1807 (N_1807,N_525,N_77);
or U1808 (N_1808,N_912,N_500);
nand U1809 (N_1809,N_303,N_961);
nand U1810 (N_1810,N_908,N_419);
or U1811 (N_1811,N_301,N_116);
or U1812 (N_1812,N_534,N_59);
and U1813 (N_1813,N_210,N_807);
or U1814 (N_1814,N_536,N_930);
nor U1815 (N_1815,N_256,N_687);
and U1816 (N_1816,N_890,N_402);
or U1817 (N_1817,N_573,N_590);
and U1818 (N_1818,N_359,N_171);
nor U1819 (N_1819,N_779,N_845);
nor U1820 (N_1820,N_387,N_990);
and U1821 (N_1821,N_665,N_517);
and U1822 (N_1822,N_100,N_503);
or U1823 (N_1823,N_389,N_3);
nor U1824 (N_1824,N_922,N_916);
and U1825 (N_1825,N_37,N_400);
and U1826 (N_1826,N_19,N_6);
and U1827 (N_1827,N_810,N_324);
nand U1828 (N_1828,N_260,N_796);
or U1829 (N_1829,N_322,N_153);
nor U1830 (N_1830,N_335,N_185);
or U1831 (N_1831,N_540,N_567);
and U1832 (N_1832,N_390,N_486);
nor U1833 (N_1833,N_609,N_595);
nor U1834 (N_1834,N_894,N_78);
nor U1835 (N_1835,N_133,N_306);
nor U1836 (N_1836,N_504,N_86);
or U1837 (N_1837,N_243,N_736);
or U1838 (N_1838,N_530,N_9);
nand U1839 (N_1839,N_996,N_78);
and U1840 (N_1840,N_19,N_635);
nor U1841 (N_1841,N_320,N_10);
nor U1842 (N_1842,N_454,N_358);
nand U1843 (N_1843,N_330,N_817);
nand U1844 (N_1844,N_634,N_229);
or U1845 (N_1845,N_903,N_803);
nor U1846 (N_1846,N_328,N_642);
and U1847 (N_1847,N_454,N_9);
and U1848 (N_1848,N_79,N_421);
nor U1849 (N_1849,N_575,N_275);
nand U1850 (N_1850,N_921,N_408);
or U1851 (N_1851,N_948,N_982);
or U1852 (N_1852,N_359,N_155);
and U1853 (N_1853,N_624,N_625);
and U1854 (N_1854,N_117,N_696);
or U1855 (N_1855,N_325,N_58);
or U1856 (N_1856,N_21,N_558);
nor U1857 (N_1857,N_326,N_140);
or U1858 (N_1858,N_783,N_596);
nor U1859 (N_1859,N_499,N_619);
nor U1860 (N_1860,N_823,N_363);
and U1861 (N_1861,N_629,N_166);
nand U1862 (N_1862,N_748,N_248);
or U1863 (N_1863,N_4,N_304);
or U1864 (N_1864,N_421,N_870);
nand U1865 (N_1865,N_782,N_346);
nand U1866 (N_1866,N_770,N_743);
nand U1867 (N_1867,N_366,N_126);
and U1868 (N_1868,N_447,N_555);
and U1869 (N_1869,N_477,N_324);
nand U1870 (N_1870,N_118,N_269);
and U1871 (N_1871,N_801,N_840);
nand U1872 (N_1872,N_955,N_51);
and U1873 (N_1873,N_457,N_942);
nand U1874 (N_1874,N_384,N_955);
nor U1875 (N_1875,N_4,N_142);
nand U1876 (N_1876,N_121,N_120);
or U1877 (N_1877,N_801,N_550);
nand U1878 (N_1878,N_259,N_777);
and U1879 (N_1879,N_337,N_893);
or U1880 (N_1880,N_797,N_189);
or U1881 (N_1881,N_242,N_949);
and U1882 (N_1882,N_493,N_275);
nor U1883 (N_1883,N_142,N_690);
or U1884 (N_1884,N_483,N_634);
nand U1885 (N_1885,N_827,N_665);
nand U1886 (N_1886,N_192,N_50);
and U1887 (N_1887,N_532,N_106);
nand U1888 (N_1888,N_987,N_195);
nor U1889 (N_1889,N_696,N_738);
nand U1890 (N_1890,N_727,N_328);
and U1891 (N_1891,N_849,N_443);
and U1892 (N_1892,N_656,N_856);
nand U1893 (N_1893,N_9,N_941);
nand U1894 (N_1894,N_658,N_814);
or U1895 (N_1895,N_580,N_237);
nor U1896 (N_1896,N_877,N_49);
or U1897 (N_1897,N_455,N_492);
nor U1898 (N_1898,N_24,N_736);
and U1899 (N_1899,N_978,N_166);
and U1900 (N_1900,N_3,N_96);
and U1901 (N_1901,N_613,N_212);
or U1902 (N_1902,N_106,N_838);
nor U1903 (N_1903,N_920,N_690);
and U1904 (N_1904,N_537,N_745);
and U1905 (N_1905,N_232,N_993);
nand U1906 (N_1906,N_261,N_9);
nand U1907 (N_1907,N_494,N_78);
nand U1908 (N_1908,N_357,N_183);
nor U1909 (N_1909,N_737,N_258);
and U1910 (N_1910,N_450,N_941);
or U1911 (N_1911,N_359,N_642);
nor U1912 (N_1912,N_812,N_988);
nand U1913 (N_1913,N_931,N_621);
nand U1914 (N_1914,N_662,N_558);
nor U1915 (N_1915,N_900,N_328);
nand U1916 (N_1916,N_223,N_620);
nand U1917 (N_1917,N_142,N_841);
or U1918 (N_1918,N_307,N_360);
nor U1919 (N_1919,N_451,N_881);
nor U1920 (N_1920,N_705,N_125);
or U1921 (N_1921,N_335,N_377);
or U1922 (N_1922,N_404,N_160);
nand U1923 (N_1923,N_187,N_768);
and U1924 (N_1924,N_728,N_998);
nand U1925 (N_1925,N_737,N_207);
and U1926 (N_1926,N_70,N_669);
nor U1927 (N_1927,N_350,N_79);
or U1928 (N_1928,N_647,N_806);
or U1929 (N_1929,N_938,N_307);
and U1930 (N_1930,N_829,N_400);
nor U1931 (N_1931,N_451,N_804);
or U1932 (N_1932,N_489,N_571);
nor U1933 (N_1933,N_313,N_312);
xnor U1934 (N_1934,N_884,N_652);
nor U1935 (N_1935,N_466,N_282);
nand U1936 (N_1936,N_75,N_752);
or U1937 (N_1937,N_344,N_479);
nand U1938 (N_1938,N_549,N_931);
and U1939 (N_1939,N_126,N_894);
and U1940 (N_1940,N_694,N_137);
nor U1941 (N_1941,N_435,N_978);
or U1942 (N_1942,N_160,N_57);
and U1943 (N_1943,N_897,N_215);
nor U1944 (N_1944,N_767,N_49);
and U1945 (N_1945,N_508,N_505);
nor U1946 (N_1946,N_638,N_617);
and U1947 (N_1947,N_659,N_564);
xnor U1948 (N_1948,N_151,N_416);
or U1949 (N_1949,N_394,N_75);
or U1950 (N_1950,N_283,N_463);
or U1951 (N_1951,N_584,N_140);
nand U1952 (N_1952,N_469,N_817);
nand U1953 (N_1953,N_642,N_994);
or U1954 (N_1954,N_224,N_706);
and U1955 (N_1955,N_432,N_474);
or U1956 (N_1956,N_645,N_224);
nand U1957 (N_1957,N_559,N_242);
nand U1958 (N_1958,N_441,N_279);
nor U1959 (N_1959,N_974,N_831);
nand U1960 (N_1960,N_129,N_338);
nand U1961 (N_1961,N_224,N_57);
nand U1962 (N_1962,N_356,N_354);
or U1963 (N_1963,N_809,N_405);
nand U1964 (N_1964,N_284,N_594);
nand U1965 (N_1965,N_104,N_974);
and U1966 (N_1966,N_917,N_411);
or U1967 (N_1967,N_919,N_352);
and U1968 (N_1968,N_404,N_702);
or U1969 (N_1969,N_699,N_48);
and U1970 (N_1970,N_614,N_708);
and U1971 (N_1971,N_404,N_619);
nand U1972 (N_1972,N_351,N_815);
or U1973 (N_1973,N_498,N_178);
and U1974 (N_1974,N_520,N_851);
nor U1975 (N_1975,N_796,N_507);
and U1976 (N_1976,N_721,N_420);
and U1977 (N_1977,N_958,N_669);
nand U1978 (N_1978,N_984,N_128);
nand U1979 (N_1979,N_332,N_626);
or U1980 (N_1980,N_104,N_795);
nor U1981 (N_1981,N_527,N_759);
or U1982 (N_1982,N_268,N_547);
nor U1983 (N_1983,N_696,N_962);
nand U1984 (N_1984,N_291,N_712);
and U1985 (N_1985,N_165,N_846);
and U1986 (N_1986,N_365,N_492);
nor U1987 (N_1987,N_466,N_581);
nand U1988 (N_1988,N_96,N_385);
nand U1989 (N_1989,N_365,N_736);
nor U1990 (N_1990,N_313,N_852);
or U1991 (N_1991,N_702,N_585);
and U1992 (N_1992,N_529,N_30);
and U1993 (N_1993,N_233,N_631);
nor U1994 (N_1994,N_167,N_910);
and U1995 (N_1995,N_474,N_741);
and U1996 (N_1996,N_198,N_674);
or U1997 (N_1997,N_618,N_284);
or U1998 (N_1998,N_372,N_725);
nor U1999 (N_1999,N_906,N_313);
nor U2000 (N_2000,N_1051,N_1810);
and U2001 (N_2001,N_1589,N_1876);
or U2002 (N_2002,N_1634,N_1282);
nor U2003 (N_2003,N_1826,N_1885);
and U2004 (N_2004,N_1555,N_1667);
or U2005 (N_2005,N_1846,N_1857);
nand U2006 (N_2006,N_1519,N_1686);
nand U2007 (N_2007,N_1259,N_1475);
nor U2008 (N_2008,N_1099,N_1266);
nand U2009 (N_2009,N_1668,N_1595);
or U2010 (N_2010,N_1756,N_1640);
or U2011 (N_2011,N_1116,N_1448);
and U2012 (N_2012,N_1804,N_1045);
nand U2013 (N_2013,N_1146,N_1186);
nand U2014 (N_2014,N_1687,N_1527);
and U2015 (N_2015,N_1495,N_1500);
nand U2016 (N_2016,N_1506,N_1446);
and U2017 (N_2017,N_1101,N_1866);
and U2018 (N_2018,N_1931,N_1729);
or U2019 (N_2019,N_1755,N_1977);
and U2020 (N_2020,N_1856,N_1759);
nor U2021 (N_2021,N_1894,N_1078);
nor U2022 (N_2022,N_1463,N_1928);
or U2023 (N_2023,N_1158,N_1651);
and U2024 (N_2024,N_1516,N_1210);
and U2025 (N_2025,N_1181,N_1537);
xor U2026 (N_2026,N_1538,N_1498);
nor U2027 (N_2027,N_1434,N_1414);
and U2028 (N_2028,N_1823,N_1194);
nand U2029 (N_2029,N_1901,N_1874);
and U2030 (N_2030,N_1150,N_1298);
or U2031 (N_2031,N_1441,N_1075);
and U2032 (N_2032,N_1166,N_1530);
and U2033 (N_2033,N_1867,N_1945);
and U2034 (N_2034,N_1552,N_1284);
nor U2035 (N_2035,N_1641,N_1923);
or U2036 (N_2036,N_1163,N_1717);
nand U2037 (N_2037,N_1321,N_1239);
or U2038 (N_2038,N_1018,N_1100);
or U2039 (N_2039,N_1649,N_1616);
nor U2040 (N_2040,N_1534,N_1432);
nand U2041 (N_2041,N_1511,N_1997);
or U2042 (N_2042,N_1108,N_1048);
or U2043 (N_2043,N_1365,N_1533);
nor U2044 (N_2044,N_1522,N_1270);
nor U2045 (N_2045,N_1470,N_1111);
nor U2046 (N_2046,N_1016,N_1491);
nand U2047 (N_2047,N_1773,N_1573);
nand U2048 (N_2048,N_1629,N_1788);
and U2049 (N_2049,N_1157,N_1395);
xnor U2050 (N_2050,N_1574,N_1221);
and U2051 (N_2051,N_1676,N_1057);
nor U2052 (N_2052,N_1747,N_1501);
or U2053 (N_2053,N_1135,N_1251);
or U2054 (N_2054,N_1912,N_1103);
and U2055 (N_2055,N_1179,N_1208);
nand U2056 (N_2056,N_1424,N_1827);
nor U2057 (N_2057,N_1204,N_1480);
or U2058 (N_2058,N_1647,N_1658);
nand U2059 (N_2059,N_1828,N_1681);
and U2060 (N_2060,N_1152,N_1155);
and U2061 (N_2061,N_1785,N_1577);
nand U2062 (N_2062,N_1122,N_1611);
nand U2063 (N_2063,N_1899,N_1026);
and U2064 (N_2064,N_1496,N_1292);
nor U2065 (N_2065,N_1043,N_1585);
or U2066 (N_2066,N_1308,N_1198);
nand U2067 (N_2067,N_1570,N_1864);
and U2068 (N_2068,N_1303,N_1503);
nand U2069 (N_2069,N_1737,N_1098);
and U2070 (N_2070,N_1701,N_1921);
nand U2071 (N_2071,N_1515,N_1934);
nor U2072 (N_2072,N_1213,N_1887);
or U2073 (N_2073,N_1401,N_1932);
nand U2074 (N_2074,N_1345,N_1721);
nor U2075 (N_2075,N_1294,N_1529);
nand U2076 (N_2076,N_1030,N_1169);
nand U2077 (N_2077,N_1201,N_1052);
nor U2078 (N_2078,N_1964,N_1246);
nor U2079 (N_2079,N_1691,N_1300);
nand U2080 (N_2080,N_1224,N_1015);
or U2081 (N_2081,N_1286,N_1021);
nand U2082 (N_2082,N_1644,N_1685);
and U2083 (N_2083,N_1722,N_1268);
and U2084 (N_2084,N_1514,N_1006);
nand U2085 (N_2085,N_1718,N_1258);
nor U2086 (N_2086,N_1064,N_1073);
nand U2087 (N_2087,N_1630,N_1397);
nor U2088 (N_2088,N_1865,N_1407);
and U2089 (N_2089,N_1130,N_1709);
or U2090 (N_2090,N_1188,N_1202);
or U2091 (N_2091,N_1940,N_1764);
and U2092 (N_2092,N_1507,N_1614);
xnor U2093 (N_2093,N_1843,N_1364);
or U2094 (N_2094,N_1551,N_1013);
or U2095 (N_2095,N_1907,N_1148);
nor U2096 (N_2096,N_1657,N_1915);
nand U2097 (N_2097,N_1707,N_1133);
nor U2098 (N_2098,N_1623,N_1217);
nor U2099 (N_2099,N_1334,N_1588);
nand U2100 (N_2100,N_1765,N_1746);
nor U2101 (N_2101,N_1858,N_1047);
nand U2102 (N_2102,N_1770,N_1390);
nand U2103 (N_2103,N_1139,N_1184);
or U2104 (N_2104,N_1170,N_1162);
or U2105 (N_2105,N_1502,N_1235);
nand U2106 (N_2106,N_1732,N_1461);
or U2107 (N_2107,N_1484,N_1083);
or U2108 (N_2108,N_1063,N_1466);
xor U2109 (N_2109,N_1325,N_1009);
nor U2110 (N_2110,N_1489,N_1674);
or U2111 (N_2111,N_1338,N_1068);
nand U2112 (N_2112,N_1607,N_1118);
or U2113 (N_2113,N_1102,N_1256);
nand U2114 (N_2114,N_1924,N_1145);
or U2115 (N_2115,N_1656,N_1022);
nand U2116 (N_2116,N_1766,N_1975);
or U2117 (N_2117,N_1689,N_1771);
nand U2118 (N_2118,N_1886,N_1632);
or U2119 (N_2119,N_1842,N_1479);
and U2120 (N_2120,N_1835,N_1058);
nand U2121 (N_2121,N_1206,N_1743);
nand U2122 (N_2122,N_1911,N_1159);
or U2123 (N_2123,N_1378,N_1851);
nor U2124 (N_2124,N_1214,N_1565);
and U2125 (N_2125,N_1177,N_1933);
or U2126 (N_2126,N_1387,N_1309);
nand U2127 (N_2127,N_1703,N_1175);
and U2128 (N_2128,N_1592,N_1394);
or U2129 (N_2129,N_1539,N_1796);
nand U2130 (N_2130,N_1591,N_1829);
nor U2131 (N_2131,N_1947,N_1076);
nor U2132 (N_2132,N_1279,N_1343);
nand U2133 (N_2133,N_1178,N_1392);
and U2134 (N_2134,N_1643,N_1723);
or U2135 (N_2135,N_1207,N_1580);
nand U2136 (N_2136,N_1458,N_1922);
nand U2137 (N_2137,N_1767,N_1220);
and U2138 (N_2138,N_1091,N_1606);
nor U2139 (N_2139,N_1447,N_1289);
and U2140 (N_2140,N_1748,N_1322);
and U2141 (N_2141,N_1879,N_1031);
nor U2142 (N_2142,N_1330,N_1077);
and U2143 (N_2143,N_1939,N_1242);
and U2144 (N_2144,N_1187,N_1627);
or U2145 (N_2145,N_1594,N_1705);
and U2146 (N_2146,N_1085,N_1994);
nor U2147 (N_2147,N_1902,N_1818);
nand U2148 (N_2148,N_1859,N_1191);
and U2149 (N_2149,N_1961,N_1136);
nor U2150 (N_2150,N_1344,N_1001);
or U2151 (N_2151,N_1472,N_1340);
or U2152 (N_2152,N_1750,N_1895);
and U2153 (N_2153,N_1457,N_1348);
or U2154 (N_2154,N_1598,N_1602);
nand U2155 (N_2155,N_1973,N_1149);
nand U2156 (N_2156,N_1557,N_1793);
nor U2157 (N_2157,N_1854,N_1084);
nand U2158 (N_2158,N_1596,N_1693);
and U2159 (N_2159,N_1549,N_1688);
nand U2160 (N_2160,N_1897,N_1942);
or U2161 (N_2161,N_1209,N_1014);
or U2162 (N_2162,N_1850,N_1413);
or U2163 (N_2163,N_1304,N_1482);
nand U2164 (N_2164,N_1107,N_1059);
nor U2165 (N_2165,N_1054,N_1636);
or U2166 (N_2166,N_1996,N_1508);
nor U2167 (N_2167,N_1036,N_1544);
nor U2168 (N_2168,N_1254,N_1028);
or U2169 (N_2169,N_1978,N_1128);
nand U2170 (N_2170,N_1852,N_1760);
nor U2171 (N_2171,N_1231,N_1740);
or U2172 (N_2172,N_1582,N_1357);
or U2173 (N_2173,N_1613,N_1359);
nor U2174 (N_2174,N_1749,N_1391);
nor U2175 (N_2175,N_1679,N_1488);
nor U2176 (N_2176,N_1728,N_1665);
and U2177 (N_2177,N_1069,N_1467);
and U2178 (N_2178,N_1991,N_1797);
or U2179 (N_2179,N_1444,N_1301);
nand U2180 (N_2180,N_1427,N_1393);
xor U2181 (N_2181,N_1443,N_1267);
nor U2182 (N_2182,N_1056,N_1790);
or U2183 (N_2183,N_1180,N_1757);
and U2184 (N_2184,N_1848,N_1377);
or U2185 (N_2185,N_1238,N_1985);
nor U2186 (N_2186,N_1541,N_1801);
or U2187 (N_2187,N_1237,N_1984);
nor U2188 (N_2188,N_1074,N_1786);
or U2189 (N_2189,N_1405,N_1954);
nand U2190 (N_2190,N_1117,N_1873);
nor U2191 (N_2191,N_1123,N_1370);
or U2192 (N_2192,N_1219,N_1455);
nor U2193 (N_2193,N_1981,N_1174);
or U2194 (N_2194,N_1477,N_1090);
nand U2195 (N_2195,N_1240,N_1497);
or U2196 (N_2196,N_1037,N_1442);
nand U2197 (N_2197,N_1412,N_1937);
nor U2198 (N_2198,N_1868,N_1271);
nand U2199 (N_2199,N_1185,N_1664);
and U2200 (N_2200,N_1811,N_1039);
nand U2201 (N_2201,N_1715,N_1941);
nand U2202 (N_2202,N_1971,N_1892);
nor U2203 (N_2203,N_1670,N_1350);
and U2204 (N_2204,N_1232,N_1426);
nand U2205 (N_2205,N_1366,N_1548);
nand U2206 (N_2206,N_1654,N_1568);
or U2207 (N_2207,N_1200,N_1165);
or U2208 (N_2208,N_1635,N_1144);
nor U2209 (N_2209,N_1540,N_1904);
or U2210 (N_2210,N_1459,N_1983);
or U2211 (N_2211,N_1418,N_1281);
or U2212 (N_2212,N_1542,N_1355);
or U2213 (N_2213,N_1019,N_1545);
nand U2214 (N_2214,N_1411,N_1735);
nor U2215 (N_2215,N_1269,N_1840);
or U2216 (N_2216,N_1361,N_1326);
or U2217 (N_2217,N_1253,N_1381);
nor U2218 (N_2218,N_1203,N_1678);
nor U2219 (N_2219,N_1010,N_1314);
and U2220 (N_2220,N_1341,N_1716);
and U2221 (N_2221,N_1929,N_1347);
nor U2222 (N_2222,N_1936,N_1410);
nor U2223 (N_2223,N_1280,N_1215);
and U2224 (N_2224,N_1306,N_1035);
nand U2225 (N_2225,N_1926,N_1097);
nor U2226 (N_2226,N_1862,N_1317);
nor U2227 (N_2227,N_1608,N_1105);
nand U2228 (N_2228,N_1638,N_1734);
or U2229 (N_2229,N_1822,N_1673);
or U2230 (N_2230,N_1171,N_1011);
nor U2231 (N_2231,N_1379,N_1569);
or U2232 (N_2232,N_1262,N_1680);
or U2233 (N_2233,N_1875,N_1336);
or U2234 (N_2234,N_1421,N_1216);
or U2235 (N_2235,N_1814,N_1986);
nand U2236 (N_2236,N_1369,N_1917);
and U2237 (N_2237,N_1012,N_1137);
nand U2238 (N_2238,N_1968,N_1966);
and U2239 (N_2239,N_1134,N_1621);
nor U2240 (N_2240,N_1250,N_1744);
and U2241 (N_2241,N_1683,N_1830);
or U2242 (N_2242,N_1662,N_1324);
nand U2243 (N_2243,N_1249,N_1261);
nor U2244 (N_2244,N_1147,N_1566);
and U2245 (N_2245,N_1910,N_1383);
or U2246 (N_2246,N_1331,N_1433);
or U2247 (N_2247,N_1727,N_1535);
or U2248 (N_2248,N_1310,N_1699);
nor U2249 (N_2249,N_1724,N_1197);
and U2250 (N_2250,N_1095,N_1730);
or U2251 (N_2251,N_1478,N_1774);
nand U2252 (N_2252,N_1252,N_1575);
and U2253 (N_2253,N_1863,N_1979);
and U2254 (N_2254,N_1999,N_1692);
nor U2255 (N_2255,N_1299,N_1311);
or U2256 (N_2256,N_1233,N_1581);
nor U2257 (N_2257,N_1297,N_1655);
nand U2258 (N_2258,N_1944,N_1504);
nand U2259 (N_2259,N_1532,N_1802);
or U2260 (N_2260,N_1599,N_1474);
nand U2261 (N_2261,N_1229,N_1871);
or U2262 (N_2262,N_1510,N_1243);
or U2263 (N_2263,N_1946,N_1618);
and U2264 (N_2264,N_1493,N_1275);
nand U2265 (N_2265,N_1189,N_1520);
nand U2266 (N_2266,N_1769,N_1451);
or U2267 (N_2267,N_1113,N_1002);
and U2268 (N_2268,N_1485,N_1562);
and U2269 (N_2269,N_1440,N_1499);
or U2270 (N_2270,N_1168,N_1800);
or U2271 (N_2271,N_1260,N_1088);
nor U2272 (N_2272,N_1104,N_1962);
or U2273 (N_2273,N_1367,N_1612);
or U2274 (N_2274,N_1572,N_1024);
nor U2275 (N_2275,N_1878,N_1263);
nor U2276 (N_2276,N_1791,N_1845);
nand U2277 (N_2277,N_1758,N_1682);
nor U2278 (N_2278,N_1353,N_1639);
or U2279 (N_2279,N_1245,N_1898);
or U2280 (N_2280,N_1645,N_1909);
nor U2281 (N_2281,N_1454,N_1005);
xnor U2282 (N_2282,N_1720,N_1141);
or U2283 (N_2283,N_1888,N_1761);
nand U2284 (N_2284,N_1388,N_1777);
or U2285 (N_2285,N_1425,N_1704);
nor U2286 (N_2286,N_1559,N_1951);
or U2287 (N_2287,N_1935,N_1960);
and U2288 (N_2288,N_1402,N_1833);
and U2289 (N_2289,N_1053,N_1409);
nand U2290 (N_2290,N_1416,N_1093);
and U2291 (N_2291,N_1349,N_1337);
nand U2292 (N_2292,N_1631,N_1576);
nor U2293 (N_2293,N_1481,N_1193);
nor U2294 (N_2294,N_1697,N_1109);
nand U2295 (N_2295,N_1041,N_1046);
and U2296 (N_2296,N_1956,N_1661);
and U2297 (N_2297,N_1452,N_1615);
or U2298 (N_2298,N_1372,N_1399);
nand U2299 (N_2299,N_1832,N_1998);
nand U2300 (N_2300,N_1558,N_1380);
or U2301 (N_2301,N_1505,N_1164);
nor U2302 (N_2302,N_1603,N_1694);
nand U2303 (N_2303,N_1140,N_1523);
or U2304 (N_2304,N_1625,N_1988);
nor U2305 (N_2305,N_1597,N_1070);
and U2306 (N_2306,N_1020,N_1494);
nor U2307 (N_2307,N_1072,N_1420);
nand U2308 (N_2308,N_1354,N_1247);
and U2309 (N_2309,N_1087,N_1736);
nor U2310 (N_2310,N_1738,N_1439);
nor U2311 (N_2311,N_1719,N_1438);
and U2312 (N_2312,N_1445,N_1619);
nor U2313 (N_2313,N_1652,N_1419);
or U2314 (N_2314,N_1669,N_1806);
nor U2315 (N_2315,N_1908,N_1449);
and U2316 (N_2316,N_1821,N_1787);
nor U2317 (N_2317,N_1029,N_1700);
or U2318 (N_2318,N_1244,N_1483);
or U2319 (N_2319,N_1007,N_1992);
or U2320 (N_2320,N_1436,N_1872);
nor U2321 (N_2321,N_1406,N_1891);
and U2322 (N_2322,N_1115,N_1172);
or U2323 (N_2323,N_1546,N_1125);
nand U2324 (N_2324,N_1027,N_1958);
nor U2325 (N_2325,N_1847,N_1733);
nand U2326 (N_2326,N_1154,N_1663);
and U2327 (N_2327,N_1695,N_1339);
nor U2328 (N_2328,N_1450,N_1653);
and U2329 (N_2329,N_1905,N_1008);
and U2330 (N_2330,N_1831,N_1536);
and U2331 (N_2331,N_1745,N_1696);
or U2332 (N_2332,N_1079,N_1437);
or U2333 (N_2333,N_1110,N_1609);
and U2334 (N_2334,N_1342,N_1295);
nor U2335 (N_2335,N_1291,N_1817);
or U2336 (N_2336,N_1763,N_1086);
nor U2337 (N_2337,N_1429,N_1792);
xor U2338 (N_2338,N_1023,N_1274);
or U2339 (N_2339,N_1230,N_1624);
nand U2340 (N_2340,N_1222,N_1335);
nor U2341 (N_2341,N_1741,N_1080);
or U2342 (N_2342,N_1313,N_1302);
and U2343 (N_2343,N_1468,N_1976);
nor U2344 (N_2344,N_1553,N_1363);
nor U2345 (N_2345,N_1151,N_1990);
nand U2346 (N_2346,N_1593,N_1803);
or U2347 (N_2347,N_1605,N_1784);
or U2348 (N_2348,N_1586,N_1969);
nor U2349 (N_2349,N_1509,N_1358);
and U2350 (N_2350,N_1285,N_1841);
and U2351 (N_2351,N_1967,N_1453);
nor U2352 (N_2352,N_1199,N_1706);
nand U2353 (N_2353,N_1889,N_1880);
and U2354 (N_2354,N_1916,N_1430);
and U2355 (N_2355,N_1671,N_1556);
or U2356 (N_2356,N_1089,N_1067);
and U2357 (N_2357,N_1659,N_1526);
and U2358 (N_2358,N_1849,N_1726);
and U2359 (N_2359,N_1752,N_1277);
and U2360 (N_2360,N_1400,N_1081);
nand U2361 (N_2361,N_1754,N_1000);
or U2362 (N_2362,N_1328,N_1914);
nor U2363 (N_2363,N_1352,N_1211);
or U2364 (N_2364,N_1512,N_1838);
nor U2365 (N_2365,N_1290,N_1315);
nor U2366 (N_2366,N_1517,N_1617);
nand U2367 (N_2367,N_1781,N_1604);
or U2368 (N_2368,N_1183,N_1861);
and U2369 (N_2369,N_1628,N_1778);
nand U2370 (N_2370,N_1799,N_1869);
nor U2371 (N_2371,N_1808,N_1476);
nand U2372 (N_2372,N_1124,N_1877);
and U2373 (N_2373,N_1906,N_1316);
nand U2374 (N_2374,N_1368,N_1900);
nand U2375 (N_2375,N_1273,N_1789);
and U2376 (N_2376,N_1226,N_1257);
nand U2377 (N_2377,N_1710,N_1825);
or U2378 (N_2378,N_1798,N_1223);
nor U2379 (N_2379,N_1296,N_1712);
nand U2380 (N_2380,N_1396,N_1196);
or U2381 (N_2381,N_1373,N_1600);
and U2382 (N_2382,N_1106,N_1783);
and U2383 (N_2383,N_1742,N_1650);
or U2384 (N_2384,N_1356,N_1044);
and U2385 (N_2385,N_1528,N_1132);
and U2386 (N_2386,N_1092,N_1903);
or U2387 (N_2387,N_1236,N_1038);
and U2388 (N_2388,N_1953,N_1884);
nor U2389 (N_2389,N_1004,N_1610);
nand U2390 (N_2390,N_1398,N_1839);
nor U2391 (N_2391,N_1795,N_1672);
nand U2392 (N_2392,N_1970,N_1531);
or U2393 (N_2393,N_1153,N_1061);
nand U2394 (N_2394,N_1836,N_1571);
nand U2395 (N_2395,N_1648,N_1173);
nand U2396 (N_2396,N_1431,N_1417);
nand U2397 (N_2397,N_1702,N_1469);
and U2398 (N_2398,N_1456,N_1927);
nor U2399 (N_2399,N_1307,N_1711);
and U2400 (N_2400,N_1982,N_1049);
and U2401 (N_2401,N_1374,N_1234);
nor U2402 (N_2402,N_1415,N_1312);
nand U2403 (N_2403,N_1385,N_1739);
nor U2404 (N_2404,N_1882,N_1042);
nor U2405 (N_2405,N_1351,N_1096);
nand U2406 (N_2406,N_1460,N_1805);
nor U2407 (N_2407,N_1003,N_1815);
nand U2408 (N_2408,N_1666,N_1794);
and U2409 (N_2409,N_1143,N_1779);
nand U2410 (N_2410,N_1813,N_1032);
or U2411 (N_2411,N_1065,N_1423);
nor U2412 (N_2412,N_1950,N_1190);
and U2413 (N_2413,N_1930,N_1870);
nor U2414 (N_2414,N_1131,N_1142);
and U2415 (N_2415,N_1384,N_1428);
or U2416 (N_2416,N_1112,N_1816);
and U2417 (N_2417,N_1563,N_1225);
and U2418 (N_2418,N_1464,N_1050);
or U2419 (N_2419,N_1974,N_1462);
nand U2420 (N_2420,N_1082,N_1126);
or U2421 (N_2421,N_1218,N_1473);
xnor U2422 (N_2422,N_1195,N_1435);
and U2423 (N_2423,N_1637,N_1287);
and U2424 (N_2424,N_1775,N_1952);
nand U2425 (N_2425,N_1919,N_1033);
nor U2426 (N_2426,N_1318,N_1993);
nand U2427 (N_2427,N_1060,N_1066);
and U2428 (N_2428,N_1062,N_1772);
nand U2429 (N_2429,N_1893,N_1276);
or U2430 (N_2430,N_1731,N_1319);
nand U2431 (N_2431,N_1837,N_1642);
and U2432 (N_2432,N_1896,N_1255);
nor U2433 (N_2433,N_1389,N_1809);
or U2434 (N_2434,N_1492,N_1853);
or U2435 (N_2435,N_1776,N_1288);
or U2436 (N_2436,N_1708,N_1513);
nand U2437 (N_2437,N_1040,N_1965);
or U2438 (N_2438,N_1957,N_1583);
nor U2439 (N_2439,N_1989,N_1332);
and U2440 (N_2440,N_1228,N_1995);
or U2441 (N_2441,N_1881,N_1360);
nor U2442 (N_2442,N_1943,N_1860);
nor U2443 (N_2443,N_1713,N_1844);
or U2444 (N_2444,N_1980,N_1182);
nor U2445 (N_2445,N_1622,N_1584);
or U2446 (N_2446,N_1329,N_1205);
nand U2447 (N_2447,N_1465,N_1959);
and U2448 (N_2448,N_1264,N_1626);
or U2449 (N_2449,N_1684,N_1633);
and U2450 (N_2450,N_1855,N_1820);
or U2451 (N_2451,N_1547,N_1471);
nand U2452 (N_2452,N_1768,N_1987);
nor U2453 (N_2453,N_1554,N_1212);
or U2454 (N_2454,N_1578,N_1293);
nor U2455 (N_2455,N_1807,N_1017);
nand U2456 (N_2456,N_1375,N_1386);
or U2457 (N_2457,N_1127,N_1120);
nor U2458 (N_2458,N_1883,N_1119);
nand U2459 (N_2459,N_1955,N_1620);
and U2460 (N_2460,N_1422,N_1346);
nand U2461 (N_2461,N_1949,N_1371);
and U2462 (N_2462,N_1920,N_1579);
or U2463 (N_2463,N_1819,N_1590);
or U2464 (N_2464,N_1780,N_1241);
and U2465 (N_2465,N_1138,N_1521);
nor U2466 (N_2466,N_1675,N_1824);
or U2467 (N_2467,N_1561,N_1834);
nor U2468 (N_2468,N_1490,N_1913);
or U2469 (N_2469,N_1963,N_1751);
nor U2470 (N_2470,N_1567,N_1972);
nor U2471 (N_2471,N_1725,N_1278);
or U2472 (N_2472,N_1265,N_1025);
nand U2473 (N_2473,N_1550,N_1129);
or U2474 (N_2474,N_1918,N_1156);
or U2475 (N_2475,N_1524,N_1034);
nand U2476 (N_2476,N_1320,N_1646);
xor U2477 (N_2477,N_1925,N_1121);
nand U2478 (N_2478,N_1690,N_1248);
and U2479 (N_2479,N_1055,N_1938);
nand U2480 (N_2480,N_1890,N_1192);
xor U2481 (N_2481,N_1408,N_1071);
or U2482 (N_2482,N_1404,N_1714);
nand U2483 (N_2483,N_1362,N_1094);
and U2484 (N_2484,N_1376,N_1167);
or U2485 (N_2485,N_1305,N_1948);
and U2486 (N_2486,N_1753,N_1161);
nand U2487 (N_2487,N_1812,N_1698);
or U2488 (N_2488,N_1518,N_1176);
and U2489 (N_2489,N_1587,N_1227);
nor U2490 (N_2490,N_1543,N_1160);
nor U2491 (N_2491,N_1560,N_1601);
nor U2492 (N_2492,N_1782,N_1762);
and U2493 (N_2493,N_1403,N_1487);
nor U2494 (N_2494,N_1272,N_1382);
nand U2495 (N_2495,N_1660,N_1677);
nor U2496 (N_2496,N_1327,N_1525);
or U2497 (N_2497,N_1486,N_1333);
or U2498 (N_2498,N_1564,N_1323);
nor U2499 (N_2499,N_1114,N_1283);
nand U2500 (N_2500,N_1989,N_1959);
or U2501 (N_2501,N_1614,N_1616);
nor U2502 (N_2502,N_1211,N_1408);
nand U2503 (N_2503,N_1173,N_1146);
and U2504 (N_2504,N_1622,N_1631);
nand U2505 (N_2505,N_1691,N_1379);
or U2506 (N_2506,N_1197,N_1622);
and U2507 (N_2507,N_1024,N_1239);
and U2508 (N_2508,N_1643,N_1429);
nor U2509 (N_2509,N_1004,N_1094);
and U2510 (N_2510,N_1809,N_1781);
and U2511 (N_2511,N_1323,N_1400);
nand U2512 (N_2512,N_1342,N_1556);
and U2513 (N_2513,N_1018,N_1349);
and U2514 (N_2514,N_1235,N_1879);
or U2515 (N_2515,N_1680,N_1699);
nand U2516 (N_2516,N_1827,N_1571);
nor U2517 (N_2517,N_1380,N_1967);
or U2518 (N_2518,N_1270,N_1443);
nand U2519 (N_2519,N_1184,N_1783);
nand U2520 (N_2520,N_1188,N_1893);
nor U2521 (N_2521,N_1840,N_1602);
and U2522 (N_2522,N_1234,N_1861);
or U2523 (N_2523,N_1335,N_1813);
and U2524 (N_2524,N_1056,N_1678);
and U2525 (N_2525,N_1637,N_1996);
or U2526 (N_2526,N_1252,N_1641);
and U2527 (N_2527,N_1130,N_1600);
nand U2528 (N_2528,N_1758,N_1300);
nand U2529 (N_2529,N_1170,N_1115);
nor U2530 (N_2530,N_1227,N_1179);
nand U2531 (N_2531,N_1066,N_1394);
nand U2532 (N_2532,N_1677,N_1156);
and U2533 (N_2533,N_1341,N_1080);
nand U2534 (N_2534,N_1842,N_1247);
and U2535 (N_2535,N_1097,N_1406);
or U2536 (N_2536,N_1965,N_1717);
or U2537 (N_2537,N_1864,N_1712);
or U2538 (N_2538,N_1957,N_1641);
nor U2539 (N_2539,N_1951,N_1030);
nor U2540 (N_2540,N_1738,N_1301);
or U2541 (N_2541,N_1800,N_1532);
nor U2542 (N_2542,N_1727,N_1042);
and U2543 (N_2543,N_1497,N_1646);
nor U2544 (N_2544,N_1512,N_1998);
and U2545 (N_2545,N_1286,N_1906);
or U2546 (N_2546,N_1317,N_1942);
nand U2547 (N_2547,N_1167,N_1633);
and U2548 (N_2548,N_1749,N_1078);
or U2549 (N_2549,N_1313,N_1062);
nand U2550 (N_2550,N_1503,N_1866);
or U2551 (N_2551,N_1794,N_1081);
or U2552 (N_2552,N_1265,N_1678);
nand U2553 (N_2553,N_1468,N_1330);
nor U2554 (N_2554,N_1014,N_1020);
or U2555 (N_2555,N_1109,N_1645);
nor U2556 (N_2556,N_1063,N_1972);
or U2557 (N_2557,N_1230,N_1350);
nor U2558 (N_2558,N_1886,N_1821);
or U2559 (N_2559,N_1305,N_1403);
nor U2560 (N_2560,N_1873,N_1298);
and U2561 (N_2561,N_1834,N_1723);
nor U2562 (N_2562,N_1135,N_1539);
and U2563 (N_2563,N_1987,N_1709);
nand U2564 (N_2564,N_1880,N_1062);
nor U2565 (N_2565,N_1939,N_1772);
and U2566 (N_2566,N_1126,N_1694);
nor U2567 (N_2567,N_1377,N_1209);
or U2568 (N_2568,N_1764,N_1346);
nor U2569 (N_2569,N_1290,N_1143);
and U2570 (N_2570,N_1860,N_1826);
and U2571 (N_2571,N_1789,N_1064);
and U2572 (N_2572,N_1124,N_1908);
or U2573 (N_2573,N_1550,N_1225);
nor U2574 (N_2574,N_1046,N_1030);
nor U2575 (N_2575,N_1112,N_1081);
xnor U2576 (N_2576,N_1209,N_1198);
nor U2577 (N_2577,N_1779,N_1743);
and U2578 (N_2578,N_1064,N_1947);
or U2579 (N_2579,N_1724,N_1247);
nand U2580 (N_2580,N_1573,N_1984);
nand U2581 (N_2581,N_1823,N_1286);
and U2582 (N_2582,N_1726,N_1222);
nand U2583 (N_2583,N_1301,N_1056);
or U2584 (N_2584,N_1939,N_1846);
nand U2585 (N_2585,N_1032,N_1278);
nand U2586 (N_2586,N_1103,N_1512);
nand U2587 (N_2587,N_1988,N_1576);
nor U2588 (N_2588,N_1148,N_1484);
nor U2589 (N_2589,N_1234,N_1907);
or U2590 (N_2590,N_1193,N_1338);
nand U2591 (N_2591,N_1849,N_1488);
nor U2592 (N_2592,N_1893,N_1086);
nand U2593 (N_2593,N_1532,N_1746);
or U2594 (N_2594,N_1818,N_1109);
nor U2595 (N_2595,N_1027,N_1694);
or U2596 (N_2596,N_1657,N_1906);
nor U2597 (N_2597,N_1433,N_1554);
or U2598 (N_2598,N_1652,N_1424);
nor U2599 (N_2599,N_1183,N_1743);
and U2600 (N_2600,N_1692,N_1051);
nor U2601 (N_2601,N_1090,N_1529);
nand U2602 (N_2602,N_1219,N_1988);
nand U2603 (N_2603,N_1551,N_1239);
and U2604 (N_2604,N_1120,N_1904);
or U2605 (N_2605,N_1200,N_1191);
xnor U2606 (N_2606,N_1023,N_1506);
and U2607 (N_2607,N_1069,N_1669);
and U2608 (N_2608,N_1170,N_1673);
and U2609 (N_2609,N_1298,N_1697);
or U2610 (N_2610,N_1082,N_1267);
nor U2611 (N_2611,N_1139,N_1224);
or U2612 (N_2612,N_1679,N_1641);
nand U2613 (N_2613,N_1643,N_1089);
nand U2614 (N_2614,N_1196,N_1350);
and U2615 (N_2615,N_1234,N_1865);
and U2616 (N_2616,N_1609,N_1757);
nor U2617 (N_2617,N_1424,N_1560);
or U2618 (N_2618,N_1729,N_1103);
nor U2619 (N_2619,N_1285,N_1518);
nor U2620 (N_2620,N_1475,N_1717);
nor U2621 (N_2621,N_1362,N_1699);
nor U2622 (N_2622,N_1026,N_1822);
or U2623 (N_2623,N_1886,N_1970);
nand U2624 (N_2624,N_1171,N_1029);
nand U2625 (N_2625,N_1491,N_1774);
or U2626 (N_2626,N_1241,N_1927);
nand U2627 (N_2627,N_1447,N_1930);
or U2628 (N_2628,N_1179,N_1622);
nand U2629 (N_2629,N_1783,N_1667);
nand U2630 (N_2630,N_1612,N_1479);
nor U2631 (N_2631,N_1556,N_1050);
nor U2632 (N_2632,N_1663,N_1841);
nor U2633 (N_2633,N_1370,N_1789);
nor U2634 (N_2634,N_1960,N_1941);
and U2635 (N_2635,N_1003,N_1302);
or U2636 (N_2636,N_1524,N_1258);
and U2637 (N_2637,N_1351,N_1926);
and U2638 (N_2638,N_1677,N_1600);
or U2639 (N_2639,N_1591,N_1625);
or U2640 (N_2640,N_1785,N_1926);
xnor U2641 (N_2641,N_1816,N_1762);
or U2642 (N_2642,N_1384,N_1790);
or U2643 (N_2643,N_1283,N_1801);
nor U2644 (N_2644,N_1668,N_1852);
or U2645 (N_2645,N_1600,N_1402);
nor U2646 (N_2646,N_1108,N_1130);
nor U2647 (N_2647,N_1610,N_1128);
and U2648 (N_2648,N_1383,N_1293);
or U2649 (N_2649,N_1292,N_1959);
and U2650 (N_2650,N_1784,N_1244);
nand U2651 (N_2651,N_1928,N_1385);
nand U2652 (N_2652,N_1246,N_1628);
nand U2653 (N_2653,N_1271,N_1014);
nand U2654 (N_2654,N_1842,N_1578);
or U2655 (N_2655,N_1004,N_1321);
nand U2656 (N_2656,N_1125,N_1131);
nor U2657 (N_2657,N_1882,N_1114);
nand U2658 (N_2658,N_1753,N_1267);
nor U2659 (N_2659,N_1929,N_1683);
or U2660 (N_2660,N_1534,N_1393);
or U2661 (N_2661,N_1126,N_1597);
or U2662 (N_2662,N_1783,N_1641);
and U2663 (N_2663,N_1138,N_1227);
or U2664 (N_2664,N_1270,N_1416);
or U2665 (N_2665,N_1123,N_1685);
nand U2666 (N_2666,N_1969,N_1962);
and U2667 (N_2667,N_1191,N_1083);
or U2668 (N_2668,N_1737,N_1269);
nor U2669 (N_2669,N_1058,N_1935);
nor U2670 (N_2670,N_1550,N_1294);
or U2671 (N_2671,N_1065,N_1676);
or U2672 (N_2672,N_1838,N_1345);
nor U2673 (N_2673,N_1778,N_1744);
xor U2674 (N_2674,N_1390,N_1513);
or U2675 (N_2675,N_1053,N_1022);
or U2676 (N_2676,N_1841,N_1019);
nand U2677 (N_2677,N_1966,N_1578);
or U2678 (N_2678,N_1822,N_1767);
nand U2679 (N_2679,N_1469,N_1972);
or U2680 (N_2680,N_1433,N_1218);
nor U2681 (N_2681,N_1043,N_1194);
nor U2682 (N_2682,N_1499,N_1155);
nor U2683 (N_2683,N_1721,N_1170);
nand U2684 (N_2684,N_1111,N_1183);
nor U2685 (N_2685,N_1110,N_1743);
nor U2686 (N_2686,N_1529,N_1172);
or U2687 (N_2687,N_1096,N_1409);
nand U2688 (N_2688,N_1452,N_1332);
or U2689 (N_2689,N_1375,N_1849);
nand U2690 (N_2690,N_1998,N_1768);
nand U2691 (N_2691,N_1927,N_1321);
nor U2692 (N_2692,N_1819,N_1069);
nand U2693 (N_2693,N_1286,N_1536);
and U2694 (N_2694,N_1985,N_1888);
nor U2695 (N_2695,N_1918,N_1229);
nor U2696 (N_2696,N_1645,N_1615);
and U2697 (N_2697,N_1932,N_1985);
nor U2698 (N_2698,N_1118,N_1215);
and U2699 (N_2699,N_1535,N_1369);
nor U2700 (N_2700,N_1608,N_1042);
nand U2701 (N_2701,N_1133,N_1817);
nand U2702 (N_2702,N_1423,N_1927);
and U2703 (N_2703,N_1072,N_1902);
nor U2704 (N_2704,N_1052,N_1850);
nand U2705 (N_2705,N_1375,N_1121);
nand U2706 (N_2706,N_1082,N_1931);
nor U2707 (N_2707,N_1582,N_1677);
nand U2708 (N_2708,N_1303,N_1052);
and U2709 (N_2709,N_1476,N_1716);
nor U2710 (N_2710,N_1547,N_1066);
or U2711 (N_2711,N_1934,N_1062);
nor U2712 (N_2712,N_1761,N_1369);
nand U2713 (N_2713,N_1808,N_1874);
or U2714 (N_2714,N_1756,N_1042);
and U2715 (N_2715,N_1645,N_1642);
and U2716 (N_2716,N_1212,N_1536);
and U2717 (N_2717,N_1534,N_1735);
nand U2718 (N_2718,N_1979,N_1281);
or U2719 (N_2719,N_1609,N_1462);
or U2720 (N_2720,N_1781,N_1711);
nand U2721 (N_2721,N_1308,N_1220);
nand U2722 (N_2722,N_1142,N_1111);
or U2723 (N_2723,N_1882,N_1580);
or U2724 (N_2724,N_1086,N_1519);
nor U2725 (N_2725,N_1216,N_1276);
nor U2726 (N_2726,N_1933,N_1145);
or U2727 (N_2727,N_1030,N_1919);
and U2728 (N_2728,N_1959,N_1522);
or U2729 (N_2729,N_1260,N_1663);
or U2730 (N_2730,N_1773,N_1944);
and U2731 (N_2731,N_1402,N_1478);
or U2732 (N_2732,N_1041,N_1901);
or U2733 (N_2733,N_1039,N_1071);
nand U2734 (N_2734,N_1095,N_1243);
nor U2735 (N_2735,N_1180,N_1564);
nor U2736 (N_2736,N_1672,N_1607);
or U2737 (N_2737,N_1617,N_1492);
nand U2738 (N_2738,N_1485,N_1825);
nor U2739 (N_2739,N_1163,N_1693);
or U2740 (N_2740,N_1343,N_1271);
nor U2741 (N_2741,N_1792,N_1557);
nand U2742 (N_2742,N_1112,N_1601);
nor U2743 (N_2743,N_1307,N_1565);
nor U2744 (N_2744,N_1782,N_1662);
nand U2745 (N_2745,N_1628,N_1755);
or U2746 (N_2746,N_1003,N_1152);
nand U2747 (N_2747,N_1322,N_1037);
and U2748 (N_2748,N_1128,N_1852);
nand U2749 (N_2749,N_1348,N_1688);
nor U2750 (N_2750,N_1561,N_1385);
and U2751 (N_2751,N_1376,N_1721);
nand U2752 (N_2752,N_1951,N_1304);
nand U2753 (N_2753,N_1873,N_1223);
or U2754 (N_2754,N_1646,N_1741);
nor U2755 (N_2755,N_1912,N_1478);
nor U2756 (N_2756,N_1389,N_1146);
and U2757 (N_2757,N_1135,N_1491);
or U2758 (N_2758,N_1940,N_1700);
and U2759 (N_2759,N_1370,N_1733);
and U2760 (N_2760,N_1866,N_1520);
nand U2761 (N_2761,N_1881,N_1749);
and U2762 (N_2762,N_1785,N_1844);
nand U2763 (N_2763,N_1093,N_1008);
nor U2764 (N_2764,N_1612,N_1099);
nor U2765 (N_2765,N_1503,N_1977);
or U2766 (N_2766,N_1211,N_1592);
or U2767 (N_2767,N_1052,N_1040);
nor U2768 (N_2768,N_1466,N_1432);
and U2769 (N_2769,N_1410,N_1325);
nand U2770 (N_2770,N_1675,N_1683);
nor U2771 (N_2771,N_1189,N_1461);
nand U2772 (N_2772,N_1050,N_1596);
or U2773 (N_2773,N_1533,N_1714);
nand U2774 (N_2774,N_1530,N_1671);
and U2775 (N_2775,N_1983,N_1390);
nor U2776 (N_2776,N_1006,N_1596);
and U2777 (N_2777,N_1149,N_1734);
or U2778 (N_2778,N_1759,N_1928);
or U2779 (N_2779,N_1062,N_1770);
or U2780 (N_2780,N_1137,N_1860);
or U2781 (N_2781,N_1953,N_1337);
and U2782 (N_2782,N_1591,N_1463);
nand U2783 (N_2783,N_1609,N_1192);
nor U2784 (N_2784,N_1792,N_1709);
and U2785 (N_2785,N_1734,N_1517);
and U2786 (N_2786,N_1331,N_1462);
nand U2787 (N_2787,N_1738,N_1919);
and U2788 (N_2788,N_1014,N_1658);
and U2789 (N_2789,N_1071,N_1085);
nor U2790 (N_2790,N_1812,N_1119);
nor U2791 (N_2791,N_1081,N_1936);
and U2792 (N_2792,N_1931,N_1064);
nand U2793 (N_2793,N_1242,N_1123);
nor U2794 (N_2794,N_1615,N_1432);
and U2795 (N_2795,N_1690,N_1795);
nand U2796 (N_2796,N_1184,N_1872);
or U2797 (N_2797,N_1039,N_1308);
and U2798 (N_2798,N_1640,N_1441);
nand U2799 (N_2799,N_1610,N_1570);
nand U2800 (N_2800,N_1698,N_1330);
nor U2801 (N_2801,N_1954,N_1867);
nand U2802 (N_2802,N_1868,N_1786);
or U2803 (N_2803,N_1141,N_1942);
nor U2804 (N_2804,N_1674,N_1711);
nor U2805 (N_2805,N_1608,N_1726);
or U2806 (N_2806,N_1966,N_1793);
or U2807 (N_2807,N_1684,N_1678);
or U2808 (N_2808,N_1188,N_1085);
and U2809 (N_2809,N_1704,N_1365);
and U2810 (N_2810,N_1686,N_1206);
nor U2811 (N_2811,N_1012,N_1769);
and U2812 (N_2812,N_1721,N_1726);
and U2813 (N_2813,N_1422,N_1918);
nand U2814 (N_2814,N_1843,N_1112);
nand U2815 (N_2815,N_1124,N_1112);
and U2816 (N_2816,N_1334,N_1655);
nor U2817 (N_2817,N_1942,N_1182);
or U2818 (N_2818,N_1115,N_1276);
and U2819 (N_2819,N_1584,N_1592);
nor U2820 (N_2820,N_1208,N_1188);
nor U2821 (N_2821,N_1903,N_1381);
or U2822 (N_2822,N_1559,N_1668);
nor U2823 (N_2823,N_1032,N_1874);
or U2824 (N_2824,N_1601,N_1924);
nand U2825 (N_2825,N_1641,N_1593);
xor U2826 (N_2826,N_1394,N_1817);
nor U2827 (N_2827,N_1998,N_1551);
and U2828 (N_2828,N_1539,N_1203);
and U2829 (N_2829,N_1161,N_1196);
nand U2830 (N_2830,N_1491,N_1752);
or U2831 (N_2831,N_1926,N_1636);
and U2832 (N_2832,N_1981,N_1819);
nand U2833 (N_2833,N_1324,N_1298);
or U2834 (N_2834,N_1410,N_1845);
nor U2835 (N_2835,N_1523,N_1598);
nor U2836 (N_2836,N_1087,N_1428);
and U2837 (N_2837,N_1914,N_1012);
or U2838 (N_2838,N_1983,N_1160);
nor U2839 (N_2839,N_1275,N_1877);
or U2840 (N_2840,N_1936,N_1484);
nor U2841 (N_2841,N_1284,N_1402);
xnor U2842 (N_2842,N_1136,N_1939);
and U2843 (N_2843,N_1223,N_1292);
nor U2844 (N_2844,N_1129,N_1646);
or U2845 (N_2845,N_1347,N_1111);
and U2846 (N_2846,N_1234,N_1060);
and U2847 (N_2847,N_1061,N_1544);
and U2848 (N_2848,N_1978,N_1027);
nand U2849 (N_2849,N_1108,N_1435);
nor U2850 (N_2850,N_1264,N_1818);
nand U2851 (N_2851,N_1186,N_1894);
xnor U2852 (N_2852,N_1928,N_1560);
nand U2853 (N_2853,N_1923,N_1142);
or U2854 (N_2854,N_1368,N_1543);
nor U2855 (N_2855,N_1725,N_1371);
nand U2856 (N_2856,N_1268,N_1805);
nand U2857 (N_2857,N_1964,N_1200);
nor U2858 (N_2858,N_1234,N_1160);
and U2859 (N_2859,N_1620,N_1396);
nor U2860 (N_2860,N_1644,N_1097);
nor U2861 (N_2861,N_1674,N_1020);
nor U2862 (N_2862,N_1534,N_1531);
nor U2863 (N_2863,N_1245,N_1418);
or U2864 (N_2864,N_1610,N_1685);
nor U2865 (N_2865,N_1541,N_1136);
nand U2866 (N_2866,N_1222,N_1701);
xor U2867 (N_2867,N_1803,N_1195);
or U2868 (N_2868,N_1384,N_1069);
and U2869 (N_2869,N_1435,N_1081);
or U2870 (N_2870,N_1012,N_1033);
nand U2871 (N_2871,N_1242,N_1869);
or U2872 (N_2872,N_1454,N_1822);
nand U2873 (N_2873,N_1211,N_1180);
nand U2874 (N_2874,N_1311,N_1709);
and U2875 (N_2875,N_1921,N_1512);
nand U2876 (N_2876,N_1658,N_1230);
and U2877 (N_2877,N_1290,N_1759);
and U2878 (N_2878,N_1835,N_1578);
nand U2879 (N_2879,N_1666,N_1473);
nand U2880 (N_2880,N_1562,N_1691);
nor U2881 (N_2881,N_1587,N_1249);
nand U2882 (N_2882,N_1089,N_1613);
or U2883 (N_2883,N_1546,N_1427);
nand U2884 (N_2884,N_1574,N_1539);
and U2885 (N_2885,N_1070,N_1445);
nand U2886 (N_2886,N_1496,N_1344);
nand U2887 (N_2887,N_1539,N_1343);
or U2888 (N_2888,N_1170,N_1360);
nor U2889 (N_2889,N_1948,N_1314);
nor U2890 (N_2890,N_1588,N_1570);
nor U2891 (N_2891,N_1748,N_1234);
nor U2892 (N_2892,N_1135,N_1594);
nand U2893 (N_2893,N_1732,N_1799);
nand U2894 (N_2894,N_1898,N_1728);
nand U2895 (N_2895,N_1529,N_1339);
nor U2896 (N_2896,N_1568,N_1389);
nand U2897 (N_2897,N_1276,N_1041);
nor U2898 (N_2898,N_1301,N_1288);
and U2899 (N_2899,N_1865,N_1962);
nand U2900 (N_2900,N_1958,N_1307);
or U2901 (N_2901,N_1006,N_1325);
nand U2902 (N_2902,N_1823,N_1181);
and U2903 (N_2903,N_1150,N_1911);
nor U2904 (N_2904,N_1166,N_1498);
and U2905 (N_2905,N_1211,N_1426);
nor U2906 (N_2906,N_1257,N_1087);
or U2907 (N_2907,N_1204,N_1748);
nand U2908 (N_2908,N_1226,N_1468);
and U2909 (N_2909,N_1726,N_1660);
nand U2910 (N_2910,N_1005,N_1240);
nor U2911 (N_2911,N_1567,N_1533);
nor U2912 (N_2912,N_1606,N_1478);
nand U2913 (N_2913,N_1303,N_1851);
and U2914 (N_2914,N_1899,N_1502);
and U2915 (N_2915,N_1606,N_1146);
nand U2916 (N_2916,N_1205,N_1455);
or U2917 (N_2917,N_1348,N_1557);
and U2918 (N_2918,N_1403,N_1066);
nand U2919 (N_2919,N_1320,N_1241);
nand U2920 (N_2920,N_1522,N_1152);
nand U2921 (N_2921,N_1989,N_1587);
and U2922 (N_2922,N_1549,N_1646);
nor U2923 (N_2923,N_1810,N_1807);
nand U2924 (N_2924,N_1539,N_1948);
and U2925 (N_2925,N_1206,N_1606);
nand U2926 (N_2926,N_1210,N_1639);
nor U2927 (N_2927,N_1668,N_1951);
or U2928 (N_2928,N_1890,N_1911);
nand U2929 (N_2929,N_1790,N_1281);
or U2930 (N_2930,N_1679,N_1871);
nand U2931 (N_2931,N_1115,N_1303);
nor U2932 (N_2932,N_1067,N_1478);
nand U2933 (N_2933,N_1332,N_1680);
and U2934 (N_2934,N_1636,N_1107);
nand U2935 (N_2935,N_1892,N_1053);
nor U2936 (N_2936,N_1674,N_1865);
or U2937 (N_2937,N_1426,N_1997);
nor U2938 (N_2938,N_1437,N_1862);
nand U2939 (N_2939,N_1815,N_1441);
or U2940 (N_2940,N_1238,N_1056);
and U2941 (N_2941,N_1550,N_1614);
nand U2942 (N_2942,N_1173,N_1706);
nor U2943 (N_2943,N_1735,N_1671);
or U2944 (N_2944,N_1113,N_1313);
nand U2945 (N_2945,N_1283,N_1161);
or U2946 (N_2946,N_1637,N_1134);
nor U2947 (N_2947,N_1046,N_1168);
and U2948 (N_2948,N_1093,N_1818);
nand U2949 (N_2949,N_1674,N_1834);
or U2950 (N_2950,N_1669,N_1202);
nand U2951 (N_2951,N_1071,N_1702);
and U2952 (N_2952,N_1760,N_1674);
or U2953 (N_2953,N_1280,N_1877);
or U2954 (N_2954,N_1411,N_1507);
nor U2955 (N_2955,N_1976,N_1764);
and U2956 (N_2956,N_1278,N_1335);
and U2957 (N_2957,N_1219,N_1890);
nor U2958 (N_2958,N_1261,N_1059);
nor U2959 (N_2959,N_1861,N_1037);
nor U2960 (N_2960,N_1091,N_1212);
nand U2961 (N_2961,N_1403,N_1565);
nor U2962 (N_2962,N_1978,N_1135);
nand U2963 (N_2963,N_1839,N_1243);
xnor U2964 (N_2964,N_1908,N_1093);
or U2965 (N_2965,N_1099,N_1528);
or U2966 (N_2966,N_1670,N_1615);
nand U2967 (N_2967,N_1942,N_1861);
and U2968 (N_2968,N_1753,N_1231);
or U2969 (N_2969,N_1467,N_1296);
and U2970 (N_2970,N_1656,N_1521);
nor U2971 (N_2971,N_1500,N_1450);
nand U2972 (N_2972,N_1067,N_1482);
nor U2973 (N_2973,N_1261,N_1410);
nor U2974 (N_2974,N_1111,N_1604);
or U2975 (N_2975,N_1133,N_1150);
nand U2976 (N_2976,N_1213,N_1676);
and U2977 (N_2977,N_1795,N_1536);
nand U2978 (N_2978,N_1289,N_1475);
nor U2979 (N_2979,N_1612,N_1839);
or U2980 (N_2980,N_1966,N_1641);
or U2981 (N_2981,N_1897,N_1766);
or U2982 (N_2982,N_1689,N_1763);
nand U2983 (N_2983,N_1487,N_1559);
xnor U2984 (N_2984,N_1268,N_1663);
or U2985 (N_2985,N_1523,N_1350);
or U2986 (N_2986,N_1798,N_1688);
nand U2987 (N_2987,N_1023,N_1298);
or U2988 (N_2988,N_1678,N_1111);
and U2989 (N_2989,N_1941,N_1647);
and U2990 (N_2990,N_1763,N_1578);
nor U2991 (N_2991,N_1353,N_1978);
and U2992 (N_2992,N_1505,N_1741);
nor U2993 (N_2993,N_1274,N_1526);
or U2994 (N_2994,N_1332,N_1905);
nand U2995 (N_2995,N_1789,N_1456);
nand U2996 (N_2996,N_1602,N_1300);
or U2997 (N_2997,N_1240,N_1825);
nor U2998 (N_2998,N_1030,N_1140);
or U2999 (N_2999,N_1454,N_1492);
nor U3000 (N_3000,N_2627,N_2528);
and U3001 (N_3001,N_2955,N_2920);
nor U3002 (N_3002,N_2663,N_2435);
or U3003 (N_3003,N_2999,N_2762);
and U3004 (N_3004,N_2283,N_2691);
nand U3005 (N_3005,N_2374,N_2657);
nand U3006 (N_3006,N_2436,N_2182);
nor U3007 (N_3007,N_2839,N_2797);
nand U3008 (N_3008,N_2269,N_2926);
nor U3009 (N_3009,N_2055,N_2879);
nand U3010 (N_3010,N_2613,N_2469);
or U3011 (N_3011,N_2750,N_2619);
or U3012 (N_3012,N_2466,N_2136);
or U3013 (N_3013,N_2796,N_2725);
and U3014 (N_3014,N_2502,N_2395);
nand U3015 (N_3015,N_2591,N_2217);
or U3016 (N_3016,N_2792,N_2549);
or U3017 (N_3017,N_2571,N_2337);
and U3018 (N_3018,N_2253,N_2565);
nor U3019 (N_3019,N_2876,N_2525);
and U3020 (N_3020,N_2574,N_2851);
or U3021 (N_3021,N_2302,N_2806);
or U3022 (N_3022,N_2458,N_2633);
and U3023 (N_3023,N_2317,N_2365);
nor U3024 (N_3024,N_2264,N_2594);
nand U3025 (N_3025,N_2043,N_2980);
and U3026 (N_3026,N_2780,N_2867);
nand U3027 (N_3027,N_2626,N_2054);
and U3028 (N_3028,N_2501,N_2494);
or U3029 (N_3029,N_2397,N_2389);
or U3030 (N_3030,N_2804,N_2786);
or U3031 (N_3031,N_2900,N_2148);
or U3032 (N_3032,N_2758,N_2120);
nor U3033 (N_3033,N_2831,N_2991);
and U3034 (N_3034,N_2498,N_2767);
nand U3035 (N_3035,N_2297,N_2132);
nor U3036 (N_3036,N_2260,N_2238);
or U3037 (N_3037,N_2412,N_2500);
nor U3038 (N_3038,N_2930,N_2721);
or U3039 (N_3039,N_2551,N_2966);
nor U3040 (N_3040,N_2661,N_2172);
or U3041 (N_3041,N_2603,N_2381);
nand U3042 (N_3042,N_2356,N_2899);
and U3043 (N_3043,N_2883,N_2101);
or U3044 (N_3044,N_2401,N_2474);
and U3045 (N_3045,N_2735,N_2402);
nand U3046 (N_3046,N_2219,N_2905);
or U3047 (N_3047,N_2104,N_2184);
nand U3048 (N_3048,N_2933,N_2962);
or U3049 (N_3049,N_2250,N_2138);
nor U3050 (N_3050,N_2270,N_2959);
or U3051 (N_3051,N_2592,N_2413);
and U3052 (N_3052,N_2378,N_2188);
and U3053 (N_3053,N_2830,N_2433);
nor U3054 (N_3054,N_2340,N_2373);
or U3055 (N_3055,N_2785,N_2858);
or U3056 (N_3056,N_2979,N_2271);
nand U3057 (N_3057,N_2699,N_2004);
and U3058 (N_3058,N_2802,N_2376);
xor U3059 (N_3059,N_2214,N_2307);
nand U3060 (N_3060,N_2838,N_2958);
nor U3061 (N_3061,N_2601,N_2090);
nor U3062 (N_3062,N_2994,N_2712);
nor U3063 (N_3063,N_2470,N_2202);
nor U3064 (N_3064,N_2332,N_2970);
or U3065 (N_3065,N_2022,N_2825);
nor U3066 (N_3066,N_2514,N_2097);
nand U3067 (N_3067,N_2150,N_2616);
and U3068 (N_3068,N_2504,N_2468);
nand U3069 (N_3069,N_2372,N_2559);
nor U3070 (N_3070,N_2940,N_2461);
nor U3071 (N_3071,N_2308,N_2153);
or U3072 (N_3072,N_2485,N_2367);
and U3073 (N_3073,N_2885,N_2612);
or U3074 (N_3074,N_2639,N_2724);
nor U3075 (N_3075,N_2487,N_2464);
nand U3076 (N_3076,N_2718,N_2027);
or U3077 (N_3077,N_2456,N_2342);
nand U3078 (N_3078,N_2204,N_2956);
nand U3079 (N_3079,N_2019,N_2985);
nor U3080 (N_3080,N_2625,N_2366);
nor U3081 (N_3081,N_2322,N_2040);
and U3082 (N_3082,N_2477,N_2998);
or U3083 (N_3083,N_2617,N_2508);
nor U3084 (N_3084,N_2646,N_2535);
and U3085 (N_3085,N_2465,N_2775);
or U3086 (N_3086,N_2254,N_2223);
nor U3087 (N_3087,N_2781,N_2803);
and U3088 (N_3088,N_2490,N_2945);
nor U3089 (N_3089,N_2768,N_2629);
nand U3090 (N_3090,N_2163,N_2094);
nor U3091 (N_3091,N_2935,N_2137);
and U3092 (N_3092,N_2537,N_2563);
nand U3093 (N_3093,N_2632,N_2353);
or U3094 (N_3094,N_2276,N_2908);
or U3095 (N_3095,N_2904,N_2773);
or U3096 (N_3096,N_2131,N_2700);
and U3097 (N_3097,N_2392,N_2868);
nand U3098 (N_3098,N_2201,N_2406);
or U3099 (N_3099,N_2808,N_2751);
and U3100 (N_3100,N_2309,N_2690);
and U3101 (N_3101,N_2578,N_2769);
nor U3102 (N_3102,N_2482,N_2074);
and U3103 (N_3103,N_2647,N_2369);
nor U3104 (N_3104,N_2357,N_2720);
nand U3105 (N_3105,N_2305,N_2007);
nor U3106 (N_3106,N_2987,N_2403);
and U3107 (N_3107,N_2348,N_2967);
nor U3108 (N_3108,N_2258,N_2496);
nor U3109 (N_3109,N_2414,N_2493);
nand U3110 (N_3110,N_2070,N_2957);
nand U3111 (N_3111,N_2067,N_2584);
or U3112 (N_3112,N_2239,N_2748);
nand U3113 (N_3113,N_2261,N_2705);
nand U3114 (N_3114,N_2451,N_2836);
nand U3115 (N_3115,N_2562,N_2282);
or U3116 (N_3116,N_2000,N_2810);
and U3117 (N_3117,N_2244,N_2198);
or U3118 (N_3118,N_2512,N_2986);
or U3119 (N_3119,N_2794,N_2637);
nand U3120 (N_3120,N_2375,N_2636);
and U3121 (N_3121,N_2763,N_2916);
nand U3122 (N_3122,N_2734,N_2864);
and U3123 (N_3123,N_2950,N_2942);
nor U3124 (N_3124,N_2921,N_2227);
nor U3125 (N_3125,N_2284,N_2078);
or U3126 (N_3126,N_2206,N_2462);
nor U3127 (N_3127,N_2896,N_2823);
or U3128 (N_3128,N_2641,N_2278);
and U3129 (N_3129,N_2852,N_2850);
or U3130 (N_3130,N_2427,N_2121);
and U3131 (N_3131,N_2404,N_2973);
and U3132 (N_3132,N_2252,N_2515);
and U3133 (N_3133,N_2939,N_2848);
nand U3134 (N_3134,N_2505,N_2558);
or U3135 (N_3135,N_2678,N_2066);
or U3136 (N_3136,N_2303,N_2053);
and U3137 (N_3137,N_2918,N_2113);
and U3138 (N_3138,N_2285,N_2706);
and U3139 (N_3139,N_2405,N_2051);
nor U3140 (N_3140,N_2795,N_2901);
and U3141 (N_3141,N_2936,N_2096);
or U3142 (N_3142,N_2886,N_2506);
nor U3143 (N_3143,N_2221,N_2207);
nor U3144 (N_3144,N_2683,N_2550);
or U3145 (N_3145,N_2503,N_2368);
nand U3146 (N_3146,N_2228,N_2640);
and U3147 (N_3147,N_2527,N_2715);
nor U3148 (N_3148,N_2299,N_2952);
nor U3149 (N_3149,N_2892,N_2906);
nand U3150 (N_3150,N_2419,N_2710);
or U3151 (N_3151,N_2915,N_2866);
or U3152 (N_3152,N_2013,N_2453);
xnor U3153 (N_3153,N_2789,N_2679);
xor U3154 (N_3154,N_2573,N_2776);
nand U3155 (N_3155,N_2263,N_2924);
nand U3156 (N_3156,N_2649,N_2701);
nand U3157 (N_3157,N_2151,N_2437);
nand U3158 (N_3158,N_2960,N_2621);
nor U3159 (N_3159,N_2364,N_2449);
nor U3160 (N_3160,N_2604,N_2726);
or U3161 (N_3161,N_2077,N_2118);
or U3162 (N_3162,N_2107,N_2814);
nor U3163 (N_3163,N_2658,N_2542);
and U3164 (N_3164,N_2877,N_2544);
or U3165 (N_3165,N_2166,N_2492);
and U3166 (N_3166,N_2393,N_2079);
or U3167 (N_3167,N_2688,N_2672);
and U3168 (N_3168,N_2519,N_2801);
nor U3169 (N_3169,N_2783,N_2106);
nor U3170 (N_3170,N_2215,N_2511);
nor U3171 (N_3171,N_2034,N_2241);
nand U3172 (N_3172,N_2233,N_2919);
nand U3173 (N_3173,N_2418,N_2310);
and U3174 (N_3174,N_2031,N_2992);
nand U3175 (N_3175,N_2593,N_2175);
nor U3176 (N_3176,N_2092,N_2362);
nor U3177 (N_3177,N_2122,N_2532);
or U3178 (N_3178,N_2267,N_2727);
nand U3179 (N_3179,N_2881,N_2390);
nor U3180 (N_3180,N_2125,N_2430);
or U3181 (N_3181,N_2387,N_2028);
or U3182 (N_3182,N_2196,N_2912);
nand U3183 (N_3183,N_2197,N_2460);
and U3184 (N_3184,N_2846,N_2420);
nand U3185 (N_3185,N_2618,N_2115);
or U3186 (N_3186,N_2878,N_2272);
and U3187 (N_3187,N_2731,N_2909);
nor U3188 (N_3188,N_2320,N_2447);
nand U3189 (N_3189,N_2495,N_2609);
or U3190 (N_3190,N_2161,N_2290);
nor U3191 (N_3191,N_2334,N_2638);
and U3192 (N_3192,N_2692,N_2583);
nand U3193 (N_3193,N_2388,N_2772);
or U3194 (N_3194,N_2399,N_2898);
and U3195 (N_3195,N_2713,N_2854);
or U3196 (N_3196,N_2743,N_2127);
and U3197 (N_3197,N_2730,N_2704);
and U3198 (N_3198,N_2738,N_2664);
or U3199 (N_3199,N_2010,N_2656);
nand U3200 (N_3200,N_2124,N_2099);
or U3201 (N_3201,N_2765,N_2448);
nor U3202 (N_3202,N_2651,N_2360);
nor U3203 (N_3203,N_2383,N_2990);
nor U3204 (N_3204,N_2614,N_2821);
nand U3205 (N_3205,N_2220,N_2602);
or U3206 (N_3206,N_2741,N_2133);
nor U3207 (N_3207,N_2585,N_2666);
nor U3208 (N_3208,N_2819,N_2554);
or U3209 (N_3209,N_2063,N_2024);
nor U3210 (N_3210,N_2109,N_2863);
and U3211 (N_3211,N_2524,N_2379);
nor U3212 (N_3212,N_2655,N_2209);
nand U3213 (N_3213,N_2586,N_2072);
or U3214 (N_3214,N_2178,N_2319);
or U3215 (N_3215,N_2428,N_2590);
and U3216 (N_3216,N_2681,N_2662);
xnor U3217 (N_3217,N_2513,N_2050);
nand U3218 (N_3218,N_2415,N_2711);
nand U3219 (N_3219,N_2893,N_2280);
or U3220 (N_3220,N_2164,N_2287);
and U3221 (N_3221,N_2871,N_2032);
nor U3222 (N_3222,N_2680,N_2907);
nor U3223 (N_3223,N_2300,N_2351);
and U3224 (N_3224,N_2169,N_2739);
and U3225 (N_3225,N_2384,N_2103);
and U3226 (N_3226,N_2306,N_2294);
nor U3227 (N_3227,N_2003,N_2702);
nand U3228 (N_3228,N_2296,N_2949);
nor U3229 (N_3229,N_2870,N_2954);
or U3230 (N_3230,N_2203,N_2245);
nand U3231 (N_3231,N_2882,N_2934);
nor U3232 (N_3232,N_2443,N_2095);
or U3233 (N_3233,N_2273,N_2579);
or U3234 (N_3234,N_2927,N_2039);
nor U3235 (N_3235,N_2671,N_2110);
nor U3236 (N_3236,N_2564,N_2518);
nor U3237 (N_3237,N_2432,N_2938);
nor U3238 (N_3238,N_2820,N_2665);
and U3239 (N_3239,N_2048,N_2326);
and U3240 (N_3240,N_2976,N_2242);
and U3241 (N_3241,N_2860,N_2128);
nand U3242 (N_3242,N_2811,N_2234);
and U3243 (N_3243,N_2536,N_2006);
or U3244 (N_3244,N_2526,N_2277);
nor U3245 (N_3245,N_2422,N_2445);
nor U3246 (N_3246,N_2472,N_2195);
or U3247 (N_3247,N_2246,N_2771);
nand U3248 (N_3248,N_2538,N_2130);
nand U3249 (N_3249,N_2540,N_2723);
or U3250 (N_3250,N_2480,N_2589);
and U3251 (N_3251,N_2257,N_2793);
nor U3252 (N_3252,N_2098,N_2757);
nor U3253 (N_3253,N_2483,N_2622);
and U3254 (N_3254,N_2624,N_2611);
nand U3255 (N_3255,N_2328,N_2676);
nor U3256 (N_3256,N_2732,N_2989);
and U3257 (N_3257,N_2889,N_2961);
or U3258 (N_3258,N_2210,N_2600);
nor U3259 (N_3259,N_2016,N_2547);
nor U3260 (N_3260,N_2965,N_2174);
and U3261 (N_3261,N_2696,N_2479);
nor U3262 (N_3262,N_2291,N_2910);
and U3263 (N_3263,N_2782,N_2440);
or U3264 (N_3264,N_2813,N_2737);
nand U3265 (N_3265,N_2798,N_2828);
nand U3266 (N_3266,N_2343,N_2510);
and U3267 (N_3267,N_2971,N_2231);
or U3268 (N_3268,N_2969,N_2902);
nor U3269 (N_3269,N_2396,N_2005);
nand U3270 (N_3270,N_2145,N_2807);
nor U3271 (N_3271,N_2059,N_2069);
nor U3272 (N_3272,N_2972,N_2753);
nand U3273 (N_3273,N_2596,N_2628);
nand U3274 (N_3274,N_2186,N_2111);
nand U3275 (N_3275,N_2832,N_2568);
nor U3276 (N_3276,N_2685,N_2385);
and U3277 (N_3277,N_2035,N_2324);
nor U3278 (N_3278,N_2083,N_2358);
nand U3279 (N_3279,N_2996,N_2194);
nand U3280 (N_3280,N_2312,N_2824);
or U3281 (N_3281,N_2635,N_2517);
nor U3282 (N_3282,N_2327,N_2088);
and U3283 (N_3283,N_2709,N_2314);
nor U3284 (N_3284,N_2108,N_2543);
nor U3285 (N_3285,N_2191,N_2890);
nand U3286 (N_3286,N_2076,N_2650);
and U3287 (N_3287,N_2084,N_2684);
nor U3288 (N_3288,N_2862,N_2471);
nor U3289 (N_3289,N_2352,N_2315);
nor U3290 (N_3290,N_2249,N_2922);
and U3291 (N_3291,N_2382,N_2599);
or U3292 (N_3292,N_2499,N_2761);
nand U3293 (N_3293,N_2259,N_2759);
nor U3294 (N_3294,N_2149,N_2873);
and U3295 (N_3295,N_2895,N_2642);
or U3296 (N_3296,N_2817,N_2157);
or U3297 (N_3297,N_2714,N_2189);
or U3298 (N_3298,N_2323,N_2350);
nor U3299 (N_3299,N_2086,N_2744);
nor U3300 (N_3300,N_2648,N_2114);
nor U3301 (N_3301,N_2330,N_2615);
and U3302 (N_3302,N_2398,N_2667);
or U3303 (N_3303,N_2064,N_2968);
nand U3304 (N_3304,N_2911,N_2682);
and U3305 (N_3305,N_2693,N_2778);
nor U3306 (N_3306,N_2236,N_2339);
nor U3307 (N_3307,N_2446,N_2229);
or U3308 (N_3308,N_2187,N_2116);
nand U3309 (N_3309,N_2875,N_2335);
and U3310 (N_3310,N_2903,N_2588);
or U3311 (N_3311,N_2347,N_2747);
and U3312 (N_3312,N_2791,N_2859);
nor U3313 (N_3313,N_2497,N_2833);
or U3314 (N_3314,N_2974,N_2481);
nor U3315 (N_3315,N_2520,N_2318);
and U3316 (N_3316,N_2719,N_2837);
or U3317 (N_3317,N_2799,N_2716);
nand U3318 (N_3318,N_2809,N_2861);
nand U3319 (N_3319,N_2756,N_2183);
or U3320 (N_3320,N_2224,N_2643);
and U3321 (N_3321,N_2377,N_2018);
nor U3322 (N_3322,N_2030,N_2673);
nand U3323 (N_3323,N_2995,N_2298);
or U3324 (N_3324,N_2452,N_2065);
nand U3325 (N_3325,N_2689,N_2391);
nor U3326 (N_3326,N_2555,N_2587);
nor U3327 (N_3327,N_2015,N_2286);
and U3328 (N_3328,N_2255,N_2946);
or U3329 (N_3329,N_2556,N_2192);
nor U3330 (N_3330,N_2193,N_2361);
nand U3331 (N_3331,N_2230,N_2595);
nor U3332 (N_3332,N_2251,N_2522);
nor U3333 (N_3333,N_2533,N_2222);
nor U3334 (N_3334,N_2425,N_2698);
or U3335 (N_3335,N_2087,N_2677);
and U3336 (N_3336,N_2226,N_2552);
or U3337 (N_3337,N_2329,N_2407);
or U3338 (N_3338,N_2770,N_2888);
and U3339 (N_3339,N_2156,N_2014);
nor U3340 (N_3340,N_2185,N_2438);
and U3341 (N_3341,N_2232,N_2333);
and U3342 (N_3342,N_2017,N_2659);
and U3343 (N_3343,N_2042,N_2026);
and U3344 (N_3344,N_2235,N_2075);
or U3345 (N_3345,N_2884,N_2044);
nand U3346 (N_3346,N_2722,N_2855);
and U3347 (N_3347,N_2580,N_2135);
nand U3348 (N_3348,N_2887,N_2993);
xor U3349 (N_3349,N_2341,N_2311);
or U3350 (N_3350,N_2872,N_2717);
and U3351 (N_3351,N_2177,N_2355);
and U3352 (N_3352,N_2205,N_2816);
nor U3353 (N_3353,N_2331,N_2047);
and U3354 (N_3354,N_2213,N_2755);
nand U3355 (N_3355,N_2478,N_2708);
or U3356 (N_3356,N_2129,N_2844);
or U3357 (N_3357,N_2410,N_2598);
and U3358 (N_3358,N_2293,N_2507);
nor U3359 (N_3359,N_2171,N_2948);
and U3360 (N_3360,N_2874,N_2301);
or U3361 (N_3361,N_2812,N_2694);
and U3362 (N_3362,N_2845,N_2764);
nand U3363 (N_3363,N_2695,N_2847);
and U3364 (N_3364,N_2141,N_2321);
nor U3365 (N_3365,N_2349,N_2857);
and U3366 (N_3366,N_2788,N_2008);
nand U3367 (N_3367,N_2931,N_2036);
xnor U3368 (N_3368,N_2325,N_2733);
or U3369 (N_3369,N_2707,N_2068);
or U3370 (N_3370,N_2434,N_2237);
and U3371 (N_3371,N_2400,N_2416);
or U3372 (N_3372,N_2645,N_2144);
and U3373 (N_3373,N_2046,N_2200);
nor U3374 (N_3374,N_2009,N_2045);
and U3375 (N_3375,N_2081,N_2212);
or U3376 (N_3376,N_2160,N_2162);
nand U3377 (N_3377,N_2338,N_2279);
and U3378 (N_3378,N_2652,N_2476);
nand U3379 (N_3379,N_2243,N_2581);
and U3380 (N_3380,N_2091,N_2167);
nor U3381 (N_3381,N_2644,N_2021);
or U3382 (N_3382,N_2582,N_2787);
and U3383 (N_3383,N_2539,N_2869);
nor U3384 (N_3384,N_2292,N_2728);
nand U3385 (N_3385,N_2266,N_2442);
nor U3386 (N_3386,N_2488,N_2923);
or U3387 (N_3387,N_2165,N_2057);
or U3388 (N_3388,N_2981,N_2181);
nand U3389 (N_3389,N_2853,N_2608);
nor U3390 (N_3390,N_2216,N_2313);
nand U3391 (N_3391,N_2439,N_2729);
nor U3392 (N_3392,N_2937,N_2849);
nand U3393 (N_3393,N_2208,N_2450);
or U3394 (N_3394,N_2553,N_2033);
and U3395 (N_3395,N_2545,N_2423);
nor U3396 (N_3396,N_2566,N_2557);
or U3397 (N_3397,N_2168,N_2978);
or U3398 (N_3398,N_2176,N_2509);
nor U3399 (N_3399,N_2630,N_2843);
and U3400 (N_3400,N_2093,N_2179);
and U3401 (N_3401,N_2371,N_2199);
nand U3402 (N_3402,N_2605,N_2800);
or U3403 (N_3403,N_2105,N_2170);
nand U3404 (N_3404,N_2012,N_2675);
nand U3405 (N_3405,N_2152,N_2982);
or U3406 (N_3406,N_2570,N_2117);
or U3407 (N_3407,N_2288,N_2606);
and U3408 (N_3408,N_2459,N_2745);
or U3409 (N_3409,N_2546,N_2475);
and U3410 (N_3410,N_2597,N_2248);
and U3411 (N_3411,N_2572,N_2523);
or U3412 (N_3412,N_2548,N_2917);
nand U3413 (N_3413,N_2247,N_2180);
nand U3414 (N_3414,N_2211,N_2444);
nand U3415 (N_3415,N_2346,N_2023);
nor U3416 (N_3416,N_2411,N_2240);
nor U3417 (N_3417,N_2218,N_2818);
or U3418 (N_3418,N_2142,N_2073);
nand U3419 (N_3419,N_2058,N_2085);
and U3420 (N_3420,N_2473,N_2686);
nand U3421 (N_3421,N_2029,N_2560);
and U3422 (N_3422,N_2463,N_2275);
nor U3423 (N_3423,N_2654,N_2941);
nor U3424 (N_3424,N_2426,N_2489);
nor U3425 (N_3425,N_2736,N_2359);
nand U3426 (N_3426,N_2703,N_2674);
nand U3427 (N_3427,N_2486,N_2052);
nand U3428 (N_3428,N_2964,N_2295);
or U3429 (N_3429,N_2623,N_2281);
nand U3430 (N_3430,N_2944,N_2457);
nand U3431 (N_3431,N_2607,N_2576);
nand U3432 (N_3432,N_2740,N_2268);
or U3433 (N_3433,N_2467,N_2669);
and U3434 (N_3434,N_2408,N_2380);
and U3435 (N_3435,N_2766,N_2894);
or U3436 (N_3436,N_2687,N_2947);
or U3437 (N_3437,N_2037,N_2827);
and U3438 (N_3438,N_2134,N_2225);
nor U3439 (N_3439,N_2529,N_2455);
or U3440 (N_3440,N_2190,N_2943);
and U3441 (N_3441,N_2610,N_2424);
or U3442 (N_3442,N_2577,N_2336);
xor U3443 (N_3443,N_2746,N_2856);
or U3444 (N_3444,N_2670,N_2575);
or U3445 (N_3445,N_2530,N_2089);
nand U3446 (N_3446,N_2567,N_2173);
or U3447 (N_3447,N_2822,N_2140);
nand U3448 (N_3448,N_2119,N_2805);
nor U3449 (N_3449,N_2421,N_2897);
or U3450 (N_3450,N_2790,N_2441);
or U3451 (N_3451,N_2123,N_2020);
nor U3452 (N_3452,N_2060,N_2865);
or U3453 (N_3453,N_2988,N_2760);
or U3454 (N_3454,N_2061,N_2561);
and U3455 (N_3455,N_2344,N_2913);
nor U3456 (N_3456,N_2011,N_2953);
and U3457 (N_3457,N_2001,N_2880);
and U3458 (N_3458,N_2779,N_2159);
xor U3459 (N_3459,N_2826,N_2742);
and U3460 (N_3460,N_2262,N_2102);
nor U3461 (N_3461,N_2840,N_2997);
and U3462 (N_3462,N_2491,N_2914);
or U3463 (N_3463,N_2394,N_2038);
and U3464 (N_3464,N_2049,N_2975);
nor U3465 (N_3465,N_2631,N_2154);
and U3466 (N_3466,N_2345,N_2041);
and U3467 (N_3467,N_2158,N_2784);
nand U3468 (N_3468,N_2835,N_2521);
or U3469 (N_3469,N_2082,N_2409);
nor U3470 (N_3470,N_2925,N_2531);
nand U3471 (N_3471,N_2634,N_2929);
and U3472 (N_3472,N_2370,N_2025);
nor U3473 (N_3473,N_2080,N_2891);
or U3474 (N_3474,N_2256,N_2752);
nor U3475 (N_3475,N_2147,N_2146);
and U3476 (N_3476,N_2289,N_2126);
nand U3477 (N_3477,N_2983,N_2951);
nand U3478 (N_3478,N_2620,N_2274);
nor U3479 (N_3479,N_2541,N_2056);
or U3480 (N_3480,N_2100,N_2431);
or U3481 (N_3481,N_2928,N_2932);
nor U3482 (N_3482,N_2815,N_2354);
or U3483 (N_3483,N_2386,N_2363);
and U3484 (N_3484,N_2841,N_2454);
nor U3485 (N_3485,N_2143,N_2516);
nor U3486 (N_3486,N_2139,N_2777);
or U3487 (N_3487,N_2304,N_2984);
nor U3488 (N_3488,N_2668,N_2749);
and U3489 (N_3489,N_2484,N_2569);
nand U3490 (N_3490,N_2071,N_2963);
nor U3491 (N_3491,N_2653,N_2660);
or U3492 (N_3492,N_2829,N_2834);
and U3493 (N_3493,N_2002,N_2429);
nand U3494 (N_3494,N_2697,N_2977);
nand U3495 (N_3495,N_2155,N_2842);
and U3496 (N_3496,N_2316,N_2062);
and U3497 (N_3497,N_2265,N_2774);
nor U3498 (N_3498,N_2112,N_2534);
or U3499 (N_3499,N_2417,N_2754);
or U3500 (N_3500,N_2572,N_2284);
nand U3501 (N_3501,N_2726,N_2045);
or U3502 (N_3502,N_2734,N_2865);
nand U3503 (N_3503,N_2027,N_2335);
nand U3504 (N_3504,N_2752,N_2367);
and U3505 (N_3505,N_2920,N_2904);
or U3506 (N_3506,N_2700,N_2978);
or U3507 (N_3507,N_2188,N_2010);
or U3508 (N_3508,N_2045,N_2976);
nand U3509 (N_3509,N_2140,N_2473);
nand U3510 (N_3510,N_2600,N_2120);
nand U3511 (N_3511,N_2761,N_2137);
and U3512 (N_3512,N_2252,N_2196);
nor U3513 (N_3513,N_2678,N_2796);
or U3514 (N_3514,N_2696,N_2023);
nor U3515 (N_3515,N_2573,N_2908);
nand U3516 (N_3516,N_2066,N_2136);
nand U3517 (N_3517,N_2189,N_2209);
nor U3518 (N_3518,N_2165,N_2325);
nand U3519 (N_3519,N_2165,N_2512);
nor U3520 (N_3520,N_2131,N_2265);
or U3521 (N_3521,N_2004,N_2515);
nor U3522 (N_3522,N_2643,N_2472);
and U3523 (N_3523,N_2318,N_2477);
and U3524 (N_3524,N_2881,N_2039);
nand U3525 (N_3525,N_2021,N_2375);
and U3526 (N_3526,N_2095,N_2983);
or U3527 (N_3527,N_2845,N_2028);
nor U3528 (N_3528,N_2774,N_2608);
or U3529 (N_3529,N_2053,N_2270);
or U3530 (N_3530,N_2958,N_2193);
nor U3531 (N_3531,N_2363,N_2613);
and U3532 (N_3532,N_2712,N_2622);
nand U3533 (N_3533,N_2409,N_2961);
nor U3534 (N_3534,N_2157,N_2169);
nor U3535 (N_3535,N_2648,N_2721);
nand U3536 (N_3536,N_2120,N_2160);
or U3537 (N_3537,N_2035,N_2427);
nand U3538 (N_3538,N_2318,N_2279);
nand U3539 (N_3539,N_2156,N_2828);
nor U3540 (N_3540,N_2463,N_2621);
and U3541 (N_3541,N_2695,N_2529);
or U3542 (N_3542,N_2878,N_2488);
nand U3543 (N_3543,N_2578,N_2745);
nor U3544 (N_3544,N_2380,N_2711);
or U3545 (N_3545,N_2465,N_2362);
and U3546 (N_3546,N_2013,N_2243);
and U3547 (N_3547,N_2141,N_2767);
and U3548 (N_3548,N_2004,N_2424);
nand U3549 (N_3549,N_2057,N_2024);
or U3550 (N_3550,N_2126,N_2016);
nand U3551 (N_3551,N_2268,N_2691);
nor U3552 (N_3552,N_2877,N_2429);
and U3553 (N_3553,N_2138,N_2453);
nor U3554 (N_3554,N_2886,N_2456);
nor U3555 (N_3555,N_2117,N_2464);
and U3556 (N_3556,N_2357,N_2586);
and U3557 (N_3557,N_2244,N_2547);
and U3558 (N_3558,N_2359,N_2030);
nor U3559 (N_3559,N_2010,N_2721);
nand U3560 (N_3560,N_2165,N_2579);
nand U3561 (N_3561,N_2724,N_2578);
and U3562 (N_3562,N_2682,N_2756);
nand U3563 (N_3563,N_2420,N_2638);
or U3564 (N_3564,N_2094,N_2633);
nand U3565 (N_3565,N_2534,N_2614);
nor U3566 (N_3566,N_2067,N_2226);
or U3567 (N_3567,N_2044,N_2604);
nand U3568 (N_3568,N_2388,N_2909);
xor U3569 (N_3569,N_2547,N_2635);
nor U3570 (N_3570,N_2550,N_2196);
and U3571 (N_3571,N_2935,N_2256);
nor U3572 (N_3572,N_2003,N_2292);
or U3573 (N_3573,N_2062,N_2019);
or U3574 (N_3574,N_2339,N_2283);
nor U3575 (N_3575,N_2432,N_2095);
nand U3576 (N_3576,N_2657,N_2882);
nand U3577 (N_3577,N_2516,N_2624);
or U3578 (N_3578,N_2571,N_2490);
xnor U3579 (N_3579,N_2127,N_2748);
nand U3580 (N_3580,N_2736,N_2026);
nor U3581 (N_3581,N_2279,N_2016);
or U3582 (N_3582,N_2263,N_2225);
xor U3583 (N_3583,N_2133,N_2676);
or U3584 (N_3584,N_2315,N_2870);
nor U3585 (N_3585,N_2461,N_2229);
or U3586 (N_3586,N_2676,N_2532);
and U3587 (N_3587,N_2959,N_2043);
nor U3588 (N_3588,N_2319,N_2759);
and U3589 (N_3589,N_2771,N_2495);
xnor U3590 (N_3590,N_2079,N_2471);
nor U3591 (N_3591,N_2829,N_2417);
or U3592 (N_3592,N_2718,N_2473);
nor U3593 (N_3593,N_2967,N_2680);
or U3594 (N_3594,N_2493,N_2833);
or U3595 (N_3595,N_2924,N_2611);
nor U3596 (N_3596,N_2606,N_2221);
nand U3597 (N_3597,N_2319,N_2440);
nand U3598 (N_3598,N_2735,N_2580);
and U3599 (N_3599,N_2285,N_2935);
and U3600 (N_3600,N_2757,N_2564);
nand U3601 (N_3601,N_2067,N_2095);
nor U3602 (N_3602,N_2920,N_2921);
and U3603 (N_3603,N_2570,N_2483);
nand U3604 (N_3604,N_2631,N_2860);
nand U3605 (N_3605,N_2396,N_2009);
nor U3606 (N_3606,N_2523,N_2602);
nor U3607 (N_3607,N_2988,N_2301);
nand U3608 (N_3608,N_2179,N_2431);
nor U3609 (N_3609,N_2804,N_2774);
and U3610 (N_3610,N_2307,N_2628);
nand U3611 (N_3611,N_2755,N_2813);
and U3612 (N_3612,N_2403,N_2020);
nand U3613 (N_3613,N_2506,N_2412);
nor U3614 (N_3614,N_2744,N_2861);
or U3615 (N_3615,N_2003,N_2045);
nor U3616 (N_3616,N_2796,N_2730);
nand U3617 (N_3617,N_2745,N_2630);
nor U3618 (N_3618,N_2858,N_2966);
nand U3619 (N_3619,N_2470,N_2087);
or U3620 (N_3620,N_2132,N_2844);
and U3621 (N_3621,N_2966,N_2082);
nor U3622 (N_3622,N_2848,N_2891);
nand U3623 (N_3623,N_2372,N_2601);
nor U3624 (N_3624,N_2367,N_2820);
or U3625 (N_3625,N_2281,N_2728);
nand U3626 (N_3626,N_2530,N_2323);
nor U3627 (N_3627,N_2415,N_2703);
nor U3628 (N_3628,N_2871,N_2463);
and U3629 (N_3629,N_2385,N_2813);
and U3630 (N_3630,N_2842,N_2977);
nand U3631 (N_3631,N_2822,N_2701);
nor U3632 (N_3632,N_2440,N_2607);
or U3633 (N_3633,N_2619,N_2843);
nand U3634 (N_3634,N_2017,N_2679);
and U3635 (N_3635,N_2873,N_2443);
nor U3636 (N_3636,N_2174,N_2393);
nand U3637 (N_3637,N_2248,N_2108);
nand U3638 (N_3638,N_2128,N_2561);
or U3639 (N_3639,N_2776,N_2691);
nor U3640 (N_3640,N_2478,N_2153);
nand U3641 (N_3641,N_2946,N_2612);
nand U3642 (N_3642,N_2180,N_2782);
nor U3643 (N_3643,N_2392,N_2387);
and U3644 (N_3644,N_2669,N_2458);
nor U3645 (N_3645,N_2528,N_2468);
or U3646 (N_3646,N_2246,N_2540);
nand U3647 (N_3647,N_2702,N_2613);
or U3648 (N_3648,N_2634,N_2829);
or U3649 (N_3649,N_2131,N_2628);
or U3650 (N_3650,N_2820,N_2471);
nor U3651 (N_3651,N_2893,N_2686);
nand U3652 (N_3652,N_2393,N_2944);
nand U3653 (N_3653,N_2230,N_2952);
nor U3654 (N_3654,N_2964,N_2300);
nand U3655 (N_3655,N_2149,N_2872);
nor U3656 (N_3656,N_2561,N_2920);
or U3657 (N_3657,N_2427,N_2520);
or U3658 (N_3658,N_2856,N_2801);
and U3659 (N_3659,N_2192,N_2151);
and U3660 (N_3660,N_2607,N_2632);
nor U3661 (N_3661,N_2577,N_2684);
or U3662 (N_3662,N_2806,N_2244);
nor U3663 (N_3663,N_2035,N_2161);
or U3664 (N_3664,N_2736,N_2527);
and U3665 (N_3665,N_2142,N_2275);
and U3666 (N_3666,N_2249,N_2423);
nor U3667 (N_3667,N_2066,N_2504);
nand U3668 (N_3668,N_2328,N_2710);
nor U3669 (N_3669,N_2343,N_2368);
nor U3670 (N_3670,N_2531,N_2287);
or U3671 (N_3671,N_2667,N_2790);
or U3672 (N_3672,N_2713,N_2560);
and U3673 (N_3673,N_2828,N_2041);
xor U3674 (N_3674,N_2201,N_2640);
nand U3675 (N_3675,N_2176,N_2415);
and U3676 (N_3676,N_2072,N_2258);
nor U3677 (N_3677,N_2503,N_2954);
or U3678 (N_3678,N_2619,N_2988);
or U3679 (N_3679,N_2114,N_2661);
nor U3680 (N_3680,N_2100,N_2005);
and U3681 (N_3681,N_2558,N_2253);
nor U3682 (N_3682,N_2280,N_2112);
and U3683 (N_3683,N_2167,N_2484);
and U3684 (N_3684,N_2684,N_2346);
and U3685 (N_3685,N_2627,N_2769);
or U3686 (N_3686,N_2960,N_2508);
nor U3687 (N_3687,N_2236,N_2704);
nor U3688 (N_3688,N_2204,N_2305);
or U3689 (N_3689,N_2329,N_2591);
nor U3690 (N_3690,N_2145,N_2172);
nor U3691 (N_3691,N_2096,N_2807);
nor U3692 (N_3692,N_2456,N_2118);
and U3693 (N_3693,N_2508,N_2411);
nand U3694 (N_3694,N_2983,N_2669);
or U3695 (N_3695,N_2671,N_2588);
or U3696 (N_3696,N_2637,N_2094);
and U3697 (N_3697,N_2936,N_2483);
nor U3698 (N_3698,N_2707,N_2184);
nor U3699 (N_3699,N_2516,N_2282);
and U3700 (N_3700,N_2581,N_2197);
and U3701 (N_3701,N_2692,N_2026);
or U3702 (N_3702,N_2353,N_2629);
nand U3703 (N_3703,N_2531,N_2699);
or U3704 (N_3704,N_2704,N_2240);
or U3705 (N_3705,N_2051,N_2188);
nor U3706 (N_3706,N_2461,N_2652);
nand U3707 (N_3707,N_2914,N_2572);
nor U3708 (N_3708,N_2091,N_2896);
or U3709 (N_3709,N_2799,N_2379);
nand U3710 (N_3710,N_2707,N_2776);
nand U3711 (N_3711,N_2316,N_2404);
or U3712 (N_3712,N_2369,N_2324);
nand U3713 (N_3713,N_2619,N_2484);
nor U3714 (N_3714,N_2906,N_2159);
or U3715 (N_3715,N_2172,N_2684);
and U3716 (N_3716,N_2505,N_2103);
nand U3717 (N_3717,N_2391,N_2628);
nand U3718 (N_3718,N_2888,N_2418);
nand U3719 (N_3719,N_2083,N_2690);
nand U3720 (N_3720,N_2340,N_2004);
nand U3721 (N_3721,N_2261,N_2454);
or U3722 (N_3722,N_2625,N_2963);
nor U3723 (N_3723,N_2511,N_2778);
nor U3724 (N_3724,N_2719,N_2173);
nor U3725 (N_3725,N_2097,N_2686);
or U3726 (N_3726,N_2859,N_2739);
or U3727 (N_3727,N_2275,N_2144);
nand U3728 (N_3728,N_2075,N_2957);
and U3729 (N_3729,N_2815,N_2401);
nor U3730 (N_3730,N_2961,N_2482);
or U3731 (N_3731,N_2980,N_2293);
and U3732 (N_3732,N_2012,N_2610);
or U3733 (N_3733,N_2962,N_2540);
and U3734 (N_3734,N_2028,N_2968);
nand U3735 (N_3735,N_2510,N_2042);
or U3736 (N_3736,N_2976,N_2582);
and U3737 (N_3737,N_2804,N_2464);
nor U3738 (N_3738,N_2035,N_2148);
nand U3739 (N_3739,N_2754,N_2239);
or U3740 (N_3740,N_2184,N_2190);
and U3741 (N_3741,N_2219,N_2408);
or U3742 (N_3742,N_2196,N_2240);
and U3743 (N_3743,N_2314,N_2777);
or U3744 (N_3744,N_2450,N_2811);
and U3745 (N_3745,N_2210,N_2991);
and U3746 (N_3746,N_2922,N_2351);
and U3747 (N_3747,N_2801,N_2649);
nor U3748 (N_3748,N_2060,N_2557);
nor U3749 (N_3749,N_2766,N_2416);
nand U3750 (N_3750,N_2258,N_2767);
nand U3751 (N_3751,N_2164,N_2933);
or U3752 (N_3752,N_2696,N_2056);
nor U3753 (N_3753,N_2502,N_2408);
nor U3754 (N_3754,N_2421,N_2943);
nor U3755 (N_3755,N_2282,N_2296);
and U3756 (N_3756,N_2782,N_2486);
xor U3757 (N_3757,N_2650,N_2765);
nor U3758 (N_3758,N_2099,N_2274);
and U3759 (N_3759,N_2685,N_2925);
and U3760 (N_3760,N_2816,N_2293);
or U3761 (N_3761,N_2479,N_2029);
and U3762 (N_3762,N_2018,N_2032);
or U3763 (N_3763,N_2618,N_2227);
nor U3764 (N_3764,N_2266,N_2965);
nor U3765 (N_3765,N_2807,N_2375);
or U3766 (N_3766,N_2705,N_2877);
and U3767 (N_3767,N_2626,N_2552);
and U3768 (N_3768,N_2547,N_2684);
nand U3769 (N_3769,N_2913,N_2685);
nor U3770 (N_3770,N_2733,N_2646);
nand U3771 (N_3771,N_2829,N_2049);
and U3772 (N_3772,N_2230,N_2783);
and U3773 (N_3773,N_2216,N_2660);
nand U3774 (N_3774,N_2732,N_2150);
nand U3775 (N_3775,N_2147,N_2117);
or U3776 (N_3776,N_2265,N_2679);
nand U3777 (N_3777,N_2536,N_2801);
or U3778 (N_3778,N_2449,N_2278);
nand U3779 (N_3779,N_2069,N_2848);
or U3780 (N_3780,N_2493,N_2200);
nor U3781 (N_3781,N_2028,N_2704);
nand U3782 (N_3782,N_2345,N_2504);
nand U3783 (N_3783,N_2615,N_2181);
or U3784 (N_3784,N_2742,N_2786);
nand U3785 (N_3785,N_2703,N_2067);
nor U3786 (N_3786,N_2648,N_2129);
xnor U3787 (N_3787,N_2580,N_2292);
or U3788 (N_3788,N_2767,N_2147);
and U3789 (N_3789,N_2830,N_2532);
and U3790 (N_3790,N_2125,N_2877);
or U3791 (N_3791,N_2638,N_2240);
or U3792 (N_3792,N_2778,N_2889);
and U3793 (N_3793,N_2413,N_2378);
nor U3794 (N_3794,N_2844,N_2802);
nor U3795 (N_3795,N_2139,N_2250);
nor U3796 (N_3796,N_2556,N_2387);
nor U3797 (N_3797,N_2403,N_2039);
and U3798 (N_3798,N_2060,N_2900);
nor U3799 (N_3799,N_2919,N_2359);
or U3800 (N_3800,N_2306,N_2570);
nor U3801 (N_3801,N_2419,N_2178);
and U3802 (N_3802,N_2054,N_2844);
or U3803 (N_3803,N_2331,N_2283);
or U3804 (N_3804,N_2683,N_2240);
nor U3805 (N_3805,N_2275,N_2672);
or U3806 (N_3806,N_2360,N_2987);
nand U3807 (N_3807,N_2097,N_2117);
nor U3808 (N_3808,N_2547,N_2478);
nand U3809 (N_3809,N_2237,N_2856);
nand U3810 (N_3810,N_2000,N_2540);
nand U3811 (N_3811,N_2665,N_2244);
or U3812 (N_3812,N_2868,N_2533);
nor U3813 (N_3813,N_2330,N_2321);
and U3814 (N_3814,N_2939,N_2055);
or U3815 (N_3815,N_2523,N_2396);
and U3816 (N_3816,N_2222,N_2401);
or U3817 (N_3817,N_2246,N_2864);
nor U3818 (N_3818,N_2364,N_2315);
nor U3819 (N_3819,N_2461,N_2689);
or U3820 (N_3820,N_2691,N_2510);
nand U3821 (N_3821,N_2625,N_2174);
and U3822 (N_3822,N_2158,N_2254);
nor U3823 (N_3823,N_2675,N_2829);
or U3824 (N_3824,N_2689,N_2458);
and U3825 (N_3825,N_2090,N_2341);
nand U3826 (N_3826,N_2172,N_2734);
or U3827 (N_3827,N_2357,N_2127);
nor U3828 (N_3828,N_2528,N_2508);
and U3829 (N_3829,N_2451,N_2326);
or U3830 (N_3830,N_2941,N_2704);
nand U3831 (N_3831,N_2280,N_2191);
and U3832 (N_3832,N_2847,N_2623);
nor U3833 (N_3833,N_2857,N_2023);
nor U3834 (N_3834,N_2732,N_2877);
and U3835 (N_3835,N_2522,N_2834);
and U3836 (N_3836,N_2361,N_2584);
nand U3837 (N_3837,N_2623,N_2751);
nor U3838 (N_3838,N_2818,N_2019);
nand U3839 (N_3839,N_2429,N_2021);
nand U3840 (N_3840,N_2634,N_2811);
and U3841 (N_3841,N_2264,N_2784);
or U3842 (N_3842,N_2128,N_2489);
or U3843 (N_3843,N_2914,N_2100);
or U3844 (N_3844,N_2316,N_2729);
nand U3845 (N_3845,N_2499,N_2335);
nand U3846 (N_3846,N_2023,N_2741);
or U3847 (N_3847,N_2266,N_2867);
and U3848 (N_3848,N_2030,N_2136);
nor U3849 (N_3849,N_2171,N_2626);
and U3850 (N_3850,N_2175,N_2928);
or U3851 (N_3851,N_2112,N_2038);
nand U3852 (N_3852,N_2249,N_2903);
or U3853 (N_3853,N_2718,N_2693);
nor U3854 (N_3854,N_2506,N_2553);
or U3855 (N_3855,N_2659,N_2728);
nor U3856 (N_3856,N_2887,N_2682);
nand U3857 (N_3857,N_2795,N_2445);
or U3858 (N_3858,N_2618,N_2476);
and U3859 (N_3859,N_2401,N_2232);
nand U3860 (N_3860,N_2130,N_2524);
or U3861 (N_3861,N_2589,N_2578);
or U3862 (N_3862,N_2182,N_2882);
and U3863 (N_3863,N_2216,N_2056);
nor U3864 (N_3864,N_2078,N_2119);
and U3865 (N_3865,N_2438,N_2260);
and U3866 (N_3866,N_2427,N_2490);
nand U3867 (N_3867,N_2740,N_2481);
nor U3868 (N_3868,N_2935,N_2436);
and U3869 (N_3869,N_2871,N_2648);
or U3870 (N_3870,N_2443,N_2104);
nor U3871 (N_3871,N_2241,N_2785);
and U3872 (N_3872,N_2219,N_2803);
nand U3873 (N_3873,N_2332,N_2560);
or U3874 (N_3874,N_2425,N_2307);
and U3875 (N_3875,N_2994,N_2764);
or U3876 (N_3876,N_2677,N_2049);
nand U3877 (N_3877,N_2580,N_2991);
nor U3878 (N_3878,N_2804,N_2266);
nor U3879 (N_3879,N_2459,N_2657);
nor U3880 (N_3880,N_2617,N_2396);
and U3881 (N_3881,N_2811,N_2593);
xor U3882 (N_3882,N_2847,N_2148);
or U3883 (N_3883,N_2999,N_2961);
or U3884 (N_3884,N_2972,N_2765);
nand U3885 (N_3885,N_2643,N_2599);
nand U3886 (N_3886,N_2171,N_2340);
nor U3887 (N_3887,N_2878,N_2149);
nand U3888 (N_3888,N_2456,N_2193);
nand U3889 (N_3889,N_2936,N_2951);
nor U3890 (N_3890,N_2043,N_2893);
nor U3891 (N_3891,N_2857,N_2822);
or U3892 (N_3892,N_2695,N_2966);
nand U3893 (N_3893,N_2729,N_2216);
or U3894 (N_3894,N_2154,N_2596);
or U3895 (N_3895,N_2207,N_2526);
and U3896 (N_3896,N_2066,N_2932);
and U3897 (N_3897,N_2502,N_2377);
or U3898 (N_3898,N_2233,N_2495);
nor U3899 (N_3899,N_2546,N_2809);
nor U3900 (N_3900,N_2296,N_2939);
nand U3901 (N_3901,N_2225,N_2511);
and U3902 (N_3902,N_2468,N_2199);
and U3903 (N_3903,N_2102,N_2005);
or U3904 (N_3904,N_2754,N_2447);
or U3905 (N_3905,N_2888,N_2780);
nor U3906 (N_3906,N_2688,N_2640);
nor U3907 (N_3907,N_2820,N_2755);
or U3908 (N_3908,N_2278,N_2880);
or U3909 (N_3909,N_2076,N_2137);
nand U3910 (N_3910,N_2535,N_2052);
and U3911 (N_3911,N_2739,N_2078);
nand U3912 (N_3912,N_2517,N_2894);
or U3913 (N_3913,N_2422,N_2828);
nand U3914 (N_3914,N_2926,N_2936);
nand U3915 (N_3915,N_2847,N_2629);
or U3916 (N_3916,N_2505,N_2820);
and U3917 (N_3917,N_2632,N_2342);
nor U3918 (N_3918,N_2303,N_2097);
nand U3919 (N_3919,N_2122,N_2430);
nand U3920 (N_3920,N_2730,N_2625);
and U3921 (N_3921,N_2751,N_2555);
and U3922 (N_3922,N_2705,N_2610);
nand U3923 (N_3923,N_2817,N_2968);
and U3924 (N_3924,N_2319,N_2249);
nand U3925 (N_3925,N_2881,N_2492);
nand U3926 (N_3926,N_2502,N_2323);
nor U3927 (N_3927,N_2065,N_2772);
nor U3928 (N_3928,N_2389,N_2127);
nand U3929 (N_3929,N_2540,N_2889);
or U3930 (N_3930,N_2743,N_2864);
nand U3931 (N_3931,N_2144,N_2356);
and U3932 (N_3932,N_2569,N_2365);
nor U3933 (N_3933,N_2986,N_2882);
nand U3934 (N_3934,N_2800,N_2739);
nor U3935 (N_3935,N_2196,N_2717);
nor U3936 (N_3936,N_2933,N_2647);
nand U3937 (N_3937,N_2781,N_2879);
or U3938 (N_3938,N_2517,N_2996);
and U3939 (N_3939,N_2200,N_2902);
nor U3940 (N_3940,N_2062,N_2348);
or U3941 (N_3941,N_2891,N_2306);
or U3942 (N_3942,N_2686,N_2464);
nand U3943 (N_3943,N_2172,N_2464);
or U3944 (N_3944,N_2257,N_2692);
nor U3945 (N_3945,N_2652,N_2065);
and U3946 (N_3946,N_2212,N_2414);
or U3947 (N_3947,N_2725,N_2521);
or U3948 (N_3948,N_2156,N_2314);
and U3949 (N_3949,N_2543,N_2252);
and U3950 (N_3950,N_2642,N_2785);
nand U3951 (N_3951,N_2669,N_2740);
or U3952 (N_3952,N_2710,N_2017);
nor U3953 (N_3953,N_2004,N_2630);
nor U3954 (N_3954,N_2172,N_2305);
nand U3955 (N_3955,N_2880,N_2594);
nand U3956 (N_3956,N_2918,N_2727);
nor U3957 (N_3957,N_2334,N_2445);
nand U3958 (N_3958,N_2831,N_2560);
or U3959 (N_3959,N_2120,N_2731);
nor U3960 (N_3960,N_2327,N_2890);
and U3961 (N_3961,N_2914,N_2066);
or U3962 (N_3962,N_2313,N_2496);
or U3963 (N_3963,N_2392,N_2309);
nor U3964 (N_3964,N_2200,N_2639);
and U3965 (N_3965,N_2868,N_2197);
nand U3966 (N_3966,N_2710,N_2248);
or U3967 (N_3967,N_2298,N_2748);
nor U3968 (N_3968,N_2527,N_2983);
or U3969 (N_3969,N_2075,N_2242);
or U3970 (N_3970,N_2297,N_2711);
or U3971 (N_3971,N_2665,N_2483);
or U3972 (N_3972,N_2233,N_2214);
or U3973 (N_3973,N_2538,N_2447);
nand U3974 (N_3974,N_2837,N_2056);
nor U3975 (N_3975,N_2129,N_2238);
nor U3976 (N_3976,N_2271,N_2673);
nor U3977 (N_3977,N_2405,N_2558);
and U3978 (N_3978,N_2557,N_2153);
or U3979 (N_3979,N_2440,N_2770);
and U3980 (N_3980,N_2068,N_2448);
nor U3981 (N_3981,N_2798,N_2670);
nand U3982 (N_3982,N_2843,N_2764);
nand U3983 (N_3983,N_2537,N_2078);
nor U3984 (N_3984,N_2061,N_2420);
or U3985 (N_3985,N_2555,N_2233);
and U3986 (N_3986,N_2182,N_2541);
nor U3987 (N_3987,N_2151,N_2093);
or U3988 (N_3988,N_2153,N_2928);
and U3989 (N_3989,N_2632,N_2120);
nor U3990 (N_3990,N_2635,N_2131);
nand U3991 (N_3991,N_2485,N_2669);
nand U3992 (N_3992,N_2313,N_2638);
nand U3993 (N_3993,N_2081,N_2442);
or U3994 (N_3994,N_2137,N_2922);
or U3995 (N_3995,N_2659,N_2368);
and U3996 (N_3996,N_2940,N_2387);
or U3997 (N_3997,N_2286,N_2631);
and U3998 (N_3998,N_2639,N_2076);
nor U3999 (N_3999,N_2680,N_2874);
nor U4000 (N_4000,N_3804,N_3172);
or U4001 (N_4001,N_3671,N_3328);
nor U4002 (N_4002,N_3104,N_3673);
nor U4003 (N_4003,N_3806,N_3921);
and U4004 (N_4004,N_3748,N_3811);
or U4005 (N_4005,N_3600,N_3091);
and U4006 (N_4006,N_3959,N_3621);
nand U4007 (N_4007,N_3617,N_3374);
nand U4008 (N_4008,N_3335,N_3842);
or U4009 (N_4009,N_3611,N_3247);
nor U4010 (N_4010,N_3991,N_3119);
nand U4011 (N_4011,N_3239,N_3730);
nand U4012 (N_4012,N_3325,N_3356);
nor U4013 (N_4013,N_3776,N_3114);
nand U4014 (N_4014,N_3364,N_3565);
or U4015 (N_4015,N_3296,N_3917);
nand U4016 (N_4016,N_3821,N_3362);
nor U4017 (N_4017,N_3238,N_3805);
nand U4018 (N_4018,N_3376,N_3354);
nor U4019 (N_4019,N_3420,N_3851);
nand U4020 (N_4020,N_3942,N_3192);
or U4021 (N_4021,N_3778,N_3840);
nand U4022 (N_4022,N_3297,N_3405);
nor U4023 (N_4023,N_3200,N_3225);
nand U4024 (N_4024,N_3530,N_3594);
and U4025 (N_4025,N_3483,N_3843);
or U4026 (N_4026,N_3450,N_3021);
nor U4027 (N_4027,N_3359,N_3146);
or U4028 (N_4028,N_3886,N_3504);
or U4029 (N_4029,N_3694,N_3506);
or U4030 (N_4030,N_3198,N_3844);
or U4031 (N_4031,N_3222,N_3683);
nor U4032 (N_4032,N_3976,N_3800);
nor U4033 (N_4033,N_3363,N_3705);
nor U4034 (N_4034,N_3562,N_3144);
nor U4035 (N_4035,N_3478,N_3718);
nand U4036 (N_4036,N_3260,N_3466);
and U4037 (N_4037,N_3881,N_3672);
nand U4038 (N_4038,N_3603,N_3217);
or U4039 (N_4039,N_3625,N_3221);
or U4040 (N_4040,N_3722,N_3736);
nor U4041 (N_4041,N_3532,N_3677);
and U4042 (N_4042,N_3922,N_3717);
nor U4043 (N_4043,N_3801,N_3965);
or U4044 (N_4044,N_3001,N_3946);
nor U4045 (N_4045,N_3610,N_3524);
and U4046 (N_4046,N_3556,N_3659);
nand U4047 (N_4047,N_3589,N_3243);
or U4048 (N_4048,N_3505,N_3387);
and U4049 (N_4049,N_3518,N_3174);
nor U4050 (N_4050,N_3384,N_3095);
and U4051 (N_4051,N_3162,N_3230);
nand U4052 (N_4052,N_3510,N_3007);
or U4053 (N_4053,N_3111,N_3741);
and U4054 (N_4054,N_3866,N_3960);
nand U4055 (N_4055,N_3400,N_3978);
nand U4056 (N_4056,N_3915,N_3094);
nand U4057 (N_4057,N_3955,N_3645);
nand U4058 (N_4058,N_3861,N_3334);
and U4059 (N_4059,N_3947,N_3244);
nand U4060 (N_4060,N_3381,N_3477);
nor U4061 (N_4061,N_3775,N_3495);
nor U4062 (N_4062,N_3046,N_3008);
nor U4063 (N_4063,N_3907,N_3648);
nand U4064 (N_4064,N_3852,N_3912);
nor U4065 (N_4065,N_3352,N_3981);
and U4066 (N_4066,N_3267,N_3544);
or U4067 (N_4067,N_3612,N_3409);
and U4068 (N_4068,N_3952,N_3257);
nor U4069 (N_4069,N_3427,N_3263);
nor U4070 (N_4070,N_3256,N_3794);
nand U4071 (N_4071,N_3576,N_3768);
nor U4072 (N_4072,N_3487,N_3330);
nand U4073 (N_4073,N_3874,N_3536);
nor U4074 (N_4074,N_3754,N_3807);
nand U4075 (N_4075,N_3925,N_3766);
and U4076 (N_4076,N_3074,N_3780);
xnor U4077 (N_4077,N_3398,N_3106);
nor U4078 (N_4078,N_3879,N_3786);
nor U4079 (N_4079,N_3446,N_3460);
nor U4080 (N_4080,N_3469,N_3595);
nor U4081 (N_4081,N_3697,N_3346);
nand U4082 (N_4082,N_3023,N_3666);
and U4083 (N_4083,N_3945,N_3178);
nand U4084 (N_4084,N_3644,N_3854);
or U4085 (N_4085,N_3411,N_3143);
nor U4086 (N_4086,N_3931,N_3517);
nand U4087 (N_4087,N_3867,N_3785);
and U4088 (N_4088,N_3492,N_3846);
and U4089 (N_4089,N_3079,N_3231);
or U4090 (N_4090,N_3739,N_3509);
and U4091 (N_4091,N_3097,N_3549);
and U4092 (N_4092,N_3271,N_3077);
and U4093 (N_4093,N_3122,N_3120);
nor U4094 (N_4094,N_3541,N_3326);
or U4095 (N_4095,N_3015,N_3216);
nor U4096 (N_4096,N_3289,N_3215);
nor U4097 (N_4097,N_3848,N_3656);
nand U4098 (N_4098,N_3660,N_3132);
nor U4099 (N_4099,N_3455,N_3447);
nor U4100 (N_4100,N_3641,N_3634);
and U4101 (N_4101,N_3068,N_3784);
nand U4102 (N_4102,N_3553,N_3471);
and U4103 (N_4103,N_3745,N_3966);
and U4104 (N_4104,N_3485,N_3017);
or U4105 (N_4105,N_3674,N_3304);
or U4106 (N_4106,N_3397,N_3164);
nor U4107 (N_4107,N_3484,N_3278);
and U4108 (N_4108,N_3570,N_3926);
nor U4109 (N_4109,N_3252,N_3935);
and U4110 (N_4110,N_3474,N_3668);
nand U4111 (N_4111,N_3615,N_3614);
nand U4112 (N_4112,N_3072,N_3743);
and U4113 (N_4113,N_3712,N_3368);
or U4114 (N_4114,N_3765,N_3961);
nor U4115 (N_4115,N_3512,N_3708);
nor U4116 (N_4116,N_3526,N_3853);
nor U4117 (N_4117,N_3761,N_3317);
or U4118 (N_4118,N_3457,N_3949);
and U4119 (N_4119,N_3914,N_3431);
or U4120 (N_4120,N_3451,N_3151);
or U4121 (N_4121,N_3987,N_3756);
nor U4122 (N_4122,N_3859,N_3901);
nand U4123 (N_4123,N_3191,N_3481);
or U4124 (N_4124,N_3895,N_3695);
and U4125 (N_4125,N_3378,N_3386);
nor U4126 (N_4126,N_3994,N_3070);
or U4127 (N_4127,N_3419,N_3041);
nor U4128 (N_4128,N_3054,N_3274);
nand U4129 (N_4129,N_3607,N_3664);
or U4130 (N_4130,N_3031,N_3270);
or U4131 (N_4131,N_3599,N_3577);
nor U4132 (N_4132,N_3367,N_3004);
nor U4133 (N_4133,N_3489,N_3803);
nor U4134 (N_4134,N_3989,N_3442);
and U4135 (N_4135,N_3219,N_3875);
and U4136 (N_4136,N_3788,N_3878);
and U4137 (N_4137,N_3266,N_3284);
nor U4138 (N_4138,N_3321,N_3944);
xor U4139 (N_4139,N_3196,N_3643);
and U4140 (N_4140,N_3033,N_3308);
or U4141 (N_4141,N_3262,N_3968);
and U4142 (N_4142,N_3523,N_3189);
or U4143 (N_4143,N_3623,N_3099);
or U4144 (N_4144,N_3402,N_3578);
nor U4145 (N_4145,N_3019,N_3676);
and U4146 (N_4146,N_3793,N_3691);
or U4147 (N_4147,N_3444,N_3721);
or U4148 (N_4148,N_3531,N_3349);
or U4149 (N_4149,N_3476,N_3956);
nor U4150 (N_4150,N_3201,N_3105);
nand U4151 (N_4151,N_3566,N_3662);
nand U4152 (N_4152,N_3314,N_3865);
and U4153 (N_4153,N_3085,N_3294);
nand U4154 (N_4154,N_3388,N_3628);
nand U4155 (N_4155,N_3288,N_3665);
nor U4156 (N_4156,N_3302,N_3109);
or U4157 (N_4157,N_3205,N_3439);
nor U4158 (N_4158,N_3626,N_3351);
nand U4159 (N_4159,N_3064,N_3152);
nor U4160 (N_4160,N_3924,N_3995);
nand U4161 (N_4161,N_3988,N_3930);
and U4162 (N_4162,N_3604,N_3060);
and U4163 (N_4163,N_3096,N_3018);
xnor U4164 (N_4164,N_3501,N_3579);
and U4165 (N_4165,N_3605,N_3592);
nand U4166 (N_4166,N_3882,N_3424);
nand U4167 (N_4167,N_3365,N_3908);
or U4168 (N_4168,N_3430,N_3309);
nor U4169 (N_4169,N_3713,N_3796);
nand U4170 (N_4170,N_3860,N_3893);
nand U4171 (N_4171,N_3627,N_3188);
nand U4172 (N_4172,N_3048,N_3682);
nand U4173 (N_4173,N_3134,N_3598);
or U4174 (N_4174,N_3343,N_3909);
or U4175 (N_4175,N_3287,N_3993);
nor U4176 (N_4176,N_3214,N_3732);
nand U4177 (N_4177,N_3437,N_3724);
nor U4178 (N_4178,N_3468,N_3283);
nand U4179 (N_4179,N_3902,N_3417);
nand U4180 (N_4180,N_3453,N_3654);
nor U4181 (N_4181,N_3957,N_3183);
and U4182 (N_4182,N_3830,N_3539);
or U4183 (N_4183,N_3783,N_3373);
and U4184 (N_4184,N_3515,N_3696);
and U4185 (N_4185,N_3273,N_3903);
or U4186 (N_4186,N_3080,N_3160);
nor U4187 (N_4187,N_3226,N_3000);
nor U4188 (N_4188,N_3552,N_3422);
or U4189 (N_4189,N_3651,N_3452);
and U4190 (N_4190,N_3545,N_3876);
nand U4191 (N_4191,N_3781,N_3371);
nor U4192 (N_4192,N_3503,N_3449);
and U4193 (N_4193,N_3818,N_3149);
and U4194 (N_4194,N_3202,N_3413);
or U4195 (N_4195,N_3850,N_3832);
xor U4196 (N_4196,N_3138,N_3891);
nand U4197 (N_4197,N_3954,N_3538);
nor U4198 (N_4198,N_3631,N_3207);
nor U4199 (N_4199,N_3958,N_3224);
nor U4200 (N_4200,N_3797,N_3281);
nor U4201 (N_4201,N_3382,N_3653);
nand U4202 (N_4202,N_3573,N_3734);
nand U4203 (N_4203,N_3337,N_3986);
nor U4204 (N_4204,N_3035,N_3084);
or U4205 (N_4205,N_3435,N_3974);
nand U4206 (N_4206,N_3764,N_3689);
nor U4207 (N_4207,N_3999,N_3970);
nor U4208 (N_4208,N_3458,N_3277);
and U4209 (N_4209,N_3575,N_3155);
or U4210 (N_4210,N_3596,N_3749);
nor U4211 (N_4211,N_3904,N_3779);
or U4212 (N_4212,N_3475,N_3066);
or U4213 (N_4213,N_3341,N_3153);
nand U4214 (N_4214,N_3300,N_3928);
nand U4215 (N_4215,N_3632,N_3649);
and U4216 (N_4216,N_3480,N_3496);
or U4217 (N_4217,N_3147,N_3071);
and U4218 (N_4218,N_3586,N_3923);
nand U4219 (N_4219,N_3332,N_3898);
and U4220 (N_4220,N_3385,N_3310);
or U4221 (N_4221,N_3513,N_3112);
and U4222 (N_4222,N_3655,N_3900);
and U4223 (N_4223,N_3150,N_3839);
nand U4224 (N_4224,N_3107,N_3440);
nand U4225 (N_4225,N_3003,N_3434);
or U4226 (N_4226,N_3208,N_3522);
and U4227 (N_4227,N_3939,N_3009);
nor U4228 (N_4228,N_3264,N_3050);
nand U4229 (N_4229,N_3175,N_3295);
or U4230 (N_4230,N_3199,N_3103);
nor U4231 (N_4231,N_3421,N_3519);
and U4232 (N_4232,N_3311,N_3640);
and U4233 (N_4233,N_3407,N_3809);
or U4234 (N_4234,N_3168,N_3681);
and U4235 (N_4235,N_3529,N_3158);
and U4236 (N_4236,N_3789,N_3973);
and U4237 (N_4237,N_3657,N_3353);
nand U4238 (N_4238,N_3248,N_3316);
and U4239 (N_4239,N_3011,N_3992);
nand U4240 (N_4240,N_3241,N_3312);
nand U4241 (N_4241,N_3240,N_3772);
and U4242 (N_4242,N_3456,N_3203);
and U4243 (N_4243,N_3318,N_3763);
nand U4244 (N_4244,N_3652,N_3377);
nand U4245 (N_4245,N_3838,N_3045);
and U4246 (N_4246,N_3165,N_3129);
nand U4247 (N_4247,N_3620,N_3030);
nand U4248 (N_4248,N_3616,N_3752);
and U4249 (N_4249,N_3394,N_3016);
or U4250 (N_4250,N_3024,N_3885);
or U4251 (N_4251,N_3299,N_3227);
nor U4252 (N_4252,N_3428,N_3380);
or U4253 (N_4253,N_3497,N_3771);
and U4254 (N_4254,N_3889,N_3005);
or U4255 (N_4255,N_3498,N_3507);
xor U4256 (N_4256,N_3344,N_3193);
and U4257 (N_4257,N_3292,N_3719);
nand U4258 (N_4258,N_3395,N_3327);
nor U4259 (N_4259,N_3399,N_3322);
or U4260 (N_4260,N_3290,N_3044);
nor U4261 (N_4261,N_3790,N_3727);
and U4262 (N_4262,N_3494,N_3379);
xor U4263 (N_4263,N_3213,N_3823);
nor U4264 (N_4264,N_3361,N_3233);
nor U4265 (N_4265,N_3390,N_3829);
nand U4266 (N_4266,N_3675,N_3305);
or U4267 (N_4267,N_3116,N_3569);
nor U4268 (N_4268,N_3769,N_3658);
nand U4269 (N_4269,N_3454,N_3688);
nor U4270 (N_4270,N_3306,N_3169);
or U4271 (N_4271,N_3985,N_3819);
nor U4272 (N_4272,N_3602,N_3619);
nand U4273 (N_4273,N_3557,N_3548);
nor U4274 (N_4274,N_3527,N_3459);
nand U4275 (N_4275,N_3740,N_3043);
xor U4276 (N_4276,N_3108,N_3432);
nor U4277 (N_4277,N_3747,N_3093);
nand U4278 (N_4278,N_3661,N_3088);
or U4279 (N_4279,N_3063,N_3342);
and U4280 (N_4280,N_3733,N_3329);
and U4281 (N_4281,N_3511,N_3690);
or U4282 (N_4282,N_3467,N_3971);
and U4283 (N_4283,N_3841,N_3464);
nor U4284 (N_4284,N_3010,N_3156);
nor U4285 (N_4285,N_3246,N_3687);
nor U4286 (N_4286,N_3036,N_3404);
nand U4287 (N_4287,N_3767,N_3593);
and U4288 (N_4288,N_3698,N_3699);
nand U4289 (N_4289,N_3934,N_3177);
or U4290 (N_4290,N_3581,N_3822);
or U4291 (N_4291,N_3237,N_3126);
or U4292 (N_4292,N_3835,N_3117);
nor U4293 (N_4293,N_3462,N_3418);
or U4294 (N_4294,N_3590,N_3037);
nand U4295 (N_4295,N_3190,N_3613);
and U4296 (N_4296,N_3679,N_3731);
nor U4297 (N_4297,N_3194,N_3113);
nor U4298 (N_4298,N_3686,N_3269);
or U4299 (N_4299,N_3555,N_3684);
nor U4300 (N_4300,N_3121,N_3759);
and U4301 (N_4301,N_3574,N_3738);
nor U4302 (N_4302,N_3998,N_3546);
or U4303 (N_4303,N_3067,N_3415);
nand U4304 (N_4304,N_3663,N_3392);
and U4305 (N_4305,N_3836,N_3040);
and U4306 (N_4306,N_3816,N_3642);
and U4307 (N_4307,N_3338,N_3218);
and U4308 (N_4308,N_3187,N_3488);
or U4309 (N_4309,N_3814,N_3052);
nor U4310 (N_4310,N_3167,N_3212);
nand U4311 (N_4311,N_3813,N_3782);
nand U4312 (N_4312,N_3880,N_3090);
or U4313 (N_4313,N_3173,N_3065);
nand U4314 (N_4314,N_3393,N_3209);
and U4315 (N_4315,N_3564,N_3856);
nand U4316 (N_4316,N_3285,N_3597);
or U4317 (N_4317,N_3127,N_3307);
nor U4318 (N_4318,N_3938,N_3086);
nor U4319 (N_4319,N_3022,N_3396);
and U4320 (N_4320,N_3972,N_3375);
and U4321 (N_4321,N_3228,N_3249);
or U4322 (N_4322,N_3825,N_3716);
nor U4323 (N_4323,N_3637,N_3013);
or U4324 (N_4324,N_3268,N_3810);
or U4325 (N_4325,N_3416,N_3056);
nor U4326 (N_4326,N_3251,N_3502);
or U4327 (N_4327,N_3855,N_3936);
nand U4328 (N_4328,N_3824,N_3963);
and U4329 (N_4329,N_3707,N_3558);
or U4330 (N_4330,N_3493,N_3962);
nor U4331 (N_4331,N_3984,N_3331);
nand U4332 (N_4332,N_3834,N_3812);
and U4333 (N_4333,N_3704,N_3533);
and U4334 (N_4334,N_3242,N_3370);
and U4335 (N_4335,N_3758,N_3873);
and U4336 (N_4336,N_3953,N_3608);
nor U4337 (N_4337,N_3014,N_3951);
and U4338 (N_4338,N_3369,N_3516);
nand U4339 (N_4339,N_3943,N_3845);
nand U4340 (N_4340,N_3279,N_3130);
nor U4341 (N_4341,N_3058,N_3723);
nand U4342 (N_4342,N_3142,N_3047);
nor U4343 (N_4343,N_3755,N_3042);
nor U4344 (N_4344,N_3685,N_3123);
nand U4345 (N_4345,N_3906,N_3588);
nand U4346 (N_4346,N_3049,N_3195);
and U4347 (N_4347,N_3061,N_3700);
or U4348 (N_4348,N_3913,N_3884);
or U4349 (N_4349,N_3403,N_3161);
and U4350 (N_4350,N_3787,N_3235);
nor U4351 (N_4351,N_3864,N_3355);
nor U4352 (N_4352,N_3678,N_3583);
nor U4353 (N_4353,N_3870,N_3735);
and U4354 (N_4354,N_3124,N_3982);
or U4355 (N_4355,N_3791,N_3537);
and U4356 (N_4356,N_3892,N_3975);
or U4357 (N_4357,N_3115,N_3486);
nand U4358 (N_4358,N_3350,N_3443);
nand U4359 (N_4359,N_3647,N_3750);
nor U4360 (N_4360,N_3542,N_3896);
nand U4361 (N_4361,N_3171,N_3323);
or U4362 (N_4362,N_3911,N_3265);
nor U4363 (N_4363,N_3983,N_3441);
xor U4364 (N_4364,N_3133,N_3833);
or U4365 (N_4365,N_3345,N_3473);
and U4366 (N_4366,N_3587,N_3639);
nand U4367 (N_4367,N_3919,N_3101);
nor U4368 (N_4368,N_3372,N_3002);
nand U4369 (N_4369,N_3026,N_3157);
or U4370 (N_4370,N_3210,N_3128);
nand U4371 (N_4371,N_3726,N_3820);
or U4372 (N_4372,N_3751,N_3163);
or U4373 (N_4373,N_3087,N_3280);
nand U4374 (N_4374,N_3899,N_3858);
or U4375 (N_4375,N_3720,N_3559);
or U4376 (N_4376,N_3701,N_3039);
and U4377 (N_4377,N_3714,N_3082);
and U4378 (N_4378,N_3897,N_3508);
and U4379 (N_4379,N_3319,N_3358);
or U4380 (N_4380,N_3591,N_3412);
nor U4381 (N_4381,N_3461,N_3561);
and U4382 (N_4382,N_3742,N_3131);
or U4383 (N_4383,N_3336,N_3141);
and U4384 (N_4384,N_3028,N_3470);
xor U4385 (N_4385,N_3872,N_3465);
and U4386 (N_4386,N_3258,N_3990);
nor U4387 (N_4387,N_3932,N_3871);
and U4388 (N_4388,N_3137,N_3706);
nor U4389 (N_4389,N_3229,N_3827);
and U4390 (N_4390,N_3702,N_3646);
or U4391 (N_4391,N_3737,N_3159);
nand U4392 (N_4392,N_3948,N_3996);
or U4393 (N_4393,N_3680,N_3798);
nor U4394 (N_4394,N_3560,N_3521);
and U4395 (N_4395,N_3291,N_3964);
nor U4396 (N_4396,N_3525,N_3633);
or U4397 (N_4397,N_3206,N_3831);
nand U4398 (N_4398,N_3282,N_3933);
or U4399 (N_4399,N_3298,N_3499);
and U4400 (N_4400,N_3448,N_3012);
nand U4401 (N_4401,N_3918,N_3170);
nand U4402 (N_4402,N_3426,N_3715);
or U4403 (N_4403,N_3979,N_3083);
and U4404 (N_4404,N_3053,N_3554);
nor U4405 (N_4405,N_3550,N_3606);
nand U4406 (N_4406,N_3223,N_3757);
nor U4407 (N_4407,N_3937,N_3255);
and U4408 (N_4408,N_3941,N_3808);
or U4409 (N_4409,N_3629,N_3261);
or U4410 (N_4410,N_3463,N_3940);
nor U4411 (N_4411,N_3630,N_3069);
and U4412 (N_4412,N_3601,N_3006);
or U4413 (N_4413,N_3092,N_3817);
and U4414 (N_4414,N_3073,N_3910);
or U4415 (N_4415,N_3275,N_3916);
and U4416 (N_4416,N_3760,N_3650);
nor U4417 (N_4417,N_3883,N_3245);
and U4418 (N_4418,N_3792,N_3770);
nand U4419 (N_4419,N_3746,N_3089);
and U4420 (N_4420,N_3977,N_3773);
or U4421 (N_4421,N_3204,N_3032);
nand U4422 (N_4422,N_3389,N_3181);
nor U4423 (N_4423,N_3410,N_3877);
nand U4424 (N_4424,N_3472,N_3479);
or U4425 (N_4425,N_3980,N_3967);
nor U4426 (N_4426,N_3888,N_3445);
nand U4427 (N_4427,N_3847,N_3391);
or U4428 (N_4428,N_3815,N_3438);
and U4429 (N_4429,N_3837,N_3849);
and U4430 (N_4430,N_3176,N_3366);
nor U4431 (N_4431,N_3692,N_3585);
nor U4432 (N_4432,N_3076,N_3075);
nand U4433 (N_4433,N_3693,N_3051);
or U4434 (N_4434,N_3333,N_3535);
and U4435 (N_4435,N_3857,N_3638);
nand U4436 (N_4436,N_3211,N_3669);
or U4437 (N_4437,N_3055,N_3868);
or U4438 (N_4438,N_3293,N_3324);
and U4439 (N_4439,N_3154,N_3250);
or U4440 (N_4440,N_3762,N_3140);
and U4441 (N_4441,N_3774,N_3711);
and U4442 (N_4442,N_3185,N_3348);
or U4443 (N_4443,N_3514,N_3490);
and U4444 (N_4444,N_3618,N_3220);
nand U4445 (N_4445,N_3667,N_3034);
and U4446 (N_4446,N_3887,N_3347);
and U4447 (N_4447,N_3166,N_3433);
nor U4448 (N_4448,N_3020,N_3286);
nand U4449 (N_4449,N_3828,N_3062);
and U4450 (N_4450,N_3950,N_3254);
nor U4451 (N_4451,N_3551,N_3777);
or U4452 (N_4452,N_3038,N_3184);
and U4453 (N_4453,N_3025,N_3997);
and U4454 (N_4454,N_3236,N_3744);
or U4455 (N_4455,N_3862,N_3182);
nor U4456 (N_4456,N_3425,N_3572);
nand U4457 (N_4457,N_3423,N_3622);
nand U4458 (N_4458,N_3401,N_3029);
and U4459 (N_4459,N_3582,N_3795);
nor U4460 (N_4460,N_3929,N_3110);
and U4461 (N_4461,N_3315,N_3584);
nor U4462 (N_4462,N_3609,N_3436);
and U4463 (N_4463,N_3118,N_3969);
nor U4464 (N_4464,N_3528,N_3301);
nand U4465 (N_4465,N_3429,N_3753);
or U4466 (N_4466,N_3234,N_3081);
nand U4467 (N_4467,N_3568,N_3135);
nor U4468 (N_4468,N_3179,N_3078);
and U4469 (N_4469,N_3100,N_3920);
nor U4470 (N_4470,N_3408,N_3197);
and U4471 (N_4471,N_3894,N_3547);
and U4472 (N_4472,N_3057,N_3482);
nor U4473 (N_4473,N_3339,N_3563);
or U4474 (N_4474,N_3313,N_3725);
nand U4475 (N_4475,N_3571,N_3580);
nand U4476 (N_4476,N_3728,N_3635);
and U4477 (N_4477,N_3905,N_3272);
and U4478 (N_4478,N_3383,N_3059);
nor U4479 (N_4479,N_3320,N_3276);
nor U4480 (N_4480,N_3232,N_3406);
xor U4481 (N_4481,N_3148,N_3624);
nand U4482 (N_4482,N_3710,N_3180);
or U4483 (N_4483,N_3799,N_3709);
nor U4484 (N_4484,N_3136,N_3125);
and U4485 (N_4485,N_3491,N_3102);
nor U4486 (N_4486,N_3567,N_3543);
nor U4487 (N_4487,N_3098,N_3259);
nor U4488 (N_4488,N_3139,N_3360);
nor U4489 (N_4489,N_3500,N_3703);
nor U4490 (N_4490,N_3357,N_3729);
nand U4491 (N_4491,N_3670,N_3927);
nand U4492 (N_4492,N_3826,N_3869);
nand U4493 (N_4493,N_3340,N_3890);
and U4494 (N_4494,N_3186,N_3520);
and U4495 (N_4495,N_3414,N_3540);
or U4496 (N_4496,N_3145,N_3636);
and U4497 (N_4497,N_3253,N_3027);
nor U4498 (N_4498,N_3303,N_3534);
nor U4499 (N_4499,N_3802,N_3863);
and U4500 (N_4500,N_3152,N_3146);
or U4501 (N_4501,N_3530,N_3601);
nand U4502 (N_4502,N_3997,N_3299);
and U4503 (N_4503,N_3773,N_3711);
and U4504 (N_4504,N_3104,N_3040);
nor U4505 (N_4505,N_3626,N_3490);
nor U4506 (N_4506,N_3802,N_3897);
nand U4507 (N_4507,N_3754,N_3844);
nand U4508 (N_4508,N_3458,N_3083);
nor U4509 (N_4509,N_3334,N_3299);
nand U4510 (N_4510,N_3842,N_3846);
and U4511 (N_4511,N_3965,N_3010);
nand U4512 (N_4512,N_3196,N_3996);
nor U4513 (N_4513,N_3087,N_3832);
nor U4514 (N_4514,N_3046,N_3440);
or U4515 (N_4515,N_3496,N_3162);
nand U4516 (N_4516,N_3450,N_3354);
nand U4517 (N_4517,N_3250,N_3823);
and U4518 (N_4518,N_3807,N_3266);
and U4519 (N_4519,N_3354,N_3715);
nor U4520 (N_4520,N_3255,N_3105);
nor U4521 (N_4521,N_3436,N_3225);
or U4522 (N_4522,N_3469,N_3860);
nor U4523 (N_4523,N_3627,N_3853);
and U4524 (N_4524,N_3610,N_3715);
nand U4525 (N_4525,N_3436,N_3937);
nor U4526 (N_4526,N_3599,N_3653);
nor U4527 (N_4527,N_3591,N_3430);
nand U4528 (N_4528,N_3599,N_3623);
nor U4529 (N_4529,N_3582,N_3751);
or U4530 (N_4530,N_3824,N_3819);
nand U4531 (N_4531,N_3272,N_3812);
nand U4532 (N_4532,N_3335,N_3256);
nand U4533 (N_4533,N_3713,N_3743);
xor U4534 (N_4534,N_3012,N_3770);
and U4535 (N_4535,N_3127,N_3328);
or U4536 (N_4536,N_3547,N_3422);
nor U4537 (N_4537,N_3378,N_3599);
nor U4538 (N_4538,N_3064,N_3949);
or U4539 (N_4539,N_3806,N_3119);
and U4540 (N_4540,N_3321,N_3647);
nor U4541 (N_4541,N_3790,N_3541);
and U4542 (N_4542,N_3290,N_3437);
and U4543 (N_4543,N_3420,N_3973);
and U4544 (N_4544,N_3619,N_3329);
or U4545 (N_4545,N_3866,N_3369);
and U4546 (N_4546,N_3516,N_3536);
or U4547 (N_4547,N_3236,N_3594);
and U4548 (N_4548,N_3690,N_3220);
or U4549 (N_4549,N_3555,N_3694);
nand U4550 (N_4550,N_3944,N_3380);
nand U4551 (N_4551,N_3263,N_3076);
nand U4552 (N_4552,N_3274,N_3420);
or U4553 (N_4553,N_3348,N_3731);
nor U4554 (N_4554,N_3534,N_3726);
or U4555 (N_4555,N_3698,N_3665);
nor U4556 (N_4556,N_3731,N_3439);
or U4557 (N_4557,N_3270,N_3579);
nand U4558 (N_4558,N_3476,N_3417);
nand U4559 (N_4559,N_3495,N_3262);
or U4560 (N_4560,N_3792,N_3553);
nor U4561 (N_4561,N_3944,N_3582);
or U4562 (N_4562,N_3532,N_3997);
xor U4563 (N_4563,N_3311,N_3908);
nand U4564 (N_4564,N_3728,N_3663);
nor U4565 (N_4565,N_3378,N_3662);
nand U4566 (N_4566,N_3191,N_3126);
and U4567 (N_4567,N_3232,N_3448);
nand U4568 (N_4568,N_3548,N_3638);
nor U4569 (N_4569,N_3135,N_3011);
nand U4570 (N_4570,N_3799,N_3029);
nor U4571 (N_4571,N_3661,N_3027);
and U4572 (N_4572,N_3077,N_3621);
nor U4573 (N_4573,N_3567,N_3074);
nor U4574 (N_4574,N_3674,N_3220);
or U4575 (N_4575,N_3617,N_3090);
and U4576 (N_4576,N_3417,N_3545);
or U4577 (N_4577,N_3770,N_3874);
and U4578 (N_4578,N_3019,N_3170);
or U4579 (N_4579,N_3322,N_3335);
nand U4580 (N_4580,N_3881,N_3845);
nand U4581 (N_4581,N_3249,N_3351);
and U4582 (N_4582,N_3610,N_3079);
nor U4583 (N_4583,N_3259,N_3950);
nand U4584 (N_4584,N_3279,N_3975);
nand U4585 (N_4585,N_3191,N_3510);
nand U4586 (N_4586,N_3824,N_3922);
nor U4587 (N_4587,N_3121,N_3784);
nand U4588 (N_4588,N_3306,N_3788);
and U4589 (N_4589,N_3039,N_3166);
nor U4590 (N_4590,N_3969,N_3866);
or U4591 (N_4591,N_3282,N_3184);
and U4592 (N_4592,N_3898,N_3689);
or U4593 (N_4593,N_3179,N_3546);
nand U4594 (N_4594,N_3778,N_3665);
or U4595 (N_4595,N_3852,N_3156);
and U4596 (N_4596,N_3700,N_3617);
nand U4597 (N_4597,N_3408,N_3776);
or U4598 (N_4598,N_3508,N_3643);
or U4599 (N_4599,N_3277,N_3538);
and U4600 (N_4600,N_3946,N_3979);
and U4601 (N_4601,N_3884,N_3728);
and U4602 (N_4602,N_3533,N_3012);
nor U4603 (N_4603,N_3192,N_3104);
nor U4604 (N_4604,N_3515,N_3313);
and U4605 (N_4605,N_3225,N_3016);
and U4606 (N_4606,N_3290,N_3007);
and U4607 (N_4607,N_3944,N_3782);
and U4608 (N_4608,N_3548,N_3091);
xnor U4609 (N_4609,N_3789,N_3463);
and U4610 (N_4610,N_3204,N_3114);
nor U4611 (N_4611,N_3055,N_3001);
and U4612 (N_4612,N_3211,N_3631);
nand U4613 (N_4613,N_3128,N_3268);
nand U4614 (N_4614,N_3091,N_3176);
and U4615 (N_4615,N_3348,N_3009);
or U4616 (N_4616,N_3500,N_3699);
nor U4617 (N_4617,N_3813,N_3089);
or U4618 (N_4618,N_3719,N_3303);
nand U4619 (N_4619,N_3445,N_3900);
nor U4620 (N_4620,N_3992,N_3247);
nor U4621 (N_4621,N_3111,N_3206);
nor U4622 (N_4622,N_3980,N_3135);
nor U4623 (N_4623,N_3645,N_3639);
or U4624 (N_4624,N_3567,N_3958);
nor U4625 (N_4625,N_3239,N_3684);
or U4626 (N_4626,N_3551,N_3966);
nor U4627 (N_4627,N_3558,N_3854);
and U4628 (N_4628,N_3315,N_3425);
or U4629 (N_4629,N_3976,N_3377);
nand U4630 (N_4630,N_3060,N_3618);
and U4631 (N_4631,N_3998,N_3441);
nand U4632 (N_4632,N_3439,N_3334);
nor U4633 (N_4633,N_3166,N_3509);
nand U4634 (N_4634,N_3379,N_3490);
and U4635 (N_4635,N_3989,N_3934);
and U4636 (N_4636,N_3010,N_3834);
or U4637 (N_4637,N_3980,N_3294);
nor U4638 (N_4638,N_3048,N_3487);
nor U4639 (N_4639,N_3590,N_3721);
nand U4640 (N_4640,N_3985,N_3976);
nand U4641 (N_4641,N_3653,N_3725);
or U4642 (N_4642,N_3670,N_3628);
nor U4643 (N_4643,N_3421,N_3838);
nor U4644 (N_4644,N_3628,N_3352);
nor U4645 (N_4645,N_3108,N_3877);
nand U4646 (N_4646,N_3906,N_3581);
nor U4647 (N_4647,N_3437,N_3601);
nor U4648 (N_4648,N_3743,N_3749);
or U4649 (N_4649,N_3976,N_3164);
nand U4650 (N_4650,N_3304,N_3885);
nand U4651 (N_4651,N_3774,N_3208);
nor U4652 (N_4652,N_3239,N_3383);
or U4653 (N_4653,N_3210,N_3380);
nor U4654 (N_4654,N_3813,N_3295);
nor U4655 (N_4655,N_3818,N_3030);
or U4656 (N_4656,N_3597,N_3609);
or U4657 (N_4657,N_3151,N_3677);
or U4658 (N_4658,N_3439,N_3352);
or U4659 (N_4659,N_3574,N_3175);
and U4660 (N_4660,N_3191,N_3885);
nor U4661 (N_4661,N_3707,N_3404);
nor U4662 (N_4662,N_3960,N_3482);
nor U4663 (N_4663,N_3983,N_3994);
and U4664 (N_4664,N_3205,N_3004);
or U4665 (N_4665,N_3224,N_3812);
nand U4666 (N_4666,N_3658,N_3881);
or U4667 (N_4667,N_3415,N_3262);
and U4668 (N_4668,N_3817,N_3512);
nand U4669 (N_4669,N_3210,N_3807);
nand U4670 (N_4670,N_3761,N_3753);
or U4671 (N_4671,N_3947,N_3422);
nor U4672 (N_4672,N_3610,N_3011);
or U4673 (N_4673,N_3399,N_3241);
and U4674 (N_4674,N_3126,N_3159);
nand U4675 (N_4675,N_3612,N_3319);
and U4676 (N_4676,N_3626,N_3818);
or U4677 (N_4677,N_3473,N_3077);
and U4678 (N_4678,N_3997,N_3818);
or U4679 (N_4679,N_3852,N_3421);
xor U4680 (N_4680,N_3673,N_3762);
nor U4681 (N_4681,N_3207,N_3524);
or U4682 (N_4682,N_3811,N_3618);
or U4683 (N_4683,N_3103,N_3976);
and U4684 (N_4684,N_3031,N_3687);
or U4685 (N_4685,N_3025,N_3392);
nand U4686 (N_4686,N_3881,N_3907);
nor U4687 (N_4687,N_3446,N_3184);
nor U4688 (N_4688,N_3341,N_3514);
nor U4689 (N_4689,N_3042,N_3214);
or U4690 (N_4690,N_3521,N_3015);
xnor U4691 (N_4691,N_3529,N_3106);
or U4692 (N_4692,N_3029,N_3357);
or U4693 (N_4693,N_3280,N_3418);
nor U4694 (N_4694,N_3749,N_3660);
and U4695 (N_4695,N_3046,N_3309);
or U4696 (N_4696,N_3405,N_3330);
nand U4697 (N_4697,N_3800,N_3881);
nand U4698 (N_4698,N_3299,N_3901);
and U4699 (N_4699,N_3823,N_3113);
nand U4700 (N_4700,N_3631,N_3135);
nor U4701 (N_4701,N_3361,N_3177);
or U4702 (N_4702,N_3701,N_3316);
or U4703 (N_4703,N_3493,N_3558);
and U4704 (N_4704,N_3419,N_3012);
and U4705 (N_4705,N_3610,N_3560);
or U4706 (N_4706,N_3495,N_3657);
or U4707 (N_4707,N_3116,N_3586);
or U4708 (N_4708,N_3362,N_3001);
nand U4709 (N_4709,N_3326,N_3963);
nand U4710 (N_4710,N_3463,N_3232);
or U4711 (N_4711,N_3254,N_3295);
and U4712 (N_4712,N_3775,N_3550);
nor U4713 (N_4713,N_3173,N_3054);
nor U4714 (N_4714,N_3228,N_3361);
and U4715 (N_4715,N_3384,N_3379);
nor U4716 (N_4716,N_3244,N_3103);
or U4717 (N_4717,N_3024,N_3493);
and U4718 (N_4718,N_3987,N_3830);
and U4719 (N_4719,N_3768,N_3001);
nor U4720 (N_4720,N_3815,N_3700);
and U4721 (N_4721,N_3159,N_3400);
or U4722 (N_4722,N_3533,N_3033);
nand U4723 (N_4723,N_3405,N_3782);
and U4724 (N_4724,N_3794,N_3002);
and U4725 (N_4725,N_3778,N_3431);
nand U4726 (N_4726,N_3882,N_3866);
nor U4727 (N_4727,N_3171,N_3428);
nand U4728 (N_4728,N_3747,N_3847);
nand U4729 (N_4729,N_3975,N_3019);
nor U4730 (N_4730,N_3320,N_3740);
and U4731 (N_4731,N_3590,N_3100);
or U4732 (N_4732,N_3701,N_3583);
and U4733 (N_4733,N_3804,N_3451);
or U4734 (N_4734,N_3638,N_3056);
or U4735 (N_4735,N_3860,N_3273);
and U4736 (N_4736,N_3025,N_3445);
nor U4737 (N_4737,N_3616,N_3853);
nor U4738 (N_4738,N_3046,N_3330);
nand U4739 (N_4739,N_3595,N_3719);
and U4740 (N_4740,N_3877,N_3587);
nand U4741 (N_4741,N_3825,N_3568);
and U4742 (N_4742,N_3628,N_3189);
nand U4743 (N_4743,N_3261,N_3120);
and U4744 (N_4744,N_3508,N_3373);
and U4745 (N_4745,N_3884,N_3549);
xnor U4746 (N_4746,N_3607,N_3243);
and U4747 (N_4747,N_3843,N_3937);
or U4748 (N_4748,N_3422,N_3658);
nor U4749 (N_4749,N_3216,N_3981);
and U4750 (N_4750,N_3870,N_3637);
nand U4751 (N_4751,N_3977,N_3684);
nand U4752 (N_4752,N_3198,N_3793);
nand U4753 (N_4753,N_3420,N_3146);
or U4754 (N_4754,N_3224,N_3657);
and U4755 (N_4755,N_3922,N_3082);
nand U4756 (N_4756,N_3056,N_3182);
and U4757 (N_4757,N_3356,N_3910);
nor U4758 (N_4758,N_3328,N_3195);
nor U4759 (N_4759,N_3230,N_3473);
nor U4760 (N_4760,N_3039,N_3798);
or U4761 (N_4761,N_3082,N_3068);
nor U4762 (N_4762,N_3978,N_3116);
nor U4763 (N_4763,N_3521,N_3738);
nand U4764 (N_4764,N_3735,N_3668);
nor U4765 (N_4765,N_3864,N_3395);
or U4766 (N_4766,N_3495,N_3342);
or U4767 (N_4767,N_3935,N_3855);
nand U4768 (N_4768,N_3101,N_3344);
nand U4769 (N_4769,N_3271,N_3093);
nor U4770 (N_4770,N_3069,N_3852);
nor U4771 (N_4771,N_3330,N_3853);
and U4772 (N_4772,N_3248,N_3966);
and U4773 (N_4773,N_3416,N_3909);
and U4774 (N_4774,N_3269,N_3150);
or U4775 (N_4775,N_3219,N_3197);
nand U4776 (N_4776,N_3883,N_3491);
nor U4777 (N_4777,N_3536,N_3902);
nor U4778 (N_4778,N_3636,N_3369);
and U4779 (N_4779,N_3106,N_3078);
and U4780 (N_4780,N_3290,N_3180);
and U4781 (N_4781,N_3257,N_3116);
nand U4782 (N_4782,N_3267,N_3346);
or U4783 (N_4783,N_3377,N_3793);
nor U4784 (N_4784,N_3603,N_3149);
nor U4785 (N_4785,N_3480,N_3179);
and U4786 (N_4786,N_3106,N_3692);
nor U4787 (N_4787,N_3992,N_3403);
nor U4788 (N_4788,N_3227,N_3843);
nor U4789 (N_4789,N_3492,N_3772);
or U4790 (N_4790,N_3385,N_3615);
nand U4791 (N_4791,N_3391,N_3329);
nor U4792 (N_4792,N_3899,N_3956);
nand U4793 (N_4793,N_3412,N_3467);
nor U4794 (N_4794,N_3242,N_3500);
or U4795 (N_4795,N_3766,N_3116);
nor U4796 (N_4796,N_3299,N_3590);
and U4797 (N_4797,N_3348,N_3991);
or U4798 (N_4798,N_3106,N_3879);
or U4799 (N_4799,N_3462,N_3842);
nor U4800 (N_4800,N_3465,N_3818);
or U4801 (N_4801,N_3731,N_3880);
or U4802 (N_4802,N_3706,N_3427);
nand U4803 (N_4803,N_3791,N_3161);
or U4804 (N_4804,N_3503,N_3008);
and U4805 (N_4805,N_3904,N_3186);
and U4806 (N_4806,N_3087,N_3163);
nor U4807 (N_4807,N_3812,N_3790);
and U4808 (N_4808,N_3297,N_3113);
nand U4809 (N_4809,N_3924,N_3390);
nand U4810 (N_4810,N_3446,N_3594);
nor U4811 (N_4811,N_3446,N_3121);
nand U4812 (N_4812,N_3440,N_3198);
and U4813 (N_4813,N_3487,N_3740);
or U4814 (N_4814,N_3700,N_3144);
or U4815 (N_4815,N_3090,N_3087);
or U4816 (N_4816,N_3740,N_3516);
nand U4817 (N_4817,N_3500,N_3636);
nor U4818 (N_4818,N_3437,N_3665);
nand U4819 (N_4819,N_3156,N_3918);
nor U4820 (N_4820,N_3024,N_3853);
and U4821 (N_4821,N_3630,N_3910);
nor U4822 (N_4822,N_3661,N_3290);
nor U4823 (N_4823,N_3538,N_3461);
nor U4824 (N_4824,N_3106,N_3599);
xor U4825 (N_4825,N_3972,N_3567);
or U4826 (N_4826,N_3357,N_3108);
or U4827 (N_4827,N_3429,N_3395);
or U4828 (N_4828,N_3807,N_3046);
nor U4829 (N_4829,N_3027,N_3717);
and U4830 (N_4830,N_3164,N_3765);
nor U4831 (N_4831,N_3033,N_3077);
nand U4832 (N_4832,N_3336,N_3095);
nand U4833 (N_4833,N_3849,N_3654);
nor U4834 (N_4834,N_3654,N_3278);
or U4835 (N_4835,N_3556,N_3117);
and U4836 (N_4836,N_3032,N_3857);
nand U4837 (N_4837,N_3144,N_3069);
and U4838 (N_4838,N_3586,N_3946);
nor U4839 (N_4839,N_3711,N_3044);
or U4840 (N_4840,N_3496,N_3178);
or U4841 (N_4841,N_3886,N_3149);
or U4842 (N_4842,N_3736,N_3116);
nor U4843 (N_4843,N_3349,N_3731);
nor U4844 (N_4844,N_3133,N_3729);
nand U4845 (N_4845,N_3617,N_3216);
nand U4846 (N_4846,N_3399,N_3642);
nand U4847 (N_4847,N_3564,N_3440);
and U4848 (N_4848,N_3164,N_3564);
nand U4849 (N_4849,N_3168,N_3350);
and U4850 (N_4850,N_3654,N_3047);
or U4851 (N_4851,N_3372,N_3765);
and U4852 (N_4852,N_3812,N_3419);
and U4853 (N_4853,N_3061,N_3454);
nand U4854 (N_4854,N_3633,N_3202);
and U4855 (N_4855,N_3348,N_3547);
and U4856 (N_4856,N_3259,N_3775);
nor U4857 (N_4857,N_3700,N_3955);
nor U4858 (N_4858,N_3806,N_3984);
or U4859 (N_4859,N_3026,N_3284);
and U4860 (N_4860,N_3248,N_3291);
or U4861 (N_4861,N_3389,N_3618);
and U4862 (N_4862,N_3447,N_3266);
and U4863 (N_4863,N_3304,N_3107);
and U4864 (N_4864,N_3974,N_3337);
xor U4865 (N_4865,N_3504,N_3933);
nor U4866 (N_4866,N_3401,N_3333);
nand U4867 (N_4867,N_3167,N_3441);
nor U4868 (N_4868,N_3862,N_3333);
and U4869 (N_4869,N_3139,N_3399);
or U4870 (N_4870,N_3533,N_3886);
or U4871 (N_4871,N_3933,N_3215);
nor U4872 (N_4872,N_3706,N_3388);
nor U4873 (N_4873,N_3874,N_3498);
and U4874 (N_4874,N_3285,N_3779);
and U4875 (N_4875,N_3172,N_3643);
nor U4876 (N_4876,N_3363,N_3055);
and U4877 (N_4877,N_3764,N_3536);
or U4878 (N_4878,N_3979,N_3637);
nor U4879 (N_4879,N_3814,N_3741);
nor U4880 (N_4880,N_3712,N_3143);
nand U4881 (N_4881,N_3258,N_3168);
or U4882 (N_4882,N_3036,N_3014);
or U4883 (N_4883,N_3771,N_3257);
nor U4884 (N_4884,N_3695,N_3629);
nand U4885 (N_4885,N_3261,N_3732);
nand U4886 (N_4886,N_3829,N_3083);
and U4887 (N_4887,N_3268,N_3334);
and U4888 (N_4888,N_3472,N_3888);
nand U4889 (N_4889,N_3921,N_3987);
and U4890 (N_4890,N_3457,N_3099);
nor U4891 (N_4891,N_3759,N_3558);
nand U4892 (N_4892,N_3111,N_3684);
xnor U4893 (N_4893,N_3730,N_3531);
and U4894 (N_4894,N_3797,N_3885);
or U4895 (N_4895,N_3824,N_3964);
or U4896 (N_4896,N_3476,N_3792);
or U4897 (N_4897,N_3161,N_3087);
and U4898 (N_4898,N_3123,N_3775);
nor U4899 (N_4899,N_3755,N_3571);
and U4900 (N_4900,N_3799,N_3579);
and U4901 (N_4901,N_3179,N_3827);
nor U4902 (N_4902,N_3249,N_3606);
nor U4903 (N_4903,N_3185,N_3679);
or U4904 (N_4904,N_3935,N_3669);
and U4905 (N_4905,N_3140,N_3590);
or U4906 (N_4906,N_3386,N_3086);
and U4907 (N_4907,N_3698,N_3798);
nand U4908 (N_4908,N_3041,N_3347);
nand U4909 (N_4909,N_3721,N_3017);
or U4910 (N_4910,N_3264,N_3881);
or U4911 (N_4911,N_3070,N_3703);
nor U4912 (N_4912,N_3493,N_3000);
or U4913 (N_4913,N_3657,N_3785);
and U4914 (N_4914,N_3016,N_3317);
and U4915 (N_4915,N_3381,N_3765);
nand U4916 (N_4916,N_3971,N_3594);
and U4917 (N_4917,N_3584,N_3586);
nand U4918 (N_4918,N_3190,N_3903);
and U4919 (N_4919,N_3087,N_3365);
and U4920 (N_4920,N_3142,N_3497);
or U4921 (N_4921,N_3112,N_3282);
and U4922 (N_4922,N_3671,N_3133);
and U4923 (N_4923,N_3728,N_3890);
nand U4924 (N_4924,N_3480,N_3619);
nor U4925 (N_4925,N_3881,N_3093);
nor U4926 (N_4926,N_3673,N_3819);
or U4927 (N_4927,N_3713,N_3807);
or U4928 (N_4928,N_3841,N_3495);
nand U4929 (N_4929,N_3622,N_3662);
nor U4930 (N_4930,N_3570,N_3478);
and U4931 (N_4931,N_3504,N_3518);
and U4932 (N_4932,N_3021,N_3685);
and U4933 (N_4933,N_3014,N_3073);
nand U4934 (N_4934,N_3283,N_3874);
nor U4935 (N_4935,N_3993,N_3378);
or U4936 (N_4936,N_3180,N_3001);
nor U4937 (N_4937,N_3404,N_3149);
nand U4938 (N_4938,N_3464,N_3220);
or U4939 (N_4939,N_3978,N_3067);
or U4940 (N_4940,N_3309,N_3745);
and U4941 (N_4941,N_3019,N_3006);
or U4942 (N_4942,N_3932,N_3962);
or U4943 (N_4943,N_3871,N_3956);
nand U4944 (N_4944,N_3921,N_3626);
nand U4945 (N_4945,N_3937,N_3174);
and U4946 (N_4946,N_3124,N_3397);
and U4947 (N_4947,N_3242,N_3861);
or U4948 (N_4948,N_3905,N_3872);
and U4949 (N_4949,N_3228,N_3095);
and U4950 (N_4950,N_3716,N_3031);
nand U4951 (N_4951,N_3705,N_3011);
and U4952 (N_4952,N_3653,N_3957);
and U4953 (N_4953,N_3603,N_3510);
nor U4954 (N_4954,N_3120,N_3940);
and U4955 (N_4955,N_3467,N_3205);
nor U4956 (N_4956,N_3529,N_3150);
and U4957 (N_4957,N_3912,N_3590);
or U4958 (N_4958,N_3786,N_3238);
nor U4959 (N_4959,N_3343,N_3819);
nor U4960 (N_4960,N_3226,N_3342);
nor U4961 (N_4961,N_3778,N_3854);
nor U4962 (N_4962,N_3238,N_3044);
nand U4963 (N_4963,N_3754,N_3441);
or U4964 (N_4964,N_3562,N_3881);
and U4965 (N_4965,N_3307,N_3688);
and U4966 (N_4966,N_3183,N_3927);
and U4967 (N_4967,N_3395,N_3212);
nor U4968 (N_4968,N_3477,N_3215);
or U4969 (N_4969,N_3212,N_3024);
and U4970 (N_4970,N_3826,N_3060);
nand U4971 (N_4971,N_3051,N_3562);
nor U4972 (N_4972,N_3698,N_3159);
or U4973 (N_4973,N_3582,N_3838);
and U4974 (N_4974,N_3850,N_3629);
nor U4975 (N_4975,N_3860,N_3843);
nor U4976 (N_4976,N_3840,N_3902);
nand U4977 (N_4977,N_3715,N_3816);
and U4978 (N_4978,N_3607,N_3911);
or U4979 (N_4979,N_3559,N_3262);
nand U4980 (N_4980,N_3680,N_3685);
and U4981 (N_4981,N_3095,N_3706);
nand U4982 (N_4982,N_3391,N_3713);
nor U4983 (N_4983,N_3200,N_3226);
nor U4984 (N_4984,N_3079,N_3212);
and U4985 (N_4985,N_3386,N_3366);
nand U4986 (N_4986,N_3949,N_3422);
nand U4987 (N_4987,N_3392,N_3073);
or U4988 (N_4988,N_3627,N_3446);
or U4989 (N_4989,N_3677,N_3763);
or U4990 (N_4990,N_3070,N_3825);
or U4991 (N_4991,N_3833,N_3395);
and U4992 (N_4992,N_3335,N_3995);
nand U4993 (N_4993,N_3730,N_3801);
xor U4994 (N_4994,N_3460,N_3940);
or U4995 (N_4995,N_3246,N_3106);
and U4996 (N_4996,N_3389,N_3721);
nand U4997 (N_4997,N_3528,N_3950);
nor U4998 (N_4998,N_3354,N_3966);
or U4999 (N_4999,N_3560,N_3252);
nor UO_0 (O_0,N_4709,N_4404);
nor UO_1 (O_1,N_4148,N_4436);
nand UO_2 (O_2,N_4648,N_4592);
nand UO_3 (O_3,N_4261,N_4501);
and UO_4 (O_4,N_4217,N_4460);
nand UO_5 (O_5,N_4800,N_4132);
nor UO_6 (O_6,N_4517,N_4389);
nand UO_7 (O_7,N_4376,N_4854);
nand UO_8 (O_8,N_4933,N_4793);
nand UO_9 (O_9,N_4452,N_4200);
nand UO_10 (O_10,N_4246,N_4368);
or UO_11 (O_11,N_4081,N_4852);
or UO_12 (O_12,N_4659,N_4600);
xor UO_13 (O_13,N_4455,N_4073);
or UO_14 (O_14,N_4543,N_4866);
or UO_15 (O_15,N_4882,N_4536);
or UO_16 (O_16,N_4486,N_4042);
or UO_17 (O_17,N_4115,N_4177);
nand UO_18 (O_18,N_4191,N_4916);
nand UO_19 (O_19,N_4730,N_4128);
or UO_20 (O_20,N_4379,N_4274);
nand UO_21 (O_21,N_4290,N_4606);
nand UO_22 (O_22,N_4817,N_4974);
or UO_23 (O_23,N_4696,N_4245);
and UO_24 (O_24,N_4045,N_4848);
or UO_25 (O_25,N_4305,N_4049);
nor UO_26 (O_26,N_4399,N_4041);
and UO_27 (O_27,N_4375,N_4756);
or UO_28 (O_28,N_4677,N_4385);
or UO_29 (O_29,N_4578,N_4503);
and UO_30 (O_30,N_4064,N_4237);
xor UO_31 (O_31,N_4388,N_4990);
nand UO_32 (O_32,N_4509,N_4872);
nor UO_33 (O_33,N_4597,N_4845);
nor UO_34 (O_34,N_4370,N_4180);
and UO_35 (O_35,N_4322,N_4704);
and UO_36 (O_36,N_4475,N_4133);
nor UO_37 (O_37,N_4153,N_4921);
or UO_38 (O_38,N_4646,N_4474);
nor UO_39 (O_39,N_4230,N_4363);
or UO_40 (O_40,N_4482,N_4136);
or UO_41 (O_41,N_4028,N_4037);
or UO_42 (O_42,N_4855,N_4637);
and UO_43 (O_43,N_4173,N_4770);
xnor UO_44 (O_44,N_4613,N_4241);
or UO_45 (O_45,N_4601,N_4579);
nand UO_46 (O_46,N_4896,N_4825);
and UO_47 (O_47,N_4863,N_4391);
or UO_48 (O_48,N_4956,N_4465);
and UO_49 (O_49,N_4072,N_4157);
or UO_50 (O_50,N_4694,N_4428);
and UO_51 (O_51,N_4183,N_4731);
nor UO_52 (O_52,N_4095,N_4006);
nor UO_53 (O_53,N_4398,N_4676);
nand UO_54 (O_54,N_4627,N_4955);
or UO_55 (O_55,N_4668,N_4821);
or UO_56 (O_56,N_4270,N_4277);
and UO_57 (O_57,N_4186,N_4221);
nor UO_58 (O_58,N_4726,N_4492);
nor UO_59 (O_59,N_4479,N_4044);
nor UO_60 (O_60,N_4522,N_4788);
nor UO_61 (O_61,N_4351,N_4602);
or UO_62 (O_62,N_4093,N_4423);
and UO_63 (O_63,N_4435,N_4117);
nor UO_64 (O_64,N_4617,N_4745);
nor UO_65 (O_65,N_4887,N_4387);
nand UO_66 (O_66,N_4378,N_4170);
and UO_67 (O_67,N_4961,N_4958);
nand UO_68 (O_68,N_4406,N_4689);
or UO_69 (O_69,N_4569,N_4764);
and UO_70 (O_70,N_4877,N_4316);
nor UO_71 (O_71,N_4498,N_4437);
nor UO_72 (O_72,N_4315,N_4488);
and UO_73 (O_73,N_4997,N_4101);
nor UO_74 (O_74,N_4758,N_4598);
nand UO_75 (O_75,N_4496,N_4381);
or UO_76 (O_76,N_4714,N_4767);
and UO_77 (O_77,N_4557,N_4131);
nor UO_78 (O_78,N_4619,N_4596);
nand UO_79 (O_79,N_4140,N_4586);
nand UO_80 (O_80,N_4297,N_4213);
nor UO_81 (O_81,N_4506,N_4001);
nor UO_82 (O_82,N_4996,N_4122);
nor UO_83 (O_83,N_4841,N_4218);
nand UO_84 (O_84,N_4220,N_4829);
or UO_85 (O_85,N_4727,N_4471);
nand UO_86 (O_86,N_4830,N_4338);
nand UO_87 (O_87,N_4105,N_4765);
nor UO_88 (O_88,N_4738,N_4296);
nor UO_89 (O_89,N_4806,N_4559);
and UO_90 (O_90,N_4026,N_4312);
and UO_91 (O_91,N_4693,N_4250);
nand UO_92 (O_92,N_4584,N_4831);
nor UO_93 (O_93,N_4654,N_4636);
nand UO_94 (O_94,N_4743,N_4047);
nand UO_95 (O_95,N_4755,N_4761);
or UO_96 (O_96,N_4440,N_4130);
or UO_97 (O_97,N_4525,N_4941);
nor UO_98 (O_98,N_4068,N_4906);
nand UO_99 (O_99,N_4334,N_4741);
nor UO_100 (O_100,N_4361,N_4035);
or UO_101 (O_101,N_4080,N_4329);
nor UO_102 (O_102,N_4902,N_4840);
nor UO_103 (O_103,N_4141,N_4138);
or UO_104 (O_104,N_4104,N_4123);
nor UO_105 (O_105,N_4989,N_4909);
or UO_106 (O_106,N_4228,N_4345);
nor UO_107 (O_107,N_4642,N_4701);
or UO_108 (O_108,N_4348,N_4832);
and UO_109 (O_109,N_4552,N_4930);
nand UO_110 (O_110,N_4110,N_4069);
or UO_111 (O_111,N_4566,N_4703);
nand UO_112 (O_112,N_4928,N_4350);
or UO_113 (O_113,N_4332,N_4807);
nor UO_114 (O_114,N_4339,N_4317);
nor UO_115 (O_115,N_4175,N_4667);
nor UO_116 (O_116,N_4669,N_4447);
nor UO_117 (O_117,N_4960,N_4702);
or UO_118 (O_118,N_4898,N_4808);
and UO_119 (O_119,N_4534,N_4926);
nand UO_120 (O_120,N_4327,N_4034);
and UO_121 (O_121,N_4193,N_4612);
nor UO_122 (O_122,N_4202,N_4744);
nor UO_123 (O_123,N_4635,N_4463);
or UO_124 (O_124,N_4735,N_4698);
nor UO_125 (O_125,N_4976,N_4024);
nand UO_126 (O_126,N_4528,N_4574);
nor UO_127 (O_127,N_4897,N_4413);
and UO_128 (O_128,N_4889,N_4448);
nand UO_129 (O_129,N_4000,N_4092);
and UO_130 (O_130,N_4979,N_4288);
and UO_131 (O_131,N_4320,N_4734);
nor UO_132 (O_132,N_4993,N_4847);
and UO_133 (O_133,N_4480,N_4798);
nor UO_134 (O_134,N_4065,N_4539);
or UO_135 (O_135,N_4537,N_4533);
nor UO_136 (O_136,N_4039,N_4615);
nand UO_137 (O_137,N_4394,N_4003);
nand UO_138 (O_138,N_4940,N_4565);
nor UO_139 (O_139,N_4155,N_4850);
or UO_140 (O_140,N_4580,N_4127);
nand UO_141 (O_141,N_4323,N_4925);
and UO_142 (O_142,N_4776,N_4742);
or UO_143 (O_143,N_4512,N_4477);
nand UO_144 (O_144,N_4951,N_4374);
nand UO_145 (O_145,N_4022,N_4868);
nand UO_146 (O_146,N_4713,N_4293);
and UO_147 (O_147,N_4038,N_4760);
nor UO_148 (O_148,N_4723,N_4680);
or UO_149 (O_149,N_4908,N_4978);
nor UO_150 (O_150,N_4014,N_4152);
nand UO_151 (O_151,N_4091,N_4287);
xor UO_152 (O_152,N_4836,N_4025);
nor UO_153 (O_153,N_4162,N_4271);
nor UO_154 (O_154,N_4950,N_4160);
nand UO_155 (O_155,N_4273,N_4239);
nand UO_156 (O_156,N_4674,N_4185);
nand UO_157 (O_157,N_4266,N_4054);
or UO_158 (O_158,N_4188,N_4985);
and UO_159 (O_159,N_4149,N_4395);
and UO_160 (O_160,N_4733,N_4556);
or UO_161 (O_161,N_4470,N_4343);
or UO_162 (O_162,N_4912,N_4298);
nand UO_163 (O_163,N_4880,N_4113);
and UO_164 (O_164,N_4629,N_4207);
nand UO_165 (O_165,N_4823,N_4881);
and UO_166 (O_166,N_4156,N_4461);
or UO_167 (O_167,N_4519,N_4969);
and UO_168 (O_168,N_4386,N_4009);
nor UO_169 (O_169,N_4750,N_4875);
nor UO_170 (O_170,N_4728,N_4894);
nor UO_171 (O_171,N_4737,N_4822);
and UO_172 (O_172,N_4259,N_4573);
or UO_173 (O_173,N_4425,N_4178);
nor UO_174 (O_174,N_4966,N_4661);
and UO_175 (O_175,N_4545,N_4446);
nand UO_176 (O_176,N_4604,N_4513);
and UO_177 (O_177,N_4711,N_4777);
or UO_178 (O_178,N_4222,N_4546);
xor UO_179 (O_179,N_4782,N_4827);
nor UO_180 (O_180,N_4356,N_4411);
or UO_181 (O_181,N_4527,N_4524);
nand UO_182 (O_182,N_4722,N_4946);
and UO_183 (O_183,N_4520,N_4942);
or UO_184 (O_184,N_4874,N_4626);
nand UO_185 (O_185,N_4518,N_4769);
or UO_186 (O_186,N_4772,N_4063);
nor UO_187 (O_187,N_4614,N_4048);
nand UO_188 (O_188,N_4995,N_4529);
nor UO_189 (O_189,N_4640,N_4724);
nand UO_190 (O_190,N_4895,N_4489);
nor UO_191 (O_191,N_4998,N_4919);
nor UO_192 (O_192,N_4986,N_4860);
nor UO_193 (O_193,N_4576,N_4957);
and UO_194 (O_194,N_4622,N_4663);
and UO_195 (O_195,N_4004,N_4258);
and UO_196 (O_196,N_4885,N_4762);
or UO_197 (O_197,N_4008,N_4797);
or UO_198 (O_198,N_4060,N_4516);
nor UO_199 (O_199,N_4856,N_4295);
or UO_200 (O_200,N_4264,N_4352);
and UO_201 (O_201,N_4630,N_4013);
nor UO_202 (O_202,N_4493,N_4124);
nand UO_203 (O_203,N_4785,N_4359);
nor UO_204 (O_204,N_4341,N_4706);
nor UO_205 (O_205,N_4795,N_4526);
and UO_206 (O_206,N_4076,N_4262);
nor UO_207 (O_207,N_4655,N_4445);
or UO_208 (O_208,N_4253,N_4236);
and UO_209 (O_209,N_4900,N_4301);
nor UO_210 (O_210,N_4815,N_4040);
nor UO_211 (O_211,N_4784,N_4901);
and UO_212 (O_212,N_4252,N_4050);
nor UO_213 (O_213,N_4310,N_4599);
and UO_214 (O_214,N_4963,N_4420);
nand UO_215 (O_215,N_4975,N_4019);
nor UO_216 (O_216,N_4820,N_4082);
nor UO_217 (O_217,N_4248,N_4907);
nor UO_218 (O_218,N_4535,N_4981);
nor UO_219 (O_219,N_4583,N_4431);
and UO_220 (O_220,N_4144,N_4905);
nand UO_221 (O_221,N_4494,N_4947);
and UO_222 (O_222,N_4948,N_4936);
nor UO_223 (O_223,N_4109,N_4538);
nor UO_224 (O_224,N_4016,N_4125);
and UO_225 (O_225,N_4208,N_4548);
or UO_226 (O_226,N_4390,N_4229);
and UO_227 (O_227,N_4865,N_4718);
and UO_228 (O_228,N_4754,N_4134);
or UO_229 (O_229,N_4427,N_4937);
nor UO_230 (O_230,N_4588,N_4892);
and UO_231 (O_231,N_4719,N_4384);
nand UO_232 (O_232,N_4837,N_4910);
nor UO_233 (O_233,N_4555,N_4189);
and UO_234 (O_234,N_4861,N_4059);
and UO_235 (O_235,N_4439,N_4652);
xnor UO_236 (O_236,N_4883,N_4721);
nor UO_237 (O_237,N_4396,N_4198);
and UO_238 (O_238,N_4729,N_4233);
nand UO_239 (O_239,N_4254,N_4313);
or UO_240 (O_240,N_4732,N_4326);
nor UO_241 (O_241,N_4292,N_4544);
or UO_242 (O_242,N_4826,N_4839);
nand UO_243 (O_243,N_4540,N_4051);
and UO_244 (O_244,N_4999,N_4833);
or UO_245 (O_245,N_4504,N_4393);
or UO_246 (O_246,N_4416,N_4859);
nor UO_247 (O_247,N_4417,N_4547);
nor UO_248 (O_248,N_4665,N_4247);
nor UO_249 (O_249,N_4405,N_4438);
nand UO_250 (O_250,N_4285,N_4862);
nand UO_251 (O_251,N_4083,N_4176);
nor UO_252 (O_252,N_4549,N_4725);
and UO_253 (O_253,N_4814,N_4336);
nand UO_254 (O_254,N_4377,N_4349);
and UO_255 (O_255,N_4112,N_4424);
or UO_256 (O_256,N_4304,N_4542);
nand UO_257 (O_257,N_4623,N_4816);
and UO_258 (O_258,N_4720,N_4712);
nand UO_259 (O_259,N_4018,N_4952);
nor UO_260 (O_260,N_4575,N_4046);
or UO_261 (O_261,N_4799,N_4021);
or UO_262 (O_262,N_4342,N_4012);
or UO_263 (O_263,N_4276,N_4154);
nor UO_264 (O_264,N_4397,N_4914);
and UO_265 (O_265,N_4194,N_4801);
or UO_266 (O_266,N_4585,N_4904);
and UO_267 (O_267,N_4867,N_4790);
nor UO_268 (O_268,N_4410,N_4358);
or UO_269 (O_269,N_4505,N_4369);
nand UO_270 (O_270,N_4740,N_4158);
nor UO_271 (O_271,N_4682,N_4182);
or UO_272 (O_272,N_4196,N_4644);
or UO_273 (O_273,N_4871,N_4043);
nor UO_274 (O_274,N_4145,N_4927);
nor UO_275 (O_275,N_4500,N_4197);
nor UO_276 (O_276,N_4577,N_4774);
nand UO_277 (O_277,N_4949,N_4007);
nand UO_278 (O_278,N_4366,N_4562);
nor UO_279 (O_279,N_4311,N_4272);
or UO_280 (O_280,N_4834,N_4563);
or UO_281 (O_281,N_4768,N_4675);
and UO_282 (O_282,N_4100,N_4521);
or UO_283 (O_283,N_4070,N_4415);
and UO_284 (O_284,N_4650,N_4357);
or UO_285 (O_285,N_4699,N_4673);
nand UO_286 (O_286,N_4691,N_4511);
nor UO_287 (O_287,N_4325,N_4407);
nor UO_288 (O_288,N_4466,N_4473);
nor UO_289 (O_289,N_4242,N_4656);
nor UO_290 (O_290,N_4199,N_4085);
and UO_291 (O_291,N_4980,N_4057);
and UO_292 (O_292,N_4685,N_4710);
nor UO_293 (O_293,N_4094,N_4027);
nor UO_294 (O_294,N_4987,N_4697);
nor UO_295 (O_295,N_4568,N_4373);
or UO_296 (O_296,N_4204,N_4893);
nor UO_297 (O_297,N_4879,N_4809);
nor UO_298 (O_298,N_4086,N_4195);
nor UO_299 (O_299,N_4432,N_4169);
nor UO_300 (O_300,N_4052,N_4321);
nor UO_301 (O_301,N_4853,N_4608);
nand UO_302 (O_302,N_4087,N_4079);
and UO_303 (O_303,N_4736,N_4462);
nor UO_304 (O_304,N_4380,N_4911);
or UO_305 (O_305,N_4347,N_4216);
nor UO_306 (O_306,N_4005,N_4056);
nor UO_307 (O_307,N_4015,N_4616);
and UO_308 (O_308,N_4263,N_4365);
nand UO_309 (O_309,N_4625,N_4499);
or UO_310 (O_310,N_4227,N_4419);
nor UO_311 (O_311,N_4593,N_4564);
or UO_312 (O_312,N_4257,N_4286);
nand UO_313 (O_313,N_4142,N_4077);
and UO_314 (O_314,N_4683,N_4283);
or UO_315 (O_315,N_4238,N_4752);
nand UO_316 (O_316,N_4137,N_4472);
or UO_317 (O_317,N_4164,N_4794);
nor UO_318 (O_318,N_4226,N_4033);
nor UO_319 (O_319,N_4485,N_4074);
and UO_320 (O_320,N_4468,N_4402);
nand UO_321 (O_321,N_4017,N_4294);
nor UO_322 (O_322,N_4231,N_4994);
nand UO_323 (O_323,N_4959,N_4097);
nand UO_324 (O_324,N_4139,N_4591);
nand UO_325 (O_325,N_4071,N_4934);
and UO_326 (O_326,N_4571,N_4337);
or UO_327 (O_327,N_4308,N_4943);
and UO_328 (O_328,N_4553,N_4789);
nor UO_329 (O_329,N_4531,N_4884);
nand UO_330 (O_330,N_4168,N_4464);
or UO_331 (O_331,N_4458,N_4058);
nor UO_332 (O_332,N_4851,N_4203);
or UO_333 (O_333,N_4444,N_4802);
or UO_334 (O_334,N_4922,N_4633);
or UO_335 (O_335,N_4643,N_4344);
or UO_336 (O_336,N_4456,N_4849);
nand UO_337 (O_337,N_4838,N_4240);
and UO_338 (O_338,N_4314,N_4031);
or UO_339 (O_339,N_4036,N_4457);
nor UO_340 (O_340,N_4067,N_4029);
nor UO_341 (O_341,N_4747,N_4913);
nand UO_342 (O_342,N_4687,N_4753);
and UO_343 (O_343,N_4924,N_4382);
nor UO_344 (O_344,N_4269,N_4163);
nor UO_345 (O_345,N_4476,N_4988);
and UO_346 (O_346,N_4484,N_4002);
nand UO_347 (O_347,N_4915,N_4291);
or UO_348 (O_348,N_4490,N_4442);
or UO_349 (O_349,N_4641,N_4962);
or UO_350 (O_350,N_4108,N_4106);
and UO_351 (O_351,N_4099,N_4430);
nand UO_352 (O_352,N_4690,N_4030);
nor UO_353 (O_353,N_4890,N_4215);
nand UO_354 (O_354,N_4695,N_4717);
or UO_355 (O_355,N_4748,N_4126);
nand UO_356 (O_356,N_4810,N_4681);
or UO_357 (O_357,N_4692,N_4205);
and UO_358 (O_358,N_4212,N_4551);
and UO_359 (O_359,N_4716,N_4224);
or UO_360 (O_360,N_4066,N_4828);
and UO_361 (O_361,N_4467,N_4903);
and UO_362 (O_362,N_4159,N_4103);
nor UO_363 (O_363,N_4403,N_4032);
or UO_364 (O_364,N_4098,N_4605);
and UO_365 (O_365,N_4869,N_4408);
nand UO_366 (O_366,N_4118,N_4354);
and UO_367 (O_367,N_4931,N_4282);
and UO_368 (O_368,N_4920,N_4116);
or UO_369 (O_369,N_4972,N_4739);
and UO_370 (O_370,N_4624,N_4491);
nand UO_371 (O_371,N_4443,N_4102);
nand UO_372 (O_372,N_4372,N_4923);
and UO_373 (O_373,N_4166,N_4409);
or UO_374 (O_374,N_4333,N_4560);
and UO_375 (O_375,N_4842,N_4715);
nand UO_376 (O_376,N_4507,N_4595);
nand UO_377 (O_377,N_4554,N_4918);
nor UO_378 (O_378,N_4232,N_4700);
and UO_379 (O_379,N_4346,N_4984);
nor UO_380 (O_380,N_4561,N_4275);
nand UO_381 (O_381,N_4813,N_4279);
or UO_382 (O_382,N_4090,N_4223);
nor UO_383 (O_383,N_4705,N_4620);
and UO_384 (O_384,N_4660,N_4284);
nor UO_385 (O_385,N_4055,N_4020);
nand UO_386 (O_386,N_4751,N_4818);
xnor UO_387 (O_387,N_4787,N_4400);
nor UO_388 (O_388,N_4151,N_4418);
and UO_389 (O_389,N_4256,N_4331);
or UO_390 (O_390,N_4330,N_4453);
nand UO_391 (O_391,N_4119,N_4982);
and UO_392 (O_392,N_4651,N_4481);
or UO_393 (O_393,N_4010,N_4146);
and UO_394 (O_394,N_4299,N_4084);
nor UO_395 (O_395,N_4964,N_4502);
or UO_396 (O_396,N_4353,N_4174);
nand UO_397 (O_397,N_4632,N_4234);
nor UO_398 (O_398,N_4383,N_4433);
or UO_399 (O_399,N_4746,N_4983);
or UO_400 (O_400,N_4791,N_4243);
and UO_401 (O_401,N_4260,N_4819);
nor UO_402 (O_402,N_4147,N_4664);
or UO_403 (O_403,N_4558,N_4469);
nand UO_404 (O_404,N_4088,N_4679);
nand UO_405 (O_405,N_4878,N_4844);
nor UO_406 (O_406,N_4804,N_4550);
xnor UO_407 (O_407,N_4932,N_4300);
or UO_408 (O_408,N_4970,N_4251);
nor UO_409 (O_409,N_4678,N_4587);
nor UO_410 (O_410,N_4306,N_4638);
and UO_411 (O_411,N_4672,N_4945);
nor UO_412 (O_412,N_4935,N_4780);
and UO_413 (O_413,N_4572,N_4089);
nand UO_414 (O_414,N_4401,N_4590);
nor UO_415 (O_415,N_4302,N_4449);
nand UO_416 (O_416,N_4603,N_4968);
and UO_417 (O_417,N_4864,N_4666);
nand UO_418 (O_418,N_4450,N_4023);
nor UO_419 (O_419,N_4708,N_4645);
nor UO_420 (O_420,N_4581,N_4766);
or UO_421 (O_421,N_4478,N_4870);
and UO_422 (O_422,N_4340,N_4206);
nor UO_423 (O_423,N_4621,N_4487);
or UO_424 (O_424,N_4371,N_4184);
or UO_425 (O_425,N_4495,N_4135);
or UO_426 (O_426,N_4335,N_4973);
nand UO_427 (O_427,N_4451,N_4179);
and UO_428 (O_428,N_4589,N_4364);
or UO_429 (O_429,N_4779,N_4309);
and UO_430 (O_430,N_4360,N_4671);
or UO_431 (O_431,N_4759,N_4143);
and UO_432 (O_432,N_4929,N_4129);
nor UO_433 (O_433,N_4429,N_4201);
nand UO_434 (O_434,N_4053,N_4355);
or UO_435 (O_435,N_4265,N_4508);
nand UO_436 (O_436,N_4107,N_4062);
nand UO_437 (O_437,N_4209,N_4497);
nand UO_438 (O_438,N_4873,N_4459);
nand UO_439 (O_439,N_4172,N_4541);
nand UO_440 (O_440,N_4114,N_4307);
nand UO_441 (O_441,N_4594,N_4786);
or UO_442 (O_442,N_4857,N_4523);
or UO_443 (O_443,N_4888,N_4953);
or UO_444 (O_444,N_4778,N_4235);
nor UO_445 (O_445,N_4422,N_4392);
or UO_446 (O_446,N_4653,N_4362);
and UO_447 (O_447,N_4281,N_4318);
xor UO_448 (O_448,N_4210,N_4171);
or UO_449 (O_449,N_4707,N_4891);
nand UO_450 (O_450,N_4917,N_4120);
nor UO_451 (O_451,N_4639,N_4967);
nor UO_452 (O_452,N_4530,N_4570);
nand UO_453 (O_453,N_4781,N_4775);
or UO_454 (O_454,N_4670,N_4111);
nand UO_455 (O_455,N_4824,N_4662);
and UO_456 (O_456,N_4647,N_4532);
nor UO_457 (O_457,N_4658,N_4944);
and UO_458 (O_458,N_4289,N_4749);
nor UO_459 (O_459,N_4992,N_4609);
and UO_460 (O_460,N_4835,N_4244);
or UO_461 (O_461,N_4688,N_4061);
or UO_462 (O_462,N_4187,N_4167);
nor UO_463 (O_463,N_4763,N_4611);
and UO_464 (O_464,N_4886,N_4255);
nor UO_465 (O_465,N_4965,N_4514);
or UO_466 (O_466,N_4634,N_4757);
nor UO_467 (O_467,N_4214,N_4078);
nand UO_468 (O_468,N_4607,N_4225);
nor UO_469 (O_469,N_4441,N_4939);
nor UO_470 (O_470,N_4812,N_4426);
or UO_471 (O_471,N_4628,N_4267);
nor UO_472 (O_472,N_4319,N_4280);
nand UO_473 (O_473,N_4434,N_4686);
and UO_474 (O_474,N_4150,N_4783);
and UO_475 (O_475,N_4211,N_4161);
nand UO_476 (O_476,N_4421,N_4165);
and UO_477 (O_477,N_4938,N_4181);
and UO_478 (O_478,N_4991,N_4971);
nand UO_479 (O_479,N_4412,N_4771);
and UO_480 (O_480,N_4954,N_4268);
and UO_481 (O_481,N_4121,N_4510);
nand UO_482 (O_482,N_4324,N_4796);
and UO_483 (O_483,N_4303,N_4899);
or UO_484 (O_484,N_4075,N_4858);
and UO_485 (O_485,N_4582,N_4567);
or UO_486 (O_486,N_4792,N_4803);
nor UO_487 (O_487,N_4414,N_4876);
nand UO_488 (O_488,N_4483,N_4618);
or UO_489 (O_489,N_4192,N_4657);
and UO_490 (O_490,N_4610,N_4367);
nor UO_491 (O_491,N_4190,N_4011);
and UO_492 (O_492,N_4843,N_4454);
and UO_493 (O_493,N_4977,N_4811);
and UO_494 (O_494,N_4249,N_4649);
or UO_495 (O_495,N_4631,N_4219);
nor UO_496 (O_496,N_4328,N_4278);
and UO_497 (O_497,N_4684,N_4846);
and UO_498 (O_498,N_4096,N_4515);
nand UO_499 (O_499,N_4773,N_4805);
and UO_500 (O_500,N_4366,N_4370);
and UO_501 (O_501,N_4948,N_4772);
nor UO_502 (O_502,N_4272,N_4337);
xor UO_503 (O_503,N_4221,N_4456);
and UO_504 (O_504,N_4679,N_4650);
nand UO_505 (O_505,N_4222,N_4411);
and UO_506 (O_506,N_4868,N_4810);
and UO_507 (O_507,N_4893,N_4297);
nor UO_508 (O_508,N_4016,N_4940);
and UO_509 (O_509,N_4710,N_4603);
nand UO_510 (O_510,N_4587,N_4299);
or UO_511 (O_511,N_4440,N_4166);
nor UO_512 (O_512,N_4405,N_4073);
nor UO_513 (O_513,N_4037,N_4315);
nor UO_514 (O_514,N_4130,N_4874);
or UO_515 (O_515,N_4834,N_4152);
and UO_516 (O_516,N_4098,N_4182);
or UO_517 (O_517,N_4294,N_4920);
or UO_518 (O_518,N_4374,N_4014);
nor UO_519 (O_519,N_4270,N_4969);
nor UO_520 (O_520,N_4219,N_4679);
nor UO_521 (O_521,N_4013,N_4640);
nand UO_522 (O_522,N_4371,N_4187);
or UO_523 (O_523,N_4789,N_4921);
or UO_524 (O_524,N_4457,N_4833);
and UO_525 (O_525,N_4419,N_4484);
and UO_526 (O_526,N_4722,N_4826);
nor UO_527 (O_527,N_4393,N_4470);
nor UO_528 (O_528,N_4152,N_4432);
and UO_529 (O_529,N_4222,N_4049);
nand UO_530 (O_530,N_4256,N_4647);
and UO_531 (O_531,N_4263,N_4787);
or UO_532 (O_532,N_4284,N_4176);
and UO_533 (O_533,N_4738,N_4967);
xnor UO_534 (O_534,N_4852,N_4133);
nand UO_535 (O_535,N_4357,N_4870);
nand UO_536 (O_536,N_4238,N_4298);
nand UO_537 (O_537,N_4429,N_4175);
nand UO_538 (O_538,N_4730,N_4081);
and UO_539 (O_539,N_4972,N_4497);
nor UO_540 (O_540,N_4560,N_4104);
nand UO_541 (O_541,N_4695,N_4197);
and UO_542 (O_542,N_4379,N_4739);
and UO_543 (O_543,N_4989,N_4709);
nor UO_544 (O_544,N_4981,N_4709);
and UO_545 (O_545,N_4520,N_4296);
nor UO_546 (O_546,N_4327,N_4416);
nor UO_547 (O_547,N_4603,N_4530);
nor UO_548 (O_548,N_4747,N_4687);
nand UO_549 (O_549,N_4983,N_4039);
nand UO_550 (O_550,N_4181,N_4654);
nand UO_551 (O_551,N_4522,N_4100);
xor UO_552 (O_552,N_4362,N_4880);
and UO_553 (O_553,N_4440,N_4694);
nor UO_554 (O_554,N_4469,N_4220);
or UO_555 (O_555,N_4669,N_4293);
nand UO_556 (O_556,N_4188,N_4268);
nor UO_557 (O_557,N_4569,N_4972);
nand UO_558 (O_558,N_4523,N_4278);
nor UO_559 (O_559,N_4578,N_4152);
or UO_560 (O_560,N_4719,N_4382);
or UO_561 (O_561,N_4772,N_4964);
nor UO_562 (O_562,N_4963,N_4523);
and UO_563 (O_563,N_4019,N_4668);
or UO_564 (O_564,N_4642,N_4630);
nor UO_565 (O_565,N_4243,N_4174);
or UO_566 (O_566,N_4967,N_4249);
or UO_567 (O_567,N_4850,N_4840);
and UO_568 (O_568,N_4767,N_4543);
and UO_569 (O_569,N_4588,N_4372);
nand UO_570 (O_570,N_4853,N_4393);
nand UO_571 (O_571,N_4969,N_4393);
nor UO_572 (O_572,N_4248,N_4265);
and UO_573 (O_573,N_4089,N_4518);
and UO_574 (O_574,N_4392,N_4887);
nor UO_575 (O_575,N_4102,N_4158);
nand UO_576 (O_576,N_4469,N_4958);
and UO_577 (O_577,N_4684,N_4440);
nand UO_578 (O_578,N_4316,N_4842);
nand UO_579 (O_579,N_4518,N_4417);
and UO_580 (O_580,N_4877,N_4359);
nand UO_581 (O_581,N_4807,N_4314);
nand UO_582 (O_582,N_4963,N_4947);
nor UO_583 (O_583,N_4006,N_4853);
nor UO_584 (O_584,N_4491,N_4681);
nand UO_585 (O_585,N_4951,N_4237);
or UO_586 (O_586,N_4397,N_4926);
xnor UO_587 (O_587,N_4025,N_4296);
or UO_588 (O_588,N_4533,N_4189);
or UO_589 (O_589,N_4652,N_4581);
or UO_590 (O_590,N_4969,N_4353);
nand UO_591 (O_591,N_4803,N_4589);
and UO_592 (O_592,N_4610,N_4189);
nand UO_593 (O_593,N_4554,N_4960);
or UO_594 (O_594,N_4492,N_4175);
nor UO_595 (O_595,N_4022,N_4390);
nor UO_596 (O_596,N_4646,N_4795);
nand UO_597 (O_597,N_4701,N_4493);
nor UO_598 (O_598,N_4548,N_4283);
or UO_599 (O_599,N_4413,N_4701);
nand UO_600 (O_600,N_4937,N_4737);
nand UO_601 (O_601,N_4907,N_4241);
nand UO_602 (O_602,N_4352,N_4635);
nand UO_603 (O_603,N_4721,N_4148);
and UO_604 (O_604,N_4546,N_4081);
nand UO_605 (O_605,N_4919,N_4104);
and UO_606 (O_606,N_4891,N_4009);
nor UO_607 (O_607,N_4407,N_4656);
or UO_608 (O_608,N_4959,N_4645);
nand UO_609 (O_609,N_4667,N_4980);
and UO_610 (O_610,N_4456,N_4426);
nor UO_611 (O_611,N_4396,N_4924);
nand UO_612 (O_612,N_4981,N_4168);
or UO_613 (O_613,N_4622,N_4801);
and UO_614 (O_614,N_4630,N_4609);
or UO_615 (O_615,N_4824,N_4438);
nand UO_616 (O_616,N_4843,N_4631);
or UO_617 (O_617,N_4626,N_4622);
and UO_618 (O_618,N_4260,N_4962);
nor UO_619 (O_619,N_4030,N_4069);
nand UO_620 (O_620,N_4012,N_4716);
or UO_621 (O_621,N_4720,N_4913);
and UO_622 (O_622,N_4589,N_4604);
and UO_623 (O_623,N_4866,N_4101);
and UO_624 (O_624,N_4495,N_4219);
nor UO_625 (O_625,N_4651,N_4678);
nor UO_626 (O_626,N_4396,N_4863);
and UO_627 (O_627,N_4627,N_4914);
nand UO_628 (O_628,N_4861,N_4956);
nor UO_629 (O_629,N_4104,N_4882);
nand UO_630 (O_630,N_4296,N_4956);
and UO_631 (O_631,N_4954,N_4738);
nand UO_632 (O_632,N_4970,N_4225);
and UO_633 (O_633,N_4021,N_4624);
nand UO_634 (O_634,N_4431,N_4309);
and UO_635 (O_635,N_4401,N_4715);
and UO_636 (O_636,N_4972,N_4131);
or UO_637 (O_637,N_4895,N_4811);
or UO_638 (O_638,N_4009,N_4494);
or UO_639 (O_639,N_4522,N_4636);
nor UO_640 (O_640,N_4715,N_4661);
nand UO_641 (O_641,N_4875,N_4394);
nand UO_642 (O_642,N_4246,N_4625);
nor UO_643 (O_643,N_4284,N_4557);
and UO_644 (O_644,N_4942,N_4873);
or UO_645 (O_645,N_4120,N_4558);
nor UO_646 (O_646,N_4328,N_4072);
nand UO_647 (O_647,N_4766,N_4105);
nand UO_648 (O_648,N_4673,N_4876);
or UO_649 (O_649,N_4641,N_4557);
nor UO_650 (O_650,N_4176,N_4766);
or UO_651 (O_651,N_4334,N_4481);
nor UO_652 (O_652,N_4647,N_4346);
or UO_653 (O_653,N_4928,N_4803);
nor UO_654 (O_654,N_4406,N_4075);
and UO_655 (O_655,N_4361,N_4116);
or UO_656 (O_656,N_4721,N_4746);
nand UO_657 (O_657,N_4826,N_4619);
xnor UO_658 (O_658,N_4246,N_4303);
nor UO_659 (O_659,N_4102,N_4469);
or UO_660 (O_660,N_4158,N_4765);
nor UO_661 (O_661,N_4091,N_4045);
nand UO_662 (O_662,N_4559,N_4453);
and UO_663 (O_663,N_4689,N_4831);
nand UO_664 (O_664,N_4815,N_4758);
nor UO_665 (O_665,N_4955,N_4185);
and UO_666 (O_666,N_4792,N_4479);
nand UO_667 (O_667,N_4051,N_4765);
nor UO_668 (O_668,N_4812,N_4680);
nor UO_669 (O_669,N_4084,N_4025);
nor UO_670 (O_670,N_4280,N_4660);
nor UO_671 (O_671,N_4107,N_4244);
nor UO_672 (O_672,N_4731,N_4048);
and UO_673 (O_673,N_4713,N_4894);
or UO_674 (O_674,N_4162,N_4832);
nand UO_675 (O_675,N_4135,N_4624);
or UO_676 (O_676,N_4389,N_4339);
and UO_677 (O_677,N_4454,N_4466);
or UO_678 (O_678,N_4529,N_4169);
or UO_679 (O_679,N_4445,N_4908);
or UO_680 (O_680,N_4342,N_4536);
nor UO_681 (O_681,N_4807,N_4365);
or UO_682 (O_682,N_4051,N_4545);
nor UO_683 (O_683,N_4788,N_4109);
nand UO_684 (O_684,N_4095,N_4614);
and UO_685 (O_685,N_4311,N_4086);
and UO_686 (O_686,N_4530,N_4435);
or UO_687 (O_687,N_4908,N_4381);
nand UO_688 (O_688,N_4664,N_4231);
or UO_689 (O_689,N_4737,N_4575);
nand UO_690 (O_690,N_4051,N_4005);
nand UO_691 (O_691,N_4338,N_4066);
nand UO_692 (O_692,N_4888,N_4177);
nor UO_693 (O_693,N_4883,N_4485);
or UO_694 (O_694,N_4829,N_4760);
and UO_695 (O_695,N_4221,N_4539);
nor UO_696 (O_696,N_4697,N_4465);
nor UO_697 (O_697,N_4347,N_4967);
nand UO_698 (O_698,N_4445,N_4589);
and UO_699 (O_699,N_4209,N_4772);
and UO_700 (O_700,N_4620,N_4836);
nand UO_701 (O_701,N_4404,N_4581);
and UO_702 (O_702,N_4499,N_4378);
and UO_703 (O_703,N_4631,N_4076);
nor UO_704 (O_704,N_4817,N_4197);
and UO_705 (O_705,N_4979,N_4128);
nand UO_706 (O_706,N_4785,N_4854);
nand UO_707 (O_707,N_4249,N_4346);
nor UO_708 (O_708,N_4274,N_4257);
or UO_709 (O_709,N_4191,N_4460);
nor UO_710 (O_710,N_4275,N_4447);
or UO_711 (O_711,N_4681,N_4394);
or UO_712 (O_712,N_4485,N_4552);
or UO_713 (O_713,N_4818,N_4236);
or UO_714 (O_714,N_4366,N_4358);
or UO_715 (O_715,N_4463,N_4117);
nor UO_716 (O_716,N_4667,N_4784);
nor UO_717 (O_717,N_4745,N_4631);
and UO_718 (O_718,N_4941,N_4208);
and UO_719 (O_719,N_4813,N_4480);
nor UO_720 (O_720,N_4680,N_4796);
or UO_721 (O_721,N_4737,N_4302);
and UO_722 (O_722,N_4818,N_4349);
nor UO_723 (O_723,N_4061,N_4472);
nor UO_724 (O_724,N_4825,N_4935);
and UO_725 (O_725,N_4110,N_4868);
nor UO_726 (O_726,N_4589,N_4610);
xor UO_727 (O_727,N_4806,N_4482);
and UO_728 (O_728,N_4524,N_4143);
nor UO_729 (O_729,N_4571,N_4504);
nand UO_730 (O_730,N_4577,N_4153);
nand UO_731 (O_731,N_4725,N_4519);
or UO_732 (O_732,N_4013,N_4005);
nor UO_733 (O_733,N_4117,N_4004);
nand UO_734 (O_734,N_4335,N_4129);
nand UO_735 (O_735,N_4348,N_4569);
or UO_736 (O_736,N_4029,N_4049);
nor UO_737 (O_737,N_4255,N_4833);
or UO_738 (O_738,N_4526,N_4472);
or UO_739 (O_739,N_4728,N_4845);
or UO_740 (O_740,N_4629,N_4744);
nand UO_741 (O_741,N_4112,N_4193);
nor UO_742 (O_742,N_4158,N_4985);
or UO_743 (O_743,N_4620,N_4829);
nand UO_744 (O_744,N_4632,N_4789);
or UO_745 (O_745,N_4530,N_4680);
nor UO_746 (O_746,N_4404,N_4284);
and UO_747 (O_747,N_4060,N_4307);
and UO_748 (O_748,N_4347,N_4581);
and UO_749 (O_749,N_4251,N_4596);
or UO_750 (O_750,N_4502,N_4805);
and UO_751 (O_751,N_4742,N_4638);
or UO_752 (O_752,N_4149,N_4611);
nand UO_753 (O_753,N_4122,N_4519);
nand UO_754 (O_754,N_4422,N_4218);
and UO_755 (O_755,N_4713,N_4312);
nand UO_756 (O_756,N_4487,N_4272);
nand UO_757 (O_757,N_4302,N_4715);
and UO_758 (O_758,N_4411,N_4866);
nor UO_759 (O_759,N_4499,N_4194);
nor UO_760 (O_760,N_4692,N_4239);
nor UO_761 (O_761,N_4656,N_4766);
or UO_762 (O_762,N_4763,N_4398);
nor UO_763 (O_763,N_4408,N_4760);
and UO_764 (O_764,N_4741,N_4693);
or UO_765 (O_765,N_4885,N_4337);
nor UO_766 (O_766,N_4437,N_4421);
or UO_767 (O_767,N_4726,N_4741);
and UO_768 (O_768,N_4244,N_4304);
nor UO_769 (O_769,N_4555,N_4581);
and UO_770 (O_770,N_4715,N_4272);
or UO_771 (O_771,N_4703,N_4676);
and UO_772 (O_772,N_4076,N_4401);
and UO_773 (O_773,N_4016,N_4405);
nor UO_774 (O_774,N_4858,N_4516);
nor UO_775 (O_775,N_4635,N_4847);
nor UO_776 (O_776,N_4385,N_4853);
and UO_777 (O_777,N_4186,N_4789);
nand UO_778 (O_778,N_4556,N_4974);
nand UO_779 (O_779,N_4561,N_4813);
and UO_780 (O_780,N_4176,N_4130);
and UO_781 (O_781,N_4047,N_4832);
or UO_782 (O_782,N_4548,N_4335);
and UO_783 (O_783,N_4253,N_4785);
nand UO_784 (O_784,N_4942,N_4530);
and UO_785 (O_785,N_4733,N_4033);
and UO_786 (O_786,N_4436,N_4819);
nor UO_787 (O_787,N_4500,N_4772);
nand UO_788 (O_788,N_4650,N_4367);
nor UO_789 (O_789,N_4942,N_4166);
and UO_790 (O_790,N_4782,N_4552);
and UO_791 (O_791,N_4009,N_4145);
or UO_792 (O_792,N_4315,N_4394);
and UO_793 (O_793,N_4647,N_4565);
nor UO_794 (O_794,N_4625,N_4192);
or UO_795 (O_795,N_4763,N_4042);
and UO_796 (O_796,N_4709,N_4925);
nor UO_797 (O_797,N_4499,N_4740);
nor UO_798 (O_798,N_4045,N_4548);
or UO_799 (O_799,N_4004,N_4986);
nand UO_800 (O_800,N_4105,N_4255);
or UO_801 (O_801,N_4375,N_4850);
nand UO_802 (O_802,N_4377,N_4482);
and UO_803 (O_803,N_4317,N_4627);
nor UO_804 (O_804,N_4518,N_4894);
nor UO_805 (O_805,N_4512,N_4932);
and UO_806 (O_806,N_4610,N_4657);
and UO_807 (O_807,N_4324,N_4597);
and UO_808 (O_808,N_4029,N_4538);
or UO_809 (O_809,N_4504,N_4519);
nand UO_810 (O_810,N_4200,N_4906);
and UO_811 (O_811,N_4912,N_4294);
or UO_812 (O_812,N_4171,N_4968);
nand UO_813 (O_813,N_4449,N_4183);
nor UO_814 (O_814,N_4036,N_4528);
nand UO_815 (O_815,N_4282,N_4495);
and UO_816 (O_816,N_4429,N_4017);
nand UO_817 (O_817,N_4710,N_4940);
nand UO_818 (O_818,N_4216,N_4292);
nor UO_819 (O_819,N_4269,N_4031);
nand UO_820 (O_820,N_4315,N_4043);
nand UO_821 (O_821,N_4915,N_4898);
nor UO_822 (O_822,N_4240,N_4078);
nor UO_823 (O_823,N_4784,N_4401);
nand UO_824 (O_824,N_4657,N_4282);
nand UO_825 (O_825,N_4007,N_4766);
nand UO_826 (O_826,N_4061,N_4753);
and UO_827 (O_827,N_4133,N_4305);
or UO_828 (O_828,N_4308,N_4596);
and UO_829 (O_829,N_4106,N_4600);
xor UO_830 (O_830,N_4227,N_4674);
and UO_831 (O_831,N_4695,N_4102);
nor UO_832 (O_832,N_4267,N_4891);
nand UO_833 (O_833,N_4875,N_4697);
nand UO_834 (O_834,N_4912,N_4573);
or UO_835 (O_835,N_4335,N_4632);
nand UO_836 (O_836,N_4783,N_4889);
or UO_837 (O_837,N_4619,N_4618);
nand UO_838 (O_838,N_4932,N_4767);
nand UO_839 (O_839,N_4332,N_4256);
and UO_840 (O_840,N_4770,N_4465);
or UO_841 (O_841,N_4969,N_4939);
or UO_842 (O_842,N_4343,N_4115);
nor UO_843 (O_843,N_4400,N_4321);
or UO_844 (O_844,N_4749,N_4910);
nor UO_845 (O_845,N_4350,N_4732);
and UO_846 (O_846,N_4077,N_4414);
nor UO_847 (O_847,N_4135,N_4821);
nor UO_848 (O_848,N_4060,N_4270);
and UO_849 (O_849,N_4631,N_4529);
and UO_850 (O_850,N_4704,N_4026);
or UO_851 (O_851,N_4096,N_4276);
nand UO_852 (O_852,N_4429,N_4957);
or UO_853 (O_853,N_4962,N_4232);
nand UO_854 (O_854,N_4796,N_4930);
and UO_855 (O_855,N_4698,N_4649);
nand UO_856 (O_856,N_4868,N_4536);
nand UO_857 (O_857,N_4140,N_4502);
and UO_858 (O_858,N_4189,N_4266);
nor UO_859 (O_859,N_4734,N_4454);
and UO_860 (O_860,N_4133,N_4065);
nor UO_861 (O_861,N_4713,N_4032);
nand UO_862 (O_862,N_4376,N_4136);
or UO_863 (O_863,N_4023,N_4196);
nor UO_864 (O_864,N_4083,N_4716);
nand UO_865 (O_865,N_4833,N_4030);
nor UO_866 (O_866,N_4610,N_4234);
nand UO_867 (O_867,N_4527,N_4630);
nand UO_868 (O_868,N_4487,N_4470);
or UO_869 (O_869,N_4095,N_4410);
nor UO_870 (O_870,N_4411,N_4106);
nor UO_871 (O_871,N_4196,N_4666);
or UO_872 (O_872,N_4284,N_4648);
and UO_873 (O_873,N_4859,N_4253);
and UO_874 (O_874,N_4849,N_4916);
and UO_875 (O_875,N_4663,N_4671);
and UO_876 (O_876,N_4421,N_4564);
and UO_877 (O_877,N_4733,N_4141);
and UO_878 (O_878,N_4112,N_4575);
nor UO_879 (O_879,N_4672,N_4236);
nand UO_880 (O_880,N_4219,N_4227);
or UO_881 (O_881,N_4587,N_4779);
nor UO_882 (O_882,N_4479,N_4439);
and UO_883 (O_883,N_4423,N_4317);
or UO_884 (O_884,N_4386,N_4630);
xor UO_885 (O_885,N_4570,N_4677);
and UO_886 (O_886,N_4038,N_4356);
or UO_887 (O_887,N_4881,N_4048);
and UO_888 (O_888,N_4489,N_4676);
nand UO_889 (O_889,N_4438,N_4014);
and UO_890 (O_890,N_4279,N_4074);
or UO_891 (O_891,N_4309,N_4347);
and UO_892 (O_892,N_4857,N_4621);
and UO_893 (O_893,N_4954,N_4687);
nand UO_894 (O_894,N_4713,N_4100);
nor UO_895 (O_895,N_4660,N_4126);
or UO_896 (O_896,N_4453,N_4852);
nor UO_897 (O_897,N_4926,N_4836);
nand UO_898 (O_898,N_4727,N_4421);
nor UO_899 (O_899,N_4706,N_4550);
nand UO_900 (O_900,N_4239,N_4924);
or UO_901 (O_901,N_4352,N_4630);
or UO_902 (O_902,N_4102,N_4256);
nor UO_903 (O_903,N_4489,N_4047);
nand UO_904 (O_904,N_4677,N_4362);
nand UO_905 (O_905,N_4291,N_4551);
nand UO_906 (O_906,N_4674,N_4487);
nor UO_907 (O_907,N_4519,N_4922);
or UO_908 (O_908,N_4343,N_4956);
nand UO_909 (O_909,N_4205,N_4951);
and UO_910 (O_910,N_4691,N_4676);
or UO_911 (O_911,N_4063,N_4333);
nor UO_912 (O_912,N_4306,N_4102);
and UO_913 (O_913,N_4966,N_4805);
nor UO_914 (O_914,N_4854,N_4382);
or UO_915 (O_915,N_4490,N_4213);
nand UO_916 (O_916,N_4909,N_4618);
or UO_917 (O_917,N_4396,N_4901);
and UO_918 (O_918,N_4743,N_4415);
and UO_919 (O_919,N_4140,N_4663);
nor UO_920 (O_920,N_4174,N_4671);
nor UO_921 (O_921,N_4824,N_4291);
and UO_922 (O_922,N_4874,N_4625);
and UO_923 (O_923,N_4249,N_4724);
nor UO_924 (O_924,N_4252,N_4783);
and UO_925 (O_925,N_4833,N_4529);
or UO_926 (O_926,N_4164,N_4966);
and UO_927 (O_927,N_4425,N_4043);
xnor UO_928 (O_928,N_4233,N_4730);
and UO_929 (O_929,N_4898,N_4247);
and UO_930 (O_930,N_4383,N_4086);
or UO_931 (O_931,N_4969,N_4341);
nor UO_932 (O_932,N_4656,N_4118);
nand UO_933 (O_933,N_4222,N_4514);
or UO_934 (O_934,N_4841,N_4260);
and UO_935 (O_935,N_4421,N_4666);
nor UO_936 (O_936,N_4280,N_4910);
or UO_937 (O_937,N_4143,N_4787);
or UO_938 (O_938,N_4972,N_4069);
and UO_939 (O_939,N_4461,N_4613);
and UO_940 (O_940,N_4072,N_4054);
nand UO_941 (O_941,N_4845,N_4438);
and UO_942 (O_942,N_4271,N_4223);
nand UO_943 (O_943,N_4190,N_4726);
nand UO_944 (O_944,N_4887,N_4905);
or UO_945 (O_945,N_4011,N_4255);
or UO_946 (O_946,N_4096,N_4655);
or UO_947 (O_947,N_4465,N_4816);
nand UO_948 (O_948,N_4190,N_4605);
nor UO_949 (O_949,N_4266,N_4485);
or UO_950 (O_950,N_4005,N_4001);
and UO_951 (O_951,N_4593,N_4586);
nor UO_952 (O_952,N_4292,N_4982);
and UO_953 (O_953,N_4158,N_4753);
and UO_954 (O_954,N_4480,N_4304);
and UO_955 (O_955,N_4002,N_4626);
and UO_956 (O_956,N_4600,N_4898);
nor UO_957 (O_957,N_4908,N_4504);
nand UO_958 (O_958,N_4196,N_4546);
and UO_959 (O_959,N_4660,N_4024);
or UO_960 (O_960,N_4599,N_4420);
nor UO_961 (O_961,N_4782,N_4584);
and UO_962 (O_962,N_4354,N_4111);
nand UO_963 (O_963,N_4422,N_4198);
nor UO_964 (O_964,N_4020,N_4848);
nand UO_965 (O_965,N_4616,N_4596);
nor UO_966 (O_966,N_4224,N_4707);
nand UO_967 (O_967,N_4744,N_4966);
nand UO_968 (O_968,N_4885,N_4263);
nor UO_969 (O_969,N_4899,N_4184);
and UO_970 (O_970,N_4047,N_4391);
nor UO_971 (O_971,N_4746,N_4461);
or UO_972 (O_972,N_4998,N_4353);
or UO_973 (O_973,N_4433,N_4825);
nand UO_974 (O_974,N_4929,N_4263);
nand UO_975 (O_975,N_4255,N_4450);
nand UO_976 (O_976,N_4662,N_4711);
nand UO_977 (O_977,N_4331,N_4692);
nand UO_978 (O_978,N_4767,N_4043);
nand UO_979 (O_979,N_4787,N_4219);
or UO_980 (O_980,N_4478,N_4766);
nor UO_981 (O_981,N_4140,N_4505);
nor UO_982 (O_982,N_4318,N_4055);
nand UO_983 (O_983,N_4623,N_4876);
or UO_984 (O_984,N_4868,N_4919);
or UO_985 (O_985,N_4330,N_4949);
nor UO_986 (O_986,N_4536,N_4288);
or UO_987 (O_987,N_4292,N_4729);
nor UO_988 (O_988,N_4823,N_4866);
nor UO_989 (O_989,N_4792,N_4464);
and UO_990 (O_990,N_4057,N_4832);
and UO_991 (O_991,N_4118,N_4843);
nand UO_992 (O_992,N_4795,N_4554);
and UO_993 (O_993,N_4146,N_4428);
nand UO_994 (O_994,N_4277,N_4689);
nor UO_995 (O_995,N_4550,N_4892);
or UO_996 (O_996,N_4389,N_4452);
nand UO_997 (O_997,N_4516,N_4856);
nor UO_998 (O_998,N_4910,N_4177);
nand UO_999 (O_999,N_4579,N_4400);
endmodule