module basic_750_5000_1000_10_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_385,In_349);
nor U1 (N_1,In_89,In_555);
or U2 (N_2,In_97,In_678);
and U3 (N_3,In_151,In_648);
nor U4 (N_4,In_677,In_410);
nor U5 (N_5,In_531,In_647);
and U6 (N_6,In_163,In_562);
nor U7 (N_7,In_743,In_236);
or U8 (N_8,In_327,In_241);
nand U9 (N_9,In_556,In_144);
nor U10 (N_10,In_464,In_707);
xor U11 (N_11,In_153,In_21);
nand U12 (N_12,In_5,In_364);
and U13 (N_13,In_75,In_428);
nand U14 (N_14,In_246,In_563);
nor U15 (N_15,In_397,In_229);
xor U16 (N_16,In_390,In_198);
xnor U17 (N_17,In_729,In_513);
nand U18 (N_18,In_576,In_25);
xnor U19 (N_19,In_724,In_351);
and U20 (N_20,In_670,In_124);
nand U21 (N_21,In_249,In_704);
xnor U22 (N_22,In_420,In_452);
nand U23 (N_23,In_119,In_736);
nand U24 (N_24,In_67,In_95);
xor U25 (N_25,In_36,In_498);
xor U26 (N_26,In_409,In_393);
nand U27 (N_27,In_612,In_567);
and U28 (N_28,In_40,In_90);
or U29 (N_29,In_642,In_192);
nor U30 (N_30,In_356,In_721);
or U31 (N_31,In_659,In_205);
and U32 (N_32,In_731,In_184);
nor U33 (N_33,In_702,In_510);
or U34 (N_34,In_157,In_109);
or U35 (N_35,In_739,In_256);
or U36 (N_36,In_360,In_221);
xnor U37 (N_37,In_602,In_130);
nor U38 (N_38,In_2,In_311);
xnor U39 (N_39,In_175,In_744);
nand U40 (N_40,In_154,In_0);
nor U41 (N_41,In_231,In_32);
xor U42 (N_42,In_517,In_160);
and U43 (N_43,In_283,In_492);
nor U44 (N_44,In_484,In_732);
nor U45 (N_45,In_518,In_526);
or U46 (N_46,In_133,In_237);
or U47 (N_47,In_714,In_355);
nor U48 (N_48,In_347,In_346);
and U49 (N_49,In_376,In_108);
nor U50 (N_50,In_515,In_554);
nand U51 (N_51,In_323,In_511);
nor U52 (N_52,In_425,In_187);
and U53 (N_53,In_536,In_167);
nor U54 (N_54,In_613,In_651);
nor U55 (N_55,In_73,In_403);
and U56 (N_56,In_593,In_671);
nor U57 (N_57,In_131,In_315);
nor U58 (N_58,In_713,In_418);
xor U59 (N_59,In_245,In_735);
or U60 (N_60,In_462,In_685);
nand U61 (N_61,In_173,In_641);
nand U62 (N_62,In_320,In_127);
or U63 (N_63,In_551,In_111);
xor U64 (N_64,In_599,In_426);
and U65 (N_65,In_379,In_329);
and U66 (N_66,In_527,In_50);
xor U67 (N_67,In_43,In_248);
or U68 (N_68,In_91,In_206);
nor U69 (N_69,In_392,In_533);
nor U70 (N_70,In_478,In_272);
xor U71 (N_71,In_106,In_595);
nand U72 (N_72,In_440,In_645);
nor U73 (N_73,In_208,In_179);
xnor U74 (N_74,In_388,In_460);
xnor U75 (N_75,In_574,In_477);
nor U76 (N_76,In_92,In_522);
and U77 (N_77,In_569,In_530);
xnor U78 (N_78,In_34,In_170);
nand U79 (N_79,In_35,In_416);
nor U80 (N_80,In_367,In_482);
nand U81 (N_81,In_580,In_705);
xnor U82 (N_82,In_453,In_583);
nand U83 (N_83,In_15,In_667);
and U84 (N_84,In_529,In_437);
and U85 (N_85,In_74,In_597);
or U86 (N_86,In_504,In_258);
nand U87 (N_87,In_46,In_373);
nand U88 (N_88,In_299,In_471);
nand U89 (N_89,In_343,In_429);
nand U90 (N_90,In_701,In_342);
nor U91 (N_91,In_550,In_436);
and U92 (N_92,In_745,In_474);
nand U93 (N_93,In_494,In_202);
and U94 (N_94,In_284,In_718);
nor U95 (N_95,In_41,In_115);
nand U96 (N_96,In_145,In_326);
nand U97 (N_97,In_282,In_62);
or U98 (N_98,In_422,In_61);
and U99 (N_99,In_293,In_446);
and U100 (N_100,In_214,In_622);
xor U101 (N_101,In_728,In_266);
and U102 (N_102,In_278,In_480);
nor U103 (N_103,In_166,In_44);
or U104 (N_104,In_263,In_431);
and U105 (N_105,In_340,In_488);
or U106 (N_106,In_414,In_690);
nand U107 (N_107,In_570,In_521);
nor U108 (N_108,In_42,In_472);
xnor U109 (N_109,In_709,In_194);
nor U110 (N_110,In_1,In_85);
and U111 (N_111,In_582,In_372);
or U112 (N_112,In_463,In_378);
nor U113 (N_113,In_338,In_137);
or U114 (N_114,In_423,In_353);
nor U115 (N_115,In_610,In_22);
xor U116 (N_116,In_623,In_618);
xnor U117 (N_117,In_165,In_101);
and U118 (N_118,In_535,In_357);
and U119 (N_119,In_102,In_318);
nor U120 (N_120,In_696,In_455);
nor U121 (N_121,In_55,In_564);
xor U122 (N_122,In_29,In_116);
nor U123 (N_123,In_352,In_719);
or U124 (N_124,In_125,In_686);
and U125 (N_125,In_489,In_501);
and U126 (N_126,In_674,In_681);
nor U127 (N_127,In_708,In_687);
nor U128 (N_128,In_218,In_506);
nor U129 (N_129,In_121,In_395);
and U130 (N_130,In_193,In_658);
nand U131 (N_131,In_128,In_448);
nand U132 (N_132,In_621,In_335);
nor U133 (N_133,In_742,In_139);
nand U134 (N_134,In_306,In_509);
nand U135 (N_135,In_424,In_112);
nand U136 (N_136,In_209,In_331);
nand U137 (N_137,In_457,In_717);
xor U138 (N_138,In_495,In_199);
or U139 (N_139,In_300,In_740);
nand U140 (N_140,In_232,In_538);
and U141 (N_141,In_325,In_262);
xor U142 (N_142,In_485,In_662);
and U143 (N_143,In_230,In_546);
or U144 (N_144,In_666,In_552);
xnor U145 (N_145,In_454,In_224);
nor U146 (N_146,In_348,In_573);
nand U147 (N_147,In_247,In_726);
or U148 (N_148,In_432,In_496);
xnor U149 (N_149,In_142,In_60);
and U150 (N_150,In_171,In_688);
or U151 (N_151,In_358,In_223);
nor U152 (N_152,In_449,In_656);
nand U153 (N_153,In_103,In_254);
or U154 (N_154,In_211,In_534);
nand U155 (N_155,In_375,In_543);
nand U156 (N_156,In_703,In_673);
or U157 (N_157,In_11,In_277);
or U158 (N_158,In_596,In_640);
nand U159 (N_159,In_514,In_722);
nor U160 (N_160,In_313,In_628);
and U161 (N_161,In_560,In_456);
nand U162 (N_162,In_730,In_7);
xor U163 (N_163,In_606,In_191);
nor U164 (N_164,In_694,In_541);
and U165 (N_165,In_201,In_113);
or U166 (N_166,In_636,In_250);
nand U167 (N_167,In_207,In_720);
nor U168 (N_168,In_695,In_143);
nor U169 (N_169,In_684,In_324);
xor U170 (N_170,In_441,In_459);
and U171 (N_171,In_319,In_407);
and U172 (N_172,In_304,In_465);
or U173 (N_173,In_438,In_401);
and U174 (N_174,In_51,In_333);
and U175 (N_175,In_747,In_123);
nor U176 (N_176,In_734,In_575);
xor U177 (N_177,In_217,In_9);
nor U178 (N_178,In_345,In_512);
nand U179 (N_179,In_159,In_607);
or U180 (N_180,In_675,In_491);
or U181 (N_181,In_430,In_244);
nand U182 (N_182,In_68,In_156);
xor U183 (N_183,In_447,In_565);
and U184 (N_184,In_104,In_483);
nor U185 (N_185,In_174,In_56);
xnor U186 (N_186,In_627,In_408);
xnor U187 (N_187,In_99,In_136);
nor U188 (N_188,In_86,In_233);
xnor U189 (N_189,In_289,In_605);
xnor U190 (N_190,In_679,In_317);
nand U191 (N_191,In_503,In_519);
and U192 (N_192,In_391,In_261);
and U193 (N_193,In_267,In_697);
xnor U194 (N_194,In_81,In_28);
nor U195 (N_195,In_350,In_138);
nor U196 (N_196,In_65,In_365);
nand U197 (N_197,In_520,In_499);
xnor U198 (N_198,In_680,In_88);
nand U199 (N_199,In_663,In_589);
and U200 (N_200,In_322,In_332);
or U201 (N_201,In_152,In_100);
xor U202 (N_202,In_302,In_197);
xnor U203 (N_203,In_698,In_611);
nor U204 (N_204,In_490,In_181);
or U205 (N_205,In_377,In_362);
nand U206 (N_206,In_107,In_646);
or U207 (N_207,In_727,In_337);
nor U208 (N_208,In_310,In_644);
xor U209 (N_209,In_204,In_616);
xor U210 (N_210,In_638,In_203);
or U211 (N_211,In_110,In_53);
nand U212 (N_212,In_712,In_434);
or U213 (N_213,In_316,In_660);
nand U214 (N_214,In_733,In_683);
nor U215 (N_215,In_84,In_265);
nand U216 (N_216,In_445,In_126);
nand U217 (N_217,In_330,In_291);
xnor U218 (N_218,In_195,In_451);
xnor U219 (N_219,In_654,In_396);
nor U220 (N_220,In_69,In_336);
nand U221 (N_221,In_502,In_132);
xnor U222 (N_222,In_213,In_286);
and U223 (N_223,In_461,In_706);
xor U224 (N_224,In_234,In_17);
or U225 (N_225,In_587,In_711);
and U226 (N_226,In_162,In_274);
or U227 (N_227,In_30,In_52);
or U228 (N_228,In_251,In_23);
xor U229 (N_229,In_285,In_31);
nand U230 (N_230,In_94,In_279);
xor U231 (N_231,In_406,In_264);
or U232 (N_232,In_389,In_309);
nor U233 (N_233,In_295,In_83);
xor U234 (N_234,In_273,In_435);
or U235 (N_235,In_24,In_158);
or U236 (N_236,In_558,In_415);
or U237 (N_237,In_59,In_118);
nor U238 (N_238,In_450,In_633);
nand U239 (N_239,In_476,In_553);
nor U240 (N_240,In_399,In_466);
nand U241 (N_241,In_296,In_544);
xor U242 (N_242,In_269,In_693);
xnor U243 (N_243,In_585,In_172);
nand U244 (N_244,In_243,In_14);
nor U245 (N_245,In_114,In_72);
and U246 (N_246,In_182,In_668);
nor U247 (N_247,In_196,In_87);
xnor U248 (N_248,In_467,In_164);
nor U249 (N_249,In_584,In_240);
nor U250 (N_250,In_168,In_559);
nor U251 (N_251,In_470,In_242);
nor U252 (N_252,In_63,In_594);
nor U253 (N_253,In_307,In_444);
or U254 (N_254,In_412,In_228);
and U255 (N_255,In_486,In_66);
xor U256 (N_256,In_371,In_312);
or U257 (N_257,In_215,In_691);
nand U258 (N_258,In_620,In_18);
nand U259 (N_259,In_297,In_443);
and U260 (N_260,In_657,In_481);
xor U261 (N_261,In_598,In_253);
or U262 (N_262,In_614,In_652);
xor U263 (N_263,In_746,In_98);
nor U264 (N_264,In_637,In_540);
nor U265 (N_265,In_661,In_79);
xnor U266 (N_266,In_615,In_524);
xor U267 (N_267,In_417,In_148);
xor U268 (N_268,In_186,In_117);
or U269 (N_269,In_16,In_146);
nand U270 (N_270,In_542,In_58);
or U271 (N_271,In_147,In_608);
nand U272 (N_272,In_402,In_479);
or U273 (N_273,In_368,In_252);
and U274 (N_274,In_47,In_354);
and U275 (N_275,In_366,In_442);
nor U276 (N_276,In_601,In_38);
or U277 (N_277,In_287,In_624);
nor U278 (N_278,In_737,In_275);
nor U279 (N_279,In_54,In_625);
xnor U280 (N_280,In_634,In_292);
xor U281 (N_281,In_6,In_8);
or U282 (N_282,In_400,In_27);
or U283 (N_283,In_692,In_225);
nand U284 (N_284,In_643,In_141);
nand U285 (N_285,In_57,In_493);
nand U286 (N_286,In_222,In_588);
or U287 (N_287,In_571,In_568);
xnor U288 (N_288,In_71,In_321);
or U289 (N_289,In_382,In_290);
or U290 (N_290,In_689,In_458);
xnor U291 (N_291,In_155,In_268);
nor U292 (N_292,In_609,In_185);
or U293 (N_293,In_150,In_664);
nor U294 (N_294,In_178,In_586);
nand U295 (N_295,In_314,In_339);
and U296 (N_296,In_539,In_305);
nand U297 (N_297,In_129,In_619);
nor U298 (N_298,In_227,In_134);
xor U299 (N_299,In_93,In_226);
and U300 (N_300,In_547,In_183);
nor U301 (N_301,In_626,In_169);
and U302 (N_302,In_37,In_303);
nor U303 (N_303,In_255,In_120);
nand U304 (N_304,In_433,In_374);
and U305 (N_305,In_308,In_188);
or U306 (N_306,In_3,In_96);
and U307 (N_307,In_592,In_363);
nand U308 (N_308,In_149,In_655);
and U309 (N_309,In_700,In_180);
xnor U310 (N_310,In_508,In_48);
and U311 (N_311,In_591,In_653);
nand U312 (N_312,In_411,In_725);
or U313 (N_313,In_549,In_715);
or U314 (N_314,In_548,In_600);
and U315 (N_315,In_523,In_405);
and U316 (N_316,In_45,In_649);
nor U317 (N_317,In_77,In_419);
or U318 (N_318,In_238,In_259);
nand U319 (N_319,In_212,In_280);
and U320 (N_320,In_176,In_19);
nor U321 (N_321,In_545,In_64);
or U322 (N_322,In_676,In_384);
and U323 (N_323,In_26,In_682);
and U324 (N_324,In_260,In_581);
xnor U325 (N_325,In_632,In_473);
nor U326 (N_326,In_161,In_257);
nor U327 (N_327,In_383,In_672);
nand U328 (N_328,In_723,In_468);
nand U329 (N_329,In_710,In_13);
and U330 (N_330,In_216,In_344);
or U331 (N_331,In_394,In_122);
xor U332 (N_332,In_190,In_487);
nor U333 (N_333,In_572,In_639);
nand U334 (N_334,In_421,In_537);
and U335 (N_335,In_528,In_387);
nand U336 (N_336,In_220,In_525);
nand U337 (N_337,In_78,In_239);
nor U338 (N_338,In_386,In_276);
nand U339 (N_339,In_497,In_70);
xor U340 (N_340,In_4,In_271);
nor U341 (N_341,In_748,In_635);
nor U342 (N_342,In_189,In_500);
xnor U343 (N_343,In_370,In_469);
nand U344 (N_344,In_33,In_359);
xor U345 (N_345,In_413,In_235);
nor U346 (N_346,In_369,In_80);
or U347 (N_347,In_475,In_629);
nor U348 (N_348,In_578,In_381);
xor U349 (N_349,In_10,In_749);
or U350 (N_350,In_140,In_76);
xnor U351 (N_351,In_532,In_219);
xnor U352 (N_352,In_294,In_604);
and U353 (N_353,In_603,In_631);
or U354 (N_354,In_507,In_361);
and U355 (N_355,In_699,In_738);
nand U356 (N_356,In_404,In_49);
or U357 (N_357,In_341,In_328);
nand U358 (N_358,In_12,In_590);
or U359 (N_359,In_716,In_516);
nor U360 (N_360,In_505,In_105);
nor U361 (N_361,In_439,In_380);
or U362 (N_362,In_177,In_270);
nor U363 (N_363,In_665,In_566);
nor U364 (N_364,In_741,In_427);
and U365 (N_365,In_650,In_669);
and U366 (N_366,In_630,In_579);
xor U367 (N_367,In_577,In_561);
or U368 (N_368,In_20,In_301);
and U369 (N_369,In_210,In_200);
or U370 (N_370,In_82,In_39);
xnor U371 (N_371,In_617,In_288);
nand U372 (N_372,In_334,In_298);
and U373 (N_373,In_135,In_557);
or U374 (N_374,In_281,In_398);
and U375 (N_375,In_568,In_498);
nand U376 (N_376,In_339,In_32);
nor U377 (N_377,In_622,In_21);
and U378 (N_378,In_737,In_520);
and U379 (N_379,In_233,In_159);
nand U380 (N_380,In_628,In_138);
xor U381 (N_381,In_200,In_59);
nor U382 (N_382,In_565,In_351);
and U383 (N_383,In_373,In_553);
nor U384 (N_384,In_109,In_445);
nor U385 (N_385,In_360,In_209);
nand U386 (N_386,In_598,In_695);
xnor U387 (N_387,In_81,In_571);
xnor U388 (N_388,In_97,In_446);
and U389 (N_389,In_374,In_384);
nor U390 (N_390,In_32,In_160);
nand U391 (N_391,In_229,In_406);
and U392 (N_392,In_138,In_305);
nor U393 (N_393,In_682,In_262);
and U394 (N_394,In_283,In_739);
and U395 (N_395,In_604,In_709);
and U396 (N_396,In_281,In_606);
xnor U397 (N_397,In_474,In_167);
or U398 (N_398,In_76,In_203);
nor U399 (N_399,In_325,In_598);
and U400 (N_400,In_396,In_61);
and U401 (N_401,In_743,In_237);
nor U402 (N_402,In_288,In_314);
nand U403 (N_403,In_412,In_61);
and U404 (N_404,In_303,In_250);
and U405 (N_405,In_287,In_710);
nand U406 (N_406,In_56,In_468);
xnor U407 (N_407,In_702,In_323);
nor U408 (N_408,In_110,In_708);
or U409 (N_409,In_629,In_535);
nor U410 (N_410,In_441,In_309);
xor U411 (N_411,In_698,In_163);
xnor U412 (N_412,In_689,In_577);
or U413 (N_413,In_0,In_149);
or U414 (N_414,In_472,In_155);
nor U415 (N_415,In_302,In_148);
and U416 (N_416,In_639,In_132);
nor U417 (N_417,In_394,In_94);
nor U418 (N_418,In_309,In_297);
and U419 (N_419,In_693,In_661);
or U420 (N_420,In_156,In_88);
and U421 (N_421,In_689,In_722);
nand U422 (N_422,In_154,In_501);
and U423 (N_423,In_645,In_533);
or U424 (N_424,In_51,In_313);
nor U425 (N_425,In_386,In_511);
nand U426 (N_426,In_34,In_403);
xnor U427 (N_427,In_573,In_585);
xor U428 (N_428,In_315,In_31);
xor U429 (N_429,In_271,In_206);
nor U430 (N_430,In_485,In_658);
and U431 (N_431,In_521,In_723);
and U432 (N_432,In_287,In_697);
or U433 (N_433,In_556,In_359);
and U434 (N_434,In_366,In_324);
or U435 (N_435,In_642,In_641);
or U436 (N_436,In_302,In_534);
nand U437 (N_437,In_724,In_171);
and U438 (N_438,In_395,In_460);
xnor U439 (N_439,In_373,In_681);
and U440 (N_440,In_673,In_618);
and U441 (N_441,In_718,In_366);
nor U442 (N_442,In_3,In_708);
nand U443 (N_443,In_88,In_465);
and U444 (N_444,In_714,In_108);
and U445 (N_445,In_200,In_11);
and U446 (N_446,In_711,In_164);
and U447 (N_447,In_717,In_420);
and U448 (N_448,In_446,In_710);
or U449 (N_449,In_310,In_33);
nor U450 (N_450,In_665,In_348);
nor U451 (N_451,In_464,In_360);
and U452 (N_452,In_462,In_108);
nor U453 (N_453,In_25,In_374);
or U454 (N_454,In_420,In_533);
xnor U455 (N_455,In_722,In_637);
nand U456 (N_456,In_355,In_224);
and U457 (N_457,In_199,In_74);
or U458 (N_458,In_681,In_332);
nor U459 (N_459,In_24,In_429);
nor U460 (N_460,In_470,In_589);
nor U461 (N_461,In_630,In_469);
and U462 (N_462,In_359,In_745);
or U463 (N_463,In_499,In_605);
nand U464 (N_464,In_325,In_299);
or U465 (N_465,In_156,In_253);
and U466 (N_466,In_443,In_543);
and U467 (N_467,In_372,In_587);
nand U468 (N_468,In_228,In_398);
nand U469 (N_469,In_304,In_566);
or U470 (N_470,In_129,In_21);
xnor U471 (N_471,In_95,In_521);
and U472 (N_472,In_378,In_704);
or U473 (N_473,In_490,In_608);
xor U474 (N_474,In_301,In_637);
xor U475 (N_475,In_534,In_539);
or U476 (N_476,In_36,In_625);
nand U477 (N_477,In_625,In_364);
nor U478 (N_478,In_211,In_457);
nor U479 (N_479,In_78,In_664);
and U480 (N_480,In_700,In_150);
nand U481 (N_481,In_185,In_146);
nand U482 (N_482,In_100,In_196);
nand U483 (N_483,In_311,In_475);
xor U484 (N_484,In_418,In_721);
and U485 (N_485,In_513,In_337);
nor U486 (N_486,In_143,In_545);
or U487 (N_487,In_703,In_285);
and U488 (N_488,In_257,In_256);
and U489 (N_489,In_306,In_713);
xor U490 (N_490,In_307,In_117);
or U491 (N_491,In_180,In_524);
and U492 (N_492,In_325,In_54);
nor U493 (N_493,In_21,In_623);
or U494 (N_494,In_351,In_362);
nor U495 (N_495,In_349,In_191);
or U496 (N_496,In_208,In_383);
nand U497 (N_497,In_404,In_28);
nand U498 (N_498,In_243,In_300);
nand U499 (N_499,In_186,In_160);
or U500 (N_500,N_442,N_430);
nor U501 (N_501,N_77,N_449);
and U502 (N_502,N_226,N_433);
and U503 (N_503,N_376,N_141);
or U504 (N_504,N_227,N_155);
or U505 (N_505,N_56,N_211);
xnor U506 (N_506,N_159,N_216);
nor U507 (N_507,N_69,N_229);
or U508 (N_508,N_112,N_225);
or U509 (N_509,N_328,N_8);
nand U510 (N_510,N_489,N_40);
or U511 (N_511,N_438,N_395);
nor U512 (N_512,N_4,N_465);
xor U513 (N_513,N_342,N_463);
xnor U514 (N_514,N_308,N_158);
and U515 (N_515,N_235,N_70);
nor U516 (N_516,N_99,N_486);
or U517 (N_517,N_475,N_209);
and U518 (N_518,N_387,N_111);
and U519 (N_519,N_150,N_423);
or U520 (N_520,N_264,N_372);
nor U521 (N_521,N_445,N_176);
or U522 (N_522,N_300,N_9);
xnor U523 (N_523,N_31,N_467);
xnor U524 (N_524,N_139,N_146);
and U525 (N_525,N_114,N_335);
xor U526 (N_526,N_196,N_205);
nand U527 (N_527,N_237,N_456);
and U528 (N_528,N_58,N_307);
and U529 (N_529,N_393,N_137);
and U530 (N_530,N_50,N_177);
nor U531 (N_531,N_431,N_116);
and U532 (N_532,N_283,N_459);
nand U533 (N_533,N_418,N_461);
nor U534 (N_534,N_364,N_254);
and U535 (N_535,N_419,N_224);
and U536 (N_536,N_66,N_12);
xnor U537 (N_537,N_240,N_468);
xor U538 (N_538,N_101,N_331);
xnor U539 (N_539,N_106,N_219);
nand U540 (N_540,N_87,N_255);
and U541 (N_541,N_36,N_143);
nand U542 (N_542,N_194,N_276);
nand U543 (N_543,N_161,N_398);
xnor U544 (N_544,N_414,N_29);
nor U545 (N_545,N_244,N_178);
or U546 (N_546,N_274,N_166);
and U547 (N_547,N_53,N_440);
nand U548 (N_548,N_422,N_492);
and U549 (N_549,N_351,N_97);
xnor U550 (N_550,N_265,N_243);
nand U551 (N_551,N_291,N_282);
nand U552 (N_552,N_201,N_415);
xnor U553 (N_553,N_168,N_370);
nand U554 (N_554,N_96,N_491);
nor U555 (N_555,N_73,N_409);
nand U556 (N_556,N_51,N_380);
nor U557 (N_557,N_144,N_83);
xor U558 (N_558,N_470,N_91);
or U559 (N_559,N_242,N_284);
or U560 (N_560,N_295,N_251);
or U561 (N_561,N_474,N_499);
nand U562 (N_562,N_374,N_426);
or U563 (N_563,N_213,N_175);
or U564 (N_564,N_82,N_90);
nor U565 (N_565,N_234,N_454);
nand U566 (N_566,N_262,N_68);
and U567 (N_567,N_173,N_202);
nor U568 (N_568,N_340,N_30);
nand U569 (N_569,N_256,N_286);
nor U570 (N_570,N_294,N_15);
xor U571 (N_571,N_287,N_94);
or U572 (N_572,N_352,N_304);
xnor U573 (N_573,N_154,N_133);
nand U574 (N_574,N_420,N_65);
and U575 (N_575,N_306,N_93);
or U576 (N_576,N_153,N_52);
nor U577 (N_577,N_165,N_183);
nor U578 (N_578,N_182,N_359);
and U579 (N_579,N_221,N_273);
and U580 (N_580,N_488,N_441);
nand U581 (N_581,N_487,N_190);
and U582 (N_582,N_281,N_115);
xnor U583 (N_583,N_476,N_13);
nand U584 (N_584,N_483,N_267);
nor U585 (N_585,N_21,N_271);
xor U586 (N_586,N_85,N_71);
nand U587 (N_587,N_322,N_92);
nor U588 (N_588,N_394,N_45);
nand U589 (N_589,N_403,N_479);
or U590 (N_590,N_54,N_428);
or U591 (N_591,N_98,N_347);
and U592 (N_592,N_135,N_105);
and U593 (N_593,N_494,N_381);
and U594 (N_594,N_471,N_493);
nor U595 (N_595,N_390,N_130);
nand U596 (N_596,N_388,N_341);
and U597 (N_597,N_43,N_278);
nand U598 (N_598,N_206,N_32);
nand U599 (N_599,N_49,N_41);
or U600 (N_600,N_301,N_186);
and U601 (N_601,N_113,N_349);
or U602 (N_602,N_171,N_360);
nand U603 (N_603,N_411,N_373);
xnor U604 (N_604,N_314,N_356);
or U605 (N_605,N_315,N_353);
and U606 (N_606,N_95,N_263);
and U607 (N_607,N_110,N_193);
or U608 (N_608,N_1,N_18);
xor U609 (N_609,N_378,N_312);
or U610 (N_610,N_417,N_148);
nand U611 (N_611,N_246,N_446);
nand U612 (N_612,N_218,N_38);
xor U613 (N_613,N_134,N_167);
nand U614 (N_614,N_236,N_37);
or U615 (N_615,N_245,N_107);
nand U616 (N_616,N_198,N_421);
or U617 (N_617,N_19,N_76);
xnor U618 (N_618,N_402,N_371);
and U619 (N_619,N_197,N_412);
or U620 (N_620,N_129,N_89);
or U621 (N_621,N_121,N_311);
nand U622 (N_622,N_140,N_24);
nand U623 (N_623,N_406,N_103);
xnor U624 (N_624,N_354,N_270);
or U625 (N_625,N_361,N_350);
or U626 (N_626,N_207,N_313);
nor U627 (N_627,N_338,N_214);
nand U628 (N_628,N_248,N_253);
or U629 (N_629,N_60,N_252);
nand U630 (N_630,N_132,N_118);
nor U631 (N_631,N_386,N_321);
nand U632 (N_632,N_450,N_44);
nor U633 (N_633,N_337,N_138);
and U634 (N_634,N_407,N_309);
nand U635 (N_635,N_266,N_443);
and U636 (N_636,N_455,N_416);
or U637 (N_637,N_289,N_277);
xor U638 (N_638,N_170,N_310);
nor U639 (N_639,N_195,N_377);
xor U640 (N_640,N_151,N_79);
and U641 (N_641,N_128,N_27);
nor U642 (N_642,N_185,N_67);
nor U643 (N_643,N_123,N_28);
nand U644 (N_644,N_192,N_203);
and U645 (N_645,N_452,N_444);
xnor U646 (N_646,N_318,N_429);
nor U647 (N_647,N_346,N_320);
or U648 (N_648,N_391,N_34);
or U649 (N_649,N_464,N_14);
or U650 (N_650,N_482,N_292);
nand U651 (N_651,N_484,N_239);
and U652 (N_652,N_261,N_220);
and U653 (N_653,N_343,N_184);
or U654 (N_654,N_212,N_208);
and U655 (N_655,N_457,N_258);
nand U656 (N_656,N_358,N_233);
or U657 (N_657,N_180,N_327);
and U658 (N_658,N_222,N_448);
and U659 (N_659,N_247,N_339);
or U660 (N_660,N_108,N_188);
nor U661 (N_661,N_250,N_490);
or U662 (N_662,N_0,N_432);
and U663 (N_663,N_147,N_319);
xor U664 (N_664,N_120,N_157);
nand U665 (N_665,N_472,N_458);
nand U666 (N_666,N_480,N_259);
nor U667 (N_667,N_232,N_392);
and U668 (N_668,N_189,N_316);
and U669 (N_669,N_303,N_57);
nor U670 (N_670,N_33,N_109);
xnor U671 (N_671,N_136,N_437);
nand U672 (N_672,N_39,N_384);
xnor U673 (N_673,N_477,N_498);
xor U674 (N_674,N_496,N_404);
and U675 (N_675,N_163,N_149);
nand U676 (N_676,N_413,N_23);
xor U677 (N_677,N_397,N_326);
or U678 (N_678,N_344,N_174);
and U679 (N_679,N_230,N_362);
or U680 (N_680,N_305,N_187);
xnor U681 (N_681,N_334,N_401);
or U682 (N_682,N_400,N_323);
or U683 (N_683,N_325,N_399);
xor U684 (N_684,N_238,N_299);
and U685 (N_685,N_62,N_363);
or U686 (N_686,N_481,N_466);
and U687 (N_687,N_462,N_332);
nor U688 (N_688,N_86,N_22);
or U689 (N_689,N_17,N_317);
nand U690 (N_690,N_434,N_25);
nor U691 (N_691,N_425,N_279);
and U692 (N_692,N_366,N_81);
or U693 (N_693,N_64,N_88);
and U694 (N_694,N_336,N_497);
xor U695 (N_695,N_61,N_293);
or U696 (N_696,N_329,N_10);
xnor U697 (N_697,N_427,N_383);
and U698 (N_698,N_275,N_210);
and U699 (N_699,N_160,N_75);
xor U700 (N_700,N_348,N_125);
xnor U701 (N_701,N_59,N_478);
and U702 (N_702,N_389,N_48);
xor U703 (N_703,N_78,N_280);
and U704 (N_704,N_124,N_269);
or U705 (N_705,N_288,N_72);
nor U706 (N_706,N_495,N_80);
and U707 (N_707,N_126,N_42);
and U708 (N_708,N_345,N_228);
nand U709 (N_709,N_268,N_297);
and U710 (N_710,N_298,N_410);
or U711 (N_711,N_16,N_473);
nor U712 (N_712,N_302,N_324);
and U713 (N_713,N_285,N_367);
or U714 (N_714,N_5,N_257);
nor U715 (N_715,N_451,N_35);
nor U716 (N_716,N_199,N_84);
xnor U717 (N_717,N_290,N_47);
nor U718 (N_718,N_355,N_131);
xor U719 (N_719,N_382,N_122);
and U720 (N_720,N_179,N_330);
xor U721 (N_721,N_357,N_162);
nand U722 (N_722,N_368,N_215);
and U723 (N_723,N_439,N_104);
xor U724 (N_724,N_164,N_436);
or U725 (N_725,N_204,N_249);
nor U726 (N_726,N_375,N_7);
nand U727 (N_727,N_63,N_55);
and U728 (N_728,N_396,N_453);
xor U729 (N_729,N_26,N_379);
nor U730 (N_730,N_117,N_172);
nand U731 (N_731,N_6,N_100);
xor U732 (N_732,N_447,N_191);
nor U733 (N_733,N_260,N_119);
xnor U734 (N_734,N_156,N_74);
and U735 (N_735,N_223,N_424);
xor U736 (N_736,N_460,N_3);
xor U737 (N_737,N_369,N_127);
xor U738 (N_738,N_2,N_142);
nand U739 (N_739,N_46,N_485);
and U740 (N_740,N_469,N_408);
or U741 (N_741,N_217,N_145);
or U742 (N_742,N_241,N_405);
nor U743 (N_743,N_231,N_20);
nand U744 (N_744,N_11,N_385);
and U745 (N_745,N_333,N_102);
nand U746 (N_746,N_200,N_169);
or U747 (N_747,N_272,N_181);
or U748 (N_748,N_152,N_435);
nand U749 (N_749,N_296,N_365);
nor U750 (N_750,N_52,N_301);
nand U751 (N_751,N_432,N_257);
nand U752 (N_752,N_474,N_372);
xor U753 (N_753,N_420,N_53);
or U754 (N_754,N_434,N_408);
nor U755 (N_755,N_205,N_225);
or U756 (N_756,N_156,N_474);
xnor U757 (N_757,N_101,N_305);
nor U758 (N_758,N_434,N_114);
and U759 (N_759,N_187,N_475);
or U760 (N_760,N_117,N_160);
nand U761 (N_761,N_163,N_159);
and U762 (N_762,N_51,N_193);
or U763 (N_763,N_255,N_439);
and U764 (N_764,N_310,N_158);
nand U765 (N_765,N_161,N_60);
and U766 (N_766,N_64,N_267);
or U767 (N_767,N_61,N_82);
and U768 (N_768,N_424,N_484);
xnor U769 (N_769,N_408,N_209);
nand U770 (N_770,N_48,N_495);
xnor U771 (N_771,N_36,N_17);
nand U772 (N_772,N_256,N_385);
nand U773 (N_773,N_431,N_94);
xnor U774 (N_774,N_193,N_457);
nor U775 (N_775,N_174,N_325);
and U776 (N_776,N_447,N_441);
nor U777 (N_777,N_265,N_115);
or U778 (N_778,N_32,N_128);
and U779 (N_779,N_21,N_208);
xor U780 (N_780,N_273,N_432);
or U781 (N_781,N_301,N_282);
xor U782 (N_782,N_175,N_281);
xor U783 (N_783,N_60,N_438);
nor U784 (N_784,N_96,N_117);
nand U785 (N_785,N_343,N_447);
nand U786 (N_786,N_171,N_324);
xor U787 (N_787,N_114,N_348);
xor U788 (N_788,N_447,N_194);
or U789 (N_789,N_95,N_88);
and U790 (N_790,N_183,N_363);
nor U791 (N_791,N_63,N_234);
xnor U792 (N_792,N_354,N_271);
xnor U793 (N_793,N_302,N_401);
or U794 (N_794,N_193,N_493);
nand U795 (N_795,N_401,N_49);
nand U796 (N_796,N_439,N_10);
nand U797 (N_797,N_433,N_142);
and U798 (N_798,N_46,N_179);
nor U799 (N_799,N_45,N_216);
xor U800 (N_800,N_124,N_373);
nand U801 (N_801,N_306,N_406);
nor U802 (N_802,N_331,N_134);
or U803 (N_803,N_428,N_381);
or U804 (N_804,N_169,N_358);
and U805 (N_805,N_478,N_356);
xnor U806 (N_806,N_229,N_238);
xnor U807 (N_807,N_434,N_91);
and U808 (N_808,N_21,N_82);
xnor U809 (N_809,N_395,N_379);
xnor U810 (N_810,N_170,N_219);
nand U811 (N_811,N_278,N_86);
nor U812 (N_812,N_103,N_106);
or U813 (N_813,N_96,N_420);
nand U814 (N_814,N_62,N_217);
and U815 (N_815,N_284,N_429);
xor U816 (N_816,N_164,N_304);
and U817 (N_817,N_143,N_38);
and U818 (N_818,N_265,N_489);
or U819 (N_819,N_235,N_84);
xnor U820 (N_820,N_159,N_481);
nand U821 (N_821,N_362,N_222);
nor U822 (N_822,N_176,N_228);
xnor U823 (N_823,N_186,N_259);
or U824 (N_824,N_318,N_465);
nand U825 (N_825,N_10,N_231);
nand U826 (N_826,N_403,N_280);
or U827 (N_827,N_213,N_143);
or U828 (N_828,N_248,N_390);
xnor U829 (N_829,N_1,N_250);
or U830 (N_830,N_164,N_132);
and U831 (N_831,N_418,N_393);
nand U832 (N_832,N_77,N_454);
nand U833 (N_833,N_101,N_84);
nand U834 (N_834,N_213,N_337);
nor U835 (N_835,N_223,N_436);
xor U836 (N_836,N_152,N_96);
xnor U837 (N_837,N_46,N_54);
or U838 (N_838,N_166,N_254);
xnor U839 (N_839,N_483,N_128);
xnor U840 (N_840,N_348,N_230);
nand U841 (N_841,N_358,N_360);
and U842 (N_842,N_382,N_371);
nor U843 (N_843,N_304,N_74);
nand U844 (N_844,N_15,N_133);
nand U845 (N_845,N_128,N_446);
and U846 (N_846,N_8,N_498);
xnor U847 (N_847,N_225,N_111);
or U848 (N_848,N_249,N_104);
and U849 (N_849,N_355,N_440);
nor U850 (N_850,N_398,N_353);
or U851 (N_851,N_127,N_288);
or U852 (N_852,N_40,N_26);
and U853 (N_853,N_148,N_405);
xor U854 (N_854,N_337,N_3);
xor U855 (N_855,N_160,N_422);
and U856 (N_856,N_89,N_357);
nand U857 (N_857,N_245,N_320);
xor U858 (N_858,N_188,N_82);
xor U859 (N_859,N_377,N_465);
nor U860 (N_860,N_236,N_312);
xnor U861 (N_861,N_341,N_198);
nor U862 (N_862,N_472,N_278);
or U863 (N_863,N_372,N_299);
or U864 (N_864,N_30,N_243);
xor U865 (N_865,N_143,N_217);
or U866 (N_866,N_145,N_465);
or U867 (N_867,N_168,N_40);
or U868 (N_868,N_259,N_217);
nor U869 (N_869,N_174,N_153);
and U870 (N_870,N_198,N_221);
or U871 (N_871,N_71,N_160);
and U872 (N_872,N_408,N_200);
or U873 (N_873,N_305,N_159);
and U874 (N_874,N_405,N_239);
or U875 (N_875,N_185,N_321);
or U876 (N_876,N_224,N_98);
nand U877 (N_877,N_156,N_366);
xnor U878 (N_878,N_165,N_48);
and U879 (N_879,N_312,N_219);
and U880 (N_880,N_289,N_349);
and U881 (N_881,N_39,N_403);
nor U882 (N_882,N_434,N_252);
or U883 (N_883,N_65,N_484);
xor U884 (N_884,N_268,N_110);
nand U885 (N_885,N_206,N_452);
xnor U886 (N_886,N_233,N_131);
nor U887 (N_887,N_271,N_352);
xnor U888 (N_888,N_287,N_175);
nand U889 (N_889,N_372,N_374);
and U890 (N_890,N_302,N_474);
or U891 (N_891,N_453,N_482);
or U892 (N_892,N_76,N_12);
and U893 (N_893,N_274,N_109);
and U894 (N_894,N_323,N_456);
xnor U895 (N_895,N_464,N_347);
nor U896 (N_896,N_217,N_109);
nand U897 (N_897,N_143,N_244);
nor U898 (N_898,N_470,N_352);
nor U899 (N_899,N_164,N_477);
or U900 (N_900,N_116,N_313);
or U901 (N_901,N_165,N_189);
nand U902 (N_902,N_287,N_25);
and U903 (N_903,N_86,N_205);
or U904 (N_904,N_80,N_422);
and U905 (N_905,N_240,N_479);
xor U906 (N_906,N_15,N_58);
nor U907 (N_907,N_253,N_401);
nand U908 (N_908,N_102,N_315);
or U909 (N_909,N_398,N_117);
xor U910 (N_910,N_446,N_160);
nand U911 (N_911,N_153,N_411);
nor U912 (N_912,N_180,N_72);
nor U913 (N_913,N_135,N_221);
or U914 (N_914,N_171,N_434);
or U915 (N_915,N_0,N_7);
or U916 (N_916,N_143,N_468);
or U917 (N_917,N_334,N_155);
nand U918 (N_918,N_148,N_147);
nand U919 (N_919,N_437,N_30);
or U920 (N_920,N_35,N_59);
nand U921 (N_921,N_192,N_281);
xor U922 (N_922,N_391,N_237);
nor U923 (N_923,N_425,N_180);
xnor U924 (N_924,N_253,N_278);
and U925 (N_925,N_477,N_86);
or U926 (N_926,N_409,N_65);
and U927 (N_927,N_201,N_411);
nand U928 (N_928,N_333,N_281);
xnor U929 (N_929,N_206,N_444);
nand U930 (N_930,N_282,N_64);
nand U931 (N_931,N_2,N_96);
xor U932 (N_932,N_470,N_382);
or U933 (N_933,N_349,N_177);
or U934 (N_934,N_153,N_30);
and U935 (N_935,N_236,N_126);
and U936 (N_936,N_113,N_372);
or U937 (N_937,N_182,N_360);
nor U938 (N_938,N_71,N_359);
xor U939 (N_939,N_343,N_56);
and U940 (N_940,N_458,N_266);
nand U941 (N_941,N_475,N_140);
or U942 (N_942,N_145,N_344);
and U943 (N_943,N_38,N_478);
nor U944 (N_944,N_99,N_313);
xnor U945 (N_945,N_421,N_269);
nor U946 (N_946,N_479,N_211);
and U947 (N_947,N_374,N_455);
and U948 (N_948,N_266,N_127);
nor U949 (N_949,N_279,N_487);
or U950 (N_950,N_70,N_258);
nand U951 (N_951,N_379,N_487);
xor U952 (N_952,N_1,N_364);
xor U953 (N_953,N_56,N_210);
or U954 (N_954,N_204,N_351);
nor U955 (N_955,N_332,N_401);
nor U956 (N_956,N_140,N_394);
or U957 (N_957,N_180,N_264);
or U958 (N_958,N_478,N_387);
nor U959 (N_959,N_302,N_234);
xnor U960 (N_960,N_249,N_173);
or U961 (N_961,N_347,N_200);
nor U962 (N_962,N_188,N_426);
nor U963 (N_963,N_148,N_32);
nand U964 (N_964,N_316,N_321);
xor U965 (N_965,N_220,N_161);
nand U966 (N_966,N_129,N_176);
xnor U967 (N_967,N_313,N_201);
xnor U968 (N_968,N_38,N_426);
nand U969 (N_969,N_75,N_222);
and U970 (N_970,N_274,N_457);
nor U971 (N_971,N_323,N_310);
or U972 (N_972,N_426,N_201);
xor U973 (N_973,N_262,N_251);
and U974 (N_974,N_134,N_392);
nor U975 (N_975,N_110,N_140);
xnor U976 (N_976,N_369,N_275);
nor U977 (N_977,N_329,N_487);
nand U978 (N_978,N_482,N_51);
nand U979 (N_979,N_318,N_43);
or U980 (N_980,N_311,N_253);
nor U981 (N_981,N_224,N_121);
nor U982 (N_982,N_151,N_53);
or U983 (N_983,N_154,N_78);
nor U984 (N_984,N_427,N_241);
xor U985 (N_985,N_193,N_68);
or U986 (N_986,N_260,N_116);
nand U987 (N_987,N_203,N_476);
nor U988 (N_988,N_206,N_46);
nand U989 (N_989,N_254,N_472);
and U990 (N_990,N_307,N_130);
nor U991 (N_991,N_145,N_126);
and U992 (N_992,N_455,N_3);
nor U993 (N_993,N_6,N_273);
or U994 (N_994,N_102,N_149);
or U995 (N_995,N_145,N_419);
and U996 (N_996,N_405,N_379);
or U997 (N_997,N_187,N_260);
nand U998 (N_998,N_136,N_55);
or U999 (N_999,N_359,N_39);
nand U1000 (N_1000,N_878,N_966);
and U1001 (N_1001,N_730,N_663);
nand U1002 (N_1002,N_862,N_547);
nand U1003 (N_1003,N_685,N_614);
or U1004 (N_1004,N_967,N_591);
and U1005 (N_1005,N_721,N_672);
nand U1006 (N_1006,N_965,N_945);
and U1007 (N_1007,N_733,N_812);
nand U1008 (N_1008,N_610,N_856);
nand U1009 (N_1009,N_992,N_932);
or U1010 (N_1010,N_904,N_770);
and U1011 (N_1011,N_736,N_836);
and U1012 (N_1012,N_826,N_930);
or U1013 (N_1013,N_680,N_750);
and U1014 (N_1014,N_594,N_604);
nand U1015 (N_1015,N_529,N_753);
or U1016 (N_1016,N_963,N_863);
xor U1017 (N_1017,N_701,N_549);
or U1018 (N_1018,N_557,N_999);
xnor U1019 (N_1019,N_808,N_751);
xnor U1020 (N_1020,N_734,N_929);
nor U1021 (N_1021,N_789,N_786);
xor U1022 (N_1022,N_596,N_854);
xnor U1023 (N_1023,N_865,N_755);
or U1024 (N_1024,N_859,N_592);
and U1025 (N_1025,N_829,N_510);
or U1026 (N_1026,N_796,N_969);
or U1027 (N_1027,N_879,N_691);
or U1028 (N_1028,N_700,N_864);
nor U1029 (N_1029,N_937,N_565);
xnor U1030 (N_1030,N_985,N_561);
nor U1031 (N_1031,N_542,N_955);
nor U1032 (N_1032,N_778,N_743);
or U1033 (N_1033,N_689,N_928);
and U1034 (N_1034,N_913,N_900);
and U1035 (N_1035,N_538,N_909);
or U1036 (N_1036,N_705,N_961);
xnor U1037 (N_1037,N_880,N_869);
nand U1038 (N_1038,N_813,N_537);
nor U1039 (N_1039,N_754,N_946);
nand U1040 (N_1040,N_749,N_723);
and U1041 (N_1041,N_630,N_681);
or U1042 (N_1042,N_884,N_760);
nand U1043 (N_1043,N_853,N_772);
or U1044 (N_1044,N_833,N_820);
or U1045 (N_1045,N_556,N_533);
nand U1046 (N_1046,N_620,N_827);
nor U1047 (N_1047,N_883,N_745);
or U1048 (N_1048,N_534,N_922);
or U1049 (N_1049,N_997,N_634);
and U1050 (N_1050,N_741,N_803);
and U1051 (N_1051,N_668,N_500);
nor U1052 (N_1052,N_839,N_819);
nor U1053 (N_1053,N_939,N_566);
nand U1054 (N_1054,N_782,N_677);
nor U1055 (N_1055,N_920,N_524);
nor U1056 (N_1056,N_779,N_886);
or U1057 (N_1057,N_590,N_970);
nor U1058 (N_1058,N_896,N_666);
nor U1059 (N_1059,N_818,N_765);
nand U1060 (N_1060,N_665,N_676);
and U1061 (N_1061,N_673,N_553);
or U1062 (N_1062,N_872,N_956);
or U1063 (N_1063,N_866,N_960);
or U1064 (N_1064,N_692,N_647);
nand U1065 (N_1065,N_981,N_622);
and U1066 (N_1066,N_984,N_943);
or U1067 (N_1067,N_605,N_842);
nor U1068 (N_1068,N_719,N_684);
and U1069 (N_1069,N_639,N_588);
nand U1070 (N_1070,N_558,N_987);
xor U1071 (N_1071,N_693,N_756);
and U1072 (N_1072,N_846,N_546);
or U1073 (N_1073,N_821,N_570);
and U1074 (N_1074,N_897,N_977);
and U1075 (N_1075,N_964,N_942);
xnor U1076 (N_1076,N_563,N_522);
xnor U1077 (N_1077,N_933,N_916);
and U1078 (N_1078,N_927,N_528);
and U1079 (N_1079,N_514,N_508);
and U1080 (N_1080,N_575,N_517);
xor U1081 (N_1081,N_595,N_906);
nor U1082 (N_1082,N_867,N_735);
xor U1083 (N_1083,N_845,N_602);
and U1084 (N_1084,N_895,N_516);
or U1085 (N_1085,N_651,N_612);
xor U1086 (N_1086,N_994,N_697);
or U1087 (N_1087,N_747,N_674);
nand U1088 (N_1088,N_536,N_850);
or U1089 (N_1089,N_655,N_844);
nor U1090 (N_1090,N_773,N_972);
and U1091 (N_1091,N_870,N_828);
nor U1092 (N_1092,N_601,N_979);
and U1093 (N_1093,N_503,N_882);
and U1094 (N_1094,N_947,N_838);
and U1095 (N_1095,N_752,N_793);
nand U1096 (N_1096,N_824,N_840);
xor U1097 (N_1097,N_924,N_791);
or U1098 (N_1098,N_934,N_968);
xnor U1099 (N_1099,N_617,N_704);
nor U1100 (N_1100,N_706,N_628);
xnor U1101 (N_1101,N_807,N_649);
nand U1102 (N_1102,N_660,N_940);
xnor U1103 (N_1103,N_662,N_573);
or U1104 (N_1104,N_852,N_623);
or U1105 (N_1105,N_720,N_777);
or U1106 (N_1106,N_640,N_848);
or U1107 (N_1107,N_759,N_739);
nand U1108 (N_1108,N_905,N_825);
nand U1109 (N_1109,N_626,N_935);
or U1110 (N_1110,N_902,N_868);
xnor U1111 (N_1111,N_607,N_746);
or U1112 (N_1112,N_768,N_530);
and U1113 (N_1113,N_952,N_722);
nor U1114 (N_1114,N_714,N_599);
nand U1115 (N_1115,N_877,N_763);
and U1116 (N_1116,N_682,N_608);
xnor U1117 (N_1117,N_511,N_797);
and U1118 (N_1118,N_802,N_815);
nor U1119 (N_1119,N_857,N_811);
xor U1120 (N_1120,N_569,N_798);
nand U1121 (N_1121,N_502,N_769);
xnor U1122 (N_1122,N_702,N_512);
nand U1123 (N_1123,N_998,N_919);
xnor U1124 (N_1124,N_914,N_577);
xnor U1125 (N_1125,N_652,N_551);
nand U1126 (N_1126,N_703,N_771);
and U1127 (N_1127,N_788,N_726);
nor U1128 (N_1128,N_944,N_874);
and U1129 (N_1129,N_589,N_548);
nand U1130 (N_1130,N_953,N_941);
and U1131 (N_1131,N_507,N_911);
xnor U1132 (N_1132,N_579,N_995);
xor U1133 (N_1133,N_699,N_891);
and U1134 (N_1134,N_871,N_564);
nand U1135 (N_1135,N_576,N_776);
or U1136 (N_1136,N_535,N_876);
nor U1137 (N_1137,N_690,N_571);
xnor U1138 (N_1138,N_980,N_688);
xnor U1139 (N_1139,N_784,N_523);
nand U1140 (N_1140,N_526,N_731);
or U1141 (N_1141,N_657,N_695);
nand U1142 (N_1142,N_748,N_951);
and U1143 (N_1143,N_629,N_781);
nor U1144 (N_1144,N_983,N_893);
xnor U1145 (N_1145,N_910,N_832);
and U1146 (N_1146,N_949,N_525);
xor U1147 (N_1147,N_948,N_583);
or U1148 (N_1148,N_908,N_975);
nor U1149 (N_1149,N_729,N_986);
and U1150 (N_1150,N_742,N_717);
and U1151 (N_1151,N_901,N_918);
or U1152 (N_1152,N_633,N_584);
nor U1153 (N_1153,N_996,N_899);
and U1154 (N_1154,N_912,N_637);
nor U1155 (N_1155,N_613,N_635);
nor U1156 (N_1156,N_830,N_707);
and U1157 (N_1157,N_925,N_860);
and U1158 (N_1158,N_806,N_923);
nand U1159 (N_1159,N_686,N_774);
and U1160 (N_1160,N_664,N_567);
nand U1161 (N_1161,N_718,N_725);
or U1162 (N_1162,N_667,N_698);
and U1163 (N_1163,N_572,N_598);
xnor U1164 (N_1164,N_683,N_600);
and U1165 (N_1165,N_586,N_671);
nor U1166 (N_1166,N_505,N_545);
and U1167 (N_1167,N_527,N_976);
nand U1168 (N_1168,N_531,N_974);
nand U1169 (N_1169,N_767,N_632);
nor U1170 (N_1170,N_696,N_792);
and U1171 (N_1171,N_959,N_890);
nand U1172 (N_1172,N_520,N_659);
or U1173 (N_1173,N_518,N_513);
nor U1174 (N_1174,N_585,N_645);
and U1175 (N_1175,N_950,N_991);
or U1176 (N_1176,N_638,N_888);
or U1177 (N_1177,N_715,N_809);
nor U1178 (N_1178,N_728,N_843);
xnor U1179 (N_1179,N_606,N_780);
nor U1180 (N_1180,N_732,N_519);
nand U1181 (N_1181,N_917,N_938);
nand U1182 (N_1182,N_823,N_708);
nand U1183 (N_1183,N_541,N_989);
nor U1184 (N_1184,N_744,N_587);
nand U1185 (N_1185,N_795,N_624);
nor U1186 (N_1186,N_501,N_615);
or U1187 (N_1187,N_737,N_835);
and U1188 (N_1188,N_988,N_609);
nor U1189 (N_1189,N_855,N_555);
and U1190 (N_1190,N_661,N_885);
nor U1191 (N_1191,N_804,N_800);
nor U1192 (N_1192,N_709,N_578);
nand U1193 (N_1193,N_539,N_543);
nand U1194 (N_1194,N_936,N_678);
and U1195 (N_1195,N_921,N_532);
xnor U1196 (N_1196,N_816,N_957);
nand U1197 (N_1197,N_619,N_907);
or U1198 (N_1198,N_650,N_926);
or U1199 (N_1199,N_603,N_506);
or U1200 (N_1200,N_631,N_814);
xor U1201 (N_1201,N_903,N_766);
xnor U1202 (N_1202,N_787,N_711);
nand U1203 (N_1203,N_679,N_646);
nor U1204 (N_1204,N_515,N_568);
nand U1205 (N_1205,N_831,N_962);
nand U1206 (N_1206,N_611,N_574);
xnor U1207 (N_1207,N_581,N_978);
nor U1208 (N_1208,N_616,N_653);
xor U1209 (N_1209,N_849,N_550);
or U1210 (N_1210,N_799,N_582);
and U1211 (N_1211,N_562,N_670);
or U1212 (N_1212,N_873,N_982);
xor U1213 (N_1213,N_712,N_875);
or U1214 (N_1214,N_687,N_509);
nand U1215 (N_1215,N_861,N_834);
nor U1216 (N_1216,N_658,N_654);
nand U1217 (N_1217,N_675,N_847);
xor U1218 (N_1218,N_971,N_817);
or U1219 (N_1219,N_559,N_641);
or U1220 (N_1220,N_990,N_521);
or U1221 (N_1221,N_801,N_757);
nor U1222 (N_1222,N_716,N_764);
nand U1223 (N_1223,N_669,N_694);
or U1224 (N_1224,N_625,N_710);
or U1225 (N_1225,N_898,N_810);
nand U1226 (N_1226,N_627,N_644);
nor U1227 (N_1227,N_822,N_931);
and U1228 (N_1228,N_762,N_790);
nand U1229 (N_1229,N_593,N_552);
or U1230 (N_1230,N_958,N_915);
nand U1231 (N_1231,N_738,N_713);
nor U1232 (N_1232,N_892,N_794);
and U1233 (N_1233,N_805,N_540);
xnor U1234 (N_1234,N_954,N_775);
nand U1235 (N_1235,N_761,N_560);
nand U1236 (N_1236,N_727,N_993);
or U1237 (N_1237,N_785,N_643);
or U1238 (N_1238,N_841,N_973);
nor U1239 (N_1239,N_887,N_724);
and U1240 (N_1240,N_783,N_851);
and U1241 (N_1241,N_881,N_837);
xor U1242 (N_1242,N_621,N_858);
nand U1243 (N_1243,N_648,N_618);
or U1244 (N_1244,N_554,N_597);
and U1245 (N_1245,N_894,N_740);
xor U1246 (N_1246,N_889,N_580);
nor U1247 (N_1247,N_758,N_504);
nor U1248 (N_1248,N_656,N_636);
nor U1249 (N_1249,N_642,N_544);
and U1250 (N_1250,N_804,N_616);
nor U1251 (N_1251,N_722,N_798);
nand U1252 (N_1252,N_672,N_783);
nand U1253 (N_1253,N_544,N_951);
or U1254 (N_1254,N_572,N_927);
xor U1255 (N_1255,N_630,N_608);
xnor U1256 (N_1256,N_568,N_819);
or U1257 (N_1257,N_509,N_943);
and U1258 (N_1258,N_845,N_673);
xnor U1259 (N_1259,N_809,N_672);
or U1260 (N_1260,N_851,N_582);
and U1261 (N_1261,N_948,N_503);
xor U1262 (N_1262,N_739,N_721);
and U1263 (N_1263,N_724,N_706);
xor U1264 (N_1264,N_687,N_580);
nand U1265 (N_1265,N_754,N_967);
xnor U1266 (N_1266,N_966,N_673);
and U1267 (N_1267,N_912,N_533);
and U1268 (N_1268,N_824,N_979);
nand U1269 (N_1269,N_789,N_960);
nand U1270 (N_1270,N_723,N_939);
nand U1271 (N_1271,N_890,N_908);
and U1272 (N_1272,N_920,N_725);
nand U1273 (N_1273,N_886,N_500);
or U1274 (N_1274,N_576,N_970);
xnor U1275 (N_1275,N_762,N_810);
or U1276 (N_1276,N_611,N_704);
xnor U1277 (N_1277,N_886,N_923);
nor U1278 (N_1278,N_873,N_664);
xor U1279 (N_1279,N_805,N_806);
or U1280 (N_1280,N_684,N_988);
nand U1281 (N_1281,N_704,N_942);
xnor U1282 (N_1282,N_931,N_833);
nand U1283 (N_1283,N_925,N_565);
nand U1284 (N_1284,N_842,N_922);
xnor U1285 (N_1285,N_928,N_696);
nor U1286 (N_1286,N_783,N_933);
nor U1287 (N_1287,N_937,N_876);
and U1288 (N_1288,N_793,N_514);
xnor U1289 (N_1289,N_837,N_882);
nor U1290 (N_1290,N_696,N_694);
nand U1291 (N_1291,N_555,N_520);
xnor U1292 (N_1292,N_899,N_685);
xor U1293 (N_1293,N_912,N_502);
xnor U1294 (N_1294,N_609,N_830);
xnor U1295 (N_1295,N_657,N_608);
nand U1296 (N_1296,N_506,N_625);
xor U1297 (N_1297,N_865,N_946);
nand U1298 (N_1298,N_980,N_841);
nor U1299 (N_1299,N_803,N_816);
or U1300 (N_1300,N_933,N_740);
nor U1301 (N_1301,N_749,N_930);
nand U1302 (N_1302,N_690,N_937);
or U1303 (N_1303,N_724,N_691);
and U1304 (N_1304,N_936,N_722);
or U1305 (N_1305,N_844,N_821);
xnor U1306 (N_1306,N_729,N_797);
xor U1307 (N_1307,N_947,N_725);
nor U1308 (N_1308,N_909,N_984);
xnor U1309 (N_1309,N_807,N_836);
nand U1310 (N_1310,N_805,N_986);
xor U1311 (N_1311,N_826,N_848);
nand U1312 (N_1312,N_812,N_522);
xor U1313 (N_1313,N_551,N_843);
nor U1314 (N_1314,N_882,N_892);
nor U1315 (N_1315,N_939,N_724);
or U1316 (N_1316,N_779,N_984);
or U1317 (N_1317,N_967,N_574);
or U1318 (N_1318,N_567,N_599);
or U1319 (N_1319,N_613,N_738);
nand U1320 (N_1320,N_607,N_851);
xor U1321 (N_1321,N_817,N_663);
nand U1322 (N_1322,N_751,N_753);
xnor U1323 (N_1323,N_737,N_568);
nand U1324 (N_1324,N_819,N_776);
and U1325 (N_1325,N_976,N_922);
nor U1326 (N_1326,N_846,N_701);
and U1327 (N_1327,N_822,N_780);
and U1328 (N_1328,N_595,N_775);
and U1329 (N_1329,N_525,N_793);
nor U1330 (N_1330,N_977,N_952);
nor U1331 (N_1331,N_543,N_576);
nand U1332 (N_1332,N_653,N_623);
or U1333 (N_1333,N_667,N_786);
xor U1334 (N_1334,N_516,N_812);
and U1335 (N_1335,N_824,N_944);
nand U1336 (N_1336,N_948,N_684);
nand U1337 (N_1337,N_997,N_826);
xor U1338 (N_1338,N_824,N_956);
and U1339 (N_1339,N_864,N_788);
xor U1340 (N_1340,N_671,N_690);
nor U1341 (N_1341,N_926,N_974);
xnor U1342 (N_1342,N_765,N_825);
xnor U1343 (N_1343,N_547,N_916);
xor U1344 (N_1344,N_807,N_934);
and U1345 (N_1345,N_783,N_652);
nand U1346 (N_1346,N_875,N_955);
nand U1347 (N_1347,N_696,N_655);
nand U1348 (N_1348,N_841,N_750);
nand U1349 (N_1349,N_747,N_621);
xnor U1350 (N_1350,N_937,N_786);
or U1351 (N_1351,N_649,N_669);
xnor U1352 (N_1352,N_867,N_781);
xor U1353 (N_1353,N_619,N_920);
xnor U1354 (N_1354,N_566,N_724);
xor U1355 (N_1355,N_930,N_745);
and U1356 (N_1356,N_501,N_519);
and U1357 (N_1357,N_858,N_955);
nand U1358 (N_1358,N_963,N_628);
and U1359 (N_1359,N_680,N_656);
or U1360 (N_1360,N_726,N_903);
or U1361 (N_1361,N_680,N_513);
nor U1362 (N_1362,N_545,N_623);
and U1363 (N_1363,N_698,N_838);
or U1364 (N_1364,N_865,N_723);
or U1365 (N_1365,N_859,N_866);
and U1366 (N_1366,N_753,N_549);
xnor U1367 (N_1367,N_927,N_523);
and U1368 (N_1368,N_932,N_720);
nor U1369 (N_1369,N_529,N_646);
or U1370 (N_1370,N_516,N_761);
xor U1371 (N_1371,N_921,N_637);
and U1372 (N_1372,N_934,N_734);
nor U1373 (N_1373,N_725,N_997);
nor U1374 (N_1374,N_508,N_933);
nor U1375 (N_1375,N_907,N_775);
and U1376 (N_1376,N_596,N_796);
nor U1377 (N_1377,N_592,N_565);
and U1378 (N_1378,N_876,N_860);
and U1379 (N_1379,N_800,N_541);
xnor U1380 (N_1380,N_530,N_504);
and U1381 (N_1381,N_974,N_902);
xnor U1382 (N_1382,N_905,N_694);
and U1383 (N_1383,N_513,N_759);
and U1384 (N_1384,N_959,N_648);
nand U1385 (N_1385,N_653,N_586);
or U1386 (N_1386,N_819,N_756);
nor U1387 (N_1387,N_607,N_569);
and U1388 (N_1388,N_759,N_686);
and U1389 (N_1389,N_904,N_987);
nand U1390 (N_1390,N_868,N_715);
or U1391 (N_1391,N_981,N_751);
nor U1392 (N_1392,N_954,N_725);
nand U1393 (N_1393,N_887,N_749);
nand U1394 (N_1394,N_696,N_861);
nand U1395 (N_1395,N_589,N_595);
xor U1396 (N_1396,N_833,N_616);
nor U1397 (N_1397,N_722,N_647);
xor U1398 (N_1398,N_503,N_913);
xnor U1399 (N_1399,N_753,N_722);
nand U1400 (N_1400,N_796,N_570);
or U1401 (N_1401,N_815,N_503);
nand U1402 (N_1402,N_872,N_697);
nor U1403 (N_1403,N_676,N_958);
xor U1404 (N_1404,N_837,N_853);
nor U1405 (N_1405,N_990,N_980);
or U1406 (N_1406,N_806,N_672);
nand U1407 (N_1407,N_789,N_536);
nor U1408 (N_1408,N_979,N_511);
or U1409 (N_1409,N_546,N_703);
and U1410 (N_1410,N_844,N_836);
nor U1411 (N_1411,N_708,N_807);
or U1412 (N_1412,N_541,N_834);
and U1413 (N_1413,N_868,N_666);
nand U1414 (N_1414,N_657,N_765);
nor U1415 (N_1415,N_963,N_793);
and U1416 (N_1416,N_597,N_948);
xnor U1417 (N_1417,N_602,N_892);
nand U1418 (N_1418,N_863,N_954);
xor U1419 (N_1419,N_651,N_810);
or U1420 (N_1420,N_506,N_716);
nand U1421 (N_1421,N_561,N_874);
xor U1422 (N_1422,N_756,N_924);
and U1423 (N_1423,N_874,N_881);
xor U1424 (N_1424,N_744,N_556);
or U1425 (N_1425,N_840,N_573);
nor U1426 (N_1426,N_619,N_736);
or U1427 (N_1427,N_507,N_908);
xor U1428 (N_1428,N_772,N_945);
nor U1429 (N_1429,N_719,N_660);
or U1430 (N_1430,N_757,N_715);
nor U1431 (N_1431,N_672,N_514);
xor U1432 (N_1432,N_579,N_622);
or U1433 (N_1433,N_700,N_886);
nand U1434 (N_1434,N_854,N_939);
xor U1435 (N_1435,N_714,N_911);
and U1436 (N_1436,N_747,N_791);
and U1437 (N_1437,N_897,N_523);
or U1438 (N_1438,N_665,N_510);
and U1439 (N_1439,N_959,N_920);
and U1440 (N_1440,N_900,N_677);
nand U1441 (N_1441,N_793,N_857);
and U1442 (N_1442,N_571,N_930);
or U1443 (N_1443,N_813,N_774);
and U1444 (N_1444,N_951,N_813);
nor U1445 (N_1445,N_722,N_585);
nor U1446 (N_1446,N_787,N_656);
or U1447 (N_1447,N_551,N_849);
or U1448 (N_1448,N_633,N_891);
nor U1449 (N_1449,N_864,N_745);
or U1450 (N_1450,N_962,N_615);
and U1451 (N_1451,N_815,N_871);
nand U1452 (N_1452,N_727,N_745);
or U1453 (N_1453,N_947,N_877);
and U1454 (N_1454,N_622,N_949);
or U1455 (N_1455,N_667,N_948);
nor U1456 (N_1456,N_925,N_510);
and U1457 (N_1457,N_514,N_668);
nand U1458 (N_1458,N_762,N_713);
nor U1459 (N_1459,N_777,N_578);
and U1460 (N_1460,N_671,N_987);
nor U1461 (N_1461,N_555,N_950);
and U1462 (N_1462,N_700,N_914);
nand U1463 (N_1463,N_599,N_886);
xnor U1464 (N_1464,N_813,N_924);
or U1465 (N_1465,N_794,N_923);
nand U1466 (N_1466,N_868,N_712);
nand U1467 (N_1467,N_663,N_969);
xor U1468 (N_1468,N_881,N_563);
or U1469 (N_1469,N_671,N_545);
xor U1470 (N_1470,N_803,N_937);
nor U1471 (N_1471,N_648,N_779);
and U1472 (N_1472,N_605,N_506);
nor U1473 (N_1473,N_747,N_848);
and U1474 (N_1474,N_963,N_612);
and U1475 (N_1475,N_585,N_991);
and U1476 (N_1476,N_609,N_528);
or U1477 (N_1477,N_724,N_596);
nor U1478 (N_1478,N_680,N_557);
xnor U1479 (N_1479,N_820,N_598);
nor U1480 (N_1480,N_899,N_508);
and U1481 (N_1481,N_576,N_765);
nor U1482 (N_1482,N_800,N_803);
nor U1483 (N_1483,N_600,N_672);
nor U1484 (N_1484,N_977,N_712);
nand U1485 (N_1485,N_852,N_821);
xor U1486 (N_1486,N_924,N_836);
or U1487 (N_1487,N_742,N_515);
xor U1488 (N_1488,N_962,N_516);
and U1489 (N_1489,N_726,N_597);
and U1490 (N_1490,N_762,N_879);
xnor U1491 (N_1491,N_794,N_983);
and U1492 (N_1492,N_946,N_910);
or U1493 (N_1493,N_615,N_564);
and U1494 (N_1494,N_526,N_789);
and U1495 (N_1495,N_585,N_621);
xnor U1496 (N_1496,N_529,N_643);
xor U1497 (N_1497,N_645,N_633);
nor U1498 (N_1498,N_932,N_746);
and U1499 (N_1499,N_558,N_978);
and U1500 (N_1500,N_1149,N_1339);
xnor U1501 (N_1501,N_1383,N_1487);
nand U1502 (N_1502,N_1307,N_1076);
nand U1503 (N_1503,N_1277,N_1156);
or U1504 (N_1504,N_1112,N_1090);
nand U1505 (N_1505,N_1394,N_1347);
or U1506 (N_1506,N_1180,N_1051);
nand U1507 (N_1507,N_1334,N_1077);
nor U1508 (N_1508,N_1260,N_1226);
and U1509 (N_1509,N_1411,N_1315);
or U1510 (N_1510,N_1061,N_1492);
nor U1511 (N_1511,N_1225,N_1374);
nor U1512 (N_1512,N_1187,N_1441);
and U1513 (N_1513,N_1044,N_1355);
xor U1514 (N_1514,N_1367,N_1106);
and U1515 (N_1515,N_1251,N_1464);
and U1516 (N_1516,N_1167,N_1333);
nand U1517 (N_1517,N_1344,N_1454);
xnor U1518 (N_1518,N_1119,N_1489);
xnor U1519 (N_1519,N_1381,N_1165);
xnor U1520 (N_1520,N_1089,N_1181);
and U1521 (N_1521,N_1499,N_1498);
xnor U1522 (N_1522,N_1214,N_1393);
nor U1523 (N_1523,N_1128,N_1306);
nand U1524 (N_1524,N_1031,N_1436);
nand U1525 (N_1525,N_1444,N_1254);
xnor U1526 (N_1526,N_1194,N_1324);
and U1527 (N_1527,N_1271,N_1137);
and U1528 (N_1528,N_1170,N_1234);
and U1529 (N_1529,N_1257,N_1134);
and U1530 (N_1530,N_1327,N_1286);
xnor U1531 (N_1531,N_1276,N_1215);
and U1532 (N_1532,N_1268,N_1365);
nor U1533 (N_1533,N_1026,N_1266);
or U1534 (N_1534,N_1084,N_1033);
or U1535 (N_1535,N_1080,N_1486);
and U1536 (N_1536,N_1375,N_1272);
and U1537 (N_1537,N_1122,N_1485);
nor U1538 (N_1538,N_1058,N_1224);
nor U1539 (N_1539,N_1159,N_1100);
and U1540 (N_1540,N_1046,N_1064);
xnor U1541 (N_1541,N_1358,N_1263);
and U1542 (N_1542,N_1107,N_1133);
nor U1543 (N_1543,N_1113,N_1458);
xor U1544 (N_1544,N_1497,N_1346);
nand U1545 (N_1545,N_1014,N_1050);
or U1546 (N_1546,N_1378,N_1190);
and U1547 (N_1547,N_1377,N_1099);
xnor U1548 (N_1548,N_1020,N_1171);
nor U1549 (N_1549,N_1348,N_1188);
xnor U1550 (N_1550,N_1140,N_1148);
xor U1551 (N_1551,N_1261,N_1239);
nand U1552 (N_1552,N_1379,N_1125);
xor U1553 (N_1553,N_1005,N_1430);
or U1554 (N_1554,N_1070,N_1437);
or U1555 (N_1555,N_1396,N_1311);
or U1556 (N_1556,N_1059,N_1053);
nor U1557 (N_1557,N_1338,N_1491);
nand U1558 (N_1558,N_1252,N_1083);
nor U1559 (N_1559,N_1245,N_1230);
nand U1560 (N_1560,N_1326,N_1183);
nor U1561 (N_1561,N_1494,N_1223);
xnor U1562 (N_1562,N_1075,N_1270);
or U1563 (N_1563,N_1309,N_1004);
and U1564 (N_1564,N_1398,N_1343);
nor U1565 (N_1565,N_1293,N_1189);
nor U1566 (N_1566,N_1399,N_1273);
nor U1567 (N_1567,N_1483,N_1172);
xnor U1568 (N_1568,N_1397,N_1364);
or U1569 (N_1569,N_1191,N_1493);
xnor U1570 (N_1570,N_1087,N_1395);
xnor U1571 (N_1571,N_1067,N_1414);
nand U1572 (N_1572,N_1422,N_1211);
or U1573 (N_1573,N_1184,N_1221);
xor U1574 (N_1574,N_1142,N_1136);
and U1575 (N_1575,N_1299,N_1431);
nand U1576 (N_1576,N_1015,N_1417);
or U1577 (N_1577,N_1298,N_1305);
nor U1578 (N_1578,N_1030,N_1316);
xnor U1579 (N_1579,N_1247,N_1423);
or U1580 (N_1580,N_1328,N_1478);
nor U1581 (N_1581,N_1297,N_1095);
nor U1582 (N_1582,N_1363,N_1463);
nand U1583 (N_1583,N_1108,N_1448);
or U1584 (N_1584,N_1407,N_1176);
nor U1585 (N_1585,N_1175,N_1490);
or U1586 (N_1586,N_1009,N_1420);
nor U1587 (N_1587,N_1475,N_1290);
and U1588 (N_1588,N_1057,N_1291);
nor U1589 (N_1589,N_1238,N_1314);
nor U1590 (N_1590,N_1488,N_1373);
nand U1591 (N_1591,N_1025,N_1256);
xor U1592 (N_1592,N_1163,N_1473);
or U1593 (N_1593,N_1129,N_1403);
nor U1594 (N_1594,N_1081,N_1289);
nor U1595 (N_1595,N_1071,N_1242);
or U1596 (N_1596,N_1021,N_1474);
nor U1597 (N_1597,N_1233,N_1438);
nor U1598 (N_1598,N_1138,N_1069);
xnor U1599 (N_1599,N_1432,N_1453);
nand U1600 (N_1600,N_1250,N_1278);
and U1601 (N_1601,N_1151,N_1001);
nand U1602 (N_1602,N_1130,N_1351);
xor U1603 (N_1603,N_1386,N_1088);
nand U1604 (N_1604,N_1246,N_1296);
nor U1605 (N_1605,N_1390,N_1016);
xnor U1606 (N_1606,N_1078,N_1178);
nor U1607 (N_1607,N_1323,N_1472);
nor U1608 (N_1608,N_1310,N_1409);
nand U1609 (N_1609,N_1185,N_1460);
or U1610 (N_1610,N_1353,N_1337);
nor U1611 (N_1611,N_1451,N_1048);
nand U1612 (N_1612,N_1421,N_1283);
or U1613 (N_1613,N_1433,N_1418);
and U1614 (N_1614,N_1274,N_1264);
xor U1615 (N_1615,N_1415,N_1120);
nor U1616 (N_1616,N_1287,N_1153);
xor U1617 (N_1617,N_1166,N_1376);
nand U1618 (N_1618,N_1425,N_1303);
nand U1619 (N_1619,N_1332,N_1229);
nand U1620 (N_1620,N_1484,N_1204);
nor U1621 (N_1621,N_1068,N_1209);
nand U1622 (N_1622,N_1457,N_1102);
or U1623 (N_1623,N_1162,N_1199);
xor U1624 (N_1624,N_1037,N_1336);
xor U1625 (N_1625,N_1392,N_1135);
nor U1626 (N_1626,N_1419,N_1198);
xnor U1627 (N_1627,N_1219,N_1359);
nor U1628 (N_1628,N_1013,N_1321);
or U1629 (N_1629,N_1258,N_1222);
nor U1630 (N_1630,N_1007,N_1391);
nand U1631 (N_1631,N_1110,N_1426);
and U1632 (N_1632,N_1470,N_1002);
and U1633 (N_1633,N_1357,N_1207);
or U1634 (N_1634,N_1062,N_1146);
and U1635 (N_1635,N_1341,N_1202);
nand U1636 (N_1636,N_1210,N_1086);
nor U1637 (N_1637,N_1118,N_1308);
or U1638 (N_1638,N_1302,N_1294);
nor U1639 (N_1639,N_1335,N_1139);
and U1640 (N_1640,N_1479,N_1143);
nor U1641 (N_1641,N_1065,N_1220);
nand U1642 (N_1642,N_1388,N_1072);
or U1643 (N_1643,N_1228,N_1406);
nor U1644 (N_1644,N_1168,N_1400);
or U1645 (N_1645,N_1248,N_1408);
or U1646 (N_1646,N_1253,N_1012);
nor U1647 (N_1647,N_1141,N_1144);
xor U1648 (N_1648,N_1208,N_1213);
nor U1649 (N_1649,N_1269,N_1466);
xor U1650 (N_1650,N_1173,N_1132);
and U1651 (N_1651,N_1201,N_1446);
nand U1652 (N_1652,N_1301,N_1495);
xnor U1653 (N_1653,N_1360,N_1255);
nand U1654 (N_1654,N_1029,N_1197);
nand U1655 (N_1655,N_1467,N_1465);
xor U1656 (N_1656,N_1186,N_1103);
nand U1657 (N_1657,N_1325,N_1340);
nor U1658 (N_1658,N_1232,N_1055);
nor U1659 (N_1659,N_1227,N_1456);
and U1660 (N_1660,N_1054,N_1434);
and U1661 (N_1661,N_1249,N_1114);
and U1662 (N_1662,N_1182,N_1352);
xor U1663 (N_1663,N_1035,N_1109);
xnor U1664 (N_1664,N_1206,N_1104);
and U1665 (N_1665,N_1174,N_1385);
nor U1666 (N_1666,N_1350,N_1123);
xnor U1667 (N_1667,N_1482,N_1349);
nor U1668 (N_1668,N_1449,N_1006);
and U1669 (N_1669,N_1096,N_1387);
nor U1670 (N_1670,N_1049,N_1041);
nand U1671 (N_1671,N_1017,N_1022);
xnor U1672 (N_1672,N_1203,N_1366);
nor U1673 (N_1673,N_1237,N_1282);
or U1674 (N_1674,N_1469,N_1371);
xor U1675 (N_1675,N_1292,N_1085);
nand U1676 (N_1676,N_1461,N_1439);
or U1677 (N_1677,N_1200,N_1342);
or U1678 (N_1678,N_1477,N_1193);
or U1679 (N_1679,N_1169,N_1265);
nand U1680 (N_1680,N_1295,N_1042);
and U1681 (N_1681,N_1101,N_1401);
nand U1682 (N_1682,N_1313,N_1145);
xor U1683 (N_1683,N_1427,N_1056);
or U1684 (N_1684,N_1079,N_1369);
or U1685 (N_1685,N_1244,N_1428);
nand U1686 (N_1686,N_1063,N_1018);
xor U1687 (N_1687,N_1218,N_1300);
nand U1688 (N_1688,N_1445,N_1157);
nand U1689 (N_1689,N_1435,N_1150);
or U1690 (N_1690,N_1196,N_1043);
or U1691 (N_1691,N_1039,N_1032);
nor U1692 (N_1692,N_1126,N_1111);
nand U1693 (N_1693,N_1241,N_1496);
nand U1694 (N_1694,N_1288,N_1161);
or U1695 (N_1695,N_1027,N_1275);
xor U1696 (N_1696,N_1092,N_1082);
nand U1697 (N_1697,N_1382,N_1098);
xor U1698 (N_1698,N_1205,N_1236);
and U1699 (N_1699,N_1179,N_1442);
nand U1700 (N_1700,N_1094,N_1450);
nand U1701 (N_1701,N_1097,N_1052);
nand U1702 (N_1702,N_1121,N_1212);
xor U1703 (N_1703,N_1331,N_1192);
nor U1704 (N_1704,N_1195,N_1003);
and U1705 (N_1705,N_1154,N_1019);
nand U1706 (N_1706,N_1177,N_1047);
nand U1707 (N_1707,N_1317,N_1008);
nand U1708 (N_1708,N_1093,N_1416);
nor U1709 (N_1709,N_1010,N_1424);
or U1710 (N_1710,N_1354,N_1231);
nor U1711 (N_1711,N_1259,N_1024);
and U1712 (N_1712,N_1404,N_1322);
or U1713 (N_1713,N_1262,N_1452);
nor U1714 (N_1714,N_1356,N_1160);
nand U1715 (N_1715,N_1023,N_1040);
xnor U1716 (N_1716,N_1370,N_1124);
or U1717 (N_1717,N_1284,N_1455);
nor U1718 (N_1718,N_1028,N_1280);
xor U1719 (N_1719,N_1116,N_1152);
xnor U1720 (N_1720,N_1476,N_1060);
nor U1721 (N_1721,N_1368,N_1362);
nand U1722 (N_1722,N_1380,N_1320);
and U1723 (N_1723,N_1147,N_1127);
xor U1724 (N_1724,N_1345,N_1279);
nor U1725 (N_1725,N_1412,N_1447);
nor U1726 (N_1726,N_1243,N_1410);
and U1727 (N_1727,N_1240,N_1131);
nand U1728 (N_1728,N_1115,N_1384);
nand U1729 (N_1729,N_1036,N_1105);
nand U1730 (N_1730,N_1471,N_1405);
and U1731 (N_1731,N_1235,N_1480);
xnor U1732 (N_1732,N_1312,N_1329);
nand U1733 (N_1733,N_1117,N_1281);
or U1734 (N_1734,N_1440,N_1330);
and U1735 (N_1735,N_1318,N_1217);
nor U1736 (N_1736,N_1155,N_1304);
and U1737 (N_1737,N_1164,N_1011);
xor U1738 (N_1738,N_1267,N_1389);
or U1739 (N_1739,N_1216,N_1462);
xnor U1740 (N_1740,N_1038,N_1413);
and U1741 (N_1741,N_1066,N_1073);
and U1742 (N_1742,N_1034,N_1372);
xnor U1743 (N_1743,N_1091,N_1429);
nor U1744 (N_1744,N_1158,N_1481);
nand U1745 (N_1745,N_1361,N_1045);
or U1746 (N_1746,N_1459,N_1000);
or U1747 (N_1747,N_1468,N_1285);
xnor U1748 (N_1748,N_1319,N_1074);
nor U1749 (N_1749,N_1443,N_1402);
or U1750 (N_1750,N_1222,N_1221);
xor U1751 (N_1751,N_1365,N_1112);
nand U1752 (N_1752,N_1499,N_1150);
xnor U1753 (N_1753,N_1229,N_1452);
nor U1754 (N_1754,N_1179,N_1420);
nand U1755 (N_1755,N_1234,N_1380);
nand U1756 (N_1756,N_1112,N_1381);
and U1757 (N_1757,N_1215,N_1204);
xnor U1758 (N_1758,N_1373,N_1110);
nor U1759 (N_1759,N_1060,N_1289);
nand U1760 (N_1760,N_1496,N_1068);
xor U1761 (N_1761,N_1253,N_1305);
and U1762 (N_1762,N_1332,N_1392);
and U1763 (N_1763,N_1004,N_1017);
xnor U1764 (N_1764,N_1243,N_1140);
xnor U1765 (N_1765,N_1190,N_1477);
nor U1766 (N_1766,N_1399,N_1290);
and U1767 (N_1767,N_1290,N_1478);
nor U1768 (N_1768,N_1166,N_1448);
nand U1769 (N_1769,N_1348,N_1302);
nand U1770 (N_1770,N_1084,N_1011);
nor U1771 (N_1771,N_1443,N_1002);
nor U1772 (N_1772,N_1182,N_1141);
xor U1773 (N_1773,N_1386,N_1368);
nor U1774 (N_1774,N_1310,N_1391);
nand U1775 (N_1775,N_1135,N_1279);
nor U1776 (N_1776,N_1468,N_1381);
nor U1777 (N_1777,N_1309,N_1496);
nor U1778 (N_1778,N_1016,N_1287);
xor U1779 (N_1779,N_1282,N_1178);
and U1780 (N_1780,N_1318,N_1298);
xor U1781 (N_1781,N_1079,N_1171);
or U1782 (N_1782,N_1477,N_1336);
and U1783 (N_1783,N_1161,N_1265);
or U1784 (N_1784,N_1345,N_1291);
nor U1785 (N_1785,N_1415,N_1329);
xor U1786 (N_1786,N_1383,N_1351);
nand U1787 (N_1787,N_1018,N_1014);
and U1788 (N_1788,N_1280,N_1053);
and U1789 (N_1789,N_1487,N_1227);
and U1790 (N_1790,N_1456,N_1400);
nand U1791 (N_1791,N_1216,N_1033);
or U1792 (N_1792,N_1103,N_1086);
or U1793 (N_1793,N_1157,N_1012);
and U1794 (N_1794,N_1381,N_1122);
nand U1795 (N_1795,N_1313,N_1380);
nor U1796 (N_1796,N_1003,N_1165);
nor U1797 (N_1797,N_1445,N_1103);
and U1798 (N_1798,N_1467,N_1399);
and U1799 (N_1799,N_1239,N_1106);
xor U1800 (N_1800,N_1360,N_1158);
or U1801 (N_1801,N_1255,N_1127);
and U1802 (N_1802,N_1467,N_1127);
xor U1803 (N_1803,N_1176,N_1100);
nand U1804 (N_1804,N_1341,N_1472);
nor U1805 (N_1805,N_1499,N_1492);
and U1806 (N_1806,N_1040,N_1045);
nor U1807 (N_1807,N_1348,N_1360);
nand U1808 (N_1808,N_1376,N_1312);
xor U1809 (N_1809,N_1310,N_1447);
nor U1810 (N_1810,N_1278,N_1358);
and U1811 (N_1811,N_1339,N_1428);
nand U1812 (N_1812,N_1265,N_1423);
nor U1813 (N_1813,N_1205,N_1478);
and U1814 (N_1814,N_1062,N_1163);
nand U1815 (N_1815,N_1265,N_1216);
or U1816 (N_1816,N_1295,N_1071);
and U1817 (N_1817,N_1216,N_1139);
nand U1818 (N_1818,N_1338,N_1046);
nand U1819 (N_1819,N_1115,N_1294);
xor U1820 (N_1820,N_1434,N_1487);
nand U1821 (N_1821,N_1012,N_1410);
xnor U1822 (N_1822,N_1339,N_1451);
nand U1823 (N_1823,N_1038,N_1190);
nor U1824 (N_1824,N_1311,N_1093);
xnor U1825 (N_1825,N_1477,N_1025);
and U1826 (N_1826,N_1351,N_1151);
or U1827 (N_1827,N_1464,N_1326);
nand U1828 (N_1828,N_1328,N_1297);
nor U1829 (N_1829,N_1396,N_1060);
xnor U1830 (N_1830,N_1419,N_1193);
nand U1831 (N_1831,N_1313,N_1457);
xnor U1832 (N_1832,N_1348,N_1308);
and U1833 (N_1833,N_1083,N_1317);
nand U1834 (N_1834,N_1476,N_1113);
nand U1835 (N_1835,N_1429,N_1406);
nor U1836 (N_1836,N_1318,N_1090);
nand U1837 (N_1837,N_1280,N_1244);
or U1838 (N_1838,N_1282,N_1002);
nand U1839 (N_1839,N_1209,N_1336);
xor U1840 (N_1840,N_1073,N_1115);
and U1841 (N_1841,N_1185,N_1416);
or U1842 (N_1842,N_1135,N_1463);
xnor U1843 (N_1843,N_1043,N_1200);
xor U1844 (N_1844,N_1332,N_1246);
or U1845 (N_1845,N_1449,N_1430);
nand U1846 (N_1846,N_1073,N_1175);
nand U1847 (N_1847,N_1050,N_1343);
xnor U1848 (N_1848,N_1182,N_1409);
or U1849 (N_1849,N_1110,N_1291);
xnor U1850 (N_1850,N_1031,N_1411);
nor U1851 (N_1851,N_1282,N_1351);
or U1852 (N_1852,N_1434,N_1485);
nand U1853 (N_1853,N_1482,N_1403);
or U1854 (N_1854,N_1379,N_1196);
nand U1855 (N_1855,N_1138,N_1217);
nand U1856 (N_1856,N_1342,N_1432);
and U1857 (N_1857,N_1396,N_1271);
and U1858 (N_1858,N_1414,N_1039);
or U1859 (N_1859,N_1115,N_1227);
xor U1860 (N_1860,N_1442,N_1084);
and U1861 (N_1861,N_1107,N_1181);
xor U1862 (N_1862,N_1072,N_1212);
nor U1863 (N_1863,N_1000,N_1193);
and U1864 (N_1864,N_1024,N_1318);
nor U1865 (N_1865,N_1239,N_1071);
and U1866 (N_1866,N_1188,N_1431);
and U1867 (N_1867,N_1302,N_1094);
nor U1868 (N_1868,N_1400,N_1126);
xnor U1869 (N_1869,N_1246,N_1247);
nand U1870 (N_1870,N_1430,N_1131);
nor U1871 (N_1871,N_1059,N_1357);
xnor U1872 (N_1872,N_1441,N_1469);
xnor U1873 (N_1873,N_1199,N_1430);
xor U1874 (N_1874,N_1428,N_1063);
and U1875 (N_1875,N_1241,N_1037);
nor U1876 (N_1876,N_1013,N_1077);
xnor U1877 (N_1877,N_1139,N_1440);
and U1878 (N_1878,N_1339,N_1353);
nand U1879 (N_1879,N_1447,N_1123);
or U1880 (N_1880,N_1248,N_1176);
xor U1881 (N_1881,N_1456,N_1022);
xor U1882 (N_1882,N_1279,N_1011);
and U1883 (N_1883,N_1128,N_1160);
nand U1884 (N_1884,N_1390,N_1130);
xor U1885 (N_1885,N_1232,N_1498);
nand U1886 (N_1886,N_1013,N_1111);
nor U1887 (N_1887,N_1177,N_1325);
xor U1888 (N_1888,N_1186,N_1063);
xnor U1889 (N_1889,N_1437,N_1306);
or U1890 (N_1890,N_1350,N_1157);
xor U1891 (N_1891,N_1250,N_1034);
xor U1892 (N_1892,N_1335,N_1494);
and U1893 (N_1893,N_1417,N_1398);
and U1894 (N_1894,N_1198,N_1239);
nor U1895 (N_1895,N_1364,N_1498);
nand U1896 (N_1896,N_1415,N_1361);
or U1897 (N_1897,N_1280,N_1042);
and U1898 (N_1898,N_1431,N_1046);
xor U1899 (N_1899,N_1469,N_1298);
xor U1900 (N_1900,N_1298,N_1248);
and U1901 (N_1901,N_1083,N_1184);
nor U1902 (N_1902,N_1244,N_1257);
nand U1903 (N_1903,N_1339,N_1256);
nand U1904 (N_1904,N_1162,N_1131);
or U1905 (N_1905,N_1037,N_1094);
xor U1906 (N_1906,N_1295,N_1265);
nand U1907 (N_1907,N_1384,N_1162);
nor U1908 (N_1908,N_1069,N_1117);
or U1909 (N_1909,N_1244,N_1145);
and U1910 (N_1910,N_1437,N_1161);
and U1911 (N_1911,N_1153,N_1495);
and U1912 (N_1912,N_1070,N_1489);
or U1913 (N_1913,N_1458,N_1126);
nor U1914 (N_1914,N_1404,N_1293);
and U1915 (N_1915,N_1324,N_1102);
xor U1916 (N_1916,N_1074,N_1195);
xor U1917 (N_1917,N_1067,N_1173);
xor U1918 (N_1918,N_1312,N_1004);
and U1919 (N_1919,N_1290,N_1006);
nor U1920 (N_1920,N_1484,N_1347);
and U1921 (N_1921,N_1488,N_1431);
or U1922 (N_1922,N_1354,N_1485);
nor U1923 (N_1923,N_1338,N_1026);
nor U1924 (N_1924,N_1099,N_1252);
nand U1925 (N_1925,N_1214,N_1428);
and U1926 (N_1926,N_1368,N_1126);
and U1927 (N_1927,N_1086,N_1115);
nor U1928 (N_1928,N_1324,N_1308);
nand U1929 (N_1929,N_1377,N_1216);
nand U1930 (N_1930,N_1486,N_1375);
nor U1931 (N_1931,N_1278,N_1337);
nand U1932 (N_1932,N_1304,N_1377);
or U1933 (N_1933,N_1408,N_1301);
xnor U1934 (N_1934,N_1028,N_1032);
nor U1935 (N_1935,N_1025,N_1050);
or U1936 (N_1936,N_1337,N_1294);
and U1937 (N_1937,N_1451,N_1074);
or U1938 (N_1938,N_1395,N_1122);
and U1939 (N_1939,N_1344,N_1281);
nor U1940 (N_1940,N_1050,N_1172);
and U1941 (N_1941,N_1436,N_1187);
xnor U1942 (N_1942,N_1446,N_1454);
and U1943 (N_1943,N_1224,N_1029);
xnor U1944 (N_1944,N_1289,N_1396);
and U1945 (N_1945,N_1149,N_1252);
and U1946 (N_1946,N_1399,N_1250);
and U1947 (N_1947,N_1469,N_1108);
nor U1948 (N_1948,N_1022,N_1067);
nand U1949 (N_1949,N_1398,N_1256);
or U1950 (N_1950,N_1337,N_1065);
nand U1951 (N_1951,N_1300,N_1049);
nand U1952 (N_1952,N_1307,N_1410);
and U1953 (N_1953,N_1101,N_1189);
xnor U1954 (N_1954,N_1081,N_1111);
and U1955 (N_1955,N_1428,N_1147);
and U1956 (N_1956,N_1117,N_1088);
or U1957 (N_1957,N_1249,N_1062);
or U1958 (N_1958,N_1011,N_1276);
nand U1959 (N_1959,N_1098,N_1426);
or U1960 (N_1960,N_1385,N_1229);
nor U1961 (N_1961,N_1271,N_1100);
and U1962 (N_1962,N_1402,N_1332);
nor U1963 (N_1963,N_1127,N_1058);
nand U1964 (N_1964,N_1315,N_1350);
xor U1965 (N_1965,N_1483,N_1207);
or U1966 (N_1966,N_1268,N_1444);
nor U1967 (N_1967,N_1238,N_1005);
or U1968 (N_1968,N_1348,N_1159);
nor U1969 (N_1969,N_1488,N_1222);
nor U1970 (N_1970,N_1249,N_1166);
or U1971 (N_1971,N_1124,N_1110);
xnor U1972 (N_1972,N_1036,N_1038);
nor U1973 (N_1973,N_1133,N_1289);
nor U1974 (N_1974,N_1211,N_1492);
or U1975 (N_1975,N_1366,N_1015);
xor U1976 (N_1976,N_1028,N_1188);
or U1977 (N_1977,N_1347,N_1396);
xor U1978 (N_1978,N_1244,N_1458);
nand U1979 (N_1979,N_1294,N_1409);
or U1980 (N_1980,N_1061,N_1124);
nand U1981 (N_1981,N_1088,N_1165);
nor U1982 (N_1982,N_1227,N_1378);
xnor U1983 (N_1983,N_1333,N_1369);
and U1984 (N_1984,N_1076,N_1262);
and U1985 (N_1985,N_1175,N_1133);
or U1986 (N_1986,N_1302,N_1126);
nand U1987 (N_1987,N_1023,N_1121);
and U1988 (N_1988,N_1376,N_1468);
xnor U1989 (N_1989,N_1443,N_1263);
nand U1990 (N_1990,N_1316,N_1249);
xor U1991 (N_1991,N_1206,N_1277);
xnor U1992 (N_1992,N_1145,N_1123);
nand U1993 (N_1993,N_1402,N_1478);
and U1994 (N_1994,N_1235,N_1319);
nand U1995 (N_1995,N_1334,N_1115);
or U1996 (N_1996,N_1230,N_1049);
or U1997 (N_1997,N_1362,N_1033);
and U1998 (N_1998,N_1408,N_1270);
and U1999 (N_1999,N_1218,N_1306);
and U2000 (N_2000,N_1750,N_1988);
or U2001 (N_2001,N_1563,N_1534);
or U2002 (N_2002,N_1782,N_1503);
nand U2003 (N_2003,N_1533,N_1821);
xor U2004 (N_2004,N_1759,N_1764);
xor U2005 (N_2005,N_1847,N_1944);
nand U2006 (N_2006,N_1674,N_1939);
or U2007 (N_2007,N_1901,N_1514);
nand U2008 (N_2008,N_1731,N_1937);
and U2009 (N_2009,N_1915,N_1806);
xor U2010 (N_2010,N_1594,N_1729);
or U2011 (N_2011,N_1580,N_1952);
nand U2012 (N_2012,N_1926,N_1522);
nor U2013 (N_2013,N_1592,N_1740);
nand U2014 (N_2014,N_1866,N_1845);
xor U2015 (N_2015,N_1662,N_1531);
nor U2016 (N_2016,N_1921,N_1950);
and U2017 (N_2017,N_1934,N_1798);
or U2018 (N_2018,N_1653,N_1850);
nor U2019 (N_2019,N_1827,N_1936);
xor U2020 (N_2020,N_1669,N_1691);
xor U2021 (N_2021,N_1981,N_1789);
nor U2022 (N_2022,N_1718,N_1949);
nand U2023 (N_2023,N_1642,N_1733);
nand U2024 (N_2024,N_1702,N_1635);
xor U2025 (N_2025,N_1854,N_1908);
nor U2026 (N_2026,N_1838,N_1987);
xnor U2027 (N_2027,N_1896,N_1730);
or U2028 (N_2028,N_1912,N_1743);
or U2029 (N_2029,N_1626,N_1689);
nand U2030 (N_2030,N_1747,N_1556);
and U2031 (N_2031,N_1589,N_1640);
or U2032 (N_2032,N_1562,N_1871);
nand U2033 (N_2033,N_1822,N_1905);
or U2034 (N_2034,N_1787,N_1572);
and U2035 (N_2035,N_1763,N_1931);
and U2036 (N_2036,N_1946,N_1510);
nor U2037 (N_2037,N_1517,N_1852);
nor U2038 (N_2038,N_1754,N_1900);
nand U2039 (N_2039,N_1667,N_1603);
and U2040 (N_2040,N_1551,N_1656);
nand U2041 (N_2041,N_1587,N_1888);
xnor U2042 (N_2042,N_1717,N_1720);
xor U2043 (N_2043,N_1693,N_1612);
and U2044 (N_2044,N_1959,N_1625);
nand U2045 (N_2045,N_1914,N_1542);
and U2046 (N_2046,N_1855,N_1808);
nor U2047 (N_2047,N_1742,N_1723);
nor U2048 (N_2048,N_1790,N_1701);
xor U2049 (N_2049,N_1872,N_1601);
and U2050 (N_2050,N_1766,N_1868);
xnor U2051 (N_2051,N_1825,N_1507);
xor U2052 (N_2052,N_1863,N_1995);
nand U2053 (N_2053,N_1802,N_1602);
nand U2054 (N_2054,N_1728,N_1508);
xnor U2055 (N_2055,N_1620,N_1663);
nor U2056 (N_2056,N_1972,N_1834);
nor U2057 (N_2057,N_1962,N_1608);
and U2058 (N_2058,N_1967,N_1889);
and U2059 (N_2059,N_1828,N_1780);
nor U2060 (N_2060,N_1753,N_1688);
or U2061 (N_2061,N_1752,N_1918);
and U2062 (N_2062,N_1844,N_1862);
nor U2063 (N_2063,N_1772,N_1775);
nor U2064 (N_2064,N_1509,N_1664);
xnor U2065 (N_2065,N_1779,N_1873);
xor U2066 (N_2066,N_1974,N_1957);
or U2067 (N_2067,N_1706,N_1684);
nand U2068 (N_2068,N_1813,N_1577);
and U2069 (N_2069,N_1982,N_1627);
xor U2070 (N_2070,N_1874,N_1857);
and U2071 (N_2071,N_1560,N_1738);
nand U2072 (N_2072,N_1985,N_1805);
xor U2073 (N_2073,N_1800,N_1910);
or U2074 (N_2074,N_1703,N_1557);
xnor U2075 (N_2075,N_1668,N_1619);
or U2076 (N_2076,N_1709,N_1575);
nor U2077 (N_2077,N_1545,N_1628);
xor U2078 (N_2078,N_1833,N_1837);
or U2079 (N_2079,N_1726,N_1561);
nor U2080 (N_2080,N_1812,N_1593);
xor U2081 (N_2081,N_1983,N_1843);
nand U2082 (N_2082,N_1961,N_1724);
and U2083 (N_2083,N_1564,N_1788);
nand U2084 (N_2084,N_1928,N_1932);
nor U2085 (N_2085,N_1708,N_1773);
nor U2086 (N_2086,N_1999,N_1956);
nor U2087 (N_2087,N_1591,N_1906);
nand U2088 (N_2088,N_1783,N_1540);
nand U2089 (N_2089,N_1920,N_1885);
and U2090 (N_2090,N_1978,N_1527);
xnor U2091 (N_2091,N_1538,N_1735);
xor U2092 (N_2092,N_1636,N_1530);
or U2093 (N_2093,N_1511,N_1911);
xor U2094 (N_2094,N_1878,N_1922);
nand U2095 (N_2095,N_1927,N_1760);
and U2096 (N_2096,N_1588,N_1998);
xor U2097 (N_2097,N_1659,N_1795);
nand U2098 (N_2098,N_1810,N_1705);
and U2099 (N_2099,N_1630,N_1604);
or U2100 (N_2100,N_1719,N_1568);
nor U2101 (N_2101,N_1869,N_1548);
or U2102 (N_2102,N_1525,N_1675);
nor U2103 (N_2103,N_1751,N_1553);
and U2104 (N_2104,N_1597,N_1513);
or U2105 (N_2105,N_1794,N_1641);
xor U2106 (N_2106,N_1797,N_1629);
nand U2107 (N_2107,N_1973,N_1887);
xor U2108 (N_2108,N_1519,N_1660);
xor U2109 (N_2109,N_1679,N_1652);
nor U2110 (N_2110,N_1769,N_1815);
xor U2111 (N_2111,N_1930,N_1824);
and U2112 (N_2112,N_1954,N_1935);
xor U2113 (N_2113,N_1964,N_1713);
nor U2114 (N_2114,N_1610,N_1741);
and U2115 (N_2115,N_1744,N_1645);
nor U2116 (N_2116,N_1582,N_1710);
and U2117 (N_2117,N_1622,N_1785);
nor U2118 (N_2118,N_1614,N_1880);
or U2119 (N_2119,N_1638,N_1819);
xor U2120 (N_2120,N_1890,N_1774);
nor U2121 (N_2121,N_1552,N_1940);
or U2122 (N_2122,N_1683,N_1715);
and U2123 (N_2123,N_1765,N_1969);
and U2124 (N_2124,N_1598,N_1992);
xor U2125 (N_2125,N_1811,N_1585);
or U2126 (N_2126,N_1839,N_1586);
xor U2127 (N_2127,N_1929,N_1632);
nand U2128 (N_2128,N_1543,N_1875);
xor U2129 (N_2129,N_1826,N_1616);
and U2130 (N_2130,N_1804,N_1699);
or U2131 (N_2131,N_1680,N_1606);
nor U2132 (N_2132,N_1960,N_1820);
or U2133 (N_2133,N_1655,N_1695);
or U2134 (N_2134,N_1676,N_1681);
or U2135 (N_2135,N_1714,N_1971);
and U2136 (N_2136,N_1725,N_1736);
nand U2137 (N_2137,N_1853,N_1945);
or U2138 (N_2138,N_1646,N_1746);
or U2139 (N_2139,N_1512,N_1879);
or U2140 (N_2140,N_1902,N_1658);
or U2141 (N_2141,N_1696,N_1739);
xnor U2142 (N_2142,N_1623,N_1618);
nor U2143 (N_2143,N_1778,N_1803);
and U2144 (N_2144,N_1768,N_1767);
xnor U2145 (N_2145,N_1786,N_1502);
nor U2146 (N_2146,N_1707,N_1634);
nand U2147 (N_2147,N_1793,N_1516);
nor U2148 (N_2148,N_1566,N_1953);
nand U2149 (N_2149,N_1571,N_1924);
and U2150 (N_2150,N_1732,N_1919);
nor U2151 (N_2151,N_1504,N_1666);
or U2152 (N_2152,N_1980,N_1784);
nor U2153 (N_2153,N_1990,N_1947);
and U2154 (N_2154,N_1958,N_1685);
nor U2155 (N_2155,N_1609,N_1505);
and U2156 (N_2156,N_1637,N_1624);
and U2157 (N_2157,N_1671,N_1762);
or U2158 (N_2158,N_1550,N_1576);
nor U2159 (N_2159,N_1758,N_1756);
and U2160 (N_2160,N_1712,N_1633);
or U2161 (N_2161,N_1734,N_1997);
nor U2162 (N_2162,N_1565,N_1907);
nand U2163 (N_2163,N_1749,N_1864);
or U2164 (N_2164,N_1993,N_1621);
nor U2165 (N_2165,N_1835,N_1840);
nor U2166 (N_2166,N_1916,N_1535);
nor U2167 (N_2167,N_1520,N_1515);
xor U2168 (N_2168,N_1882,N_1590);
or U2169 (N_2169,N_1979,N_1996);
nor U2170 (N_2170,N_1951,N_1831);
or U2171 (N_2171,N_1851,N_1694);
nand U2172 (N_2172,N_1518,N_1941);
and U2173 (N_2173,N_1672,N_1977);
or U2174 (N_2174,N_1745,N_1865);
or U2175 (N_2175,N_1529,N_1617);
nand U2176 (N_2176,N_1599,N_1532);
nor U2177 (N_2177,N_1500,N_1748);
xor U2178 (N_2178,N_1523,N_1673);
and U2179 (N_2179,N_1541,N_1555);
and U2180 (N_2180,N_1611,N_1573);
or U2181 (N_2181,N_1860,N_1737);
and U2182 (N_2182,N_1994,N_1574);
and U2183 (N_2183,N_1700,N_1596);
xor U2184 (N_2184,N_1521,N_1923);
nand U2185 (N_2185,N_1809,N_1917);
or U2186 (N_2186,N_1841,N_1904);
or U2187 (N_2187,N_1581,N_1678);
or U2188 (N_2188,N_1955,N_1942);
nor U2189 (N_2189,N_1881,N_1651);
and U2190 (N_2190,N_1698,N_1607);
or U2191 (N_2191,N_1567,N_1799);
nor U2192 (N_2192,N_1897,N_1661);
nand U2193 (N_2193,N_1781,N_1836);
nor U2194 (N_2194,N_1579,N_1792);
and U2195 (N_2195,N_1842,N_1801);
xnor U2196 (N_2196,N_1870,N_1986);
nor U2197 (N_2197,N_1968,N_1583);
and U2198 (N_2198,N_1975,N_1970);
nand U2199 (N_2199,N_1721,N_1570);
and U2200 (N_2200,N_1816,N_1639);
nor U2201 (N_2201,N_1859,N_1861);
xnor U2202 (N_2202,N_1613,N_1755);
xor U2203 (N_2203,N_1682,N_1559);
nand U2204 (N_2204,N_1849,N_1807);
and U2205 (N_2205,N_1818,N_1697);
xor U2206 (N_2206,N_1963,N_1584);
nand U2207 (N_2207,N_1501,N_1777);
nor U2208 (N_2208,N_1692,N_1791);
nor U2209 (N_2209,N_1578,N_1814);
nand U2210 (N_2210,N_1644,N_1569);
nor U2211 (N_2211,N_1829,N_1686);
xnor U2212 (N_2212,N_1966,N_1544);
nor U2213 (N_2213,N_1605,N_1894);
or U2214 (N_2214,N_1991,N_1933);
nand U2215 (N_2215,N_1537,N_1647);
or U2216 (N_2216,N_1893,N_1976);
xnor U2217 (N_2217,N_1727,N_1711);
or U2218 (N_2218,N_1817,N_1796);
xnor U2219 (N_2219,N_1665,N_1830);
nand U2220 (N_2220,N_1776,N_1846);
nand U2221 (N_2221,N_1650,N_1506);
or U2222 (N_2222,N_1848,N_1899);
nor U2223 (N_2223,N_1867,N_1558);
xnor U2224 (N_2224,N_1895,N_1643);
nor U2225 (N_2225,N_1909,N_1877);
and U2226 (N_2226,N_1943,N_1948);
nand U2227 (N_2227,N_1539,N_1891);
nand U2228 (N_2228,N_1716,N_1761);
nor U2229 (N_2229,N_1823,N_1649);
nand U2230 (N_2230,N_1536,N_1549);
or U2231 (N_2231,N_1595,N_1722);
or U2232 (N_2232,N_1858,N_1757);
nor U2233 (N_2233,N_1600,N_1832);
and U2234 (N_2234,N_1989,N_1615);
xnor U2235 (N_2235,N_1528,N_1856);
nor U2236 (N_2236,N_1892,N_1771);
nor U2237 (N_2237,N_1690,N_1903);
nand U2238 (N_2238,N_1898,N_1704);
xnor U2239 (N_2239,N_1770,N_1657);
nor U2240 (N_2240,N_1876,N_1984);
nor U2241 (N_2241,N_1524,N_1913);
xnor U2242 (N_2242,N_1554,N_1883);
xor U2243 (N_2243,N_1965,N_1687);
nand U2244 (N_2244,N_1546,N_1886);
and U2245 (N_2245,N_1677,N_1631);
nor U2246 (N_2246,N_1670,N_1547);
xor U2247 (N_2247,N_1654,N_1648);
and U2248 (N_2248,N_1925,N_1938);
and U2249 (N_2249,N_1884,N_1526);
nand U2250 (N_2250,N_1630,N_1772);
and U2251 (N_2251,N_1867,N_1895);
and U2252 (N_2252,N_1650,N_1662);
nand U2253 (N_2253,N_1582,N_1617);
nor U2254 (N_2254,N_1518,N_1626);
xor U2255 (N_2255,N_1996,N_1890);
nor U2256 (N_2256,N_1688,N_1839);
or U2257 (N_2257,N_1853,N_1758);
and U2258 (N_2258,N_1513,N_1794);
and U2259 (N_2259,N_1979,N_1802);
xor U2260 (N_2260,N_1693,N_1898);
nor U2261 (N_2261,N_1564,N_1752);
and U2262 (N_2262,N_1790,N_1523);
or U2263 (N_2263,N_1514,N_1595);
nand U2264 (N_2264,N_1715,N_1925);
nand U2265 (N_2265,N_1739,N_1946);
or U2266 (N_2266,N_1822,N_1527);
xnor U2267 (N_2267,N_1831,N_1752);
nand U2268 (N_2268,N_1988,N_1721);
nand U2269 (N_2269,N_1618,N_1700);
nor U2270 (N_2270,N_1987,N_1757);
nor U2271 (N_2271,N_1747,N_1699);
or U2272 (N_2272,N_1731,N_1767);
nor U2273 (N_2273,N_1702,N_1657);
nand U2274 (N_2274,N_1970,N_1525);
and U2275 (N_2275,N_1917,N_1803);
nand U2276 (N_2276,N_1993,N_1958);
nor U2277 (N_2277,N_1666,N_1912);
or U2278 (N_2278,N_1568,N_1676);
nor U2279 (N_2279,N_1966,N_1943);
xnor U2280 (N_2280,N_1935,N_1956);
or U2281 (N_2281,N_1557,N_1930);
or U2282 (N_2282,N_1602,N_1969);
xnor U2283 (N_2283,N_1590,N_1862);
and U2284 (N_2284,N_1589,N_1900);
nand U2285 (N_2285,N_1855,N_1523);
xnor U2286 (N_2286,N_1652,N_1616);
nor U2287 (N_2287,N_1941,N_1813);
or U2288 (N_2288,N_1997,N_1726);
and U2289 (N_2289,N_1764,N_1689);
or U2290 (N_2290,N_1540,N_1883);
or U2291 (N_2291,N_1836,N_1910);
nor U2292 (N_2292,N_1838,N_1571);
and U2293 (N_2293,N_1643,N_1902);
nand U2294 (N_2294,N_1860,N_1584);
nand U2295 (N_2295,N_1665,N_1890);
nand U2296 (N_2296,N_1894,N_1589);
nand U2297 (N_2297,N_1515,N_1866);
nand U2298 (N_2298,N_1831,N_1989);
or U2299 (N_2299,N_1859,N_1943);
xnor U2300 (N_2300,N_1925,N_1615);
xnor U2301 (N_2301,N_1944,N_1948);
and U2302 (N_2302,N_1632,N_1569);
nor U2303 (N_2303,N_1532,N_1784);
nor U2304 (N_2304,N_1750,N_1785);
nand U2305 (N_2305,N_1878,N_1658);
or U2306 (N_2306,N_1822,N_1607);
or U2307 (N_2307,N_1614,N_1839);
or U2308 (N_2308,N_1770,N_1502);
nor U2309 (N_2309,N_1853,N_1569);
and U2310 (N_2310,N_1923,N_1984);
xor U2311 (N_2311,N_1776,N_1909);
and U2312 (N_2312,N_1559,N_1676);
and U2313 (N_2313,N_1998,N_1556);
nand U2314 (N_2314,N_1558,N_1953);
nand U2315 (N_2315,N_1654,N_1798);
and U2316 (N_2316,N_1871,N_1926);
or U2317 (N_2317,N_1960,N_1933);
xnor U2318 (N_2318,N_1640,N_1864);
and U2319 (N_2319,N_1572,N_1760);
and U2320 (N_2320,N_1846,N_1706);
or U2321 (N_2321,N_1806,N_1630);
and U2322 (N_2322,N_1713,N_1679);
xor U2323 (N_2323,N_1642,N_1833);
and U2324 (N_2324,N_1990,N_1936);
nor U2325 (N_2325,N_1859,N_1599);
nand U2326 (N_2326,N_1834,N_1874);
or U2327 (N_2327,N_1737,N_1677);
or U2328 (N_2328,N_1793,N_1609);
nor U2329 (N_2329,N_1542,N_1633);
and U2330 (N_2330,N_1991,N_1736);
xor U2331 (N_2331,N_1902,N_1627);
nor U2332 (N_2332,N_1648,N_1629);
xor U2333 (N_2333,N_1767,N_1793);
and U2334 (N_2334,N_1562,N_1734);
nand U2335 (N_2335,N_1787,N_1996);
nor U2336 (N_2336,N_1908,N_1773);
xnor U2337 (N_2337,N_1695,N_1638);
nor U2338 (N_2338,N_1795,N_1960);
nand U2339 (N_2339,N_1913,N_1569);
nand U2340 (N_2340,N_1893,N_1886);
xnor U2341 (N_2341,N_1770,N_1606);
nand U2342 (N_2342,N_1998,N_1857);
xnor U2343 (N_2343,N_1804,N_1952);
xnor U2344 (N_2344,N_1541,N_1986);
nor U2345 (N_2345,N_1859,N_1804);
and U2346 (N_2346,N_1525,N_1757);
nor U2347 (N_2347,N_1721,N_1817);
and U2348 (N_2348,N_1670,N_1694);
nand U2349 (N_2349,N_1989,N_1669);
nor U2350 (N_2350,N_1678,N_1513);
or U2351 (N_2351,N_1601,N_1963);
and U2352 (N_2352,N_1541,N_1637);
and U2353 (N_2353,N_1885,N_1788);
nor U2354 (N_2354,N_1916,N_1843);
and U2355 (N_2355,N_1749,N_1906);
xnor U2356 (N_2356,N_1869,N_1507);
xor U2357 (N_2357,N_1692,N_1726);
and U2358 (N_2358,N_1820,N_1554);
nor U2359 (N_2359,N_1505,N_1705);
or U2360 (N_2360,N_1663,N_1795);
xnor U2361 (N_2361,N_1545,N_1939);
xor U2362 (N_2362,N_1978,N_1768);
xnor U2363 (N_2363,N_1507,N_1920);
nand U2364 (N_2364,N_1892,N_1681);
nand U2365 (N_2365,N_1893,N_1729);
nand U2366 (N_2366,N_1714,N_1834);
or U2367 (N_2367,N_1898,N_1993);
xnor U2368 (N_2368,N_1980,N_1777);
xnor U2369 (N_2369,N_1889,N_1624);
or U2370 (N_2370,N_1683,N_1504);
nand U2371 (N_2371,N_1554,N_1708);
or U2372 (N_2372,N_1932,N_1804);
xor U2373 (N_2373,N_1843,N_1551);
xor U2374 (N_2374,N_1783,N_1831);
nor U2375 (N_2375,N_1686,N_1519);
xnor U2376 (N_2376,N_1931,N_1856);
or U2377 (N_2377,N_1795,N_1779);
nor U2378 (N_2378,N_1782,N_1672);
nand U2379 (N_2379,N_1723,N_1884);
nor U2380 (N_2380,N_1750,N_1843);
or U2381 (N_2381,N_1682,N_1795);
nand U2382 (N_2382,N_1536,N_1807);
and U2383 (N_2383,N_1758,N_1760);
nand U2384 (N_2384,N_1682,N_1548);
or U2385 (N_2385,N_1844,N_1781);
xnor U2386 (N_2386,N_1801,N_1967);
nor U2387 (N_2387,N_1611,N_1858);
nor U2388 (N_2388,N_1728,N_1563);
or U2389 (N_2389,N_1833,N_1989);
and U2390 (N_2390,N_1965,N_1835);
or U2391 (N_2391,N_1596,N_1937);
or U2392 (N_2392,N_1839,N_1913);
or U2393 (N_2393,N_1584,N_1576);
or U2394 (N_2394,N_1664,N_1570);
and U2395 (N_2395,N_1869,N_1742);
and U2396 (N_2396,N_1551,N_1813);
or U2397 (N_2397,N_1804,N_1808);
or U2398 (N_2398,N_1656,N_1677);
nor U2399 (N_2399,N_1529,N_1893);
xnor U2400 (N_2400,N_1987,N_1654);
xnor U2401 (N_2401,N_1729,N_1794);
and U2402 (N_2402,N_1894,N_1561);
xnor U2403 (N_2403,N_1591,N_1639);
xnor U2404 (N_2404,N_1689,N_1915);
and U2405 (N_2405,N_1752,N_1914);
and U2406 (N_2406,N_1875,N_1551);
or U2407 (N_2407,N_1592,N_1511);
and U2408 (N_2408,N_1501,N_1627);
xnor U2409 (N_2409,N_1627,N_1520);
and U2410 (N_2410,N_1770,N_1958);
nand U2411 (N_2411,N_1975,N_1512);
nand U2412 (N_2412,N_1540,N_1842);
nand U2413 (N_2413,N_1552,N_1507);
and U2414 (N_2414,N_1876,N_1918);
nor U2415 (N_2415,N_1583,N_1708);
nand U2416 (N_2416,N_1757,N_1666);
xnor U2417 (N_2417,N_1819,N_1782);
nor U2418 (N_2418,N_1781,N_1936);
nand U2419 (N_2419,N_1573,N_1586);
xor U2420 (N_2420,N_1899,N_1550);
nor U2421 (N_2421,N_1937,N_1583);
nor U2422 (N_2422,N_1753,N_1563);
nand U2423 (N_2423,N_1816,N_1582);
or U2424 (N_2424,N_1610,N_1814);
nor U2425 (N_2425,N_1621,N_1843);
and U2426 (N_2426,N_1781,N_1508);
and U2427 (N_2427,N_1584,N_1692);
xor U2428 (N_2428,N_1766,N_1728);
nand U2429 (N_2429,N_1569,N_1957);
and U2430 (N_2430,N_1816,N_1604);
nor U2431 (N_2431,N_1713,N_1932);
xnor U2432 (N_2432,N_1536,N_1905);
nor U2433 (N_2433,N_1810,N_1816);
nor U2434 (N_2434,N_1965,N_1964);
nor U2435 (N_2435,N_1997,N_1659);
nand U2436 (N_2436,N_1864,N_1906);
and U2437 (N_2437,N_1655,N_1542);
and U2438 (N_2438,N_1951,N_1888);
nor U2439 (N_2439,N_1801,N_1615);
nand U2440 (N_2440,N_1832,N_1677);
nand U2441 (N_2441,N_1784,N_1569);
xnor U2442 (N_2442,N_1785,N_1597);
nor U2443 (N_2443,N_1834,N_1504);
xnor U2444 (N_2444,N_1946,N_1807);
and U2445 (N_2445,N_1523,N_1772);
and U2446 (N_2446,N_1790,N_1784);
xor U2447 (N_2447,N_1948,N_1606);
or U2448 (N_2448,N_1714,N_1967);
nand U2449 (N_2449,N_1507,N_1956);
or U2450 (N_2450,N_1878,N_1569);
nor U2451 (N_2451,N_1838,N_1905);
or U2452 (N_2452,N_1840,N_1926);
nor U2453 (N_2453,N_1878,N_1703);
and U2454 (N_2454,N_1941,N_1867);
nor U2455 (N_2455,N_1928,N_1604);
xor U2456 (N_2456,N_1670,N_1518);
or U2457 (N_2457,N_1850,N_1546);
or U2458 (N_2458,N_1996,N_1969);
nand U2459 (N_2459,N_1896,N_1554);
xnor U2460 (N_2460,N_1956,N_1866);
nor U2461 (N_2461,N_1886,N_1787);
and U2462 (N_2462,N_1573,N_1979);
nand U2463 (N_2463,N_1684,N_1552);
nor U2464 (N_2464,N_1995,N_1717);
xor U2465 (N_2465,N_1506,N_1528);
or U2466 (N_2466,N_1659,N_1873);
or U2467 (N_2467,N_1672,N_1679);
nand U2468 (N_2468,N_1609,N_1817);
and U2469 (N_2469,N_1544,N_1805);
xnor U2470 (N_2470,N_1667,N_1676);
nand U2471 (N_2471,N_1523,N_1793);
nand U2472 (N_2472,N_1809,N_1626);
or U2473 (N_2473,N_1540,N_1832);
nor U2474 (N_2474,N_1755,N_1512);
or U2475 (N_2475,N_1613,N_1570);
xor U2476 (N_2476,N_1603,N_1713);
nand U2477 (N_2477,N_1511,N_1567);
xor U2478 (N_2478,N_1943,N_1728);
xnor U2479 (N_2479,N_1763,N_1675);
nor U2480 (N_2480,N_1661,N_1550);
xnor U2481 (N_2481,N_1861,N_1601);
and U2482 (N_2482,N_1581,N_1767);
nand U2483 (N_2483,N_1633,N_1804);
xor U2484 (N_2484,N_1995,N_1827);
nor U2485 (N_2485,N_1984,N_1750);
nor U2486 (N_2486,N_1757,N_1553);
nand U2487 (N_2487,N_1628,N_1959);
and U2488 (N_2488,N_1542,N_1734);
nand U2489 (N_2489,N_1566,N_1860);
or U2490 (N_2490,N_1790,N_1969);
nand U2491 (N_2491,N_1630,N_1943);
xor U2492 (N_2492,N_1751,N_1752);
and U2493 (N_2493,N_1903,N_1614);
nor U2494 (N_2494,N_1856,N_1956);
and U2495 (N_2495,N_1677,N_1637);
nand U2496 (N_2496,N_1685,N_1930);
nor U2497 (N_2497,N_1829,N_1895);
nand U2498 (N_2498,N_1866,N_1639);
nand U2499 (N_2499,N_1695,N_1715);
nor U2500 (N_2500,N_2067,N_2087);
xor U2501 (N_2501,N_2138,N_2425);
xor U2502 (N_2502,N_2491,N_2146);
and U2503 (N_2503,N_2160,N_2251);
nand U2504 (N_2504,N_2119,N_2113);
nand U2505 (N_2505,N_2226,N_2098);
nand U2506 (N_2506,N_2400,N_2244);
nand U2507 (N_2507,N_2132,N_2124);
or U2508 (N_2508,N_2062,N_2332);
nor U2509 (N_2509,N_2191,N_2478);
or U2510 (N_2510,N_2105,N_2014);
nor U2511 (N_2511,N_2279,N_2116);
and U2512 (N_2512,N_2430,N_2088);
or U2513 (N_2513,N_2018,N_2225);
or U2514 (N_2514,N_2338,N_2096);
nor U2515 (N_2515,N_2056,N_2083);
and U2516 (N_2516,N_2195,N_2493);
xnor U2517 (N_2517,N_2097,N_2368);
and U2518 (N_2518,N_2261,N_2084);
xnor U2519 (N_2519,N_2071,N_2199);
xnor U2520 (N_2520,N_2273,N_2416);
nand U2521 (N_2521,N_2396,N_2323);
nor U2522 (N_2522,N_2085,N_2488);
or U2523 (N_2523,N_2026,N_2398);
nand U2524 (N_2524,N_2187,N_2005);
xnor U2525 (N_2525,N_2100,N_2315);
and U2526 (N_2526,N_2209,N_2143);
xnor U2527 (N_2527,N_2412,N_2344);
and U2528 (N_2528,N_2134,N_2269);
nand U2529 (N_2529,N_2294,N_2431);
nor U2530 (N_2530,N_2079,N_2301);
or U2531 (N_2531,N_2008,N_2059);
or U2532 (N_2532,N_2043,N_2406);
and U2533 (N_2533,N_2200,N_2420);
xnor U2534 (N_2534,N_2361,N_2211);
xor U2535 (N_2535,N_2466,N_2000);
and U2536 (N_2536,N_2296,N_2122);
or U2537 (N_2537,N_2437,N_2024);
and U2538 (N_2538,N_2252,N_2287);
and U2539 (N_2539,N_2066,N_2190);
xnor U2540 (N_2540,N_2401,N_2475);
xnor U2541 (N_2541,N_2048,N_2374);
or U2542 (N_2542,N_2135,N_2417);
xor U2543 (N_2543,N_2265,N_2064);
xor U2544 (N_2544,N_2073,N_2045);
xnor U2545 (N_2545,N_2293,N_2237);
xnor U2546 (N_2546,N_2485,N_2189);
xnor U2547 (N_2547,N_2305,N_2490);
xnor U2548 (N_2548,N_2164,N_2458);
xor U2549 (N_2549,N_2214,N_2072);
nor U2550 (N_2550,N_2057,N_2384);
xnor U2551 (N_2551,N_2317,N_2013);
nand U2552 (N_2552,N_2354,N_2250);
or U2553 (N_2553,N_2445,N_2419);
nand U2554 (N_2554,N_2010,N_2314);
nand U2555 (N_2555,N_2335,N_2110);
and U2556 (N_2556,N_2223,N_2373);
nand U2557 (N_2557,N_2347,N_2175);
nor U2558 (N_2558,N_2179,N_2452);
xnor U2559 (N_2559,N_2203,N_2345);
and U2560 (N_2560,N_2463,N_2234);
and U2561 (N_2561,N_2304,N_2258);
and U2562 (N_2562,N_2140,N_2394);
and U2563 (N_2563,N_2230,N_2240);
xnor U2564 (N_2564,N_2442,N_2220);
xor U2565 (N_2565,N_2016,N_2356);
nand U2566 (N_2566,N_2102,N_2464);
xnor U2567 (N_2567,N_2242,N_2031);
and U2568 (N_2568,N_2451,N_2413);
nor U2569 (N_2569,N_2041,N_2131);
nand U2570 (N_2570,N_2217,N_2108);
nand U2571 (N_2571,N_2393,N_2241);
nor U2572 (N_2572,N_2178,N_2070);
xor U2573 (N_2573,N_2353,N_2465);
or U2574 (N_2574,N_2007,N_2228);
or U2575 (N_2575,N_2243,N_2063);
xor U2576 (N_2576,N_2263,N_2144);
xnor U2577 (N_2577,N_2205,N_2290);
or U2578 (N_2578,N_2486,N_2415);
or U2579 (N_2579,N_2389,N_2403);
and U2580 (N_2580,N_2029,N_2471);
and U2581 (N_2581,N_2081,N_2065);
nand U2582 (N_2582,N_2327,N_2499);
or U2583 (N_2583,N_2111,N_2280);
and U2584 (N_2584,N_2362,N_2307);
and U2585 (N_2585,N_2422,N_2109);
xor U2586 (N_2586,N_2216,N_2391);
nor U2587 (N_2587,N_2245,N_2208);
nand U2588 (N_2588,N_2408,N_2174);
nand U2589 (N_2589,N_2274,N_2038);
nor U2590 (N_2590,N_2002,N_2232);
xor U2591 (N_2591,N_2346,N_2318);
nor U2592 (N_2592,N_2027,N_2473);
nand U2593 (N_2593,N_2341,N_2333);
nand U2594 (N_2594,N_2297,N_2104);
and U2595 (N_2595,N_2162,N_2141);
nor U2596 (N_2596,N_2308,N_2103);
or U2597 (N_2597,N_2054,N_2120);
xor U2598 (N_2598,N_2061,N_2494);
xor U2599 (N_2599,N_2192,N_2198);
nand U2600 (N_2600,N_2432,N_2249);
or U2601 (N_2601,N_2435,N_2363);
and U2602 (N_2602,N_2311,N_2246);
and U2603 (N_2603,N_2371,N_2260);
and U2604 (N_2604,N_2278,N_2201);
nand U2605 (N_2605,N_2316,N_2348);
or U2606 (N_2606,N_2276,N_2227);
nor U2607 (N_2607,N_2414,N_2009);
nor U2608 (N_2608,N_2309,N_2441);
and U2609 (N_2609,N_2476,N_2028);
nand U2610 (N_2610,N_2117,N_2331);
xnor U2611 (N_2611,N_2106,N_2044);
nor U2612 (N_2612,N_2447,N_2042);
nor U2613 (N_2613,N_2453,N_2090);
xor U2614 (N_2614,N_2277,N_2112);
nor U2615 (N_2615,N_2154,N_2367);
nor U2616 (N_2616,N_2325,N_2129);
xor U2617 (N_2617,N_2236,N_2051);
nand U2618 (N_2618,N_2372,N_2218);
nand U2619 (N_2619,N_2019,N_2456);
nand U2620 (N_2620,N_2498,N_2349);
nand U2621 (N_2621,N_2259,N_2186);
nand U2622 (N_2622,N_2350,N_2233);
xor U2623 (N_2623,N_2376,N_2310);
nor U2624 (N_2624,N_2411,N_2180);
and U2625 (N_2625,N_2383,N_2188);
xor U2626 (N_2626,N_2182,N_2221);
nor U2627 (N_2627,N_2262,N_2254);
nand U2628 (N_2628,N_2365,N_2155);
and U2629 (N_2629,N_2171,N_2428);
nand U2630 (N_2630,N_2388,N_2324);
nor U2631 (N_2631,N_2282,N_2337);
and U2632 (N_2632,N_2101,N_2358);
xor U2633 (N_2633,N_2046,N_2118);
xor U2634 (N_2634,N_2424,N_2012);
nor U2635 (N_2635,N_2001,N_2484);
or U2636 (N_2636,N_2421,N_2352);
xor U2637 (N_2637,N_2397,N_2379);
nand U2638 (N_2638,N_2257,N_2446);
xor U2639 (N_2639,N_2342,N_2093);
xnor U2640 (N_2640,N_2266,N_2480);
nand U2641 (N_2641,N_2039,N_2288);
and U2642 (N_2642,N_2213,N_2015);
or U2643 (N_2643,N_2040,N_2099);
xnor U2644 (N_2644,N_2443,N_2074);
and U2645 (N_2645,N_2137,N_2395);
nor U2646 (N_2646,N_2239,N_2272);
or U2647 (N_2647,N_2334,N_2444);
nor U2648 (N_2648,N_2482,N_2173);
xnor U2649 (N_2649,N_2436,N_2434);
nand U2650 (N_2650,N_2461,N_2405);
nor U2651 (N_2651,N_2433,N_2380);
nor U2652 (N_2652,N_2459,N_2210);
or U2653 (N_2653,N_2483,N_2360);
or U2654 (N_2654,N_2133,N_2387);
or U2655 (N_2655,N_2336,N_2247);
xnor U2656 (N_2656,N_2091,N_2364);
nor U2657 (N_2657,N_2429,N_2033);
xnor U2658 (N_2658,N_2238,N_2080);
or U2659 (N_2659,N_2145,N_2060);
nand U2660 (N_2660,N_2130,N_2271);
nand U2661 (N_2661,N_2219,N_2298);
xor U2662 (N_2662,N_2340,N_2303);
nand U2663 (N_2663,N_2017,N_2114);
nand U2664 (N_2664,N_2121,N_2055);
nor U2665 (N_2665,N_2032,N_2047);
nand U2666 (N_2666,N_2256,N_2231);
xnor U2667 (N_2667,N_2163,N_2177);
or U2668 (N_2668,N_2150,N_2169);
xor U2669 (N_2669,N_2194,N_2127);
nor U2670 (N_2670,N_2184,N_2082);
or U2671 (N_2671,N_2495,N_2496);
xor U2672 (N_2672,N_2284,N_2455);
xor U2673 (N_2673,N_2181,N_2193);
and U2674 (N_2674,N_2107,N_2022);
and U2675 (N_2675,N_2479,N_2215);
or U2676 (N_2676,N_2440,N_2390);
and U2677 (N_2677,N_2165,N_2075);
or U2678 (N_2678,N_2086,N_2438);
or U2679 (N_2679,N_2196,N_2283);
or U2680 (N_2680,N_2222,N_2460);
and U2681 (N_2681,N_2248,N_2281);
xor U2682 (N_2682,N_2370,N_2004);
or U2683 (N_2683,N_2381,N_2030);
nand U2684 (N_2684,N_2185,N_2168);
xor U2685 (N_2685,N_2142,N_2253);
xnor U2686 (N_2686,N_2123,N_2212);
and U2687 (N_2687,N_2094,N_2462);
and U2688 (N_2688,N_2025,N_2404);
nand U2689 (N_2689,N_2170,N_2302);
or U2690 (N_2690,N_2295,N_2300);
and U2691 (N_2691,N_2407,N_2052);
nand U2692 (N_2692,N_2003,N_2357);
nand U2693 (N_2693,N_2322,N_2439);
or U2694 (N_2694,N_2126,N_2158);
or U2695 (N_2695,N_2313,N_2312);
nand U2696 (N_2696,N_2448,N_2021);
xnor U2697 (N_2697,N_2204,N_2399);
nor U2698 (N_2698,N_2006,N_2343);
nand U2699 (N_2699,N_2267,N_2469);
and U2700 (N_2700,N_2377,N_2151);
xnor U2701 (N_2701,N_2050,N_2139);
and U2702 (N_2702,N_2034,N_2382);
nand U2703 (N_2703,N_2092,N_2418);
or U2704 (N_2704,N_2049,N_2229);
and U2705 (N_2705,N_2076,N_2197);
xnor U2706 (N_2706,N_2449,N_2176);
or U2707 (N_2707,N_2023,N_2264);
nand U2708 (N_2708,N_2069,N_2078);
and U2709 (N_2709,N_2206,N_2329);
xor U2710 (N_2710,N_2147,N_2474);
or U2711 (N_2711,N_2423,N_2077);
nor U2712 (N_2712,N_2156,N_2068);
and U2713 (N_2713,N_2351,N_2157);
nor U2714 (N_2714,N_2489,N_2454);
or U2715 (N_2715,N_2089,N_2320);
nor U2716 (N_2716,N_2053,N_2450);
nand U2717 (N_2717,N_2328,N_2224);
xor U2718 (N_2718,N_2286,N_2481);
xor U2719 (N_2719,N_2035,N_2319);
xor U2720 (N_2720,N_2159,N_2402);
or U2721 (N_2721,N_2306,N_2153);
nor U2722 (N_2722,N_2020,N_2235);
nor U2723 (N_2723,N_2148,N_2472);
nand U2724 (N_2724,N_2292,N_2299);
or U2725 (N_2725,N_2477,N_2410);
nor U2726 (N_2726,N_2369,N_2275);
or U2727 (N_2727,N_2161,N_2385);
and U2728 (N_2728,N_2011,N_2375);
xor U2729 (N_2729,N_2321,N_2285);
and U2730 (N_2730,N_2289,N_2427);
or U2731 (N_2731,N_2378,N_2392);
nand U2732 (N_2732,N_2470,N_2202);
xor U2733 (N_2733,N_2409,N_2128);
or U2734 (N_2734,N_2457,N_2339);
and U2735 (N_2735,N_2037,N_2136);
or U2736 (N_2736,N_2207,N_2036);
and U2737 (N_2737,N_2468,N_2291);
nand U2738 (N_2738,N_2115,N_2330);
and U2739 (N_2739,N_2255,N_2125);
and U2740 (N_2740,N_2166,N_2492);
and U2741 (N_2741,N_2426,N_2326);
xor U2742 (N_2742,N_2487,N_2058);
and U2743 (N_2743,N_2366,N_2270);
xor U2744 (N_2744,N_2149,N_2386);
or U2745 (N_2745,N_2183,N_2497);
nand U2746 (N_2746,N_2152,N_2172);
or U2747 (N_2747,N_2268,N_2355);
and U2748 (N_2748,N_2467,N_2359);
nor U2749 (N_2749,N_2095,N_2167);
nand U2750 (N_2750,N_2164,N_2451);
or U2751 (N_2751,N_2315,N_2340);
nand U2752 (N_2752,N_2327,N_2210);
and U2753 (N_2753,N_2498,N_2148);
nor U2754 (N_2754,N_2011,N_2447);
or U2755 (N_2755,N_2222,N_2388);
and U2756 (N_2756,N_2171,N_2306);
xor U2757 (N_2757,N_2126,N_2141);
or U2758 (N_2758,N_2120,N_2041);
xor U2759 (N_2759,N_2308,N_2239);
nand U2760 (N_2760,N_2353,N_2089);
nand U2761 (N_2761,N_2375,N_2337);
nand U2762 (N_2762,N_2404,N_2153);
and U2763 (N_2763,N_2261,N_2488);
or U2764 (N_2764,N_2280,N_2000);
and U2765 (N_2765,N_2338,N_2000);
nor U2766 (N_2766,N_2055,N_2273);
nor U2767 (N_2767,N_2449,N_2151);
nand U2768 (N_2768,N_2007,N_2464);
xnor U2769 (N_2769,N_2260,N_2082);
nor U2770 (N_2770,N_2074,N_2101);
and U2771 (N_2771,N_2101,N_2440);
or U2772 (N_2772,N_2474,N_2055);
and U2773 (N_2773,N_2086,N_2212);
xor U2774 (N_2774,N_2089,N_2067);
or U2775 (N_2775,N_2324,N_2272);
nor U2776 (N_2776,N_2369,N_2438);
nand U2777 (N_2777,N_2248,N_2315);
nor U2778 (N_2778,N_2046,N_2105);
and U2779 (N_2779,N_2224,N_2369);
nand U2780 (N_2780,N_2399,N_2488);
nor U2781 (N_2781,N_2044,N_2458);
or U2782 (N_2782,N_2351,N_2045);
nor U2783 (N_2783,N_2215,N_2154);
xor U2784 (N_2784,N_2167,N_2130);
or U2785 (N_2785,N_2414,N_2221);
or U2786 (N_2786,N_2063,N_2272);
and U2787 (N_2787,N_2006,N_2162);
nor U2788 (N_2788,N_2123,N_2104);
nor U2789 (N_2789,N_2270,N_2236);
or U2790 (N_2790,N_2338,N_2282);
nor U2791 (N_2791,N_2436,N_2343);
or U2792 (N_2792,N_2222,N_2033);
or U2793 (N_2793,N_2288,N_2258);
xor U2794 (N_2794,N_2032,N_2218);
xnor U2795 (N_2795,N_2333,N_2012);
nand U2796 (N_2796,N_2144,N_2195);
nand U2797 (N_2797,N_2126,N_2365);
and U2798 (N_2798,N_2186,N_2087);
nand U2799 (N_2799,N_2165,N_2074);
or U2800 (N_2800,N_2031,N_2385);
nand U2801 (N_2801,N_2087,N_2016);
nand U2802 (N_2802,N_2254,N_2255);
nand U2803 (N_2803,N_2325,N_2014);
or U2804 (N_2804,N_2022,N_2301);
nor U2805 (N_2805,N_2079,N_2447);
xnor U2806 (N_2806,N_2224,N_2197);
or U2807 (N_2807,N_2244,N_2406);
nand U2808 (N_2808,N_2282,N_2465);
nand U2809 (N_2809,N_2159,N_2321);
or U2810 (N_2810,N_2347,N_2354);
nand U2811 (N_2811,N_2059,N_2403);
or U2812 (N_2812,N_2122,N_2480);
nand U2813 (N_2813,N_2239,N_2138);
and U2814 (N_2814,N_2430,N_2034);
and U2815 (N_2815,N_2207,N_2071);
or U2816 (N_2816,N_2239,N_2002);
or U2817 (N_2817,N_2347,N_2393);
nand U2818 (N_2818,N_2018,N_2486);
or U2819 (N_2819,N_2446,N_2015);
xor U2820 (N_2820,N_2395,N_2076);
and U2821 (N_2821,N_2178,N_2192);
xor U2822 (N_2822,N_2348,N_2414);
nor U2823 (N_2823,N_2065,N_2099);
nand U2824 (N_2824,N_2447,N_2359);
nand U2825 (N_2825,N_2248,N_2262);
and U2826 (N_2826,N_2495,N_2498);
nand U2827 (N_2827,N_2114,N_2134);
xor U2828 (N_2828,N_2445,N_2410);
xor U2829 (N_2829,N_2312,N_2404);
and U2830 (N_2830,N_2461,N_2040);
or U2831 (N_2831,N_2462,N_2240);
xor U2832 (N_2832,N_2358,N_2150);
nand U2833 (N_2833,N_2117,N_2305);
and U2834 (N_2834,N_2283,N_2157);
or U2835 (N_2835,N_2439,N_2343);
nand U2836 (N_2836,N_2038,N_2341);
or U2837 (N_2837,N_2332,N_2402);
nor U2838 (N_2838,N_2037,N_2099);
nor U2839 (N_2839,N_2241,N_2339);
or U2840 (N_2840,N_2042,N_2108);
nand U2841 (N_2841,N_2154,N_2298);
or U2842 (N_2842,N_2474,N_2053);
nand U2843 (N_2843,N_2437,N_2149);
nand U2844 (N_2844,N_2474,N_2266);
nor U2845 (N_2845,N_2410,N_2174);
nand U2846 (N_2846,N_2321,N_2460);
nand U2847 (N_2847,N_2376,N_2377);
nor U2848 (N_2848,N_2253,N_2185);
nand U2849 (N_2849,N_2090,N_2413);
nor U2850 (N_2850,N_2287,N_2172);
xor U2851 (N_2851,N_2309,N_2256);
and U2852 (N_2852,N_2380,N_2189);
nand U2853 (N_2853,N_2124,N_2173);
or U2854 (N_2854,N_2265,N_2250);
nor U2855 (N_2855,N_2038,N_2311);
nor U2856 (N_2856,N_2118,N_2387);
nor U2857 (N_2857,N_2355,N_2187);
or U2858 (N_2858,N_2323,N_2382);
and U2859 (N_2859,N_2373,N_2433);
or U2860 (N_2860,N_2012,N_2050);
nor U2861 (N_2861,N_2179,N_2335);
and U2862 (N_2862,N_2004,N_2089);
and U2863 (N_2863,N_2170,N_2484);
or U2864 (N_2864,N_2477,N_2397);
nand U2865 (N_2865,N_2329,N_2318);
nor U2866 (N_2866,N_2275,N_2174);
nor U2867 (N_2867,N_2304,N_2455);
xnor U2868 (N_2868,N_2177,N_2175);
or U2869 (N_2869,N_2491,N_2126);
xnor U2870 (N_2870,N_2445,N_2191);
or U2871 (N_2871,N_2374,N_2241);
xnor U2872 (N_2872,N_2362,N_2424);
nand U2873 (N_2873,N_2073,N_2130);
xnor U2874 (N_2874,N_2302,N_2243);
nand U2875 (N_2875,N_2290,N_2479);
nand U2876 (N_2876,N_2121,N_2115);
nand U2877 (N_2877,N_2391,N_2421);
nand U2878 (N_2878,N_2268,N_2426);
nor U2879 (N_2879,N_2297,N_2156);
nand U2880 (N_2880,N_2146,N_2256);
xnor U2881 (N_2881,N_2208,N_2256);
or U2882 (N_2882,N_2237,N_2177);
or U2883 (N_2883,N_2162,N_2130);
xnor U2884 (N_2884,N_2239,N_2289);
or U2885 (N_2885,N_2259,N_2326);
and U2886 (N_2886,N_2044,N_2061);
xor U2887 (N_2887,N_2276,N_2414);
and U2888 (N_2888,N_2254,N_2435);
nand U2889 (N_2889,N_2167,N_2054);
nand U2890 (N_2890,N_2067,N_2247);
xnor U2891 (N_2891,N_2180,N_2363);
or U2892 (N_2892,N_2128,N_2366);
nor U2893 (N_2893,N_2489,N_2127);
nor U2894 (N_2894,N_2318,N_2007);
xnor U2895 (N_2895,N_2142,N_2428);
xnor U2896 (N_2896,N_2219,N_2389);
and U2897 (N_2897,N_2096,N_2034);
xor U2898 (N_2898,N_2226,N_2155);
nand U2899 (N_2899,N_2024,N_2460);
or U2900 (N_2900,N_2375,N_2293);
xnor U2901 (N_2901,N_2176,N_2266);
nand U2902 (N_2902,N_2316,N_2198);
or U2903 (N_2903,N_2323,N_2058);
and U2904 (N_2904,N_2451,N_2425);
xor U2905 (N_2905,N_2065,N_2203);
and U2906 (N_2906,N_2499,N_2412);
nand U2907 (N_2907,N_2352,N_2189);
or U2908 (N_2908,N_2222,N_2137);
xor U2909 (N_2909,N_2435,N_2280);
xnor U2910 (N_2910,N_2328,N_2278);
and U2911 (N_2911,N_2416,N_2008);
xnor U2912 (N_2912,N_2245,N_2450);
xor U2913 (N_2913,N_2026,N_2312);
nor U2914 (N_2914,N_2385,N_2017);
nand U2915 (N_2915,N_2489,N_2280);
xnor U2916 (N_2916,N_2290,N_2087);
xor U2917 (N_2917,N_2220,N_2321);
nand U2918 (N_2918,N_2271,N_2458);
or U2919 (N_2919,N_2136,N_2096);
or U2920 (N_2920,N_2370,N_2421);
or U2921 (N_2921,N_2178,N_2438);
nand U2922 (N_2922,N_2216,N_2354);
nor U2923 (N_2923,N_2056,N_2400);
and U2924 (N_2924,N_2001,N_2097);
xor U2925 (N_2925,N_2452,N_2277);
nor U2926 (N_2926,N_2310,N_2481);
and U2927 (N_2927,N_2022,N_2106);
xnor U2928 (N_2928,N_2142,N_2368);
and U2929 (N_2929,N_2352,N_2195);
nand U2930 (N_2930,N_2148,N_2058);
xor U2931 (N_2931,N_2009,N_2384);
nand U2932 (N_2932,N_2490,N_2387);
nand U2933 (N_2933,N_2442,N_2117);
nor U2934 (N_2934,N_2052,N_2471);
xnor U2935 (N_2935,N_2031,N_2200);
xnor U2936 (N_2936,N_2431,N_2138);
xor U2937 (N_2937,N_2393,N_2137);
nor U2938 (N_2938,N_2048,N_2432);
nor U2939 (N_2939,N_2192,N_2349);
nor U2940 (N_2940,N_2264,N_2301);
xnor U2941 (N_2941,N_2139,N_2294);
nor U2942 (N_2942,N_2386,N_2277);
and U2943 (N_2943,N_2134,N_2103);
nand U2944 (N_2944,N_2217,N_2294);
xor U2945 (N_2945,N_2442,N_2064);
and U2946 (N_2946,N_2444,N_2427);
nor U2947 (N_2947,N_2250,N_2234);
or U2948 (N_2948,N_2479,N_2072);
and U2949 (N_2949,N_2173,N_2065);
and U2950 (N_2950,N_2491,N_2110);
xor U2951 (N_2951,N_2459,N_2297);
xor U2952 (N_2952,N_2016,N_2359);
xnor U2953 (N_2953,N_2379,N_2442);
or U2954 (N_2954,N_2365,N_2187);
nand U2955 (N_2955,N_2356,N_2116);
nor U2956 (N_2956,N_2413,N_2284);
xor U2957 (N_2957,N_2475,N_2487);
or U2958 (N_2958,N_2201,N_2337);
and U2959 (N_2959,N_2152,N_2477);
nor U2960 (N_2960,N_2069,N_2020);
nand U2961 (N_2961,N_2175,N_2443);
and U2962 (N_2962,N_2245,N_2239);
xor U2963 (N_2963,N_2171,N_2385);
nor U2964 (N_2964,N_2086,N_2147);
nand U2965 (N_2965,N_2071,N_2455);
xor U2966 (N_2966,N_2192,N_2394);
or U2967 (N_2967,N_2329,N_2317);
nand U2968 (N_2968,N_2289,N_2181);
and U2969 (N_2969,N_2159,N_2200);
nand U2970 (N_2970,N_2084,N_2208);
or U2971 (N_2971,N_2380,N_2247);
nor U2972 (N_2972,N_2248,N_2437);
nor U2973 (N_2973,N_2144,N_2140);
xor U2974 (N_2974,N_2332,N_2486);
or U2975 (N_2975,N_2209,N_2339);
xnor U2976 (N_2976,N_2052,N_2143);
nor U2977 (N_2977,N_2428,N_2033);
or U2978 (N_2978,N_2218,N_2357);
and U2979 (N_2979,N_2086,N_2299);
or U2980 (N_2980,N_2306,N_2168);
nor U2981 (N_2981,N_2034,N_2019);
and U2982 (N_2982,N_2270,N_2331);
nand U2983 (N_2983,N_2377,N_2169);
or U2984 (N_2984,N_2169,N_2434);
xnor U2985 (N_2985,N_2370,N_2334);
nor U2986 (N_2986,N_2003,N_2047);
or U2987 (N_2987,N_2064,N_2491);
nor U2988 (N_2988,N_2235,N_2107);
nor U2989 (N_2989,N_2176,N_2190);
nand U2990 (N_2990,N_2382,N_2096);
xor U2991 (N_2991,N_2261,N_2051);
xnor U2992 (N_2992,N_2218,N_2258);
and U2993 (N_2993,N_2061,N_2057);
nand U2994 (N_2994,N_2262,N_2380);
nor U2995 (N_2995,N_2197,N_2177);
xor U2996 (N_2996,N_2058,N_2291);
nor U2997 (N_2997,N_2479,N_2071);
or U2998 (N_2998,N_2366,N_2337);
xor U2999 (N_2999,N_2180,N_2276);
xor U3000 (N_3000,N_2689,N_2614);
xnor U3001 (N_3001,N_2609,N_2652);
xor U3002 (N_3002,N_2538,N_2997);
or U3003 (N_3003,N_2677,N_2845);
nor U3004 (N_3004,N_2669,N_2617);
nor U3005 (N_3005,N_2923,N_2661);
nand U3006 (N_3006,N_2968,N_2817);
and U3007 (N_3007,N_2980,N_2671);
nand U3008 (N_3008,N_2588,N_2935);
nor U3009 (N_3009,N_2673,N_2561);
nand U3010 (N_3010,N_2631,N_2909);
nor U3011 (N_3011,N_2873,N_2889);
or U3012 (N_3012,N_2762,N_2828);
nor U3013 (N_3013,N_2637,N_2535);
or U3014 (N_3014,N_2999,N_2901);
xnor U3015 (N_3015,N_2994,N_2896);
and U3016 (N_3016,N_2945,N_2589);
and U3017 (N_3017,N_2960,N_2519);
nor U3018 (N_3018,N_2773,N_2978);
and U3019 (N_3019,N_2686,N_2862);
nand U3020 (N_3020,N_2894,N_2648);
nor U3021 (N_3021,N_2606,N_2750);
and U3022 (N_3022,N_2787,N_2825);
nand U3023 (N_3023,N_2580,N_2629);
or U3024 (N_3024,N_2786,N_2914);
and U3025 (N_3025,N_2537,N_2848);
and U3026 (N_3026,N_2663,N_2760);
nand U3027 (N_3027,N_2613,N_2685);
nand U3028 (N_3028,N_2586,N_2579);
nor U3029 (N_3029,N_2619,N_2986);
and U3030 (N_3030,N_2932,N_2527);
xnor U3031 (N_3031,N_2902,N_2566);
xnor U3032 (N_3032,N_2983,N_2700);
or U3033 (N_3033,N_2584,N_2822);
nand U3034 (N_3034,N_2670,N_2951);
xnor U3035 (N_3035,N_2948,N_2805);
nand U3036 (N_3036,N_2938,N_2975);
or U3037 (N_3037,N_2747,N_2879);
or U3038 (N_3038,N_2856,N_2716);
xnor U3039 (N_3039,N_2577,N_2831);
and U3040 (N_3040,N_2912,N_2963);
or U3041 (N_3041,N_2749,N_2735);
and U3042 (N_3042,N_2859,N_2529);
and U3043 (N_3043,N_2723,N_2719);
nor U3044 (N_3044,N_2953,N_2815);
nor U3045 (N_3045,N_2849,N_2746);
nor U3046 (N_3046,N_2816,N_2811);
nand U3047 (N_3047,N_2563,N_2585);
xor U3048 (N_3048,N_2634,N_2501);
and U3049 (N_3049,N_2989,N_2868);
or U3050 (N_3050,N_2515,N_2688);
and U3051 (N_3051,N_2682,N_2984);
xor U3052 (N_3052,N_2844,N_2924);
or U3053 (N_3053,N_2581,N_2667);
xnor U3054 (N_3054,N_2572,N_2954);
xnor U3055 (N_3055,N_2630,N_2740);
or U3056 (N_3056,N_2635,N_2722);
nand U3057 (N_3057,N_2709,N_2744);
nor U3058 (N_3058,N_2647,N_2540);
xor U3059 (N_3059,N_2564,N_2644);
nand U3060 (N_3060,N_2990,N_2513);
nor U3061 (N_3061,N_2509,N_2827);
nor U3062 (N_3062,N_2737,N_2927);
and U3063 (N_3063,N_2718,N_2905);
or U3064 (N_3064,N_2866,N_2952);
or U3065 (N_3065,N_2610,N_2778);
nor U3066 (N_3066,N_2597,N_2941);
or U3067 (N_3067,N_2721,N_2955);
nor U3068 (N_3068,N_2521,N_2857);
nand U3069 (N_3069,N_2576,N_2895);
nor U3070 (N_3070,N_2777,N_2712);
and U3071 (N_3071,N_2771,N_2818);
or U3072 (N_3072,N_2690,N_2979);
xnor U3073 (N_3073,N_2824,N_2969);
and U3074 (N_3074,N_2706,N_2957);
nand U3075 (N_3075,N_2591,N_2510);
nor U3076 (N_3076,N_2594,N_2664);
nor U3077 (N_3077,N_2539,N_2803);
nand U3078 (N_3078,N_2823,N_2812);
nand U3079 (N_3079,N_2867,N_2517);
or U3080 (N_3080,N_2639,N_2885);
xnor U3081 (N_3081,N_2813,N_2720);
nand U3082 (N_3082,N_2928,N_2904);
and U3083 (N_3083,N_2869,N_2684);
or U3084 (N_3084,N_2833,N_2791);
and U3085 (N_3085,N_2583,N_2651);
and U3086 (N_3086,N_2657,N_2615);
xnor U3087 (N_3087,N_2917,N_2695);
and U3088 (N_3088,N_2679,N_2939);
nor U3089 (N_3089,N_2621,N_2769);
nand U3090 (N_3090,N_2533,N_2881);
or U3091 (N_3091,N_2626,N_2870);
nor U3092 (N_3092,N_2542,N_2708);
nor U3093 (N_3093,N_2875,N_2699);
xnor U3094 (N_3094,N_2784,N_2593);
nor U3095 (N_3095,N_2654,N_2961);
nor U3096 (N_3096,N_2692,N_2571);
or U3097 (N_3097,N_2887,N_2755);
and U3098 (N_3098,N_2906,N_2587);
and U3099 (N_3099,N_2618,N_2996);
or U3100 (N_3100,N_2544,N_2508);
xor U3101 (N_3101,N_2855,N_2506);
nor U3102 (N_3102,N_2525,N_2876);
and U3103 (N_3103,N_2764,N_2713);
nand U3104 (N_3104,N_2570,N_2920);
and U3105 (N_3105,N_2897,N_2836);
and U3106 (N_3106,N_2977,N_2925);
or U3107 (N_3107,N_2504,N_2877);
and U3108 (N_3108,N_2554,N_2810);
nor U3109 (N_3109,N_2505,N_2569);
and U3110 (N_3110,N_2582,N_2972);
xnor U3111 (N_3111,N_2809,N_2853);
xor U3112 (N_3112,N_2874,N_2789);
nor U3113 (N_3113,N_2532,N_2742);
and U3114 (N_3114,N_2780,N_2793);
nand U3115 (N_3115,N_2604,N_2886);
and U3116 (N_3116,N_2694,N_2931);
nand U3117 (N_3117,N_2611,N_2929);
xor U3118 (N_3118,N_2547,N_2512);
xnor U3119 (N_3119,N_2861,N_2832);
or U3120 (N_3120,N_2514,N_2598);
nor U3121 (N_3121,N_2846,N_2590);
or U3122 (N_3122,N_2503,N_2731);
nor U3123 (N_3123,N_2806,N_2528);
and U3124 (N_3124,N_2847,N_2625);
nor U3125 (N_3125,N_2575,N_2916);
or U3126 (N_3126,N_2600,N_2696);
and U3127 (N_3127,N_2934,N_2553);
nor U3128 (N_3128,N_2502,N_2991);
nand U3129 (N_3129,N_2943,N_2801);
or U3130 (N_3130,N_2739,N_2883);
nor U3131 (N_3131,N_2680,N_2681);
or U3132 (N_3132,N_2552,N_2641);
nor U3133 (N_3133,N_2627,N_2601);
nor U3134 (N_3134,N_2650,N_2636);
nor U3135 (N_3135,N_2985,N_2655);
and U3136 (N_3136,N_2913,N_2921);
and U3137 (N_3137,N_2702,N_2674);
xor U3138 (N_3138,N_2662,N_2633);
nor U3139 (N_3139,N_2882,N_2993);
nor U3140 (N_3140,N_2937,N_2599);
xor U3141 (N_3141,N_2820,N_2628);
or U3142 (N_3142,N_2922,N_2772);
nand U3143 (N_3143,N_2616,N_2958);
nor U3144 (N_3144,N_2888,N_2612);
or U3145 (N_3145,N_2752,N_2548);
and U3146 (N_3146,N_2918,N_2687);
or U3147 (N_3147,N_2871,N_2767);
and U3148 (N_3148,N_2843,N_2558);
nand U3149 (N_3149,N_2756,N_2776);
and U3150 (N_3150,N_2754,N_2839);
nand U3151 (N_3151,N_2522,N_2753);
xnor U3152 (N_3152,N_2946,N_2638);
xnor U3153 (N_3153,N_2562,N_2518);
and U3154 (N_3154,N_2981,N_2725);
nor U3155 (N_3155,N_2607,N_2878);
or U3156 (N_3156,N_2797,N_2524);
nor U3157 (N_3157,N_2541,N_2555);
or U3158 (N_3158,N_2704,N_2782);
nor U3159 (N_3159,N_2798,N_2693);
or U3160 (N_3160,N_2665,N_2907);
or U3161 (N_3161,N_2602,N_2872);
nor U3162 (N_3162,N_2790,N_2973);
nor U3163 (N_3163,N_2768,N_2795);
nand U3164 (N_3164,N_2947,N_2995);
nor U3165 (N_3165,N_2732,N_2523);
nand U3166 (N_3166,N_2763,N_2850);
nor U3167 (N_3167,N_2814,N_2703);
or U3168 (N_3168,N_2988,N_2944);
nor U3169 (N_3169,N_2770,N_2900);
and U3170 (N_3170,N_2534,N_2863);
nand U3171 (N_3171,N_2807,N_2864);
xor U3172 (N_3172,N_2624,N_2557);
or U3173 (N_3173,N_2892,N_2632);
nand U3174 (N_3174,N_2757,N_2730);
nand U3175 (N_3175,N_2715,N_2530);
or U3176 (N_3176,N_2835,N_2783);
and U3177 (N_3177,N_2691,N_2642);
or U3178 (N_3178,N_2837,N_2711);
or U3179 (N_3179,N_2919,N_2826);
or U3180 (N_3180,N_2974,N_2758);
or U3181 (N_3181,N_2728,N_2603);
xnor U3182 (N_3182,N_2781,N_2526);
nand U3183 (N_3183,N_2683,N_2551);
nor U3184 (N_3184,N_2851,N_2761);
and U3185 (N_3185,N_2545,N_2858);
xor U3186 (N_3186,N_2726,N_2970);
and U3187 (N_3187,N_2819,N_2841);
or U3188 (N_3188,N_2933,N_2794);
and U3189 (N_3189,N_2936,N_2656);
nor U3190 (N_3190,N_2893,N_2595);
and U3191 (N_3191,N_2516,N_2903);
and U3192 (N_3192,N_2821,N_2992);
and U3193 (N_3193,N_2500,N_2678);
nand U3194 (N_3194,N_2949,N_2792);
xnor U3195 (N_3195,N_2675,N_2574);
xnor U3196 (N_3196,N_2605,N_2727);
nand U3197 (N_3197,N_2592,N_2724);
nor U3198 (N_3198,N_2568,N_2775);
nand U3199 (N_3199,N_2880,N_2779);
nand U3200 (N_3200,N_2766,N_2842);
xor U3201 (N_3201,N_2701,N_2659);
nor U3202 (N_3202,N_2962,N_2808);
nor U3203 (N_3203,N_2898,N_2559);
nand U3204 (N_3204,N_2622,N_2976);
xnor U3205 (N_3205,N_2987,N_2910);
and U3206 (N_3206,N_2653,N_2736);
nand U3207 (N_3207,N_2799,N_2950);
nand U3208 (N_3208,N_2890,N_2560);
or U3209 (N_3209,N_2956,N_2751);
and U3210 (N_3210,N_2546,N_2891);
nand U3211 (N_3211,N_2774,N_2734);
nor U3212 (N_3212,N_2748,N_2549);
nor U3213 (N_3213,N_2998,N_2738);
or U3214 (N_3214,N_2672,N_2964);
nand U3215 (N_3215,N_2567,N_2796);
or U3216 (N_3216,N_2717,N_2930);
nand U3217 (N_3217,N_2915,N_2838);
and U3218 (N_3218,N_2865,N_2714);
xor U3219 (N_3219,N_2550,N_2965);
xor U3220 (N_3220,N_2668,N_2578);
and U3221 (N_3221,N_2658,N_2829);
and U3222 (N_3222,N_2926,N_2596);
xor U3223 (N_3223,N_2697,N_2507);
xor U3224 (N_3224,N_2834,N_2511);
nand U3225 (N_3225,N_2940,N_2710);
or U3226 (N_3226,N_2620,N_2676);
xnor U3227 (N_3227,N_2623,N_2800);
nor U3228 (N_3228,N_2698,N_2942);
or U3229 (N_3229,N_2573,N_2649);
nor U3230 (N_3230,N_2860,N_2788);
and U3231 (N_3231,N_2852,N_2556);
nor U3232 (N_3232,N_2908,N_2971);
and U3233 (N_3233,N_2840,N_2884);
nor U3234 (N_3234,N_2707,N_2608);
and U3235 (N_3235,N_2640,N_2565);
nand U3236 (N_3236,N_2743,N_2645);
xnor U3237 (N_3237,N_2520,N_2729);
nor U3238 (N_3238,N_2785,N_2531);
or U3239 (N_3239,N_2643,N_2705);
and U3240 (N_3240,N_2741,N_2536);
nand U3241 (N_3241,N_2959,N_2802);
and U3242 (N_3242,N_2660,N_2966);
or U3243 (N_3243,N_2911,N_2830);
nand U3244 (N_3244,N_2646,N_2982);
xnor U3245 (N_3245,N_2804,N_2899);
xor U3246 (N_3246,N_2759,N_2733);
nor U3247 (N_3247,N_2854,N_2745);
and U3248 (N_3248,N_2765,N_2666);
nor U3249 (N_3249,N_2967,N_2543);
xnor U3250 (N_3250,N_2881,N_2912);
and U3251 (N_3251,N_2942,N_2622);
or U3252 (N_3252,N_2856,N_2982);
nor U3253 (N_3253,N_2686,N_2759);
or U3254 (N_3254,N_2839,N_2798);
xor U3255 (N_3255,N_2965,N_2711);
xnor U3256 (N_3256,N_2858,N_2929);
xor U3257 (N_3257,N_2936,N_2741);
xnor U3258 (N_3258,N_2829,N_2999);
nand U3259 (N_3259,N_2693,N_2720);
nand U3260 (N_3260,N_2751,N_2671);
or U3261 (N_3261,N_2748,N_2657);
or U3262 (N_3262,N_2832,N_2843);
xnor U3263 (N_3263,N_2799,N_2930);
nor U3264 (N_3264,N_2987,N_2588);
nor U3265 (N_3265,N_2721,N_2646);
and U3266 (N_3266,N_2656,N_2734);
and U3267 (N_3267,N_2701,N_2520);
xnor U3268 (N_3268,N_2958,N_2528);
nand U3269 (N_3269,N_2864,N_2924);
and U3270 (N_3270,N_2855,N_2952);
or U3271 (N_3271,N_2502,N_2840);
nand U3272 (N_3272,N_2978,N_2688);
xor U3273 (N_3273,N_2673,N_2528);
nor U3274 (N_3274,N_2978,N_2679);
or U3275 (N_3275,N_2670,N_2864);
nand U3276 (N_3276,N_2829,N_2883);
nand U3277 (N_3277,N_2737,N_2957);
or U3278 (N_3278,N_2852,N_2934);
or U3279 (N_3279,N_2765,N_2726);
nand U3280 (N_3280,N_2973,N_2817);
xor U3281 (N_3281,N_2743,N_2589);
xor U3282 (N_3282,N_2880,N_2968);
and U3283 (N_3283,N_2984,N_2532);
and U3284 (N_3284,N_2860,N_2705);
nand U3285 (N_3285,N_2984,N_2793);
xnor U3286 (N_3286,N_2660,N_2851);
or U3287 (N_3287,N_2703,N_2524);
xnor U3288 (N_3288,N_2816,N_2696);
nand U3289 (N_3289,N_2901,N_2503);
and U3290 (N_3290,N_2620,N_2695);
nor U3291 (N_3291,N_2559,N_2783);
or U3292 (N_3292,N_2544,N_2626);
and U3293 (N_3293,N_2849,N_2791);
nand U3294 (N_3294,N_2702,N_2983);
and U3295 (N_3295,N_2880,N_2751);
nor U3296 (N_3296,N_2783,N_2794);
nor U3297 (N_3297,N_2793,N_2553);
xnor U3298 (N_3298,N_2918,N_2581);
nor U3299 (N_3299,N_2614,N_2505);
or U3300 (N_3300,N_2756,N_2608);
nand U3301 (N_3301,N_2733,N_2650);
nor U3302 (N_3302,N_2608,N_2745);
nand U3303 (N_3303,N_2530,N_2881);
nor U3304 (N_3304,N_2979,N_2705);
xor U3305 (N_3305,N_2512,N_2831);
nand U3306 (N_3306,N_2863,N_2884);
and U3307 (N_3307,N_2893,N_2671);
or U3308 (N_3308,N_2527,N_2821);
or U3309 (N_3309,N_2852,N_2808);
and U3310 (N_3310,N_2830,N_2642);
or U3311 (N_3311,N_2964,N_2696);
or U3312 (N_3312,N_2762,N_2515);
nand U3313 (N_3313,N_2964,N_2687);
and U3314 (N_3314,N_2720,N_2669);
or U3315 (N_3315,N_2513,N_2606);
nand U3316 (N_3316,N_2680,N_2656);
xor U3317 (N_3317,N_2893,N_2694);
nand U3318 (N_3318,N_2900,N_2767);
nand U3319 (N_3319,N_2940,N_2758);
or U3320 (N_3320,N_2667,N_2883);
nand U3321 (N_3321,N_2975,N_2912);
nand U3322 (N_3322,N_2773,N_2878);
xnor U3323 (N_3323,N_2560,N_2824);
and U3324 (N_3324,N_2688,N_2758);
nand U3325 (N_3325,N_2804,N_2947);
xnor U3326 (N_3326,N_2870,N_2602);
and U3327 (N_3327,N_2759,N_2711);
xor U3328 (N_3328,N_2703,N_2859);
nand U3329 (N_3329,N_2992,N_2746);
or U3330 (N_3330,N_2644,N_2855);
xnor U3331 (N_3331,N_2615,N_2763);
xnor U3332 (N_3332,N_2885,N_2711);
nand U3333 (N_3333,N_2646,N_2513);
and U3334 (N_3334,N_2995,N_2966);
and U3335 (N_3335,N_2549,N_2928);
xor U3336 (N_3336,N_2967,N_2718);
xor U3337 (N_3337,N_2526,N_2626);
and U3338 (N_3338,N_2575,N_2858);
and U3339 (N_3339,N_2939,N_2611);
and U3340 (N_3340,N_2972,N_2888);
nor U3341 (N_3341,N_2609,N_2779);
or U3342 (N_3342,N_2522,N_2660);
nand U3343 (N_3343,N_2742,N_2810);
xnor U3344 (N_3344,N_2713,N_2930);
or U3345 (N_3345,N_2892,N_2765);
or U3346 (N_3346,N_2949,N_2576);
nand U3347 (N_3347,N_2632,N_2960);
nor U3348 (N_3348,N_2824,N_2795);
xor U3349 (N_3349,N_2721,N_2590);
xnor U3350 (N_3350,N_2807,N_2652);
xnor U3351 (N_3351,N_2745,N_2819);
xor U3352 (N_3352,N_2562,N_2567);
nand U3353 (N_3353,N_2585,N_2947);
nand U3354 (N_3354,N_2601,N_2894);
nand U3355 (N_3355,N_2539,N_2873);
xor U3356 (N_3356,N_2697,N_2709);
xnor U3357 (N_3357,N_2741,N_2579);
or U3358 (N_3358,N_2927,N_2668);
and U3359 (N_3359,N_2728,N_2897);
nor U3360 (N_3360,N_2778,N_2756);
or U3361 (N_3361,N_2532,N_2773);
nor U3362 (N_3362,N_2939,N_2938);
or U3363 (N_3363,N_2781,N_2641);
and U3364 (N_3364,N_2807,N_2632);
or U3365 (N_3365,N_2922,N_2809);
nand U3366 (N_3366,N_2694,N_2912);
or U3367 (N_3367,N_2703,N_2760);
and U3368 (N_3368,N_2719,N_2554);
or U3369 (N_3369,N_2615,N_2891);
nor U3370 (N_3370,N_2903,N_2944);
xnor U3371 (N_3371,N_2716,N_2683);
nand U3372 (N_3372,N_2666,N_2576);
or U3373 (N_3373,N_2975,N_2594);
nand U3374 (N_3374,N_2862,N_2533);
nand U3375 (N_3375,N_2561,N_2815);
xnor U3376 (N_3376,N_2665,N_2566);
nand U3377 (N_3377,N_2938,N_2637);
xor U3378 (N_3378,N_2833,N_2778);
nor U3379 (N_3379,N_2741,N_2642);
xor U3380 (N_3380,N_2702,N_2909);
or U3381 (N_3381,N_2657,N_2602);
nand U3382 (N_3382,N_2873,N_2890);
or U3383 (N_3383,N_2755,N_2861);
and U3384 (N_3384,N_2846,N_2750);
or U3385 (N_3385,N_2516,N_2520);
nor U3386 (N_3386,N_2637,N_2750);
or U3387 (N_3387,N_2877,N_2595);
xor U3388 (N_3388,N_2788,N_2867);
nor U3389 (N_3389,N_2730,N_2752);
or U3390 (N_3390,N_2546,N_2746);
nand U3391 (N_3391,N_2966,N_2659);
and U3392 (N_3392,N_2991,N_2550);
or U3393 (N_3393,N_2543,N_2775);
nor U3394 (N_3394,N_2831,N_2631);
nor U3395 (N_3395,N_2895,N_2573);
or U3396 (N_3396,N_2669,N_2525);
nand U3397 (N_3397,N_2568,N_2841);
or U3398 (N_3398,N_2861,N_2984);
nor U3399 (N_3399,N_2665,N_2599);
or U3400 (N_3400,N_2584,N_2788);
nor U3401 (N_3401,N_2814,N_2554);
and U3402 (N_3402,N_2960,N_2929);
or U3403 (N_3403,N_2662,N_2664);
nor U3404 (N_3404,N_2975,N_2897);
and U3405 (N_3405,N_2545,N_2693);
nor U3406 (N_3406,N_2823,N_2621);
nand U3407 (N_3407,N_2786,N_2695);
or U3408 (N_3408,N_2973,N_2560);
xor U3409 (N_3409,N_2711,N_2523);
nand U3410 (N_3410,N_2673,N_2871);
xnor U3411 (N_3411,N_2920,N_2976);
nor U3412 (N_3412,N_2772,N_2965);
nor U3413 (N_3413,N_2925,N_2502);
or U3414 (N_3414,N_2726,N_2727);
and U3415 (N_3415,N_2736,N_2728);
nor U3416 (N_3416,N_2719,N_2629);
or U3417 (N_3417,N_2521,N_2941);
and U3418 (N_3418,N_2776,N_2556);
nand U3419 (N_3419,N_2916,N_2808);
nand U3420 (N_3420,N_2868,N_2725);
and U3421 (N_3421,N_2550,N_2984);
xnor U3422 (N_3422,N_2835,N_2992);
and U3423 (N_3423,N_2961,N_2997);
nand U3424 (N_3424,N_2842,N_2506);
nor U3425 (N_3425,N_2990,N_2882);
and U3426 (N_3426,N_2916,N_2680);
nand U3427 (N_3427,N_2535,N_2826);
xor U3428 (N_3428,N_2655,N_2970);
and U3429 (N_3429,N_2729,N_2944);
and U3430 (N_3430,N_2987,N_2564);
nor U3431 (N_3431,N_2585,N_2818);
nor U3432 (N_3432,N_2664,N_2640);
nor U3433 (N_3433,N_2678,N_2773);
nor U3434 (N_3434,N_2720,N_2853);
and U3435 (N_3435,N_2925,N_2987);
and U3436 (N_3436,N_2822,N_2543);
or U3437 (N_3437,N_2938,N_2879);
xor U3438 (N_3438,N_2689,N_2880);
nand U3439 (N_3439,N_2621,N_2563);
nor U3440 (N_3440,N_2886,N_2768);
and U3441 (N_3441,N_2898,N_2804);
or U3442 (N_3442,N_2713,N_2878);
or U3443 (N_3443,N_2910,N_2772);
and U3444 (N_3444,N_2672,N_2690);
and U3445 (N_3445,N_2691,N_2924);
and U3446 (N_3446,N_2589,N_2935);
nor U3447 (N_3447,N_2908,N_2848);
nand U3448 (N_3448,N_2948,N_2501);
nor U3449 (N_3449,N_2683,N_2728);
and U3450 (N_3450,N_2705,N_2745);
and U3451 (N_3451,N_2761,N_2602);
xnor U3452 (N_3452,N_2699,N_2891);
nor U3453 (N_3453,N_2773,N_2798);
xnor U3454 (N_3454,N_2958,N_2719);
and U3455 (N_3455,N_2691,N_2751);
xor U3456 (N_3456,N_2988,N_2967);
nor U3457 (N_3457,N_2513,N_2775);
xnor U3458 (N_3458,N_2657,N_2513);
or U3459 (N_3459,N_2967,N_2550);
nor U3460 (N_3460,N_2586,N_2569);
nand U3461 (N_3461,N_2528,N_2816);
or U3462 (N_3462,N_2894,N_2914);
nand U3463 (N_3463,N_2738,N_2844);
nor U3464 (N_3464,N_2943,N_2771);
nand U3465 (N_3465,N_2941,N_2799);
nor U3466 (N_3466,N_2722,N_2990);
nor U3467 (N_3467,N_2965,N_2960);
or U3468 (N_3468,N_2864,N_2630);
and U3469 (N_3469,N_2650,N_2868);
xnor U3470 (N_3470,N_2894,N_2550);
xor U3471 (N_3471,N_2959,N_2836);
nor U3472 (N_3472,N_2638,N_2948);
nand U3473 (N_3473,N_2540,N_2914);
xor U3474 (N_3474,N_2923,N_2655);
or U3475 (N_3475,N_2728,N_2922);
nor U3476 (N_3476,N_2800,N_2780);
nor U3477 (N_3477,N_2887,N_2610);
or U3478 (N_3478,N_2893,N_2736);
nand U3479 (N_3479,N_2500,N_2877);
nand U3480 (N_3480,N_2710,N_2578);
or U3481 (N_3481,N_2734,N_2906);
or U3482 (N_3482,N_2784,N_2986);
nor U3483 (N_3483,N_2523,N_2504);
xor U3484 (N_3484,N_2939,N_2553);
xnor U3485 (N_3485,N_2633,N_2720);
nor U3486 (N_3486,N_2969,N_2562);
and U3487 (N_3487,N_2818,N_2537);
or U3488 (N_3488,N_2622,N_2710);
and U3489 (N_3489,N_2666,N_2709);
or U3490 (N_3490,N_2899,N_2991);
or U3491 (N_3491,N_2957,N_2554);
or U3492 (N_3492,N_2996,N_2863);
nand U3493 (N_3493,N_2888,N_2571);
and U3494 (N_3494,N_2629,N_2635);
nand U3495 (N_3495,N_2875,N_2513);
xor U3496 (N_3496,N_2557,N_2626);
or U3497 (N_3497,N_2515,N_2514);
xnor U3498 (N_3498,N_2963,N_2687);
or U3499 (N_3499,N_2621,N_2879);
xor U3500 (N_3500,N_3034,N_3371);
nand U3501 (N_3501,N_3282,N_3068);
nand U3502 (N_3502,N_3144,N_3043);
or U3503 (N_3503,N_3079,N_3214);
nand U3504 (N_3504,N_3202,N_3404);
xnor U3505 (N_3505,N_3486,N_3397);
nor U3506 (N_3506,N_3220,N_3284);
and U3507 (N_3507,N_3415,N_3374);
nand U3508 (N_3508,N_3273,N_3003);
nand U3509 (N_3509,N_3064,N_3010);
nand U3510 (N_3510,N_3170,N_3025);
or U3511 (N_3511,N_3382,N_3014);
or U3512 (N_3512,N_3210,N_3426);
nand U3513 (N_3513,N_3256,N_3248);
and U3514 (N_3514,N_3205,N_3150);
xor U3515 (N_3515,N_3028,N_3037);
and U3516 (N_3516,N_3357,N_3339);
nand U3517 (N_3517,N_3254,N_3431);
and U3518 (N_3518,N_3302,N_3436);
nor U3519 (N_3519,N_3148,N_3005);
nand U3520 (N_3520,N_3443,N_3208);
nand U3521 (N_3521,N_3149,N_3095);
and U3522 (N_3522,N_3153,N_3324);
or U3523 (N_3523,N_3027,N_3224);
nor U3524 (N_3524,N_3447,N_3097);
and U3525 (N_3525,N_3345,N_3231);
or U3526 (N_3526,N_3127,N_3306);
nand U3527 (N_3527,N_3269,N_3152);
xnor U3528 (N_3528,N_3381,N_3230);
xor U3529 (N_3529,N_3408,N_3213);
nand U3530 (N_3530,N_3219,N_3067);
nand U3531 (N_3531,N_3180,N_3232);
or U3532 (N_3532,N_3416,N_3178);
xnor U3533 (N_3533,N_3480,N_3305);
nand U3534 (N_3534,N_3174,N_3477);
nand U3535 (N_3535,N_3196,N_3048);
xnor U3536 (N_3536,N_3359,N_3352);
xnor U3537 (N_3537,N_3234,N_3419);
xnor U3538 (N_3538,N_3361,N_3376);
or U3539 (N_3539,N_3267,N_3473);
nor U3540 (N_3540,N_3207,N_3309);
nand U3541 (N_3541,N_3294,N_3026);
or U3542 (N_3542,N_3100,N_3463);
and U3543 (N_3543,N_3413,N_3314);
and U3544 (N_3544,N_3369,N_3467);
and U3545 (N_3545,N_3159,N_3368);
nor U3546 (N_3546,N_3074,N_3249);
xor U3547 (N_3547,N_3176,N_3323);
nand U3548 (N_3548,N_3112,N_3494);
and U3549 (N_3549,N_3041,N_3163);
or U3550 (N_3550,N_3192,N_3199);
xnor U3551 (N_3551,N_3098,N_3030);
nand U3552 (N_3552,N_3360,N_3434);
nor U3553 (N_3553,N_3177,N_3185);
xor U3554 (N_3554,N_3440,N_3243);
xor U3555 (N_3555,N_3222,N_3304);
nand U3556 (N_3556,N_3044,N_3307);
or U3557 (N_3557,N_3425,N_3084);
nor U3558 (N_3558,N_3375,N_3221);
nand U3559 (N_3559,N_3091,N_3492);
or U3560 (N_3560,N_3365,N_3218);
or U3561 (N_3561,N_3423,N_3029);
xor U3562 (N_3562,N_3216,N_3490);
and U3563 (N_3563,N_3090,N_3120);
or U3564 (N_3564,N_3479,N_3040);
nor U3565 (N_3565,N_3464,N_3105);
xnor U3566 (N_3566,N_3481,N_3461);
xor U3567 (N_3567,N_3452,N_3087);
and U3568 (N_3568,N_3146,N_3069);
or U3569 (N_3569,N_3118,N_3388);
nand U3570 (N_3570,N_3266,N_3108);
nor U3571 (N_3571,N_3056,N_3168);
nor U3572 (N_3572,N_3175,N_3343);
or U3573 (N_3573,N_3387,N_3096);
and U3574 (N_3574,N_3126,N_3311);
or U3575 (N_3575,N_3061,N_3189);
xnor U3576 (N_3576,N_3341,N_3295);
and U3577 (N_3577,N_3468,N_3407);
nor U3578 (N_3578,N_3383,N_3313);
nand U3579 (N_3579,N_3346,N_3366);
nor U3580 (N_3580,N_3349,N_3156);
xor U3581 (N_3581,N_3227,N_3332);
or U3582 (N_3582,N_3330,N_3271);
nor U3583 (N_3583,N_3086,N_3342);
nand U3584 (N_3584,N_3083,N_3225);
nand U3585 (N_3585,N_3115,N_3035);
nand U3586 (N_3586,N_3011,N_3402);
or U3587 (N_3587,N_3223,N_3103);
nand U3588 (N_3588,N_3296,N_3364);
nor U3589 (N_3589,N_3321,N_3181);
and U3590 (N_3590,N_3372,N_3395);
and U3591 (N_3591,N_3102,N_3050);
and U3592 (N_3592,N_3021,N_3328);
nand U3593 (N_3593,N_3261,N_3299);
xnor U3594 (N_3594,N_3475,N_3006);
and U3595 (N_3595,N_3493,N_3457);
and U3596 (N_3596,N_3308,N_3370);
nand U3597 (N_3597,N_3496,N_3128);
and U3598 (N_3598,N_3356,N_3155);
nand U3599 (N_3599,N_3393,N_3456);
nor U3600 (N_3600,N_3184,N_3052);
nand U3601 (N_3601,N_3277,N_3186);
nor U3602 (N_3602,N_3065,N_3054);
or U3603 (N_3603,N_3350,N_3092);
xor U3604 (N_3604,N_3430,N_3264);
xnor U3605 (N_3605,N_3421,N_3179);
and U3606 (N_3606,N_3099,N_3335);
nand U3607 (N_3607,N_3110,N_3472);
nand U3608 (N_3608,N_3448,N_3228);
and U3609 (N_3609,N_3020,N_3193);
and U3610 (N_3610,N_3190,N_3251);
xor U3611 (N_3611,N_3437,N_3428);
nor U3612 (N_3612,N_3089,N_3203);
or U3613 (N_3613,N_3257,N_3031);
nand U3614 (N_3614,N_3046,N_3077);
nand U3615 (N_3615,N_3215,N_3138);
and U3616 (N_3616,N_3134,N_3389);
nor U3617 (N_3617,N_3255,N_3013);
and U3618 (N_3618,N_3182,N_3039);
and U3619 (N_3619,N_3301,N_3390);
and U3620 (N_3620,N_3094,N_3060);
nand U3621 (N_3621,N_3075,N_3137);
xnor U3622 (N_3622,N_3334,N_3133);
nor U3623 (N_3623,N_3131,N_3080);
or U3624 (N_3624,N_3462,N_3062);
xnor U3625 (N_3625,N_3449,N_3143);
nand U3626 (N_3626,N_3002,N_3378);
xnor U3627 (N_3627,N_3226,N_3275);
or U3628 (N_3628,N_3337,N_3063);
xnor U3629 (N_3629,N_3183,N_3398);
nand U3630 (N_3630,N_3057,N_3400);
nor U3631 (N_3631,N_3454,N_3088);
or U3632 (N_3632,N_3451,N_3288);
or U3633 (N_3633,N_3344,N_3217);
xnor U3634 (N_3634,N_3188,N_3459);
nand U3635 (N_3635,N_3290,N_3147);
xor U3636 (N_3636,N_3141,N_3032);
xor U3637 (N_3637,N_3292,N_3247);
nor U3638 (N_3638,N_3410,N_3236);
nand U3639 (N_3639,N_3023,N_3384);
and U3640 (N_3640,N_3417,N_3489);
nor U3641 (N_3641,N_3004,N_3445);
nor U3642 (N_3642,N_3315,N_3268);
and U3643 (N_3643,N_3386,N_3319);
nor U3644 (N_3644,N_3379,N_3326);
nor U3645 (N_3645,N_3081,N_3173);
or U3646 (N_3646,N_3336,N_3474);
nor U3647 (N_3647,N_3139,N_3238);
nor U3648 (N_3648,N_3113,N_3209);
and U3649 (N_3649,N_3198,N_3291);
nor U3650 (N_3650,N_3272,N_3201);
xor U3651 (N_3651,N_3485,N_3409);
nor U3652 (N_3652,N_3085,N_3258);
nor U3653 (N_3653,N_3466,N_3123);
or U3654 (N_3654,N_3399,N_3385);
nor U3655 (N_3655,N_3197,N_3045);
xor U3656 (N_3656,N_3121,N_3212);
xor U3657 (N_3657,N_3073,N_3262);
nor U3658 (N_3658,N_3403,N_3495);
or U3659 (N_3659,N_3154,N_3047);
and U3660 (N_3660,N_3450,N_3289);
xnor U3661 (N_3661,N_3422,N_3394);
nor U3662 (N_3662,N_3022,N_3242);
nor U3663 (N_3663,N_3009,N_3066);
xnor U3664 (N_3664,N_3132,N_3469);
nor U3665 (N_3665,N_3312,N_3274);
nor U3666 (N_3666,N_3114,N_3235);
and U3667 (N_3667,N_3245,N_3460);
nand U3668 (N_3668,N_3008,N_3482);
and U3669 (N_3669,N_3125,N_3101);
xnor U3670 (N_3670,N_3396,N_3206);
and U3671 (N_3671,N_3465,N_3444);
nand U3672 (N_3672,N_3318,N_3418);
nor U3673 (N_3673,N_3018,N_3007);
nand U3674 (N_3674,N_3191,N_3298);
or U3675 (N_3675,N_3015,N_3263);
nor U3676 (N_3676,N_3325,N_3338);
nand U3677 (N_3677,N_3082,N_3406);
or U3678 (N_3678,N_3001,N_3107);
nor U3679 (N_3679,N_3195,N_3078);
and U3680 (N_3680,N_3405,N_3471);
nand U3681 (N_3681,N_3283,N_3265);
or U3682 (N_3682,N_3252,N_3194);
xor U3683 (N_3683,N_3362,N_3287);
nand U3684 (N_3684,N_3438,N_3348);
and U3685 (N_3685,N_3420,N_3233);
nand U3686 (N_3686,N_3303,N_3355);
nor U3687 (N_3687,N_3051,N_3033);
or U3688 (N_3688,N_3498,N_3487);
nor U3689 (N_3689,N_3017,N_3171);
xnor U3690 (N_3690,N_3130,N_3049);
and U3691 (N_3691,N_3476,N_3012);
nand U3692 (N_3692,N_3237,N_3162);
or U3693 (N_3693,N_3104,N_3161);
or U3694 (N_3694,N_3122,N_3000);
and U3695 (N_3695,N_3327,N_3165);
or U3696 (N_3696,N_3446,N_3135);
xor U3697 (N_3697,N_3320,N_3453);
nor U3698 (N_3698,N_3412,N_3211);
nor U3699 (N_3699,N_3317,N_3331);
nor U3700 (N_3700,N_3136,N_3145);
nand U3701 (N_3701,N_3484,N_3363);
xnor U3702 (N_3702,N_3276,N_3491);
nand U3703 (N_3703,N_3260,N_3093);
xor U3704 (N_3704,N_3076,N_3160);
nor U3705 (N_3705,N_3240,N_3333);
xor U3706 (N_3706,N_3322,N_3310);
nor U3707 (N_3707,N_3300,N_3172);
and U3708 (N_3708,N_3455,N_3429);
xnor U3709 (N_3709,N_3111,N_3164);
xnor U3710 (N_3710,N_3187,N_3059);
xor U3711 (N_3711,N_3109,N_3279);
xor U3712 (N_3712,N_3241,N_3024);
xor U3713 (N_3713,N_3433,N_3392);
nor U3714 (N_3714,N_3278,N_3071);
nor U3715 (N_3715,N_3497,N_3347);
and U3716 (N_3716,N_3070,N_3016);
nor U3717 (N_3717,N_3157,N_3129);
or U3718 (N_3718,N_3377,N_3142);
or U3719 (N_3719,N_3250,N_3058);
or U3720 (N_3720,N_3036,N_3411);
or U3721 (N_3721,N_3151,N_3353);
or U3722 (N_3722,N_3285,N_3286);
and U3723 (N_3723,N_3380,N_3204);
xor U3724 (N_3724,N_3166,N_3038);
or U3725 (N_3725,N_3119,N_3358);
or U3726 (N_3726,N_3414,N_3293);
and U3727 (N_3727,N_3458,N_3354);
nor U3728 (N_3728,N_3200,N_3167);
nand U3729 (N_3729,N_3072,N_3391);
xor U3730 (N_3730,N_3483,N_3229);
xor U3731 (N_3731,N_3280,N_3427);
xor U3732 (N_3732,N_3470,N_3106);
nand U3733 (N_3733,N_3042,N_3401);
xor U3734 (N_3734,N_3246,N_3441);
and U3735 (N_3735,N_3439,N_3329);
or U3736 (N_3736,N_3340,N_3158);
and U3737 (N_3737,N_3117,N_3297);
xnor U3738 (N_3738,N_3281,N_3019);
or U3739 (N_3739,N_3499,N_3488);
xnor U3740 (N_3740,N_3270,N_3253);
nor U3741 (N_3741,N_3351,N_3244);
nand U3742 (N_3742,N_3367,N_3239);
nor U3743 (N_3743,N_3053,N_3140);
xor U3744 (N_3744,N_3424,N_3442);
nand U3745 (N_3745,N_3432,N_3116);
and U3746 (N_3746,N_3124,N_3316);
nand U3747 (N_3747,N_3259,N_3435);
and U3748 (N_3748,N_3373,N_3055);
and U3749 (N_3749,N_3169,N_3478);
nor U3750 (N_3750,N_3207,N_3452);
and U3751 (N_3751,N_3455,N_3018);
and U3752 (N_3752,N_3437,N_3467);
xnor U3753 (N_3753,N_3202,N_3088);
and U3754 (N_3754,N_3118,N_3285);
or U3755 (N_3755,N_3029,N_3449);
or U3756 (N_3756,N_3227,N_3180);
nor U3757 (N_3757,N_3198,N_3466);
xor U3758 (N_3758,N_3457,N_3109);
or U3759 (N_3759,N_3115,N_3269);
nor U3760 (N_3760,N_3381,N_3353);
nor U3761 (N_3761,N_3396,N_3093);
and U3762 (N_3762,N_3077,N_3389);
nor U3763 (N_3763,N_3406,N_3346);
nor U3764 (N_3764,N_3396,N_3131);
and U3765 (N_3765,N_3229,N_3478);
xor U3766 (N_3766,N_3266,N_3458);
nand U3767 (N_3767,N_3095,N_3168);
nor U3768 (N_3768,N_3416,N_3204);
nor U3769 (N_3769,N_3201,N_3181);
nor U3770 (N_3770,N_3210,N_3438);
xnor U3771 (N_3771,N_3470,N_3480);
nor U3772 (N_3772,N_3159,N_3090);
or U3773 (N_3773,N_3422,N_3078);
or U3774 (N_3774,N_3343,N_3019);
and U3775 (N_3775,N_3091,N_3261);
nor U3776 (N_3776,N_3331,N_3293);
and U3777 (N_3777,N_3082,N_3456);
nand U3778 (N_3778,N_3349,N_3341);
and U3779 (N_3779,N_3374,N_3285);
xor U3780 (N_3780,N_3095,N_3468);
nand U3781 (N_3781,N_3216,N_3289);
or U3782 (N_3782,N_3007,N_3379);
and U3783 (N_3783,N_3353,N_3138);
nand U3784 (N_3784,N_3223,N_3098);
xor U3785 (N_3785,N_3098,N_3264);
nor U3786 (N_3786,N_3267,N_3182);
and U3787 (N_3787,N_3005,N_3020);
nand U3788 (N_3788,N_3071,N_3444);
and U3789 (N_3789,N_3323,N_3124);
nor U3790 (N_3790,N_3337,N_3077);
or U3791 (N_3791,N_3158,N_3089);
nor U3792 (N_3792,N_3255,N_3155);
nand U3793 (N_3793,N_3438,N_3439);
and U3794 (N_3794,N_3360,N_3123);
or U3795 (N_3795,N_3068,N_3088);
xnor U3796 (N_3796,N_3252,N_3468);
or U3797 (N_3797,N_3105,N_3051);
nor U3798 (N_3798,N_3495,N_3198);
nor U3799 (N_3799,N_3271,N_3054);
xnor U3800 (N_3800,N_3235,N_3241);
or U3801 (N_3801,N_3334,N_3115);
and U3802 (N_3802,N_3041,N_3358);
and U3803 (N_3803,N_3163,N_3264);
and U3804 (N_3804,N_3443,N_3117);
or U3805 (N_3805,N_3030,N_3137);
xnor U3806 (N_3806,N_3169,N_3331);
and U3807 (N_3807,N_3428,N_3017);
xor U3808 (N_3808,N_3213,N_3173);
nor U3809 (N_3809,N_3459,N_3386);
nor U3810 (N_3810,N_3109,N_3104);
nand U3811 (N_3811,N_3150,N_3024);
and U3812 (N_3812,N_3017,N_3307);
nand U3813 (N_3813,N_3400,N_3024);
or U3814 (N_3814,N_3455,N_3350);
or U3815 (N_3815,N_3350,N_3353);
nand U3816 (N_3816,N_3310,N_3171);
nor U3817 (N_3817,N_3008,N_3179);
nor U3818 (N_3818,N_3331,N_3205);
nor U3819 (N_3819,N_3094,N_3010);
nor U3820 (N_3820,N_3069,N_3473);
xor U3821 (N_3821,N_3488,N_3486);
nand U3822 (N_3822,N_3433,N_3366);
nor U3823 (N_3823,N_3179,N_3395);
xor U3824 (N_3824,N_3010,N_3430);
and U3825 (N_3825,N_3085,N_3374);
or U3826 (N_3826,N_3208,N_3440);
and U3827 (N_3827,N_3369,N_3435);
and U3828 (N_3828,N_3040,N_3170);
nor U3829 (N_3829,N_3451,N_3427);
nor U3830 (N_3830,N_3342,N_3393);
xor U3831 (N_3831,N_3379,N_3071);
nand U3832 (N_3832,N_3134,N_3077);
or U3833 (N_3833,N_3256,N_3427);
or U3834 (N_3834,N_3154,N_3477);
nor U3835 (N_3835,N_3137,N_3001);
xor U3836 (N_3836,N_3413,N_3391);
and U3837 (N_3837,N_3295,N_3214);
and U3838 (N_3838,N_3081,N_3271);
nor U3839 (N_3839,N_3014,N_3092);
xnor U3840 (N_3840,N_3209,N_3026);
xor U3841 (N_3841,N_3344,N_3459);
xor U3842 (N_3842,N_3353,N_3265);
and U3843 (N_3843,N_3322,N_3425);
nor U3844 (N_3844,N_3398,N_3181);
nand U3845 (N_3845,N_3314,N_3166);
and U3846 (N_3846,N_3377,N_3417);
nor U3847 (N_3847,N_3005,N_3188);
xnor U3848 (N_3848,N_3048,N_3119);
and U3849 (N_3849,N_3449,N_3425);
nor U3850 (N_3850,N_3499,N_3018);
and U3851 (N_3851,N_3392,N_3469);
nand U3852 (N_3852,N_3495,N_3366);
or U3853 (N_3853,N_3357,N_3048);
xor U3854 (N_3854,N_3211,N_3108);
xnor U3855 (N_3855,N_3403,N_3325);
nor U3856 (N_3856,N_3159,N_3234);
nand U3857 (N_3857,N_3058,N_3331);
or U3858 (N_3858,N_3440,N_3078);
or U3859 (N_3859,N_3065,N_3157);
nor U3860 (N_3860,N_3334,N_3341);
xnor U3861 (N_3861,N_3110,N_3264);
and U3862 (N_3862,N_3304,N_3168);
and U3863 (N_3863,N_3247,N_3291);
and U3864 (N_3864,N_3371,N_3125);
nand U3865 (N_3865,N_3444,N_3461);
and U3866 (N_3866,N_3308,N_3432);
nor U3867 (N_3867,N_3219,N_3253);
or U3868 (N_3868,N_3378,N_3478);
and U3869 (N_3869,N_3259,N_3075);
nor U3870 (N_3870,N_3011,N_3260);
nand U3871 (N_3871,N_3026,N_3312);
xnor U3872 (N_3872,N_3315,N_3242);
or U3873 (N_3873,N_3064,N_3244);
nand U3874 (N_3874,N_3081,N_3042);
xor U3875 (N_3875,N_3471,N_3489);
nor U3876 (N_3876,N_3294,N_3065);
or U3877 (N_3877,N_3470,N_3051);
nor U3878 (N_3878,N_3360,N_3400);
or U3879 (N_3879,N_3202,N_3208);
nand U3880 (N_3880,N_3311,N_3323);
nor U3881 (N_3881,N_3373,N_3380);
nand U3882 (N_3882,N_3265,N_3259);
nor U3883 (N_3883,N_3310,N_3144);
nand U3884 (N_3884,N_3400,N_3303);
nor U3885 (N_3885,N_3273,N_3209);
or U3886 (N_3886,N_3294,N_3265);
nand U3887 (N_3887,N_3182,N_3103);
xnor U3888 (N_3888,N_3094,N_3281);
xor U3889 (N_3889,N_3144,N_3309);
or U3890 (N_3890,N_3381,N_3181);
nor U3891 (N_3891,N_3206,N_3033);
xnor U3892 (N_3892,N_3382,N_3142);
xnor U3893 (N_3893,N_3165,N_3388);
or U3894 (N_3894,N_3167,N_3202);
and U3895 (N_3895,N_3001,N_3380);
xnor U3896 (N_3896,N_3107,N_3000);
and U3897 (N_3897,N_3460,N_3226);
and U3898 (N_3898,N_3493,N_3236);
nand U3899 (N_3899,N_3211,N_3057);
nor U3900 (N_3900,N_3294,N_3253);
nor U3901 (N_3901,N_3144,N_3441);
and U3902 (N_3902,N_3168,N_3389);
or U3903 (N_3903,N_3050,N_3079);
xor U3904 (N_3904,N_3002,N_3017);
xnor U3905 (N_3905,N_3197,N_3357);
and U3906 (N_3906,N_3207,N_3110);
xnor U3907 (N_3907,N_3409,N_3252);
and U3908 (N_3908,N_3414,N_3291);
nor U3909 (N_3909,N_3300,N_3074);
or U3910 (N_3910,N_3118,N_3441);
and U3911 (N_3911,N_3460,N_3203);
nand U3912 (N_3912,N_3156,N_3025);
and U3913 (N_3913,N_3495,N_3011);
nand U3914 (N_3914,N_3172,N_3128);
and U3915 (N_3915,N_3425,N_3022);
nand U3916 (N_3916,N_3160,N_3091);
nor U3917 (N_3917,N_3014,N_3459);
xnor U3918 (N_3918,N_3110,N_3391);
and U3919 (N_3919,N_3158,N_3277);
nor U3920 (N_3920,N_3074,N_3220);
nor U3921 (N_3921,N_3468,N_3361);
nor U3922 (N_3922,N_3451,N_3093);
or U3923 (N_3923,N_3183,N_3361);
nor U3924 (N_3924,N_3145,N_3339);
and U3925 (N_3925,N_3402,N_3057);
nor U3926 (N_3926,N_3281,N_3343);
xnor U3927 (N_3927,N_3067,N_3497);
and U3928 (N_3928,N_3275,N_3175);
and U3929 (N_3929,N_3126,N_3049);
xor U3930 (N_3930,N_3498,N_3380);
xnor U3931 (N_3931,N_3333,N_3353);
nor U3932 (N_3932,N_3285,N_3346);
or U3933 (N_3933,N_3244,N_3160);
and U3934 (N_3934,N_3227,N_3222);
and U3935 (N_3935,N_3108,N_3341);
and U3936 (N_3936,N_3364,N_3058);
or U3937 (N_3937,N_3318,N_3097);
xnor U3938 (N_3938,N_3252,N_3202);
nor U3939 (N_3939,N_3052,N_3253);
nand U3940 (N_3940,N_3443,N_3446);
nor U3941 (N_3941,N_3128,N_3402);
nor U3942 (N_3942,N_3352,N_3223);
nand U3943 (N_3943,N_3052,N_3112);
and U3944 (N_3944,N_3352,N_3253);
nand U3945 (N_3945,N_3119,N_3153);
or U3946 (N_3946,N_3277,N_3403);
nand U3947 (N_3947,N_3020,N_3173);
and U3948 (N_3948,N_3300,N_3224);
nor U3949 (N_3949,N_3455,N_3491);
and U3950 (N_3950,N_3281,N_3438);
or U3951 (N_3951,N_3331,N_3424);
nor U3952 (N_3952,N_3247,N_3325);
nand U3953 (N_3953,N_3294,N_3176);
nand U3954 (N_3954,N_3340,N_3328);
nor U3955 (N_3955,N_3131,N_3019);
nor U3956 (N_3956,N_3337,N_3195);
and U3957 (N_3957,N_3254,N_3240);
or U3958 (N_3958,N_3200,N_3390);
or U3959 (N_3959,N_3443,N_3468);
nand U3960 (N_3960,N_3265,N_3439);
nor U3961 (N_3961,N_3163,N_3108);
and U3962 (N_3962,N_3313,N_3220);
nand U3963 (N_3963,N_3488,N_3171);
nor U3964 (N_3964,N_3108,N_3274);
and U3965 (N_3965,N_3006,N_3325);
nor U3966 (N_3966,N_3090,N_3088);
nor U3967 (N_3967,N_3423,N_3047);
or U3968 (N_3968,N_3420,N_3295);
nand U3969 (N_3969,N_3325,N_3422);
and U3970 (N_3970,N_3272,N_3279);
nor U3971 (N_3971,N_3224,N_3164);
xnor U3972 (N_3972,N_3089,N_3153);
xor U3973 (N_3973,N_3202,N_3097);
or U3974 (N_3974,N_3310,N_3038);
nor U3975 (N_3975,N_3062,N_3014);
xor U3976 (N_3976,N_3344,N_3468);
nor U3977 (N_3977,N_3459,N_3209);
or U3978 (N_3978,N_3244,N_3188);
or U3979 (N_3979,N_3318,N_3064);
xor U3980 (N_3980,N_3011,N_3404);
xor U3981 (N_3981,N_3426,N_3242);
or U3982 (N_3982,N_3473,N_3156);
or U3983 (N_3983,N_3130,N_3374);
nand U3984 (N_3984,N_3251,N_3268);
nor U3985 (N_3985,N_3333,N_3380);
and U3986 (N_3986,N_3440,N_3074);
nor U3987 (N_3987,N_3191,N_3346);
and U3988 (N_3988,N_3038,N_3058);
or U3989 (N_3989,N_3408,N_3093);
xor U3990 (N_3990,N_3288,N_3027);
nand U3991 (N_3991,N_3411,N_3254);
or U3992 (N_3992,N_3279,N_3147);
nand U3993 (N_3993,N_3226,N_3060);
and U3994 (N_3994,N_3276,N_3455);
or U3995 (N_3995,N_3180,N_3021);
or U3996 (N_3996,N_3407,N_3022);
and U3997 (N_3997,N_3404,N_3312);
nand U3998 (N_3998,N_3309,N_3013);
and U3999 (N_3999,N_3001,N_3219);
nor U4000 (N_4000,N_3564,N_3580);
nand U4001 (N_4001,N_3925,N_3825);
nor U4002 (N_4002,N_3670,N_3881);
nand U4003 (N_4003,N_3746,N_3575);
nor U4004 (N_4004,N_3877,N_3757);
nand U4005 (N_4005,N_3504,N_3762);
and U4006 (N_4006,N_3519,N_3539);
xor U4007 (N_4007,N_3926,N_3721);
nor U4008 (N_4008,N_3745,N_3584);
or U4009 (N_4009,N_3635,N_3809);
or U4010 (N_4010,N_3720,N_3694);
and U4011 (N_4011,N_3761,N_3653);
xnor U4012 (N_4012,N_3585,N_3936);
xor U4013 (N_4013,N_3513,N_3978);
nand U4014 (N_4014,N_3536,N_3606);
nand U4015 (N_4015,N_3582,N_3736);
or U4016 (N_4016,N_3544,N_3968);
or U4017 (N_4017,N_3967,N_3930);
nor U4018 (N_4018,N_3953,N_3661);
nand U4019 (N_4019,N_3971,N_3888);
nand U4020 (N_4020,N_3975,N_3916);
or U4021 (N_4021,N_3727,N_3908);
xor U4022 (N_4022,N_3867,N_3759);
and U4023 (N_4023,N_3939,N_3714);
nor U4024 (N_4024,N_3545,N_3807);
or U4025 (N_4025,N_3955,N_3501);
or U4026 (N_4026,N_3569,N_3647);
nand U4027 (N_4027,N_3943,N_3945);
and U4028 (N_4028,N_3724,N_3543);
nand U4029 (N_4029,N_3725,N_3534);
and U4030 (N_4030,N_3652,N_3834);
or U4031 (N_4031,N_3615,N_3704);
and U4032 (N_4032,N_3707,N_3567);
xnor U4033 (N_4033,N_3516,N_3904);
or U4034 (N_4034,N_3586,N_3705);
xnor U4035 (N_4035,N_3642,N_3597);
and U4036 (N_4036,N_3612,N_3716);
nand U4037 (N_4037,N_3913,N_3944);
xor U4038 (N_4038,N_3795,N_3832);
and U4039 (N_4039,N_3970,N_3894);
nor U4040 (N_4040,N_3817,N_3658);
or U4041 (N_4041,N_3682,N_3770);
nand U4042 (N_4042,N_3747,N_3677);
nor U4043 (N_4043,N_3800,N_3703);
nor U4044 (N_4044,N_3660,N_3875);
nand U4045 (N_4045,N_3787,N_3988);
xnor U4046 (N_4046,N_3692,N_3903);
nor U4047 (N_4047,N_3851,N_3644);
nor U4048 (N_4048,N_3711,N_3591);
nand U4049 (N_4049,N_3574,N_3878);
nand U4050 (N_4050,N_3909,N_3616);
nor U4051 (N_4051,N_3588,N_3884);
and U4052 (N_4052,N_3623,N_3651);
and U4053 (N_4053,N_3838,N_3897);
nor U4054 (N_4054,N_3594,N_3611);
or U4055 (N_4055,N_3932,N_3592);
nand U4056 (N_4056,N_3992,N_3781);
nor U4057 (N_4057,N_3981,N_3828);
nand U4058 (N_4058,N_3537,N_3910);
and U4059 (N_4059,N_3603,N_3928);
or U4060 (N_4060,N_3870,N_3871);
and U4061 (N_4061,N_3823,N_3608);
xor U4062 (N_4062,N_3990,N_3985);
xor U4063 (N_4063,N_3960,N_3785);
xnor U4064 (N_4064,N_3752,N_3912);
and U4065 (N_4065,N_3693,N_3958);
nand U4066 (N_4066,N_3901,N_3502);
nor U4067 (N_4067,N_3998,N_3982);
and U4068 (N_4068,N_3741,N_3850);
and U4069 (N_4069,N_3915,N_3805);
nand U4070 (N_4070,N_3627,N_3751);
nand U4071 (N_4071,N_3590,N_3510);
nor U4072 (N_4072,N_3696,N_3866);
nor U4073 (N_4073,N_3972,N_3788);
and U4074 (N_4074,N_3645,N_3523);
and U4075 (N_4075,N_3771,N_3710);
or U4076 (N_4076,N_3515,N_3654);
or U4077 (N_4077,N_3620,N_3667);
nand U4078 (N_4078,N_3622,N_3614);
xnor U4079 (N_4079,N_3893,N_3695);
nor U4080 (N_4080,N_3547,N_3835);
nand U4081 (N_4081,N_3854,N_3554);
nand U4082 (N_4082,N_3931,N_3522);
nand U4083 (N_4083,N_3768,N_3637);
and U4084 (N_4084,N_3507,N_3719);
nor U4085 (N_4085,N_3793,N_3680);
and U4086 (N_4086,N_3839,N_3605);
or U4087 (N_4087,N_3733,N_3966);
xnor U4088 (N_4088,N_3822,N_3549);
or U4089 (N_4089,N_3902,N_3646);
nor U4090 (N_4090,N_3948,N_3824);
nor U4091 (N_4091,N_3500,N_3609);
nor U4092 (N_4092,N_3869,N_3780);
or U4093 (N_4093,N_3688,N_3900);
nand U4094 (N_4094,N_3666,N_3923);
xnor U4095 (N_4095,N_3618,N_3553);
and U4096 (N_4096,N_3613,N_3775);
nor U4097 (N_4097,N_3810,N_3779);
and U4098 (N_4098,N_3621,N_3599);
nor U4099 (N_4099,N_3526,N_3865);
nor U4100 (N_4100,N_3836,N_3626);
nor U4101 (N_4101,N_3994,N_3989);
and U4102 (N_4102,N_3831,N_3540);
and U4103 (N_4103,N_3673,N_3708);
xnor U4104 (N_4104,N_3699,N_3706);
xor U4105 (N_4105,N_3701,N_3639);
nor U4106 (N_4106,N_3541,N_3528);
nand U4107 (N_4107,N_3969,N_3617);
nand U4108 (N_4108,N_3525,N_3572);
or U4109 (N_4109,N_3689,N_3718);
and U4110 (N_4110,N_3961,N_3521);
and U4111 (N_4111,N_3565,N_3734);
or U4112 (N_4112,N_3740,N_3949);
nand U4113 (N_4113,N_3940,N_3976);
xnor U4114 (N_4114,N_3550,N_3873);
nor U4115 (N_4115,N_3772,N_3520);
xor U4116 (N_4116,N_3630,N_3715);
or U4117 (N_4117,N_3907,N_3533);
and U4118 (N_4118,N_3995,N_3886);
and U4119 (N_4119,N_3722,N_3852);
xnor U4120 (N_4120,N_3937,N_3563);
xor U4121 (N_4121,N_3980,N_3959);
xor U4122 (N_4122,N_3796,N_3748);
nand U4123 (N_4123,N_3610,N_3571);
xnor U4124 (N_4124,N_3843,N_3511);
or U4125 (N_4125,N_3802,N_3655);
nand U4126 (N_4126,N_3774,N_3503);
nand U4127 (N_4127,N_3672,N_3755);
xor U4128 (N_4128,N_3678,N_3847);
or U4129 (N_4129,N_3974,N_3773);
and U4130 (N_4130,N_3794,N_3837);
nor U4131 (N_4131,N_3963,N_3636);
xnor U4132 (N_4132,N_3892,N_3538);
and U4133 (N_4133,N_3702,N_3887);
or U4134 (N_4134,N_3532,N_3786);
nand U4135 (N_4135,N_3927,N_3938);
nand U4136 (N_4136,N_3973,N_3880);
nand U4137 (N_4137,N_3987,N_3600);
xnor U4138 (N_4138,N_3531,N_3579);
and U4139 (N_4139,N_3861,N_3804);
nor U4140 (N_4140,N_3983,N_3846);
nor U4141 (N_4141,N_3864,N_3561);
nand U4142 (N_4142,N_3862,N_3849);
xnor U4143 (N_4143,N_3557,N_3763);
xnor U4144 (N_4144,N_3530,N_3941);
nand U4145 (N_4145,N_3942,N_3656);
or U4146 (N_4146,N_3629,N_3679);
xor U4147 (N_4147,N_3820,N_3924);
and U4148 (N_4148,N_3581,N_3596);
xor U4149 (N_4149,N_3950,N_3681);
or U4150 (N_4150,N_3999,N_3709);
nor U4151 (N_4151,N_3675,N_3889);
nand U4152 (N_4152,N_3638,N_3684);
and U4153 (N_4153,N_3542,N_3555);
and U4154 (N_4154,N_3598,N_3602);
nand U4155 (N_4155,N_3662,N_3643);
nor U4156 (N_4156,N_3814,N_3855);
xor U4157 (N_4157,N_3514,N_3857);
and U4158 (N_4158,N_3566,N_3568);
nor U4159 (N_4159,N_3791,N_3683);
nor U4160 (N_4160,N_3601,N_3876);
or U4161 (N_4161,N_3778,N_3535);
and U4162 (N_4162,N_3821,N_3663);
nand U4163 (N_4163,N_3595,N_3754);
xor U4164 (N_4164,N_3735,N_3765);
xor U4165 (N_4165,N_3801,N_3883);
nor U4166 (N_4166,N_3691,N_3798);
or U4167 (N_4167,N_3783,N_3641);
and U4168 (N_4168,N_3738,N_3685);
nand U4169 (N_4169,N_3979,N_3858);
and U4170 (N_4170,N_3728,N_3750);
or U4171 (N_4171,N_3593,N_3921);
and U4172 (N_4172,N_3792,N_3607);
xnor U4173 (N_4173,N_3833,N_3841);
nor U4174 (N_4174,N_3885,N_3640);
nand U4175 (N_4175,N_3844,N_3700);
and U4176 (N_4176,N_3697,N_3729);
or U4177 (N_4177,N_3856,N_3576);
or U4178 (N_4178,N_3631,N_3556);
nor U4179 (N_4179,N_3911,N_3559);
and U4180 (N_4180,N_3717,N_3946);
nand U4181 (N_4181,N_3506,N_3578);
or U4182 (N_4182,N_3845,N_3756);
or U4183 (N_4183,N_3665,N_3764);
and U4184 (N_4184,N_3997,N_3562);
and U4185 (N_4185,N_3650,N_3826);
or U4186 (N_4186,N_3984,N_3790);
nor U4187 (N_4187,N_3687,N_3782);
or U4188 (N_4188,N_3558,N_3776);
xor U4189 (N_4189,N_3753,N_3674);
and U4190 (N_4190,N_3731,N_3957);
nor U4191 (N_4191,N_3977,N_3874);
and U4192 (N_4192,N_3818,N_3777);
or U4193 (N_4193,N_3548,N_3934);
nor U4194 (N_4194,N_3905,N_3732);
nor U4195 (N_4195,N_3524,N_3829);
nand U4196 (N_4196,N_3895,N_3632);
and U4197 (N_4197,N_3784,N_3690);
nand U4198 (N_4198,N_3552,N_3604);
or U4199 (N_4199,N_3922,N_3739);
xor U4200 (N_4200,N_3758,N_3956);
xor U4201 (N_4201,N_3799,N_3742);
nand U4202 (N_4202,N_3951,N_3527);
nand U4203 (N_4203,N_3860,N_3676);
xnor U4204 (N_4204,N_3853,N_3789);
or U4205 (N_4205,N_3518,N_3917);
xor U4206 (N_4206,N_3668,N_3920);
and U4207 (N_4207,N_3749,N_3570);
nand U4208 (N_4208,N_3664,N_3624);
nor U4209 (N_4209,N_3509,N_3872);
xor U4210 (N_4210,N_3808,N_3769);
and U4211 (N_4211,N_3628,N_3819);
nor U4212 (N_4212,N_3659,N_3813);
nand U4213 (N_4213,N_3842,N_3508);
or U4214 (N_4214,N_3589,N_3906);
nor U4215 (N_4215,N_3649,N_3899);
xor U4216 (N_4216,N_3577,N_3737);
nor U4217 (N_4217,N_3767,N_3993);
and U4218 (N_4218,N_3634,N_3929);
or U4219 (N_4219,N_3898,N_3657);
and U4220 (N_4220,N_3723,N_3879);
nor U4221 (N_4221,N_3760,N_3766);
or U4222 (N_4222,N_3954,N_3648);
nand U4223 (N_4223,N_3830,N_3863);
and U4224 (N_4224,N_3868,N_3986);
nand U4225 (N_4225,N_3996,N_3848);
nor U4226 (N_4226,N_3947,N_3965);
nand U4227 (N_4227,N_3573,N_3505);
nand U4228 (N_4228,N_3812,N_3806);
xnor U4229 (N_4229,N_3583,N_3633);
and U4230 (N_4230,N_3619,N_3713);
nor U4231 (N_4231,N_3712,N_3890);
nand U4232 (N_4232,N_3859,N_3686);
xor U4233 (N_4233,N_3882,N_3744);
nor U4234 (N_4234,N_3726,N_3560);
or U4235 (N_4235,N_3811,N_3891);
xnor U4236 (N_4236,N_3962,N_3587);
nand U4237 (N_4237,N_3952,N_3517);
or U4238 (N_4238,N_3896,N_3669);
nor U4239 (N_4239,N_3803,N_3512);
and U4240 (N_4240,N_3698,N_3840);
xnor U4241 (N_4241,N_3797,N_3914);
and U4242 (N_4242,N_3815,N_3743);
xor U4243 (N_4243,N_3671,N_3827);
nor U4244 (N_4244,N_3933,N_3964);
or U4245 (N_4245,N_3935,N_3546);
and U4246 (N_4246,N_3816,N_3529);
and U4247 (N_4247,N_3625,N_3730);
nand U4248 (N_4248,N_3551,N_3991);
and U4249 (N_4249,N_3918,N_3919);
or U4250 (N_4250,N_3786,N_3712);
and U4251 (N_4251,N_3824,N_3909);
or U4252 (N_4252,N_3668,N_3713);
and U4253 (N_4253,N_3846,N_3958);
nand U4254 (N_4254,N_3944,N_3696);
xnor U4255 (N_4255,N_3879,N_3962);
nand U4256 (N_4256,N_3938,N_3505);
and U4257 (N_4257,N_3745,N_3858);
or U4258 (N_4258,N_3685,N_3706);
or U4259 (N_4259,N_3603,N_3585);
or U4260 (N_4260,N_3798,N_3717);
xnor U4261 (N_4261,N_3634,N_3575);
xor U4262 (N_4262,N_3962,N_3772);
xor U4263 (N_4263,N_3780,N_3558);
nand U4264 (N_4264,N_3813,N_3806);
nand U4265 (N_4265,N_3766,N_3726);
xnor U4266 (N_4266,N_3691,N_3657);
xor U4267 (N_4267,N_3542,N_3709);
and U4268 (N_4268,N_3718,N_3591);
or U4269 (N_4269,N_3906,N_3884);
xnor U4270 (N_4270,N_3532,N_3718);
xnor U4271 (N_4271,N_3774,N_3868);
nand U4272 (N_4272,N_3943,N_3806);
and U4273 (N_4273,N_3674,N_3980);
nor U4274 (N_4274,N_3665,N_3963);
nand U4275 (N_4275,N_3965,N_3648);
xor U4276 (N_4276,N_3516,N_3569);
nor U4277 (N_4277,N_3572,N_3697);
and U4278 (N_4278,N_3523,N_3823);
xnor U4279 (N_4279,N_3861,N_3783);
nand U4280 (N_4280,N_3508,N_3517);
nor U4281 (N_4281,N_3781,N_3811);
nor U4282 (N_4282,N_3698,N_3522);
or U4283 (N_4283,N_3502,N_3594);
xor U4284 (N_4284,N_3810,N_3840);
and U4285 (N_4285,N_3879,N_3958);
and U4286 (N_4286,N_3767,N_3990);
nor U4287 (N_4287,N_3514,N_3958);
nand U4288 (N_4288,N_3603,N_3723);
or U4289 (N_4289,N_3774,N_3962);
or U4290 (N_4290,N_3834,N_3787);
xor U4291 (N_4291,N_3812,N_3721);
or U4292 (N_4292,N_3734,N_3861);
nor U4293 (N_4293,N_3930,N_3999);
xnor U4294 (N_4294,N_3745,N_3780);
or U4295 (N_4295,N_3768,N_3930);
nor U4296 (N_4296,N_3955,N_3950);
or U4297 (N_4297,N_3662,N_3912);
nor U4298 (N_4298,N_3727,N_3569);
or U4299 (N_4299,N_3500,N_3683);
and U4300 (N_4300,N_3699,N_3609);
nand U4301 (N_4301,N_3903,N_3711);
nor U4302 (N_4302,N_3976,N_3618);
nor U4303 (N_4303,N_3608,N_3981);
xor U4304 (N_4304,N_3649,N_3975);
nor U4305 (N_4305,N_3736,N_3549);
nand U4306 (N_4306,N_3976,N_3525);
nand U4307 (N_4307,N_3673,N_3525);
nand U4308 (N_4308,N_3797,N_3712);
and U4309 (N_4309,N_3678,N_3789);
or U4310 (N_4310,N_3854,N_3664);
or U4311 (N_4311,N_3605,N_3818);
or U4312 (N_4312,N_3563,N_3503);
and U4313 (N_4313,N_3836,N_3894);
nor U4314 (N_4314,N_3699,N_3641);
nor U4315 (N_4315,N_3750,N_3576);
and U4316 (N_4316,N_3895,N_3971);
or U4317 (N_4317,N_3952,N_3970);
and U4318 (N_4318,N_3815,N_3996);
nand U4319 (N_4319,N_3618,N_3627);
nand U4320 (N_4320,N_3765,N_3566);
or U4321 (N_4321,N_3529,N_3901);
xnor U4322 (N_4322,N_3988,N_3560);
or U4323 (N_4323,N_3951,N_3782);
or U4324 (N_4324,N_3620,N_3702);
xor U4325 (N_4325,N_3558,N_3834);
xor U4326 (N_4326,N_3558,N_3818);
and U4327 (N_4327,N_3741,N_3904);
nor U4328 (N_4328,N_3744,N_3658);
nand U4329 (N_4329,N_3932,N_3750);
and U4330 (N_4330,N_3680,N_3558);
or U4331 (N_4331,N_3934,N_3859);
nor U4332 (N_4332,N_3956,N_3920);
and U4333 (N_4333,N_3648,N_3916);
xnor U4334 (N_4334,N_3741,N_3923);
and U4335 (N_4335,N_3644,N_3619);
nand U4336 (N_4336,N_3521,N_3621);
or U4337 (N_4337,N_3609,N_3665);
and U4338 (N_4338,N_3957,N_3774);
or U4339 (N_4339,N_3698,N_3667);
and U4340 (N_4340,N_3973,N_3620);
nand U4341 (N_4341,N_3917,N_3907);
and U4342 (N_4342,N_3582,N_3674);
xor U4343 (N_4343,N_3854,N_3950);
or U4344 (N_4344,N_3722,N_3668);
and U4345 (N_4345,N_3522,N_3765);
nor U4346 (N_4346,N_3813,N_3538);
or U4347 (N_4347,N_3841,N_3785);
or U4348 (N_4348,N_3577,N_3861);
xor U4349 (N_4349,N_3547,N_3505);
nor U4350 (N_4350,N_3580,N_3697);
nor U4351 (N_4351,N_3928,N_3563);
nand U4352 (N_4352,N_3514,N_3802);
and U4353 (N_4353,N_3786,N_3589);
nand U4354 (N_4354,N_3511,N_3835);
and U4355 (N_4355,N_3571,N_3751);
or U4356 (N_4356,N_3950,N_3614);
and U4357 (N_4357,N_3538,N_3592);
and U4358 (N_4358,N_3890,N_3609);
or U4359 (N_4359,N_3809,N_3717);
and U4360 (N_4360,N_3805,N_3505);
nor U4361 (N_4361,N_3622,N_3853);
nor U4362 (N_4362,N_3804,N_3736);
or U4363 (N_4363,N_3855,N_3656);
xnor U4364 (N_4364,N_3910,N_3745);
nor U4365 (N_4365,N_3534,N_3809);
and U4366 (N_4366,N_3545,N_3718);
nand U4367 (N_4367,N_3940,N_3788);
xor U4368 (N_4368,N_3698,N_3617);
nor U4369 (N_4369,N_3866,N_3561);
and U4370 (N_4370,N_3920,N_3892);
or U4371 (N_4371,N_3626,N_3517);
or U4372 (N_4372,N_3821,N_3569);
or U4373 (N_4373,N_3642,N_3803);
xor U4374 (N_4374,N_3708,N_3665);
xnor U4375 (N_4375,N_3847,N_3931);
or U4376 (N_4376,N_3677,N_3943);
nor U4377 (N_4377,N_3767,N_3659);
xnor U4378 (N_4378,N_3791,N_3711);
or U4379 (N_4379,N_3798,N_3913);
xnor U4380 (N_4380,N_3984,N_3840);
and U4381 (N_4381,N_3582,N_3745);
xor U4382 (N_4382,N_3966,N_3529);
or U4383 (N_4383,N_3628,N_3666);
nand U4384 (N_4384,N_3749,N_3859);
xor U4385 (N_4385,N_3829,N_3882);
xnor U4386 (N_4386,N_3661,N_3595);
xnor U4387 (N_4387,N_3670,N_3742);
or U4388 (N_4388,N_3748,N_3830);
nor U4389 (N_4389,N_3731,N_3794);
or U4390 (N_4390,N_3736,N_3557);
or U4391 (N_4391,N_3598,N_3735);
nor U4392 (N_4392,N_3852,N_3796);
xnor U4393 (N_4393,N_3906,N_3658);
nand U4394 (N_4394,N_3589,N_3725);
xor U4395 (N_4395,N_3886,N_3669);
and U4396 (N_4396,N_3560,N_3735);
and U4397 (N_4397,N_3742,N_3896);
and U4398 (N_4398,N_3725,N_3747);
nand U4399 (N_4399,N_3840,N_3842);
nor U4400 (N_4400,N_3926,N_3568);
and U4401 (N_4401,N_3642,N_3523);
or U4402 (N_4402,N_3867,N_3909);
or U4403 (N_4403,N_3684,N_3538);
nand U4404 (N_4404,N_3938,N_3614);
nand U4405 (N_4405,N_3938,N_3764);
nor U4406 (N_4406,N_3688,N_3969);
and U4407 (N_4407,N_3888,N_3666);
or U4408 (N_4408,N_3858,N_3821);
nor U4409 (N_4409,N_3649,N_3514);
and U4410 (N_4410,N_3976,N_3579);
xor U4411 (N_4411,N_3818,N_3973);
and U4412 (N_4412,N_3727,N_3692);
and U4413 (N_4413,N_3560,N_3605);
and U4414 (N_4414,N_3998,N_3895);
xor U4415 (N_4415,N_3681,N_3854);
or U4416 (N_4416,N_3785,N_3952);
nand U4417 (N_4417,N_3984,N_3587);
nand U4418 (N_4418,N_3750,N_3653);
and U4419 (N_4419,N_3993,N_3781);
xor U4420 (N_4420,N_3981,N_3707);
nor U4421 (N_4421,N_3806,N_3572);
or U4422 (N_4422,N_3627,N_3546);
xor U4423 (N_4423,N_3512,N_3797);
or U4424 (N_4424,N_3873,N_3816);
nor U4425 (N_4425,N_3886,N_3551);
nand U4426 (N_4426,N_3611,N_3677);
nand U4427 (N_4427,N_3944,N_3885);
xor U4428 (N_4428,N_3633,N_3922);
nand U4429 (N_4429,N_3562,N_3611);
nor U4430 (N_4430,N_3839,N_3971);
and U4431 (N_4431,N_3978,N_3852);
and U4432 (N_4432,N_3872,N_3775);
nand U4433 (N_4433,N_3947,N_3696);
nor U4434 (N_4434,N_3923,N_3985);
and U4435 (N_4435,N_3734,N_3641);
xor U4436 (N_4436,N_3715,N_3849);
nor U4437 (N_4437,N_3720,N_3750);
xor U4438 (N_4438,N_3560,N_3817);
or U4439 (N_4439,N_3819,N_3827);
nor U4440 (N_4440,N_3681,N_3685);
or U4441 (N_4441,N_3556,N_3887);
or U4442 (N_4442,N_3969,N_3598);
xnor U4443 (N_4443,N_3933,N_3568);
xor U4444 (N_4444,N_3958,N_3957);
and U4445 (N_4445,N_3900,N_3637);
or U4446 (N_4446,N_3605,N_3804);
nand U4447 (N_4447,N_3690,N_3758);
nor U4448 (N_4448,N_3763,N_3582);
xor U4449 (N_4449,N_3987,N_3583);
or U4450 (N_4450,N_3841,N_3927);
xor U4451 (N_4451,N_3914,N_3949);
and U4452 (N_4452,N_3509,N_3576);
xnor U4453 (N_4453,N_3749,N_3877);
or U4454 (N_4454,N_3996,N_3853);
or U4455 (N_4455,N_3892,N_3649);
xnor U4456 (N_4456,N_3576,N_3508);
nand U4457 (N_4457,N_3850,N_3831);
or U4458 (N_4458,N_3998,N_3577);
and U4459 (N_4459,N_3705,N_3570);
nor U4460 (N_4460,N_3567,N_3792);
xnor U4461 (N_4461,N_3670,N_3857);
nor U4462 (N_4462,N_3698,N_3902);
and U4463 (N_4463,N_3825,N_3763);
or U4464 (N_4464,N_3665,N_3911);
xnor U4465 (N_4465,N_3758,N_3764);
nand U4466 (N_4466,N_3675,N_3620);
or U4467 (N_4467,N_3724,N_3826);
or U4468 (N_4468,N_3531,N_3869);
nand U4469 (N_4469,N_3708,N_3508);
or U4470 (N_4470,N_3615,N_3946);
nand U4471 (N_4471,N_3926,N_3511);
and U4472 (N_4472,N_3966,N_3937);
nor U4473 (N_4473,N_3990,N_3977);
and U4474 (N_4474,N_3806,N_3829);
nor U4475 (N_4475,N_3708,N_3897);
nand U4476 (N_4476,N_3505,N_3960);
nor U4477 (N_4477,N_3620,N_3783);
xor U4478 (N_4478,N_3527,N_3667);
nand U4479 (N_4479,N_3897,N_3975);
or U4480 (N_4480,N_3527,N_3613);
nor U4481 (N_4481,N_3630,N_3972);
nor U4482 (N_4482,N_3501,N_3557);
nand U4483 (N_4483,N_3711,N_3949);
and U4484 (N_4484,N_3835,N_3512);
or U4485 (N_4485,N_3762,N_3711);
nand U4486 (N_4486,N_3848,N_3535);
nor U4487 (N_4487,N_3962,N_3874);
and U4488 (N_4488,N_3667,N_3945);
and U4489 (N_4489,N_3615,N_3886);
or U4490 (N_4490,N_3938,N_3554);
nor U4491 (N_4491,N_3975,N_3882);
and U4492 (N_4492,N_3913,N_3579);
nor U4493 (N_4493,N_3695,N_3503);
xnor U4494 (N_4494,N_3616,N_3522);
and U4495 (N_4495,N_3841,N_3871);
or U4496 (N_4496,N_3512,N_3870);
nand U4497 (N_4497,N_3627,N_3786);
xnor U4498 (N_4498,N_3850,N_3771);
nand U4499 (N_4499,N_3723,N_3561);
xor U4500 (N_4500,N_4390,N_4384);
xor U4501 (N_4501,N_4080,N_4392);
or U4502 (N_4502,N_4295,N_4443);
nor U4503 (N_4503,N_4374,N_4039);
and U4504 (N_4504,N_4296,N_4011);
nor U4505 (N_4505,N_4079,N_4228);
or U4506 (N_4506,N_4234,N_4439);
nor U4507 (N_4507,N_4438,N_4471);
nand U4508 (N_4508,N_4282,N_4357);
nand U4509 (N_4509,N_4403,N_4365);
nor U4510 (N_4510,N_4211,N_4152);
xor U4511 (N_4511,N_4141,N_4214);
nor U4512 (N_4512,N_4272,N_4178);
xnor U4513 (N_4513,N_4107,N_4288);
and U4514 (N_4514,N_4327,N_4358);
or U4515 (N_4515,N_4492,N_4216);
and U4516 (N_4516,N_4381,N_4275);
nor U4517 (N_4517,N_4019,N_4434);
or U4518 (N_4518,N_4078,N_4468);
nand U4519 (N_4519,N_4267,N_4205);
nand U4520 (N_4520,N_4407,N_4363);
xnor U4521 (N_4521,N_4355,N_4190);
nor U4522 (N_4522,N_4105,N_4068);
and U4523 (N_4523,N_4370,N_4281);
and U4524 (N_4524,N_4343,N_4408);
nand U4525 (N_4525,N_4171,N_4143);
nand U4526 (N_4526,N_4274,N_4353);
and U4527 (N_4527,N_4032,N_4386);
nand U4528 (N_4528,N_4454,N_4306);
xor U4529 (N_4529,N_4337,N_4473);
nor U4530 (N_4530,N_4488,N_4298);
xnor U4531 (N_4531,N_4168,N_4486);
or U4532 (N_4532,N_4360,N_4184);
nor U4533 (N_4533,N_4125,N_4478);
nor U4534 (N_4534,N_4284,N_4301);
and U4535 (N_4535,N_4110,N_4305);
xor U4536 (N_4536,N_4132,N_4015);
xor U4537 (N_4537,N_4076,N_4270);
and U4538 (N_4538,N_4003,N_4450);
and U4539 (N_4539,N_4457,N_4349);
or U4540 (N_4540,N_4200,N_4223);
and U4541 (N_4541,N_4145,N_4226);
nor U4542 (N_4542,N_4022,N_4236);
or U4543 (N_4543,N_4065,N_4163);
nand U4544 (N_4544,N_4176,N_4209);
and U4545 (N_4545,N_4120,N_4091);
xnor U4546 (N_4546,N_4302,N_4480);
and U4547 (N_4547,N_4331,N_4150);
xnor U4548 (N_4548,N_4151,N_4461);
and U4549 (N_4549,N_4098,N_4332);
or U4550 (N_4550,N_4398,N_4289);
nor U4551 (N_4551,N_4266,N_4138);
xor U4552 (N_4552,N_4241,N_4417);
and U4553 (N_4553,N_4231,N_4127);
nand U4554 (N_4554,N_4220,N_4402);
xor U4555 (N_4555,N_4293,N_4045);
nand U4556 (N_4556,N_4193,N_4207);
nand U4557 (N_4557,N_4073,N_4255);
and U4558 (N_4558,N_4056,N_4062);
nand U4559 (N_4559,N_4232,N_4013);
nand U4560 (N_4560,N_4458,N_4376);
and U4561 (N_4561,N_4257,N_4380);
xnor U4562 (N_4562,N_4169,N_4007);
xor U4563 (N_4563,N_4320,N_4042);
and U4564 (N_4564,N_4081,N_4435);
nor U4565 (N_4565,N_4005,N_4038);
or U4566 (N_4566,N_4246,N_4099);
and U4567 (N_4567,N_4428,N_4047);
and U4568 (N_4568,N_4414,N_4009);
or U4569 (N_4569,N_4044,N_4291);
nor U4570 (N_4570,N_4304,N_4177);
or U4571 (N_4571,N_4425,N_4344);
xnor U4572 (N_4572,N_4256,N_4156);
or U4573 (N_4573,N_4279,N_4496);
nand U4574 (N_4574,N_4404,N_4271);
xor U4575 (N_4575,N_4087,N_4467);
nand U4576 (N_4576,N_4033,N_4373);
and U4577 (N_4577,N_4070,N_4139);
nor U4578 (N_4578,N_4440,N_4208);
xnor U4579 (N_4579,N_4401,N_4490);
nor U4580 (N_4580,N_4411,N_4021);
or U4581 (N_4581,N_4175,N_4061);
nand U4582 (N_4582,N_4074,N_4052);
nand U4583 (N_4583,N_4122,N_4261);
or U4584 (N_4584,N_4248,N_4262);
xnor U4585 (N_4585,N_4340,N_4174);
xnor U4586 (N_4586,N_4029,N_4130);
nor U4587 (N_4587,N_4452,N_4333);
nor U4588 (N_4588,N_4335,N_4499);
nor U4589 (N_4589,N_4054,N_4329);
nor U4590 (N_4590,N_4463,N_4245);
xor U4591 (N_4591,N_4339,N_4149);
nand U4592 (N_4592,N_4476,N_4240);
xnor U4593 (N_4593,N_4194,N_4394);
nor U4594 (N_4594,N_4160,N_4451);
nand U4595 (N_4595,N_4377,N_4406);
and U4596 (N_4596,N_4067,N_4427);
nor U4597 (N_4597,N_4260,N_4325);
or U4598 (N_4598,N_4225,N_4046);
xor U4599 (N_4599,N_4183,N_4385);
and U4600 (N_4600,N_4410,N_4158);
nor U4601 (N_4601,N_4153,N_4412);
nand U4602 (N_4602,N_4126,N_4089);
xor U4603 (N_4603,N_4109,N_4104);
nand U4604 (N_4604,N_4182,N_4135);
and U4605 (N_4605,N_4375,N_4326);
nand U4606 (N_4606,N_4354,N_4244);
nand U4607 (N_4607,N_4114,N_4113);
nand U4608 (N_4608,N_4491,N_4308);
xnor U4609 (N_4609,N_4314,N_4161);
nand U4610 (N_4610,N_4484,N_4487);
xnor U4611 (N_4611,N_4229,N_4053);
xor U4612 (N_4612,N_4419,N_4187);
and U4613 (N_4613,N_4196,N_4085);
xor U4614 (N_4614,N_4263,N_4112);
xor U4615 (N_4615,N_4023,N_4323);
nor U4616 (N_4616,N_4198,N_4140);
or U4617 (N_4617,N_4278,N_4106);
nor U4618 (N_4618,N_4167,N_4215);
xor U4619 (N_4619,N_4498,N_4071);
nor U4620 (N_4620,N_4342,N_4083);
nand U4621 (N_4621,N_4133,N_4347);
nand U4622 (N_4622,N_4455,N_4268);
and U4623 (N_4623,N_4494,N_4155);
and U4624 (N_4624,N_4383,N_4460);
or U4625 (N_4625,N_4162,N_4362);
and U4626 (N_4626,N_4495,N_4064);
or U4627 (N_4627,N_4142,N_4233);
nand U4628 (N_4628,N_4418,N_4201);
nand U4629 (N_4629,N_4277,N_4453);
nand U4630 (N_4630,N_4307,N_4031);
and U4631 (N_4631,N_4103,N_4247);
or U4632 (N_4632,N_4322,N_4286);
xnor U4633 (N_4633,N_4111,N_4086);
xor U4634 (N_4634,N_4294,N_4287);
nor U4635 (N_4635,N_4059,N_4313);
and U4636 (N_4636,N_4474,N_4117);
nor U4637 (N_4637,N_4250,N_4134);
nor U4638 (N_4638,N_4433,N_4217);
nor U4639 (N_4639,N_4048,N_4422);
or U4640 (N_4640,N_4077,N_4060);
or U4641 (N_4641,N_4265,N_4049);
nand U4642 (N_4642,N_4123,N_4028);
and U4643 (N_4643,N_4129,N_4318);
nor U4644 (N_4644,N_4035,N_4400);
nand U4645 (N_4645,N_4466,N_4118);
xor U4646 (N_4646,N_4010,N_4075);
and U4647 (N_4647,N_4203,N_4324);
or U4648 (N_4648,N_4489,N_4356);
nand U4649 (N_4649,N_4227,N_4391);
xnor U4650 (N_4650,N_4379,N_4165);
xor U4651 (N_4651,N_4100,N_4396);
xnor U4652 (N_4652,N_4051,N_4025);
or U4653 (N_4653,N_4368,N_4172);
or U4654 (N_4654,N_4456,N_4020);
and U4655 (N_4655,N_4101,N_4243);
xnor U4656 (N_4656,N_4102,N_4202);
nor U4657 (N_4657,N_4413,N_4040);
or U4658 (N_4658,N_4283,N_4336);
nand U4659 (N_4659,N_4469,N_4252);
and U4660 (N_4660,N_4334,N_4470);
xor U4661 (N_4661,N_4088,N_4399);
nor U4662 (N_4662,N_4312,N_4297);
and U4663 (N_4663,N_4147,N_4222);
xor U4664 (N_4664,N_4242,N_4426);
and U4665 (N_4665,N_4210,N_4321);
nand U4666 (N_4666,N_4230,N_4382);
and U4667 (N_4667,N_4273,N_4166);
or U4668 (N_4668,N_4173,N_4280);
xnor U4669 (N_4669,N_4405,N_4027);
or U4670 (N_4670,N_4001,N_4185);
nand U4671 (N_4671,N_4254,N_4014);
xnor U4672 (N_4672,N_4371,N_4481);
xor U4673 (N_4673,N_4462,N_4094);
or U4674 (N_4674,N_4148,N_4164);
and U4675 (N_4675,N_4303,N_4206);
nor U4676 (N_4676,N_4006,N_4219);
or U4677 (N_4677,N_4179,N_4465);
xnor U4678 (N_4678,N_4437,N_4097);
nor U4679 (N_4679,N_4004,N_4115);
nor U4680 (N_4680,N_4249,N_4264);
and U4681 (N_4681,N_4072,N_4442);
nor U4682 (N_4682,N_4002,N_4195);
or U4683 (N_4683,N_4012,N_4483);
xor U4684 (N_4684,N_4181,N_4387);
nor U4685 (N_4685,N_4237,N_4366);
xor U4686 (N_4686,N_4258,N_4497);
xnor U4687 (N_4687,N_4186,N_4144);
nor U4688 (N_4688,N_4199,N_4095);
nor U4689 (N_4689,N_4204,N_4449);
xnor U4690 (N_4690,N_4180,N_4309);
or U4691 (N_4691,N_4034,N_4090);
xnor U4692 (N_4692,N_4341,N_4235);
xor U4693 (N_4693,N_4212,N_4475);
or U4694 (N_4694,N_4108,N_4397);
and U4695 (N_4695,N_4269,N_4084);
and U4696 (N_4696,N_4393,N_4436);
or U4697 (N_4697,N_4066,N_4253);
and U4698 (N_4698,N_4459,N_4285);
nor U4699 (N_4699,N_4157,N_4479);
nand U4700 (N_4700,N_4421,N_4448);
nand U4701 (N_4701,N_4119,N_4316);
or U4702 (N_4702,N_4369,N_4218);
or U4703 (N_4703,N_4050,N_4146);
and U4704 (N_4704,N_4477,N_4482);
or U4705 (N_4705,N_4063,N_4030);
nor U4706 (N_4706,N_4092,N_4300);
nor U4707 (N_4707,N_4446,N_4319);
nor U4708 (N_4708,N_4096,N_4259);
or U4709 (N_4709,N_4154,N_4359);
nand U4710 (N_4710,N_4136,N_4239);
or U4711 (N_4711,N_4213,N_4423);
or U4712 (N_4712,N_4361,N_4131);
nor U4713 (N_4713,N_4445,N_4317);
or U4714 (N_4714,N_4238,N_4159);
nand U4715 (N_4715,N_4338,N_4018);
xor U4716 (N_4716,N_4441,N_4328);
nand U4717 (N_4717,N_4082,N_4367);
nor U4718 (N_4718,N_4221,N_4430);
nor U4719 (N_4719,N_4057,N_4416);
and U4720 (N_4720,N_4008,N_4348);
or U4721 (N_4721,N_4191,N_4330);
xor U4722 (N_4722,N_4395,N_4351);
or U4723 (N_4723,N_4388,N_4409);
xor U4724 (N_4724,N_4292,N_4485);
or U4725 (N_4725,N_4299,N_4346);
nand U4726 (N_4726,N_4058,N_4378);
or U4727 (N_4727,N_4121,N_4431);
xnor U4728 (N_4728,N_4197,N_4493);
and U4729 (N_4729,N_4026,N_4124);
or U4730 (N_4730,N_4447,N_4444);
xnor U4731 (N_4731,N_4069,N_4188);
nor U4732 (N_4732,N_4350,N_4093);
nand U4733 (N_4733,N_4224,N_4016);
nor U4734 (N_4734,N_4037,N_4424);
or U4735 (N_4735,N_4192,N_4276);
nor U4736 (N_4736,N_4432,N_4315);
or U4737 (N_4737,N_4310,N_4024);
or U4738 (N_4738,N_4116,N_4345);
nand U4739 (N_4739,N_4472,N_4251);
nor U4740 (N_4740,N_4017,N_4170);
nand U4741 (N_4741,N_4189,N_4041);
xnor U4742 (N_4742,N_4036,N_4137);
or U4743 (N_4743,N_4311,N_4290);
xnor U4744 (N_4744,N_4055,N_4043);
nor U4745 (N_4745,N_4352,N_4420);
xnor U4746 (N_4746,N_4000,N_4415);
or U4747 (N_4747,N_4389,N_4372);
or U4748 (N_4748,N_4429,N_4364);
nor U4749 (N_4749,N_4128,N_4464);
nand U4750 (N_4750,N_4085,N_4251);
nand U4751 (N_4751,N_4315,N_4455);
xor U4752 (N_4752,N_4201,N_4477);
nor U4753 (N_4753,N_4193,N_4494);
xor U4754 (N_4754,N_4396,N_4082);
xor U4755 (N_4755,N_4384,N_4476);
nand U4756 (N_4756,N_4262,N_4040);
nor U4757 (N_4757,N_4486,N_4150);
xor U4758 (N_4758,N_4092,N_4492);
xnor U4759 (N_4759,N_4245,N_4203);
nand U4760 (N_4760,N_4032,N_4414);
and U4761 (N_4761,N_4230,N_4350);
xnor U4762 (N_4762,N_4061,N_4340);
or U4763 (N_4763,N_4379,N_4241);
or U4764 (N_4764,N_4318,N_4182);
and U4765 (N_4765,N_4262,N_4414);
nor U4766 (N_4766,N_4225,N_4071);
nor U4767 (N_4767,N_4499,N_4035);
xnor U4768 (N_4768,N_4456,N_4495);
nor U4769 (N_4769,N_4499,N_4458);
nor U4770 (N_4770,N_4106,N_4274);
and U4771 (N_4771,N_4147,N_4288);
xor U4772 (N_4772,N_4397,N_4445);
xnor U4773 (N_4773,N_4015,N_4427);
or U4774 (N_4774,N_4209,N_4344);
and U4775 (N_4775,N_4359,N_4365);
nand U4776 (N_4776,N_4198,N_4186);
and U4777 (N_4777,N_4095,N_4112);
nand U4778 (N_4778,N_4379,N_4338);
xor U4779 (N_4779,N_4327,N_4278);
nor U4780 (N_4780,N_4068,N_4459);
nor U4781 (N_4781,N_4100,N_4382);
or U4782 (N_4782,N_4232,N_4055);
and U4783 (N_4783,N_4044,N_4181);
nand U4784 (N_4784,N_4363,N_4250);
and U4785 (N_4785,N_4046,N_4047);
and U4786 (N_4786,N_4353,N_4383);
and U4787 (N_4787,N_4139,N_4209);
nor U4788 (N_4788,N_4134,N_4339);
nand U4789 (N_4789,N_4119,N_4252);
xnor U4790 (N_4790,N_4453,N_4151);
nand U4791 (N_4791,N_4206,N_4385);
nor U4792 (N_4792,N_4467,N_4055);
nand U4793 (N_4793,N_4274,N_4060);
xor U4794 (N_4794,N_4106,N_4165);
or U4795 (N_4795,N_4304,N_4454);
nand U4796 (N_4796,N_4206,N_4224);
or U4797 (N_4797,N_4414,N_4162);
or U4798 (N_4798,N_4132,N_4135);
and U4799 (N_4799,N_4361,N_4182);
and U4800 (N_4800,N_4062,N_4179);
xnor U4801 (N_4801,N_4391,N_4155);
xnor U4802 (N_4802,N_4276,N_4007);
xor U4803 (N_4803,N_4153,N_4042);
xor U4804 (N_4804,N_4043,N_4300);
and U4805 (N_4805,N_4295,N_4030);
and U4806 (N_4806,N_4135,N_4279);
nand U4807 (N_4807,N_4384,N_4308);
and U4808 (N_4808,N_4485,N_4174);
nor U4809 (N_4809,N_4122,N_4496);
nor U4810 (N_4810,N_4488,N_4177);
xor U4811 (N_4811,N_4461,N_4458);
and U4812 (N_4812,N_4381,N_4494);
and U4813 (N_4813,N_4242,N_4380);
nand U4814 (N_4814,N_4045,N_4068);
nand U4815 (N_4815,N_4351,N_4483);
nor U4816 (N_4816,N_4135,N_4415);
nor U4817 (N_4817,N_4408,N_4476);
xnor U4818 (N_4818,N_4320,N_4196);
or U4819 (N_4819,N_4183,N_4440);
and U4820 (N_4820,N_4470,N_4237);
nand U4821 (N_4821,N_4175,N_4024);
nand U4822 (N_4822,N_4014,N_4082);
nor U4823 (N_4823,N_4169,N_4223);
and U4824 (N_4824,N_4430,N_4402);
xor U4825 (N_4825,N_4201,N_4120);
xor U4826 (N_4826,N_4361,N_4347);
or U4827 (N_4827,N_4166,N_4389);
xor U4828 (N_4828,N_4120,N_4495);
nor U4829 (N_4829,N_4384,N_4309);
and U4830 (N_4830,N_4273,N_4361);
and U4831 (N_4831,N_4092,N_4315);
and U4832 (N_4832,N_4413,N_4313);
nor U4833 (N_4833,N_4464,N_4360);
xnor U4834 (N_4834,N_4056,N_4184);
nand U4835 (N_4835,N_4326,N_4306);
and U4836 (N_4836,N_4217,N_4317);
nand U4837 (N_4837,N_4485,N_4127);
nand U4838 (N_4838,N_4097,N_4064);
nand U4839 (N_4839,N_4402,N_4090);
nand U4840 (N_4840,N_4466,N_4490);
and U4841 (N_4841,N_4477,N_4499);
xnor U4842 (N_4842,N_4243,N_4057);
nand U4843 (N_4843,N_4448,N_4499);
xnor U4844 (N_4844,N_4440,N_4485);
xor U4845 (N_4845,N_4185,N_4097);
xor U4846 (N_4846,N_4367,N_4269);
and U4847 (N_4847,N_4094,N_4284);
and U4848 (N_4848,N_4224,N_4257);
nor U4849 (N_4849,N_4306,N_4264);
nand U4850 (N_4850,N_4227,N_4159);
nand U4851 (N_4851,N_4236,N_4124);
or U4852 (N_4852,N_4372,N_4268);
xor U4853 (N_4853,N_4493,N_4149);
nor U4854 (N_4854,N_4168,N_4017);
or U4855 (N_4855,N_4126,N_4272);
nand U4856 (N_4856,N_4259,N_4228);
xnor U4857 (N_4857,N_4224,N_4131);
or U4858 (N_4858,N_4418,N_4153);
nand U4859 (N_4859,N_4243,N_4444);
and U4860 (N_4860,N_4023,N_4372);
nand U4861 (N_4861,N_4386,N_4117);
or U4862 (N_4862,N_4466,N_4134);
nor U4863 (N_4863,N_4330,N_4079);
or U4864 (N_4864,N_4303,N_4203);
nor U4865 (N_4865,N_4008,N_4457);
xnor U4866 (N_4866,N_4421,N_4227);
nand U4867 (N_4867,N_4444,N_4302);
nor U4868 (N_4868,N_4406,N_4103);
or U4869 (N_4869,N_4120,N_4209);
nor U4870 (N_4870,N_4362,N_4036);
nor U4871 (N_4871,N_4384,N_4041);
xnor U4872 (N_4872,N_4220,N_4275);
nor U4873 (N_4873,N_4237,N_4276);
xnor U4874 (N_4874,N_4341,N_4049);
and U4875 (N_4875,N_4095,N_4053);
or U4876 (N_4876,N_4250,N_4020);
and U4877 (N_4877,N_4497,N_4164);
nor U4878 (N_4878,N_4131,N_4154);
xor U4879 (N_4879,N_4258,N_4419);
and U4880 (N_4880,N_4016,N_4491);
nor U4881 (N_4881,N_4481,N_4238);
xor U4882 (N_4882,N_4058,N_4122);
and U4883 (N_4883,N_4299,N_4498);
or U4884 (N_4884,N_4103,N_4372);
nand U4885 (N_4885,N_4414,N_4322);
nor U4886 (N_4886,N_4451,N_4433);
nand U4887 (N_4887,N_4109,N_4144);
or U4888 (N_4888,N_4146,N_4263);
or U4889 (N_4889,N_4373,N_4214);
or U4890 (N_4890,N_4169,N_4292);
xnor U4891 (N_4891,N_4399,N_4371);
and U4892 (N_4892,N_4364,N_4114);
xor U4893 (N_4893,N_4333,N_4484);
nand U4894 (N_4894,N_4428,N_4088);
or U4895 (N_4895,N_4301,N_4492);
or U4896 (N_4896,N_4441,N_4435);
or U4897 (N_4897,N_4003,N_4193);
xnor U4898 (N_4898,N_4189,N_4332);
and U4899 (N_4899,N_4291,N_4494);
or U4900 (N_4900,N_4151,N_4253);
or U4901 (N_4901,N_4229,N_4009);
or U4902 (N_4902,N_4368,N_4495);
or U4903 (N_4903,N_4187,N_4124);
and U4904 (N_4904,N_4377,N_4370);
nor U4905 (N_4905,N_4395,N_4063);
xnor U4906 (N_4906,N_4259,N_4040);
xnor U4907 (N_4907,N_4008,N_4293);
nand U4908 (N_4908,N_4268,N_4363);
and U4909 (N_4909,N_4428,N_4198);
or U4910 (N_4910,N_4001,N_4409);
nor U4911 (N_4911,N_4414,N_4448);
nor U4912 (N_4912,N_4426,N_4490);
and U4913 (N_4913,N_4433,N_4063);
nand U4914 (N_4914,N_4088,N_4454);
nor U4915 (N_4915,N_4396,N_4319);
nor U4916 (N_4916,N_4287,N_4161);
nor U4917 (N_4917,N_4181,N_4419);
nor U4918 (N_4918,N_4009,N_4201);
nor U4919 (N_4919,N_4077,N_4413);
nand U4920 (N_4920,N_4271,N_4175);
xor U4921 (N_4921,N_4367,N_4494);
nor U4922 (N_4922,N_4133,N_4061);
xnor U4923 (N_4923,N_4227,N_4363);
nor U4924 (N_4924,N_4003,N_4322);
nand U4925 (N_4925,N_4288,N_4217);
and U4926 (N_4926,N_4239,N_4020);
or U4927 (N_4927,N_4204,N_4244);
nand U4928 (N_4928,N_4424,N_4226);
xor U4929 (N_4929,N_4393,N_4242);
and U4930 (N_4930,N_4340,N_4214);
or U4931 (N_4931,N_4178,N_4030);
nor U4932 (N_4932,N_4194,N_4363);
and U4933 (N_4933,N_4227,N_4038);
or U4934 (N_4934,N_4486,N_4206);
nand U4935 (N_4935,N_4378,N_4351);
and U4936 (N_4936,N_4037,N_4244);
nor U4937 (N_4937,N_4085,N_4377);
xor U4938 (N_4938,N_4451,N_4196);
nor U4939 (N_4939,N_4242,N_4124);
or U4940 (N_4940,N_4071,N_4323);
or U4941 (N_4941,N_4420,N_4075);
nand U4942 (N_4942,N_4319,N_4429);
xnor U4943 (N_4943,N_4159,N_4046);
nor U4944 (N_4944,N_4208,N_4379);
nor U4945 (N_4945,N_4357,N_4084);
and U4946 (N_4946,N_4487,N_4251);
xnor U4947 (N_4947,N_4233,N_4089);
xnor U4948 (N_4948,N_4224,N_4479);
and U4949 (N_4949,N_4248,N_4439);
nor U4950 (N_4950,N_4325,N_4102);
and U4951 (N_4951,N_4365,N_4439);
nand U4952 (N_4952,N_4497,N_4379);
xor U4953 (N_4953,N_4176,N_4192);
and U4954 (N_4954,N_4481,N_4077);
xor U4955 (N_4955,N_4456,N_4145);
nand U4956 (N_4956,N_4046,N_4493);
and U4957 (N_4957,N_4146,N_4343);
nor U4958 (N_4958,N_4459,N_4222);
and U4959 (N_4959,N_4119,N_4351);
nand U4960 (N_4960,N_4426,N_4039);
xnor U4961 (N_4961,N_4028,N_4407);
xor U4962 (N_4962,N_4079,N_4235);
and U4963 (N_4963,N_4208,N_4391);
or U4964 (N_4964,N_4222,N_4070);
xor U4965 (N_4965,N_4248,N_4094);
xnor U4966 (N_4966,N_4195,N_4415);
nand U4967 (N_4967,N_4454,N_4323);
xnor U4968 (N_4968,N_4036,N_4263);
and U4969 (N_4969,N_4329,N_4084);
nor U4970 (N_4970,N_4209,N_4326);
and U4971 (N_4971,N_4081,N_4327);
xor U4972 (N_4972,N_4201,N_4118);
nand U4973 (N_4973,N_4358,N_4131);
and U4974 (N_4974,N_4151,N_4273);
and U4975 (N_4975,N_4013,N_4136);
xor U4976 (N_4976,N_4440,N_4144);
nor U4977 (N_4977,N_4364,N_4362);
nand U4978 (N_4978,N_4103,N_4453);
and U4979 (N_4979,N_4074,N_4004);
nor U4980 (N_4980,N_4052,N_4262);
nand U4981 (N_4981,N_4031,N_4188);
and U4982 (N_4982,N_4299,N_4292);
xor U4983 (N_4983,N_4124,N_4194);
nor U4984 (N_4984,N_4361,N_4029);
xnor U4985 (N_4985,N_4470,N_4185);
or U4986 (N_4986,N_4254,N_4336);
xor U4987 (N_4987,N_4069,N_4157);
nor U4988 (N_4988,N_4409,N_4150);
nor U4989 (N_4989,N_4072,N_4409);
nor U4990 (N_4990,N_4152,N_4008);
and U4991 (N_4991,N_4126,N_4187);
nand U4992 (N_4992,N_4489,N_4277);
or U4993 (N_4993,N_4483,N_4246);
xor U4994 (N_4994,N_4027,N_4075);
nor U4995 (N_4995,N_4456,N_4358);
or U4996 (N_4996,N_4417,N_4326);
xnor U4997 (N_4997,N_4024,N_4247);
nor U4998 (N_4998,N_4386,N_4498);
or U4999 (N_4999,N_4063,N_4432);
and UO_0 (O_0,N_4648,N_4811);
nand UO_1 (O_1,N_4623,N_4807);
nand UO_2 (O_2,N_4637,N_4676);
or UO_3 (O_3,N_4727,N_4922);
xnor UO_4 (O_4,N_4520,N_4522);
nor UO_5 (O_5,N_4611,N_4519);
nor UO_6 (O_6,N_4548,N_4614);
and UO_7 (O_7,N_4636,N_4750);
nand UO_8 (O_8,N_4918,N_4854);
or UO_9 (O_9,N_4577,N_4670);
xnor UO_10 (O_10,N_4781,N_4579);
xor UO_11 (O_11,N_4730,N_4694);
nor UO_12 (O_12,N_4596,N_4893);
or UO_13 (O_13,N_4942,N_4860);
nor UO_14 (O_14,N_4853,N_4754);
nor UO_15 (O_15,N_4945,N_4732);
xnor UO_16 (O_16,N_4952,N_4822);
or UO_17 (O_17,N_4849,N_4783);
and UO_18 (O_18,N_4937,N_4819);
and UO_19 (O_19,N_4801,N_4746);
xnor UO_20 (O_20,N_4949,N_4588);
xnor UO_21 (O_21,N_4728,N_4525);
or UO_22 (O_22,N_4724,N_4516);
nor UO_23 (O_23,N_4573,N_4771);
nand UO_24 (O_24,N_4787,N_4718);
and UO_25 (O_25,N_4609,N_4982);
xor UO_26 (O_26,N_4967,N_4668);
xor UO_27 (O_27,N_4566,N_4810);
xnor UO_28 (O_28,N_4815,N_4890);
xor UO_29 (O_29,N_4991,N_4654);
nand UO_30 (O_30,N_4747,N_4652);
nor UO_31 (O_31,N_4719,N_4831);
xor UO_32 (O_32,N_4722,N_4758);
nor UO_33 (O_33,N_4707,N_4874);
nand UO_34 (O_34,N_4954,N_4639);
nand UO_35 (O_35,N_4714,N_4761);
or UO_36 (O_36,N_4656,N_4792);
nand UO_37 (O_37,N_4773,N_4908);
xnor UO_38 (O_38,N_4552,N_4751);
and UO_39 (O_39,N_4657,N_4524);
nor UO_40 (O_40,N_4666,N_4858);
xor UO_41 (O_41,N_4635,N_4508);
xor UO_42 (O_42,N_4843,N_4820);
nor UO_43 (O_43,N_4752,N_4593);
xor UO_44 (O_44,N_4988,N_4612);
nand UO_45 (O_45,N_4560,N_4503);
nor UO_46 (O_46,N_4550,N_4790);
nand UO_47 (O_47,N_4740,N_4586);
xor UO_48 (O_48,N_4641,N_4576);
nand UO_49 (O_49,N_4646,N_4979);
or UO_50 (O_50,N_4585,N_4613);
nand UO_51 (O_51,N_4618,N_4808);
nand UO_52 (O_52,N_4821,N_4558);
or UO_53 (O_53,N_4562,N_4650);
and UO_54 (O_54,N_4603,N_4832);
xor UO_55 (O_55,N_4805,N_4546);
or UO_56 (O_56,N_4539,N_4762);
nand UO_57 (O_57,N_4534,N_4989);
and UO_58 (O_58,N_4910,N_4532);
and UO_59 (O_59,N_4536,N_4696);
xor UO_60 (O_60,N_4658,N_4745);
nor UO_61 (O_61,N_4834,N_4911);
or UO_62 (O_62,N_4994,N_4531);
nand UO_63 (O_63,N_4768,N_4541);
nor UO_64 (O_64,N_4688,N_4863);
nand UO_65 (O_65,N_4924,N_4765);
nor UO_66 (O_66,N_4710,N_4526);
or UO_67 (O_67,N_4993,N_4594);
or UO_68 (O_68,N_4926,N_4742);
and UO_69 (O_69,N_4543,N_4659);
and UO_70 (O_70,N_4587,N_4959);
and UO_71 (O_71,N_4841,N_4735);
or UO_72 (O_72,N_4923,N_4825);
or UO_73 (O_73,N_4833,N_4749);
nand UO_74 (O_74,N_4595,N_4681);
and UO_75 (O_75,N_4788,N_4844);
nand UO_76 (O_76,N_4607,N_4604);
xnor UO_77 (O_77,N_4873,N_4794);
or UO_78 (O_78,N_4615,N_4713);
xnor UO_79 (O_79,N_4517,N_4693);
nand UO_80 (O_80,N_4624,N_4806);
nand UO_81 (O_81,N_4813,N_4680);
xnor UO_82 (O_82,N_4961,N_4877);
nand UO_83 (O_83,N_4921,N_4506);
nor UO_84 (O_84,N_4823,N_4677);
and UO_85 (O_85,N_4511,N_4699);
xor UO_86 (O_86,N_4687,N_4757);
nand UO_87 (O_87,N_4628,N_4686);
xnor UO_88 (O_88,N_4592,N_4891);
and UO_89 (O_89,N_4510,N_4563);
or UO_90 (O_90,N_4556,N_4721);
or UO_91 (O_91,N_4850,N_4675);
or UO_92 (O_92,N_4845,N_4651);
and UO_93 (O_93,N_4673,N_4917);
xor UO_94 (O_94,N_4933,N_4523);
or UO_95 (O_95,N_4990,N_4929);
or UO_96 (O_96,N_4838,N_4591);
and UO_97 (O_97,N_4928,N_4800);
or UO_98 (O_98,N_4551,N_4899);
nand UO_99 (O_99,N_4947,N_4701);
xnor UO_100 (O_100,N_4744,N_4878);
nor UO_101 (O_101,N_4887,N_4888);
or UO_102 (O_102,N_4974,N_4655);
and UO_103 (O_103,N_4868,N_4976);
nor UO_104 (O_104,N_4554,N_4698);
nand UO_105 (O_105,N_4647,N_4892);
and UO_106 (O_106,N_4502,N_4570);
xnor UO_107 (O_107,N_4764,N_4731);
nor UO_108 (O_108,N_4995,N_4900);
or UO_109 (O_109,N_4644,N_4620);
or UO_110 (O_110,N_4649,N_4785);
xor UO_111 (O_111,N_4981,N_4962);
and UO_112 (O_112,N_4784,N_4739);
or UO_113 (O_113,N_4977,N_4690);
xnor UO_114 (O_114,N_4507,N_4625);
xnor UO_115 (O_115,N_4540,N_4634);
xor UO_116 (O_116,N_4711,N_4763);
and UO_117 (O_117,N_4555,N_4683);
nor UO_118 (O_118,N_4951,N_4733);
or UO_119 (O_119,N_4786,N_4934);
or UO_120 (O_120,N_4925,N_4953);
or UO_121 (O_121,N_4549,N_4679);
nand UO_122 (O_122,N_4884,N_4606);
nor UO_123 (O_123,N_4966,N_4983);
xor UO_124 (O_124,N_4766,N_4968);
nor UO_125 (O_125,N_4817,N_4716);
and UO_126 (O_126,N_4944,N_4816);
nor UO_127 (O_127,N_4941,N_4572);
nand UO_128 (O_128,N_4671,N_4564);
nand UO_129 (O_129,N_4705,N_4880);
and UO_130 (O_130,N_4772,N_4798);
and UO_131 (O_131,N_4835,N_4969);
or UO_132 (O_132,N_4920,N_4638);
nor UO_133 (O_133,N_4793,N_4528);
xnor UO_134 (O_134,N_4725,N_4950);
nor UO_135 (O_135,N_4561,N_4987);
xnor UO_136 (O_136,N_4909,N_4774);
xnor UO_137 (O_137,N_4756,N_4857);
nor UO_138 (O_138,N_4682,N_4608);
and UO_139 (O_139,N_4667,N_4779);
or UO_140 (O_140,N_4799,N_4919);
or UO_141 (O_141,N_4978,N_4598);
nor UO_142 (O_142,N_4956,N_4915);
or UO_143 (O_143,N_4839,N_4965);
xor UO_144 (O_144,N_4963,N_4847);
nand UO_145 (O_145,N_4662,N_4697);
and UO_146 (O_146,N_4871,N_4544);
xnor UO_147 (O_147,N_4867,N_4568);
xor UO_148 (O_148,N_4580,N_4984);
or UO_149 (O_149,N_4789,N_4599);
nand UO_150 (O_150,N_4859,N_4914);
and UO_151 (O_151,N_4997,N_4939);
xor UO_152 (O_152,N_4537,N_4706);
nand UO_153 (O_153,N_4881,N_4797);
xnor UO_154 (O_154,N_4582,N_4889);
or UO_155 (O_155,N_4703,N_4814);
nand UO_156 (O_156,N_4533,N_4866);
nand UO_157 (O_157,N_4896,N_4938);
nor UO_158 (O_158,N_4743,N_4804);
nor UO_159 (O_159,N_4770,N_4795);
nand UO_160 (O_160,N_4842,N_4569);
or UO_161 (O_161,N_4824,N_4898);
nor UO_162 (O_162,N_4848,N_4943);
and UO_163 (O_163,N_4940,N_4729);
xnor UO_164 (O_164,N_4791,N_4741);
or UO_165 (O_165,N_4907,N_4960);
or UO_166 (O_166,N_4602,N_4509);
and UO_167 (O_167,N_4700,N_4678);
xnor UO_168 (O_168,N_4557,N_4830);
nand UO_169 (O_169,N_4759,N_4643);
and UO_170 (O_170,N_4894,N_4882);
nand UO_171 (O_171,N_4574,N_4616);
xnor UO_172 (O_172,N_4685,N_4916);
nand UO_173 (O_173,N_4930,N_4975);
xor UO_174 (O_174,N_4645,N_4672);
and UO_175 (O_175,N_4617,N_4684);
and UO_176 (O_176,N_4674,N_4876);
xor UO_177 (O_177,N_4948,N_4905);
nor UO_178 (O_178,N_4664,N_4778);
xnor UO_179 (O_179,N_4521,N_4970);
xnor UO_180 (O_180,N_4559,N_4583);
xor UO_181 (O_181,N_4836,N_4957);
xnor UO_182 (O_182,N_4903,N_4753);
and UO_183 (O_183,N_4633,N_4581);
xor UO_184 (O_184,N_4665,N_4955);
and UO_185 (O_185,N_4709,N_4883);
or UO_186 (O_186,N_4865,N_4870);
nor UO_187 (O_187,N_4998,N_4973);
or UO_188 (O_188,N_4972,N_4780);
nand UO_189 (O_189,N_4964,N_4738);
nand UO_190 (O_190,N_4627,N_4547);
and UO_191 (O_191,N_4708,N_4601);
xnor UO_192 (O_192,N_4632,N_4837);
and UO_193 (O_193,N_4885,N_4912);
nand UO_194 (O_194,N_4589,N_4663);
and UO_195 (O_195,N_4980,N_4913);
nor UO_196 (O_196,N_4971,N_4518);
nor UO_197 (O_197,N_4535,N_4567);
nand UO_198 (O_198,N_4906,N_4512);
nor UO_199 (O_199,N_4864,N_4600);
nand UO_200 (O_200,N_4875,N_4584);
or UO_201 (O_201,N_4886,N_4902);
or UO_202 (O_202,N_4545,N_4695);
xnor UO_203 (O_203,N_4840,N_4852);
or UO_204 (O_204,N_4605,N_4737);
or UO_205 (O_205,N_4529,N_4897);
nand UO_206 (O_206,N_4515,N_4769);
nand UO_207 (O_207,N_4640,N_4826);
xnor UO_208 (O_208,N_4931,N_4879);
nand UO_209 (O_209,N_4935,N_4828);
and UO_210 (O_210,N_4755,N_4775);
nand UO_211 (O_211,N_4872,N_4527);
and UO_212 (O_212,N_4565,N_4985);
nor UO_213 (O_213,N_4501,N_4514);
or UO_214 (O_214,N_4861,N_4829);
xor UO_215 (O_215,N_4715,N_4777);
nand UO_216 (O_216,N_4631,N_4704);
or UO_217 (O_217,N_4856,N_4702);
nor UO_218 (O_218,N_4610,N_4530);
nand UO_219 (O_219,N_4927,N_4999);
xnor UO_220 (O_220,N_4736,N_4622);
nand UO_221 (O_221,N_4575,N_4803);
nor UO_222 (O_222,N_4653,N_4660);
or UO_223 (O_223,N_4796,N_4851);
nand UO_224 (O_224,N_4827,N_4691);
xor UO_225 (O_225,N_4689,N_4869);
and UO_226 (O_226,N_4500,N_4712);
or UO_227 (O_227,N_4542,N_4642);
and UO_228 (O_228,N_4597,N_4629);
nand UO_229 (O_229,N_4590,N_4513);
or UO_230 (O_230,N_4932,N_4986);
or UO_231 (O_231,N_4996,N_4782);
xor UO_232 (O_232,N_4661,N_4626);
nor UO_233 (O_233,N_4717,N_4630);
nand UO_234 (O_234,N_4992,N_4818);
xor UO_235 (O_235,N_4776,N_4619);
xnor UO_236 (O_236,N_4901,N_4862);
nor UO_237 (O_237,N_4505,N_4846);
nor UO_238 (O_238,N_4904,N_4855);
xor UO_239 (O_239,N_4895,N_4553);
xnor UO_240 (O_240,N_4748,N_4946);
xor UO_241 (O_241,N_4809,N_4621);
and UO_242 (O_242,N_4723,N_4571);
xnor UO_243 (O_243,N_4692,N_4812);
and UO_244 (O_244,N_4669,N_4767);
and UO_245 (O_245,N_4734,N_4578);
and UO_246 (O_246,N_4958,N_4538);
nor UO_247 (O_247,N_4802,N_4720);
or UO_248 (O_248,N_4504,N_4936);
or UO_249 (O_249,N_4760,N_4726);
nor UO_250 (O_250,N_4883,N_4734);
xnor UO_251 (O_251,N_4865,N_4527);
nor UO_252 (O_252,N_4575,N_4751);
nand UO_253 (O_253,N_4642,N_4655);
nand UO_254 (O_254,N_4747,N_4756);
xor UO_255 (O_255,N_4584,N_4701);
xor UO_256 (O_256,N_4883,N_4752);
or UO_257 (O_257,N_4811,N_4619);
and UO_258 (O_258,N_4752,N_4660);
and UO_259 (O_259,N_4872,N_4846);
and UO_260 (O_260,N_4685,N_4810);
nor UO_261 (O_261,N_4558,N_4833);
and UO_262 (O_262,N_4851,N_4664);
and UO_263 (O_263,N_4944,N_4557);
nand UO_264 (O_264,N_4583,N_4882);
or UO_265 (O_265,N_4802,N_4729);
and UO_266 (O_266,N_4752,N_4539);
xnor UO_267 (O_267,N_4972,N_4509);
nand UO_268 (O_268,N_4540,N_4742);
nor UO_269 (O_269,N_4616,N_4893);
or UO_270 (O_270,N_4513,N_4867);
xor UO_271 (O_271,N_4511,N_4755);
nor UO_272 (O_272,N_4547,N_4598);
xnor UO_273 (O_273,N_4576,N_4811);
xor UO_274 (O_274,N_4695,N_4857);
and UO_275 (O_275,N_4959,N_4547);
or UO_276 (O_276,N_4768,N_4910);
nor UO_277 (O_277,N_4847,N_4671);
or UO_278 (O_278,N_4662,N_4560);
xor UO_279 (O_279,N_4505,N_4867);
xor UO_280 (O_280,N_4774,N_4715);
xor UO_281 (O_281,N_4666,N_4520);
nand UO_282 (O_282,N_4812,N_4680);
nand UO_283 (O_283,N_4602,N_4886);
nor UO_284 (O_284,N_4652,N_4693);
xnor UO_285 (O_285,N_4955,N_4509);
xnor UO_286 (O_286,N_4625,N_4653);
nand UO_287 (O_287,N_4954,N_4649);
xor UO_288 (O_288,N_4759,N_4574);
nand UO_289 (O_289,N_4910,N_4675);
or UO_290 (O_290,N_4671,N_4628);
xor UO_291 (O_291,N_4597,N_4797);
nand UO_292 (O_292,N_4740,N_4513);
or UO_293 (O_293,N_4738,N_4899);
and UO_294 (O_294,N_4515,N_4619);
and UO_295 (O_295,N_4662,N_4728);
or UO_296 (O_296,N_4689,N_4873);
and UO_297 (O_297,N_4925,N_4659);
xnor UO_298 (O_298,N_4973,N_4634);
xnor UO_299 (O_299,N_4985,N_4530);
xor UO_300 (O_300,N_4918,N_4882);
nor UO_301 (O_301,N_4828,N_4721);
xor UO_302 (O_302,N_4973,N_4551);
or UO_303 (O_303,N_4885,N_4597);
xor UO_304 (O_304,N_4526,N_4696);
nand UO_305 (O_305,N_4863,N_4618);
nor UO_306 (O_306,N_4560,N_4701);
and UO_307 (O_307,N_4731,N_4726);
and UO_308 (O_308,N_4939,N_4597);
xnor UO_309 (O_309,N_4743,N_4810);
or UO_310 (O_310,N_4546,N_4640);
nand UO_311 (O_311,N_4807,N_4865);
nand UO_312 (O_312,N_4872,N_4501);
and UO_313 (O_313,N_4633,N_4527);
nand UO_314 (O_314,N_4619,N_4683);
nand UO_315 (O_315,N_4964,N_4549);
and UO_316 (O_316,N_4604,N_4901);
or UO_317 (O_317,N_4677,N_4944);
nor UO_318 (O_318,N_4720,N_4925);
nor UO_319 (O_319,N_4976,N_4714);
nand UO_320 (O_320,N_4731,N_4943);
nand UO_321 (O_321,N_4968,N_4980);
nor UO_322 (O_322,N_4888,N_4965);
nor UO_323 (O_323,N_4718,N_4902);
and UO_324 (O_324,N_4998,N_4663);
or UO_325 (O_325,N_4846,N_4754);
nor UO_326 (O_326,N_4735,N_4503);
and UO_327 (O_327,N_4936,N_4841);
and UO_328 (O_328,N_4982,N_4874);
or UO_329 (O_329,N_4683,N_4881);
or UO_330 (O_330,N_4616,N_4592);
nand UO_331 (O_331,N_4970,N_4617);
and UO_332 (O_332,N_4786,N_4505);
nand UO_333 (O_333,N_4605,N_4858);
xnor UO_334 (O_334,N_4576,N_4580);
xor UO_335 (O_335,N_4956,N_4686);
nor UO_336 (O_336,N_4548,N_4717);
or UO_337 (O_337,N_4564,N_4979);
xor UO_338 (O_338,N_4715,N_4766);
xnor UO_339 (O_339,N_4541,N_4986);
xor UO_340 (O_340,N_4687,N_4588);
nand UO_341 (O_341,N_4508,N_4633);
nor UO_342 (O_342,N_4632,N_4652);
nor UO_343 (O_343,N_4857,N_4874);
or UO_344 (O_344,N_4676,N_4666);
nand UO_345 (O_345,N_4581,N_4513);
and UO_346 (O_346,N_4839,N_4665);
nor UO_347 (O_347,N_4917,N_4944);
and UO_348 (O_348,N_4590,N_4682);
and UO_349 (O_349,N_4644,N_4616);
and UO_350 (O_350,N_4658,N_4756);
or UO_351 (O_351,N_4513,N_4511);
or UO_352 (O_352,N_4740,N_4894);
nand UO_353 (O_353,N_4686,N_4734);
nor UO_354 (O_354,N_4824,N_4593);
nor UO_355 (O_355,N_4857,N_4513);
nor UO_356 (O_356,N_4707,N_4755);
or UO_357 (O_357,N_4870,N_4767);
nand UO_358 (O_358,N_4773,N_4641);
nor UO_359 (O_359,N_4845,N_4929);
xnor UO_360 (O_360,N_4639,N_4562);
xnor UO_361 (O_361,N_4615,N_4921);
nand UO_362 (O_362,N_4598,N_4559);
or UO_363 (O_363,N_4765,N_4992);
or UO_364 (O_364,N_4922,N_4730);
nor UO_365 (O_365,N_4985,N_4877);
and UO_366 (O_366,N_4797,N_4869);
nor UO_367 (O_367,N_4793,N_4530);
nor UO_368 (O_368,N_4862,N_4983);
or UO_369 (O_369,N_4545,N_4630);
xnor UO_370 (O_370,N_4822,N_4507);
nor UO_371 (O_371,N_4714,N_4688);
and UO_372 (O_372,N_4587,N_4784);
nor UO_373 (O_373,N_4634,N_4982);
xor UO_374 (O_374,N_4668,N_4645);
xor UO_375 (O_375,N_4949,N_4763);
xor UO_376 (O_376,N_4797,N_4784);
nand UO_377 (O_377,N_4569,N_4595);
or UO_378 (O_378,N_4567,N_4637);
nand UO_379 (O_379,N_4733,N_4868);
and UO_380 (O_380,N_4786,N_4501);
and UO_381 (O_381,N_4666,N_4541);
and UO_382 (O_382,N_4752,N_4766);
nand UO_383 (O_383,N_4843,N_4534);
nor UO_384 (O_384,N_4689,N_4921);
nand UO_385 (O_385,N_4893,N_4833);
nand UO_386 (O_386,N_4591,N_4561);
nor UO_387 (O_387,N_4991,N_4634);
and UO_388 (O_388,N_4890,N_4512);
xnor UO_389 (O_389,N_4884,N_4874);
and UO_390 (O_390,N_4546,N_4680);
and UO_391 (O_391,N_4755,N_4615);
or UO_392 (O_392,N_4849,N_4658);
and UO_393 (O_393,N_4945,N_4604);
xnor UO_394 (O_394,N_4746,N_4567);
or UO_395 (O_395,N_4941,N_4769);
or UO_396 (O_396,N_4748,N_4685);
nor UO_397 (O_397,N_4783,N_4510);
or UO_398 (O_398,N_4876,N_4652);
and UO_399 (O_399,N_4675,N_4572);
nand UO_400 (O_400,N_4844,N_4905);
or UO_401 (O_401,N_4854,N_4824);
or UO_402 (O_402,N_4693,N_4935);
xor UO_403 (O_403,N_4914,N_4621);
xnor UO_404 (O_404,N_4605,N_4991);
nand UO_405 (O_405,N_4867,N_4665);
or UO_406 (O_406,N_4525,N_4565);
nor UO_407 (O_407,N_4616,N_4786);
xnor UO_408 (O_408,N_4557,N_4553);
xor UO_409 (O_409,N_4906,N_4789);
nand UO_410 (O_410,N_4561,N_4813);
xor UO_411 (O_411,N_4668,N_4946);
nor UO_412 (O_412,N_4797,N_4862);
xor UO_413 (O_413,N_4937,N_4531);
or UO_414 (O_414,N_4983,N_4809);
nor UO_415 (O_415,N_4823,N_4826);
and UO_416 (O_416,N_4641,N_4958);
nand UO_417 (O_417,N_4580,N_4533);
or UO_418 (O_418,N_4717,N_4761);
or UO_419 (O_419,N_4872,N_4671);
nand UO_420 (O_420,N_4507,N_4823);
or UO_421 (O_421,N_4521,N_4943);
nand UO_422 (O_422,N_4717,N_4887);
or UO_423 (O_423,N_4721,N_4699);
nand UO_424 (O_424,N_4925,N_4892);
or UO_425 (O_425,N_4625,N_4704);
or UO_426 (O_426,N_4903,N_4931);
xor UO_427 (O_427,N_4955,N_4510);
nand UO_428 (O_428,N_4687,N_4750);
and UO_429 (O_429,N_4524,N_4652);
and UO_430 (O_430,N_4961,N_4980);
or UO_431 (O_431,N_4742,N_4639);
and UO_432 (O_432,N_4714,N_4890);
nor UO_433 (O_433,N_4900,N_4880);
nor UO_434 (O_434,N_4673,N_4832);
or UO_435 (O_435,N_4841,N_4502);
and UO_436 (O_436,N_4889,N_4898);
or UO_437 (O_437,N_4729,N_4722);
and UO_438 (O_438,N_4855,N_4556);
xnor UO_439 (O_439,N_4886,N_4638);
nand UO_440 (O_440,N_4662,N_4827);
and UO_441 (O_441,N_4618,N_4609);
xnor UO_442 (O_442,N_4792,N_4556);
xnor UO_443 (O_443,N_4676,N_4882);
or UO_444 (O_444,N_4515,N_4906);
nor UO_445 (O_445,N_4743,N_4744);
nand UO_446 (O_446,N_4689,N_4714);
nand UO_447 (O_447,N_4935,N_4502);
or UO_448 (O_448,N_4679,N_4822);
or UO_449 (O_449,N_4905,N_4779);
xnor UO_450 (O_450,N_4504,N_4594);
xor UO_451 (O_451,N_4522,N_4640);
and UO_452 (O_452,N_4879,N_4751);
and UO_453 (O_453,N_4820,N_4534);
xnor UO_454 (O_454,N_4744,N_4857);
or UO_455 (O_455,N_4657,N_4850);
or UO_456 (O_456,N_4965,N_4533);
nor UO_457 (O_457,N_4561,N_4727);
or UO_458 (O_458,N_4688,N_4929);
or UO_459 (O_459,N_4919,N_4653);
nor UO_460 (O_460,N_4556,N_4649);
and UO_461 (O_461,N_4894,N_4518);
nand UO_462 (O_462,N_4946,N_4595);
or UO_463 (O_463,N_4783,N_4708);
xor UO_464 (O_464,N_4612,N_4516);
nand UO_465 (O_465,N_4904,N_4736);
nor UO_466 (O_466,N_4967,N_4812);
nand UO_467 (O_467,N_4870,N_4629);
nor UO_468 (O_468,N_4588,N_4688);
nand UO_469 (O_469,N_4674,N_4843);
xor UO_470 (O_470,N_4534,N_4911);
xnor UO_471 (O_471,N_4826,N_4540);
and UO_472 (O_472,N_4911,N_4709);
nor UO_473 (O_473,N_4907,N_4606);
or UO_474 (O_474,N_4581,N_4731);
nand UO_475 (O_475,N_4724,N_4554);
or UO_476 (O_476,N_4870,N_4974);
or UO_477 (O_477,N_4543,N_4685);
or UO_478 (O_478,N_4623,N_4990);
and UO_479 (O_479,N_4827,N_4745);
and UO_480 (O_480,N_4916,N_4878);
xnor UO_481 (O_481,N_4764,N_4807);
and UO_482 (O_482,N_4649,N_4610);
nor UO_483 (O_483,N_4939,N_4569);
nor UO_484 (O_484,N_4511,N_4529);
nor UO_485 (O_485,N_4750,N_4923);
or UO_486 (O_486,N_4981,N_4834);
nor UO_487 (O_487,N_4755,N_4963);
nand UO_488 (O_488,N_4840,N_4936);
and UO_489 (O_489,N_4837,N_4738);
xnor UO_490 (O_490,N_4861,N_4952);
nand UO_491 (O_491,N_4590,N_4915);
nor UO_492 (O_492,N_4656,N_4534);
or UO_493 (O_493,N_4665,N_4623);
xnor UO_494 (O_494,N_4863,N_4708);
or UO_495 (O_495,N_4669,N_4665);
nand UO_496 (O_496,N_4907,N_4992);
or UO_497 (O_497,N_4692,N_4565);
xnor UO_498 (O_498,N_4537,N_4758);
xnor UO_499 (O_499,N_4594,N_4780);
nand UO_500 (O_500,N_4790,N_4838);
nor UO_501 (O_501,N_4679,N_4513);
or UO_502 (O_502,N_4796,N_4872);
nand UO_503 (O_503,N_4661,N_4531);
nand UO_504 (O_504,N_4797,N_4515);
or UO_505 (O_505,N_4848,N_4803);
or UO_506 (O_506,N_4641,N_4750);
or UO_507 (O_507,N_4943,N_4835);
and UO_508 (O_508,N_4700,N_4605);
xnor UO_509 (O_509,N_4692,N_4534);
nor UO_510 (O_510,N_4711,N_4929);
xor UO_511 (O_511,N_4811,N_4522);
xor UO_512 (O_512,N_4794,N_4757);
or UO_513 (O_513,N_4503,N_4703);
nand UO_514 (O_514,N_4734,N_4887);
nand UO_515 (O_515,N_4531,N_4993);
nand UO_516 (O_516,N_4916,N_4711);
xor UO_517 (O_517,N_4931,N_4564);
xor UO_518 (O_518,N_4854,N_4993);
or UO_519 (O_519,N_4987,N_4861);
xnor UO_520 (O_520,N_4560,N_4616);
nand UO_521 (O_521,N_4727,N_4620);
or UO_522 (O_522,N_4641,N_4670);
xor UO_523 (O_523,N_4516,N_4985);
nor UO_524 (O_524,N_4854,N_4722);
or UO_525 (O_525,N_4861,N_4795);
nand UO_526 (O_526,N_4949,N_4753);
nor UO_527 (O_527,N_4877,N_4620);
nor UO_528 (O_528,N_4677,N_4979);
nor UO_529 (O_529,N_4526,N_4562);
xnor UO_530 (O_530,N_4923,N_4770);
and UO_531 (O_531,N_4983,N_4969);
nand UO_532 (O_532,N_4787,N_4826);
and UO_533 (O_533,N_4771,N_4821);
and UO_534 (O_534,N_4945,N_4927);
nor UO_535 (O_535,N_4741,N_4841);
nor UO_536 (O_536,N_4646,N_4937);
or UO_537 (O_537,N_4741,N_4734);
nor UO_538 (O_538,N_4565,N_4573);
xnor UO_539 (O_539,N_4907,N_4880);
nand UO_540 (O_540,N_4637,N_4719);
nor UO_541 (O_541,N_4932,N_4935);
nor UO_542 (O_542,N_4633,N_4841);
nand UO_543 (O_543,N_4862,N_4722);
nand UO_544 (O_544,N_4765,N_4908);
nor UO_545 (O_545,N_4795,N_4527);
or UO_546 (O_546,N_4713,N_4566);
and UO_547 (O_547,N_4860,N_4821);
and UO_548 (O_548,N_4682,N_4551);
nor UO_549 (O_549,N_4617,N_4959);
nand UO_550 (O_550,N_4706,N_4508);
and UO_551 (O_551,N_4913,N_4905);
or UO_552 (O_552,N_4530,N_4643);
and UO_553 (O_553,N_4719,N_4755);
xor UO_554 (O_554,N_4760,N_4516);
and UO_555 (O_555,N_4592,N_4848);
nand UO_556 (O_556,N_4996,N_4642);
nor UO_557 (O_557,N_4901,N_4800);
xnor UO_558 (O_558,N_4773,N_4668);
nor UO_559 (O_559,N_4575,N_4968);
nor UO_560 (O_560,N_4613,N_4817);
nor UO_561 (O_561,N_4659,N_4737);
or UO_562 (O_562,N_4558,N_4988);
nand UO_563 (O_563,N_4672,N_4799);
xor UO_564 (O_564,N_4524,N_4765);
nand UO_565 (O_565,N_4523,N_4944);
xnor UO_566 (O_566,N_4895,N_4747);
xnor UO_567 (O_567,N_4580,N_4975);
or UO_568 (O_568,N_4986,N_4935);
nand UO_569 (O_569,N_4640,N_4648);
and UO_570 (O_570,N_4939,N_4760);
and UO_571 (O_571,N_4934,N_4847);
xor UO_572 (O_572,N_4604,N_4574);
nand UO_573 (O_573,N_4569,N_4809);
xor UO_574 (O_574,N_4568,N_4790);
nand UO_575 (O_575,N_4513,N_4926);
and UO_576 (O_576,N_4876,N_4797);
xor UO_577 (O_577,N_4822,N_4908);
xor UO_578 (O_578,N_4716,N_4904);
and UO_579 (O_579,N_4542,N_4628);
nand UO_580 (O_580,N_4756,N_4930);
and UO_581 (O_581,N_4974,N_4988);
nor UO_582 (O_582,N_4606,N_4715);
xor UO_583 (O_583,N_4603,N_4655);
or UO_584 (O_584,N_4553,N_4736);
nor UO_585 (O_585,N_4845,N_4932);
or UO_586 (O_586,N_4524,N_4799);
nand UO_587 (O_587,N_4893,N_4673);
or UO_588 (O_588,N_4862,N_4919);
and UO_589 (O_589,N_4824,N_4682);
and UO_590 (O_590,N_4964,N_4654);
or UO_591 (O_591,N_4772,N_4750);
xnor UO_592 (O_592,N_4740,N_4767);
or UO_593 (O_593,N_4666,N_4837);
nor UO_594 (O_594,N_4516,N_4586);
xnor UO_595 (O_595,N_4741,N_4773);
and UO_596 (O_596,N_4970,N_4701);
or UO_597 (O_597,N_4842,N_4824);
xor UO_598 (O_598,N_4988,N_4683);
xnor UO_599 (O_599,N_4827,N_4550);
nand UO_600 (O_600,N_4833,N_4661);
nor UO_601 (O_601,N_4629,N_4918);
and UO_602 (O_602,N_4856,N_4638);
and UO_603 (O_603,N_4648,N_4873);
xnor UO_604 (O_604,N_4968,N_4872);
xor UO_605 (O_605,N_4741,N_4788);
nor UO_606 (O_606,N_4536,N_4524);
nand UO_607 (O_607,N_4954,N_4613);
xnor UO_608 (O_608,N_4675,N_4826);
or UO_609 (O_609,N_4864,N_4739);
nand UO_610 (O_610,N_4864,N_4894);
nor UO_611 (O_611,N_4664,N_4759);
or UO_612 (O_612,N_4936,N_4861);
or UO_613 (O_613,N_4597,N_4582);
nor UO_614 (O_614,N_4814,N_4506);
xnor UO_615 (O_615,N_4958,N_4956);
xnor UO_616 (O_616,N_4658,N_4525);
nor UO_617 (O_617,N_4566,N_4947);
xor UO_618 (O_618,N_4685,N_4998);
or UO_619 (O_619,N_4854,N_4991);
xor UO_620 (O_620,N_4616,N_4844);
nor UO_621 (O_621,N_4516,N_4633);
or UO_622 (O_622,N_4622,N_4621);
nor UO_623 (O_623,N_4559,N_4989);
or UO_624 (O_624,N_4593,N_4724);
xnor UO_625 (O_625,N_4600,N_4869);
nand UO_626 (O_626,N_4993,N_4675);
or UO_627 (O_627,N_4759,N_4573);
nand UO_628 (O_628,N_4802,N_4857);
and UO_629 (O_629,N_4848,N_4890);
xnor UO_630 (O_630,N_4931,N_4670);
and UO_631 (O_631,N_4692,N_4949);
xor UO_632 (O_632,N_4708,N_4786);
and UO_633 (O_633,N_4861,N_4713);
nor UO_634 (O_634,N_4822,N_4766);
nor UO_635 (O_635,N_4710,N_4633);
xor UO_636 (O_636,N_4803,N_4669);
or UO_637 (O_637,N_4911,N_4896);
nor UO_638 (O_638,N_4984,N_4518);
xor UO_639 (O_639,N_4599,N_4990);
nor UO_640 (O_640,N_4830,N_4789);
and UO_641 (O_641,N_4811,N_4506);
xor UO_642 (O_642,N_4885,N_4690);
nor UO_643 (O_643,N_4974,N_4720);
nand UO_644 (O_644,N_4768,N_4526);
or UO_645 (O_645,N_4611,N_4576);
xnor UO_646 (O_646,N_4797,N_4828);
nor UO_647 (O_647,N_4593,N_4704);
nor UO_648 (O_648,N_4644,N_4935);
nor UO_649 (O_649,N_4708,N_4778);
or UO_650 (O_650,N_4501,N_4643);
nor UO_651 (O_651,N_4683,N_4688);
nor UO_652 (O_652,N_4526,N_4632);
and UO_653 (O_653,N_4924,N_4889);
and UO_654 (O_654,N_4790,N_4697);
nand UO_655 (O_655,N_4513,N_4610);
and UO_656 (O_656,N_4591,N_4545);
or UO_657 (O_657,N_4963,N_4536);
nor UO_658 (O_658,N_4820,N_4866);
nor UO_659 (O_659,N_4979,N_4996);
xor UO_660 (O_660,N_4944,N_4774);
nand UO_661 (O_661,N_4836,N_4841);
and UO_662 (O_662,N_4898,N_4949);
xor UO_663 (O_663,N_4714,N_4985);
nor UO_664 (O_664,N_4540,N_4822);
xnor UO_665 (O_665,N_4616,N_4962);
xnor UO_666 (O_666,N_4655,N_4746);
and UO_667 (O_667,N_4598,N_4557);
or UO_668 (O_668,N_4824,N_4503);
nor UO_669 (O_669,N_4633,N_4997);
or UO_670 (O_670,N_4709,N_4604);
nor UO_671 (O_671,N_4738,N_4737);
or UO_672 (O_672,N_4541,N_4599);
and UO_673 (O_673,N_4958,N_4784);
or UO_674 (O_674,N_4513,N_4654);
nor UO_675 (O_675,N_4925,N_4924);
nand UO_676 (O_676,N_4937,N_4855);
xnor UO_677 (O_677,N_4747,N_4944);
or UO_678 (O_678,N_4958,N_4886);
and UO_679 (O_679,N_4785,N_4584);
nand UO_680 (O_680,N_4818,N_4664);
nor UO_681 (O_681,N_4569,N_4950);
nand UO_682 (O_682,N_4516,N_4504);
nor UO_683 (O_683,N_4806,N_4640);
xor UO_684 (O_684,N_4576,N_4583);
or UO_685 (O_685,N_4623,N_4849);
xnor UO_686 (O_686,N_4731,N_4639);
nand UO_687 (O_687,N_4676,N_4786);
xnor UO_688 (O_688,N_4844,N_4631);
nand UO_689 (O_689,N_4852,N_4950);
nand UO_690 (O_690,N_4516,N_4530);
and UO_691 (O_691,N_4569,N_4801);
xor UO_692 (O_692,N_4548,N_4792);
and UO_693 (O_693,N_4788,N_4790);
and UO_694 (O_694,N_4933,N_4682);
nor UO_695 (O_695,N_4854,N_4965);
xnor UO_696 (O_696,N_4583,N_4702);
xor UO_697 (O_697,N_4743,N_4775);
or UO_698 (O_698,N_4727,N_4596);
and UO_699 (O_699,N_4719,N_4738);
xor UO_700 (O_700,N_4883,N_4919);
xor UO_701 (O_701,N_4749,N_4817);
and UO_702 (O_702,N_4695,N_4647);
and UO_703 (O_703,N_4897,N_4744);
nor UO_704 (O_704,N_4885,N_4775);
and UO_705 (O_705,N_4661,N_4812);
and UO_706 (O_706,N_4737,N_4951);
or UO_707 (O_707,N_4989,N_4580);
and UO_708 (O_708,N_4719,N_4777);
nor UO_709 (O_709,N_4612,N_4509);
nor UO_710 (O_710,N_4808,N_4901);
xor UO_711 (O_711,N_4705,N_4871);
nand UO_712 (O_712,N_4530,N_4722);
or UO_713 (O_713,N_4768,N_4669);
and UO_714 (O_714,N_4878,N_4680);
or UO_715 (O_715,N_4966,N_4642);
nand UO_716 (O_716,N_4876,N_4528);
and UO_717 (O_717,N_4728,N_4614);
xnor UO_718 (O_718,N_4886,N_4795);
or UO_719 (O_719,N_4757,N_4776);
and UO_720 (O_720,N_4511,N_4708);
xor UO_721 (O_721,N_4973,N_4520);
nor UO_722 (O_722,N_4916,N_4665);
and UO_723 (O_723,N_4946,N_4788);
nor UO_724 (O_724,N_4949,N_4694);
or UO_725 (O_725,N_4796,N_4631);
or UO_726 (O_726,N_4662,N_4932);
and UO_727 (O_727,N_4576,N_4520);
xor UO_728 (O_728,N_4838,N_4871);
nand UO_729 (O_729,N_4826,N_4653);
nand UO_730 (O_730,N_4593,N_4741);
or UO_731 (O_731,N_4725,N_4631);
xnor UO_732 (O_732,N_4668,N_4731);
or UO_733 (O_733,N_4738,N_4644);
xor UO_734 (O_734,N_4738,N_4518);
or UO_735 (O_735,N_4582,N_4807);
xor UO_736 (O_736,N_4827,N_4697);
xor UO_737 (O_737,N_4612,N_4976);
or UO_738 (O_738,N_4605,N_4750);
or UO_739 (O_739,N_4857,N_4698);
xnor UO_740 (O_740,N_4816,N_4657);
and UO_741 (O_741,N_4741,N_4798);
xor UO_742 (O_742,N_4858,N_4930);
nand UO_743 (O_743,N_4962,N_4708);
xnor UO_744 (O_744,N_4966,N_4844);
nor UO_745 (O_745,N_4685,N_4537);
and UO_746 (O_746,N_4940,N_4636);
nand UO_747 (O_747,N_4521,N_4650);
nand UO_748 (O_748,N_4957,N_4558);
nand UO_749 (O_749,N_4853,N_4633);
nand UO_750 (O_750,N_4651,N_4743);
or UO_751 (O_751,N_4996,N_4828);
or UO_752 (O_752,N_4753,N_4927);
nor UO_753 (O_753,N_4949,N_4985);
or UO_754 (O_754,N_4723,N_4977);
or UO_755 (O_755,N_4629,N_4527);
and UO_756 (O_756,N_4920,N_4943);
nor UO_757 (O_757,N_4956,N_4838);
xor UO_758 (O_758,N_4682,N_4806);
xor UO_759 (O_759,N_4910,N_4697);
nor UO_760 (O_760,N_4517,N_4928);
and UO_761 (O_761,N_4901,N_4993);
nor UO_762 (O_762,N_4672,N_4768);
nor UO_763 (O_763,N_4610,N_4795);
or UO_764 (O_764,N_4545,N_4511);
or UO_765 (O_765,N_4741,N_4727);
xnor UO_766 (O_766,N_4974,N_4764);
or UO_767 (O_767,N_4586,N_4869);
or UO_768 (O_768,N_4536,N_4931);
or UO_769 (O_769,N_4830,N_4746);
nor UO_770 (O_770,N_4950,N_4658);
nor UO_771 (O_771,N_4502,N_4922);
nor UO_772 (O_772,N_4952,N_4617);
or UO_773 (O_773,N_4982,N_4944);
nor UO_774 (O_774,N_4707,N_4832);
and UO_775 (O_775,N_4896,N_4525);
and UO_776 (O_776,N_4769,N_4857);
xnor UO_777 (O_777,N_4861,N_4831);
or UO_778 (O_778,N_4576,N_4813);
or UO_779 (O_779,N_4513,N_4886);
xor UO_780 (O_780,N_4896,N_4839);
nor UO_781 (O_781,N_4916,N_4533);
or UO_782 (O_782,N_4625,N_4548);
nand UO_783 (O_783,N_4838,N_4821);
nor UO_784 (O_784,N_4716,N_4886);
nand UO_785 (O_785,N_4872,N_4621);
or UO_786 (O_786,N_4541,N_4634);
and UO_787 (O_787,N_4890,N_4520);
nand UO_788 (O_788,N_4611,N_4973);
or UO_789 (O_789,N_4834,N_4892);
xnor UO_790 (O_790,N_4948,N_4655);
and UO_791 (O_791,N_4625,N_4813);
nor UO_792 (O_792,N_4545,N_4586);
nand UO_793 (O_793,N_4932,N_4771);
xor UO_794 (O_794,N_4621,N_4602);
or UO_795 (O_795,N_4685,N_4922);
nor UO_796 (O_796,N_4930,N_4535);
or UO_797 (O_797,N_4727,N_4591);
nor UO_798 (O_798,N_4731,N_4585);
nand UO_799 (O_799,N_4720,N_4573);
xor UO_800 (O_800,N_4726,N_4555);
and UO_801 (O_801,N_4636,N_4923);
nand UO_802 (O_802,N_4775,N_4835);
and UO_803 (O_803,N_4827,N_4985);
nand UO_804 (O_804,N_4608,N_4975);
nand UO_805 (O_805,N_4584,N_4709);
or UO_806 (O_806,N_4661,N_4697);
or UO_807 (O_807,N_4648,N_4901);
nand UO_808 (O_808,N_4795,N_4809);
nor UO_809 (O_809,N_4813,N_4607);
and UO_810 (O_810,N_4679,N_4751);
and UO_811 (O_811,N_4819,N_4933);
xor UO_812 (O_812,N_4641,N_4603);
xnor UO_813 (O_813,N_4715,N_4611);
or UO_814 (O_814,N_4746,N_4908);
xor UO_815 (O_815,N_4576,N_4861);
nand UO_816 (O_816,N_4828,N_4501);
or UO_817 (O_817,N_4535,N_4768);
nor UO_818 (O_818,N_4859,N_4770);
or UO_819 (O_819,N_4739,N_4922);
xnor UO_820 (O_820,N_4526,N_4734);
and UO_821 (O_821,N_4729,N_4688);
or UO_822 (O_822,N_4701,N_4923);
or UO_823 (O_823,N_4957,N_4605);
nor UO_824 (O_824,N_4900,N_4516);
xnor UO_825 (O_825,N_4732,N_4626);
and UO_826 (O_826,N_4690,N_4623);
or UO_827 (O_827,N_4707,N_4699);
or UO_828 (O_828,N_4641,N_4596);
and UO_829 (O_829,N_4560,N_4683);
nand UO_830 (O_830,N_4730,N_4803);
or UO_831 (O_831,N_4943,N_4967);
xnor UO_832 (O_832,N_4882,N_4960);
nor UO_833 (O_833,N_4566,N_4637);
nand UO_834 (O_834,N_4939,N_4728);
xnor UO_835 (O_835,N_4641,N_4743);
nand UO_836 (O_836,N_4844,N_4782);
or UO_837 (O_837,N_4914,N_4804);
nand UO_838 (O_838,N_4810,N_4655);
nand UO_839 (O_839,N_4522,N_4796);
nor UO_840 (O_840,N_4761,N_4786);
xor UO_841 (O_841,N_4567,N_4983);
nand UO_842 (O_842,N_4998,N_4541);
xor UO_843 (O_843,N_4991,N_4665);
or UO_844 (O_844,N_4976,N_4700);
and UO_845 (O_845,N_4864,N_4839);
or UO_846 (O_846,N_4991,N_4843);
nor UO_847 (O_847,N_4756,N_4758);
and UO_848 (O_848,N_4603,N_4622);
or UO_849 (O_849,N_4924,N_4572);
and UO_850 (O_850,N_4935,N_4737);
xnor UO_851 (O_851,N_4634,N_4898);
xnor UO_852 (O_852,N_4731,N_4537);
and UO_853 (O_853,N_4885,N_4849);
and UO_854 (O_854,N_4980,N_4669);
nor UO_855 (O_855,N_4785,N_4520);
xnor UO_856 (O_856,N_4689,N_4737);
nand UO_857 (O_857,N_4701,N_4615);
and UO_858 (O_858,N_4871,N_4663);
xnor UO_859 (O_859,N_4711,N_4787);
nor UO_860 (O_860,N_4738,N_4923);
and UO_861 (O_861,N_4624,N_4920);
nand UO_862 (O_862,N_4510,N_4932);
xnor UO_863 (O_863,N_4597,N_4679);
and UO_864 (O_864,N_4979,N_4593);
nor UO_865 (O_865,N_4573,N_4803);
nor UO_866 (O_866,N_4811,N_4692);
nand UO_867 (O_867,N_4809,N_4779);
nor UO_868 (O_868,N_4628,N_4858);
xnor UO_869 (O_869,N_4933,N_4518);
or UO_870 (O_870,N_4553,N_4826);
nand UO_871 (O_871,N_4967,N_4745);
or UO_872 (O_872,N_4540,N_4627);
and UO_873 (O_873,N_4977,N_4974);
or UO_874 (O_874,N_4723,N_4532);
or UO_875 (O_875,N_4991,N_4938);
and UO_876 (O_876,N_4514,N_4546);
or UO_877 (O_877,N_4672,N_4729);
or UO_878 (O_878,N_4760,N_4764);
xor UO_879 (O_879,N_4864,N_4715);
xnor UO_880 (O_880,N_4805,N_4596);
nor UO_881 (O_881,N_4510,N_4893);
and UO_882 (O_882,N_4524,N_4530);
or UO_883 (O_883,N_4858,N_4791);
or UO_884 (O_884,N_4542,N_4961);
xnor UO_885 (O_885,N_4707,N_4691);
xor UO_886 (O_886,N_4521,N_4987);
nor UO_887 (O_887,N_4656,N_4678);
or UO_888 (O_888,N_4764,N_4501);
nor UO_889 (O_889,N_4632,N_4860);
nand UO_890 (O_890,N_4666,N_4776);
or UO_891 (O_891,N_4856,N_4724);
or UO_892 (O_892,N_4665,N_4660);
nor UO_893 (O_893,N_4831,N_4559);
nor UO_894 (O_894,N_4776,N_4508);
nor UO_895 (O_895,N_4858,N_4937);
or UO_896 (O_896,N_4721,N_4516);
nand UO_897 (O_897,N_4528,N_4860);
xnor UO_898 (O_898,N_4731,N_4684);
xnor UO_899 (O_899,N_4847,N_4775);
or UO_900 (O_900,N_4695,N_4569);
and UO_901 (O_901,N_4671,N_4565);
nor UO_902 (O_902,N_4610,N_4963);
xor UO_903 (O_903,N_4704,N_4678);
nand UO_904 (O_904,N_4663,N_4869);
nor UO_905 (O_905,N_4660,N_4563);
nor UO_906 (O_906,N_4510,N_4552);
nand UO_907 (O_907,N_4632,N_4646);
nand UO_908 (O_908,N_4889,N_4550);
or UO_909 (O_909,N_4759,N_4719);
nand UO_910 (O_910,N_4707,N_4891);
xnor UO_911 (O_911,N_4886,N_4937);
and UO_912 (O_912,N_4607,N_4868);
nand UO_913 (O_913,N_4980,N_4826);
nand UO_914 (O_914,N_4749,N_4737);
xnor UO_915 (O_915,N_4874,N_4681);
nor UO_916 (O_916,N_4603,N_4789);
or UO_917 (O_917,N_4946,N_4933);
or UO_918 (O_918,N_4975,N_4687);
nor UO_919 (O_919,N_4908,N_4504);
or UO_920 (O_920,N_4946,N_4613);
and UO_921 (O_921,N_4801,N_4719);
or UO_922 (O_922,N_4539,N_4657);
or UO_923 (O_923,N_4784,N_4708);
or UO_924 (O_924,N_4825,N_4771);
xnor UO_925 (O_925,N_4933,N_4642);
nand UO_926 (O_926,N_4592,N_4504);
nand UO_927 (O_927,N_4763,N_4671);
and UO_928 (O_928,N_4735,N_4720);
or UO_929 (O_929,N_4934,N_4770);
xor UO_930 (O_930,N_4616,N_4627);
nand UO_931 (O_931,N_4512,N_4893);
xnor UO_932 (O_932,N_4729,N_4742);
nand UO_933 (O_933,N_4585,N_4755);
and UO_934 (O_934,N_4906,N_4713);
and UO_935 (O_935,N_4844,N_4674);
nand UO_936 (O_936,N_4509,N_4988);
nor UO_937 (O_937,N_4745,N_4778);
and UO_938 (O_938,N_4583,N_4859);
nor UO_939 (O_939,N_4539,N_4644);
nor UO_940 (O_940,N_4548,N_4559);
xnor UO_941 (O_941,N_4614,N_4771);
nand UO_942 (O_942,N_4862,N_4534);
nand UO_943 (O_943,N_4592,N_4963);
nand UO_944 (O_944,N_4985,N_4707);
nand UO_945 (O_945,N_4807,N_4749);
nor UO_946 (O_946,N_4961,N_4740);
and UO_947 (O_947,N_4571,N_4768);
nand UO_948 (O_948,N_4944,N_4525);
or UO_949 (O_949,N_4996,N_4690);
and UO_950 (O_950,N_4984,N_4623);
nor UO_951 (O_951,N_4856,N_4886);
nand UO_952 (O_952,N_4792,N_4964);
nor UO_953 (O_953,N_4601,N_4701);
or UO_954 (O_954,N_4872,N_4865);
xnor UO_955 (O_955,N_4548,N_4876);
nor UO_956 (O_956,N_4942,N_4540);
nand UO_957 (O_957,N_4586,N_4604);
and UO_958 (O_958,N_4709,N_4560);
or UO_959 (O_959,N_4828,N_4705);
nor UO_960 (O_960,N_4972,N_4565);
nand UO_961 (O_961,N_4591,N_4758);
and UO_962 (O_962,N_4691,N_4532);
or UO_963 (O_963,N_4813,N_4719);
or UO_964 (O_964,N_4674,N_4782);
and UO_965 (O_965,N_4629,N_4951);
nand UO_966 (O_966,N_4722,N_4831);
xnor UO_967 (O_967,N_4558,N_4765);
nor UO_968 (O_968,N_4782,N_4861);
xnor UO_969 (O_969,N_4547,N_4541);
or UO_970 (O_970,N_4968,N_4871);
or UO_971 (O_971,N_4921,N_4736);
nand UO_972 (O_972,N_4892,N_4526);
nand UO_973 (O_973,N_4808,N_4955);
xor UO_974 (O_974,N_4757,N_4591);
nand UO_975 (O_975,N_4570,N_4568);
xor UO_976 (O_976,N_4535,N_4503);
or UO_977 (O_977,N_4527,N_4528);
and UO_978 (O_978,N_4978,N_4953);
or UO_979 (O_979,N_4988,N_4987);
and UO_980 (O_980,N_4939,N_4853);
xnor UO_981 (O_981,N_4827,N_4705);
nand UO_982 (O_982,N_4959,N_4522);
nor UO_983 (O_983,N_4860,N_4789);
and UO_984 (O_984,N_4681,N_4792);
nand UO_985 (O_985,N_4603,N_4708);
xnor UO_986 (O_986,N_4705,N_4591);
and UO_987 (O_987,N_4883,N_4783);
and UO_988 (O_988,N_4519,N_4938);
nor UO_989 (O_989,N_4817,N_4567);
and UO_990 (O_990,N_4925,N_4962);
nor UO_991 (O_991,N_4837,N_4818);
and UO_992 (O_992,N_4778,N_4513);
xor UO_993 (O_993,N_4977,N_4800);
nor UO_994 (O_994,N_4944,N_4999);
nand UO_995 (O_995,N_4760,N_4945);
nor UO_996 (O_996,N_4606,N_4802);
nor UO_997 (O_997,N_4671,N_4655);
or UO_998 (O_998,N_4514,N_4549);
and UO_999 (O_999,N_4585,N_4720);
endmodule