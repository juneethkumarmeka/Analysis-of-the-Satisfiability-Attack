module basic_2500_25000_3000_10_levels_1xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_1864,In_397);
nor U1 (N_1,In_2092,In_1869);
nand U2 (N_2,In_962,In_2016);
and U3 (N_3,In_1513,In_690);
or U4 (N_4,In_225,In_1371);
and U5 (N_5,In_1730,In_1650);
and U6 (N_6,In_266,In_971);
or U7 (N_7,In_2177,In_1305);
or U8 (N_8,In_929,In_1937);
and U9 (N_9,In_226,In_1638);
nand U10 (N_10,In_1161,In_240);
nor U11 (N_11,In_1091,In_2326);
nor U12 (N_12,In_2347,In_2135);
nor U13 (N_13,In_1659,In_370);
or U14 (N_14,In_374,In_1732);
nor U15 (N_15,In_783,In_2007);
nand U16 (N_16,In_100,In_1183);
or U17 (N_17,In_1539,In_1466);
or U18 (N_18,In_1546,In_1706);
or U19 (N_19,In_1278,In_1609);
nand U20 (N_20,In_1023,In_277);
and U21 (N_21,In_221,In_2172);
or U22 (N_22,In_2445,In_585);
nand U23 (N_23,In_259,In_711);
or U24 (N_24,In_981,In_1399);
or U25 (N_25,In_2272,In_2428);
or U26 (N_26,In_1890,In_338);
nand U27 (N_27,In_552,In_562);
nand U28 (N_28,In_373,In_1345);
or U29 (N_29,In_747,In_748);
nand U30 (N_30,In_1806,In_1655);
nand U31 (N_31,In_601,In_671);
xnor U32 (N_32,In_1042,In_120);
and U33 (N_33,In_2478,In_1716);
nor U34 (N_34,In_2076,In_1497);
or U35 (N_35,In_1179,In_459);
or U36 (N_36,In_368,In_1772);
or U37 (N_37,In_996,In_1576);
nor U38 (N_38,In_464,In_1290);
nand U39 (N_39,In_1435,In_1191);
and U40 (N_40,In_1571,In_1248);
nand U41 (N_41,In_2382,In_251);
nor U42 (N_42,In_1250,In_43);
nand U43 (N_43,In_1858,In_1383);
xnor U44 (N_44,In_175,In_124);
or U45 (N_45,In_36,In_2063);
and U46 (N_46,In_1851,In_2417);
or U47 (N_47,In_219,In_188);
or U48 (N_48,In_1284,In_1657);
or U49 (N_49,In_1620,In_183);
nor U50 (N_50,In_1796,In_692);
or U51 (N_51,In_1781,In_2137);
or U52 (N_52,In_454,In_730);
or U53 (N_53,In_2247,In_233);
nand U54 (N_54,In_1619,In_1985);
nor U55 (N_55,In_2253,In_1264);
or U56 (N_56,In_1591,In_56);
or U57 (N_57,In_384,In_2388);
nor U58 (N_58,In_1164,In_1564);
or U59 (N_59,In_32,In_1963);
nor U60 (N_60,In_1559,In_1681);
and U61 (N_61,In_903,In_1477);
and U62 (N_62,In_2334,In_1958);
or U63 (N_63,In_631,In_1319);
nor U64 (N_64,In_2472,In_2147);
or U65 (N_65,In_656,In_2165);
and U66 (N_66,In_223,In_1334);
nor U67 (N_67,In_1308,In_639);
nor U68 (N_68,In_1240,In_1063);
and U69 (N_69,In_797,In_13);
and U70 (N_70,In_1606,In_1805);
nand U71 (N_71,In_1004,In_289);
or U72 (N_72,In_621,In_1432);
nor U73 (N_73,In_589,In_1346);
nor U74 (N_74,In_130,In_1569);
nor U75 (N_75,In_1793,In_238);
or U76 (N_76,In_295,In_1932);
or U77 (N_77,In_1670,In_2364);
or U78 (N_78,In_2006,In_791);
and U79 (N_79,In_1203,In_1131);
nor U80 (N_80,In_307,In_779);
nor U81 (N_81,In_1975,In_2050);
and U82 (N_82,In_1066,In_170);
nor U83 (N_83,In_1364,In_2127);
or U84 (N_84,In_570,In_157);
and U85 (N_85,In_1133,In_1615);
or U86 (N_86,In_1162,In_2237);
nor U87 (N_87,In_495,In_1763);
and U88 (N_88,In_2228,In_1443);
nor U89 (N_89,In_1385,In_992);
nand U90 (N_90,In_2318,In_1007);
nand U91 (N_91,In_342,In_1151);
or U92 (N_92,In_990,In_960);
nor U93 (N_93,In_818,In_148);
and U94 (N_94,In_1511,In_719);
nand U95 (N_95,In_152,In_54);
nor U96 (N_96,In_921,In_2460);
or U97 (N_97,In_574,In_1704);
or U98 (N_98,In_239,In_389);
nor U99 (N_99,In_1418,In_1515);
nand U100 (N_100,In_624,In_1033);
or U101 (N_101,In_407,In_61);
nor U102 (N_102,In_2216,In_242);
and U103 (N_103,In_683,In_1724);
nand U104 (N_104,In_1981,In_1922);
nand U105 (N_105,In_109,In_1380);
nand U106 (N_106,In_1524,In_1617);
or U107 (N_107,In_1697,In_1865);
nor U108 (N_108,In_1715,In_198);
or U109 (N_109,In_288,In_619);
nand U110 (N_110,In_846,In_2363);
nor U111 (N_111,In_1895,In_1901);
or U112 (N_112,In_1542,In_1229);
and U113 (N_113,In_1573,In_670);
and U114 (N_114,In_2110,In_97);
nor U115 (N_115,In_1288,In_1748);
or U116 (N_116,In_667,In_1430);
and U117 (N_117,In_1834,In_1351);
nand U118 (N_118,In_2181,In_1253);
nand U119 (N_119,In_83,In_2391);
nand U120 (N_120,In_2360,In_2011);
or U121 (N_121,In_1123,In_1701);
nor U122 (N_122,In_1084,In_1882);
or U123 (N_123,In_39,In_880);
nor U124 (N_124,In_1487,In_1);
nand U125 (N_125,In_1787,In_526);
and U126 (N_126,In_1832,In_73);
nand U127 (N_127,In_882,In_432);
and U128 (N_128,In_972,In_901);
and U129 (N_129,In_1900,In_2134);
or U130 (N_130,In_914,In_916);
or U131 (N_131,In_1077,In_2190);
nor U132 (N_132,In_2107,In_125);
nand U133 (N_133,In_2257,In_1983);
nand U134 (N_134,In_1098,In_2030);
nor U135 (N_135,In_1978,In_227);
and U136 (N_136,In_1809,In_2087);
nand U137 (N_137,In_1570,In_1794);
or U138 (N_138,In_773,In_387);
or U139 (N_139,In_792,In_1790);
nor U140 (N_140,In_1829,In_2234);
or U141 (N_141,In_1441,In_272);
nand U142 (N_142,In_69,In_1445);
nor U143 (N_143,In_2071,In_948);
and U144 (N_144,In_2383,In_2402);
nor U145 (N_145,In_451,In_287);
or U146 (N_146,In_320,In_1109);
and U147 (N_147,In_807,In_34);
nand U148 (N_148,In_2200,In_367);
nand U149 (N_149,In_1447,In_231);
nor U150 (N_150,In_560,In_1255);
or U151 (N_151,In_2404,In_1930);
nand U152 (N_152,In_1647,In_1977);
nor U153 (N_153,In_1625,In_1616);
nand U154 (N_154,In_1957,In_164);
nand U155 (N_155,In_991,In_1299);
nor U156 (N_156,In_510,In_2466);
or U157 (N_157,In_472,In_733);
or U158 (N_158,In_1982,In_2225);
and U159 (N_159,In_923,In_1686);
nor U160 (N_160,In_2311,In_1661);
and U161 (N_161,In_486,In_2273);
nand U162 (N_162,In_1674,In_1744);
nor U163 (N_163,In_98,In_2343);
nand U164 (N_164,In_2114,In_86);
nor U165 (N_165,In_870,In_831);
or U166 (N_166,In_662,In_892);
and U167 (N_167,In_2152,In_1537);
nand U168 (N_168,In_162,In_1948);
nor U169 (N_169,In_1106,In_2043);
and U170 (N_170,In_1283,In_1685);
nor U171 (N_171,In_2124,In_1516);
nor U172 (N_172,In_197,In_610);
or U173 (N_173,In_1672,In_160);
nor U174 (N_174,In_720,In_550);
or U175 (N_175,In_1618,In_84);
or U176 (N_176,In_1665,In_1044);
and U177 (N_177,In_1700,In_246);
and U178 (N_178,In_524,In_2157);
or U179 (N_179,In_1262,In_902);
nand U180 (N_180,In_814,In_134);
and U181 (N_181,In_952,In_825);
or U182 (N_182,In_268,In_2297);
nor U183 (N_183,In_504,In_1558);
nand U184 (N_184,In_1773,In_493);
nand U185 (N_185,In_715,In_412);
nor U186 (N_186,In_2299,In_2375);
nand U187 (N_187,In_1759,In_453);
nor U188 (N_188,In_81,In_1074);
nor U189 (N_189,In_2229,In_1272);
or U190 (N_190,In_523,In_563);
or U191 (N_191,In_1354,In_2386);
nor U192 (N_192,In_1145,In_1696);
nor U193 (N_193,In_1816,In_508);
nor U194 (N_194,In_638,In_1928);
nand U195 (N_195,In_1879,In_2132);
nand U196 (N_196,In_1608,In_2);
and U197 (N_197,In_885,In_520);
or U198 (N_198,In_1104,In_806);
or U199 (N_199,In_2487,In_1636);
nor U200 (N_200,In_2396,In_2118);
nand U201 (N_201,In_1518,In_1118);
or U202 (N_202,In_2119,In_1474);
or U203 (N_203,In_444,In_995);
nand U204 (N_204,In_1215,In_1398);
and U205 (N_205,In_1968,In_385);
and U206 (N_206,In_851,In_2056);
nor U207 (N_207,In_1753,In_1552);
nor U208 (N_208,In_2395,In_271);
nand U209 (N_209,In_993,In_2091);
nor U210 (N_210,In_703,In_1875);
nor U211 (N_211,In_787,In_729);
or U212 (N_212,In_299,In_1232);
nand U213 (N_213,In_2032,In_2207);
nand U214 (N_214,In_1989,In_429);
and U215 (N_215,In_745,In_1810);
nor U216 (N_216,In_297,In_2268);
nor U217 (N_217,In_1596,In_376);
or U218 (N_218,In_1874,In_1973);
and U219 (N_219,In_2451,In_2389);
nor U220 (N_220,In_717,In_2325);
or U221 (N_221,In_150,In_980);
and U222 (N_222,In_114,In_1916);
nor U223 (N_223,In_666,In_1111);
nand U224 (N_224,In_616,In_1572);
and U225 (N_225,In_635,In_131);
nor U226 (N_226,In_313,In_2185);
nor U227 (N_227,In_1312,In_153);
or U228 (N_228,In_1872,In_461);
or U229 (N_229,In_55,In_1610);
and U230 (N_230,In_538,In_1330);
or U231 (N_231,In_2488,In_2312);
nor U232 (N_232,In_201,In_1999);
nor U233 (N_233,In_516,In_534);
nor U234 (N_234,In_127,In_1757);
nor U235 (N_235,In_539,In_2085);
and U236 (N_236,In_784,In_1736);
or U237 (N_237,In_2189,In_1451);
nand U238 (N_238,In_2427,In_680);
and U239 (N_239,In_191,In_326);
or U240 (N_240,In_819,In_2143);
or U241 (N_241,In_2133,In_2154);
and U242 (N_242,In_2010,In_1483);
nand U243 (N_243,In_1835,In_613);
xnor U244 (N_244,In_840,In_1208);
nor U245 (N_245,In_1538,In_1194);
or U246 (N_246,In_2463,In_304);
and U247 (N_247,In_2204,In_1413);
or U248 (N_248,In_1857,In_741);
nand U249 (N_249,In_281,In_132);
nor U250 (N_250,In_1406,In_1000);
and U251 (N_251,In_1574,In_884);
and U252 (N_252,In_859,In_190);
nand U253 (N_253,In_1940,In_1603);
nor U254 (N_254,In_2289,In_2102);
nand U255 (N_255,In_1493,In_1236);
and U256 (N_256,In_1517,In_2313);
nand U257 (N_257,In_9,In_408);
and U258 (N_258,In_514,In_1219);
nand U259 (N_259,In_1627,In_1450);
and U260 (N_260,In_1138,In_30);
nand U261 (N_261,In_1465,In_509);
nand U262 (N_262,In_310,In_1951);
nor U263 (N_263,In_1727,In_1070);
nor U264 (N_264,In_323,In_511);
nand U265 (N_265,In_536,In_1935);
nand U266 (N_266,In_2298,In_1011);
and U267 (N_267,In_2150,In_1801);
nor U268 (N_268,In_1101,In_2418);
nor U269 (N_269,In_1550,In_581);
or U270 (N_270,In_2355,In_1494);
nand U271 (N_271,In_1257,In_260);
or U272 (N_272,In_1306,In_2285);
xnor U273 (N_273,In_2014,In_1231);
nand U274 (N_274,In_1268,In_890);
nor U275 (N_275,In_11,In_1235);
or U276 (N_276,In_928,In_87);
nor U277 (N_277,In_702,In_1047);
and U278 (N_278,In_1291,In_2286);
nand U279 (N_279,In_1313,In_177);
nor U280 (N_280,In_2049,In_742);
nor U281 (N_281,In_1375,In_1397);
and U282 (N_282,In_2136,In_1854);
and U283 (N_283,In_518,In_426);
nor U284 (N_284,In_2483,In_835);
or U285 (N_285,In_2038,In_2155);
or U286 (N_286,In_77,In_2479);
nand U287 (N_287,In_52,In_433);
or U288 (N_288,In_448,In_126);
or U289 (N_289,In_2354,In_1143);
nand U290 (N_290,In_1277,In_1522);
nor U291 (N_291,In_1448,In_1863);
nor U292 (N_292,In_2057,In_1745);
and U293 (N_293,In_668,In_1648);
nand U294 (N_294,In_2405,In_1357);
nor U295 (N_295,In_920,In_1839);
nand U296 (N_296,In_1592,In_1640);
nor U297 (N_297,In_490,In_1234);
nand U298 (N_298,In_1961,In_2440);
or U299 (N_299,In_2142,In_2276);
nor U300 (N_300,In_909,In_1969);
xnor U301 (N_301,In_521,In_1327);
nor U302 (N_302,In_2371,In_1153);
nor U303 (N_303,In_1919,In_1896);
nand U304 (N_304,In_1034,In_123);
nor U305 (N_305,In_826,In_1256);
nand U306 (N_306,In_1274,In_634);
or U307 (N_307,In_643,In_476);
and U308 (N_308,In_2464,In_1669);
nor U309 (N_309,In_1386,In_1915);
nor U310 (N_310,In_1423,In_1035);
or U311 (N_311,In_70,In_193);
xnor U312 (N_312,In_2351,In_1452);
or U313 (N_313,In_2446,In_2040);
or U314 (N_314,In_1113,In_161);
or U315 (N_315,In_793,In_1006);
or U316 (N_316,In_894,In_630);
nor U317 (N_317,In_1032,In_595);
nand U318 (N_318,In_2356,In_1988);
and U319 (N_319,In_1979,In_1280);
and U320 (N_320,In_1873,In_2481);
or U321 (N_321,In_1583,In_984);
and U322 (N_322,In_414,In_652);
or U323 (N_323,In_2047,In_422);
nand U324 (N_324,In_2473,In_1238);
nor U325 (N_325,In_383,In_942);
nand U326 (N_326,In_1827,In_1929);
nand U327 (N_327,In_1960,In_1848);
nor U328 (N_328,In_1742,In_1623);
or U329 (N_329,In_258,In_1944);
and U330 (N_330,In_1843,In_839);
or U331 (N_331,In_889,In_2455);
nor U332 (N_332,In_1218,In_2384);
and U333 (N_333,In_381,In_1883);
nor U334 (N_334,In_1938,In_1720);
nor U335 (N_335,In_1855,In_1422);
and U336 (N_336,In_21,In_1712);
or U337 (N_337,In_1764,In_1769);
nand U338 (N_338,In_1927,In_12);
and U339 (N_339,In_1575,In_1393);
or U340 (N_340,In_1404,In_485);
and U341 (N_341,In_76,In_2103);
and U342 (N_342,In_2274,In_1693);
nand U343 (N_343,In_28,In_480);
or U344 (N_344,In_722,In_2227);
nand U345 (N_345,In_1714,In_1633);
or U346 (N_346,In_1867,In_419);
nor U347 (N_347,In_1076,In_2453);
and U348 (N_348,In_2240,In_1970);
nor U349 (N_349,In_2302,In_762);
or U350 (N_350,In_1318,In_2097);
nand U351 (N_351,In_663,In_1439);
or U352 (N_352,In_1285,In_274);
nand U353 (N_353,In_554,In_20);
or U354 (N_354,In_1239,In_1156);
and U355 (N_355,In_1329,In_2209);
nor U356 (N_356,In_107,In_1590);
and U357 (N_357,In_973,In_1136);
nand U358 (N_358,In_1557,In_915);
nor U359 (N_359,In_1389,In_1949);
or U360 (N_360,In_1196,In_405);
nand U361 (N_361,In_1833,In_2376);
and U362 (N_362,In_640,In_1335);
nand U363 (N_363,In_2116,In_887);
and U364 (N_364,In_802,In_700);
and U365 (N_365,In_2020,In_2176);
and U366 (N_366,In_592,In_515);
nand U367 (N_367,In_1130,In_632);
and U368 (N_368,In_2146,In_2160);
nor U369 (N_369,In_473,In_404);
nor U370 (N_370,In_140,In_232);
and U371 (N_371,In_2018,In_89);
and U372 (N_372,In_388,In_1826);
or U373 (N_373,In_2454,In_1582);
nand U374 (N_374,In_1519,In_675);
nor U375 (N_375,In_1824,In_857);
nor U376 (N_376,In_596,In_2490);
xnor U377 (N_377,In_1611,In_401);
and U378 (N_378,In_2013,In_2284);
or U379 (N_379,In_1918,In_2443);
and U380 (N_380,In_1342,In_1946);
nand U381 (N_381,In_1222,In_608);
and U382 (N_382,In_1129,In_540);
nand U383 (N_383,In_881,In_533);
and U384 (N_384,In_1103,In_1456);
nor U385 (N_385,In_2084,In_757);
or U386 (N_386,In_1225,In_1767);
nor U387 (N_387,In_1967,In_760);
nor U388 (N_388,In_910,In_415);
nand U389 (N_389,In_1770,In_349);
and U390 (N_390,In_1671,In_1437);
and U391 (N_391,In_2476,In_1749);
and U392 (N_392,In_471,In_1293);
nor U393 (N_393,In_2075,In_2264);
or U394 (N_394,In_1039,In_1015);
or U395 (N_395,In_2163,In_458);
and U396 (N_396,In_559,In_63);
and U397 (N_397,In_1260,In_185);
or U398 (N_398,In_1626,In_1237);
and U399 (N_399,In_1069,In_254);
or U400 (N_400,In_1026,In_1534);
nor U401 (N_401,In_1921,In_128);
xnor U402 (N_402,In_208,In_2290);
and U403 (N_403,In_1217,In_2497);
or U404 (N_404,In_364,In_450);
nor U405 (N_405,In_424,In_2051);
nand U406 (N_406,In_979,In_2361);
nor U407 (N_407,In_617,In_1054);
nand U408 (N_408,In_936,In_462);
nor U409 (N_409,In_2438,In_1602);
or U410 (N_410,In_1458,In_1726);
nor U411 (N_411,In_1295,In_333);
and U412 (N_412,In_525,In_598);
or U413 (N_413,In_1001,In_1838);
nor U414 (N_414,In_241,In_2205);
or U415 (N_415,In_328,In_347);
or U416 (N_416,In_35,In_1646);
or U417 (N_417,In_1190,In_314);
nor U418 (N_418,In_824,In_174);
nor U419 (N_419,In_2482,In_312);
and U420 (N_420,In_869,In_2230);
nor U421 (N_421,In_1666,In_138);
or U422 (N_422,In_2241,In_877);
or U423 (N_423,In_2309,In_1897);
nand U424 (N_424,In_2465,In_1475);
nor U425 (N_425,In_15,In_1544);
and U426 (N_426,In_1529,In_113);
nor U427 (N_427,In_586,In_82);
or U428 (N_428,In_2235,In_2031);
nand U429 (N_429,In_1316,In_1504);
nor U430 (N_430,In_576,In_940);
nor U431 (N_431,In_360,In_119);
nand U432 (N_432,In_1642,In_1846);
nand U433 (N_433,In_1003,In_265);
and U434 (N_434,In_2278,In_315);
nand U435 (N_435,In_2198,In_1349);
nand U436 (N_436,In_336,In_1741);
or U437 (N_437,In_409,In_532);
and U438 (N_438,In_758,In_772);
and U439 (N_439,In_1689,In_529);
and U440 (N_440,In_676,In_205);
nand U441 (N_441,In_1792,In_1783);
nand U442 (N_442,In_755,In_122);
or U443 (N_443,In_431,In_1321);
nand U444 (N_444,In_214,In_457);
or U445 (N_445,In_737,In_1024);
nand U446 (N_446,In_445,In_1990);
and U447 (N_447,In_2158,In_1269);
xnor U448 (N_448,In_1680,In_832);
and U449 (N_449,In_446,In_1579);
or U450 (N_450,In_256,In_398);
nand U451 (N_451,In_568,In_939);
and U452 (N_452,In_479,In_1859);
nand U453 (N_453,In_19,In_1333);
nor U454 (N_454,In_1678,In_1547);
nand U455 (N_455,In_1812,In_1514);
nand U456 (N_456,In_217,In_1739);
or U457 (N_457,In_830,In_842);
or U458 (N_458,In_1980,In_1079);
nand U459 (N_459,In_146,In_2022);
nand U460 (N_460,In_925,In_1473);
nor U461 (N_461,In_544,In_1315);
nand U462 (N_462,In_606,In_994);
or U463 (N_463,In_513,In_121);
and U464 (N_464,In_1297,In_2183);
or U465 (N_465,In_1431,In_449);
and U466 (N_466,In_1540,In_911);
and U467 (N_467,In_1841,In_2288);
nand U468 (N_468,In_660,In_474);
nor U469 (N_469,In_1703,In_611);
nor U470 (N_470,In_2421,In_924);
and U471 (N_471,In_1226,In_1141);
nand U472 (N_472,In_1391,In_1907);
nand U473 (N_473,In_1411,In_1852);
or U474 (N_474,In_2109,In_584);
nand U475 (N_475,In_477,In_466);
nor U476 (N_476,In_2435,In_1180);
or U477 (N_477,In_305,In_2162);
nand U478 (N_478,In_764,In_1267);
and U479 (N_479,In_402,In_1148);
nand U480 (N_480,In_1762,In_578);
nor U481 (N_481,In_329,In_961);
nand U482 (N_482,In_337,In_1067);
nor U483 (N_483,In_2398,In_1994);
nand U484 (N_484,In_341,In_956);
and U485 (N_485,In_2457,In_2104);
nor U486 (N_486,In_1728,In_1566);
xor U487 (N_487,In_917,In_3);
and U488 (N_488,In_1709,In_1228);
nor U489 (N_489,In_1014,In_603);
and U490 (N_490,In_951,In_2002);
or U491 (N_491,In_1630,In_1362);
nor U492 (N_492,In_1637,In_224);
nand U493 (N_493,In_2046,In_1690);
and U494 (N_494,In_235,In_535);
or U495 (N_495,In_423,In_1056);
nor U496 (N_496,In_2399,In_1193);
nor U497 (N_497,In_1213,In_350);
nor U498 (N_498,In_2180,In_1811);
and U499 (N_499,In_487,In_59);
or U500 (N_500,In_905,In_798);
and U501 (N_501,In_853,In_1013);
nor U502 (N_502,In_1581,In_1653);
nor U503 (N_503,In_196,In_580);
nor U504 (N_504,In_2098,In_2432);
nand U505 (N_505,In_352,In_937);
nor U506 (N_506,In_1292,In_332);
nand U507 (N_507,In_657,In_1645);
nor U508 (N_508,In_800,In_2462);
and U509 (N_509,In_58,In_99);
or U510 (N_510,In_2159,In_1005);
nand U511 (N_511,In_1296,In_967);
and U512 (N_512,In_263,In_1395);
and U513 (N_513,In_2221,In_1045);
and U514 (N_514,In_276,In_2425);
and U515 (N_515,In_1503,In_1607);
and U516 (N_516,In_2436,In_1541);
and U517 (N_517,In_117,In_2292);
and U518 (N_518,In_1998,In_843);
nand U519 (N_519,In_1055,In_1365);
or U520 (N_520,In_421,In_605);
nand U521 (N_521,In_1556,In_1083);
nand U522 (N_522,In_456,In_1825);
and U523 (N_523,In_1945,In_2251);
nor U524 (N_524,In_2077,In_180);
or U525 (N_525,In_1107,In_249);
nand U526 (N_526,In_173,In_1830);
and U527 (N_527,In_854,In_2359);
or U528 (N_528,In_2308,In_2217);
nand U529 (N_529,In_2148,In_1894);
nor U530 (N_530,In_1476,In_5);
or U531 (N_531,In_1100,In_1181);
and U532 (N_532,In_655,In_1172);
nor U533 (N_533,In_597,In_618);
or U534 (N_534,In_1481,In_1797);
nand U535 (N_535,In_751,In_1382);
and U536 (N_536,In_803,In_2452);
nor U537 (N_537,In_873,In_858);
nand U538 (N_538,In_2414,In_904);
nor U539 (N_539,In_2449,In_2305);
nand U540 (N_540,In_2362,In_1303);
and U541 (N_541,In_2317,In_844);
or U542 (N_542,In_2271,In_1102);
nor U543 (N_543,In_2263,In_96);
or U544 (N_544,In_182,In_105);
and U545 (N_545,In_2044,In_1040);
nor U546 (N_546,In_496,In_1245);
nand U547 (N_547,In_575,In_253);
nor U548 (N_548,In_665,In_2331);
nor U549 (N_549,In_1710,In_306);
and U550 (N_550,In_855,In_2173);
or U551 (N_551,In_2083,In_2301);
or U552 (N_552,In_1523,In_348);
nand U553 (N_553,In_2495,In_2105);
nor U554 (N_554,In_2053,In_1247);
or U555 (N_555,In_2260,In_2036);
nor U556 (N_556,In_142,In_1876);
nand U557 (N_557,In_1071,In_2416);
nor U558 (N_558,In_1317,In_1495);
or U559 (N_559,In_1807,In_1986);
nor U560 (N_560,In_878,In_796);
or U561 (N_561,In_736,In_944);
or U562 (N_562,In_2471,In_1964);
or U563 (N_563,In_1146,In_2408);
nand U564 (N_564,In_363,In_704);
or U565 (N_565,In_200,In_726);
xnor U566 (N_566,In_1030,In_252);
nand U567 (N_567,In_187,In_1307);
nor U568 (N_568,In_677,In_66);
nand U569 (N_569,In_1604,In_1567);
nand U570 (N_570,In_2339,In_434);
nor U571 (N_571,In_2149,In_759);
or U572 (N_572,In_2210,In_1018);
or U573 (N_573,In_1535,In_1729);
and U574 (N_574,In_926,In_1294);
nand U575 (N_575,In_1584,In_502);
and U576 (N_576,In_294,In_2485);
nand U577 (N_577,In_2059,In_522);
or U578 (N_578,In_1713,In_647);
or U579 (N_579,In_2277,In_1880);
nand U580 (N_580,In_1251,In_1675);
nand U581 (N_581,In_270,In_1010);
nor U582 (N_582,In_1482,In_51);
or U583 (N_583,In_1530,In_969);
and U584 (N_584,In_171,In_821);
nor U585 (N_585,In_2125,In_27);
or U586 (N_586,In_1221,In_2496);
nand U587 (N_587,In_1421,In_1428);
and U588 (N_588,In_594,In_1282);
and U589 (N_589,In_1127,In_2151);
or U590 (N_590,In_699,In_2067);
and U591 (N_591,In_1597,In_379);
nor U592 (N_592,In_324,In_790);
nand U593 (N_593,In_590,In_1588);
and U594 (N_594,In_2178,In_1170);
or U595 (N_595,In_788,In_2259);
or U596 (N_596,In_2400,In_2291);
or U597 (N_597,In_25,In_137);
or U598 (N_598,In_2349,In_1112);
nor U599 (N_599,In_2358,In_1933);
nor U600 (N_600,In_2412,In_1536);
and U601 (N_601,In_727,In_118);
nor U602 (N_602,In_2099,In_499);
nor U603 (N_603,In_425,In_648);
nor U604 (N_604,In_1580,In_406);
or U605 (N_605,In_1195,In_1388);
and U606 (N_606,In_732,In_228);
nor U607 (N_607,In_319,In_1962);
nor U608 (N_608,In_2035,In_1302);
nor U609 (N_609,In_2431,In_285);
nand U610 (N_610,In_1008,In_469);
nand U611 (N_611,In_2467,In_172);
nand U612 (N_612,In_1440,In_1427);
and U613 (N_613,In_192,In_2281);
and U614 (N_614,In_1878,In_528);
nor U615 (N_615,In_2215,In_1198);
nand U616 (N_616,In_1691,In_2034);
or U617 (N_617,In_2244,In_1201);
nand U618 (N_618,In_420,In_1419);
and U619 (N_619,In_1174,In_1777);
nand U620 (N_620,In_735,In_988);
and U621 (N_621,In_970,In_556);
nand U622 (N_622,In_1931,In_430);
nand U623 (N_623,In_1017,In_1132);
and U624 (N_624,In_463,In_317);
nor U625 (N_625,In_1068,In_1038);
nor U626 (N_626,In_1698,In_527);
or U627 (N_627,In_1993,In_1224);
and U628 (N_628,In_1454,In_963);
nor U629 (N_629,In_876,In_1095);
nand U630 (N_630,In_67,In_1358);
nand U631 (N_631,In_817,In_2374);
or U632 (N_632,In_1124,In_2045);
and U633 (N_633,In_38,In_1683);
and U634 (N_634,In_2008,In_441);
and U635 (N_635,In_1363,In_2403);
or U636 (N_636,In_1688,In_1025);
nor U637 (N_637,In_860,In_1150);
or U638 (N_638,In_1622,In_957);
nor U639 (N_639,In_1836,In_1585);
nand U640 (N_640,In_1120,In_169);
or U641 (N_641,In_391,In_1959);
nor U642 (N_642,In_1155,In_1434);
or U643 (N_643,In_2069,In_357);
and U644 (N_644,In_2037,In_212);
or U645 (N_645,In_93,In_2064);
or U646 (N_646,In_1800,In_1754);
and U647 (N_647,In_1370,In_1078);
nor U648 (N_648,In_799,In_2211);
nor U649 (N_649,In_1134,In_1913);
and U650 (N_650,In_922,In_931);
nor U651 (N_651,In_841,In_2082);
or U652 (N_652,In_809,In_579);
nor U653 (N_653,In_2423,In_1737);
and U654 (N_654,In_959,In_65);
or U655 (N_655,In_88,In_1485);
and U656 (N_656,In_1097,In_1254);
nand U657 (N_657,In_1813,In_2366);
nor U658 (N_658,In_607,In_686);
nor U659 (N_659,In_2306,In_135);
and U660 (N_660,In_1021,In_1722);
and U661 (N_661,In_2321,In_1230);
nor U662 (N_662,In_2441,In_1080);
nand U663 (N_663,In_1206,In_1725);
and U664 (N_664,In_2261,In_1490);
and U665 (N_665,In_2319,In_92);
nor U666 (N_666,In_1462,In_1776);
or U667 (N_667,In_1847,In_558);
or U668 (N_668,In_681,In_1271);
nand U669 (N_669,In_1808,In_998);
nand U670 (N_670,In_1205,In_335);
or U671 (N_671,In_255,In_1692);
nand U672 (N_672,In_1601,In_2101);
xnor U673 (N_673,In_280,In_261);
nor U674 (N_674,In_1220,In_1840);
nor U675 (N_675,In_1649,In_761);
or U676 (N_676,In_1891,In_2459);
nor U677 (N_677,In_678,In_436);
nand U678 (N_678,In_701,In_2390);
nand U679 (N_679,In_1974,In_2304);
nor U680 (N_680,In_1548,In_410);
nor U681 (N_681,In_1184,In_1176);
or U682 (N_682,In_330,In_672);
xor U683 (N_683,In_1105,In_2074);
nor U684 (N_684,In_2269,In_264);
and U685 (N_685,In_1664,In_2005);
and U686 (N_686,In_974,In_356);
nand U687 (N_687,In_1089,In_2129);
and U688 (N_688,In_1906,In_229);
nand U689 (N_689,In_600,In_1934);
nand U690 (N_690,In_339,In_2236);
nand U691 (N_691,In_2139,In_1721);
nand U692 (N_692,In_1702,In_369);
nand U693 (N_693,In_1244,In_749);
nand U694 (N_694,In_2174,In_1415);
nor U695 (N_695,In_2144,In_1022);
nor U696 (N_696,In_2434,In_151);
nor U697 (N_697,In_2324,In_2262);
nand U698 (N_698,In_1192,In_932);
or U699 (N_699,In_1275,In_1992);
and U700 (N_700,In_1803,In_1502);
and U701 (N_701,In_1860,In_1509);
nor U702 (N_702,In_1378,In_629);
or U703 (N_703,In_203,In_1470);
and U704 (N_704,In_1861,In_2029);
nand U705 (N_705,In_2484,In_1322);
nor U706 (N_706,In_2410,In_1199);
nand U707 (N_707,In_2387,In_116);
nand U708 (N_708,In_1043,In_1243);
or U709 (N_709,In_1041,In_637);
and U710 (N_710,In_359,In_1241);
nor U711 (N_711,In_1075,In_709);
and U712 (N_712,In_2131,In_2232);
nand U713 (N_713,In_2238,In_1568);
and U714 (N_714,In_1455,In_1778);
nand U715 (N_715,In_1426,In_947);
nand U716 (N_716,In_2213,In_62);
nor U717 (N_717,In_1200,In_673);
or U718 (N_718,In_1149,In_497);
nand U719 (N_719,In_1289,In_864);
nor U720 (N_720,In_1178,In_7);
or U721 (N_721,In_286,In_1367);
nand U722 (N_722,In_688,In_2081);
nor U723 (N_723,In_1799,In_2368);
or U724 (N_724,In_1694,In_1050);
or U725 (N_725,In_2348,In_615);
and U726 (N_726,In_0,In_2090);
nor U727 (N_727,In_1612,In_777);
and U728 (N_728,In_2433,In_2033);
and U729 (N_729,In_782,In_1795);
or U730 (N_730,In_1966,In_1058);
and U731 (N_731,In_650,In_143);
and U732 (N_732,In_1939,In_1379);
nand U733 (N_733,In_2186,In_2474);
and U734 (N_734,In_1121,In_1708);
nor U735 (N_735,In_1886,In_245);
and U736 (N_736,In_2019,In_2065);
nor U737 (N_737,In_1920,In_321);
nand U738 (N_738,In_90,In_1212);
nor U739 (N_739,In_1273,In_492);
nor U740 (N_740,In_366,In_220);
and U741 (N_741,In_1500,In_1818);
nor U742 (N_742,In_500,In_1387);
nor U743 (N_743,In_543,In_2342);
and U744 (N_744,In_2369,In_1892);
or U745 (N_745,In_2224,In_1837);
nor U746 (N_746,In_1845,In_353);
and U747 (N_747,In_2429,In_1286);
nor U748 (N_748,In_2015,In_75);
or U749 (N_749,In_1774,In_2254);
nor U750 (N_750,In_1361,In_1420);
nor U751 (N_751,In_309,In_1012);
and U752 (N_752,In_1788,In_2258);
nor U753 (N_753,In_1266,In_867);
or U754 (N_754,In_1750,In_1887);
nor U755 (N_755,In_250,In_1562);
nor U756 (N_756,In_768,In_2197);
and U757 (N_757,In_934,In_756);
xor U758 (N_758,In_918,In_1209);
nor U759 (N_759,In_2367,In_17);
nand U760 (N_760,In_1002,In_1154);
nor U761 (N_761,In_2280,In_1644);
nand U762 (N_762,In_1492,In_1344);
or U763 (N_763,In_1971,In_2267);
nor U764 (N_764,In_1325,In_1261);
or U765 (N_765,In_111,In_1941);
and U766 (N_766,In_1392,In_769);
nor U767 (N_767,In_1459,In_612);
and U768 (N_768,In_852,In_2168);
or U769 (N_769,In_1377,In_375);
or U770 (N_770,In_837,In_750);
nand U771 (N_771,In_1339,In_1128);
nor U772 (N_772,In_413,In_1073);
nand U773 (N_773,In_1888,In_1908);
or U774 (N_774,In_1301,In_14);
nor U775 (N_775,In_541,In_2123);
nor U776 (N_776,In_862,In_318);
or U777 (N_777,In_2279,In_2492);
and U778 (N_778,In_181,In_997);
or U779 (N_779,In_2320,In_2191);
or U780 (N_780,In_1791,In_2491);
nor U781 (N_781,In_1372,In_778);
and U782 (N_782,In_1520,In_470);
nor U783 (N_783,In_2265,In_834);
nor U784 (N_784,In_298,In_765);
nor U785 (N_785,In_1893,In_2346);
nand U786 (N_786,In_872,In_1997);
nand U787 (N_787,In_930,In_625);
nor U788 (N_788,In_1287,In_2214);
nand U789 (N_789,In_1186,In_2009);
xor U790 (N_790,In_102,In_16);
nand U791 (N_791,In_284,In_411);
or U792 (N_792,In_2249,In_1403);
nor U793 (N_793,In_2001,In_900);
nand U794 (N_794,In_2231,In_438);
or U795 (N_795,In_2499,In_1090);
nand U796 (N_796,In_1175,In_1578);
nand U797 (N_797,In_2397,In_744);
nand U798 (N_798,In_2128,In_1605);
or U799 (N_799,In_178,In_1505);
and U800 (N_800,In_1396,In_708);
nor U801 (N_801,In_2072,In_1819);
xnor U802 (N_802,In_1281,In_2239);
or U803 (N_803,In_716,In_2470);
nor U804 (N_804,In_475,In_1009);
nand U805 (N_805,In_2089,In_658);
or U806 (N_806,In_1912,In_1065);
and U807 (N_807,In_2025,In_718);
nand U808 (N_808,In_18,In_2328);
nor U809 (N_809,In_159,In_498);
and U810 (N_810,In_1031,In_1782);
and U811 (N_811,In_2079,In_2250);
or U812 (N_812,In_566,In_2307);
nor U813 (N_813,In_943,In_674);
or U814 (N_814,In_1853,In_1533);
nor U815 (N_815,In_687,In_1554);
and U816 (N_816,In_293,In_1328);
nand U817 (N_817,In_440,In_1384);
or U818 (N_818,In_679,In_505);
and U819 (N_819,In_685,In_1755);
or U820 (N_820,In_1587,In_1457);
nand U821 (N_821,In_1323,In_1352);
or U822 (N_822,In_1765,In_1923);
nor U823 (N_823,In_1189,In_975);
and U824 (N_824,In_1216,In_1168);
or U825 (N_825,In_1488,In_447);
nand U826 (N_826,In_623,In_695);
and U827 (N_827,In_743,In_561);
nor U828 (N_828,In_935,In_2444);
and U829 (N_829,In_195,In_2179);
xor U830 (N_830,In_1259,In_207);
and U831 (N_831,In_1673,In_2458);
nand U832 (N_832,In_378,In_354);
nand U833 (N_833,In_129,In_507);
nand U834 (N_834,In_1850,In_941);
xor U835 (N_835,In_1496,In_1510);
and U836 (N_836,In_1719,In_465);
xor U837 (N_837,In_577,In_2223);
nand U838 (N_838,In_494,In_1924);
nor U839 (N_839,In_1756,In_206);
or U840 (N_840,In_1718,In_1429);
or U841 (N_841,In_1499,In_1166);
or U842 (N_842,In_1324,In_244);
nor U843 (N_843,In_2344,In_399);
or U844 (N_844,In_1233,In_435);
and U845 (N_845,In_689,In_176);
nand U846 (N_846,In_753,In_1137);
nor U847 (N_847,In_1775,In_2322);
nand U848 (N_848,In_91,In_2138);
nand U849 (N_849,In_2182,In_949);
and U850 (N_850,In_115,In_2203);
nand U851 (N_851,In_1249,In_1336);
nand U852 (N_852,In_893,In_1051);
and U853 (N_853,In_548,In_1207);
and U854 (N_854,In_820,In_555);
nand U855 (N_855,In_977,In_1817);
nand U856 (N_856,In_776,In_94);
nor U857 (N_857,In_723,In_1560);
or U858 (N_858,In_2222,In_481);
and U859 (N_859,In_1489,In_1780);
or U860 (N_860,In_1815,In_728);
nor U861 (N_861,In_1185,In_10);
nor U862 (N_862,In_1972,In_898);
xor U863 (N_863,In_891,In_856);
xnor U864 (N_864,In_1996,In_582);
nor U865 (N_865,In_1453,In_2422);
nor U866 (N_866,In_2468,In_344);
nand U867 (N_867,In_2420,In_1468);
nor U868 (N_868,In_48,In_1258);
nand U869 (N_869,In_243,In_763);
and U870 (N_870,In_866,In_1140);
nand U871 (N_871,In_1480,In_1871);
or U872 (N_872,In_112,In_2245);
nor U873 (N_873,In_644,In_1545);
nand U874 (N_874,In_2252,In_1169);
or U875 (N_875,In_2336,In_801);
or U876 (N_876,In_725,In_2012);
nand U877 (N_877,In_2169,In_1731);
nor U878 (N_878,In_1723,In_428);
nand U879 (N_879,In_37,In_2394);
or U880 (N_880,In_883,In_1758);
nand U881 (N_881,In_1831,In_400);
or U882 (N_882,In_976,In_6);
nand U883 (N_883,In_1048,In_752);
and U884 (N_884,In_1991,In_641);
nand U885 (N_885,In_1469,In_2195);
and U886 (N_886,In_1746,In_2003);
and U887 (N_887,In_296,In_868);
or U888 (N_888,In_248,In_896);
nor U889 (N_889,In_847,In_569);
nand U890 (N_890,In_706,In_302);
or U891 (N_891,In_1093,In_1862);
nand U892 (N_892,In_2380,In_2426);
nor U893 (N_893,In_2329,In_488);
and U894 (N_894,In_1634,In_2199);
nor U895 (N_895,In_1914,In_2447);
or U896 (N_896,In_216,In_1311);
and U897 (N_897,In_147,In_1211);
or U898 (N_898,In_2000,In_340);
and U899 (N_899,In_1472,In_1072);
or U900 (N_900,In_714,In_1160);
nand U901 (N_901,In_1823,In_144);
or U902 (N_902,In_2041,In_427);
nor U903 (N_903,In_2270,In_1019);
or U904 (N_904,In_2068,In_71);
or U905 (N_905,In_2086,In_443);
nor U906 (N_906,In_546,In_1821);
nor U907 (N_907,In_2218,In_1117);
nor U908 (N_908,In_1092,In_565);
nor U909 (N_909,In_2192,In_1464);
and U910 (N_910,In_204,In_895);
and U911 (N_911,In_1171,In_1408);
nor U912 (N_912,In_1820,In_1414);
nor U913 (N_913,In_2442,In_2161);
or U914 (N_914,In_31,In_72);
nor U915 (N_915,In_1433,In_279);
and U916 (N_916,In_372,In_850);
and U917 (N_917,In_325,In_2494);
nand U918 (N_918,In_1159,In_865);
nand U919 (N_919,In_184,In_1635);
or U920 (N_920,In_1643,In_609);
and U921 (N_921,In_1052,In_871);
or U922 (N_922,In_938,In_1096);
nor U923 (N_923,In_1521,In_417);
nand U924 (N_924,In_273,In_955);
nor U925 (N_925,In_642,In_2379);
nand U926 (N_926,In_1081,In_1600);
nor U927 (N_927,In_628,In_1555);
nor U928 (N_928,In_1786,In_2337);
nand U929 (N_929,In_2256,In_879);
nand U930 (N_930,In_1086,In_571);
nand U931 (N_931,In_1210,In_53);
or U932 (N_932,In_2187,In_1956);
nor U933 (N_933,In_1953,In_2021);
nor U934 (N_934,In_1125,In_2080);
nand U935 (N_935,In_2477,In_1114);
nor U936 (N_936,In_1687,In_1467);
nand U937 (N_937,In_2248,In_2106);
nand U938 (N_938,In_2112,In_442);
and U939 (N_939,In_57,In_553);
nor U940 (N_940,In_1214,In_2055);
and U941 (N_941,In_346,In_2316);
and U942 (N_942,In_300,In_770);
nor U943 (N_943,In_395,In_2370);
and U944 (N_944,In_167,In_1270);
nor U945 (N_945,In_622,In_41);
nor U946 (N_946,In_2126,In_620);
and U947 (N_947,In_1508,In_1331);
nand U948 (N_948,In_1347,In_1501);
nand U949 (N_949,In_2372,In_2048);
and U950 (N_950,In_2345,In_2120);
and U951 (N_951,In_2314,In_950);
and U952 (N_952,In_636,In_386);
xor U953 (N_953,In_1276,In_645);
nor U954 (N_954,In_1663,In_1549);
or U955 (N_955,In_301,In_1512);
nor U956 (N_956,In_1613,In_1373);
and U957 (N_957,In_45,In_1899);
nor U958 (N_958,In_1188,In_80);
nor U959 (N_959,In_1438,In_1828);
nor U960 (N_960,In_2352,In_290);
nor U961 (N_961,In_1881,In_2188);
nor U962 (N_962,In_2220,In_2283);
or U963 (N_963,In_1119,In_816);
or U964 (N_964,In_987,In_766);
or U965 (N_965,In_154,In_1925);
nor U966 (N_966,In_371,In_2437);
nand U967 (N_967,In_754,In_740);
nand U968 (N_968,In_1027,In_602);
or U969 (N_969,In_2130,In_786);
nor U970 (N_970,In_908,In_845);
nand U971 (N_971,In_836,In_278);
and U972 (N_972,In_713,In_1394);
or U973 (N_973,In_912,In_1595);
or U974 (N_974,In_2357,In_651);
nor U975 (N_975,In_2246,In_2255);
or U976 (N_976,In_1561,In_95);
nand U977 (N_977,In_355,In_1926);
or U978 (N_978,In_501,In_2498);
or U979 (N_979,In_731,In_247);
nand U980 (N_980,In_179,In_2335);
and U981 (N_981,In_1965,In_828);
nor U982 (N_982,In_2088,In_982);
or U983 (N_983,In_452,In_2170);
and U984 (N_984,In_163,In_199);
nand U985 (N_985,In_1676,In_1842);
and U986 (N_986,In_780,In_1016);
nand U987 (N_987,In_1173,In_345);
or U988 (N_988,In_985,In_1374);
and U989 (N_989,In_365,In_158);
nor U990 (N_990,In_168,In_721);
nand U991 (N_991,In_215,In_394);
and U992 (N_992,In_1695,In_390);
nor U993 (N_993,In_583,In_999);
nand U994 (N_994,In_1461,In_44);
or U995 (N_995,In_2073,In_1656);
or U996 (N_996,In_1064,In_1116);
or U997 (N_997,In_202,In_416);
nor U998 (N_998,In_2061,In_1870);
nand U999 (N_999,In_808,In_1390);
nor U1000 (N_1000,In_2078,In_604);
nor U1001 (N_1001,In_1528,In_308);
and U1002 (N_1002,In_1157,In_49);
or U1003 (N_1003,In_1621,In_1761);
nor U1004 (N_1004,In_2194,In_1632);
and U1005 (N_1005,In_403,In_2373);
and U1006 (N_1006,In_906,In_257);
nor U1007 (N_1007,In_1532,In_1527);
nor U1008 (N_1008,In_2052,In_1525);
and U1009 (N_1009,In_2226,In_2365);
or U1010 (N_1010,In_145,In_2340);
nand U1011 (N_1011,In_1341,In_1902);
nor U1012 (N_1012,In_1223,In_1658);
nand U1013 (N_1013,In_822,In_964);
or U1014 (N_1014,In_1798,In_1300);
nand U1015 (N_1015,In_455,In_1954);
or U1016 (N_1016,In_2027,In_1020);
and U1017 (N_1017,In_2208,In_506);
and U1018 (N_1018,In_933,In_1771);
nand U1019 (N_1019,In_738,In_1152);
nand U1020 (N_1020,In_653,In_1057);
nand U1021 (N_1021,In_907,In_698);
nand U1022 (N_1022,In_771,In_1785);
nand U1023 (N_1023,In_104,In_863);
or U1024 (N_1024,In_1227,In_155);
and U1025 (N_1025,In_396,In_2303);
nand U1026 (N_1026,In_2353,In_2201);
nor U1027 (N_1027,In_2385,In_2094);
xor U1028 (N_1028,In_2350,In_303);
or U1029 (N_1029,In_156,In_572);
nor U1030 (N_1030,In_283,In_311);
nor U1031 (N_1031,In_669,In_1400);
and U1032 (N_1032,In_2042,In_2212);
nand U1033 (N_1033,In_2175,In_1460);
and U1034 (N_1034,In_1631,In_1577);
nor U1035 (N_1035,In_1866,In_1740);
nor U1036 (N_1036,In_2323,In_1436);
and U1037 (N_1037,In_1099,In_2184);
nor U1038 (N_1038,In_2282,In_139);
nor U1039 (N_1039,In_2164,In_23);
or U1040 (N_1040,In_2293,In_47);
nor U1041 (N_1041,In_2095,In_1407);
or U1042 (N_1042,In_2219,In_1784);
nand U1043 (N_1043,In_705,In_530);
and U1044 (N_1044,In_1144,In_1629);
and U1045 (N_1045,In_2141,In_22);
and U1046 (N_1046,In_322,In_291);
and U1047 (N_1047,In_1158,In_739);
and U1048 (N_1048,In_1733,In_2202);
or U1049 (N_1049,In_710,In_812);
and U1050 (N_1050,In_2461,In_1088);
and U1051 (N_1051,In_358,In_2243);
or U1052 (N_1052,In_1320,In_1804);
nand U1053 (N_1053,In_1110,In_986);
or U1054 (N_1054,In_2341,In_1424);
and U1055 (N_1055,In_141,In_953);
or U1056 (N_1056,In_781,In_1350);
nand U1057 (N_1057,In_517,In_133);
nor U1058 (N_1058,In_40,In_2377);
and U1059 (N_1059,In_1061,In_2300);
or U1060 (N_1060,In_237,In_42);
nand U1061 (N_1061,In_24,In_382);
nor U1062 (N_1062,In_1856,In_794);
nor U1063 (N_1063,In_1654,In_2486);
nand U1064 (N_1064,In_1884,In_1165);
nor U1065 (N_1065,In_1668,In_1376);
nor U1066 (N_1066,In_2004,In_1182);
or U1067 (N_1067,In_1551,In_1094);
nor U1068 (N_1068,In_1639,In_875);
and U1069 (N_1069,In_886,In_946);
and U1070 (N_1070,In_810,In_1526);
and U1071 (N_1071,In_437,In_478);
nand U1072 (N_1072,In_2480,In_1987);
or U1073 (N_1073,In_2469,In_211);
nor U1074 (N_1074,In_2242,In_805);
or U1075 (N_1075,In_573,In_1402);
nand U1076 (N_1076,In_545,In_2100);
or U1077 (N_1077,In_1624,In_1743);
or U1078 (N_1078,In_1917,In_1814);
nor U1079 (N_1079,In_2338,In_1142);
nor U1080 (N_1080,In_2266,In_2196);
nand U1081 (N_1081,In_149,In_789);
or U1082 (N_1082,In_1108,In_874);
and U1083 (N_1083,In_1310,In_1768);
and U1084 (N_1084,In_1401,In_899);
nand U1085 (N_1085,In_654,In_1705);
or U1086 (N_1086,In_1425,In_1135);
nand U1087 (N_1087,In_1479,In_2295);
nor U1088 (N_1088,In_1868,In_1599);
or U1089 (N_1089,In_627,In_2378);
or U1090 (N_1090,In_1366,In_2058);
nand U1091 (N_1091,In_2424,In_1028);
and U1092 (N_1092,In_2206,In_1471);
nor U1093 (N_1093,In_483,In_591);
nor U1094 (N_1094,In_482,In_351);
and U1095 (N_1095,In_599,In_848);
or U1096 (N_1096,In_564,In_1309);
nor U1097 (N_1097,In_1995,In_1484);
and U1098 (N_1098,In_2327,In_2381);
nor U1099 (N_1099,In_804,In_2028);
nand U1100 (N_1100,In_664,In_811);
nand U1101 (N_1101,In_1263,In_331);
nor U1102 (N_1102,In_1734,In_1586);
or U1103 (N_1103,In_1062,In_1844);
nand U1104 (N_1104,In_2093,In_1565);
nand U1105 (N_1105,In_2167,In_468);
nand U1106 (N_1106,In_829,In_85);
nand U1107 (N_1107,In_1381,In_1717);
or U1108 (N_1108,In_2411,In_696);
nand U1109 (N_1109,In_1340,In_795);
nand U1110 (N_1110,In_1589,In_1735);
nand U1111 (N_1111,In_1849,In_1822);
or U1112 (N_1112,In_78,In_1442);
and U1113 (N_1113,In_60,In_927);
and U1114 (N_1114,In_1369,In_2060);
or U1115 (N_1115,In_1711,In_2294);
nand U1116 (N_1116,In_74,In_547);
or U1117 (N_1117,In_833,In_282);
and U1118 (N_1118,In_1059,In_1593);
nor U1119 (N_1119,In_1082,In_1594);
and U1120 (N_1120,In_724,In_103);
nor U1121 (N_1121,In_712,In_2117);
nor U1122 (N_1122,In_1976,In_1360);
nor U1123 (N_1123,In_1679,In_1355);
nor U1124 (N_1124,In_1641,In_1197);
and U1125 (N_1125,In_2062,In_194);
or U1126 (N_1126,In_775,In_888);
or U1127 (N_1127,In_377,In_218);
nand U1128 (N_1128,In_1279,In_1598);
and U1129 (N_1129,In_1337,In_68);
or U1130 (N_1130,In_2413,In_2156);
nor U1131 (N_1131,In_2024,In_1936);
or U1132 (N_1132,In_1486,In_1177);
and U1133 (N_1133,In_236,In_230);
and U1134 (N_1134,In_691,In_1553);
and U1135 (N_1135,In_1126,In_484);
nor U1136 (N_1136,In_2153,In_2039);
or U1137 (N_1137,In_2415,In_1304);
nor U1138 (N_1138,In_343,In_1332);
or U1139 (N_1139,In_968,In_2096);
and U1140 (N_1140,In_1122,In_1651);
and U1141 (N_1141,In_1910,In_1087);
nand U1142 (N_1142,In_292,In_614);
nand U1143 (N_1143,In_2493,In_2475);
nand U1144 (N_1144,In_2054,In_697);
nor U1145 (N_1145,In_1903,In_557);
and U1146 (N_1146,In_1955,In_361);
or U1147 (N_1147,In_2108,In_588);
xnor U1148 (N_1148,In_2450,In_29);
nor U1149 (N_1149,In_2122,In_1506);
nor U1150 (N_1150,In_1898,In_334);
and U1151 (N_1151,In_537,In_746);
nand U1152 (N_1152,In_1682,In_2193);
or U1153 (N_1153,In_626,In_2066);
or U1154 (N_1154,In_2489,In_110);
and U1155 (N_1155,In_1036,In_1707);
and U1156 (N_1156,In_1298,In_2333);
and U1157 (N_1157,In_380,In_919);
and U1158 (N_1158,In_2115,In_1802);
nand U1159 (N_1159,In_1163,In_213);
or U1160 (N_1160,In_551,In_8);
or U1161 (N_1161,In_64,In_1952);
nor U1162 (N_1162,In_1139,In_1498);
nor U1163 (N_1163,In_734,In_1343);
nand U1164 (N_1164,In_1943,In_1049);
or U1165 (N_1165,In_1760,In_2409);
and U1166 (N_1166,In_1037,In_707);
nand U1167 (N_1167,In_50,In_1677);
nand U1168 (N_1168,In_1053,In_2456);
or U1169 (N_1169,In_785,In_659);
or U1170 (N_1170,In_593,In_2023);
and U1171 (N_1171,In_838,In_2401);
and U1172 (N_1172,In_1628,In_1684);
nand U1173 (N_1173,In_646,In_682);
nand U1174 (N_1174,In_813,In_209);
or U1175 (N_1175,In_815,In_989);
or U1176 (N_1176,In_269,In_2145);
nor U1177 (N_1177,In_1416,In_2407);
nand U1178 (N_1178,In_1531,In_1085);
and U1179 (N_1179,In_503,In_1752);
or U1180 (N_1180,In_2275,In_2121);
nand U1181 (N_1181,In_2233,In_489);
and U1182 (N_1182,In_362,In_392);
or U1183 (N_1183,In_1660,In_1405);
nor U1184 (N_1184,In_1368,In_684);
nand U1185 (N_1185,In_1242,In_1246);
nand U1186 (N_1186,In_1614,In_1779);
and U1187 (N_1187,In_1909,In_189);
nor U1188 (N_1188,In_1167,In_2070);
and U1189 (N_1189,In_661,In_2406);
or U1190 (N_1190,In_2330,In_1652);
or U1191 (N_1191,In_1202,In_2296);
or U1192 (N_1192,In_222,In_1563);
nor U1193 (N_1193,In_2430,In_33);
nand U1194 (N_1194,In_108,In_1942);
nor U1195 (N_1195,In_694,In_1314);
nand U1196 (N_1196,In_542,In_774);
nand U1197 (N_1197,In_1478,In_1699);
nor U1198 (N_1198,In_2113,In_1252);
and U1199 (N_1199,In_1444,In_1491);
or U1200 (N_1200,In_1950,In_1446);
nor U1201 (N_1201,In_1147,In_2140);
nor U1202 (N_1202,In_587,In_2393);
and U1203 (N_1203,In_1029,In_1046);
nand U1204 (N_1204,In_46,In_2166);
nand U1205 (N_1205,In_767,In_327);
nor U1206 (N_1206,In_945,In_978);
and U1207 (N_1207,In_467,In_439);
nor U1208 (N_1208,In_861,In_2448);
and U1209 (N_1209,In_2419,In_954);
or U1210 (N_1210,In_2171,In_567);
or U1211 (N_1211,In_983,In_1904);
nand U1212 (N_1212,In_1885,In_79);
or U1213 (N_1213,In_316,In_512);
and U1214 (N_1214,In_460,In_418);
nor U1215 (N_1215,In_186,In_1507);
or U1216 (N_1216,In_1747,In_2310);
nor U1217 (N_1217,In_165,In_1326);
nor U1218 (N_1218,In_106,In_913);
nor U1219 (N_1219,In_1751,In_2026);
and U1220 (N_1220,In_1060,In_101);
nand U1221 (N_1221,In_1905,In_1265);
and U1222 (N_1222,In_965,In_649);
or U1223 (N_1223,In_1359,In_958);
nand U1224 (N_1224,In_393,In_849);
and U1225 (N_1225,In_1911,In_1417);
and U1226 (N_1226,In_267,In_1409);
nor U1227 (N_1227,In_136,In_1204);
nand U1228 (N_1228,In_1187,In_1412);
or U1229 (N_1229,In_1356,In_1984);
or U1230 (N_1230,In_2332,In_2439);
and U1231 (N_1231,In_2315,In_26);
nand U1232 (N_1232,In_1877,In_2017);
nand U1233 (N_1233,In_234,In_1115);
or U1234 (N_1234,In_519,In_897);
or U1235 (N_1235,In_827,In_2111);
and U1236 (N_1236,In_1353,In_2392);
nor U1237 (N_1237,In_1463,In_549);
nand U1238 (N_1238,In_166,In_2287);
and U1239 (N_1239,In_1789,In_1348);
and U1240 (N_1240,In_262,In_4);
nor U1241 (N_1241,In_1766,In_1667);
and U1242 (N_1242,In_1543,In_1449);
or U1243 (N_1243,In_823,In_693);
and U1244 (N_1244,In_1947,In_633);
and U1245 (N_1245,In_1889,In_966);
and U1246 (N_1246,In_1662,In_275);
nand U1247 (N_1247,In_1338,In_491);
and U1248 (N_1248,In_1738,In_1410);
nand U1249 (N_1249,In_210,In_531);
and U1250 (N_1250,In_1900,In_2117);
nand U1251 (N_1251,In_870,In_1391);
nor U1252 (N_1252,In_425,In_2389);
nand U1253 (N_1253,In_724,In_38);
nor U1254 (N_1254,In_1218,In_1235);
or U1255 (N_1255,In_1306,In_366);
nor U1256 (N_1256,In_884,In_2055);
nor U1257 (N_1257,In_102,In_1091);
and U1258 (N_1258,In_2021,In_133);
or U1259 (N_1259,In_1361,In_1852);
nor U1260 (N_1260,In_1130,In_2347);
nand U1261 (N_1261,In_2336,In_562);
nand U1262 (N_1262,In_1050,In_304);
and U1263 (N_1263,In_1033,In_1150);
nor U1264 (N_1264,In_100,In_369);
or U1265 (N_1265,In_1861,In_2017);
or U1266 (N_1266,In_743,In_2140);
and U1267 (N_1267,In_1849,In_448);
or U1268 (N_1268,In_1206,In_691);
nand U1269 (N_1269,In_278,In_1663);
and U1270 (N_1270,In_1068,In_1222);
or U1271 (N_1271,In_197,In_1021);
and U1272 (N_1272,In_1112,In_832);
or U1273 (N_1273,In_972,In_2130);
nor U1274 (N_1274,In_1627,In_1411);
nand U1275 (N_1275,In_73,In_900);
or U1276 (N_1276,In_2399,In_528);
or U1277 (N_1277,In_1180,In_2122);
xnor U1278 (N_1278,In_1615,In_777);
and U1279 (N_1279,In_1580,In_14);
nor U1280 (N_1280,In_1867,In_1396);
nand U1281 (N_1281,In_1784,In_1028);
and U1282 (N_1282,In_194,In_2067);
or U1283 (N_1283,In_1684,In_609);
nand U1284 (N_1284,In_2139,In_1391);
nand U1285 (N_1285,In_1972,In_1051);
or U1286 (N_1286,In_890,In_1651);
or U1287 (N_1287,In_2098,In_2024);
or U1288 (N_1288,In_1018,In_421);
nand U1289 (N_1289,In_862,In_2327);
nor U1290 (N_1290,In_226,In_1758);
nand U1291 (N_1291,In_997,In_2116);
nand U1292 (N_1292,In_338,In_222);
nor U1293 (N_1293,In_405,In_1730);
nand U1294 (N_1294,In_1411,In_438);
and U1295 (N_1295,In_462,In_1577);
nor U1296 (N_1296,In_1965,In_1944);
nor U1297 (N_1297,In_703,In_1936);
nand U1298 (N_1298,In_387,In_1950);
or U1299 (N_1299,In_1113,In_460);
or U1300 (N_1300,In_1471,In_190);
nor U1301 (N_1301,In_364,In_1673);
and U1302 (N_1302,In_694,In_488);
or U1303 (N_1303,In_1795,In_1571);
nand U1304 (N_1304,In_2473,In_887);
nand U1305 (N_1305,In_2019,In_2460);
nor U1306 (N_1306,In_941,In_2149);
nor U1307 (N_1307,In_2307,In_1696);
nor U1308 (N_1308,In_2162,In_2026);
or U1309 (N_1309,In_1331,In_1715);
nand U1310 (N_1310,In_193,In_218);
or U1311 (N_1311,In_464,In_1829);
xor U1312 (N_1312,In_1412,In_176);
nor U1313 (N_1313,In_1900,In_260);
or U1314 (N_1314,In_2458,In_2219);
and U1315 (N_1315,In_2148,In_1264);
or U1316 (N_1316,In_2235,In_2206);
nor U1317 (N_1317,In_14,In_136);
or U1318 (N_1318,In_2214,In_2200);
or U1319 (N_1319,In_228,In_644);
or U1320 (N_1320,In_2190,In_1983);
or U1321 (N_1321,In_1887,In_1986);
nand U1322 (N_1322,In_2454,In_1393);
or U1323 (N_1323,In_553,In_2046);
or U1324 (N_1324,In_117,In_889);
nand U1325 (N_1325,In_1593,In_303);
and U1326 (N_1326,In_1077,In_2368);
and U1327 (N_1327,In_990,In_1566);
nand U1328 (N_1328,In_2184,In_567);
nor U1329 (N_1329,In_172,In_737);
nand U1330 (N_1330,In_76,In_198);
and U1331 (N_1331,In_2177,In_1593);
nand U1332 (N_1332,In_181,In_2023);
and U1333 (N_1333,In_111,In_1251);
nor U1334 (N_1334,In_859,In_1229);
and U1335 (N_1335,In_2282,In_375);
nand U1336 (N_1336,In_795,In_1379);
nor U1337 (N_1337,In_1099,In_928);
and U1338 (N_1338,In_798,In_770);
and U1339 (N_1339,In_1511,In_2463);
nor U1340 (N_1340,In_1980,In_1717);
or U1341 (N_1341,In_1921,In_1982);
nand U1342 (N_1342,In_943,In_561);
nand U1343 (N_1343,In_2164,In_313);
and U1344 (N_1344,In_1207,In_190);
nor U1345 (N_1345,In_2176,In_257);
nor U1346 (N_1346,In_1821,In_472);
or U1347 (N_1347,In_2129,In_624);
or U1348 (N_1348,In_2358,In_2090);
and U1349 (N_1349,In_975,In_836);
nand U1350 (N_1350,In_45,In_331);
or U1351 (N_1351,In_541,In_257);
and U1352 (N_1352,In_801,In_1816);
and U1353 (N_1353,In_2263,In_2476);
nand U1354 (N_1354,In_763,In_449);
nor U1355 (N_1355,In_905,In_1185);
or U1356 (N_1356,In_592,In_1663);
or U1357 (N_1357,In_1288,In_1080);
nor U1358 (N_1358,In_2150,In_255);
nand U1359 (N_1359,In_308,In_2072);
nand U1360 (N_1360,In_235,In_412);
and U1361 (N_1361,In_1391,In_1193);
or U1362 (N_1362,In_799,In_2425);
and U1363 (N_1363,In_2492,In_514);
nand U1364 (N_1364,In_944,In_1911);
nand U1365 (N_1365,In_2398,In_1074);
and U1366 (N_1366,In_677,In_1500);
or U1367 (N_1367,In_192,In_232);
or U1368 (N_1368,In_317,In_645);
and U1369 (N_1369,In_1810,In_1762);
or U1370 (N_1370,In_2423,In_1424);
nand U1371 (N_1371,In_401,In_2151);
nand U1372 (N_1372,In_638,In_2458);
nand U1373 (N_1373,In_298,In_2300);
nand U1374 (N_1374,In_1371,In_1607);
or U1375 (N_1375,In_1881,In_1231);
or U1376 (N_1376,In_1305,In_2127);
nor U1377 (N_1377,In_1474,In_569);
and U1378 (N_1378,In_2045,In_745);
or U1379 (N_1379,In_963,In_2150);
or U1380 (N_1380,In_552,In_145);
and U1381 (N_1381,In_1809,In_1841);
and U1382 (N_1382,In_1198,In_136);
nor U1383 (N_1383,In_188,In_612);
or U1384 (N_1384,In_1984,In_1104);
and U1385 (N_1385,In_465,In_1016);
nand U1386 (N_1386,In_99,In_1024);
and U1387 (N_1387,In_704,In_392);
nand U1388 (N_1388,In_1963,In_624);
nand U1389 (N_1389,In_916,In_669);
and U1390 (N_1390,In_2259,In_1431);
nand U1391 (N_1391,In_1598,In_1593);
and U1392 (N_1392,In_1309,In_878);
or U1393 (N_1393,In_1105,In_1973);
nor U1394 (N_1394,In_59,In_2311);
nand U1395 (N_1395,In_1839,In_942);
and U1396 (N_1396,In_1706,In_2365);
nand U1397 (N_1397,In_528,In_612);
or U1398 (N_1398,In_1526,In_1715);
nor U1399 (N_1399,In_697,In_120);
and U1400 (N_1400,In_2439,In_1463);
nor U1401 (N_1401,In_764,In_1067);
and U1402 (N_1402,In_1104,In_529);
or U1403 (N_1403,In_248,In_1058);
and U1404 (N_1404,In_2189,In_1655);
or U1405 (N_1405,In_1883,In_1637);
and U1406 (N_1406,In_1920,In_642);
nand U1407 (N_1407,In_880,In_1178);
and U1408 (N_1408,In_527,In_2348);
nor U1409 (N_1409,In_1958,In_1185);
and U1410 (N_1410,In_1215,In_1249);
or U1411 (N_1411,In_1177,In_1965);
and U1412 (N_1412,In_589,In_412);
nor U1413 (N_1413,In_934,In_2442);
nor U1414 (N_1414,In_2424,In_591);
or U1415 (N_1415,In_2089,In_779);
nor U1416 (N_1416,In_1476,In_860);
or U1417 (N_1417,In_1283,In_619);
nand U1418 (N_1418,In_767,In_1499);
xnor U1419 (N_1419,In_1905,In_757);
nor U1420 (N_1420,In_2258,In_1169);
nor U1421 (N_1421,In_1273,In_2205);
nor U1422 (N_1422,In_227,In_2454);
nand U1423 (N_1423,In_1936,In_2243);
nor U1424 (N_1424,In_2095,In_493);
or U1425 (N_1425,In_2391,In_2192);
and U1426 (N_1426,In_1303,In_1178);
nand U1427 (N_1427,In_1800,In_1159);
nand U1428 (N_1428,In_2370,In_2156);
or U1429 (N_1429,In_1196,In_2138);
and U1430 (N_1430,In_1890,In_1963);
nand U1431 (N_1431,In_1118,In_691);
nand U1432 (N_1432,In_355,In_319);
and U1433 (N_1433,In_1784,In_383);
nor U1434 (N_1434,In_2235,In_1246);
nand U1435 (N_1435,In_1478,In_2491);
and U1436 (N_1436,In_1348,In_1016);
and U1437 (N_1437,In_2263,In_1235);
or U1438 (N_1438,In_638,In_884);
nand U1439 (N_1439,In_1580,In_914);
and U1440 (N_1440,In_751,In_711);
nor U1441 (N_1441,In_2368,In_60);
or U1442 (N_1442,In_100,In_1705);
or U1443 (N_1443,In_2105,In_1052);
nor U1444 (N_1444,In_15,In_1854);
and U1445 (N_1445,In_2200,In_1001);
nor U1446 (N_1446,In_1028,In_715);
nor U1447 (N_1447,In_1009,In_1288);
and U1448 (N_1448,In_904,In_1227);
nor U1449 (N_1449,In_2172,In_1397);
nor U1450 (N_1450,In_425,In_558);
nand U1451 (N_1451,In_1711,In_77);
and U1452 (N_1452,In_40,In_492);
or U1453 (N_1453,In_1451,In_2149);
nand U1454 (N_1454,In_1734,In_1892);
and U1455 (N_1455,In_1151,In_2407);
nor U1456 (N_1456,In_1563,In_2329);
nor U1457 (N_1457,In_101,In_2424);
and U1458 (N_1458,In_481,In_1767);
nor U1459 (N_1459,In_253,In_1634);
or U1460 (N_1460,In_2404,In_936);
nand U1461 (N_1461,In_1829,In_2176);
nor U1462 (N_1462,In_2128,In_1777);
or U1463 (N_1463,In_1280,In_1816);
nand U1464 (N_1464,In_2385,In_1231);
nor U1465 (N_1465,In_1283,In_2025);
nand U1466 (N_1466,In_622,In_651);
nor U1467 (N_1467,In_2132,In_165);
nor U1468 (N_1468,In_979,In_95);
or U1469 (N_1469,In_757,In_1877);
nand U1470 (N_1470,In_1012,In_1238);
or U1471 (N_1471,In_166,In_1345);
and U1472 (N_1472,In_955,In_566);
and U1473 (N_1473,In_445,In_1307);
nand U1474 (N_1474,In_195,In_1492);
nor U1475 (N_1475,In_268,In_1146);
and U1476 (N_1476,In_1928,In_2059);
and U1477 (N_1477,In_2214,In_1569);
nor U1478 (N_1478,In_691,In_214);
nor U1479 (N_1479,In_2083,In_642);
xnor U1480 (N_1480,In_62,In_550);
nand U1481 (N_1481,In_940,In_1197);
or U1482 (N_1482,In_758,In_1020);
nor U1483 (N_1483,In_632,In_168);
nor U1484 (N_1484,In_747,In_1516);
and U1485 (N_1485,In_1803,In_2069);
and U1486 (N_1486,In_1281,In_1968);
and U1487 (N_1487,In_175,In_2334);
nor U1488 (N_1488,In_1637,In_1407);
or U1489 (N_1489,In_1846,In_2129);
or U1490 (N_1490,In_1660,In_1341);
or U1491 (N_1491,In_1819,In_680);
nor U1492 (N_1492,In_1976,In_1315);
and U1493 (N_1493,In_33,In_234);
and U1494 (N_1494,In_228,In_1501);
or U1495 (N_1495,In_1863,In_1390);
nand U1496 (N_1496,In_1041,In_1824);
nand U1497 (N_1497,In_2339,In_837);
nor U1498 (N_1498,In_1168,In_1669);
or U1499 (N_1499,In_1793,In_1924);
nand U1500 (N_1500,In_21,In_1262);
nor U1501 (N_1501,In_2137,In_2444);
or U1502 (N_1502,In_793,In_1070);
nand U1503 (N_1503,In_323,In_1224);
or U1504 (N_1504,In_1584,In_1725);
nor U1505 (N_1505,In_529,In_1342);
nor U1506 (N_1506,In_648,In_1611);
and U1507 (N_1507,In_1222,In_2000);
nand U1508 (N_1508,In_2386,In_2378);
xnor U1509 (N_1509,In_1754,In_1219);
nand U1510 (N_1510,In_265,In_1720);
nand U1511 (N_1511,In_989,In_1744);
nor U1512 (N_1512,In_139,In_665);
and U1513 (N_1513,In_3,In_2196);
and U1514 (N_1514,In_1660,In_258);
or U1515 (N_1515,In_1770,In_344);
and U1516 (N_1516,In_785,In_1029);
and U1517 (N_1517,In_2074,In_2338);
and U1518 (N_1518,In_209,In_1635);
and U1519 (N_1519,In_2031,In_2018);
nor U1520 (N_1520,In_433,In_1908);
nor U1521 (N_1521,In_51,In_2148);
nand U1522 (N_1522,In_870,In_97);
or U1523 (N_1523,In_2495,In_2445);
nand U1524 (N_1524,In_1577,In_818);
nor U1525 (N_1525,In_1389,In_1152);
nor U1526 (N_1526,In_1637,In_23);
or U1527 (N_1527,In_1997,In_767);
nor U1528 (N_1528,In_911,In_551);
and U1529 (N_1529,In_163,In_307);
and U1530 (N_1530,In_1661,In_794);
nand U1531 (N_1531,In_1511,In_2136);
nor U1532 (N_1532,In_1495,In_780);
nor U1533 (N_1533,In_1434,In_395);
nor U1534 (N_1534,In_1266,In_1794);
nand U1535 (N_1535,In_195,In_1637);
nand U1536 (N_1536,In_1248,In_938);
nor U1537 (N_1537,In_1365,In_896);
or U1538 (N_1538,In_314,In_1479);
and U1539 (N_1539,In_300,In_2225);
or U1540 (N_1540,In_822,In_1472);
nand U1541 (N_1541,In_1327,In_999);
nor U1542 (N_1542,In_1314,In_2194);
nand U1543 (N_1543,In_2278,In_108);
nand U1544 (N_1544,In_2382,In_2090);
nand U1545 (N_1545,In_679,In_1453);
and U1546 (N_1546,In_1750,In_333);
and U1547 (N_1547,In_619,In_2414);
or U1548 (N_1548,In_1948,In_1081);
xor U1549 (N_1549,In_942,In_755);
and U1550 (N_1550,In_2341,In_241);
and U1551 (N_1551,In_1477,In_776);
or U1552 (N_1552,In_92,In_354);
nand U1553 (N_1553,In_1481,In_1916);
and U1554 (N_1554,In_113,In_315);
and U1555 (N_1555,In_1532,In_1663);
nor U1556 (N_1556,In_135,In_1802);
or U1557 (N_1557,In_821,In_40);
or U1558 (N_1558,In_566,In_1844);
nand U1559 (N_1559,In_1335,In_1931);
and U1560 (N_1560,In_617,In_1669);
nand U1561 (N_1561,In_2309,In_1163);
and U1562 (N_1562,In_1587,In_968);
nor U1563 (N_1563,In_986,In_1334);
nor U1564 (N_1564,In_1547,In_2295);
nor U1565 (N_1565,In_456,In_2485);
nor U1566 (N_1566,In_1999,In_2057);
nor U1567 (N_1567,In_2352,In_1298);
nor U1568 (N_1568,In_1970,In_446);
nor U1569 (N_1569,In_423,In_1092);
nand U1570 (N_1570,In_2395,In_1360);
and U1571 (N_1571,In_1503,In_192);
nor U1572 (N_1572,In_1207,In_1752);
nand U1573 (N_1573,In_1621,In_761);
or U1574 (N_1574,In_754,In_509);
or U1575 (N_1575,In_1837,In_2097);
nor U1576 (N_1576,In_895,In_656);
nor U1577 (N_1577,In_468,In_1692);
or U1578 (N_1578,In_2243,In_352);
or U1579 (N_1579,In_1741,In_2464);
nand U1580 (N_1580,In_1274,In_1701);
nor U1581 (N_1581,In_628,In_1434);
and U1582 (N_1582,In_1314,In_347);
or U1583 (N_1583,In_2259,In_1731);
or U1584 (N_1584,In_1104,In_169);
and U1585 (N_1585,In_1979,In_2168);
nor U1586 (N_1586,In_116,In_1984);
or U1587 (N_1587,In_2058,In_1553);
nor U1588 (N_1588,In_239,In_824);
nor U1589 (N_1589,In_1520,In_2357);
and U1590 (N_1590,In_1822,In_1218);
nor U1591 (N_1591,In_1524,In_1698);
nand U1592 (N_1592,In_2211,In_1752);
nand U1593 (N_1593,In_544,In_537);
and U1594 (N_1594,In_279,In_1982);
or U1595 (N_1595,In_915,In_1054);
nand U1596 (N_1596,In_2253,In_408);
nor U1597 (N_1597,In_2218,In_2477);
and U1598 (N_1598,In_2387,In_1760);
or U1599 (N_1599,In_1486,In_331);
and U1600 (N_1600,In_873,In_1686);
nor U1601 (N_1601,In_1885,In_1144);
nand U1602 (N_1602,In_463,In_2494);
or U1603 (N_1603,In_2012,In_248);
nand U1604 (N_1604,In_1097,In_147);
or U1605 (N_1605,In_60,In_1993);
or U1606 (N_1606,In_889,In_493);
nor U1607 (N_1607,In_1788,In_1220);
nand U1608 (N_1608,In_1742,In_71);
and U1609 (N_1609,In_1587,In_2208);
nand U1610 (N_1610,In_1415,In_948);
nand U1611 (N_1611,In_765,In_714);
nand U1612 (N_1612,In_1429,In_198);
nor U1613 (N_1613,In_1352,In_2442);
nor U1614 (N_1614,In_628,In_1742);
nand U1615 (N_1615,In_1973,In_2184);
nor U1616 (N_1616,In_2458,In_2008);
nand U1617 (N_1617,In_1201,In_721);
nand U1618 (N_1618,In_361,In_118);
nor U1619 (N_1619,In_2263,In_1801);
nor U1620 (N_1620,In_1857,In_2386);
nand U1621 (N_1621,In_1960,In_588);
nor U1622 (N_1622,In_1895,In_1084);
nor U1623 (N_1623,In_926,In_595);
or U1624 (N_1624,In_2142,In_2263);
or U1625 (N_1625,In_2438,In_2465);
and U1626 (N_1626,In_2377,In_2164);
nor U1627 (N_1627,In_2030,In_1958);
nor U1628 (N_1628,In_245,In_2105);
or U1629 (N_1629,In_1593,In_2346);
or U1630 (N_1630,In_1864,In_368);
and U1631 (N_1631,In_2054,In_175);
nor U1632 (N_1632,In_2240,In_744);
and U1633 (N_1633,In_849,In_719);
and U1634 (N_1634,In_2273,In_2340);
nor U1635 (N_1635,In_1,In_1216);
nor U1636 (N_1636,In_1503,In_1942);
nor U1637 (N_1637,In_1861,In_467);
nand U1638 (N_1638,In_812,In_2368);
and U1639 (N_1639,In_2348,In_346);
nor U1640 (N_1640,In_1267,In_1374);
or U1641 (N_1641,In_238,In_1949);
or U1642 (N_1642,In_42,In_2324);
nand U1643 (N_1643,In_2207,In_993);
nand U1644 (N_1644,In_2015,In_322);
nand U1645 (N_1645,In_1724,In_2150);
xor U1646 (N_1646,In_1836,In_2036);
and U1647 (N_1647,In_561,In_993);
nor U1648 (N_1648,In_1216,In_2247);
nor U1649 (N_1649,In_710,In_1980);
nand U1650 (N_1650,In_1888,In_161);
nand U1651 (N_1651,In_453,In_147);
or U1652 (N_1652,In_2281,In_271);
nand U1653 (N_1653,In_2393,In_118);
and U1654 (N_1654,In_310,In_1738);
nand U1655 (N_1655,In_2412,In_514);
nor U1656 (N_1656,In_1222,In_396);
nor U1657 (N_1657,In_2436,In_914);
nor U1658 (N_1658,In_880,In_1333);
or U1659 (N_1659,In_2433,In_2395);
nand U1660 (N_1660,In_658,In_1580);
and U1661 (N_1661,In_255,In_2227);
or U1662 (N_1662,In_2494,In_60);
and U1663 (N_1663,In_1836,In_1407);
nor U1664 (N_1664,In_637,In_668);
nor U1665 (N_1665,In_520,In_2296);
and U1666 (N_1666,In_1882,In_2045);
or U1667 (N_1667,In_91,In_2064);
nand U1668 (N_1668,In_1659,In_924);
nand U1669 (N_1669,In_2270,In_617);
or U1670 (N_1670,In_246,In_597);
nand U1671 (N_1671,In_580,In_512);
and U1672 (N_1672,In_1845,In_1931);
and U1673 (N_1673,In_133,In_339);
nor U1674 (N_1674,In_1294,In_480);
and U1675 (N_1675,In_1335,In_1081);
and U1676 (N_1676,In_1061,In_1176);
nand U1677 (N_1677,In_1960,In_2237);
nand U1678 (N_1678,In_1687,In_175);
nor U1679 (N_1679,In_1057,In_1099);
and U1680 (N_1680,In_1714,In_86);
or U1681 (N_1681,In_244,In_196);
or U1682 (N_1682,In_1792,In_372);
nor U1683 (N_1683,In_1365,In_1931);
or U1684 (N_1684,In_460,In_1402);
or U1685 (N_1685,In_29,In_1047);
and U1686 (N_1686,In_2446,In_719);
or U1687 (N_1687,In_2172,In_1545);
or U1688 (N_1688,In_80,In_833);
and U1689 (N_1689,In_2408,In_2149);
and U1690 (N_1690,In_371,In_23);
and U1691 (N_1691,In_427,In_1253);
nor U1692 (N_1692,In_793,In_1847);
nand U1693 (N_1693,In_189,In_272);
or U1694 (N_1694,In_1645,In_1131);
nand U1695 (N_1695,In_2200,In_1272);
nand U1696 (N_1696,In_1404,In_927);
nor U1697 (N_1697,In_2375,In_322);
nor U1698 (N_1698,In_1277,In_245);
and U1699 (N_1699,In_559,In_738);
xor U1700 (N_1700,In_1631,In_1599);
xnor U1701 (N_1701,In_727,In_2351);
and U1702 (N_1702,In_352,In_4);
and U1703 (N_1703,In_1202,In_791);
and U1704 (N_1704,In_1547,In_2005);
or U1705 (N_1705,In_844,In_1791);
nand U1706 (N_1706,In_1747,In_608);
nand U1707 (N_1707,In_1998,In_199);
or U1708 (N_1708,In_261,In_1099);
nor U1709 (N_1709,In_2491,In_1328);
or U1710 (N_1710,In_2217,In_55);
and U1711 (N_1711,In_858,In_576);
and U1712 (N_1712,In_1054,In_1175);
or U1713 (N_1713,In_1966,In_1760);
and U1714 (N_1714,In_1803,In_1337);
nand U1715 (N_1715,In_157,In_976);
and U1716 (N_1716,In_1040,In_2251);
and U1717 (N_1717,In_488,In_996);
or U1718 (N_1718,In_243,In_1936);
and U1719 (N_1719,In_979,In_1681);
and U1720 (N_1720,In_1410,In_2295);
nand U1721 (N_1721,In_1875,In_997);
nand U1722 (N_1722,In_171,In_2290);
or U1723 (N_1723,In_1187,In_2408);
nand U1724 (N_1724,In_1833,In_1321);
nand U1725 (N_1725,In_312,In_1270);
and U1726 (N_1726,In_1032,In_565);
or U1727 (N_1727,In_1587,In_1961);
and U1728 (N_1728,In_1716,In_2205);
and U1729 (N_1729,In_886,In_2315);
nor U1730 (N_1730,In_1818,In_1565);
or U1731 (N_1731,In_1460,In_1567);
or U1732 (N_1732,In_498,In_1675);
or U1733 (N_1733,In_2273,In_1312);
nand U1734 (N_1734,In_1409,In_201);
nor U1735 (N_1735,In_637,In_2132);
nor U1736 (N_1736,In_70,In_2191);
and U1737 (N_1737,In_2107,In_995);
nand U1738 (N_1738,In_2342,In_983);
nor U1739 (N_1739,In_1396,In_607);
or U1740 (N_1740,In_824,In_2269);
and U1741 (N_1741,In_2277,In_779);
nand U1742 (N_1742,In_1637,In_1009);
or U1743 (N_1743,In_1299,In_591);
nand U1744 (N_1744,In_140,In_777);
and U1745 (N_1745,In_1026,In_1987);
nand U1746 (N_1746,In_1338,In_2479);
or U1747 (N_1747,In_1846,In_1033);
nand U1748 (N_1748,In_1850,In_1982);
nor U1749 (N_1749,In_327,In_381);
nor U1750 (N_1750,In_1474,In_323);
or U1751 (N_1751,In_1307,In_2411);
and U1752 (N_1752,In_32,In_526);
nor U1753 (N_1753,In_1994,In_2132);
and U1754 (N_1754,In_883,In_1594);
nor U1755 (N_1755,In_794,In_463);
nand U1756 (N_1756,In_2129,In_157);
nor U1757 (N_1757,In_1778,In_507);
or U1758 (N_1758,In_1976,In_981);
and U1759 (N_1759,In_1324,In_1450);
nand U1760 (N_1760,In_1825,In_883);
nand U1761 (N_1761,In_551,In_1986);
and U1762 (N_1762,In_1229,In_1971);
or U1763 (N_1763,In_304,In_236);
and U1764 (N_1764,In_16,In_1563);
and U1765 (N_1765,In_2195,In_1296);
nand U1766 (N_1766,In_211,In_1965);
and U1767 (N_1767,In_1924,In_881);
nor U1768 (N_1768,In_2314,In_775);
nor U1769 (N_1769,In_426,In_37);
or U1770 (N_1770,In_1386,In_1694);
nand U1771 (N_1771,In_459,In_1345);
and U1772 (N_1772,In_2347,In_23);
nand U1773 (N_1773,In_2344,In_1768);
or U1774 (N_1774,In_796,In_2244);
or U1775 (N_1775,In_1121,In_749);
nor U1776 (N_1776,In_1361,In_1516);
or U1777 (N_1777,In_489,In_2002);
or U1778 (N_1778,In_160,In_709);
and U1779 (N_1779,In_739,In_1201);
and U1780 (N_1780,In_891,In_1863);
and U1781 (N_1781,In_2289,In_2224);
or U1782 (N_1782,In_2419,In_2087);
or U1783 (N_1783,In_1170,In_1890);
nand U1784 (N_1784,In_2194,In_448);
and U1785 (N_1785,In_729,In_1658);
nand U1786 (N_1786,In_1951,In_1549);
nand U1787 (N_1787,In_1222,In_2413);
nand U1788 (N_1788,In_1025,In_2004);
nor U1789 (N_1789,In_2061,In_1668);
or U1790 (N_1790,In_663,In_283);
nand U1791 (N_1791,In_1342,In_2387);
nor U1792 (N_1792,In_82,In_1397);
nand U1793 (N_1793,In_431,In_1824);
and U1794 (N_1794,In_1979,In_1071);
nand U1795 (N_1795,In_539,In_1682);
or U1796 (N_1796,In_1045,In_1010);
or U1797 (N_1797,In_1721,In_1292);
and U1798 (N_1798,In_2081,In_2262);
nand U1799 (N_1799,In_1120,In_819);
and U1800 (N_1800,In_2452,In_1869);
or U1801 (N_1801,In_1178,In_1026);
nor U1802 (N_1802,In_310,In_1915);
and U1803 (N_1803,In_226,In_1493);
or U1804 (N_1804,In_1879,In_306);
and U1805 (N_1805,In_723,In_559);
or U1806 (N_1806,In_902,In_2044);
or U1807 (N_1807,In_2333,In_2089);
nand U1808 (N_1808,In_2167,In_1151);
nor U1809 (N_1809,In_1304,In_2470);
nand U1810 (N_1810,In_1525,In_55);
xor U1811 (N_1811,In_696,In_114);
nor U1812 (N_1812,In_23,In_2482);
or U1813 (N_1813,In_1014,In_1642);
nand U1814 (N_1814,In_2133,In_1875);
or U1815 (N_1815,In_647,In_2209);
or U1816 (N_1816,In_1894,In_1995);
and U1817 (N_1817,In_1981,In_2419);
or U1818 (N_1818,In_1697,In_1675);
nand U1819 (N_1819,In_1136,In_388);
nand U1820 (N_1820,In_1626,In_2193);
nor U1821 (N_1821,In_689,In_649);
nor U1822 (N_1822,In_550,In_2496);
and U1823 (N_1823,In_786,In_1083);
or U1824 (N_1824,In_1082,In_26);
and U1825 (N_1825,In_2455,In_1134);
and U1826 (N_1826,In_806,In_1766);
nand U1827 (N_1827,In_1590,In_867);
and U1828 (N_1828,In_135,In_1275);
or U1829 (N_1829,In_2073,In_599);
nor U1830 (N_1830,In_838,In_1588);
nor U1831 (N_1831,In_1244,In_1172);
nor U1832 (N_1832,In_2188,In_956);
or U1833 (N_1833,In_1877,In_333);
nand U1834 (N_1834,In_538,In_2395);
or U1835 (N_1835,In_344,In_1917);
nand U1836 (N_1836,In_917,In_906);
nand U1837 (N_1837,In_603,In_788);
and U1838 (N_1838,In_1665,In_1234);
or U1839 (N_1839,In_1215,In_1617);
nand U1840 (N_1840,In_741,In_702);
and U1841 (N_1841,In_1974,In_2192);
and U1842 (N_1842,In_929,In_1494);
nor U1843 (N_1843,In_1232,In_1883);
nor U1844 (N_1844,In_189,In_597);
nor U1845 (N_1845,In_2457,In_273);
nor U1846 (N_1846,In_142,In_669);
nor U1847 (N_1847,In_274,In_881);
nand U1848 (N_1848,In_571,In_128);
or U1849 (N_1849,In_2067,In_365);
and U1850 (N_1850,In_944,In_454);
and U1851 (N_1851,In_675,In_2173);
or U1852 (N_1852,In_383,In_1249);
and U1853 (N_1853,In_45,In_1506);
and U1854 (N_1854,In_727,In_888);
nor U1855 (N_1855,In_1024,In_1984);
or U1856 (N_1856,In_855,In_506);
and U1857 (N_1857,In_1272,In_821);
or U1858 (N_1858,In_1895,In_810);
nor U1859 (N_1859,In_2327,In_1075);
nor U1860 (N_1860,In_2011,In_266);
nand U1861 (N_1861,In_1333,In_2474);
nor U1862 (N_1862,In_1058,In_562);
and U1863 (N_1863,In_699,In_765);
nand U1864 (N_1864,In_54,In_1654);
or U1865 (N_1865,In_67,In_1318);
and U1866 (N_1866,In_2282,In_330);
nor U1867 (N_1867,In_629,In_1032);
nand U1868 (N_1868,In_800,In_393);
nor U1869 (N_1869,In_2353,In_1960);
nand U1870 (N_1870,In_261,In_157);
and U1871 (N_1871,In_1781,In_2095);
nand U1872 (N_1872,In_1401,In_1737);
or U1873 (N_1873,In_2196,In_2373);
or U1874 (N_1874,In_1198,In_564);
or U1875 (N_1875,In_51,In_2493);
and U1876 (N_1876,In_1194,In_1196);
nor U1877 (N_1877,In_2333,In_1128);
nand U1878 (N_1878,In_922,In_1744);
or U1879 (N_1879,In_375,In_451);
or U1880 (N_1880,In_689,In_1603);
and U1881 (N_1881,In_339,In_1385);
nand U1882 (N_1882,In_306,In_1843);
or U1883 (N_1883,In_2023,In_1668);
nand U1884 (N_1884,In_403,In_128);
nand U1885 (N_1885,In_528,In_2488);
or U1886 (N_1886,In_844,In_997);
or U1887 (N_1887,In_53,In_1655);
or U1888 (N_1888,In_1580,In_484);
or U1889 (N_1889,In_1427,In_558);
nor U1890 (N_1890,In_1173,In_180);
nand U1891 (N_1891,In_1585,In_1707);
nor U1892 (N_1892,In_1853,In_1326);
and U1893 (N_1893,In_2269,In_1608);
and U1894 (N_1894,In_1270,In_2435);
and U1895 (N_1895,In_1197,In_977);
or U1896 (N_1896,In_2482,In_1103);
and U1897 (N_1897,In_2312,In_1287);
or U1898 (N_1898,In_597,In_366);
or U1899 (N_1899,In_1973,In_1506);
or U1900 (N_1900,In_2347,In_2038);
nor U1901 (N_1901,In_665,In_2295);
and U1902 (N_1902,In_1721,In_1817);
nor U1903 (N_1903,In_605,In_75);
or U1904 (N_1904,In_17,In_505);
or U1905 (N_1905,In_1374,In_1786);
nand U1906 (N_1906,In_2324,In_1393);
or U1907 (N_1907,In_1294,In_409);
nor U1908 (N_1908,In_1699,In_290);
nand U1909 (N_1909,In_451,In_321);
nand U1910 (N_1910,In_1330,In_373);
nor U1911 (N_1911,In_570,In_1117);
nor U1912 (N_1912,In_599,In_1237);
nand U1913 (N_1913,In_2464,In_2019);
and U1914 (N_1914,In_1598,In_334);
nand U1915 (N_1915,In_232,In_634);
nand U1916 (N_1916,In_750,In_85);
nor U1917 (N_1917,In_686,In_1546);
nand U1918 (N_1918,In_1783,In_2259);
nand U1919 (N_1919,In_294,In_1550);
nor U1920 (N_1920,In_13,In_1925);
nor U1921 (N_1921,In_327,In_120);
or U1922 (N_1922,In_505,In_638);
or U1923 (N_1923,In_2400,In_1947);
or U1924 (N_1924,In_2311,In_2101);
nor U1925 (N_1925,In_1982,In_1284);
nor U1926 (N_1926,In_1588,In_73);
nand U1927 (N_1927,In_522,In_512);
and U1928 (N_1928,In_658,In_2273);
and U1929 (N_1929,In_2202,In_223);
or U1930 (N_1930,In_376,In_804);
or U1931 (N_1931,In_1120,In_862);
and U1932 (N_1932,In_2259,In_1730);
or U1933 (N_1933,In_2328,In_761);
and U1934 (N_1934,In_1422,In_2186);
and U1935 (N_1935,In_2344,In_1439);
or U1936 (N_1936,In_2285,In_2289);
or U1937 (N_1937,In_438,In_671);
nor U1938 (N_1938,In_199,In_2135);
and U1939 (N_1939,In_731,In_661);
or U1940 (N_1940,In_1819,In_768);
or U1941 (N_1941,In_1464,In_1685);
nor U1942 (N_1942,In_2180,In_660);
and U1943 (N_1943,In_1974,In_414);
nand U1944 (N_1944,In_1358,In_1736);
nand U1945 (N_1945,In_2114,In_538);
or U1946 (N_1946,In_1230,In_1712);
or U1947 (N_1947,In_1205,In_1170);
nor U1948 (N_1948,In_465,In_1115);
nor U1949 (N_1949,In_1007,In_110);
or U1950 (N_1950,In_116,In_1297);
nor U1951 (N_1951,In_983,In_1274);
or U1952 (N_1952,In_1939,In_1579);
nand U1953 (N_1953,In_804,In_855);
nand U1954 (N_1954,In_553,In_1197);
and U1955 (N_1955,In_595,In_1104);
nand U1956 (N_1956,In_274,In_1228);
and U1957 (N_1957,In_2036,In_2310);
nor U1958 (N_1958,In_574,In_1836);
nor U1959 (N_1959,In_81,In_263);
and U1960 (N_1960,In_1894,In_1433);
and U1961 (N_1961,In_1814,In_2233);
nand U1962 (N_1962,In_218,In_1295);
and U1963 (N_1963,In_2470,In_1986);
and U1964 (N_1964,In_1515,In_1884);
nor U1965 (N_1965,In_430,In_102);
or U1966 (N_1966,In_746,In_2409);
and U1967 (N_1967,In_1022,In_119);
nor U1968 (N_1968,In_493,In_2176);
and U1969 (N_1969,In_137,In_319);
xnor U1970 (N_1970,In_1110,In_1291);
and U1971 (N_1971,In_2380,In_2327);
or U1972 (N_1972,In_2187,In_1101);
and U1973 (N_1973,In_2122,In_76);
and U1974 (N_1974,In_2152,In_2138);
and U1975 (N_1975,In_1317,In_1959);
and U1976 (N_1976,In_2182,In_1412);
nor U1977 (N_1977,In_759,In_1821);
nor U1978 (N_1978,In_162,In_1079);
or U1979 (N_1979,In_67,In_776);
or U1980 (N_1980,In_2100,In_2271);
nor U1981 (N_1981,In_994,In_2296);
nor U1982 (N_1982,In_1207,In_1573);
and U1983 (N_1983,In_1317,In_2028);
or U1984 (N_1984,In_1821,In_1651);
nand U1985 (N_1985,In_415,In_179);
nor U1986 (N_1986,In_1768,In_1950);
or U1987 (N_1987,In_1086,In_2070);
or U1988 (N_1988,In_118,In_2425);
or U1989 (N_1989,In_1383,In_2168);
and U1990 (N_1990,In_2147,In_2055);
nor U1991 (N_1991,In_1993,In_490);
nor U1992 (N_1992,In_960,In_385);
or U1993 (N_1993,In_1067,In_907);
and U1994 (N_1994,In_1363,In_1912);
nand U1995 (N_1995,In_3,In_1118);
nand U1996 (N_1996,In_756,In_2312);
or U1997 (N_1997,In_1980,In_1000);
or U1998 (N_1998,In_1994,In_290);
and U1999 (N_1999,In_1431,In_2463);
or U2000 (N_2000,In_1073,In_307);
or U2001 (N_2001,In_1098,In_1776);
nand U2002 (N_2002,In_1643,In_1548);
nor U2003 (N_2003,In_713,In_383);
nand U2004 (N_2004,In_2339,In_1706);
or U2005 (N_2005,In_1412,In_1832);
or U2006 (N_2006,In_329,In_2259);
and U2007 (N_2007,In_279,In_2271);
nor U2008 (N_2008,In_1830,In_411);
xor U2009 (N_2009,In_2032,In_1384);
and U2010 (N_2010,In_245,In_471);
nor U2011 (N_2011,In_259,In_1867);
or U2012 (N_2012,In_1349,In_1541);
or U2013 (N_2013,In_1220,In_2477);
nand U2014 (N_2014,In_1335,In_2285);
and U2015 (N_2015,In_1381,In_366);
and U2016 (N_2016,In_1791,In_1424);
nor U2017 (N_2017,In_1021,In_1811);
nor U2018 (N_2018,In_1754,In_1875);
nor U2019 (N_2019,In_2293,In_1196);
and U2020 (N_2020,In_1872,In_246);
nor U2021 (N_2021,In_2069,In_22);
nor U2022 (N_2022,In_2020,In_1946);
or U2023 (N_2023,In_1536,In_831);
or U2024 (N_2024,In_1172,In_519);
and U2025 (N_2025,In_2432,In_991);
and U2026 (N_2026,In_180,In_2003);
nand U2027 (N_2027,In_2253,In_217);
xor U2028 (N_2028,In_1743,In_2331);
or U2029 (N_2029,In_2470,In_1565);
or U2030 (N_2030,In_524,In_1934);
nor U2031 (N_2031,In_1764,In_1394);
or U2032 (N_2032,In_1569,In_297);
nand U2033 (N_2033,In_1832,In_2354);
nand U2034 (N_2034,In_967,In_1458);
nor U2035 (N_2035,In_2451,In_196);
and U2036 (N_2036,In_2161,In_1086);
nor U2037 (N_2037,In_346,In_1160);
and U2038 (N_2038,In_2464,In_1031);
nand U2039 (N_2039,In_722,In_1774);
and U2040 (N_2040,In_1791,In_149);
nor U2041 (N_2041,In_1249,In_2182);
nand U2042 (N_2042,In_1027,In_1324);
nor U2043 (N_2043,In_2384,In_1190);
and U2044 (N_2044,In_1167,In_1986);
or U2045 (N_2045,In_1076,In_1386);
nor U2046 (N_2046,In_1604,In_1287);
or U2047 (N_2047,In_824,In_1486);
nor U2048 (N_2048,In_1736,In_1802);
and U2049 (N_2049,In_1379,In_309);
nand U2050 (N_2050,In_1682,In_1632);
and U2051 (N_2051,In_86,In_1867);
nand U2052 (N_2052,In_2077,In_2238);
xnor U2053 (N_2053,In_1279,In_1032);
nand U2054 (N_2054,In_1544,In_1607);
and U2055 (N_2055,In_1961,In_2265);
nand U2056 (N_2056,In_971,In_942);
and U2057 (N_2057,In_966,In_1147);
or U2058 (N_2058,In_2210,In_1027);
or U2059 (N_2059,In_2298,In_2421);
and U2060 (N_2060,In_1171,In_710);
xnor U2061 (N_2061,In_674,In_1840);
or U2062 (N_2062,In_1048,In_570);
or U2063 (N_2063,In_1958,In_711);
and U2064 (N_2064,In_1009,In_302);
nand U2065 (N_2065,In_1607,In_1688);
and U2066 (N_2066,In_2473,In_741);
nor U2067 (N_2067,In_367,In_1704);
nand U2068 (N_2068,In_1284,In_1577);
nand U2069 (N_2069,In_2369,In_69);
nand U2070 (N_2070,In_1447,In_717);
or U2071 (N_2071,In_708,In_2341);
and U2072 (N_2072,In_1727,In_1316);
and U2073 (N_2073,In_106,In_333);
or U2074 (N_2074,In_2325,In_2411);
and U2075 (N_2075,In_1728,In_1433);
and U2076 (N_2076,In_191,In_1006);
and U2077 (N_2077,In_850,In_1061);
nand U2078 (N_2078,In_1719,In_1483);
or U2079 (N_2079,In_2088,In_1719);
and U2080 (N_2080,In_1973,In_1178);
nor U2081 (N_2081,In_1309,In_2403);
nand U2082 (N_2082,In_1751,In_1582);
nor U2083 (N_2083,In_2029,In_553);
or U2084 (N_2084,In_1037,In_593);
nor U2085 (N_2085,In_450,In_1547);
nor U2086 (N_2086,In_1661,In_1221);
nor U2087 (N_2087,In_1398,In_2075);
and U2088 (N_2088,In_1960,In_1618);
nand U2089 (N_2089,In_1751,In_551);
and U2090 (N_2090,In_1016,In_1227);
nand U2091 (N_2091,In_1022,In_878);
and U2092 (N_2092,In_441,In_1528);
and U2093 (N_2093,In_997,In_2405);
or U2094 (N_2094,In_1630,In_2466);
nand U2095 (N_2095,In_455,In_1686);
nand U2096 (N_2096,In_2449,In_1820);
and U2097 (N_2097,In_1325,In_2390);
nor U2098 (N_2098,In_1925,In_155);
and U2099 (N_2099,In_157,In_557);
nand U2100 (N_2100,In_1255,In_2129);
nor U2101 (N_2101,In_677,In_2016);
nand U2102 (N_2102,In_1831,In_1530);
nand U2103 (N_2103,In_869,In_985);
xnor U2104 (N_2104,In_791,In_1911);
and U2105 (N_2105,In_356,In_1362);
nand U2106 (N_2106,In_1595,In_1021);
nor U2107 (N_2107,In_65,In_542);
and U2108 (N_2108,In_1796,In_1251);
nor U2109 (N_2109,In_2475,In_183);
and U2110 (N_2110,In_1176,In_226);
nand U2111 (N_2111,In_2142,In_1269);
nor U2112 (N_2112,In_939,In_1430);
nor U2113 (N_2113,In_1064,In_877);
and U2114 (N_2114,In_1687,In_191);
nand U2115 (N_2115,In_1741,In_1785);
nand U2116 (N_2116,In_1734,In_2492);
and U2117 (N_2117,In_127,In_2311);
or U2118 (N_2118,In_508,In_1421);
and U2119 (N_2119,In_2059,In_2418);
nor U2120 (N_2120,In_70,In_1584);
nand U2121 (N_2121,In_750,In_197);
or U2122 (N_2122,In_1638,In_1986);
or U2123 (N_2123,In_784,In_228);
and U2124 (N_2124,In_490,In_1659);
nand U2125 (N_2125,In_2272,In_1360);
and U2126 (N_2126,In_168,In_2444);
nor U2127 (N_2127,In_2328,In_948);
nor U2128 (N_2128,In_1017,In_330);
nor U2129 (N_2129,In_796,In_385);
nand U2130 (N_2130,In_1869,In_2088);
nand U2131 (N_2131,In_1478,In_1679);
nor U2132 (N_2132,In_1764,In_367);
nor U2133 (N_2133,In_1166,In_2275);
or U2134 (N_2134,In_1831,In_1016);
nor U2135 (N_2135,In_1852,In_2445);
or U2136 (N_2136,In_89,In_2194);
nor U2137 (N_2137,In_1120,In_1441);
nor U2138 (N_2138,In_529,In_2289);
and U2139 (N_2139,In_736,In_2419);
or U2140 (N_2140,In_1009,In_169);
nand U2141 (N_2141,In_707,In_1138);
nand U2142 (N_2142,In_2253,In_1451);
nor U2143 (N_2143,In_971,In_1859);
or U2144 (N_2144,In_2388,In_1225);
nor U2145 (N_2145,In_2261,In_1075);
nor U2146 (N_2146,In_2042,In_1487);
nor U2147 (N_2147,In_92,In_801);
nor U2148 (N_2148,In_1365,In_2278);
nor U2149 (N_2149,In_715,In_1508);
nand U2150 (N_2150,In_2413,In_1385);
and U2151 (N_2151,In_86,In_2473);
or U2152 (N_2152,In_1936,In_275);
nand U2153 (N_2153,In_488,In_617);
and U2154 (N_2154,In_2279,In_1967);
nand U2155 (N_2155,In_654,In_1627);
nor U2156 (N_2156,In_1489,In_1612);
nand U2157 (N_2157,In_2183,In_256);
and U2158 (N_2158,In_2047,In_208);
nor U2159 (N_2159,In_2242,In_292);
nor U2160 (N_2160,In_914,In_582);
and U2161 (N_2161,In_1914,In_1261);
and U2162 (N_2162,In_2342,In_1715);
and U2163 (N_2163,In_1012,In_1706);
nand U2164 (N_2164,In_861,In_876);
nand U2165 (N_2165,In_568,In_2200);
nor U2166 (N_2166,In_824,In_575);
nor U2167 (N_2167,In_487,In_1907);
nand U2168 (N_2168,In_1559,In_793);
nand U2169 (N_2169,In_1850,In_530);
nand U2170 (N_2170,In_2075,In_91);
nand U2171 (N_2171,In_481,In_227);
nand U2172 (N_2172,In_1939,In_913);
and U2173 (N_2173,In_1309,In_1745);
and U2174 (N_2174,In_1519,In_1958);
and U2175 (N_2175,In_976,In_1756);
nand U2176 (N_2176,In_1163,In_1677);
or U2177 (N_2177,In_2001,In_667);
and U2178 (N_2178,In_874,In_1091);
or U2179 (N_2179,In_1296,In_630);
or U2180 (N_2180,In_1806,In_311);
nor U2181 (N_2181,In_998,In_1079);
nand U2182 (N_2182,In_1648,In_1671);
or U2183 (N_2183,In_1450,In_214);
and U2184 (N_2184,In_1382,In_1776);
nor U2185 (N_2185,In_1423,In_2385);
and U2186 (N_2186,In_1202,In_2096);
or U2187 (N_2187,In_490,In_451);
and U2188 (N_2188,In_809,In_1512);
and U2189 (N_2189,In_2449,In_1054);
nand U2190 (N_2190,In_1093,In_961);
nor U2191 (N_2191,In_1275,In_395);
nor U2192 (N_2192,In_1262,In_840);
nor U2193 (N_2193,In_2081,In_1244);
nand U2194 (N_2194,In_449,In_1826);
and U2195 (N_2195,In_385,In_915);
and U2196 (N_2196,In_1659,In_2011);
nand U2197 (N_2197,In_1179,In_948);
nand U2198 (N_2198,In_1981,In_575);
nand U2199 (N_2199,In_18,In_2391);
nor U2200 (N_2200,In_945,In_1822);
and U2201 (N_2201,In_99,In_752);
nor U2202 (N_2202,In_1755,In_793);
nor U2203 (N_2203,In_2198,In_2180);
or U2204 (N_2204,In_1291,In_959);
nand U2205 (N_2205,In_2058,In_170);
nand U2206 (N_2206,In_1281,In_775);
or U2207 (N_2207,In_1395,In_2142);
nor U2208 (N_2208,In_1691,In_2412);
nand U2209 (N_2209,In_2459,In_2296);
nand U2210 (N_2210,In_1390,In_442);
nor U2211 (N_2211,In_1516,In_125);
nand U2212 (N_2212,In_1646,In_1480);
and U2213 (N_2213,In_2390,In_340);
nor U2214 (N_2214,In_596,In_1610);
or U2215 (N_2215,In_1376,In_268);
nor U2216 (N_2216,In_1529,In_1583);
or U2217 (N_2217,In_2340,In_157);
nand U2218 (N_2218,In_1802,In_482);
or U2219 (N_2219,In_2109,In_2307);
and U2220 (N_2220,In_418,In_835);
or U2221 (N_2221,In_456,In_119);
nor U2222 (N_2222,In_1126,In_1255);
nand U2223 (N_2223,In_1842,In_1089);
and U2224 (N_2224,In_1653,In_984);
nor U2225 (N_2225,In_1843,In_798);
nor U2226 (N_2226,In_1893,In_2092);
nand U2227 (N_2227,In_41,In_351);
nand U2228 (N_2228,In_2129,In_138);
or U2229 (N_2229,In_1325,In_562);
or U2230 (N_2230,In_212,In_337);
or U2231 (N_2231,In_2000,In_2232);
and U2232 (N_2232,In_988,In_24);
or U2233 (N_2233,In_723,In_1797);
or U2234 (N_2234,In_2067,In_753);
or U2235 (N_2235,In_504,In_1194);
nor U2236 (N_2236,In_1422,In_526);
and U2237 (N_2237,In_968,In_2099);
nor U2238 (N_2238,In_2162,In_815);
or U2239 (N_2239,In_2360,In_1449);
nand U2240 (N_2240,In_545,In_773);
and U2241 (N_2241,In_1429,In_952);
nor U2242 (N_2242,In_298,In_2226);
nor U2243 (N_2243,In_2330,In_2146);
or U2244 (N_2244,In_112,In_2160);
or U2245 (N_2245,In_1653,In_416);
nand U2246 (N_2246,In_2424,In_1349);
nand U2247 (N_2247,In_1125,In_2456);
or U2248 (N_2248,In_2313,In_604);
nor U2249 (N_2249,In_229,In_1482);
and U2250 (N_2250,In_988,In_22);
nand U2251 (N_2251,In_1535,In_457);
nor U2252 (N_2252,In_1407,In_327);
xor U2253 (N_2253,In_1127,In_2193);
or U2254 (N_2254,In_1454,In_710);
nor U2255 (N_2255,In_990,In_2249);
nor U2256 (N_2256,In_1455,In_1006);
xnor U2257 (N_2257,In_1776,In_1364);
or U2258 (N_2258,In_1539,In_371);
nand U2259 (N_2259,In_1694,In_1597);
nand U2260 (N_2260,In_1570,In_1179);
nand U2261 (N_2261,In_157,In_490);
or U2262 (N_2262,In_1054,In_1009);
or U2263 (N_2263,In_1726,In_2111);
nand U2264 (N_2264,In_1044,In_463);
nand U2265 (N_2265,In_1098,In_1952);
or U2266 (N_2266,In_899,In_642);
nand U2267 (N_2267,In_162,In_1235);
xor U2268 (N_2268,In_1210,In_1181);
and U2269 (N_2269,In_78,In_2201);
nor U2270 (N_2270,In_1372,In_1468);
nand U2271 (N_2271,In_1128,In_2422);
nand U2272 (N_2272,In_2447,In_1825);
nand U2273 (N_2273,In_746,In_318);
or U2274 (N_2274,In_989,In_2201);
nand U2275 (N_2275,In_912,In_1393);
nor U2276 (N_2276,In_2386,In_350);
nand U2277 (N_2277,In_1472,In_2306);
or U2278 (N_2278,In_1820,In_1762);
and U2279 (N_2279,In_1289,In_720);
or U2280 (N_2280,In_1919,In_1929);
or U2281 (N_2281,In_2468,In_2034);
nor U2282 (N_2282,In_1385,In_1703);
or U2283 (N_2283,In_1609,In_464);
or U2284 (N_2284,In_1517,In_1747);
or U2285 (N_2285,In_1627,In_2134);
and U2286 (N_2286,In_1283,In_1346);
nor U2287 (N_2287,In_1122,In_652);
nor U2288 (N_2288,In_242,In_40);
nor U2289 (N_2289,In_2469,In_930);
or U2290 (N_2290,In_756,In_1062);
nor U2291 (N_2291,In_1247,In_2489);
nand U2292 (N_2292,In_190,In_1244);
or U2293 (N_2293,In_2035,In_768);
or U2294 (N_2294,In_2252,In_1924);
xnor U2295 (N_2295,In_504,In_1694);
nor U2296 (N_2296,In_2333,In_1520);
nand U2297 (N_2297,In_2025,In_247);
or U2298 (N_2298,In_2490,In_1316);
xnor U2299 (N_2299,In_1728,In_1816);
nand U2300 (N_2300,In_2001,In_2084);
nor U2301 (N_2301,In_1386,In_182);
or U2302 (N_2302,In_264,In_1009);
or U2303 (N_2303,In_325,In_2215);
or U2304 (N_2304,In_2391,In_403);
and U2305 (N_2305,In_600,In_826);
nor U2306 (N_2306,In_2398,In_376);
nor U2307 (N_2307,In_177,In_634);
or U2308 (N_2308,In_505,In_2249);
nand U2309 (N_2309,In_23,In_1699);
or U2310 (N_2310,In_240,In_1213);
nand U2311 (N_2311,In_995,In_1430);
or U2312 (N_2312,In_705,In_1306);
or U2313 (N_2313,In_2189,In_2353);
nand U2314 (N_2314,In_1464,In_1569);
and U2315 (N_2315,In_1067,In_301);
nor U2316 (N_2316,In_920,In_2132);
and U2317 (N_2317,In_1579,In_1684);
nor U2318 (N_2318,In_1131,In_1993);
nor U2319 (N_2319,In_1769,In_40);
nand U2320 (N_2320,In_1801,In_1743);
and U2321 (N_2321,In_394,In_1982);
or U2322 (N_2322,In_1677,In_1561);
nor U2323 (N_2323,In_1334,In_1838);
or U2324 (N_2324,In_1489,In_1076);
and U2325 (N_2325,In_1032,In_1512);
and U2326 (N_2326,In_1201,In_2469);
and U2327 (N_2327,In_1972,In_1922);
or U2328 (N_2328,In_766,In_2022);
nor U2329 (N_2329,In_1039,In_16);
or U2330 (N_2330,In_1674,In_1319);
and U2331 (N_2331,In_1795,In_850);
or U2332 (N_2332,In_679,In_1395);
and U2333 (N_2333,In_2109,In_1677);
xnor U2334 (N_2334,In_852,In_828);
nand U2335 (N_2335,In_1591,In_339);
nand U2336 (N_2336,In_185,In_491);
or U2337 (N_2337,In_179,In_2023);
or U2338 (N_2338,In_1734,In_716);
nand U2339 (N_2339,In_870,In_1941);
nor U2340 (N_2340,In_869,In_1228);
nand U2341 (N_2341,In_1517,In_513);
or U2342 (N_2342,In_931,In_1926);
and U2343 (N_2343,In_354,In_1361);
or U2344 (N_2344,In_1128,In_2008);
or U2345 (N_2345,In_2307,In_680);
nor U2346 (N_2346,In_996,In_1361);
or U2347 (N_2347,In_230,In_33);
and U2348 (N_2348,In_2359,In_1175);
and U2349 (N_2349,In_1099,In_1543);
and U2350 (N_2350,In_2300,In_1410);
nand U2351 (N_2351,In_2377,In_2171);
nor U2352 (N_2352,In_1867,In_511);
nor U2353 (N_2353,In_533,In_666);
or U2354 (N_2354,In_248,In_1059);
nand U2355 (N_2355,In_957,In_1255);
nor U2356 (N_2356,In_381,In_1200);
nor U2357 (N_2357,In_767,In_415);
nand U2358 (N_2358,In_2396,In_645);
or U2359 (N_2359,In_1703,In_1981);
nand U2360 (N_2360,In_688,In_732);
nand U2361 (N_2361,In_96,In_241);
nor U2362 (N_2362,In_1369,In_1234);
or U2363 (N_2363,In_1172,In_457);
and U2364 (N_2364,In_25,In_1292);
or U2365 (N_2365,In_585,In_43);
nor U2366 (N_2366,In_11,In_2293);
nand U2367 (N_2367,In_1553,In_2265);
nand U2368 (N_2368,In_1161,In_971);
and U2369 (N_2369,In_2498,In_287);
and U2370 (N_2370,In_2029,In_1403);
nor U2371 (N_2371,In_2143,In_844);
nand U2372 (N_2372,In_512,In_1188);
nor U2373 (N_2373,In_1116,In_2039);
or U2374 (N_2374,In_1279,In_1938);
nor U2375 (N_2375,In_2418,In_1369);
and U2376 (N_2376,In_378,In_2442);
nand U2377 (N_2377,In_2249,In_507);
nand U2378 (N_2378,In_2336,In_1536);
or U2379 (N_2379,In_1218,In_1992);
nor U2380 (N_2380,In_2013,In_1194);
nor U2381 (N_2381,In_2490,In_1737);
or U2382 (N_2382,In_1881,In_175);
and U2383 (N_2383,In_379,In_1807);
and U2384 (N_2384,In_461,In_1846);
or U2385 (N_2385,In_681,In_1806);
and U2386 (N_2386,In_1103,In_1307);
nor U2387 (N_2387,In_1613,In_576);
nand U2388 (N_2388,In_702,In_1337);
xnor U2389 (N_2389,In_1158,In_1500);
nor U2390 (N_2390,In_2403,In_932);
or U2391 (N_2391,In_1776,In_102);
nor U2392 (N_2392,In_1513,In_1160);
or U2393 (N_2393,In_2226,In_1206);
or U2394 (N_2394,In_919,In_901);
or U2395 (N_2395,In_981,In_2345);
and U2396 (N_2396,In_1361,In_1645);
nand U2397 (N_2397,In_500,In_729);
nand U2398 (N_2398,In_2296,In_1961);
nand U2399 (N_2399,In_1910,In_1767);
nor U2400 (N_2400,In_2064,In_1408);
nand U2401 (N_2401,In_170,In_949);
nor U2402 (N_2402,In_2185,In_1589);
or U2403 (N_2403,In_819,In_347);
and U2404 (N_2404,In_581,In_2144);
and U2405 (N_2405,In_61,In_2269);
and U2406 (N_2406,In_2105,In_2382);
nand U2407 (N_2407,In_1848,In_2346);
or U2408 (N_2408,In_1644,In_1024);
nand U2409 (N_2409,In_529,In_1571);
or U2410 (N_2410,In_1956,In_1055);
and U2411 (N_2411,In_47,In_1091);
and U2412 (N_2412,In_206,In_2344);
nand U2413 (N_2413,In_1543,In_1855);
or U2414 (N_2414,In_1085,In_842);
nor U2415 (N_2415,In_1159,In_1576);
nor U2416 (N_2416,In_2107,In_1757);
and U2417 (N_2417,In_2085,In_176);
or U2418 (N_2418,In_1307,In_364);
or U2419 (N_2419,In_412,In_569);
nor U2420 (N_2420,In_947,In_310);
and U2421 (N_2421,In_470,In_306);
nand U2422 (N_2422,In_1768,In_2090);
nor U2423 (N_2423,In_1154,In_8);
or U2424 (N_2424,In_2330,In_946);
nand U2425 (N_2425,In_1267,In_2140);
nand U2426 (N_2426,In_24,In_1574);
and U2427 (N_2427,In_1081,In_2162);
nand U2428 (N_2428,In_2139,In_2203);
xnor U2429 (N_2429,In_834,In_1300);
nand U2430 (N_2430,In_2106,In_566);
or U2431 (N_2431,In_1848,In_2092);
nand U2432 (N_2432,In_669,In_29);
nor U2433 (N_2433,In_1768,In_2225);
nor U2434 (N_2434,In_357,In_2180);
nor U2435 (N_2435,In_1606,In_2109);
or U2436 (N_2436,In_1562,In_346);
nor U2437 (N_2437,In_1364,In_730);
or U2438 (N_2438,In_2437,In_1503);
and U2439 (N_2439,In_541,In_44);
nand U2440 (N_2440,In_1876,In_377);
nor U2441 (N_2441,In_718,In_1689);
or U2442 (N_2442,In_1354,In_634);
and U2443 (N_2443,In_1971,In_333);
or U2444 (N_2444,In_2470,In_1761);
or U2445 (N_2445,In_1058,In_1087);
or U2446 (N_2446,In_1534,In_2398);
or U2447 (N_2447,In_2139,In_2166);
or U2448 (N_2448,In_2461,In_231);
nor U2449 (N_2449,In_416,In_747);
nor U2450 (N_2450,In_1534,In_1433);
or U2451 (N_2451,In_983,In_479);
nor U2452 (N_2452,In_2026,In_489);
nand U2453 (N_2453,In_755,In_1435);
or U2454 (N_2454,In_866,In_2307);
nand U2455 (N_2455,In_108,In_1138);
or U2456 (N_2456,In_962,In_876);
or U2457 (N_2457,In_1168,In_2067);
or U2458 (N_2458,In_326,In_1037);
nor U2459 (N_2459,In_2201,In_1171);
or U2460 (N_2460,In_1496,In_673);
and U2461 (N_2461,In_1407,In_235);
nor U2462 (N_2462,In_2342,In_2421);
nand U2463 (N_2463,In_800,In_2014);
nand U2464 (N_2464,In_2246,In_1061);
and U2465 (N_2465,In_2096,In_145);
nand U2466 (N_2466,In_252,In_1287);
and U2467 (N_2467,In_96,In_758);
and U2468 (N_2468,In_556,In_786);
nand U2469 (N_2469,In_492,In_1103);
and U2470 (N_2470,In_2001,In_483);
nand U2471 (N_2471,In_2214,In_1869);
nand U2472 (N_2472,In_2042,In_2173);
nor U2473 (N_2473,In_1674,In_1897);
nor U2474 (N_2474,In_2294,In_167);
xor U2475 (N_2475,In_596,In_1241);
nand U2476 (N_2476,In_2170,In_596);
xor U2477 (N_2477,In_1668,In_2484);
nor U2478 (N_2478,In_1781,In_1121);
nand U2479 (N_2479,In_1878,In_710);
or U2480 (N_2480,In_378,In_230);
nand U2481 (N_2481,In_1506,In_1748);
or U2482 (N_2482,In_2102,In_1994);
nor U2483 (N_2483,In_2301,In_860);
nand U2484 (N_2484,In_976,In_285);
or U2485 (N_2485,In_2426,In_109);
and U2486 (N_2486,In_1688,In_266);
nand U2487 (N_2487,In_1748,In_2101);
nand U2488 (N_2488,In_1935,In_2191);
nor U2489 (N_2489,In_2267,In_1981);
or U2490 (N_2490,In_731,In_1502);
nand U2491 (N_2491,In_1439,In_107);
nand U2492 (N_2492,In_283,In_110);
nor U2493 (N_2493,In_352,In_1186);
or U2494 (N_2494,In_1871,In_1687);
nand U2495 (N_2495,In_2002,In_1982);
and U2496 (N_2496,In_1331,In_1938);
and U2497 (N_2497,In_1323,In_1854);
or U2498 (N_2498,In_1116,In_1885);
or U2499 (N_2499,In_2040,In_813);
or U2500 (N_2500,N_27,N_444);
or U2501 (N_2501,N_1632,N_118);
and U2502 (N_2502,N_2402,N_500);
and U2503 (N_2503,N_1221,N_377);
xor U2504 (N_2504,N_2054,N_668);
nand U2505 (N_2505,N_15,N_369);
or U2506 (N_2506,N_1556,N_1521);
or U2507 (N_2507,N_1623,N_215);
and U2508 (N_2508,N_623,N_2274);
or U2509 (N_2509,N_345,N_399);
nor U2510 (N_2510,N_2077,N_539);
nand U2511 (N_2511,N_2017,N_565);
or U2512 (N_2512,N_2168,N_2134);
or U2513 (N_2513,N_419,N_516);
nand U2514 (N_2514,N_1537,N_933);
nand U2515 (N_2515,N_819,N_848);
nor U2516 (N_2516,N_2418,N_1726);
or U2517 (N_2517,N_275,N_1797);
or U2518 (N_2518,N_645,N_2465);
nor U2519 (N_2519,N_1772,N_1816);
nand U2520 (N_2520,N_553,N_10);
nand U2521 (N_2521,N_2308,N_1123);
and U2522 (N_2522,N_1652,N_1165);
nand U2523 (N_2523,N_2412,N_2140);
or U2524 (N_2524,N_1211,N_296);
nor U2525 (N_2525,N_1826,N_420);
xnor U2526 (N_2526,N_899,N_2087);
or U2527 (N_2527,N_380,N_976);
nand U2528 (N_2528,N_1151,N_2332);
nor U2529 (N_2529,N_1161,N_134);
nor U2530 (N_2530,N_1377,N_656);
and U2531 (N_2531,N_418,N_2003);
or U2532 (N_2532,N_1666,N_1212);
and U2533 (N_2533,N_1692,N_1576);
nand U2534 (N_2534,N_1155,N_909);
or U2535 (N_2535,N_403,N_2157);
and U2536 (N_2536,N_2027,N_1599);
nand U2537 (N_2537,N_1657,N_1718);
or U2538 (N_2538,N_2137,N_1146);
nor U2539 (N_2539,N_1822,N_1837);
or U2540 (N_2540,N_635,N_586);
nor U2541 (N_2541,N_889,N_1964);
or U2542 (N_2542,N_35,N_147);
nand U2543 (N_2543,N_2059,N_1640);
and U2544 (N_2544,N_1915,N_942);
and U2545 (N_2545,N_1827,N_1887);
nor U2546 (N_2546,N_96,N_1598);
and U2547 (N_2547,N_626,N_1960);
or U2548 (N_2548,N_1954,N_491);
nor U2549 (N_2549,N_1566,N_1935);
nand U2550 (N_2550,N_852,N_1651);
nor U2551 (N_2551,N_1564,N_965);
and U2552 (N_2552,N_2067,N_2147);
and U2553 (N_2553,N_1514,N_995);
and U2554 (N_2554,N_785,N_524);
and U2555 (N_2555,N_2490,N_1268);
and U2556 (N_2556,N_192,N_2117);
or U2557 (N_2557,N_1644,N_466);
nand U2558 (N_2558,N_2433,N_2251);
and U2559 (N_2559,N_218,N_1531);
nand U2560 (N_2560,N_636,N_238);
or U2561 (N_2561,N_1364,N_347);
or U2562 (N_2562,N_1490,N_1908);
and U2563 (N_2563,N_319,N_1398);
or U2564 (N_2564,N_2124,N_764);
nand U2565 (N_2565,N_1804,N_2065);
nor U2566 (N_2566,N_2101,N_73);
and U2567 (N_2567,N_1931,N_1806);
and U2568 (N_2568,N_2411,N_203);
nor U2569 (N_2569,N_2301,N_484);
or U2570 (N_2570,N_1451,N_61);
or U2571 (N_2571,N_2061,N_430);
nor U2572 (N_2572,N_915,N_564);
nor U2573 (N_2573,N_139,N_1747);
or U2574 (N_2574,N_1259,N_1344);
nand U2575 (N_2575,N_996,N_1184);
or U2576 (N_2576,N_727,N_2189);
nand U2577 (N_2577,N_962,N_1883);
nand U2578 (N_2578,N_1140,N_537);
nand U2579 (N_2579,N_2241,N_2007);
nor U2580 (N_2580,N_1167,N_2123);
nor U2581 (N_2581,N_879,N_724);
and U2582 (N_2582,N_1064,N_1730);
or U2583 (N_2583,N_721,N_1955);
nor U2584 (N_2584,N_1049,N_258);
nor U2585 (N_2585,N_922,N_1611);
or U2586 (N_2586,N_281,N_446);
nor U2587 (N_2587,N_1499,N_1130);
or U2588 (N_2588,N_1902,N_1823);
and U2589 (N_2589,N_2161,N_458);
nor U2590 (N_2590,N_2291,N_1909);
nand U2591 (N_2591,N_2139,N_227);
nand U2592 (N_2592,N_2230,N_1810);
nand U2593 (N_2593,N_2342,N_1843);
nor U2594 (N_2594,N_712,N_1817);
nor U2595 (N_2595,N_1443,N_983);
nand U2596 (N_2596,N_285,N_2167);
nand U2597 (N_2597,N_1467,N_2);
and U2598 (N_2598,N_1127,N_2459);
or U2599 (N_2599,N_1223,N_905);
nor U2600 (N_2600,N_577,N_2265);
nand U2601 (N_2601,N_1191,N_1974);
nand U2602 (N_2602,N_287,N_1097);
nor U2603 (N_2603,N_990,N_1449);
or U2604 (N_2604,N_711,N_1343);
nand U2605 (N_2605,N_1688,N_985);
nand U2606 (N_2606,N_1716,N_177);
nor U2607 (N_2607,N_1637,N_638);
nor U2608 (N_2608,N_1865,N_1094);
or U2609 (N_2609,N_706,N_563);
and U2610 (N_2610,N_988,N_24);
or U2611 (N_2611,N_360,N_1335);
nand U2612 (N_2612,N_2401,N_1358);
and U2613 (N_2613,N_2309,N_2238);
nand U2614 (N_2614,N_286,N_836);
and U2615 (N_2615,N_137,N_1348);
or U2616 (N_2616,N_1007,N_1356);
nand U2617 (N_2617,N_2306,N_621);
nor U2618 (N_2618,N_986,N_2200);
nor U2619 (N_2619,N_2322,N_2236);
nor U2620 (N_2620,N_796,N_1524);
and U2621 (N_2621,N_1267,N_2389);
nor U2622 (N_2622,N_2129,N_291);
and U2623 (N_2623,N_2081,N_1395);
and U2624 (N_2624,N_546,N_1543);
nand U2625 (N_2625,N_1781,N_2156);
or U2626 (N_2626,N_1107,N_517);
nand U2627 (N_2627,N_662,N_1800);
and U2628 (N_2628,N_219,N_1316);
and U2629 (N_2629,N_1446,N_1108);
nor U2630 (N_2630,N_876,N_1409);
or U2631 (N_2631,N_1145,N_17);
and U2632 (N_2632,N_1081,N_1733);
and U2633 (N_2633,N_812,N_1572);
nor U2634 (N_2634,N_186,N_1619);
or U2635 (N_2635,N_261,N_1676);
or U2636 (N_2636,N_1687,N_1038);
or U2637 (N_2637,N_2034,N_1088);
or U2638 (N_2638,N_1922,N_1670);
and U2639 (N_2639,N_1828,N_36);
nand U2640 (N_2640,N_1735,N_1602);
nor U2641 (N_2641,N_1755,N_1963);
or U2642 (N_2642,N_2467,N_1427);
nor U2643 (N_2643,N_200,N_1054);
nor U2644 (N_2644,N_110,N_2035);
nand U2645 (N_2645,N_1762,N_970);
or U2646 (N_2646,N_750,N_1095);
and U2647 (N_2647,N_921,N_181);
or U2648 (N_2648,N_2142,N_95);
and U2649 (N_2649,N_1557,N_20);
nand U2650 (N_2650,N_28,N_531);
and U2651 (N_2651,N_325,N_2350);
or U2652 (N_2652,N_896,N_1340);
or U2653 (N_2653,N_861,N_698);
nor U2654 (N_2654,N_2240,N_805);
or U2655 (N_2655,N_1043,N_741);
nor U2656 (N_2656,N_867,N_734);
or U2657 (N_2657,N_1789,N_2296);
or U2658 (N_2658,N_23,N_1455);
and U2659 (N_2659,N_1590,N_1250);
and U2660 (N_2660,N_1143,N_806);
nand U2661 (N_2661,N_143,N_1737);
nand U2662 (N_2662,N_434,N_590);
nand U2663 (N_2663,N_1849,N_189);
nand U2664 (N_2664,N_2425,N_777);
and U2665 (N_2665,N_1885,N_297);
nor U2666 (N_2666,N_1276,N_1222);
nand U2667 (N_2667,N_328,N_1037);
or U2668 (N_2668,N_766,N_1525);
nand U2669 (N_2669,N_824,N_2318);
nand U2670 (N_2670,N_1458,N_119);
nor U2671 (N_2671,N_1082,N_1937);
nor U2672 (N_2672,N_1175,N_860);
nor U2673 (N_2673,N_30,N_1397);
nor U2674 (N_2674,N_2434,N_1080);
and U2675 (N_2675,N_210,N_199);
nor U2676 (N_2676,N_1195,N_1306);
and U2677 (N_2677,N_594,N_1560);
and U2678 (N_2678,N_1649,N_1493);
and U2679 (N_2679,N_1967,N_1717);
and U2680 (N_2680,N_904,N_1292);
and U2681 (N_2681,N_865,N_1880);
nor U2682 (N_2682,N_1854,N_59);
nor U2683 (N_2683,N_2400,N_1923);
nand U2684 (N_2684,N_846,N_2000);
and U2685 (N_2685,N_87,N_2305);
nand U2686 (N_2686,N_613,N_787);
and U2687 (N_2687,N_1264,N_1940);
nor U2688 (N_2688,N_966,N_1575);
and U2689 (N_2689,N_929,N_994);
or U2690 (N_2690,N_2187,N_88);
nor U2691 (N_2691,N_1247,N_1392);
or U2692 (N_2692,N_1901,N_1630);
nor U2693 (N_2693,N_1607,N_2404);
or U2694 (N_2694,N_1579,N_1819);
nor U2695 (N_2695,N_923,N_982);
and U2696 (N_2696,N_2232,N_483);
or U2697 (N_2697,N_1313,N_1594);
or U2698 (N_2698,N_2104,N_1179);
or U2699 (N_2699,N_574,N_173);
nor U2700 (N_2700,N_804,N_2310);
nor U2701 (N_2701,N_823,N_495);
and U2702 (N_2702,N_841,N_1180);
and U2703 (N_2703,N_522,N_1702);
and U2704 (N_2704,N_1078,N_302);
nor U2705 (N_2705,N_295,N_2431);
nor U2706 (N_2706,N_1609,N_2358);
or U2707 (N_2707,N_1798,N_1552);
nand U2708 (N_2708,N_365,N_2136);
nor U2709 (N_2709,N_1034,N_25);
nor U2710 (N_2710,N_148,N_1587);
or U2711 (N_2711,N_2354,N_2385);
and U2712 (N_2712,N_1787,N_2046);
and U2713 (N_2713,N_1378,N_1041);
and U2714 (N_2714,N_478,N_1251);
nand U2715 (N_2715,N_1706,N_1658);
nand U2716 (N_2716,N_920,N_2337);
or U2717 (N_2717,N_161,N_2379);
nor U2718 (N_2718,N_1421,N_2103);
nor U2719 (N_2719,N_121,N_737);
and U2720 (N_2720,N_1021,N_2351);
nand U2721 (N_2721,N_687,N_2284);
and U2722 (N_2722,N_2100,N_1947);
or U2723 (N_2723,N_2392,N_672);
and U2724 (N_2724,N_1426,N_2215);
xor U2725 (N_2725,N_575,N_1907);
nor U2726 (N_2726,N_2254,N_315);
nor U2727 (N_2727,N_649,N_2173);
nor U2728 (N_2728,N_1488,N_1842);
nor U2729 (N_2729,N_1945,N_443);
and U2730 (N_2730,N_75,N_2032);
nand U2731 (N_2731,N_1695,N_1998);
and U2732 (N_2732,N_1711,N_624);
and U2733 (N_2733,N_1515,N_1198);
or U2734 (N_2734,N_2255,N_2464);
and U2735 (N_2735,N_2393,N_578);
nor U2736 (N_2736,N_12,N_34);
nand U2737 (N_2737,N_414,N_1573);
nand U2738 (N_2738,N_1784,N_1836);
nor U2739 (N_2739,N_2093,N_1805);
nand U2740 (N_2740,N_320,N_1910);
nand U2741 (N_2741,N_1148,N_1675);
nor U2742 (N_2742,N_941,N_957);
or U2743 (N_2743,N_1445,N_1696);
and U2744 (N_2744,N_332,N_1990);
or U2745 (N_2745,N_1079,N_1385);
or U2746 (N_2746,N_1612,N_1035);
or U2747 (N_2747,N_887,N_2458);
nand U2748 (N_2748,N_640,N_870);
nand U2749 (N_2749,N_1319,N_324);
and U2750 (N_2750,N_1355,N_632);
nand U2751 (N_2751,N_748,N_1163);
nand U2752 (N_2752,N_888,N_1884);
and U2753 (N_2753,N_1989,N_445);
xnor U2754 (N_2754,N_386,N_2057);
or U2755 (N_2755,N_664,N_267);
nor U2756 (N_2756,N_1156,N_19);
or U2757 (N_2757,N_784,N_1848);
nand U2758 (N_2758,N_1371,N_2462);
and U2759 (N_2759,N_1863,N_1765);
or U2760 (N_2760,N_2207,N_1460);
nor U2761 (N_2761,N_317,N_1601);
and U2762 (N_2762,N_2429,N_1424);
nor U2763 (N_2763,N_2118,N_2323);
nor U2764 (N_2764,N_205,N_503);
nand U2765 (N_2765,N_908,N_1568);
and U2766 (N_2766,N_2245,N_417);
and U2767 (N_2767,N_874,N_26);
or U2768 (N_2768,N_481,N_81);
or U2769 (N_2769,N_1086,N_112);
nor U2770 (N_2770,N_550,N_1986);
and U2771 (N_2771,N_840,N_385);
nand U2772 (N_2772,N_460,N_329);
and U2773 (N_2773,N_1879,N_1480);
nor U2774 (N_2774,N_2158,N_164);
or U2775 (N_2775,N_2126,N_609);
and U2776 (N_2776,N_1769,N_556);
nor U2777 (N_2777,N_811,N_1932);
nor U2778 (N_2778,N_641,N_1677);
nand U2779 (N_2779,N_371,N_1824);
or U2780 (N_2780,N_396,N_442);
nor U2781 (N_2781,N_1509,N_997);
or U2782 (N_2782,N_92,N_1122);
or U2783 (N_2783,N_1739,N_765);
nand U2784 (N_2784,N_740,N_1936);
or U2785 (N_2785,N_601,N_871);
nand U2786 (N_2786,N_881,N_1431);
nand U2787 (N_2787,N_1109,N_1691);
or U2788 (N_2788,N_1239,N_1604);
or U2789 (N_2789,N_2098,N_381);
nand U2790 (N_2790,N_2013,N_337);
nor U2791 (N_2791,N_1825,N_843);
nor U2792 (N_2792,N_2028,N_1278);
nand U2793 (N_2793,N_470,N_45);
or U2794 (N_2794,N_694,N_447);
and U2795 (N_2795,N_2381,N_1315);
nand U2796 (N_2796,N_1948,N_138);
nand U2797 (N_2797,N_2273,N_1890);
or U2798 (N_2798,N_2179,N_1384);
nand U2799 (N_2799,N_1025,N_2492);
nor U2800 (N_2800,N_1501,N_2446);
or U2801 (N_2801,N_2441,N_1668);
or U2802 (N_2802,N_2432,N_2440);
or U2803 (N_2803,N_1994,N_18);
and U2804 (N_2804,N_1699,N_487);
or U2805 (N_2805,N_2498,N_65);
nor U2806 (N_2806,N_648,N_1969);
nand U2807 (N_2807,N_492,N_1000);
and U2808 (N_2808,N_1546,N_1526);
nand U2809 (N_2809,N_2494,N_428);
nand U2810 (N_2810,N_400,N_663);
nand U2811 (N_2811,N_695,N_171);
or U2812 (N_2812,N_2072,N_815);
nor U2813 (N_2813,N_1654,N_1172);
nand U2814 (N_2814,N_2399,N_1406);
nor U2815 (N_2815,N_828,N_1856);
nor U2816 (N_2816,N_2470,N_1206);
nand U2817 (N_2817,N_555,N_589);
and U2818 (N_2818,N_1513,N_1655);
and U2819 (N_2819,N_616,N_1162);
or U2820 (N_2820,N_105,N_989);
nor U2821 (N_2821,N_977,N_1063);
or U2822 (N_2822,N_141,N_2019);
and U2823 (N_2823,N_1149,N_2331);
and U2824 (N_2824,N_1775,N_72);
or U2825 (N_2825,N_1917,N_1820);
nor U2826 (N_2826,N_1983,N_469);
nand U2827 (N_2827,N_390,N_407);
and U2828 (N_2828,N_1510,N_1382);
nor U2829 (N_2829,N_2480,N_591);
or U2830 (N_2830,N_13,N_1438);
or U2831 (N_2831,N_2461,N_475);
nor U2832 (N_2832,N_2010,N_751);
nand U2833 (N_2833,N_859,N_2218);
or U2834 (N_2834,N_439,N_2338);
and U2835 (N_2835,N_1815,N_212);
or U2836 (N_2836,N_1582,N_1190);
nand U2837 (N_2837,N_2194,N_1920);
nor U2838 (N_2838,N_596,N_64);
nand U2839 (N_2839,N_731,N_2293);
or U2840 (N_2840,N_236,N_1299);
nor U2841 (N_2841,N_827,N_1927);
or U2842 (N_2842,N_1567,N_2479);
nor U2843 (N_2843,N_2279,N_50);
nand U2844 (N_2844,N_2031,N_1921);
nand U2845 (N_2845,N_704,N_2085);
and U2846 (N_2846,N_728,N_1878);
xor U2847 (N_2847,N_2290,N_1485);
nand U2848 (N_2848,N_508,N_2112);
and U2849 (N_2849,N_167,N_674);
and U2850 (N_2850,N_1158,N_2324);
and U2851 (N_2851,N_2343,N_1024);
nor U2852 (N_2852,N_1432,N_2030);
xor U2853 (N_2853,N_1653,N_1913);
nor U2854 (N_2854,N_154,N_1011);
nand U2855 (N_2855,N_2113,N_845);
or U2856 (N_2856,N_82,N_778);
or U2857 (N_2857,N_1408,N_321);
and U2858 (N_2858,N_1896,N_1099);
nand U2859 (N_2859,N_802,N_2415);
or U2860 (N_2860,N_1217,N_204);
and U2861 (N_2861,N_2280,N_561);
and U2862 (N_2862,N_2396,N_607);
nor U2863 (N_2863,N_1183,N_2233);
and U2864 (N_2864,N_697,N_2210);
nor U2865 (N_2865,N_2130,N_615);
or U2866 (N_2866,N_1850,N_1282);
nand U2867 (N_2867,N_851,N_552);
nand U2868 (N_2868,N_630,N_2481);
and U2869 (N_2869,N_1115,N_981);
nor U2870 (N_2870,N_1214,N_357);
and U2871 (N_2871,N_1229,N_758);
nand U2872 (N_2872,N_467,N_1864);
or U2873 (N_2873,N_2105,N_683);
or U2874 (N_2874,N_1366,N_145);
nand U2875 (N_2875,N_1561,N_196);
or U2876 (N_2876,N_1578,N_1574);
xnor U2877 (N_2877,N_1996,N_1357);
nand U2878 (N_2878,N_1293,N_2363);
nor U2879 (N_2879,N_776,N_979);
and U2880 (N_2880,N_1629,N_974);
and U2881 (N_2881,N_1110,N_625);
nor U2882 (N_2882,N_643,N_2227);
nor U2883 (N_2883,N_1396,N_432);
and U2884 (N_2884,N_2212,N_1656);
xnor U2885 (N_2885,N_1465,N_1502);
nor U2886 (N_2886,N_898,N_1372);
nor U2887 (N_2887,N_1703,N_441);
nor U2888 (N_2888,N_2313,N_1202);
nor U2889 (N_2889,N_2430,N_506);
nand U2890 (N_2890,N_2316,N_1142);
or U2891 (N_2891,N_256,N_125);
nand U2892 (N_2892,N_2048,N_1489);
nor U2893 (N_2893,N_2082,N_2219);
and U2894 (N_2894,N_333,N_1059);
or U2895 (N_2895,N_251,N_426);
and U2896 (N_2896,N_1724,N_1219);
or U2897 (N_2897,N_1006,N_2473);
or U2898 (N_2898,N_1709,N_1633);
or U2899 (N_2899,N_1417,N_991);
and U2900 (N_2900,N_661,N_2277);
nor U2901 (N_2901,N_1550,N_1121);
or U2902 (N_2902,N_1470,N_1616);
and U2903 (N_2903,N_462,N_1428);
nand U2904 (N_2904,N_583,N_1416);
nor U2905 (N_2905,N_1518,N_2149);
and U2906 (N_2906,N_2224,N_1591);
nand U2907 (N_2907,N_844,N_1814);
nand U2908 (N_2908,N_5,N_311);
or U2909 (N_2909,N_891,N_1138);
nand U2910 (N_2910,N_1708,N_2190);
nor U2911 (N_2911,N_1533,N_1694);
and U2912 (N_2912,N_2336,N_700);
or U2913 (N_2913,N_2202,N_207);
and U2914 (N_2914,N_310,N_1505);
nand U2915 (N_2915,N_1205,N_2371);
or U2916 (N_2916,N_33,N_789);
nor U2917 (N_2917,N_193,N_1734);
and U2918 (N_2918,N_1131,N_2246);
or U2919 (N_2919,N_1862,N_937);
nor U2920 (N_2920,N_2300,N_2199);
or U2921 (N_2921,N_2299,N_1453);
nor U2922 (N_2922,N_980,N_1437);
nand U2923 (N_2923,N_2203,N_1005);
nand U2924 (N_2924,N_2420,N_397);
nor U2925 (N_2925,N_2269,N_2133);
nand U2926 (N_2926,N_1341,N_330);
nor U2927 (N_2927,N_2115,N_998);
nand U2928 (N_2928,N_2042,N_1643);
nand U2929 (N_2929,N_1628,N_352);
and U2930 (N_2930,N_886,N_1022);
and U2931 (N_2931,N_1646,N_464);
or U2932 (N_2932,N_652,N_1106);
and U2933 (N_2933,N_1727,N_1273);
or U2934 (N_2934,N_919,N_2406);
nor U2935 (N_2935,N_169,N_1089);
or U2936 (N_2936,N_2275,N_1196);
and U2937 (N_2937,N_80,N_975);
or U2938 (N_2938,N_1622,N_1295);
or U2939 (N_2939,N_43,N_717);
and U2940 (N_2940,N_653,N_158);
nor U2941 (N_2941,N_705,N_1995);
nand U2942 (N_2942,N_1980,N_1203);
nor U2943 (N_2943,N_1867,N_1301);
nor U2944 (N_2944,N_437,N_1855);
nand U2945 (N_2945,N_903,N_2395);
and U2946 (N_2946,N_1271,N_1234);
nor U2947 (N_2947,N_832,N_755);
nand U2948 (N_2948,N_1066,N_71);
and U2949 (N_2949,N_378,N_2315);
and U2950 (N_2950,N_1905,N_538);
and U2951 (N_2951,N_1351,N_1484);
or U2952 (N_2952,N_1984,N_1725);
nand U2953 (N_2953,N_1197,N_350);
and U2954 (N_2954,N_1053,N_2008);
or U2955 (N_2955,N_725,N_2195);
or U2956 (N_2956,N_2049,N_584);
nand U2957 (N_2957,N_912,N_1710);
nand U2958 (N_2958,N_2029,N_1997);
nor U2959 (N_2959,N_1238,N_2497);
and U2960 (N_2960,N_1736,N_2486);
nand U2961 (N_2961,N_2416,N_2225);
nor U2962 (N_2962,N_140,N_91);
nor U2963 (N_2963,N_108,N_1635);
nor U2964 (N_2964,N_1926,N_739);
or U2965 (N_2965,N_1152,N_452);
nor U2966 (N_2966,N_754,N_526);
xor U2967 (N_2967,N_402,N_160);
or U2968 (N_2968,N_1390,N_2272);
nand U2969 (N_2969,N_1128,N_1934);
and U2970 (N_2970,N_1585,N_1311);
and U2971 (N_2971,N_1471,N_2078);
or U2972 (N_2972,N_2159,N_2214);
and U2973 (N_2973,N_566,N_334);
or U2974 (N_2974,N_322,N_1407);
xnor U2975 (N_2975,N_132,N_969);
nand U2976 (N_2976,N_1778,N_298);
or U2977 (N_2977,N_31,N_883);
or U2978 (N_2978,N_106,N_2005);
nor U2979 (N_2979,N_1215,N_1410);
and U2980 (N_2980,N_1853,N_797);
xor U2981 (N_2981,N_1388,N_2022);
and U2982 (N_2982,N_2009,N_480);
and U2983 (N_2983,N_1729,N_367);
and U2984 (N_2984,N_703,N_849);
nor U2985 (N_2985,N_1845,N_2438);
or U2986 (N_2986,N_1678,N_1260);
nor U2987 (N_2987,N_2346,N_2033);
and U2988 (N_2988,N_567,N_1768);
and U2989 (N_2989,N_128,N_55);
nand U2990 (N_2990,N_1500,N_289);
nand U2991 (N_2991,N_628,N_463);
or U2992 (N_2992,N_608,N_1009);
nor U2993 (N_2993,N_1369,N_2347);
or U2994 (N_2994,N_2261,N_8);
nor U2995 (N_2995,N_304,N_2483);
and U2996 (N_2996,N_2015,N_2319);
nand U2997 (N_2997,N_1044,N_1199);
and U2998 (N_2998,N_1999,N_1096);
and U2999 (N_2999,N_1182,N_1617);
nor U3000 (N_3000,N_2169,N_280);
nand U3001 (N_3001,N_2355,N_1791);
nand U3002 (N_3002,N_234,N_2160);
nand U3003 (N_3003,N_175,N_2307);
nor U3004 (N_3004,N_52,N_425);
or U3005 (N_3005,N_2119,N_1770);
and U3006 (N_3006,N_1120,N_2239);
nor U3007 (N_3007,N_149,N_1783);
and U3008 (N_3008,N_1930,N_2079);
nand U3009 (N_3009,N_2417,N_1051);
nand U3010 (N_3010,N_2452,N_1661);
and U3011 (N_3011,N_6,N_512);
or U3012 (N_3012,N_1608,N_1134);
nor U3013 (N_3013,N_472,N_1244);
nor U3014 (N_3014,N_1425,N_489);
nand U3015 (N_3015,N_681,N_1365);
nand U3016 (N_3016,N_2468,N_44);
or U3017 (N_3017,N_2234,N_479);
and U3018 (N_3018,N_1101,N_2256);
nand U3019 (N_3019,N_1627,N_326);
nor U3020 (N_3020,N_340,N_1168);
and U3021 (N_3021,N_809,N_1338);
nand U3022 (N_3022,N_1209,N_1474);
or U3023 (N_3023,N_792,N_958);
or U3024 (N_3024,N_1660,N_545);
nor U3025 (N_3025,N_927,N_2055);
nand U3026 (N_3026,N_675,N_1394);
nor U3027 (N_3027,N_1400,N_1329);
nand U3028 (N_3028,N_429,N_2180);
nor U3029 (N_3029,N_216,N_422);
or U3030 (N_3030,N_2171,N_1799);
nand U3031 (N_3031,N_1801,N_2356);
nor U3032 (N_3032,N_1283,N_274);
and U3033 (N_3033,N_1452,N_1634);
nor U3034 (N_3034,N_2349,N_14);
nand U3035 (N_3035,N_2360,N_1777);
and U3036 (N_3036,N_781,N_499);
nor U3037 (N_3037,N_2127,N_37);
nor U3038 (N_3038,N_1869,N_934);
and U3039 (N_3039,N_74,N_1565);
nor U3040 (N_3040,N_928,N_948);
and U3041 (N_3041,N_1056,N_2089);
and U3042 (N_3042,N_2083,N_1322);
nand U3043 (N_3043,N_372,N_1188);
nand U3044 (N_3044,N_551,N_932);
and U3045 (N_3045,N_42,N_901);
nand U3046 (N_3046,N_264,N_1133);
nor U3047 (N_3047,N_2177,N_246);
and U3048 (N_3048,N_2334,N_1174);
and U3049 (N_3049,N_1528,N_1411);
and U3050 (N_3050,N_1118,N_972);
and U3051 (N_3051,N_1979,N_1893);
nand U3052 (N_3052,N_745,N_292);
or U3053 (N_3053,N_943,N_486);
nand U3054 (N_3054,N_2150,N_2053);
nand U3055 (N_3055,N_1918,N_202);
and U3056 (N_3056,N_1705,N_129);
and U3057 (N_3057,N_1257,N_1636);
nand U3058 (N_3058,N_956,N_293);
or U3059 (N_3059,N_877,N_678);
nand U3060 (N_3060,N_2128,N_671);
nand U3061 (N_3061,N_834,N_1559);
xor U3062 (N_3062,N_1423,N_1262);
nand U3063 (N_3063,N_2038,N_2437);
or U3064 (N_3064,N_254,N_2264);
or U3065 (N_3065,N_1898,N_973);
and U3066 (N_3066,N_2253,N_1642);
nor U3067 (N_3067,N_391,N_992);
nor U3068 (N_3068,N_1912,N_1779);
and U3069 (N_3069,N_1650,N_1686);
and U3070 (N_3070,N_1792,N_89);
or U3071 (N_3071,N_497,N_2326);
or U3072 (N_3072,N_2228,N_944);
nand U3073 (N_3073,N_1889,N_122);
and U3074 (N_3074,N_2320,N_2155);
or U3075 (N_3075,N_2397,N_1712);
nand U3076 (N_3076,N_156,N_351);
nor U3077 (N_3077,N_1857,N_1418);
and U3078 (N_3078,N_1925,N_1040);
or U3079 (N_3079,N_309,N_2243);
or U3080 (N_3080,N_252,N_894);
or U3081 (N_3081,N_1753,N_2178);
and U3082 (N_3082,N_90,N_1227);
nor U3083 (N_3083,N_1665,N_642);
or U3084 (N_3084,N_2110,N_1332);
and U3085 (N_3085,N_2353,N_709);
and U3086 (N_3086,N_895,N_1263);
nor U3087 (N_3087,N_1403,N_2281);
and U3088 (N_3088,N_1373,N_631);
and U3089 (N_3089,N_2023,N_339);
nor U3090 (N_3090,N_1065,N_810);
or U3091 (N_3091,N_1284,N_971);
or U3092 (N_3092,N_2044,N_2466);
nor U3093 (N_3093,N_78,N_2176);
and U3094 (N_3094,N_97,N_902);
nor U3095 (N_3095,N_690,N_762);
and U3096 (N_3096,N_245,N_2317);
or U3097 (N_3097,N_1129,N_1952);
or U3098 (N_3098,N_1200,N_1220);
nand U3099 (N_3099,N_1057,N_1639);
or U3100 (N_3100,N_501,N_1210);
and U3101 (N_3101,N_1113,N_1742);
or U3102 (N_3102,N_1583,N_1468);
or U3103 (N_3103,N_768,N_1874);
or U3104 (N_3104,N_2040,N_2493);
nor U3105 (N_3105,N_1353,N_1046);
nor U3106 (N_3106,N_1914,N_960);
and U3107 (N_3107,N_1968,N_1136);
and U3108 (N_3108,N_135,N_782);
or U3109 (N_3109,N_255,N_1977);
nand U3110 (N_3110,N_1176,N_1897);
and U3111 (N_3111,N_98,N_1192);
nor U3112 (N_3112,N_2052,N_2476);
and U3113 (N_3113,N_1303,N_165);
or U3114 (N_3114,N_159,N_1389);
or U3115 (N_3115,N_1457,N_1962);
and U3116 (N_3116,N_162,N_4);
nor U3117 (N_3117,N_788,N_814);
or U3118 (N_3118,N_1087,N_1571);
or U3119 (N_3119,N_411,N_598);
nor U3120 (N_3120,N_906,N_1255);
nor U3121 (N_3121,N_1307,N_1071);
or U3122 (N_3122,N_614,N_1933);
and U3123 (N_3123,N_510,N_498);
and U3124 (N_3124,N_779,N_2114);
and U3125 (N_3125,N_1281,N_799);
and U3126 (N_3126,N_1846,N_2063);
or U3127 (N_3127,N_370,N_2444);
nand U3128 (N_3128,N_606,N_1405);
nor U3129 (N_3129,N_2454,N_1462);
and U3130 (N_3130,N_2002,N_1744);
and U3131 (N_3131,N_1434,N_465);
nand U3132 (N_3132,N_2201,N_1669);
and U3133 (N_3133,N_468,N_2378);
and U3134 (N_3134,N_84,N_240);
nand U3135 (N_3135,N_406,N_47);
and U3136 (N_3136,N_729,N_423);
and U3137 (N_3137,N_247,N_1906);
nor U3138 (N_3138,N_243,N_1216);
nor U3139 (N_3139,N_416,N_1361);
nor U3140 (N_3140,N_2367,N_892);
nor U3141 (N_3141,N_1834,N_16);
nand U3142 (N_3142,N_837,N_1254);
nand U3143 (N_3143,N_1667,N_2384);
nor U3144 (N_3144,N_507,N_244);
and U3145 (N_3145,N_576,N_2436);
nor U3146 (N_3146,N_2448,N_1596);
nor U3147 (N_3147,N_1645,N_1439);
or U3148 (N_3148,N_1868,N_2365);
nor U3149 (N_3149,N_1350,N_1697);
nor U3150 (N_3150,N_228,N_1334);
and U3151 (N_3151,N_2182,N_677);
or U3152 (N_3152,N_2191,N_1504);
nor U3153 (N_3153,N_914,N_1558);
nor U3154 (N_3154,N_1886,N_774);
and U3155 (N_3155,N_2152,N_76);
or U3156 (N_3156,N_890,N_2036);
or U3157 (N_3157,N_2143,N_1472);
nor U3158 (N_3158,N_1626,N_2186);
and U3159 (N_3159,N_1756,N_21);
nor U3160 (N_3160,N_820,N_346);
nand U3161 (N_3161,N_808,N_1758);
or U3162 (N_3162,N_176,N_2193);
or U3163 (N_3163,N_1833,N_272);
or U3164 (N_3164,N_1252,N_825);
nand U3165 (N_3165,N_2455,N_450);
or U3166 (N_3166,N_1750,N_1683);
nor U3167 (N_3167,N_1105,N_595);
and U3168 (N_3168,N_1551,N_1320);
nor U3169 (N_3169,N_67,N_211);
or U3170 (N_3170,N_716,N_1562);
or U3171 (N_3171,N_669,N_1008);
nand U3172 (N_3172,N_363,N_126);
nor U3173 (N_3173,N_2388,N_2226);
and U3174 (N_3174,N_693,N_1720);
or U3175 (N_3175,N_673,N_83);
or U3176 (N_3176,N_952,N_2447);
nand U3177 (N_3177,N_651,N_884);
nor U3178 (N_3178,N_253,N_2428);
nand U3179 (N_3179,N_257,N_573);
nor U3180 (N_3180,N_830,N_786);
nor U3181 (N_3181,N_2321,N_2145);
xor U3182 (N_3182,N_1987,N_1847);
and U3183 (N_3183,N_713,N_770);
nand U3184 (N_3184,N_155,N_1871);
and U3185 (N_3185,N_682,N_1852);
nand U3186 (N_3186,N_622,N_1363);
or U3187 (N_3187,N_448,N_1305);
and U3188 (N_3188,N_514,N_2086);
nand U3189 (N_3189,N_847,N_2080);
or U3190 (N_3190,N_93,N_1224);
and U3191 (N_3191,N_1116,N_2341);
nor U3192 (N_3192,N_1530,N_527);
or U3193 (N_3193,N_1153,N_1185);
nand U3194 (N_3194,N_686,N_471);
nor U3195 (N_3195,N_144,N_2267);
or U3196 (N_3196,N_354,N_1336);
and U3197 (N_3197,N_1018,N_2407);
nor U3198 (N_3198,N_736,N_1304);
and U3199 (N_3199,N_1872,N_2376);
or U3200 (N_3200,N_1554,N_1290);
and U3201 (N_3201,N_451,N_835);
nor U3202 (N_3202,N_1519,N_117);
or U3203 (N_3203,N_1698,N_230);
or U3204 (N_3204,N_599,N_1256);
and U3205 (N_3205,N_1597,N_2165);
nor U3206 (N_3206,N_1641,N_1542);
or U3207 (N_3207,N_1939,N_1821);
and U3208 (N_3208,N_60,N_1137);
nand U3209 (N_3209,N_1570,N_2469);
nor U3210 (N_3210,N_2163,N_1141);
or U3211 (N_3211,N_2237,N_178);
nand U3212 (N_3212,N_967,N_54);
nand U3213 (N_3213,N_2423,N_1548);
nor U3214 (N_3214,N_1535,N_1166);
nor U3215 (N_3215,N_232,N_1840);
or U3216 (N_3216,N_1296,N_1068);
nor U3217 (N_3217,N_1589,N_2120);
nor U3218 (N_3218,N_1838,N_107);
nor U3219 (N_3219,N_842,N_1859);
or U3220 (N_3220,N_1039,N_1782);
or U3221 (N_3221,N_2174,N_2047);
and U3222 (N_3222,N_1072,N_1988);
and U3223 (N_3223,N_1061,N_57);
or U3224 (N_3224,N_111,N_826);
nor U3225 (N_3225,N_1581,N_2285);
nand U3226 (N_3226,N_1595,N_38);
and U3227 (N_3227,N_123,N_1052);
nor U3228 (N_3228,N_548,N_917);
or U3229 (N_3229,N_2102,N_2183);
or U3230 (N_3230,N_897,N_1337);
or U3231 (N_3231,N_109,N_250);
and U3232 (N_3232,N_679,N_866);
and U3233 (N_3233,N_2056,N_1045);
and U3234 (N_3234,N_494,N_1790);
nor U3235 (N_3235,N_1444,N_1246);
nor U3236 (N_3236,N_582,N_1966);
and U3237 (N_3237,N_2244,N_213);
nor U3238 (N_3238,N_1312,N_560);
and U3239 (N_3239,N_769,N_49);
and U3240 (N_3240,N_999,N_2312);
nor U3241 (N_3241,N_1342,N_1208);
and U3242 (N_3242,N_1701,N_1728);
and U3243 (N_3243,N_1436,N_1684);
or U3244 (N_3244,N_336,N_277);
nor U3245 (N_3245,N_1461,N_341);
and U3246 (N_3246,N_2491,N_1985);
nand U3247 (N_3247,N_39,N_2252);
nand U3248 (N_3248,N_744,N_2097);
or U3249 (N_3249,N_493,N_1359);
nand U3250 (N_3250,N_2220,N_1830);
and U3251 (N_3251,N_720,N_2456);
nor U3252 (N_3252,N_1613,N_900);
nand U3253 (N_3253,N_831,N_1492);
nand U3254 (N_3254,N_1620,N_1013);
nor U3255 (N_3255,N_699,N_1555);
nor U3256 (N_3256,N_726,N_1091);
and U3257 (N_3257,N_1938,N_1959);
nor U3258 (N_3258,N_2460,N_1415);
nand U3259 (N_3259,N_485,N_2146);
and U3260 (N_3260,N_627,N_1139);
and U3261 (N_3261,N_2108,N_558);
nand U3262 (N_3262,N_511,N_1807);
or U3263 (N_3263,N_231,N_667);
nand U3264 (N_3264,N_1346,N_2141);
or U3265 (N_3265,N_654,N_1508);
or U3266 (N_3266,N_666,N_1347);
and U3267 (N_3267,N_759,N_133);
nand U3268 (N_3268,N_1147,N_525);
and U3269 (N_3269,N_2278,N_2025);
or U3270 (N_3270,N_2472,N_1982);
nand U3271 (N_3271,N_1272,N_938);
nor U3272 (N_3272,N_2068,N_646);
or U3273 (N_3273,N_1181,N_1261);
and U3274 (N_3274,N_283,N_1333);
nor U3275 (N_3275,N_343,N_2096);
nor U3276 (N_3276,N_1473,N_1248);
nor U3277 (N_3277,N_1456,N_276);
or U3278 (N_3278,N_1788,N_359);
or U3279 (N_3279,N_1861,N_1682);
nand U3280 (N_3280,N_2495,N_1506);
nand U3281 (N_3281,N_619,N_1159);
or U3282 (N_3282,N_1092,N_2289);
nand U3283 (N_3283,N_1903,N_2205);
and U3284 (N_3284,N_356,N_536);
nor U3285 (N_3285,N_2424,N_1536);
nand U3286 (N_3286,N_1387,N_94);
nor U3287 (N_3287,N_839,N_1186);
or U3288 (N_3288,N_303,N_361);
nand U3289 (N_3289,N_2014,N_1029);
nand U3290 (N_3290,N_1527,N_2394);
nor U3291 (N_3291,N_1615,N_1380);
or U3292 (N_3292,N_1475,N_543);
nand U3293 (N_3293,N_344,N_103);
and U3294 (N_3294,N_1318,N_562);
and U3295 (N_3295,N_1793,N_1279);
nand U3296 (N_3296,N_1478,N_1230);
nor U3297 (N_3297,N_1760,N_1813);
nor U3298 (N_3298,N_771,N_1391);
nor U3299 (N_3299,N_1073,N_70);
and U3300 (N_3300,N_2297,N_1370);
and U3301 (N_3301,N_541,N_1873);
nor U3302 (N_3302,N_1839,N_2421);
nor U3303 (N_3303,N_680,N_1638);
nand U3304 (N_3304,N_1614,N_338);
nor U3305 (N_3305,N_2192,N_637);
or U3306 (N_3306,N_2386,N_1228);
nand U3307 (N_3307,N_780,N_2362);
nand U3308 (N_3308,N_1098,N_634);
or U3309 (N_3309,N_2018,N_1876);
or U3310 (N_3310,N_719,N_1420);
or U3311 (N_3311,N_1266,N_882);
nor U3312 (N_3312,N_1412,N_1844);
nor U3313 (N_3313,N_104,N_335);
and U3314 (N_3314,N_2478,N_9);
nor U3315 (N_3315,N_312,N_1715);
or U3316 (N_3316,N_197,N_453);
or U3317 (N_3317,N_1911,N_821);
nand U3318 (N_3318,N_2172,N_1719);
or U3319 (N_3319,N_41,N_1647);
nor U3320 (N_3320,N_1811,N_659);
or U3321 (N_3321,N_1189,N_327);
or U3322 (N_3322,N_1077,N_2325);
nor U3323 (N_3323,N_1012,N_858);
and U3324 (N_3324,N_323,N_1067);
and U3325 (N_3325,N_916,N_689);
nor U3326 (N_3326,N_1992,N_1961);
or U3327 (N_3327,N_603,N_1941);
and U3328 (N_3328,N_1740,N_1360);
or U3329 (N_3329,N_2075,N_1624);
nand U3330 (N_3330,N_2196,N_658);
and U3331 (N_3331,N_409,N_150);
nor U3332 (N_3332,N_29,N_735);
nor U3333 (N_3333,N_1763,N_523);
and U3334 (N_3334,N_760,N_410);
and U3335 (N_3335,N_413,N_875);
or U3336 (N_3336,N_2229,N_2099);
and U3337 (N_3337,N_2069,N_925);
nor U3338 (N_3338,N_1464,N_801);
or U3339 (N_3339,N_1060,N_2304);
nand U3340 (N_3340,N_743,N_602);
nor U3341 (N_3341,N_1204,N_440);
or U3342 (N_3342,N_893,N_2107);
or U3343 (N_3343,N_353,N_2294);
nor U3344 (N_3344,N_1076,N_1243);
or U3345 (N_3345,N_1331,N_790);
and U3346 (N_3346,N_557,N_1386);
and U3347 (N_3347,N_1036,N_1144);
nor U3348 (N_3348,N_2335,N_696);
nand U3349 (N_3349,N_191,N_2131);
nand U3350 (N_3350,N_1956,N_157);
nand U3351 (N_3351,N_1310,N_220);
and U3352 (N_3352,N_1891,N_174);
and U3353 (N_3353,N_63,N_209);
nand U3354 (N_3354,N_504,N_182);
or U3355 (N_3355,N_1,N_1083);
and U3356 (N_3356,N_1368,N_168);
nor U3357 (N_3357,N_1447,N_362);
nand U3358 (N_3358,N_1659,N_532);
and U3359 (N_3359,N_1330,N_2004);
and U3360 (N_3360,N_2154,N_1308);
and U3361 (N_3361,N_457,N_2361);
nor U3362 (N_3362,N_542,N_733);
or U3363 (N_3363,N_554,N_954);
nand U3364 (N_3364,N_963,N_146);
and U3365 (N_3365,N_2039,N_1981);
or U3366 (N_3366,N_1592,N_1732);
and U3367 (N_3367,N_455,N_872);
xnor U3368 (N_3368,N_2148,N_1808);
nand U3369 (N_3369,N_2208,N_271);
nor U3370 (N_3370,N_1454,N_2377);
nand U3371 (N_3371,N_48,N_1606);
nor U3372 (N_3372,N_2050,N_2135);
nand U3373 (N_3373,N_136,N_2216);
and U3374 (N_3374,N_2062,N_803);
nand U3375 (N_3375,N_1497,N_142);
nand U3376 (N_3376,N_249,N_723);
and U3377 (N_3377,N_2153,N_2164);
nor U3378 (N_3378,N_505,N_1942);
nor U3379 (N_3379,N_284,N_730);
or U3380 (N_3380,N_949,N_1731);
nor U3381 (N_3381,N_2398,N_2181);
nor U3382 (N_3382,N_163,N_130);
or U3383 (N_3383,N_1253,N_2463);
nor U3384 (N_3384,N_1381,N_408);
nand U3385 (N_3385,N_2374,N_2314);
or U3386 (N_3386,N_2211,N_2016);
nand U3387 (N_3387,N_1831,N_1047);
and U3388 (N_3388,N_746,N_1523);
or U3389 (N_3389,N_1754,N_1245);
and U3390 (N_3390,N_2410,N_384);
or U3391 (N_3391,N_710,N_331);
nand U3392 (N_3392,N_2475,N_2166);
and U3393 (N_3393,N_2288,N_1401);
nor U3394 (N_3394,N_1588,N_40);
and U3395 (N_3395,N_714,N_807);
and U3396 (N_3396,N_1766,N_223);
or U3397 (N_3397,N_795,N_1469);
nand U3398 (N_3398,N_2286,N_1780);
or U3399 (N_3399,N_270,N_833);
nand U3400 (N_3400,N_1916,N_863);
nor U3401 (N_3401,N_862,N_1539);
or U3402 (N_3402,N_1503,N_1544);
and U3403 (N_3403,N_1795,N_2001);
and U3404 (N_3404,N_2064,N_1419);
and U3405 (N_3405,N_1714,N_1476);
nand U3406 (N_3406,N_2344,N_1631);
and U3407 (N_3407,N_1707,N_2443);
and U3408 (N_3408,N_229,N_1680);
nor U3409 (N_3409,N_1786,N_588);
nand U3410 (N_3410,N_685,N_1111);
nor U3411 (N_3411,N_2058,N_1402);
nand U3412 (N_3412,N_1976,N_950);
nand U3413 (N_3413,N_1028,N_1949);
and U3414 (N_3414,N_568,N_1553);
or U3415 (N_3415,N_1441,N_856);
or U3416 (N_3416,N_1538,N_388);
or U3417 (N_3417,N_1662,N_1430);
or U3418 (N_3418,N_692,N_1383);
nand U3419 (N_3419,N_1679,N_1818);
and U3420 (N_3420,N_482,N_1213);
nand U3421 (N_3421,N_2248,N_1177);
nand U3422 (N_3422,N_1953,N_1802);
and U3423 (N_3423,N_1399,N_2283);
nand U3424 (N_3424,N_2427,N_1157);
nor U3425 (N_3425,N_1745,N_349);
nor U3426 (N_3426,N_102,N_2387);
nor U3427 (N_3427,N_1033,N_918);
nand U3428 (N_3428,N_300,N_152);
nor U3429 (N_3429,N_854,N_1300);
or U3430 (N_3430,N_0,N_1055);
nand U3431 (N_3431,N_2184,N_850);
and U3432 (N_3432,N_940,N_931);
or U3433 (N_3433,N_1674,N_2144);
and U3434 (N_3434,N_2408,N_570);
nand U3435 (N_3435,N_1170,N_1090);
nand U3436 (N_3436,N_2024,N_1015);
or U3437 (N_3437,N_1103,N_1442);
or U3438 (N_3438,N_1761,N_2380);
nor U3439 (N_3439,N_2037,N_2084);
or U3440 (N_3440,N_1114,N_2329);
and U3441 (N_3441,N_2073,N_1746);
or U3442 (N_3442,N_1882,N_1748);
nor U3443 (N_3443,N_533,N_1314);
xor U3444 (N_3444,N_1031,N_1738);
xor U3445 (N_3445,N_1413,N_1017);
and U3446 (N_3446,N_579,N_530);
nand U3447 (N_3447,N_822,N_2422);
and U3448 (N_3448,N_1904,N_1970);
and U3449 (N_3449,N_124,N_1541);
and U3450 (N_3450,N_395,N_911);
nor U3451 (N_3451,N_355,N_2383);
nor U3452 (N_3452,N_1440,N_398);
and U3453 (N_3453,N_2066,N_1841);
or U3454 (N_3454,N_2262,N_800);
and U3455 (N_3455,N_2204,N_521);
nor U3456 (N_3456,N_1362,N_1280);
nand U3457 (N_3457,N_1625,N_1759);
and U3458 (N_3458,N_655,N_1194);
or U3459 (N_3459,N_2247,N_959);
nand U3460 (N_3460,N_1580,N_77);
or U3461 (N_3461,N_2151,N_1093);
nand U3462 (N_3462,N_2287,N_1429);
or U3463 (N_3463,N_732,N_2041);
xor U3464 (N_3464,N_978,N_1352);
nand U3465 (N_3465,N_113,N_2327);
and U3466 (N_3466,N_1529,N_509);
and U3467 (N_3467,N_2043,N_597);
or U3468 (N_3468,N_376,N_593);
or U3469 (N_3469,N_282,N_2094);
nor U3470 (N_3470,N_620,N_1773);
nor U3471 (N_3471,N_2328,N_936);
nand U3472 (N_3472,N_534,N_2026);
nand U3473 (N_3473,N_1771,N_1483);
and U3474 (N_3474,N_1258,N_670);
nand U3475 (N_3475,N_1002,N_2175);
and U3476 (N_3476,N_853,N_515);
and U3477 (N_3477,N_2071,N_1743);
and U3478 (N_3478,N_1374,N_1102);
nand U3479 (N_3479,N_241,N_513);
and U3480 (N_3480,N_366,N_657);
and U3481 (N_3481,N_235,N_459);
or U3482 (N_3482,N_1232,N_2197);
or U3483 (N_3483,N_187,N_1178);
nand U3484 (N_3484,N_206,N_518);
nor U3485 (N_3485,N_1367,N_1605);
and U3486 (N_3486,N_1870,N_559);
nor U3487 (N_3487,N_1124,N_2090);
and U3488 (N_3488,N_1023,N_798);
nor U3489 (N_3489,N_955,N_600);
nor U3490 (N_3490,N_1950,N_2271);
nand U3491 (N_3491,N_427,N_1349);
nand U3492 (N_3492,N_1899,N_2260);
nand U3493 (N_3493,N_2345,N_2414);
and U3494 (N_3494,N_1671,N_1577);
nor U3495 (N_3495,N_1858,N_1171);
nor U3496 (N_3496,N_2330,N_738);
and U3497 (N_3497,N_2132,N_2045);
nand U3498 (N_3498,N_375,N_2450);
nand U3499 (N_3499,N_885,N_1235);
nand U3500 (N_3500,N_951,N_308);
and U3501 (N_3501,N_2250,N_1586);
or U3502 (N_3502,N_1540,N_436);
and U3503 (N_3503,N_2382,N_421);
and U3504 (N_3504,N_1294,N_2368);
and U3505 (N_3505,N_1003,N_405);
or U3506 (N_3506,N_1971,N_2348);
or U3507 (N_3507,N_1919,N_1241);
and U3508 (N_3508,N_924,N_188);
nor U3509 (N_3509,N_1603,N_2170);
or U3510 (N_3510,N_1242,N_1563);
nand U3511 (N_3511,N_260,N_1048);
or U3512 (N_3512,N_2257,N_639);
or U3513 (N_3513,N_1302,N_69);
or U3514 (N_3514,N_1112,N_1160);
or U3515 (N_3515,N_1693,N_1298);
nor U3516 (N_3516,N_1991,N_2070);
nand U3517 (N_3517,N_2372,N_572);
or U3518 (N_3518,N_629,N_1713);
or U3519 (N_3519,N_166,N_454);
nor U3520 (N_3520,N_1723,N_294);
nor U3521 (N_3521,N_1327,N_1965);
nand U3522 (N_3522,N_2298,N_198);
nor U3523 (N_3523,N_585,N_2409);
and U3524 (N_3524,N_502,N_1975);
or U3525 (N_3525,N_647,N_1532);
or U3526 (N_3526,N_816,N_1275);
and U3527 (N_3527,N_1104,N_1317);
nor U3528 (N_3528,N_431,N_569);
or U3529 (N_3529,N_2266,N_2076);
nand U3530 (N_3530,N_2249,N_2453);
or U3531 (N_3531,N_587,N_1498);
nand U3532 (N_3532,N_387,N_939);
nand U3533 (N_3533,N_520,N_1477);
nand U3534 (N_3534,N_1285,N_101);
and U3535 (N_3535,N_2217,N_1119);
nor U3536 (N_3536,N_611,N_2333);
or U3537 (N_3537,N_873,N_1972);
nor U3538 (N_3538,N_1721,N_2403);
and U3539 (N_3539,N_1325,N_767);
nand U3540 (N_3540,N_1062,N_314);
or U3541 (N_3541,N_1495,N_32);
or U3542 (N_3542,N_773,N_1240);
nand U3543 (N_3543,N_829,N_299);
or U3544 (N_3544,N_262,N_2485);
nand U3545 (N_3545,N_389,N_1001);
and U3546 (N_3546,N_2373,N_46);
or U3547 (N_3547,N_1010,N_2391);
nand U3548 (N_3548,N_2445,N_435);
or U3549 (N_3549,N_2021,N_11);
nor U3550 (N_3550,N_1032,N_1881);
nand U3551 (N_3551,N_183,N_2357);
nand U3552 (N_3552,N_68,N_519);
nor U3553 (N_3553,N_127,N_2340);
or U3554 (N_3554,N_404,N_438);
nor U3555 (N_3555,N_763,N_179);
xor U3556 (N_3556,N_412,N_1004);
and U3557 (N_3557,N_1757,N_813);
and U3558 (N_3558,N_1339,N_2116);
nand U3559 (N_3559,N_1117,N_214);
nor U3560 (N_3560,N_2375,N_1681);
nand U3561 (N_3561,N_1100,N_1274);
and U3562 (N_3562,N_1450,N_2242);
nor U3563 (N_3563,N_794,N_424);
nand U3564 (N_3564,N_263,N_1075);
or U3565 (N_3565,N_747,N_358);
or U3566 (N_3566,N_1835,N_259);
nor U3567 (N_3567,N_702,N_2222);
or U3568 (N_3568,N_1448,N_783);
nor U3569 (N_3569,N_1479,N_1900);
or U3570 (N_3570,N_1225,N_935);
nor U3571 (N_3571,N_1866,N_2074);
and U3572 (N_3572,N_1809,N_342);
nor U3573 (N_3573,N_757,N_1375);
and U3574 (N_3574,N_1481,N_753);
nand U3575 (N_3575,N_2020,N_305);
and U3576 (N_3576,N_1020,N_1026);
nand U3577 (N_3577,N_2258,N_2484);
nor U3578 (N_3578,N_461,N_749);
nor U3579 (N_3579,N_946,N_544);
nor U3580 (N_3580,N_279,N_217);
nand U3581 (N_3581,N_1741,N_791);
and U3582 (N_3582,N_401,N_2051);
and U3583 (N_3583,N_2303,N_1875);
nor U3584 (N_3584,N_1764,N_592);
or U3585 (N_3585,N_1796,N_1265);
nor U3586 (N_3586,N_318,N_868);
nor U3587 (N_3587,N_1321,N_1751);
nand U3588 (N_3588,N_1832,N_1135);
xnor U3589 (N_3589,N_2442,N_2435);
nand U3590 (N_3590,N_1892,N_225);
nand U3591 (N_3591,N_857,N_1496);
nor U3592 (N_3592,N_99,N_2419);
and U3593 (N_3593,N_3,N_1328);
nand U3594 (N_3594,N_1685,N_1672);
nand U3595 (N_3595,N_1511,N_1042);
or U3596 (N_3596,N_772,N_1767);
and U3597 (N_3597,N_496,N_131);
nand U3598 (N_3598,N_1154,N_1749);
nor U3599 (N_3599,N_2359,N_53);
nand U3600 (N_3600,N_1928,N_1610);
nand U3601 (N_3601,N_2449,N_2477);
and U3602 (N_3602,N_2496,N_268);
nand U3603 (N_3603,N_691,N_1414);
nand U3604 (N_3604,N_2339,N_1016);
and U3605 (N_3605,N_581,N_1877);
nand U3606 (N_3606,N_761,N_393);
nor U3607 (N_3607,N_718,N_1648);
nand U3608 (N_3608,N_151,N_1584);
and U3609 (N_3609,N_618,N_266);
or U3610 (N_3610,N_1704,N_2263);
nor U3611 (N_3611,N_817,N_650);
and U3612 (N_3612,N_374,N_1459);
and U3613 (N_3613,N_1978,N_2213);
or U3614 (N_3614,N_301,N_1569);
nand U3615 (N_3615,N_1664,N_2292);
nor U3616 (N_3616,N_383,N_2482);
and U3617 (N_3617,N_1169,N_474);
nand U3618 (N_3618,N_2457,N_456);
nor U3619 (N_3619,N_1074,N_1226);
and U3620 (N_3620,N_2106,N_701);
nor U3621 (N_3621,N_1323,N_490);
or U3622 (N_3622,N_1277,N_1058);
nor U3623 (N_3623,N_617,N_1309);
and U3624 (N_3624,N_968,N_2413);
or U3625 (N_3625,N_1973,N_2276);
nor U3626 (N_3626,N_1466,N_2011);
and U3627 (N_3627,N_2295,N_549);
and U3628 (N_3628,N_290,N_2426);
nand U3629 (N_3629,N_1173,N_273);
and U3630 (N_3630,N_1236,N_1520);
nand U3631 (N_3631,N_612,N_58);
nor U3632 (N_3632,N_855,N_547);
nand U3633 (N_3633,N_265,N_1486);
xor U3634 (N_3634,N_1069,N_1785);
or U3635 (N_3635,N_184,N_1700);
nand U3636 (N_3636,N_433,N_1993);
nor U3637 (N_3637,N_708,N_633);
nand U3638 (N_3638,N_987,N_1132);
or U3639 (N_3639,N_1794,N_208);
nand U3640 (N_3640,N_2499,N_2390);
nor U3641 (N_3641,N_1291,N_2091);
nor U3642 (N_3642,N_2221,N_476);
nor U3643 (N_3643,N_2370,N_1233);
and U3644 (N_3644,N_1376,N_115);
or U3645 (N_3645,N_477,N_529);
and U3646 (N_3646,N_1435,N_1270);
or U3647 (N_3647,N_1354,N_2125);
nor U3648 (N_3648,N_221,N_2439);
nand U3649 (N_3649,N_1482,N_910);
nand U3650 (N_3650,N_1288,N_864);
nand U3651 (N_3651,N_1125,N_1201);
nor U3652 (N_3652,N_2122,N_1326);
nand U3653 (N_3653,N_1237,N_2109);
and U3654 (N_3654,N_1929,N_2209);
nor U3655 (N_3655,N_1289,N_153);
and U3656 (N_3656,N_348,N_1673);
nand U3657 (N_3657,N_170,N_1324);
and U3658 (N_3658,N_2092,N_1516);
xor U3659 (N_3659,N_379,N_313);
or U3660 (N_3660,N_239,N_1621);
and U3661 (N_3661,N_316,N_2471);
nand U3662 (N_3662,N_878,N_1894);
nand U3663 (N_3663,N_373,N_1269);
and U3664 (N_3664,N_22,N_1860);
nor U3665 (N_3665,N_237,N_7);
nor U3666 (N_3666,N_288,N_660);
and U3667 (N_3667,N_880,N_2352);
nor U3668 (N_3668,N_1463,N_226);
nand U3669 (N_3669,N_528,N_1600);
and U3670 (N_3670,N_1851,N_488);
or U3671 (N_3671,N_1297,N_2235);
nand U3672 (N_3672,N_1164,N_201);
nand U3673 (N_3673,N_2369,N_85);
nand U3674 (N_3674,N_2088,N_644);
or U3675 (N_3675,N_1545,N_2268);
and U3676 (N_3676,N_1084,N_1050);
or U3677 (N_3677,N_930,N_1776);
nor U3678 (N_3678,N_1404,N_1433);
nand U3679 (N_3679,N_1019,N_2231);
and U3680 (N_3680,N_1287,N_2198);
nor U3681 (N_3681,N_2282,N_1689);
nor U3682 (N_3682,N_2060,N_62);
and U3683 (N_3683,N_1957,N_610);
and U3684 (N_3684,N_1193,N_233);
and U3685 (N_3685,N_172,N_1774);
or U3686 (N_3686,N_1085,N_2111);
nor U3687 (N_3687,N_2474,N_1187);
or U3688 (N_3688,N_120,N_676);
nand U3689 (N_3689,N_1491,N_913);
or U3690 (N_3690,N_604,N_382);
or U3691 (N_3691,N_1014,N_926);
nand U3692 (N_3692,N_1507,N_100);
nand U3693 (N_3693,N_86,N_1924);
nor U3694 (N_3694,N_1379,N_79);
nor U3695 (N_3695,N_1888,N_2366);
and U3696 (N_3696,N_945,N_2405);
or U3697 (N_3697,N_1812,N_869);
and U3698 (N_3698,N_993,N_1752);
nand U3699 (N_3699,N_775,N_394);
and U3700 (N_3700,N_1207,N_688);
nor U3701 (N_3701,N_269,N_1895);
nor U3702 (N_3702,N_1618,N_2095);
and U3703 (N_3703,N_1722,N_368);
nor U3704 (N_3704,N_114,N_1946);
nor U3705 (N_3705,N_1422,N_180);
and U3706 (N_3706,N_415,N_306);
nand U3707 (N_3707,N_278,N_953);
nor U3708 (N_3708,N_742,N_838);
and U3709 (N_3709,N_947,N_1150);
or U3710 (N_3710,N_2223,N_242);
nor U3711 (N_3711,N_1218,N_2364);
or U3712 (N_3712,N_2206,N_1249);
or U3713 (N_3713,N_984,N_793);
nand U3714 (N_3714,N_1690,N_307);
and U3715 (N_3715,N_194,N_1126);
nor U3716 (N_3716,N_1517,N_1027);
nor U3717 (N_3717,N_605,N_1593);
or U3718 (N_3718,N_66,N_1951);
nor U3719 (N_3719,N_571,N_665);
and U3720 (N_3720,N_684,N_1070);
nor U3721 (N_3721,N_392,N_248);
nand U3722 (N_3722,N_364,N_1829);
xor U3723 (N_3723,N_2138,N_195);
and U3724 (N_3724,N_1534,N_2302);
and U3725 (N_3725,N_185,N_707);
or U3726 (N_3726,N_2012,N_2311);
and U3727 (N_3727,N_535,N_2259);
and U3728 (N_3728,N_190,N_961);
nand U3729 (N_3729,N_756,N_116);
or U3730 (N_3730,N_2488,N_2270);
nand U3731 (N_3731,N_1803,N_449);
and U3732 (N_3732,N_222,N_818);
or U3733 (N_3733,N_2451,N_715);
nor U3734 (N_3734,N_1231,N_540);
nand U3735 (N_3735,N_1494,N_1549);
and U3736 (N_3736,N_722,N_51);
nand U3737 (N_3737,N_1547,N_1286);
or U3738 (N_3738,N_2006,N_1030);
nor U3739 (N_3739,N_1345,N_1487);
nand U3740 (N_3740,N_964,N_1393);
or U3741 (N_3741,N_2185,N_1944);
nor U3742 (N_3742,N_1512,N_1663);
nand U3743 (N_3743,N_224,N_2162);
and U3744 (N_3744,N_2489,N_2487);
nand U3745 (N_3745,N_2188,N_2121);
nor U3746 (N_3746,N_1943,N_580);
nor U3747 (N_3747,N_907,N_1958);
nand U3748 (N_3748,N_752,N_473);
nand U3749 (N_3749,N_56,N_1522);
nor U3750 (N_3750,N_642,N_2255);
nor U3751 (N_3751,N_1509,N_627);
and U3752 (N_3752,N_2368,N_307);
nand U3753 (N_3753,N_2329,N_1528);
nor U3754 (N_3754,N_1654,N_1534);
nor U3755 (N_3755,N_171,N_2491);
and U3756 (N_3756,N_492,N_1704);
nor U3757 (N_3757,N_1228,N_1265);
and U3758 (N_3758,N_1743,N_1857);
and U3759 (N_3759,N_2188,N_1763);
nand U3760 (N_3760,N_1128,N_2128);
nor U3761 (N_3761,N_1780,N_1561);
and U3762 (N_3762,N_1103,N_307);
or U3763 (N_3763,N_1031,N_646);
or U3764 (N_3764,N_656,N_140);
nand U3765 (N_3765,N_2484,N_1654);
or U3766 (N_3766,N_2465,N_72);
nand U3767 (N_3767,N_1043,N_869);
or U3768 (N_3768,N_2372,N_1846);
and U3769 (N_3769,N_792,N_706);
nor U3770 (N_3770,N_1122,N_2276);
and U3771 (N_3771,N_1331,N_1268);
nand U3772 (N_3772,N_816,N_654);
nor U3773 (N_3773,N_1695,N_819);
and U3774 (N_3774,N_753,N_401);
and U3775 (N_3775,N_1576,N_2447);
or U3776 (N_3776,N_315,N_1931);
or U3777 (N_3777,N_1002,N_1310);
and U3778 (N_3778,N_1555,N_2345);
nand U3779 (N_3779,N_2224,N_319);
nand U3780 (N_3780,N_1442,N_2469);
nand U3781 (N_3781,N_1135,N_1788);
nand U3782 (N_3782,N_2150,N_1502);
xor U3783 (N_3783,N_302,N_2219);
nor U3784 (N_3784,N_1234,N_144);
nand U3785 (N_3785,N_225,N_549);
or U3786 (N_3786,N_145,N_413);
nor U3787 (N_3787,N_1063,N_337);
xor U3788 (N_3788,N_465,N_1022);
nor U3789 (N_3789,N_1075,N_1697);
nor U3790 (N_3790,N_1361,N_1004);
or U3791 (N_3791,N_1371,N_2257);
or U3792 (N_3792,N_2486,N_38);
or U3793 (N_3793,N_2085,N_1708);
nor U3794 (N_3794,N_945,N_2059);
or U3795 (N_3795,N_741,N_1875);
or U3796 (N_3796,N_750,N_2225);
nand U3797 (N_3797,N_520,N_981);
nor U3798 (N_3798,N_1472,N_1579);
and U3799 (N_3799,N_1045,N_1201);
nor U3800 (N_3800,N_294,N_624);
nor U3801 (N_3801,N_2234,N_853);
or U3802 (N_3802,N_198,N_302);
nor U3803 (N_3803,N_714,N_250);
nor U3804 (N_3804,N_2420,N_447);
and U3805 (N_3805,N_1678,N_1900);
and U3806 (N_3806,N_2102,N_1628);
or U3807 (N_3807,N_2184,N_280);
nand U3808 (N_3808,N_1370,N_1955);
nand U3809 (N_3809,N_787,N_1589);
nand U3810 (N_3810,N_1269,N_2480);
nand U3811 (N_3811,N_14,N_566);
or U3812 (N_3812,N_1538,N_1419);
and U3813 (N_3813,N_1849,N_884);
or U3814 (N_3814,N_1176,N_1179);
or U3815 (N_3815,N_398,N_123);
or U3816 (N_3816,N_1615,N_409);
or U3817 (N_3817,N_2224,N_1011);
nor U3818 (N_3818,N_2368,N_1180);
nand U3819 (N_3819,N_1573,N_2095);
and U3820 (N_3820,N_744,N_1467);
and U3821 (N_3821,N_485,N_2105);
and U3822 (N_3822,N_1695,N_1662);
nand U3823 (N_3823,N_1811,N_2267);
and U3824 (N_3824,N_1590,N_685);
and U3825 (N_3825,N_1528,N_1473);
and U3826 (N_3826,N_403,N_2212);
nand U3827 (N_3827,N_1009,N_138);
nor U3828 (N_3828,N_467,N_1619);
or U3829 (N_3829,N_56,N_293);
or U3830 (N_3830,N_2023,N_832);
and U3831 (N_3831,N_867,N_1557);
nand U3832 (N_3832,N_768,N_2173);
nor U3833 (N_3833,N_407,N_287);
nand U3834 (N_3834,N_201,N_2496);
and U3835 (N_3835,N_426,N_1248);
or U3836 (N_3836,N_244,N_94);
nor U3837 (N_3837,N_522,N_76);
nand U3838 (N_3838,N_2199,N_1728);
xnor U3839 (N_3839,N_205,N_1048);
or U3840 (N_3840,N_1294,N_351);
or U3841 (N_3841,N_1913,N_1271);
nor U3842 (N_3842,N_2380,N_1892);
nor U3843 (N_3843,N_1015,N_1148);
and U3844 (N_3844,N_571,N_462);
nor U3845 (N_3845,N_664,N_549);
or U3846 (N_3846,N_1655,N_1828);
and U3847 (N_3847,N_221,N_88);
and U3848 (N_3848,N_156,N_2414);
or U3849 (N_3849,N_1303,N_1539);
or U3850 (N_3850,N_1563,N_1486);
and U3851 (N_3851,N_1722,N_1154);
and U3852 (N_3852,N_2009,N_2027);
nand U3853 (N_3853,N_1407,N_640);
or U3854 (N_3854,N_1964,N_1318);
and U3855 (N_3855,N_2200,N_1884);
nor U3856 (N_3856,N_1109,N_1876);
nand U3857 (N_3857,N_1876,N_304);
nand U3858 (N_3858,N_1699,N_1758);
or U3859 (N_3859,N_1272,N_2124);
or U3860 (N_3860,N_1229,N_1281);
nor U3861 (N_3861,N_1145,N_2050);
nor U3862 (N_3862,N_156,N_699);
nand U3863 (N_3863,N_2362,N_1462);
and U3864 (N_3864,N_1167,N_1561);
or U3865 (N_3865,N_1087,N_1934);
nand U3866 (N_3866,N_1526,N_2039);
nor U3867 (N_3867,N_173,N_2430);
or U3868 (N_3868,N_870,N_1648);
or U3869 (N_3869,N_217,N_1815);
nor U3870 (N_3870,N_421,N_1668);
and U3871 (N_3871,N_144,N_1712);
xnor U3872 (N_3872,N_2357,N_472);
or U3873 (N_3873,N_1515,N_146);
or U3874 (N_3874,N_2041,N_2314);
or U3875 (N_3875,N_591,N_469);
and U3876 (N_3876,N_1061,N_431);
and U3877 (N_3877,N_1782,N_1318);
nand U3878 (N_3878,N_2122,N_2332);
and U3879 (N_3879,N_1837,N_805);
nor U3880 (N_3880,N_1042,N_1519);
and U3881 (N_3881,N_525,N_1089);
xnor U3882 (N_3882,N_2214,N_1253);
nor U3883 (N_3883,N_595,N_2196);
and U3884 (N_3884,N_1496,N_1150);
nand U3885 (N_3885,N_678,N_796);
and U3886 (N_3886,N_1858,N_1595);
nor U3887 (N_3887,N_2141,N_1440);
or U3888 (N_3888,N_1828,N_933);
or U3889 (N_3889,N_1255,N_1351);
nand U3890 (N_3890,N_513,N_780);
nand U3891 (N_3891,N_1933,N_1471);
nor U3892 (N_3892,N_1169,N_2208);
and U3893 (N_3893,N_702,N_899);
xnor U3894 (N_3894,N_1338,N_1858);
or U3895 (N_3895,N_587,N_474);
or U3896 (N_3896,N_2315,N_1467);
nand U3897 (N_3897,N_2396,N_726);
nor U3898 (N_3898,N_714,N_1917);
nor U3899 (N_3899,N_1233,N_1216);
nor U3900 (N_3900,N_2384,N_207);
nor U3901 (N_3901,N_1691,N_741);
or U3902 (N_3902,N_1756,N_1740);
or U3903 (N_3903,N_1558,N_2217);
nand U3904 (N_3904,N_401,N_2124);
or U3905 (N_3905,N_2332,N_1561);
nor U3906 (N_3906,N_1829,N_1530);
and U3907 (N_3907,N_974,N_772);
or U3908 (N_3908,N_2089,N_1571);
or U3909 (N_3909,N_45,N_1995);
or U3910 (N_3910,N_560,N_2173);
nand U3911 (N_3911,N_954,N_111);
nor U3912 (N_3912,N_1043,N_2089);
nor U3913 (N_3913,N_2448,N_747);
or U3914 (N_3914,N_1918,N_2373);
nor U3915 (N_3915,N_1795,N_502);
nand U3916 (N_3916,N_2259,N_1864);
nor U3917 (N_3917,N_1078,N_1266);
or U3918 (N_3918,N_112,N_1972);
or U3919 (N_3919,N_1608,N_2195);
or U3920 (N_3920,N_1208,N_958);
nor U3921 (N_3921,N_1,N_1532);
and U3922 (N_3922,N_2483,N_224);
and U3923 (N_3923,N_1837,N_1986);
or U3924 (N_3924,N_1994,N_357);
or U3925 (N_3925,N_1651,N_1286);
or U3926 (N_3926,N_560,N_1339);
nor U3927 (N_3927,N_307,N_240);
nand U3928 (N_3928,N_1103,N_1308);
and U3929 (N_3929,N_971,N_517);
nor U3930 (N_3930,N_1953,N_1101);
nand U3931 (N_3931,N_1228,N_972);
or U3932 (N_3932,N_1321,N_2496);
or U3933 (N_3933,N_755,N_2023);
or U3934 (N_3934,N_2310,N_55);
nor U3935 (N_3935,N_1044,N_2293);
or U3936 (N_3936,N_851,N_1007);
nand U3937 (N_3937,N_1703,N_1872);
nand U3938 (N_3938,N_797,N_167);
nand U3939 (N_3939,N_2379,N_2433);
nor U3940 (N_3940,N_1510,N_1573);
and U3941 (N_3941,N_2054,N_1692);
and U3942 (N_3942,N_1716,N_375);
nor U3943 (N_3943,N_1564,N_2354);
nor U3944 (N_3944,N_360,N_1942);
nor U3945 (N_3945,N_73,N_2475);
and U3946 (N_3946,N_767,N_772);
nand U3947 (N_3947,N_538,N_1658);
nor U3948 (N_3948,N_481,N_196);
nor U3949 (N_3949,N_2220,N_1496);
or U3950 (N_3950,N_495,N_2337);
or U3951 (N_3951,N_868,N_1922);
nand U3952 (N_3952,N_582,N_1738);
or U3953 (N_3953,N_855,N_1798);
nor U3954 (N_3954,N_2384,N_2069);
nand U3955 (N_3955,N_351,N_2271);
and U3956 (N_3956,N_787,N_49);
or U3957 (N_3957,N_2424,N_920);
nor U3958 (N_3958,N_1680,N_2135);
nor U3959 (N_3959,N_2320,N_142);
nor U3960 (N_3960,N_141,N_603);
and U3961 (N_3961,N_1302,N_2142);
nand U3962 (N_3962,N_94,N_993);
and U3963 (N_3963,N_2108,N_1946);
nor U3964 (N_3964,N_922,N_1212);
or U3965 (N_3965,N_264,N_240);
nand U3966 (N_3966,N_1202,N_2282);
nor U3967 (N_3967,N_1619,N_2326);
and U3968 (N_3968,N_756,N_910);
nand U3969 (N_3969,N_2015,N_2260);
or U3970 (N_3970,N_332,N_908);
or U3971 (N_3971,N_921,N_1505);
and U3972 (N_3972,N_2086,N_1541);
nand U3973 (N_3973,N_1453,N_1563);
and U3974 (N_3974,N_1010,N_1931);
nand U3975 (N_3975,N_772,N_1902);
nor U3976 (N_3976,N_2411,N_159);
and U3977 (N_3977,N_486,N_325);
nor U3978 (N_3978,N_171,N_2293);
or U3979 (N_3979,N_2289,N_1392);
and U3980 (N_3980,N_1323,N_1422);
nor U3981 (N_3981,N_1381,N_768);
nand U3982 (N_3982,N_707,N_66);
nand U3983 (N_3983,N_2346,N_1421);
nand U3984 (N_3984,N_68,N_252);
or U3985 (N_3985,N_1431,N_1250);
nor U3986 (N_3986,N_936,N_1580);
or U3987 (N_3987,N_1283,N_1204);
and U3988 (N_3988,N_584,N_1512);
and U3989 (N_3989,N_1528,N_952);
or U3990 (N_3990,N_1823,N_1027);
or U3991 (N_3991,N_168,N_2014);
nor U3992 (N_3992,N_1886,N_718);
or U3993 (N_3993,N_1954,N_194);
and U3994 (N_3994,N_1119,N_1567);
and U3995 (N_3995,N_2340,N_1637);
or U3996 (N_3996,N_2130,N_2223);
nand U3997 (N_3997,N_108,N_881);
nand U3998 (N_3998,N_1609,N_1448);
nand U3999 (N_3999,N_865,N_159);
nand U4000 (N_4000,N_45,N_538);
and U4001 (N_4001,N_32,N_2147);
and U4002 (N_4002,N_527,N_1069);
nor U4003 (N_4003,N_828,N_1044);
or U4004 (N_4004,N_1619,N_1090);
nand U4005 (N_4005,N_50,N_1873);
nand U4006 (N_4006,N_657,N_2426);
nor U4007 (N_4007,N_700,N_882);
or U4008 (N_4008,N_1652,N_2053);
nand U4009 (N_4009,N_2277,N_1088);
and U4010 (N_4010,N_2496,N_674);
nor U4011 (N_4011,N_656,N_1700);
or U4012 (N_4012,N_126,N_802);
nor U4013 (N_4013,N_1406,N_632);
or U4014 (N_4014,N_2330,N_512);
or U4015 (N_4015,N_1878,N_993);
nor U4016 (N_4016,N_1148,N_1448);
xor U4017 (N_4017,N_930,N_148);
or U4018 (N_4018,N_312,N_1770);
nand U4019 (N_4019,N_1441,N_1256);
nor U4020 (N_4020,N_1452,N_197);
nand U4021 (N_4021,N_89,N_2055);
nand U4022 (N_4022,N_1738,N_2186);
or U4023 (N_4023,N_2397,N_435);
nor U4024 (N_4024,N_1197,N_684);
or U4025 (N_4025,N_1258,N_1214);
nor U4026 (N_4026,N_1865,N_1368);
nor U4027 (N_4027,N_593,N_1245);
or U4028 (N_4028,N_2464,N_190);
and U4029 (N_4029,N_450,N_1056);
and U4030 (N_4030,N_1364,N_1178);
nand U4031 (N_4031,N_1881,N_402);
nor U4032 (N_4032,N_1021,N_1978);
and U4033 (N_4033,N_562,N_1814);
and U4034 (N_4034,N_1134,N_2159);
and U4035 (N_4035,N_1212,N_75);
or U4036 (N_4036,N_512,N_1557);
nand U4037 (N_4037,N_528,N_1993);
or U4038 (N_4038,N_1854,N_2293);
nor U4039 (N_4039,N_1081,N_825);
and U4040 (N_4040,N_2082,N_2180);
nor U4041 (N_4041,N_2274,N_1030);
or U4042 (N_4042,N_2424,N_1369);
and U4043 (N_4043,N_2295,N_1130);
or U4044 (N_4044,N_1079,N_2435);
or U4045 (N_4045,N_411,N_129);
nand U4046 (N_4046,N_1932,N_156);
nor U4047 (N_4047,N_1679,N_219);
or U4048 (N_4048,N_950,N_1506);
and U4049 (N_4049,N_2314,N_785);
and U4050 (N_4050,N_23,N_2074);
or U4051 (N_4051,N_2419,N_2047);
and U4052 (N_4052,N_601,N_1206);
or U4053 (N_4053,N_955,N_1836);
nor U4054 (N_4054,N_1242,N_570);
and U4055 (N_4055,N_1863,N_1555);
nand U4056 (N_4056,N_1191,N_697);
and U4057 (N_4057,N_1774,N_1074);
nand U4058 (N_4058,N_1034,N_288);
nand U4059 (N_4059,N_865,N_1746);
or U4060 (N_4060,N_1943,N_1156);
nand U4061 (N_4061,N_291,N_222);
and U4062 (N_4062,N_2231,N_1423);
nand U4063 (N_4063,N_1145,N_797);
and U4064 (N_4064,N_665,N_975);
and U4065 (N_4065,N_1343,N_605);
nor U4066 (N_4066,N_2499,N_1217);
nor U4067 (N_4067,N_2481,N_365);
nor U4068 (N_4068,N_466,N_2002);
nand U4069 (N_4069,N_458,N_2288);
and U4070 (N_4070,N_1466,N_183);
and U4071 (N_4071,N_2302,N_2203);
nand U4072 (N_4072,N_1908,N_1798);
or U4073 (N_4073,N_2303,N_876);
and U4074 (N_4074,N_356,N_1549);
nand U4075 (N_4075,N_1990,N_1371);
or U4076 (N_4076,N_2062,N_2291);
and U4077 (N_4077,N_100,N_1399);
nor U4078 (N_4078,N_1071,N_1162);
and U4079 (N_4079,N_940,N_901);
and U4080 (N_4080,N_1858,N_195);
or U4081 (N_4081,N_833,N_67);
or U4082 (N_4082,N_2294,N_949);
and U4083 (N_4083,N_1679,N_1290);
nand U4084 (N_4084,N_943,N_1290);
nand U4085 (N_4085,N_1806,N_1025);
or U4086 (N_4086,N_734,N_1058);
nor U4087 (N_4087,N_818,N_1785);
or U4088 (N_4088,N_377,N_1573);
and U4089 (N_4089,N_1298,N_2056);
and U4090 (N_4090,N_137,N_413);
nand U4091 (N_4091,N_1734,N_1524);
nor U4092 (N_4092,N_433,N_1533);
nor U4093 (N_4093,N_835,N_838);
nand U4094 (N_4094,N_2247,N_730);
nor U4095 (N_4095,N_631,N_1178);
and U4096 (N_4096,N_813,N_2320);
nor U4097 (N_4097,N_788,N_1295);
and U4098 (N_4098,N_1611,N_856);
or U4099 (N_4099,N_656,N_502);
or U4100 (N_4100,N_1553,N_1494);
nor U4101 (N_4101,N_1679,N_765);
nand U4102 (N_4102,N_2107,N_51);
nand U4103 (N_4103,N_1219,N_2165);
and U4104 (N_4104,N_767,N_67);
nand U4105 (N_4105,N_257,N_10);
nor U4106 (N_4106,N_1422,N_2302);
nand U4107 (N_4107,N_1054,N_425);
and U4108 (N_4108,N_271,N_2290);
and U4109 (N_4109,N_264,N_774);
nand U4110 (N_4110,N_2306,N_1334);
xor U4111 (N_4111,N_1294,N_2463);
or U4112 (N_4112,N_852,N_1477);
nor U4113 (N_4113,N_566,N_424);
nor U4114 (N_4114,N_1608,N_2335);
or U4115 (N_4115,N_1504,N_1897);
or U4116 (N_4116,N_623,N_1220);
nand U4117 (N_4117,N_1970,N_136);
or U4118 (N_4118,N_738,N_39);
nor U4119 (N_4119,N_1586,N_2147);
or U4120 (N_4120,N_1688,N_2345);
and U4121 (N_4121,N_2202,N_2311);
and U4122 (N_4122,N_1267,N_2050);
nand U4123 (N_4123,N_1646,N_1260);
nor U4124 (N_4124,N_1385,N_2407);
or U4125 (N_4125,N_1578,N_1245);
nand U4126 (N_4126,N_2006,N_216);
nor U4127 (N_4127,N_932,N_1084);
nand U4128 (N_4128,N_1719,N_2184);
nand U4129 (N_4129,N_2431,N_252);
or U4130 (N_4130,N_1390,N_1320);
nand U4131 (N_4131,N_146,N_1690);
and U4132 (N_4132,N_828,N_513);
nand U4133 (N_4133,N_1790,N_1882);
and U4134 (N_4134,N_952,N_438);
or U4135 (N_4135,N_1028,N_1120);
and U4136 (N_4136,N_1287,N_1590);
or U4137 (N_4137,N_1598,N_1515);
or U4138 (N_4138,N_1304,N_1994);
and U4139 (N_4139,N_26,N_256);
nand U4140 (N_4140,N_1098,N_1870);
and U4141 (N_4141,N_420,N_1736);
nand U4142 (N_4142,N_806,N_1498);
nand U4143 (N_4143,N_2400,N_2403);
or U4144 (N_4144,N_919,N_1026);
or U4145 (N_4145,N_730,N_1133);
and U4146 (N_4146,N_1252,N_1539);
nor U4147 (N_4147,N_2233,N_2287);
and U4148 (N_4148,N_1655,N_1588);
and U4149 (N_4149,N_1650,N_166);
nor U4150 (N_4150,N_1433,N_2249);
nor U4151 (N_4151,N_806,N_550);
or U4152 (N_4152,N_1406,N_218);
or U4153 (N_4153,N_1425,N_1535);
nand U4154 (N_4154,N_1461,N_583);
nor U4155 (N_4155,N_262,N_1505);
nand U4156 (N_4156,N_326,N_2047);
and U4157 (N_4157,N_414,N_492);
nor U4158 (N_4158,N_1601,N_1858);
nor U4159 (N_4159,N_444,N_877);
nor U4160 (N_4160,N_597,N_58);
nand U4161 (N_4161,N_70,N_1268);
nand U4162 (N_4162,N_1953,N_79);
nand U4163 (N_4163,N_1920,N_2090);
or U4164 (N_4164,N_327,N_1682);
or U4165 (N_4165,N_567,N_1637);
nor U4166 (N_4166,N_1946,N_1786);
and U4167 (N_4167,N_2408,N_2348);
or U4168 (N_4168,N_1486,N_1525);
or U4169 (N_4169,N_1924,N_1726);
and U4170 (N_4170,N_750,N_1663);
or U4171 (N_4171,N_353,N_1694);
and U4172 (N_4172,N_1165,N_2227);
nor U4173 (N_4173,N_2405,N_2017);
and U4174 (N_4174,N_1180,N_1086);
nor U4175 (N_4175,N_243,N_343);
nor U4176 (N_4176,N_448,N_2264);
nand U4177 (N_4177,N_1566,N_2211);
or U4178 (N_4178,N_846,N_650);
nand U4179 (N_4179,N_861,N_80);
and U4180 (N_4180,N_425,N_2196);
nand U4181 (N_4181,N_1690,N_2334);
or U4182 (N_4182,N_1113,N_1998);
or U4183 (N_4183,N_1140,N_995);
and U4184 (N_4184,N_2219,N_2065);
and U4185 (N_4185,N_1385,N_1630);
nor U4186 (N_4186,N_2418,N_1406);
or U4187 (N_4187,N_943,N_2392);
or U4188 (N_4188,N_359,N_1696);
and U4189 (N_4189,N_2442,N_2321);
and U4190 (N_4190,N_1256,N_170);
nand U4191 (N_4191,N_1775,N_1295);
nand U4192 (N_4192,N_847,N_242);
and U4193 (N_4193,N_696,N_2438);
nor U4194 (N_4194,N_1123,N_907);
and U4195 (N_4195,N_485,N_2402);
and U4196 (N_4196,N_423,N_1726);
or U4197 (N_4197,N_573,N_1691);
and U4198 (N_4198,N_140,N_2232);
or U4199 (N_4199,N_723,N_476);
and U4200 (N_4200,N_653,N_558);
and U4201 (N_4201,N_574,N_1768);
nand U4202 (N_4202,N_1851,N_678);
nand U4203 (N_4203,N_2098,N_1276);
or U4204 (N_4204,N_1614,N_403);
nor U4205 (N_4205,N_1259,N_2190);
nand U4206 (N_4206,N_1645,N_2171);
or U4207 (N_4207,N_2266,N_818);
and U4208 (N_4208,N_1367,N_2126);
nor U4209 (N_4209,N_1523,N_1492);
and U4210 (N_4210,N_969,N_1810);
nor U4211 (N_4211,N_913,N_1416);
nor U4212 (N_4212,N_1562,N_764);
and U4213 (N_4213,N_1268,N_80);
and U4214 (N_4214,N_200,N_1573);
and U4215 (N_4215,N_1157,N_2250);
or U4216 (N_4216,N_2181,N_68);
or U4217 (N_4217,N_1150,N_1359);
and U4218 (N_4218,N_1947,N_2011);
nand U4219 (N_4219,N_2463,N_2205);
xnor U4220 (N_4220,N_429,N_923);
or U4221 (N_4221,N_1042,N_2323);
or U4222 (N_4222,N_217,N_309);
and U4223 (N_4223,N_2058,N_366);
or U4224 (N_4224,N_662,N_1846);
or U4225 (N_4225,N_788,N_1129);
and U4226 (N_4226,N_370,N_182);
nand U4227 (N_4227,N_720,N_664);
nor U4228 (N_4228,N_1493,N_1880);
or U4229 (N_4229,N_1591,N_2457);
or U4230 (N_4230,N_673,N_1484);
nand U4231 (N_4231,N_1250,N_1589);
nor U4232 (N_4232,N_1094,N_2068);
and U4233 (N_4233,N_485,N_1092);
nor U4234 (N_4234,N_1935,N_1580);
nor U4235 (N_4235,N_1938,N_1025);
or U4236 (N_4236,N_2389,N_932);
nor U4237 (N_4237,N_1489,N_542);
or U4238 (N_4238,N_2456,N_2464);
or U4239 (N_4239,N_837,N_1952);
or U4240 (N_4240,N_2252,N_2212);
or U4241 (N_4241,N_2490,N_1818);
nor U4242 (N_4242,N_991,N_1386);
xnor U4243 (N_4243,N_1342,N_948);
nand U4244 (N_4244,N_1410,N_1565);
nor U4245 (N_4245,N_1970,N_2473);
and U4246 (N_4246,N_472,N_2317);
and U4247 (N_4247,N_1123,N_144);
nand U4248 (N_4248,N_1680,N_333);
or U4249 (N_4249,N_496,N_467);
and U4250 (N_4250,N_150,N_1139);
and U4251 (N_4251,N_1847,N_2081);
or U4252 (N_4252,N_1629,N_2274);
nor U4253 (N_4253,N_1797,N_1402);
or U4254 (N_4254,N_2491,N_1330);
nand U4255 (N_4255,N_231,N_1683);
or U4256 (N_4256,N_686,N_354);
nand U4257 (N_4257,N_633,N_1107);
nand U4258 (N_4258,N_1684,N_610);
nand U4259 (N_4259,N_2206,N_1017);
nor U4260 (N_4260,N_547,N_788);
nor U4261 (N_4261,N_1746,N_462);
nor U4262 (N_4262,N_2158,N_2206);
or U4263 (N_4263,N_2270,N_1244);
or U4264 (N_4264,N_454,N_1531);
nand U4265 (N_4265,N_1033,N_1604);
nor U4266 (N_4266,N_980,N_1936);
and U4267 (N_4267,N_1582,N_1774);
nor U4268 (N_4268,N_739,N_794);
and U4269 (N_4269,N_66,N_2116);
nor U4270 (N_4270,N_908,N_1090);
and U4271 (N_4271,N_1816,N_653);
and U4272 (N_4272,N_1788,N_306);
nor U4273 (N_4273,N_1331,N_728);
nand U4274 (N_4274,N_146,N_1762);
nand U4275 (N_4275,N_2424,N_369);
nand U4276 (N_4276,N_1357,N_2235);
nor U4277 (N_4277,N_282,N_2314);
nand U4278 (N_4278,N_1466,N_721);
and U4279 (N_4279,N_2299,N_1823);
xor U4280 (N_4280,N_1717,N_1145);
nand U4281 (N_4281,N_161,N_1915);
and U4282 (N_4282,N_1023,N_3);
nor U4283 (N_4283,N_603,N_493);
nor U4284 (N_4284,N_671,N_298);
nand U4285 (N_4285,N_855,N_1026);
xnor U4286 (N_4286,N_2289,N_371);
nand U4287 (N_4287,N_2023,N_639);
and U4288 (N_4288,N_607,N_32);
and U4289 (N_4289,N_1605,N_1596);
nor U4290 (N_4290,N_402,N_1301);
or U4291 (N_4291,N_1707,N_1458);
nor U4292 (N_4292,N_1571,N_954);
and U4293 (N_4293,N_1969,N_1777);
nor U4294 (N_4294,N_219,N_2020);
nor U4295 (N_4295,N_1553,N_2288);
nand U4296 (N_4296,N_920,N_27);
and U4297 (N_4297,N_2359,N_1633);
nor U4298 (N_4298,N_1130,N_2148);
nand U4299 (N_4299,N_2287,N_65);
nand U4300 (N_4300,N_428,N_704);
or U4301 (N_4301,N_1909,N_1976);
nand U4302 (N_4302,N_2286,N_1612);
and U4303 (N_4303,N_1209,N_812);
nor U4304 (N_4304,N_257,N_2084);
and U4305 (N_4305,N_1537,N_1035);
nor U4306 (N_4306,N_693,N_1719);
and U4307 (N_4307,N_1166,N_1687);
nor U4308 (N_4308,N_2496,N_699);
nor U4309 (N_4309,N_2138,N_2320);
nor U4310 (N_4310,N_2003,N_74);
and U4311 (N_4311,N_1781,N_2028);
nor U4312 (N_4312,N_1978,N_722);
or U4313 (N_4313,N_149,N_1397);
and U4314 (N_4314,N_285,N_1170);
nor U4315 (N_4315,N_2347,N_481);
nand U4316 (N_4316,N_1517,N_112);
nor U4317 (N_4317,N_1799,N_1938);
or U4318 (N_4318,N_2205,N_1324);
nor U4319 (N_4319,N_608,N_1041);
nand U4320 (N_4320,N_1061,N_67);
nor U4321 (N_4321,N_1635,N_94);
and U4322 (N_4322,N_2150,N_1053);
or U4323 (N_4323,N_578,N_1686);
and U4324 (N_4324,N_1457,N_572);
or U4325 (N_4325,N_228,N_82);
and U4326 (N_4326,N_1297,N_378);
and U4327 (N_4327,N_2347,N_2147);
nor U4328 (N_4328,N_2026,N_22);
nor U4329 (N_4329,N_1845,N_945);
xor U4330 (N_4330,N_1437,N_2258);
nor U4331 (N_4331,N_1580,N_2246);
and U4332 (N_4332,N_1814,N_984);
nand U4333 (N_4333,N_1869,N_852);
nor U4334 (N_4334,N_620,N_2120);
or U4335 (N_4335,N_1546,N_1627);
xor U4336 (N_4336,N_1476,N_801);
nand U4337 (N_4337,N_45,N_1268);
nand U4338 (N_4338,N_960,N_2138);
nand U4339 (N_4339,N_44,N_2347);
nand U4340 (N_4340,N_2244,N_1087);
or U4341 (N_4341,N_511,N_781);
or U4342 (N_4342,N_570,N_1944);
nand U4343 (N_4343,N_1160,N_1302);
and U4344 (N_4344,N_863,N_1331);
and U4345 (N_4345,N_358,N_1417);
and U4346 (N_4346,N_1583,N_1561);
nand U4347 (N_4347,N_749,N_728);
and U4348 (N_4348,N_1671,N_1494);
xnor U4349 (N_4349,N_2038,N_1174);
nor U4350 (N_4350,N_224,N_234);
nand U4351 (N_4351,N_1887,N_2468);
nor U4352 (N_4352,N_818,N_1148);
and U4353 (N_4353,N_477,N_158);
or U4354 (N_4354,N_470,N_750);
or U4355 (N_4355,N_1354,N_1952);
or U4356 (N_4356,N_818,N_2239);
and U4357 (N_4357,N_272,N_2372);
nor U4358 (N_4358,N_306,N_1896);
nor U4359 (N_4359,N_357,N_2002);
nor U4360 (N_4360,N_1581,N_2277);
or U4361 (N_4361,N_292,N_1826);
nand U4362 (N_4362,N_2015,N_1116);
nand U4363 (N_4363,N_486,N_1650);
and U4364 (N_4364,N_765,N_1165);
nand U4365 (N_4365,N_715,N_2154);
nand U4366 (N_4366,N_367,N_845);
nand U4367 (N_4367,N_695,N_1214);
or U4368 (N_4368,N_807,N_969);
or U4369 (N_4369,N_2345,N_969);
and U4370 (N_4370,N_2356,N_1084);
and U4371 (N_4371,N_1528,N_929);
and U4372 (N_4372,N_81,N_116);
and U4373 (N_4373,N_1809,N_181);
and U4374 (N_4374,N_2246,N_57);
nor U4375 (N_4375,N_1583,N_200);
nor U4376 (N_4376,N_992,N_230);
and U4377 (N_4377,N_1553,N_2239);
nand U4378 (N_4378,N_192,N_2416);
or U4379 (N_4379,N_1467,N_509);
nand U4380 (N_4380,N_334,N_2381);
nand U4381 (N_4381,N_2315,N_1424);
and U4382 (N_4382,N_2282,N_2299);
or U4383 (N_4383,N_121,N_1374);
nand U4384 (N_4384,N_1730,N_2038);
and U4385 (N_4385,N_1848,N_982);
nor U4386 (N_4386,N_378,N_2353);
and U4387 (N_4387,N_2375,N_2079);
nor U4388 (N_4388,N_860,N_1509);
nand U4389 (N_4389,N_1230,N_769);
and U4390 (N_4390,N_2137,N_2007);
or U4391 (N_4391,N_711,N_259);
and U4392 (N_4392,N_919,N_534);
and U4393 (N_4393,N_2099,N_1926);
nor U4394 (N_4394,N_1651,N_1584);
nor U4395 (N_4395,N_1631,N_1387);
and U4396 (N_4396,N_1107,N_345);
nor U4397 (N_4397,N_2487,N_256);
nand U4398 (N_4398,N_1817,N_134);
and U4399 (N_4399,N_604,N_870);
and U4400 (N_4400,N_1595,N_2085);
nand U4401 (N_4401,N_12,N_1866);
nand U4402 (N_4402,N_2293,N_2294);
nand U4403 (N_4403,N_1988,N_383);
xnor U4404 (N_4404,N_1040,N_2337);
nand U4405 (N_4405,N_1298,N_2271);
or U4406 (N_4406,N_1472,N_837);
or U4407 (N_4407,N_1147,N_2005);
or U4408 (N_4408,N_1885,N_2102);
or U4409 (N_4409,N_1104,N_2214);
nor U4410 (N_4410,N_759,N_1549);
and U4411 (N_4411,N_1365,N_1359);
nor U4412 (N_4412,N_831,N_129);
or U4413 (N_4413,N_1993,N_674);
and U4414 (N_4414,N_1249,N_1494);
and U4415 (N_4415,N_393,N_426);
and U4416 (N_4416,N_727,N_375);
and U4417 (N_4417,N_193,N_2402);
or U4418 (N_4418,N_1301,N_1286);
or U4419 (N_4419,N_1061,N_739);
and U4420 (N_4420,N_549,N_2322);
nor U4421 (N_4421,N_1359,N_874);
nor U4422 (N_4422,N_2318,N_56);
or U4423 (N_4423,N_1737,N_712);
nor U4424 (N_4424,N_1958,N_2040);
and U4425 (N_4425,N_1901,N_2294);
nand U4426 (N_4426,N_1316,N_2293);
nor U4427 (N_4427,N_1335,N_1729);
nor U4428 (N_4428,N_1873,N_1451);
xnor U4429 (N_4429,N_1632,N_734);
nand U4430 (N_4430,N_1222,N_953);
nor U4431 (N_4431,N_808,N_456);
and U4432 (N_4432,N_1311,N_1216);
or U4433 (N_4433,N_2275,N_553);
or U4434 (N_4434,N_2235,N_2266);
nand U4435 (N_4435,N_440,N_1144);
nand U4436 (N_4436,N_1678,N_647);
nor U4437 (N_4437,N_521,N_112);
or U4438 (N_4438,N_428,N_943);
and U4439 (N_4439,N_733,N_1881);
nor U4440 (N_4440,N_1573,N_1660);
and U4441 (N_4441,N_1781,N_96);
nand U4442 (N_4442,N_1459,N_1772);
or U4443 (N_4443,N_2299,N_43);
and U4444 (N_4444,N_2346,N_671);
and U4445 (N_4445,N_674,N_2175);
nand U4446 (N_4446,N_1094,N_683);
nor U4447 (N_4447,N_129,N_1670);
and U4448 (N_4448,N_1486,N_1448);
nor U4449 (N_4449,N_1573,N_290);
xnor U4450 (N_4450,N_1294,N_655);
nor U4451 (N_4451,N_1478,N_2292);
or U4452 (N_4452,N_1292,N_143);
or U4453 (N_4453,N_1253,N_405);
nor U4454 (N_4454,N_343,N_237);
nor U4455 (N_4455,N_2085,N_284);
and U4456 (N_4456,N_2121,N_2034);
nor U4457 (N_4457,N_865,N_553);
and U4458 (N_4458,N_543,N_1948);
or U4459 (N_4459,N_2245,N_1281);
nor U4460 (N_4460,N_335,N_2036);
nor U4461 (N_4461,N_1662,N_1242);
nor U4462 (N_4462,N_1884,N_10);
nor U4463 (N_4463,N_154,N_2491);
nor U4464 (N_4464,N_718,N_1650);
and U4465 (N_4465,N_828,N_1262);
nor U4466 (N_4466,N_1351,N_823);
nand U4467 (N_4467,N_1534,N_776);
nand U4468 (N_4468,N_217,N_1623);
and U4469 (N_4469,N_138,N_1132);
and U4470 (N_4470,N_1320,N_2315);
and U4471 (N_4471,N_481,N_285);
or U4472 (N_4472,N_1395,N_864);
nor U4473 (N_4473,N_114,N_800);
or U4474 (N_4474,N_1083,N_817);
nor U4475 (N_4475,N_295,N_2037);
or U4476 (N_4476,N_519,N_1378);
and U4477 (N_4477,N_2476,N_1009);
and U4478 (N_4478,N_562,N_2263);
or U4479 (N_4479,N_1657,N_2068);
nor U4480 (N_4480,N_1058,N_1280);
and U4481 (N_4481,N_1646,N_1858);
and U4482 (N_4482,N_1061,N_807);
or U4483 (N_4483,N_1352,N_1165);
or U4484 (N_4484,N_1858,N_1859);
nor U4485 (N_4485,N_2241,N_591);
nand U4486 (N_4486,N_1575,N_242);
nand U4487 (N_4487,N_1360,N_2145);
and U4488 (N_4488,N_1720,N_1675);
and U4489 (N_4489,N_1768,N_2493);
nor U4490 (N_4490,N_27,N_1910);
or U4491 (N_4491,N_359,N_2356);
or U4492 (N_4492,N_1386,N_356);
and U4493 (N_4493,N_2379,N_1873);
or U4494 (N_4494,N_1866,N_1305);
nor U4495 (N_4495,N_259,N_1905);
and U4496 (N_4496,N_811,N_175);
and U4497 (N_4497,N_822,N_2196);
nor U4498 (N_4498,N_1477,N_182);
nor U4499 (N_4499,N_1991,N_848);
nand U4500 (N_4500,N_2335,N_1318);
nand U4501 (N_4501,N_894,N_1767);
nor U4502 (N_4502,N_414,N_1614);
or U4503 (N_4503,N_1119,N_1159);
or U4504 (N_4504,N_1324,N_580);
and U4505 (N_4505,N_1362,N_2232);
nand U4506 (N_4506,N_1463,N_444);
and U4507 (N_4507,N_1665,N_2371);
and U4508 (N_4508,N_1265,N_170);
or U4509 (N_4509,N_441,N_1804);
nand U4510 (N_4510,N_1745,N_1832);
nor U4511 (N_4511,N_1409,N_1286);
or U4512 (N_4512,N_1170,N_1508);
nand U4513 (N_4513,N_241,N_476);
and U4514 (N_4514,N_681,N_2370);
nor U4515 (N_4515,N_2232,N_1884);
nand U4516 (N_4516,N_2421,N_349);
or U4517 (N_4517,N_1172,N_1822);
nor U4518 (N_4518,N_2111,N_1901);
and U4519 (N_4519,N_190,N_1270);
nor U4520 (N_4520,N_1526,N_670);
nand U4521 (N_4521,N_2239,N_1399);
and U4522 (N_4522,N_324,N_1233);
nor U4523 (N_4523,N_2098,N_132);
and U4524 (N_4524,N_2483,N_43);
nand U4525 (N_4525,N_804,N_938);
or U4526 (N_4526,N_900,N_1293);
or U4527 (N_4527,N_470,N_1993);
and U4528 (N_4528,N_2341,N_2114);
nor U4529 (N_4529,N_11,N_237);
and U4530 (N_4530,N_866,N_1671);
and U4531 (N_4531,N_449,N_39);
nand U4532 (N_4532,N_929,N_345);
nand U4533 (N_4533,N_1944,N_1144);
nand U4534 (N_4534,N_596,N_368);
nand U4535 (N_4535,N_2076,N_713);
nand U4536 (N_4536,N_2176,N_891);
nor U4537 (N_4537,N_1400,N_2484);
nor U4538 (N_4538,N_687,N_2354);
nand U4539 (N_4539,N_1839,N_2445);
nand U4540 (N_4540,N_1527,N_1193);
and U4541 (N_4541,N_1965,N_2438);
nor U4542 (N_4542,N_2175,N_1291);
nor U4543 (N_4543,N_57,N_52);
nor U4544 (N_4544,N_2321,N_1338);
nand U4545 (N_4545,N_1349,N_2380);
nand U4546 (N_4546,N_2106,N_489);
and U4547 (N_4547,N_467,N_1638);
nor U4548 (N_4548,N_1383,N_2378);
nand U4549 (N_4549,N_444,N_577);
nand U4550 (N_4550,N_592,N_346);
or U4551 (N_4551,N_1086,N_96);
or U4552 (N_4552,N_1868,N_1051);
and U4553 (N_4553,N_1872,N_1208);
and U4554 (N_4554,N_25,N_286);
or U4555 (N_4555,N_827,N_376);
nand U4556 (N_4556,N_2386,N_2090);
nor U4557 (N_4557,N_1807,N_153);
nand U4558 (N_4558,N_74,N_1927);
or U4559 (N_4559,N_1505,N_1037);
or U4560 (N_4560,N_1632,N_67);
nor U4561 (N_4561,N_759,N_33);
nor U4562 (N_4562,N_735,N_55);
or U4563 (N_4563,N_1370,N_151);
or U4564 (N_4564,N_1106,N_160);
and U4565 (N_4565,N_187,N_68);
and U4566 (N_4566,N_419,N_613);
nand U4567 (N_4567,N_136,N_2147);
nand U4568 (N_4568,N_141,N_420);
xor U4569 (N_4569,N_254,N_2180);
nand U4570 (N_4570,N_188,N_2144);
nor U4571 (N_4571,N_653,N_2443);
and U4572 (N_4572,N_1410,N_1515);
nand U4573 (N_4573,N_666,N_627);
nand U4574 (N_4574,N_1177,N_1691);
or U4575 (N_4575,N_1765,N_1398);
nand U4576 (N_4576,N_531,N_1199);
nor U4577 (N_4577,N_865,N_210);
or U4578 (N_4578,N_2068,N_1075);
nand U4579 (N_4579,N_876,N_486);
nor U4580 (N_4580,N_1027,N_990);
and U4581 (N_4581,N_2223,N_675);
and U4582 (N_4582,N_91,N_1629);
nand U4583 (N_4583,N_1264,N_1628);
nor U4584 (N_4584,N_1702,N_305);
or U4585 (N_4585,N_2000,N_467);
nand U4586 (N_4586,N_168,N_762);
and U4587 (N_4587,N_1020,N_503);
or U4588 (N_4588,N_150,N_1807);
and U4589 (N_4589,N_323,N_1828);
nor U4590 (N_4590,N_1782,N_2199);
nand U4591 (N_4591,N_844,N_418);
and U4592 (N_4592,N_2109,N_2385);
nor U4593 (N_4593,N_2335,N_546);
and U4594 (N_4594,N_1189,N_2276);
and U4595 (N_4595,N_1433,N_1712);
or U4596 (N_4596,N_998,N_932);
nor U4597 (N_4597,N_159,N_1734);
nand U4598 (N_4598,N_165,N_18);
nand U4599 (N_4599,N_1744,N_2172);
nor U4600 (N_4600,N_364,N_2076);
nor U4601 (N_4601,N_2367,N_543);
nor U4602 (N_4602,N_448,N_289);
and U4603 (N_4603,N_1695,N_1796);
and U4604 (N_4604,N_2041,N_2266);
nor U4605 (N_4605,N_1586,N_825);
and U4606 (N_4606,N_2491,N_853);
nand U4607 (N_4607,N_220,N_148);
nor U4608 (N_4608,N_1935,N_1203);
nor U4609 (N_4609,N_1328,N_2278);
nor U4610 (N_4610,N_1539,N_1326);
and U4611 (N_4611,N_1016,N_2354);
nand U4612 (N_4612,N_716,N_935);
or U4613 (N_4613,N_1775,N_62);
and U4614 (N_4614,N_948,N_2303);
nor U4615 (N_4615,N_871,N_929);
nand U4616 (N_4616,N_2223,N_2109);
nand U4617 (N_4617,N_1877,N_950);
xor U4618 (N_4618,N_2183,N_2113);
or U4619 (N_4619,N_252,N_140);
nor U4620 (N_4620,N_1442,N_1217);
nor U4621 (N_4621,N_50,N_2028);
and U4622 (N_4622,N_1929,N_1222);
or U4623 (N_4623,N_445,N_2005);
nand U4624 (N_4624,N_1842,N_708);
and U4625 (N_4625,N_23,N_2468);
nand U4626 (N_4626,N_1625,N_520);
nand U4627 (N_4627,N_967,N_124);
nand U4628 (N_4628,N_1027,N_1874);
and U4629 (N_4629,N_1813,N_1603);
or U4630 (N_4630,N_637,N_1513);
nand U4631 (N_4631,N_1860,N_864);
nor U4632 (N_4632,N_2385,N_357);
nand U4633 (N_4633,N_296,N_1795);
and U4634 (N_4634,N_1491,N_1239);
and U4635 (N_4635,N_319,N_2190);
and U4636 (N_4636,N_49,N_1218);
nand U4637 (N_4637,N_746,N_310);
nor U4638 (N_4638,N_254,N_870);
nor U4639 (N_4639,N_1239,N_2461);
or U4640 (N_4640,N_696,N_472);
and U4641 (N_4641,N_1249,N_1691);
or U4642 (N_4642,N_2103,N_1286);
nand U4643 (N_4643,N_2272,N_2017);
or U4644 (N_4644,N_1886,N_1460);
nor U4645 (N_4645,N_664,N_223);
or U4646 (N_4646,N_28,N_144);
xnor U4647 (N_4647,N_795,N_2436);
nor U4648 (N_4648,N_645,N_1262);
nand U4649 (N_4649,N_2024,N_1882);
nand U4650 (N_4650,N_991,N_1380);
nor U4651 (N_4651,N_191,N_99);
nand U4652 (N_4652,N_736,N_1098);
xor U4653 (N_4653,N_688,N_78);
and U4654 (N_4654,N_55,N_1085);
nand U4655 (N_4655,N_2487,N_1565);
nor U4656 (N_4656,N_1119,N_498);
or U4657 (N_4657,N_477,N_1993);
nand U4658 (N_4658,N_1186,N_2380);
and U4659 (N_4659,N_23,N_781);
nor U4660 (N_4660,N_2176,N_1824);
and U4661 (N_4661,N_1216,N_2266);
and U4662 (N_4662,N_914,N_2097);
and U4663 (N_4663,N_803,N_374);
nand U4664 (N_4664,N_1335,N_1451);
nand U4665 (N_4665,N_458,N_1910);
nand U4666 (N_4666,N_2017,N_513);
nor U4667 (N_4667,N_1345,N_1924);
nor U4668 (N_4668,N_307,N_1987);
and U4669 (N_4669,N_310,N_1781);
nor U4670 (N_4670,N_1291,N_1479);
nor U4671 (N_4671,N_600,N_1215);
nand U4672 (N_4672,N_666,N_1039);
and U4673 (N_4673,N_950,N_1612);
and U4674 (N_4674,N_2436,N_1273);
nor U4675 (N_4675,N_1818,N_928);
or U4676 (N_4676,N_2097,N_2175);
or U4677 (N_4677,N_31,N_1760);
or U4678 (N_4678,N_1922,N_634);
nand U4679 (N_4679,N_979,N_1967);
and U4680 (N_4680,N_2325,N_212);
nor U4681 (N_4681,N_2074,N_1673);
and U4682 (N_4682,N_786,N_1104);
and U4683 (N_4683,N_1824,N_564);
and U4684 (N_4684,N_955,N_2006);
nor U4685 (N_4685,N_794,N_167);
or U4686 (N_4686,N_1286,N_805);
or U4687 (N_4687,N_1460,N_1706);
and U4688 (N_4688,N_212,N_2093);
nor U4689 (N_4689,N_124,N_290);
or U4690 (N_4690,N_591,N_1429);
or U4691 (N_4691,N_371,N_2089);
nand U4692 (N_4692,N_1327,N_1682);
or U4693 (N_4693,N_1103,N_1551);
and U4694 (N_4694,N_936,N_1485);
nand U4695 (N_4695,N_1741,N_305);
nor U4696 (N_4696,N_536,N_1312);
and U4697 (N_4697,N_1900,N_2270);
nor U4698 (N_4698,N_2267,N_394);
and U4699 (N_4699,N_271,N_290);
and U4700 (N_4700,N_1721,N_1722);
and U4701 (N_4701,N_1169,N_2156);
nand U4702 (N_4702,N_1973,N_92);
and U4703 (N_4703,N_785,N_320);
nand U4704 (N_4704,N_1187,N_2166);
or U4705 (N_4705,N_2404,N_1811);
nor U4706 (N_4706,N_120,N_1469);
nand U4707 (N_4707,N_2452,N_1789);
nor U4708 (N_4708,N_1969,N_1241);
and U4709 (N_4709,N_1953,N_1941);
or U4710 (N_4710,N_2268,N_2253);
nor U4711 (N_4711,N_1201,N_1074);
or U4712 (N_4712,N_1355,N_830);
nand U4713 (N_4713,N_249,N_428);
nor U4714 (N_4714,N_260,N_387);
and U4715 (N_4715,N_1619,N_931);
nor U4716 (N_4716,N_533,N_844);
nor U4717 (N_4717,N_384,N_1572);
nand U4718 (N_4718,N_2269,N_2078);
nand U4719 (N_4719,N_211,N_2231);
nor U4720 (N_4720,N_1180,N_192);
nand U4721 (N_4721,N_1036,N_2409);
nor U4722 (N_4722,N_797,N_1484);
and U4723 (N_4723,N_1254,N_1484);
nor U4724 (N_4724,N_870,N_2110);
nand U4725 (N_4725,N_2332,N_1396);
nor U4726 (N_4726,N_399,N_245);
and U4727 (N_4727,N_1206,N_313);
nor U4728 (N_4728,N_1196,N_1580);
or U4729 (N_4729,N_2403,N_2426);
nand U4730 (N_4730,N_1262,N_1434);
nand U4731 (N_4731,N_1100,N_407);
and U4732 (N_4732,N_969,N_1658);
nand U4733 (N_4733,N_1942,N_2078);
or U4734 (N_4734,N_14,N_1721);
nand U4735 (N_4735,N_1360,N_781);
or U4736 (N_4736,N_1115,N_600);
or U4737 (N_4737,N_691,N_2213);
or U4738 (N_4738,N_931,N_1318);
or U4739 (N_4739,N_403,N_990);
or U4740 (N_4740,N_1635,N_2176);
nor U4741 (N_4741,N_1324,N_873);
nor U4742 (N_4742,N_181,N_208);
nor U4743 (N_4743,N_529,N_2127);
nor U4744 (N_4744,N_1437,N_825);
nand U4745 (N_4745,N_1506,N_1856);
nor U4746 (N_4746,N_1113,N_689);
and U4747 (N_4747,N_591,N_1522);
nor U4748 (N_4748,N_732,N_2192);
or U4749 (N_4749,N_1572,N_1742);
or U4750 (N_4750,N_542,N_1356);
or U4751 (N_4751,N_1991,N_846);
and U4752 (N_4752,N_2377,N_1238);
or U4753 (N_4753,N_783,N_1824);
or U4754 (N_4754,N_1510,N_1289);
and U4755 (N_4755,N_317,N_214);
or U4756 (N_4756,N_220,N_1821);
nor U4757 (N_4757,N_389,N_247);
nand U4758 (N_4758,N_1456,N_2243);
nor U4759 (N_4759,N_104,N_1681);
or U4760 (N_4760,N_1356,N_1773);
and U4761 (N_4761,N_2092,N_680);
and U4762 (N_4762,N_162,N_1721);
and U4763 (N_4763,N_1876,N_2481);
nor U4764 (N_4764,N_379,N_1415);
and U4765 (N_4765,N_1168,N_17);
or U4766 (N_4766,N_1615,N_1087);
and U4767 (N_4767,N_617,N_869);
xnor U4768 (N_4768,N_177,N_1773);
and U4769 (N_4769,N_1047,N_793);
and U4770 (N_4770,N_401,N_415);
nand U4771 (N_4771,N_917,N_1012);
or U4772 (N_4772,N_2455,N_863);
or U4773 (N_4773,N_1862,N_1153);
and U4774 (N_4774,N_232,N_2440);
nor U4775 (N_4775,N_1214,N_133);
nand U4776 (N_4776,N_176,N_2364);
nand U4777 (N_4777,N_324,N_98);
and U4778 (N_4778,N_924,N_1653);
nor U4779 (N_4779,N_1521,N_1015);
and U4780 (N_4780,N_384,N_114);
or U4781 (N_4781,N_1213,N_502);
nor U4782 (N_4782,N_495,N_2087);
or U4783 (N_4783,N_1307,N_1026);
nor U4784 (N_4784,N_2293,N_308);
nand U4785 (N_4785,N_941,N_423);
and U4786 (N_4786,N_188,N_1572);
or U4787 (N_4787,N_397,N_1185);
or U4788 (N_4788,N_1118,N_1061);
or U4789 (N_4789,N_825,N_538);
and U4790 (N_4790,N_1345,N_1294);
nand U4791 (N_4791,N_2156,N_101);
and U4792 (N_4792,N_2442,N_799);
or U4793 (N_4793,N_1820,N_1483);
and U4794 (N_4794,N_102,N_1707);
nand U4795 (N_4795,N_1419,N_953);
nor U4796 (N_4796,N_999,N_2096);
xnor U4797 (N_4797,N_1543,N_263);
nand U4798 (N_4798,N_1694,N_204);
nor U4799 (N_4799,N_2269,N_478);
or U4800 (N_4800,N_34,N_2454);
nor U4801 (N_4801,N_2200,N_2383);
nor U4802 (N_4802,N_1606,N_2015);
nand U4803 (N_4803,N_328,N_1520);
and U4804 (N_4804,N_1328,N_1031);
and U4805 (N_4805,N_2271,N_65);
and U4806 (N_4806,N_1781,N_1153);
and U4807 (N_4807,N_1048,N_121);
nand U4808 (N_4808,N_2264,N_36);
nor U4809 (N_4809,N_2209,N_800);
nor U4810 (N_4810,N_773,N_1596);
nand U4811 (N_4811,N_1848,N_1999);
and U4812 (N_4812,N_2051,N_500);
or U4813 (N_4813,N_2161,N_1450);
or U4814 (N_4814,N_634,N_154);
nor U4815 (N_4815,N_2384,N_1224);
or U4816 (N_4816,N_1494,N_2482);
nor U4817 (N_4817,N_920,N_2083);
and U4818 (N_4818,N_1281,N_1973);
nand U4819 (N_4819,N_47,N_1413);
and U4820 (N_4820,N_1277,N_2208);
xor U4821 (N_4821,N_887,N_1605);
nand U4822 (N_4822,N_2363,N_1915);
nand U4823 (N_4823,N_1320,N_1309);
and U4824 (N_4824,N_2033,N_1047);
and U4825 (N_4825,N_1070,N_1127);
nand U4826 (N_4826,N_2261,N_1496);
or U4827 (N_4827,N_1003,N_520);
and U4828 (N_4828,N_2473,N_1612);
or U4829 (N_4829,N_169,N_2231);
nand U4830 (N_4830,N_1481,N_414);
nand U4831 (N_4831,N_1881,N_638);
nand U4832 (N_4832,N_263,N_26);
and U4833 (N_4833,N_1421,N_2312);
nand U4834 (N_4834,N_29,N_1414);
nor U4835 (N_4835,N_1612,N_290);
nor U4836 (N_4836,N_960,N_322);
nand U4837 (N_4837,N_339,N_1416);
nand U4838 (N_4838,N_2420,N_630);
nor U4839 (N_4839,N_694,N_2396);
and U4840 (N_4840,N_277,N_576);
or U4841 (N_4841,N_1583,N_312);
and U4842 (N_4842,N_1838,N_1180);
nand U4843 (N_4843,N_596,N_2062);
or U4844 (N_4844,N_1972,N_576);
nor U4845 (N_4845,N_116,N_723);
or U4846 (N_4846,N_848,N_1921);
nor U4847 (N_4847,N_2181,N_1864);
nand U4848 (N_4848,N_1671,N_350);
and U4849 (N_4849,N_1353,N_271);
nand U4850 (N_4850,N_566,N_2233);
or U4851 (N_4851,N_2214,N_477);
nor U4852 (N_4852,N_1036,N_424);
and U4853 (N_4853,N_1068,N_2271);
nand U4854 (N_4854,N_499,N_2434);
nand U4855 (N_4855,N_1782,N_496);
nand U4856 (N_4856,N_1317,N_760);
nand U4857 (N_4857,N_1604,N_1288);
and U4858 (N_4858,N_1121,N_261);
nor U4859 (N_4859,N_143,N_472);
and U4860 (N_4860,N_240,N_1579);
or U4861 (N_4861,N_1520,N_1176);
xnor U4862 (N_4862,N_1012,N_605);
nor U4863 (N_4863,N_299,N_2402);
nor U4864 (N_4864,N_247,N_349);
nor U4865 (N_4865,N_667,N_915);
or U4866 (N_4866,N_65,N_418);
and U4867 (N_4867,N_2066,N_1652);
nand U4868 (N_4868,N_619,N_644);
nor U4869 (N_4869,N_1420,N_659);
or U4870 (N_4870,N_871,N_2162);
or U4871 (N_4871,N_30,N_847);
or U4872 (N_4872,N_2134,N_2174);
xnor U4873 (N_4873,N_1220,N_893);
or U4874 (N_4874,N_2079,N_1805);
nand U4875 (N_4875,N_2423,N_511);
or U4876 (N_4876,N_1743,N_1004);
or U4877 (N_4877,N_2460,N_148);
nor U4878 (N_4878,N_2221,N_689);
nand U4879 (N_4879,N_1993,N_1252);
and U4880 (N_4880,N_612,N_1583);
or U4881 (N_4881,N_41,N_73);
and U4882 (N_4882,N_1549,N_2144);
or U4883 (N_4883,N_2254,N_1443);
nor U4884 (N_4884,N_573,N_218);
nor U4885 (N_4885,N_1489,N_871);
and U4886 (N_4886,N_1536,N_1289);
or U4887 (N_4887,N_560,N_1383);
and U4888 (N_4888,N_1580,N_926);
nor U4889 (N_4889,N_575,N_1005);
or U4890 (N_4890,N_1763,N_1250);
or U4891 (N_4891,N_2094,N_2477);
and U4892 (N_4892,N_559,N_2224);
nor U4893 (N_4893,N_1415,N_1784);
and U4894 (N_4894,N_1758,N_0);
nor U4895 (N_4895,N_908,N_2024);
and U4896 (N_4896,N_1418,N_1856);
or U4897 (N_4897,N_635,N_2456);
nand U4898 (N_4898,N_1243,N_148);
or U4899 (N_4899,N_632,N_1944);
or U4900 (N_4900,N_2114,N_1283);
nand U4901 (N_4901,N_932,N_2340);
and U4902 (N_4902,N_1494,N_580);
nand U4903 (N_4903,N_1101,N_2207);
nand U4904 (N_4904,N_1441,N_26);
or U4905 (N_4905,N_18,N_387);
or U4906 (N_4906,N_231,N_1093);
nor U4907 (N_4907,N_1428,N_2224);
or U4908 (N_4908,N_297,N_528);
or U4909 (N_4909,N_2258,N_934);
or U4910 (N_4910,N_2173,N_1639);
nand U4911 (N_4911,N_1770,N_991);
or U4912 (N_4912,N_1155,N_1661);
nand U4913 (N_4913,N_2066,N_2355);
nor U4914 (N_4914,N_419,N_1602);
nand U4915 (N_4915,N_862,N_2104);
or U4916 (N_4916,N_1269,N_1599);
or U4917 (N_4917,N_306,N_2144);
nand U4918 (N_4918,N_1036,N_1277);
or U4919 (N_4919,N_1781,N_839);
nand U4920 (N_4920,N_1313,N_366);
nor U4921 (N_4921,N_2492,N_2148);
nor U4922 (N_4922,N_1401,N_2444);
nand U4923 (N_4923,N_2336,N_710);
and U4924 (N_4924,N_2029,N_1091);
or U4925 (N_4925,N_1563,N_1424);
nand U4926 (N_4926,N_644,N_829);
and U4927 (N_4927,N_1929,N_1368);
or U4928 (N_4928,N_2181,N_2064);
nand U4929 (N_4929,N_355,N_1621);
or U4930 (N_4930,N_1924,N_1900);
nand U4931 (N_4931,N_1264,N_251);
and U4932 (N_4932,N_1916,N_844);
nor U4933 (N_4933,N_1348,N_799);
nand U4934 (N_4934,N_1503,N_1061);
and U4935 (N_4935,N_97,N_209);
nor U4936 (N_4936,N_2078,N_2140);
nor U4937 (N_4937,N_1189,N_1296);
nand U4938 (N_4938,N_20,N_2427);
or U4939 (N_4939,N_950,N_133);
nor U4940 (N_4940,N_2373,N_256);
and U4941 (N_4941,N_1850,N_397);
or U4942 (N_4942,N_715,N_1862);
nand U4943 (N_4943,N_1174,N_15);
or U4944 (N_4944,N_2210,N_1825);
and U4945 (N_4945,N_297,N_2032);
or U4946 (N_4946,N_2086,N_2026);
nand U4947 (N_4947,N_1603,N_1737);
nor U4948 (N_4948,N_1141,N_499);
nor U4949 (N_4949,N_41,N_935);
nand U4950 (N_4950,N_1122,N_263);
nand U4951 (N_4951,N_2064,N_714);
nand U4952 (N_4952,N_917,N_448);
and U4953 (N_4953,N_1246,N_2091);
nor U4954 (N_4954,N_543,N_729);
or U4955 (N_4955,N_414,N_2123);
or U4956 (N_4956,N_830,N_803);
or U4957 (N_4957,N_2367,N_2202);
nand U4958 (N_4958,N_1246,N_2084);
nand U4959 (N_4959,N_1023,N_1393);
nand U4960 (N_4960,N_2198,N_216);
xor U4961 (N_4961,N_1020,N_319);
or U4962 (N_4962,N_2302,N_939);
nand U4963 (N_4963,N_573,N_114);
and U4964 (N_4964,N_737,N_966);
or U4965 (N_4965,N_1124,N_705);
nand U4966 (N_4966,N_1208,N_396);
or U4967 (N_4967,N_2191,N_2303);
nand U4968 (N_4968,N_1622,N_1261);
nor U4969 (N_4969,N_482,N_918);
nor U4970 (N_4970,N_1119,N_2260);
and U4971 (N_4971,N_1642,N_818);
nor U4972 (N_4972,N_761,N_1771);
and U4973 (N_4973,N_1214,N_1159);
or U4974 (N_4974,N_2436,N_2406);
nand U4975 (N_4975,N_823,N_931);
nor U4976 (N_4976,N_1343,N_1741);
nand U4977 (N_4977,N_2317,N_660);
and U4978 (N_4978,N_2209,N_939);
nor U4979 (N_4979,N_2106,N_1452);
or U4980 (N_4980,N_67,N_1381);
or U4981 (N_4981,N_870,N_415);
nor U4982 (N_4982,N_638,N_976);
nor U4983 (N_4983,N_266,N_1814);
and U4984 (N_4984,N_78,N_1044);
nand U4985 (N_4985,N_1777,N_2006);
or U4986 (N_4986,N_1656,N_1712);
or U4987 (N_4987,N_2326,N_1874);
and U4988 (N_4988,N_2156,N_708);
or U4989 (N_4989,N_1018,N_1379);
nor U4990 (N_4990,N_605,N_1502);
or U4991 (N_4991,N_777,N_1551);
and U4992 (N_4992,N_2249,N_354);
and U4993 (N_4993,N_1831,N_68);
or U4994 (N_4994,N_2063,N_2498);
nor U4995 (N_4995,N_978,N_710);
and U4996 (N_4996,N_1203,N_1318);
and U4997 (N_4997,N_1696,N_1744);
xor U4998 (N_4998,N_1911,N_1015);
and U4999 (N_4999,N_1436,N_1444);
nor U5000 (N_5000,N_4495,N_4494);
or U5001 (N_5001,N_3307,N_4938);
and U5002 (N_5002,N_4208,N_4270);
or U5003 (N_5003,N_4618,N_3083);
nand U5004 (N_5004,N_3508,N_3536);
xnor U5005 (N_5005,N_3708,N_4247);
nand U5006 (N_5006,N_3197,N_3850);
or U5007 (N_5007,N_4934,N_3893);
and U5008 (N_5008,N_4070,N_4811);
or U5009 (N_5009,N_4133,N_3745);
or U5010 (N_5010,N_3973,N_4988);
nand U5011 (N_5011,N_2657,N_4281);
or U5012 (N_5012,N_4765,N_2810);
and U5013 (N_5013,N_4752,N_2641);
or U5014 (N_5014,N_4172,N_4457);
and U5015 (N_5015,N_2608,N_4604);
nor U5016 (N_5016,N_4864,N_3749);
nor U5017 (N_5017,N_4061,N_4499);
nand U5018 (N_5018,N_4942,N_3626);
nand U5019 (N_5019,N_3776,N_4388);
or U5020 (N_5020,N_3930,N_4092);
nand U5021 (N_5021,N_2639,N_4478);
or U5022 (N_5022,N_3814,N_4330);
or U5023 (N_5023,N_3562,N_4547);
and U5024 (N_5024,N_4939,N_2527);
nor U5025 (N_5025,N_4305,N_3060);
xnor U5026 (N_5026,N_2865,N_4375);
or U5027 (N_5027,N_2552,N_3951);
and U5028 (N_5028,N_3681,N_3057);
and U5029 (N_5029,N_2854,N_4719);
nand U5030 (N_5030,N_2522,N_3333);
nand U5031 (N_5031,N_3996,N_4687);
nor U5032 (N_5032,N_2794,N_4932);
or U5033 (N_5033,N_4455,N_4782);
nand U5034 (N_5034,N_2572,N_3637);
nand U5035 (N_5035,N_3670,N_4698);
nor U5036 (N_5036,N_3542,N_2895);
and U5037 (N_5037,N_2846,N_2856);
or U5038 (N_5038,N_3963,N_3938);
or U5039 (N_5039,N_2908,N_2693);
and U5040 (N_5040,N_3134,N_3486);
or U5041 (N_5041,N_3774,N_4084);
nor U5042 (N_5042,N_4037,N_3877);
and U5043 (N_5043,N_2947,N_3650);
and U5044 (N_5044,N_4737,N_4404);
nand U5045 (N_5045,N_2610,N_4717);
nand U5046 (N_5046,N_4417,N_3808);
and U5047 (N_5047,N_3202,N_4574);
or U5048 (N_5048,N_4053,N_4371);
or U5049 (N_5049,N_4958,N_3099);
and U5050 (N_5050,N_4738,N_2537);
or U5051 (N_5051,N_2560,N_2642);
and U5052 (N_5052,N_3147,N_3062);
nand U5053 (N_5053,N_3361,N_3857);
nand U5054 (N_5054,N_4729,N_3932);
and U5055 (N_5055,N_2937,N_4658);
nand U5056 (N_5056,N_4855,N_3087);
nor U5057 (N_5057,N_4215,N_3530);
and U5058 (N_5058,N_2832,N_3610);
or U5059 (N_5059,N_3009,N_4905);
nand U5060 (N_5060,N_4653,N_2899);
nand U5061 (N_5061,N_2807,N_2729);
or U5062 (N_5062,N_4400,N_3594);
and U5063 (N_5063,N_2583,N_4397);
nand U5064 (N_5064,N_4901,N_3621);
and U5065 (N_5065,N_4413,N_3402);
and U5066 (N_5066,N_4832,N_3565);
nor U5067 (N_5067,N_4586,N_3622);
or U5068 (N_5068,N_2573,N_4209);
nand U5069 (N_5069,N_2600,N_4394);
nor U5070 (N_5070,N_3515,N_3678);
and U5071 (N_5071,N_3546,N_4088);
nand U5072 (N_5072,N_2556,N_4861);
or U5073 (N_5073,N_4761,N_2933);
nor U5074 (N_5074,N_3751,N_4881);
and U5075 (N_5075,N_4333,N_3509);
or U5076 (N_5076,N_3547,N_3107);
or U5077 (N_5077,N_3810,N_3500);
nor U5078 (N_5078,N_3700,N_3685);
or U5079 (N_5079,N_4667,N_4205);
or U5080 (N_5080,N_4476,N_4140);
and U5081 (N_5081,N_3686,N_3200);
and U5082 (N_5082,N_3394,N_4530);
nor U5083 (N_5083,N_2944,N_3868);
or U5084 (N_5084,N_3525,N_4122);
or U5085 (N_5085,N_4844,N_3431);
or U5086 (N_5086,N_2667,N_2523);
and U5087 (N_5087,N_3615,N_4091);
or U5088 (N_5088,N_3955,N_3252);
nor U5089 (N_5089,N_3108,N_2844);
and U5090 (N_5090,N_4664,N_3886);
nor U5091 (N_5091,N_3958,N_3653);
and U5092 (N_5092,N_3150,N_2890);
nor U5093 (N_5093,N_4021,N_3370);
and U5094 (N_5094,N_4633,N_2765);
nor U5095 (N_5095,N_2542,N_4927);
and U5096 (N_5096,N_3258,N_4976);
nor U5097 (N_5097,N_4789,N_3033);
nor U5098 (N_5098,N_3855,N_4242);
nor U5099 (N_5099,N_4280,N_4343);
nand U5100 (N_5100,N_2670,N_4526);
nor U5101 (N_5101,N_3701,N_3986);
nor U5102 (N_5102,N_4080,N_4451);
nor U5103 (N_5103,N_4012,N_2823);
nor U5104 (N_5104,N_3226,N_3605);
nor U5105 (N_5105,N_4358,N_3702);
xor U5106 (N_5106,N_2697,N_4943);
and U5107 (N_5107,N_3350,N_4297);
nor U5108 (N_5108,N_4331,N_2849);
and U5109 (N_5109,N_3987,N_2809);
nor U5110 (N_5110,N_4899,N_3948);
nor U5111 (N_5111,N_3335,N_4403);
nand U5112 (N_5112,N_2688,N_3941);
or U5113 (N_5113,N_4121,N_4860);
nand U5114 (N_5114,N_2742,N_2645);
or U5115 (N_5115,N_2804,N_4059);
and U5116 (N_5116,N_4800,N_4273);
nand U5117 (N_5117,N_4060,N_2718);
or U5118 (N_5118,N_3095,N_4655);
nand U5119 (N_5119,N_3505,N_3295);
nand U5120 (N_5120,N_3121,N_4481);
nor U5121 (N_5121,N_4046,N_4148);
or U5122 (N_5122,N_2633,N_4833);
nand U5123 (N_5123,N_4598,N_2623);
nand U5124 (N_5124,N_2748,N_3916);
nand U5125 (N_5125,N_3204,N_4852);
and U5126 (N_5126,N_2978,N_4533);
or U5127 (N_5127,N_2516,N_2601);
nor U5128 (N_5128,N_3102,N_3097);
or U5129 (N_5129,N_4848,N_2784);
or U5130 (N_5130,N_3053,N_3597);
and U5131 (N_5131,N_4056,N_4113);
nand U5132 (N_5132,N_3796,N_3429);
nand U5133 (N_5133,N_4029,N_2827);
nor U5134 (N_5134,N_3929,N_3110);
nand U5135 (N_5135,N_2781,N_4415);
or U5136 (N_5136,N_4773,N_3477);
nor U5137 (N_5137,N_4685,N_4111);
and U5138 (N_5138,N_3544,N_3193);
nand U5139 (N_5139,N_2607,N_3199);
nor U5140 (N_5140,N_3704,N_4985);
nand U5141 (N_5141,N_4585,N_3391);
and U5142 (N_5142,N_3705,N_2932);
nor U5143 (N_5143,N_3762,N_3408);
nor U5144 (N_5144,N_4469,N_4026);
nand U5145 (N_5145,N_2584,N_4191);
or U5146 (N_5146,N_3464,N_4069);
nand U5147 (N_5147,N_3367,N_3981);
nand U5148 (N_5148,N_2617,N_2689);
nand U5149 (N_5149,N_3235,N_4880);
nor U5150 (N_5150,N_3209,N_3261);
nand U5151 (N_5151,N_3876,N_2538);
nand U5152 (N_5152,N_3922,N_2761);
or U5153 (N_5153,N_3791,N_2826);
and U5154 (N_5154,N_2997,N_3523);
nand U5155 (N_5155,N_4704,N_4039);
nor U5156 (N_5156,N_4776,N_3711);
nor U5157 (N_5157,N_2758,N_2732);
or U5158 (N_5158,N_4551,N_4941);
nor U5159 (N_5159,N_3553,N_2529);
and U5160 (N_5160,N_4108,N_4110);
nor U5161 (N_5161,N_3510,N_4434);
nand U5162 (N_5162,N_3139,N_4758);
xor U5163 (N_5163,N_2636,N_4344);
nor U5164 (N_5164,N_3441,N_3342);
nor U5165 (N_5165,N_2963,N_3723);
and U5166 (N_5166,N_3819,N_4202);
nand U5167 (N_5167,N_3504,N_2614);
nor U5168 (N_5168,N_2582,N_2549);
nand U5169 (N_5169,N_2707,N_2575);
nor U5170 (N_5170,N_2665,N_2676);
nand U5171 (N_5171,N_2650,N_2915);
nand U5172 (N_5172,N_4853,N_4194);
nor U5173 (N_5173,N_3625,N_4185);
nor U5174 (N_5174,N_2692,N_3640);
or U5175 (N_5175,N_4360,N_2816);
nor U5176 (N_5176,N_4563,N_4335);
nand U5177 (N_5177,N_2727,N_4078);
nand U5178 (N_5178,N_4623,N_3502);
nor U5179 (N_5179,N_3690,N_4957);
nor U5180 (N_5180,N_4326,N_3444);
or U5181 (N_5181,N_2672,N_2593);
nor U5182 (N_5182,N_4570,N_4702);
nand U5183 (N_5183,N_3919,N_3560);
and U5184 (N_5184,N_4724,N_4525);
nand U5185 (N_5185,N_4695,N_3215);
nor U5186 (N_5186,N_4614,N_4238);
nand U5187 (N_5187,N_2730,N_3806);
and U5188 (N_5188,N_3914,N_4236);
nor U5189 (N_5189,N_3218,N_2561);
and U5190 (N_5190,N_3960,N_3338);
and U5191 (N_5191,N_4176,N_4747);
nor U5192 (N_5192,N_3365,N_4278);
nor U5193 (N_5193,N_2803,N_3142);
or U5194 (N_5194,N_4458,N_3660);
nand U5195 (N_5195,N_4341,N_3943);
or U5196 (N_5196,N_3341,N_2666);
nor U5197 (N_5197,N_3779,N_3082);
nor U5198 (N_5198,N_4302,N_4418);
and U5199 (N_5199,N_4014,N_3664);
nor U5200 (N_5200,N_4592,N_3761);
or U5201 (N_5201,N_4402,N_3128);
nor U5202 (N_5202,N_3122,N_3120);
nand U5203 (N_5203,N_3381,N_3976);
or U5204 (N_5204,N_3752,N_2864);
or U5205 (N_5205,N_2753,N_4309);
and U5206 (N_5206,N_4240,N_2514);
nor U5207 (N_5207,N_3130,N_4625);
and U5208 (N_5208,N_4025,N_4186);
and U5209 (N_5209,N_4733,N_3773);
or U5210 (N_5210,N_4541,N_3856);
or U5211 (N_5211,N_4249,N_3399);
nand U5212 (N_5212,N_4783,N_4619);
or U5213 (N_5213,N_4293,N_4267);
or U5214 (N_5214,N_4696,N_3063);
nor U5215 (N_5215,N_4116,N_3915);
nand U5216 (N_5216,N_2926,N_3470);
nand U5217 (N_5217,N_2589,N_3067);
nand U5218 (N_5218,N_4079,N_4534);
or U5219 (N_5219,N_4157,N_3116);
or U5220 (N_5220,N_3173,N_4561);
xor U5221 (N_5221,N_3568,N_4809);
or U5222 (N_5222,N_3931,N_2935);
nand U5223 (N_5223,N_4726,N_4143);
and U5224 (N_5224,N_2694,N_3729);
nor U5225 (N_5225,N_4223,N_2562);
or U5226 (N_5226,N_4031,N_3840);
or U5227 (N_5227,N_4363,N_4874);
or U5228 (N_5228,N_2988,N_4973);
nand U5229 (N_5229,N_3927,N_4154);
nor U5230 (N_5230,N_2924,N_4916);
or U5231 (N_5231,N_4003,N_2546);
nand U5232 (N_5232,N_3165,N_3074);
nand U5233 (N_5233,N_2540,N_2961);
and U5234 (N_5234,N_2681,N_4219);
or U5235 (N_5235,N_4032,N_2559);
nand U5236 (N_5236,N_3160,N_4791);
and U5237 (N_5237,N_4107,N_3482);
nor U5238 (N_5238,N_3599,N_3171);
nor U5239 (N_5239,N_4828,N_3356);
nand U5240 (N_5240,N_3574,N_2837);
nor U5241 (N_5241,N_4347,N_3100);
nand U5242 (N_5242,N_3999,N_3225);
nand U5243 (N_5243,N_2504,N_3946);
nor U5244 (N_5244,N_3240,N_3835);
or U5245 (N_5245,N_4180,N_4395);
or U5246 (N_5246,N_3519,N_4544);
nor U5247 (N_5247,N_2543,N_4411);
nor U5248 (N_5248,N_3006,N_4638);
or U5249 (N_5249,N_2717,N_3680);
nor U5250 (N_5250,N_2945,N_2515);
and U5251 (N_5251,N_2792,N_3939);
xnor U5252 (N_5252,N_4306,N_2889);
and U5253 (N_5253,N_2622,N_2796);
or U5254 (N_5254,N_4230,N_4595);
nand U5255 (N_5255,N_3124,N_3149);
nor U5256 (N_5256,N_4668,N_3741);
nor U5257 (N_5257,N_3188,N_4264);
and U5258 (N_5258,N_3957,N_2946);
nor U5259 (N_5259,N_3011,N_3414);
nand U5260 (N_5260,N_2592,N_4956);
nor U5261 (N_5261,N_2825,N_4073);
or U5262 (N_5262,N_4651,N_3129);
nor U5263 (N_5263,N_4991,N_4231);
or U5264 (N_5264,N_2913,N_4989);
and U5265 (N_5265,N_3086,N_2747);
and U5266 (N_5266,N_2801,N_3382);
and U5267 (N_5267,N_4010,N_3459);
nand U5268 (N_5268,N_4671,N_4682);
nor U5269 (N_5269,N_3112,N_4642);
or U5270 (N_5270,N_2594,N_4296);
or U5271 (N_5271,N_4516,N_2891);
nand U5272 (N_5272,N_3529,N_2595);
and U5273 (N_5273,N_2776,N_3205);
nand U5274 (N_5274,N_4020,N_4362);
or U5275 (N_5275,N_4596,N_4322);
nor U5276 (N_5276,N_3816,N_4139);
or U5277 (N_5277,N_4398,N_3353);
nor U5278 (N_5278,N_4117,N_3019);
or U5279 (N_5279,N_2661,N_4568);
nor U5280 (N_5280,N_4894,N_3201);
and U5281 (N_5281,N_4022,N_4156);
or U5282 (N_5282,N_3123,N_2558);
nor U5283 (N_5283,N_2914,N_4166);
nand U5284 (N_5284,N_3588,N_3170);
and U5285 (N_5285,N_4774,N_3954);
nand U5286 (N_5286,N_2513,N_4199);
nand U5287 (N_5287,N_3712,N_4211);
nor U5288 (N_5288,N_2786,N_2840);
nand U5289 (N_5289,N_3027,N_4510);
and U5290 (N_5290,N_3883,N_4064);
nand U5291 (N_5291,N_4300,N_3595);
or U5292 (N_5292,N_2526,N_4262);
or U5293 (N_5293,N_4688,N_4519);
and U5294 (N_5294,N_3054,N_4907);
nor U5295 (N_5295,N_3179,N_4858);
or U5296 (N_5296,N_4244,N_4963);
and U5297 (N_5297,N_2568,N_4162);
or U5298 (N_5298,N_2957,N_3318);
nor U5299 (N_5299,N_4981,N_3163);
nand U5300 (N_5300,N_2848,N_4491);
nor U5301 (N_5301,N_4882,N_3551);
nor U5302 (N_5302,N_4556,N_3432);
or U5303 (N_5303,N_2948,N_2964);
or U5304 (N_5304,N_3646,N_3611);
and U5305 (N_5305,N_2956,N_4727);
and U5306 (N_5306,N_3113,N_3265);
nor U5307 (N_5307,N_4888,N_4239);
and U5308 (N_5308,N_2643,N_3892);
nand U5309 (N_5309,N_4466,N_2738);
nand U5310 (N_5310,N_4065,N_3784);
and U5311 (N_5311,N_4871,N_4674);
and U5312 (N_5312,N_2887,N_4127);
or U5313 (N_5313,N_4016,N_3238);
xnor U5314 (N_5314,N_4788,N_3190);
or U5315 (N_5315,N_4441,N_4569);
nor U5316 (N_5316,N_3048,N_3224);
nor U5317 (N_5317,N_4316,N_4097);
nor U5318 (N_5318,N_2524,N_3496);
nand U5319 (N_5319,N_4703,N_4299);
or U5320 (N_5320,N_4986,N_3347);
or U5321 (N_5321,N_4757,N_2658);
or U5322 (N_5322,N_4178,N_3041);
or U5323 (N_5323,N_3879,N_4233);
nand U5324 (N_5324,N_2519,N_4898);
and U5325 (N_5325,N_4929,N_4198);
nand U5326 (N_5326,N_4334,N_3627);
or U5327 (N_5327,N_2774,N_2866);
nand U5328 (N_5328,N_4390,N_4801);
nand U5329 (N_5329,N_3782,N_2669);
and U5330 (N_5330,N_4196,N_4489);
and U5331 (N_5331,N_3305,N_4967);
nand U5332 (N_5332,N_4826,N_3586);
and U5333 (N_5333,N_2749,N_3550);
nor U5334 (N_5334,N_4301,N_4849);
or U5335 (N_5335,N_4896,N_4804);
or U5336 (N_5336,N_3268,N_4132);
and U5337 (N_5337,N_2879,N_4323);
and U5338 (N_5338,N_3308,N_2858);
nand U5339 (N_5339,N_4036,N_4921);
and U5340 (N_5340,N_2752,N_3366);
nor U5341 (N_5341,N_3903,N_3507);
nor U5342 (N_5342,N_4475,N_4550);
nor U5343 (N_5343,N_3316,N_2777);
and U5344 (N_5344,N_4537,N_4593);
or U5345 (N_5345,N_4850,N_2842);
nand U5346 (N_5346,N_4517,N_3178);
and U5347 (N_5347,N_2716,N_4803);
or U5348 (N_5348,N_4226,N_3639);
nand U5349 (N_5349,N_3321,N_3346);
or U5350 (N_5350,N_2971,N_4536);
nor U5351 (N_5351,N_4251,N_3406);
and U5352 (N_5352,N_3056,N_4017);
nor U5353 (N_5353,N_3239,N_3183);
and U5354 (N_5354,N_3259,N_3925);
nand U5355 (N_5355,N_2847,N_4617);
and U5356 (N_5356,N_2505,N_3719);
nand U5357 (N_5357,N_3401,N_4409);
and U5358 (N_5358,N_2812,N_2570);
nor U5359 (N_5359,N_4446,N_2567);
or U5360 (N_5360,N_4778,N_2881);
or U5361 (N_5361,N_2511,N_4189);
nor U5362 (N_5362,N_3263,N_4318);
nand U5363 (N_5363,N_4159,N_4220);
or U5364 (N_5364,N_4500,N_4548);
nand U5365 (N_5365,N_2757,N_4203);
nand U5366 (N_5366,N_3602,N_4980);
and U5367 (N_5367,N_2684,N_3029);
nand U5368 (N_5368,N_4275,N_2628);
and U5369 (N_5369,N_2664,N_4573);
or U5370 (N_5370,N_3880,N_3888);
nor U5371 (N_5371,N_2852,N_3952);
or U5372 (N_5372,N_4532,N_4968);
or U5373 (N_5373,N_3833,N_3917);
nand U5374 (N_5374,N_2800,N_4171);
nor U5375 (N_5375,N_2877,N_4120);
xnor U5376 (N_5376,N_2934,N_2950);
nor U5377 (N_5377,N_2867,N_3805);
nand U5378 (N_5378,N_4665,N_4339);
or U5379 (N_5379,N_2714,N_3001);
or U5380 (N_5380,N_2701,N_4373);
nand U5381 (N_5381,N_4700,N_4405);
or U5382 (N_5382,N_2532,N_3978);
and U5383 (N_5383,N_4279,N_4201);
nor U5384 (N_5384,N_3077,N_4155);
nand U5385 (N_5385,N_4915,N_3728);
nor U5386 (N_5386,N_3244,N_4576);
nor U5387 (N_5387,N_4520,N_3021);
or U5388 (N_5388,N_2634,N_4830);
and U5389 (N_5389,N_2949,N_4386);
and U5390 (N_5390,N_2986,N_3002);
or U5391 (N_5391,N_4448,N_3609);
nor U5392 (N_5392,N_3407,N_3320);
nand U5393 (N_5393,N_4009,N_2618);
or U5394 (N_5394,N_3266,N_4184);
and U5395 (N_5395,N_4790,N_3528);
nor U5396 (N_5396,N_3596,N_4987);
and U5397 (N_5397,N_3870,N_2577);
nor U5398 (N_5398,N_3484,N_4304);
or U5399 (N_5399,N_2942,N_2735);
nor U5400 (N_5400,N_2951,N_3334);
or U5401 (N_5401,N_3293,N_2720);
nand U5402 (N_5402,N_3968,N_2544);
nor U5403 (N_5403,N_4340,N_2647);
or U5404 (N_5404,N_3272,N_3884);
nand U5405 (N_5405,N_3374,N_4786);
or U5406 (N_5406,N_3590,N_2909);
nand U5407 (N_5407,N_2506,N_3720);
or U5408 (N_5408,N_4690,N_3468);
nand U5409 (N_5409,N_2687,N_4128);
and U5410 (N_5410,N_2911,N_4506);
or U5411 (N_5411,N_4608,N_2649);
and U5412 (N_5412,N_3022,N_3688);
nand U5413 (N_5413,N_3329,N_3827);
or U5414 (N_5414,N_4214,N_2553);
and U5415 (N_5415,N_4253,N_3993);
nand U5416 (N_5416,N_4952,N_3772);
nand U5417 (N_5417,N_4669,N_3289);
nand U5418 (N_5418,N_2706,N_2868);
and U5419 (N_5419,N_3288,N_3157);
nor U5420 (N_5420,N_2962,N_4497);
and U5421 (N_5421,N_4337,N_2928);
or U5422 (N_5422,N_3658,N_4450);
nand U5423 (N_5423,N_3094,N_3101);
and U5424 (N_5424,N_3659,N_4422);
nand U5425 (N_5425,N_3878,N_3456);
nand U5426 (N_5426,N_3378,N_2766);
nand U5427 (N_5427,N_4854,N_2695);
nor U5428 (N_5428,N_4490,N_3575);
nand U5429 (N_5429,N_4435,N_4524);
nor U5430 (N_5430,N_4762,N_3859);
and U5431 (N_5431,N_4935,N_3354);
nor U5432 (N_5432,N_4540,N_4886);
nor U5433 (N_5433,N_3065,N_3449);
nand U5434 (N_5434,N_4207,N_2973);
nand U5435 (N_5435,N_3801,N_4683);
or U5436 (N_5436,N_3742,N_3994);
or U5437 (N_5437,N_4924,N_2859);
and U5438 (N_5438,N_2900,N_2631);
or U5439 (N_5439,N_3831,N_4163);
and U5440 (N_5440,N_2824,N_4911);
nor U5441 (N_5441,N_2958,N_4057);
and U5442 (N_5442,N_4964,N_2822);
and U5443 (N_5443,N_3256,N_3052);
or U5444 (N_5444,N_4232,N_4391);
nand U5445 (N_5445,N_4875,N_4884);
nor U5446 (N_5446,N_3618,N_4355);
or U5447 (N_5447,N_4751,N_4705);
or U5448 (N_5448,N_2883,N_3455);
or U5449 (N_5449,N_3699,N_4217);
nor U5450 (N_5450,N_4770,N_3298);
and U5451 (N_5451,N_4842,N_4425);
nor U5452 (N_5452,N_4480,N_3781);
nand U5453 (N_5453,N_3386,N_3073);
nand U5454 (N_5454,N_4427,N_3039);
nor U5455 (N_5455,N_2920,N_3282);
nand U5456 (N_5456,N_3953,N_4173);
nand U5457 (N_5457,N_3759,N_4483);
and U5458 (N_5458,N_4796,N_4908);
and U5459 (N_5459,N_2699,N_3945);
or U5460 (N_5460,N_3349,N_4523);
nand U5461 (N_5461,N_4124,N_3559);
or U5462 (N_5462,N_4701,N_4158);
nor U5463 (N_5463,N_2968,N_3090);
and U5464 (N_5464,N_2975,N_3848);
and U5465 (N_5465,N_2789,N_3898);
nand U5466 (N_5466,N_3376,N_4841);
and U5467 (N_5467,N_3750,N_3445);
and U5468 (N_5468,N_4815,N_2870);
or U5469 (N_5469,N_3079,N_2502);
and U5470 (N_5470,N_3398,N_3617);
and U5471 (N_5471,N_3206,N_4867);
nand U5472 (N_5472,N_4027,N_3393);
nor U5473 (N_5473,N_3436,N_4603);
and U5474 (N_5474,N_2712,N_4807);
or U5475 (N_5475,N_2686,N_2901);
nand U5476 (N_5476,N_3194,N_4282);
and U5477 (N_5477,N_2989,N_2835);
or U5478 (N_5478,N_3890,N_4077);
and U5479 (N_5479,N_3585,N_3013);
nand U5480 (N_5480,N_3623,N_4145);
and U5481 (N_5481,N_4799,N_4678);
or U5482 (N_5482,N_3311,N_3531);
nand U5483 (N_5483,N_4925,N_4130);
or U5484 (N_5484,N_3234,N_4384);
or U5485 (N_5485,N_4177,N_4153);
nor U5486 (N_5486,N_4948,N_4063);
nor U5487 (N_5487,N_4954,N_3304);
nor U5488 (N_5488,N_3718,N_3975);
nor U5489 (N_5489,N_4484,N_3292);
or U5490 (N_5490,N_3744,N_2813);
and U5491 (N_5491,N_3404,N_4744);
nor U5492 (N_5492,N_3989,N_4136);
nor U5493 (N_5493,N_4718,N_3988);
nand U5494 (N_5494,N_4873,N_4138);
nor U5495 (N_5495,N_4558,N_3854);
or U5496 (N_5496,N_3322,N_4464);
or U5497 (N_5497,N_4643,N_3005);
nand U5498 (N_5498,N_4930,N_4917);
or U5499 (N_5499,N_3426,N_3191);
nor U5500 (N_5500,N_3245,N_3900);
nor U5501 (N_5501,N_4094,N_3689);
nor U5502 (N_5502,N_4661,N_4182);
nor U5503 (N_5503,N_3863,N_2967);
nand U5504 (N_5504,N_3522,N_4732);
or U5505 (N_5505,N_3760,N_2981);
nand U5506 (N_5506,N_3984,N_3461);
and U5507 (N_5507,N_2996,N_3332);
and U5508 (N_5508,N_4950,N_4473);
nand U5509 (N_5509,N_2534,N_3126);
nor U5510 (N_5510,N_4099,N_3400);
and U5511 (N_5511,N_4463,N_4715);
nor U5512 (N_5512,N_3387,N_4338);
nand U5513 (N_5513,N_4147,N_4539);
nand U5514 (N_5514,N_3545,N_3807);
nor U5515 (N_5515,N_4443,N_4920);
nor U5516 (N_5516,N_2736,N_4112);
nand U5517 (N_5517,N_2551,N_3246);
nand U5518 (N_5518,N_3379,N_4931);
nand U5519 (N_5519,N_2763,N_3891);
or U5520 (N_5520,N_4529,N_3800);
nor U5521 (N_5521,N_3319,N_4759);
or U5522 (N_5522,N_3228,N_4181);
and U5523 (N_5523,N_3707,N_3841);
and U5524 (N_5524,N_2501,N_4090);
or U5525 (N_5525,N_3476,N_3254);
nor U5526 (N_5526,N_3260,N_4599);
and U5527 (N_5527,N_3587,N_4294);
nand U5528 (N_5528,N_3140,N_3710);
and U5529 (N_5529,N_4246,N_4221);
and U5530 (N_5530,N_3222,N_3730);
nand U5531 (N_5531,N_3000,N_4439);
and U5532 (N_5532,N_4487,N_3276);
or U5533 (N_5533,N_3115,N_2569);
or U5534 (N_5534,N_3044,N_4834);
nor U5535 (N_5535,N_4847,N_3328);
and U5536 (N_5536,N_3576,N_4572);
nand U5537 (N_5537,N_2638,N_3264);
or U5538 (N_5538,N_4381,N_4314);
nand U5539 (N_5539,N_3411,N_2843);
and U5540 (N_5540,N_4997,N_2905);
nor U5541 (N_5541,N_3675,N_4083);
and U5542 (N_5542,N_3495,N_2711);
nor U5543 (N_5543,N_4327,N_4357);
and U5544 (N_5544,N_2850,N_3836);
and U5545 (N_5545,N_3642,N_4276);
and U5546 (N_5546,N_3861,N_4440);
nor U5547 (N_5547,N_3306,N_4000);
or U5548 (N_5548,N_4471,N_4252);
nand U5549 (N_5549,N_2733,N_3489);
xnor U5550 (N_5550,N_3068,N_3154);
nand U5551 (N_5551,N_3300,N_4319);
nor U5552 (N_5552,N_3098,N_3907);
or U5553 (N_5553,N_2744,N_4292);
or U5554 (N_5554,N_3210,N_3631);
nor U5555 (N_5555,N_3790,N_2795);
nand U5556 (N_5556,N_4308,N_2705);
or U5557 (N_5557,N_4190,N_3488);
nand U5558 (N_5558,N_4597,N_3133);
and U5559 (N_5559,N_2679,N_2960);
and U5560 (N_5560,N_3716,N_3158);
or U5561 (N_5561,N_3629,N_3942);
and U5562 (N_5562,N_3969,N_4709);
and U5563 (N_5563,N_4712,N_3340);
nor U5564 (N_5564,N_4002,N_3249);
and U5565 (N_5565,N_2972,N_3051);
nand U5566 (N_5566,N_4258,N_3604);
nand U5567 (N_5567,N_4001,N_3153);
nor U5568 (N_5568,N_3416,N_2836);
nor U5569 (N_5569,N_4295,N_2713);
nor U5570 (N_5570,N_3974,N_3267);
nand U5571 (N_5571,N_3851,N_4164);
nor U5572 (N_5572,N_4310,N_4071);
or U5573 (N_5573,N_2880,N_3947);
and U5574 (N_5574,N_4554,N_3480);
and U5575 (N_5575,N_4169,N_4351);
or U5576 (N_5576,N_3487,N_4485);
nand U5577 (N_5577,N_3460,N_3345);
or U5578 (N_5578,N_2839,N_4256);
and U5579 (N_5579,N_2979,N_4605);
and U5580 (N_5580,N_3748,N_4923);
nand U5581 (N_5581,N_4602,N_3817);
nand U5582 (N_5582,N_2992,N_4566);
nor U5583 (N_5583,N_3563,N_4795);
and U5584 (N_5584,N_4011,N_3015);
nand U5585 (N_5585,N_2910,N_3668);
nand U5586 (N_5586,N_4691,N_4660);
nor U5587 (N_5587,N_4160,N_4959);
or U5588 (N_5588,N_3117,N_3135);
nand U5589 (N_5589,N_4419,N_4414);
and U5590 (N_5590,N_4714,N_4889);
nor U5591 (N_5591,N_3286,N_3799);
or U5592 (N_5592,N_2700,N_4937);
or U5593 (N_5593,N_4656,N_2547);
xor U5594 (N_5594,N_3926,N_4735);
nand U5595 (N_5595,N_4686,N_2646);
and U5596 (N_5596,N_4429,N_3895);
or U5597 (N_5597,N_3294,N_4421);
and U5598 (N_5598,N_3765,N_3450);
nand U5599 (N_5599,N_4454,N_2609);
nor U5600 (N_5600,N_3657,N_4066);
nor U5601 (N_5601,N_2509,N_3182);
or U5602 (N_5602,N_4802,N_3151);
and U5603 (N_5603,N_3679,N_3503);
or U5604 (N_5604,N_2977,N_4103);
nor U5605 (N_5605,N_4562,N_3887);
or U5606 (N_5606,N_4129,N_4058);
nand U5607 (N_5607,N_4105,N_3755);
nand U5608 (N_5608,N_2674,N_3091);
and U5609 (N_5609,N_3966,N_2535);
or U5610 (N_5610,N_4983,N_4352);
nor U5611 (N_5611,N_4552,N_3207);
and U5612 (N_5612,N_3148,N_4777);
and U5613 (N_5613,N_4449,N_4407);
nand U5614 (N_5614,N_3633,N_4459);
nand U5615 (N_5615,N_2663,N_2806);
nor U5616 (N_5616,N_3549,N_3314);
and U5617 (N_5617,N_3770,N_4798);
nor U5618 (N_5618,N_3192,N_3008);
and U5619 (N_5619,N_4168,N_3369);
and U5620 (N_5620,N_3018,N_2861);
or U5621 (N_5621,N_3832,N_4269);
and U5622 (N_5622,N_4359,N_3119);
and U5623 (N_5623,N_4518,N_3336);
nor U5624 (N_5624,N_4028,N_4406);
nor U5625 (N_5625,N_3666,N_2896);
xnor U5626 (N_5626,N_2851,N_3023);
nand U5627 (N_5627,N_4609,N_4047);
and U5628 (N_5628,N_4349,N_4613);
nand U5629 (N_5629,N_4627,N_4502);
nand U5630 (N_5630,N_3684,N_3991);
and U5631 (N_5631,N_4412,N_3233);
and U5632 (N_5632,N_3669,N_4645);
or U5633 (N_5633,N_2869,N_4637);
and U5634 (N_5634,N_4823,N_3392);
or U5635 (N_5635,N_4792,N_4965);
nor U5636 (N_5636,N_4794,N_3721);
nand U5637 (N_5637,N_4042,N_4994);
nand U5638 (N_5638,N_2970,N_4468);
and U5639 (N_5639,N_3934,N_3351);
and U5640 (N_5640,N_3327,N_2723);
nand U5641 (N_5641,N_4141,N_4673);
nor U5642 (N_5642,N_3046,N_4034);
or U5643 (N_5643,N_4571,N_2775);
and U5644 (N_5644,N_2919,N_4836);
nand U5645 (N_5645,N_3483,N_3004);
and U5646 (N_5646,N_3080,N_4423);
or U5647 (N_5647,N_4722,N_3906);
and U5648 (N_5648,N_4461,N_2517);
nand U5649 (N_5649,N_4303,N_4175);
nand U5650 (N_5650,N_3965,N_4150);
and U5651 (N_5651,N_4290,N_4006);
nor U5652 (N_5652,N_4767,N_2797);
and U5653 (N_5653,N_3904,N_4342);
or U5654 (N_5654,N_3830,N_3352);
and U5655 (N_5655,N_2885,N_3372);
nor U5656 (N_5656,N_4962,N_2904);
nand U5657 (N_5657,N_3435,N_4912);
or U5658 (N_5658,N_3452,N_3490);
or U5659 (N_5659,N_3084,N_4813);
or U5660 (N_5660,N_3853,N_2725);
nor U5661 (N_5661,N_4462,N_3180);
or U5662 (N_5662,N_3527,N_4332);
and U5663 (N_5663,N_4174,N_2635);
nor U5664 (N_5664,N_2651,N_3746);
or U5665 (N_5665,N_4708,N_3198);
nand U5666 (N_5666,N_2925,N_4675);
nand U5667 (N_5667,N_3383,N_3440);
or U5668 (N_5668,N_4693,N_3255);
nand U5669 (N_5669,N_4559,N_2721);
and U5670 (N_5670,N_4616,N_4877);
and U5671 (N_5671,N_4565,N_4234);
and U5672 (N_5672,N_4452,N_2764);
nand U5673 (N_5673,N_4775,N_2939);
and U5674 (N_5674,N_3902,N_4816);
nor U5675 (N_5675,N_3257,N_4606);
or U5676 (N_5676,N_3012,N_3377);
nor U5677 (N_5677,N_3715,N_2871);
nand U5678 (N_5678,N_2838,N_2627);
nor U5679 (N_5679,N_2811,N_4317);
nor U5680 (N_5680,N_3035,N_2878);
and U5681 (N_5681,N_4346,N_2653);
and U5682 (N_5682,N_3203,N_4081);
nor U5683 (N_5683,N_3824,N_3231);
and U5684 (N_5684,N_3105,N_4271);
or U5685 (N_5685,N_4639,N_3982);
or U5686 (N_5686,N_2654,N_4814);
and U5687 (N_5687,N_4152,N_3025);
and U5688 (N_5688,N_3092,N_4243);
or U5689 (N_5689,N_4051,N_4410);
nand U5690 (N_5690,N_3823,N_2805);
and U5691 (N_5691,N_3324,N_3722);
nor U5692 (N_5692,N_3433,N_4577);
nor U5693 (N_5693,N_3537,N_4101);
nor U5694 (N_5694,N_3913,N_3874);
nand U5695 (N_5695,N_2872,N_3425);
nand U5696 (N_5696,N_2918,N_4862);
nand U5697 (N_5697,N_2966,N_4622);
nand U5698 (N_5698,N_4694,N_4878);
nor U5699 (N_5699,N_3843,N_3076);
nor U5700 (N_5700,N_4748,N_3127);
nor U5701 (N_5701,N_4947,N_3248);
nor U5702 (N_5702,N_3787,N_2599);
and U5703 (N_5703,N_2508,N_3038);
or U5704 (N_5704,N_2820,N_3959);
or U5705 (N_5705,N_2974,N_3270);
or U5706 (N_5706,N_2585,N_4456);
nand U5707 (N_5707,N_3794,N_3277);
or U5708 (N_5708,N_3608,N_3437);
and U5709 (N_5709,N_3571,N_3804);
or U5710 (N_5710,N_3555,N_3427);
nand U5711 (N_5711,N_4940,N_4119);
nand U5712 (N_5712,N_2845,N_3663);
nand U5713 (N_5713,N_4100,N_3162);
and U5714 (N_5714,N_3737,N_3592);
nand U5715 (N_5715,N_4743,N_4692);
nand U5716 (N_5716,N_4052,N_2750);
nor U5717 (N_5717,N_3457,N_4549);
nand U5718 (N_5718,N_2903,N_3598);
nor U5719 (N_5719,N_3463,N_4313);
or U5720 (N_5720,N_3439,N_3072);
and U5721 (N_5721,N_2930,N_2912);
or U5722 (N_5722,N_2652,N_2853);
and U5723 (N_5723,N_4289,N_4706);
nor U5724 (N_5724,N_3901,N_3873);
and U5725 (N_5725,N_2576,N_4235);
nor U5726 (N_5726,N_3667,N_4067);
and U5727 (N_5727,N_4266,N_3924);
and U5728 (N_5728,N_4123,N_3578);
nand U5729 (N_5729,N_4222,N_4629);
or U5730 (N_5730,N_4325,N_3141);
or U5731 (N_5731,N_2655,N_2612);
or U5732 (N_5732,N_2888,N_3434);
and U5733 (N_5733,N_4453,N_3287);
nor U5734 (N_5734,N_4900,N_4068);
or U5735 (N_5735,N_3032,N_3656);
xor U5736 (N_5736,N_3665,N_4089);
or U5737 (N_5737,N_3413,N_4049);
nor U5738 (N_5738,N_2510,N_4131);
nor U5739 (N_5739,N_3714,N_3299);
or U5740 (N_5740,N_4035,N_4442);
nor U5741 (N_5741,N_3513,N_3921);
or U5742 (N_5742,N_3521,N_3727);
or U5743 (N_5743,N_4805,N_3059);
and U5744 (N_5744,N_2581,N_4531);
and U5745 (N_5745,N_4496,N_4969);
and U5746 (N_5746,N_4644,N_4507);
and U5747 (N_5747,N_3395,N_3373);
nor U5748 (N_5748,N_2680,N_4218);
or U5749 (N_5749,N_2611,N_3174);
nor U5750 (N_5750,N_3451,N_3849);
or U5751 (N_5751,N_3216,N_4227);
or U5752 (N_5752,N_3359,N_4007);
nand U5753 (N_5753,N_4872,N_3343);
and U5754 (N_5754,N_4379,N_4567);
nor U5755 (N_5755,N_3767,N_4354);
nor U5756 (N_5756,N_4955,N_4263);
or U5757 (N_5757,N_3410,N_4096);
nand U5758 (N_5758,N_3725,N_3514);
nor U5759 (N_5759,N_4024,N_3992);
or U5760 (N_5760,N_2525,N_2662);
nand U5761 (N_5761,N_2726,N_3743);
and U5762 (N_5762,N_3227,N_4324);
or U5763 (N_5763,N_4255,N_3894);
nor U5764 (N_5764,N_3302,N_4482);
or U5765 (N_5765,N_2671,N_2528);
nand U5766 (N_5766,N_2921,N_2999);
nand U5767 (N_5767,N_2993,N_3543);
nand U5768 (N_5768,N_3539,N_4018);
nor U5769 (N_5769,N_4560,N_4200);
or U5770 (N_5770,N_4897,N_2983);
or U5771 (N_5771,N_3236,N_3882);
nor U5772 (N_5772,N_4161,N_4615);
nor U5773 (N_5773,N_4812,N_3462);
and U5774 (N_5774,N_3905,N_3250);
nand U5775 (N_5775,N_2644,N_3066);
nor U5776 (N_5776,N_2724,N_2814);
or U5777 (N_5777,N_4589,N_3499);
nand U5778 (N_5778,N_3971,N_3283);
or U5779 (N_5779,N_3498,N_4498);
xnor U5780 (N_5780,N_4307,N_4040);
and U5781 (N_5781,N_4546,N_2965);
nand U5782 (N_5782,N_4731,N_3803);
and U5783 (N_5783,N_3818,N_3132);
and U5784 (N_5784,N_4144,N_3017);
nor U5785 (N_5785,N_4320,N_3793);
nor U5786 (N_5786,N_2916,N_4628);
and U5787 (N_5787,N_4728,N_4492);
or U5788 (N_5788,N_3385,N_3753);
nor U5789 (N_5789,N_4806,N_3242);
or U5790 (N_5790,N_4684,N_3756);
and U5791 (N_5791,N_4730,N_4509);
nor U5792 (N_5792,N_3420,N_4254);
xor U5793 (N_5793,N_2507,N_4260);
and U5794 (N_5794,N_4835,N_4015);
nand U5795 (N_5795,N_2521,N_4846);
or U5796 (N_5796,N_3269,N_3405);
and U5797 (N_5797,N_4328,N_4914);
nor U5798 (N_5798,N_4508,N_3593);
or U5799 (N_5799,N_3262,N_3071);
and U5800 (N_5800,N_3047,N_3424);
or U5801 (N_5801,N_4165,N_4192);
and U5802 (N_5802,N_3070,N_3775);
and U5803 (N_5803,N_3187,N_2941);
nor U5804 (N_5804,N_4433,N_3475);
and U5805 (N_5805,N_4903,N_3601);
and U5806 (N_5806,N_3364,N_3858);
and U5807 (N_5807,N_2530,N_3443);
and U5808 (N_5808,N_2500,N_3673);
nand U5809 (N_5809,N_3355,N_4513);
and U5810 (N_5810,N_2685,N_4868);
and U5811 (N_5811,N_2787,N_4401);
nor U5812 (N_5812,N_3839,N_3186);
or U5813 (N_5813,N_4072,N_3466);
or U5814 (N_5814,N_4356,N_2923);
or U5815 (N_5815,N_4380,N_2785);
and U5816 (N_5816,N_4474,N_4721);
nand U5817 (N_5817,N_3144,N_3348);
and U5818 (N_5818,N_4624,N_4102);
or U5819 (N_5819,N_3368,N_4740);
nor U5820 (N_5820,N_2917,N_4364);
nor U5821 (N_5821,N_2799,N_3613);
or U5822 (N_5822,N_4374,N_3865);
and U5823 (N_5823,N_2602,N_4023);
nand U5824 (N_5824,N_3176,N_2994);
or U5825 (N_5825,N_4245,N_4634);
nor U5826 (N_5826,N_3281,N_4710);
and U5827 (N_5827,N_2554,N_3644);
or U5828 (N_5828,N_3897,N_2876);
or U5829 (N_5829,N_3778,N_4810);
and U5830 (N_5830,N_3694,N_3875);
nand U5831 (N_5831,N_4662,N_4392);
nor U5832 (N_5832,N_4756,N_3344);
and U5833 (N_5833,N_4652,N_3494);
or U5834 (N_5834,N_3384,N_4635);
or U5835 (N_5835,N_3279,N_3687);
nor U5836 (N_5836,N_4564,N_3196);
and U5837 (N_5837,N_3811,N_4445);
or U5838 (N_5838,N_4135,N_3970);
nand U5839 (N_5839,N_4820,N_4237);
and U5840 (N_5840,N_2605,N_3310);
or U5841 (N_5841,N_2790,N_4467);
nand U5842 (N_5842,N_4048,N_3607);
nand U5843 (N_5843,N_4367,N_4975);
or U5844 (N_5844,N_3583,N_4366);
nor U5845 (N_5845,N_2755,N_4870);
or U5846 (N_5846,N_2541,N_2615);
nand U5847 (N_5847,N_4115,N_4626);
and U5848 (N_5848,N_2863,N_4741);
or U5849 (N_5849,N_2616,N_3491);
nor U5850 (N_5850,N_3860,N_2683);
nor U5851 (N_5851,N_4753,N_4829);
and U5852 (N_5852,N_2734,N_4372);
nor U5853 (N_5853,N_4885,N_4118);
or U5854 (N_5854,N_4447,N_3866);
and U5855 (N_5855,N_2656,N_3573);
and U5856 (N_5856,N_4972,N_2557);
nand U5857 (N_5857,N_2802,N_2767);
nor U5858 (N_5858,N_3069,N_3661);
nor U5859 (N_5859,N_4851,N_3554);
or U5860 (N_5860,N_4666,N_2708);
or U5861 (N_5861,N_2660,N_3428);
or U5862 (N_5862,N_3172,N_3212);
and U5863 (N_5863,N_2620,N_3652);
or U5864 (N_5864,N_2746,N_3889);
or U5865 (N_5865,N_2613,N_2762);
and U5866 (N_5866,N_4378,N_3733);
nor U5867 (N_5867,N_4636,N_4771);
nand U5868 (N_5868,N_2927,N_2985);
and U5869 (N_5869,N_4216,N_3738);
or U5870 (N_5870,N_4109,N_4430);
nand U5871 (N_5871,N_3454,N_3768);
nand U5872 (N_5872,N_4098,N_4887);
or U5873 (N_5873,N_4134,N_3789);
nand U5874 (N_5874,N_3271,N_4583);
nor U5875 (N_5875,N_3695,N_4167);
nor U5876 (N_5876,N_3677,N_3213);
or U5877 (N_5877,N_4312,N_3995);
or U5878 (N_5878,N_3492,N_3109);
or U5879 (N_5879,N_4960,N_4892);
and U5880 (N_5880,N_4953,N_3990);
nand U5881 (N_5881,N_4677,N_2821);
nand U5882 (N_5882,N_2731,N_2860);
nand U5883 (N_5883,N_3217,N_2675);
or U5884 (N_5884,N_2637,N_3713);
or U5885 (N_5885,N_3003,N_3195);
or U5886 (N_5886,N_3478,N_3612);
and U5887 (N_5887,N_4579,N_3662);
nor U5888 (N_5888,N_4993,N_2640);
and U5889 (N_5889,N_3088,N_2819);
nand U5890 (N_5890,N_3747,N_3820);
and U5891 (N_5891,N_3780,N_3055);
and U5892 (N_5892,N_4315,N_4857);
nor U5893 (N_5893,N_4866,N_2907);
nor U5894 (N_5894,N_4676,N_4149);
nor U5895 (N_5895,N_3655,N_3438);
or U5896 (N_5896,N_3166,N_3828);
nor U5897 (N_5897,N_3548,N_3223);
nor U5898 (N_5898,N_4183,N_4734);
nand U5899 (N_5899,N_3014,N_4272);
and U5900 (N_5900,N_3754,N_3896);
and U5901 (N_5901,N_2648,N_3221);
and U5902 (N_5902,N_2884,N_3998);
nand U5903 (N_5903,N_3448,N_2678);
nand U5904 (N_5904,N_2555,N_4904);
nand U5905 (N_5905,N_3763,N_4350);
nand U5906 (N_5906,N_3371,N_3089);
and U5907 (N_5907,N_4085,N_3331);
nor U5908 (N_5908,N_2959,N_3532);
and U5909 (N_5909,N_4982,N_4647);
and U5910 (N_5910,N_3278,N_3111);
nand U5911 (N_5911,N_4557,N_4707);
and U5912 (N_5912,N_4250,N_2929);
and U5913 (N_5913,N_2586,N_2829);
or U5914 (N_5914,N_4465,N_4268);
nand U5915 (N_5915,N_2793,N_4336);
and U5916 (N_5916,N_4768,N_4584);
and U5917 (N_5917,N_2817,N_4389);
nand U5918 (N_5918,N_4213,N_2564);
nor U5919 (N_5919,N_3950,N_3409);
or U5920 (N_5920,N_3758,N_3520);
and U5921 (N_5921,N_2536,N_2808);
and U5922 (N_5922,N_4444,N_2606);
or U5923 (N_5923,N_3511,N_2882);
nor U5924 (N_5924,N_3651,N_4891);
and U5925 (N_5925,N_2574,N_4212);
and U5926 (N_5926,N_4764,N_2754);
nand U5927 (N_5927,N_3125,N_4631);
and U5928 (N_5928,N_3317,N_3184);
or U5929 (N_5929,N_4736,N_3412);
nand U5930 (N_5930,N_4863,N_3566);
and U5931 (N_5931,N_3229,N_4062);
nor U5932 (N_5932,N_2936,N_3852);
nor U5933 (N_5933,N_3577,N_3415);
and U5934 (N_5934,N_2831,N_4286);
or U5935 (N_5935,N_3654,N_2520);
and U5936 (N_5936,N_3977,N_3936);
and U5937 (N_5937,N_4460,N_3326);
nand U5938 (N_5938,N_4784,N_4146);
nor U5939 (N_5939,N_4206,N_4946);
and U5940 (N_5940,N_4895,N_4521);
or U5941 (N_5941,N_2703,N_2984);
xor U5942 (N_5942,N_3159,N_3164);
and U5943 (N_5943,N_3358,N_3556);
nor U5944 (N_5944,N_4890,N_2830);
and U5945 (N_5945,N_4679,N_3812);
or U5946 (N_5946,N_2892,N_4781);
and U5947 (N_5947,N_3649,N_4588);
and U5948 (N_5948,N_4995,N_3815);
nor U5949 (N_5949,N_3337,N_3706);
nand U5950 (N_5950,N_3493,N_4689);
nand U5951 (N_5951,N_3638,N_4725);
or U5952 (N_5952,N_3997,N_3869);
or U5953 (N_5953,N_2629,N_4511);
nor U5954 (N_5954,N_3469,N_3798);
or U5955 (N_5955,N_3937,N_2798);
or U5956 (N_5956,N_4843,N_3682);
nor U5957 (N_5957,N_3620,N_4961);
or U5958 (N_5958,N_3131,N_4488);
and U5959 (N_5959,N_3421,N_4287);
or U5960 (N_5960,N_3881,N_3692);
xor U5961 (N_5961,N_3189,N_3303);
or U5962 (N_5962,N_4879,N_3672);
or U5963 (N_5963,N_3584,N_3582);
nand U5964 (N_5964,N_4093,N_3636);
nand U5965 (N_5965,N_3785,N_4699);
or U5966 (N_5966,N_3388,N_2953);
and U5967 (N_5967,N_4004,N_3864);
and U5968 (N_5968,N_3580,N_2940);
or U5969 (N_5969,N_2955,N_2715);
nand U5970 (N_5970,N_2874,N_4045);
or U5971 (N_5971,N_2815,N_3847);
or U5972 (N_5972,N_2673,N_3717);
or U5973 (N_5973,N_3786,N_4720);
or U5974 (N_5974,N_4818,N_3323);
nor U5975 (N_5975,N_3028,N_3572);
and U5976 (N_5976,N_3284,N_3275);
nand U5977 (N_5977,N_3569,N_4979);
nand U5978 (N_5978,N_4087,N_4545);
or U5979 (N_5979,N_4104,N_4142);
nor U5980 (N_5980,N_4361,N_3274);
xor U5981 (N_5981,N_4228,N_4612);
and U5982 (N_5982,N_4114,N_2677);
or U5983 (N_5983,N_3016,N_2625);
and U5984 (N_5984,N_3430,N_2739);
and U5985 (N_5985,N_2603,N_2931);
and U5986 (N_5986,N_3418,N_4856);
nand U5987 (N_5987,N_4408,N_4438);
nor U5988 (N_5988,N_3230,N_4074);
nand U5989 (N_5989,N_3506,N_4772);
and U5990 (N_5990,N_3872,N_3911);
or U5991 (N_5991,N_2998,N_4038);
and U5992 (N_5992,N_3766,N_3036);
nor U5993 (N_5993,N_4257,N_4348);
xnor U5994 (N_5994,N_2566,N_3809);
nand U5995 (N_5995,N_3783,N_3155);
or U5996 (N_5996,N_3634,N_4076);
or U5997 (N_5997,N_4195,N_3757);
and U5998 (N_5998,N_2982,N_2893);
nand U5999 (N_5999,N_3979,N_4426);
or U6000 (N_6000,N_4424,N_3535);
and U6001 (N_6001,N_2741,N_3724);
and U6002 (N_6002,N_4600,N_4365);
or U6003 (N_6003,N_3247,N_4428);
nand U6004 (N_6004,N_4838,N_4578);
nand U6005 (N_6005,N_4261,N_3674);
or U6006 (N_6006,N_4670,N_4277);
or U6007 (N_6007,N_3918,N_4193);
nand U6008 (N_6008,N_2782,N_2771);
and U6009 (N_6009,N_3726,N_4951);
or U6010 (N_6010,N_4043,N_3453);
and U6011 (N_6011,N_4387,N_3614);
nor U6012 (N_6012,N_2780,N_3423);
or U6013 (N_6013,N_3867,N_3910);
and U6014 (N_6014,N_3380,N_3697);
nand U6015 (N_6015,N_4876,N_3237);
nand U6016 (N_6016,N_3834,N_2571);
or U6017 (N_6017,N_4345,N_4291);
and U6018 (N_6018,N_3558,N_3251);
or U6019 (N_6019,N_2772,N_3375);
or U6020 (N_6020,N_2659,N_2563);
nand U6021 (N_6021,N_3777,N_4376);
nand U6022 (N_6022,N_4288,N_2597);
and U6023 (N_6023,N_2668,N_3908);
nand U6024 (N_6024,N_4369,N_3138);
or U6025 (N_6025,N_4311,N_4590);
and U6026 (N_6026,N_3829,N_4575);
or U6027 (N_6027,N_2773,N_3273);
nand U6028 (N_6028,N_3557,N_3944);
and U6029 (N_6029,N_3161,N_2728);
and U6030 (N_6030,N_3291,N_3232);
or U6031 (N_6031,N_3683,N_4044);
and U6032 (N_6032,N_4543,N_4432);
or U6033 (N_6033,N_4396,N_4657);
nor U6034 (N_6034,N_3540,N_3825);
or U6035 (N_6035,N_3175,N_4368);
nand U6036 (N_6036,N_3049,N_4944);
nor U6037 (N_6037,N_3647,N_2938);
nor U6038 (N_6038,N_4298,N_4385);
and U6039 (N_6039,N_3473,N_3635);
nand U6040 (N_6040,N_3552,N_3838);
nand U6041 (N_6041,N_4601,N_4241);
or U6042 (N_6042,N_4913,N_4837);
and U6043 (N_6043,N_3645,N_2779);
nor U6044 (N_6044,N_4607,N_2769);
and U6045 (N_6045,N_3389,N_4906);
or U6046 (N_6046,N_4470,N_3734);
xor U6047 (N_6047,N_4008,N_3043);
or U6048 (N_6048,N_3497,N_2770);
nand U6049 (N_6049,N_4760,N_3691);
nor U6050 (N_6050,N_4019,N_2737);
nand U6051 (N_6051,N_3732,N_4284);
nand U6052 (N_6052,N_4926,N_2902);
nor U6053 (N_6053,N_4821,N_4824);
nor U6054 (N_6054,N_2709,N_2743);
and U6055 (N_6055,N_3285,N_3104);
and U6056 (N_6056,N_3096,N_3181);
nor U6057 (N_6057,N_4431,N_2587);
and U6058 (N_6058,N_3253,N_4187);
nor U6059 (N_6059,N_3136,N_3933);
or U6060 (N_6060,N_2722,N_4055);
nor U6061 (N_6061,N_3600,N_3280);
or U6062 (N_6062,N_3764,N_3301);
or U6063 (N_6063,N_4005,N_4883);
and U6064 (N_6064,N_4711,N_2740);
nor U6065 (N_6065,N_2760,N_2862);
nand U6066 (N_6066,N_3842,N_3802);
nor U6067 (N_6067,N_4865,N_4493);
and U6068 (N_6068,N_3103,N_3146);
nand U6069 (N_6069,N_4893,N_2632);
or U6070 (N_6070,N_4370,N_4248);
and U6071 (N_6071,N_2855,N_3961);
nor U6072 (N_6072,N_2894,N_2604);
and U6073 (N_6073,N_3167,N_3797);
and U6074 (N_6074,N_2886,N_3363);
nand U6075 (N_6075,N_4582,N_3570);
nand U6076 (N_6076,N_3788,N_3871);
nand U6077 (N_6077,N_2873,N_3050);
or U6078 (N_6078,N_2952,N_3479);
and U6079 (N_6079,N_2778,N_4646);
nor U6080 (N_6080,N_4745,N_3541);
nand U6081 (N_6081,N_4151,N_3030);
or U6082 (N_6082,N_3703,N_4869);
nand U6083 (N_6083,N_4204,N_3561);
and U6084 (N_6084,N_2922,N_4591);
nand U6085 (N_6085,N_4086,N_3771);
nand U6086 (N_6086,N_2696,N_4594);
nor U6087 (N_6087,N_3472,N_4974);
nor U6088 (N_6088,N_3928,N_4746);
nor U6089 (N_6089,N_4229,N_4197);
nor U6090 (N_6090,N_4919,N_3844);
or U6091 (N_6091,N_4648,N_2578);
and U6092 (N_6092,N_3516,N_3693);
and U6093 (N_6093,N_4831,N_2591);
nor U6094 (N_6094,N_3481,N_3081);
or U6095 (N_6095,N_4859,N_2875);
or U6096 (N_6096,N_4909,N_3208);
or U6097 (N_6097,N_3935,N_3983);
nor U6098 (N_6098,N_3403,N_4170);
nand U6099 (N_6099,N_3632,N_4659);
nor U6100 (N_6100,N_3956,N_4621);
nor U6101 (N_6101,N_3862,N_4793);
or U6102 (N_6102,N_4902,N_3325);
nand U6103 (N_6103,N_3589,N_3517);
and U6104 (N_6104,N_2834,N_3168);
or U6105 (N_6105,N_3676,N_2943);
and U6106 (N_6106,N_2756,N_3940);
or U6107 (N_6107,N_3526,N_3143);
and U6108 (N_6108,N_3106,N_4825);
nand U6109 (N_6109,N_4377,N_3671);
and U6110 (N_6110,N_2833,N_4766);
or U6111 (N_6111,N_4265,N_3296);
nand U6112 (N_6112,N_3923,N_4936);
or U6113 (N_6113,N_4477,N_3061);
nand U6114 (N_6114,N_3603,N_3949);
nor U6115 (N_6115,N_4910,N_2565);
or U6116 (N_6116,N_3471,N_3145);
and U6117 (N_6117,N_3078,N_2590);
and U6118 (N_6118,N_3241,N_4527);
or U6119 (N_6119,N_3075,N_3909);
or U6120 (N_6120,N_3396,N_3045);
or U6121 (N_6121,N_3624,N_3628);
and U6122 (N_6122,N_4126,N_4538);
nand U6123 (N_6123,N_2579,N_4845);
or U6124 (N_6124,N_2710,N_3114);
nand U6125 (N_6125,N_3739,N_3579);
nand U6126 (N_6126,N_4382,N_3446);
nand U6127 (N_6127,N_2621,N_3920);
and U6128 (N_6128,N_4050,N_2991);
or U6129 (N_6129,N_4501,N_4992);
or U6130 (N_6130,N_4420,N_4188);
nand U6131 (N_6131,N_4797,N_3792);
and U6132 (N_6132,N_4966,N_3846);
nand U6133 (N_6133,N_4535,N_4949);
nor U6134 (N_6134,N_4285,N_4779);
nand U6135 (N_6135,N_4095,N_3795);
nand U6136 (N_6136,N_3026,N_3698);
or U6137 (N_6137,N_4393,N_3822);
nand U6138 (N_6138,N_3533,N_4654);
and U6139 (N_6139,N_4486,N_4649);
or U6140 (N_6140,N_3360,N_2702);
or U6141 (N_6141,N_4522,N_3912);
or U6142 (N_6142,N_2704,N_2987);
and U6143 (N_6143,N_4739,N_4840);
or U6144 (N_6144,N_3417,N_4274);
nor U6145 (N_6145,N_3058,N_3769);
or U6146 (N_6146,N_4998,N_4723);
nor U6147 (N_6147,N_3709,N_4713);
nand U6148 (N_6148,N_3243,N_4075);
or U6149 (N_6149,N_4054,N_4632);
nor U6150 (N_6150,N_4697,N_3007);
and U6151 (N_6151,N_3821,N_2897);
nor U6152 (N_6152,N_4512,N_4321);
nand U6153 (N_6153,N_3512,N_3185);
or U6154 (N_6154,N_4978,N_2682);
nor U6155 (N_6155,N_3641,N_3219);
nand U6156 (N_6156,N_3312,N_2768);
nand U6157 (N_6157,N_2751,N_2995);
nand U6158 (N_6158,N_3313,N_4504);
and U6159 (N_6159,N_4399,N_3010);
and U6160 (N_6160,N_4581,N_4137);
and U6161 (N_6161,N_3740,N_4436);
nand U6162 (N_6162,N_3315,N_4179);
and U6163 (N_6163,N_4928,N_2548);
and U6164 (N_6164,N_4125,N_2619);
and U6165 (N_6165,N_4225,N_4990);
nor U6166 (N_6166,N_3362,N_2969);
nor U6167 (N_6167,N_2691,N_4472);
and U6168 (N_6168,N_4528,N_4839);
nand U6169 (N_6169,N_2624,N_4827);
and U6170 (N_6170,N_3037,N_2759);
nand U6171 (N_6171,N_4984,N_2533);
nor U6172 (N_6172,N_2550,N_3731);
and U6173 (N_6173,N_2818,N_3538);
nor U6174 (N_6174,N_3447,N_3964);
and U6175 (N_6175,N_4542,N_4650);
nand U6176 (N_6176,N_2745,N_4580);
or U6177 (N_6177,N_4977,N_3220);
and U6178 (N_6178,N_2630,N_3422);
nand U6179 (N_6179,N_4640,N_3085);
and U6180 (N_6180,N_4013,N_4611);
and U6181 (N_6181,N_4610,N_2512);
nor U6182 (N_6182,N_3837,N_4755);
nor U6183 (N_6183,N_4933,N_4224);
nor U6184 (N_6184,N_2580,N_3024);
nor U6185 (N_6185,N_3813,N_2596);
nor U6186 (N_6186,N_4514,N_2788);
nand U6187 (N_6187,N_4503,N_2690);
nand U6188 (N_6188,N_3064,N_3330);
nand U6189 (N_6189,N_4641,N_4437);
nand U6190 (N_6190,N_4680,N_3591);
nor U6191 (N_6191,N_4630,N_3518);
and U6192 (N_6192,N_2598,N_4416);
nand U6193 (N_6193,N_4750,N_4819);
nor U6194 (N_6194,N_3020,N_4587);
or U6195 (N_6195,N_4259,N_3214);
nor U6196 (N_6196,N_4971,N_3826);
or U6197 (N_6197,N_3643,N_3972);
and U6198 (N_6198,N_4383,N_3619);
or U6199 (N_6199,N_2990,N_4945);
nand U6200 (N_6200,N_3152,N_4769);
nand U6201 (N_6201,N_4970,N_3736);
nor U6202 (N_6202,N_3581,N_3093);
nand U6203 (N_6203,N_3606,N_3501);
nand U6204 (N_6204,N_3034,N_3290);
and U6205 (N_6205,N_4553,N_4030);
nand U6206 (N_6206,N_4787,N_3419);
and U6207 (N_6207,N_3442,N_4780);
nand U6208 (N_6208,N_4210,N_3137);
or U6209 (N_6209,N_4785,N_3339);
and U6210 (N_6210,N_3390,N_4082);
xor U6211 (N_6211,N_3899,N_3040);
nand U6212 (N_6212,N_2980,N_4283);
nor U6213 (N_6213,N_2898,N_3648);
and U6214 (N_6214,N_2531,N_4822);
or U6215 (N_6215,N_3567,N_3397);
nand U6216 (N_6216,N_3967,N_2503);
xor U6217 (N_6217,N_3042,N_4808);
and U6218 (N_6218,N_4505,N_3177);
or U6219 (N_6219,N_4555,N_4353);
and U6220 (N_6220,N_3534,N_3735);
nand U6221 (N_6221,N_3458,N_4716);
nor U6222 (N_6222,N_3474,N_4329);
nor U6223 (N_6223,N_4999,N_3696);
or U6224 (N_6224,N_4479,N_4663);
nor U6225 (N_6225,N_2791,N_4681);
nor U6226 (N_6226,N_3465,N_3169);
nand U6227 (N_6227,N_3118,N_2954);
nand U6228 (N_6228,N_4515,N_2719);
nor U6229 (N_6229,N_3980,N_2783);
nand U6230 (N_6230,N_4763,N_3309);
nor U6231 (N_6231,N_3485,N_4817);
nor U6232 (N_6232,N_2698,N_2976);
nor U6233 (N_6233,N_4106,N_2828);
and U6234 (N_6234,N_2906,N_4672);
nor U6235 (N_6235,N_2518,N_3630);
nand U6236 (N_6236,N_4620,N_2626);
nor U6237 (N_6237,N_3564,N_4996);
xor U6238 (N_6238,N_4749,N_3524);
nor U6239 (N_6239,N_3031,N_3985);
or U6240 (N_6240,N_2539,N_4041);
or U6241 (N_6241,N_3357,N_3962);
or U6242 (N_6242,N_4754,N_2841);
and U6243 (N_6243,N_3467,N_3845);
or U6244 (N_6244,N_3211,N_2545);
or U6245 (N_6245,N_4033,N_2857);
nor U6246 (N_6246,N_2588,N_3885);
nand U6247 (N_6247,N_3616,N_3156);
and U6248 (N_6248,N_3297,N_4922);
nand U6249 (N_6249,N_4742,N_4918);
or U6250 (N_6250,N_2593,N_4952);
nand U6251 (N_6251,N_4005,N_3230);
and U6252 (N_6252,N_4215,N_4155);
or U6253 (N_6253,N_3672,N_3635);
nor U6254 (N_6254,N_4669,N_4665);
nand U6255 (N_6255,N_4408,N_3926);
nor U6256 (N_6256,N_4543,N_3519);
and U6257 (N_6257,N_4945,N_4630);
nand U6258 (N_6258,N_3605,N_4864);
nor U6259 (N_6259,N_4653,N_3687);
nor U6260 (N_6260,N_4180,N_3434);
nor U6261 (N_6261,N_3037,N_2570);
and U6262 (N_6262,N_4910,N_4273);
and U6263 (N_6263,N_2527,N_4106);
or U6264 (N_6264,N_4935,N_4927);
and U6265 (N_6265,N_2678,N_3128);
nand U6266 (N_6266,N_4722,N_3163);
and U6267 (N_6267,N_4452,N_3258);
nand U6268 (N_6268,N_4064,N_2918);
or U6269 (N_6269,N_3336,N_4551);
or U6270 (N_6270,N_3560,N_3518);
nor U6271 (N_6271,N_3740,N_4693);
nand U6272 (N_6272,N_2507,N_3342);
or U6273 (N_6273,N_3546,N_2537);
or U6274 (N_6274,N_4755,N_3735);
nor U6275 (N_6275,N_4342,N_4812);
nand U6276 (N_6276,N_4074,N_2810);
or U6277 (N_6277,N_2947,N_4455);
and U6278 (N_6278,N_2538,N_2961);
and U6279 (N_6279,N_4273,N_4098);
or U6280 (N_6280,N_3309,N_2926);
nand U6281 (N_6281,N_4020,N_3155);
nor U6282 (N_6282,N_3831,N_3537);
or U6283 (N_6283,N_4810,N_4853);
or U6284 (N_6284,N_4901,N_3207);
and U6285 (N_6285,N_4391,N_4540);
nand U6286 (N_6286,N_2595,N_4185);
and U6287 (N_6287,N_4956,N_2718);
nor U6288 (N_6288,N_2736,N_4861);
and U6289 (N_6289,N_3862,N_3346);
or U6290 (N_6290,N_3461,N_4239);
and U6291 (N_6291,N_2751,N_3706);
or U6292 (N_6292,N_4337,N_2503);
nand U6293 (N_6293,N_3211,N_3049);
and U6294 (N_6294,N_3262,N_3541);
and U6295 (N_6295,N_4562,N_3456);
nand U6296 (N_6296,N_4449,N_3237);
or U6297 (N_6297,N_4843,N_4333);
or U6298 (N_6298,N_3204,N_3219);
nor U6299 (N_6299,N_4764,N_2536);
nor U6300 (N_6300,N_3018,N_2742);
or U6301 (N_6301,N_3795,N_4894);
and U6302 (N_6302,N_3188,N_2905);
or U6303 (N_6303,N_2996,N_3392);
or U6304 (N_6304,N_3104,N_3713);
and U6305 (N_6305,N_2905,N_3771);
and U6306 (N_6306,N_2746,N_4205);
nand U6307 (N_6307,N_3949,N_2697);
nor U6308 (N_6308,N_3197,N_3811);
nand U6309 (N_6309,N_3923,N_3551);
and U6310 (N_6310,N_4583,N_3266);
nor U6311 (N_6311,N_2523,N_3043);
nor U6312 (N_6312,N_3030,N_2566);
and U6313 (N_6313,N_3680,N_4052);
nor U6314 (N_6314,N_4088,N_3780);
or U6315 (N_6315,N_2557,N_4181);
nor U6316 (N_6316,N_4010,N_4468);
nand U6317 (N_6317,N_3197,N_4575);
nor U6318 (N_6318,N_3457,N_2873);
xnor U6319 (N_6319,N_2938,N_3987);
and U6320 (N_6320,N_3854,N_2535);
nor U6321 (N_6321,N_3542,N_3212);
nor U6322 (N_6322,N_2858,N_2771);
nand U6323 (N_6323,N_2815,N_3832);
nor U6324 (N_6324,N_3683,N_2903);
nor U6325 (N_6325,N_4023,N_3337);
and U6326 (N_6326,N_2982,N_3153);
and U6327 (N_6327,N_2990,N_3936);
nor U6328 (N_6328,N_3163,N_2938);
nor U6329 (N_6329,N_2852,N_3617);
nand U6330 (N_6330,N_4800,N_3033);
nor U6331 (N_6331,N_3883,N_2777);
nor U6332 (N_6332,N_2558,N_4382);
or U6333 (N_6333,N_4419,N_4970);
nand U6334 (N_6334,N_3888,N_3639);
and U6335 (N_6335,N_2549,N_4901);
nand U6336 (N_6336,N_3688,N_2506);
and U6337 (N_6337,N_3632,N_3812);
or U6338 (N_6338,N_2888,N_3197);
or U6339 (N_6339,N_3387,N_2569);
nand U6340 (N_6340,N_3079,N_3500);
and U6341 (N_6341,N_2566,N_2948);
nor U6342 (N_6342,N_3408,N_4214);
or U6343 (N_6343,N_2577,N_4305);
xor U6344 (N_6344,N_3960,N_4998);
nor U6345 (N_6345,N_4382,N_4461);
and U6346 (N_6346,N_3142,N_4283);
or U6347 (N_6347,N_3929,N_2985);
or U6348 (N_6348,N_4919,N_4064);
and U6349 (N_6349,N_3820,N_4342);
or U6350 (N_6350,N_4875,N_4888);
nand U6351 (N_6351,N_3751,N_2890);
nor U6352 (N_6352,N_2775,N_3388);
nor U6353 (N_6353,N_2678,N_2544);
nand U6354 (N_6354,N_4331,N_2556);
or U6355 (N_6355,N_4977,N_4473);
or U6356 (N_6356,N_4158,N_4864);
or U6357 (N_6357,N_4065,N_4974);
and U6358 (N_6358,N_3709,N_2573);
nor U6359 (N_6359,N_3470,N_4444);
and U6360 (N_6360,N_4904,N_4085);
or U6361 (N_6361,N_4557,N_4662);
nand U6362 (N_6362,N_4634,N_3534);
nand U6363 (N_6363,N_2738,N_4120);
nor U6364 (N_6364,N_4422,N_3358);
and U6365 (N_6365,N_4694,N_3038);
or U6366 (N_6366,N_3461,N_3520);
or U6367 (N_6367,N_4483,N_3647);
nor U6368 (N_6368,N_4022,N_4518);
and U6369 (N_6369,N_3658,N_3240);
nand U6370 (N_6370,N_2722,N_4127);
nand U6371 (N_6371,N_3985,N_3260);
or U6372 (N_6372,N_3497,N_3566);
or U6373 (N_6373,N_4699,N_4168);
nor U6374 (N_6374,N_3798,N_4773);
nor U6375 (N_6375,N_3397,N_4993);
or U6376 (N_6376,N_2867,N_3061);
nand U6377 (N_6377,N_3228,N_3880);
nor U6378 (N_6378,N_3446,N_3029);
nor U6379 (N_6379,N_3714,N_3164);
and U6380 (N_6380,N_3604,N_3416);
nor U6381 (N_6381,N_2754,N_3742);
nand U6382 (N_6382,N_2775,N_4398);
or U6383 (N_6383,N_3764,N_4484);
and U6384 (N_6384,N_3245,N_4482);
nand U6385 (N_6385,N_3084,N_3485);
nand U6386 (N_6386,N_4736,N_3875);
and U6387 (N_6387,N_3856,N_4910);
or U6388 (N_6388,N_2689,N_3018);
nand U6389 (N_6389,N_2656,N_3463);
nor U6390 (N_6390,N_2610,N_3958);
and U6391 (N_6391,N_3214,N_4062);
and U6392 (N_6392,N_3015,N_4831);
and U6393 (N_6393,N_4131,N_4558);
and U6394 (N_6394,N_3387,N_3180);
nor U6395 (N_6395,N_3137,N_3129);
or U6396 (N_6396,N_4475,N_3087);
nor U6397 (N_6397,N_3313,N_3875);
nor U6398 (N_6398,N_2708,N_2915);
nand U6399 (N_6399,N_4388,N_4153);
or U6400 (N_6400,N_3741,N_3666);
or U6401 (N_6401,N_3251,N_4837);
and U6402 (N_6402,N_4015,N_2779);
and U6403 (N_6403,N_4586,N_3202);
nor U6404 (N_6404,N_4453,N_4342);
or U6405 (N_6405,N_2937,N_4925);
and U6406 (N_6406,N_2613,N_4140);
and U6407 (N_6407,N_3122,N_3113);
nand U6408 (N_6408,N_2865,N_4868);
or U6409 (N_6409,N_3214,N_2825);
nor U6410 (N_6410,N_2609,N_4115);
nand U6411 (N_6411,N_4587,N_4504);
nand U6412 (N_6412,N_3093,N_3403);
or U6413 (N_6413,N_4311,N_4946);
nor U6414 (N_6414,N_2896,N_4291);
nand U6415 (N_6415,N_4672,N_4215);
or U6416 (N_6416,N_4236,N_4808);
or U6417 (N_6417,N_3954,N_2629);
and U6418 (N_6418,N_3919,N_2669);
or U6419 (N_6419,N_4617,N_3129);
nor U6420 (N_6420,N_4805,N_4810);
and U6421 (N_6421,N_3112,N_4762);
or U6422 (N_6422,N_3393,N_3087);
nand U6423 (N_6423,N_2839,N_2595);
nand U6424 (N_6424,N_2667,N_3455);
and U6425 (N_6425,N_3645,N_2626);
or U6426 (N_6426,N_4080,N_3834);
or U6427 (N_6427,N_3683,N_3266);
nor U6428 (N_6428,N_2555,N_4765);
or U6429 (N_6429,N_3839,N_4214);
and U6430 (N_6430,N_3095,N_3295);
and U6431 (N_6431,N_3895,N_4575);
or U6432 (N_6432,N_2654,N_4885);
nor U6433 (N_6433,N_2624,N_3463);
nor U6434 (N_6434,N_2977,N_2649);
nor U6435 (N_6435,N_4609,N_4903);
or U6436 (N_6436,N_2994,N_3761);
nor U6437 (N_6437,N_3198,N_4772);
or U6438 (N_6438,N_4713,N_4717);
and U6439 (N_6439,N_4763,N_3726);
nor U6440 (N_6440,N_4971,N_4141);
nand U6441 (N_6441,N_4306,N_3958);
and U6442 (N_6442,N_3501,N_2808);
nand U6443 (N_6443,N_3776,N_4353);
nand U6444 (N_6444,N_2646,N_4644);
or U6445 (N_6445,N_4006,N_4113);
nor U6446 (N_6446,N_3649,N_3521);
nor U6447 (N_6447,N_2696,N_4905);
nor U6448 (N_6448,N_3519,N_2736);
or U6449 (N_6449,N_4562,N_3389);
nor U6450 (N_6450,N_3550,N_4317);
or U6451 (N_6451,N_4233,N_3336);
nor U6452 (N_6452,N_4421,N_4602);
or U6453 (N_6453,N_3792,N_4441);
nand U6454 (N_6454,N_3634,N_4003);
nand U6455 (N_6455,N_4754,N_3971);
and U6456 (N_6456,N_3778,N_4715);
nand U6457 (N_6457,N_4857,N_4281);
nor U6458 (N_6458,N_4163,N_3804);
and U6459 (N_6459,N_2869,N_3989);
and U6460 (N_6460,N_4205,N_4281);
and U6461 (N_6461,N_4736,N_3748);
nor U6462 (N_6462,N_4863,N_3029);
and U6463 (N_6463,N_2778,N_4827);
nand U6464 (N_6464,N_3919,N_2916);
or U6465 (N_6465,N_3078,N_4743);
or U6466 (N_6466,N_4091,N_4452);
or U6467 (N_6467,N_3503,N_3842);
xnor U6468 (N_6468,N_3222,N_2983);
nand U6469 (N_6469,N_4492,N_4754);
or U6470 (N_6470,N_2612,N_4108);
nor U6471 (N_6471,N_2597,N_4712);
nand U6472 (N_6472,N_3041,N_4697);
and U6473 (N_6473,N_4463,N_2756);
nor U6474 (N_6474,N_3677,N_4256);
or U6475 (N_6475,N_4895,N_4220);
nand U6476 (N_6476,N_2887,N_3688);
or U6477 (N_6477,N_2563,N_4373);
and U6478 (N_6478,N_2673,N_2765);
or U6479 (N_6479,N_4066,N_3062);
nor U6480 (N_6480,N_4919,N_3262);
and U6481 (N_6481,N_2986,N_3373);
nand U6482 (N_6482,N_4320,N_3098);
or U6483 (N_6483,N_4079,N_3401);
nand U6484 (N_6484,N_2723,N_4847);
and U6485 (N_6485,N_3263,N_3219);
nor U6486 (N_6486,N_2502,N_4163);
or U6487 (N_6487,N_3476,N_3861);
or U6488 (N_6488,N_4406,N_3215);
and U6489 (N_6489,N_2515,N_3859);
nand U6490 (N_6490,N_4449,N_3334);
or U6491 (N_6491,N_2981,N_2754);
or U6492 (N_6492,N_3783,N_2500);
and U6493 (N_6493,N_2521,N_4538);
and U6494 (N_6494,N_2530,N_4408);
and U6495 (N_6495,N_3930,N_4029);
or U6496 (N_6496,N_2775,N_3954);
xnor U6497 (N_6497,N_3633,N_4716);
nor U6498 (N_6498,N_4535,N_4132);
and U6499 (N_6499,N_2641,N_3436);
nor U6500 (N_6500,N_3300,N_3439);
nor U6501 (N_6501,N_4326,N_2714);
nor U6502 (N_6502,N_3052,N_3043);
nand U6503 (N_6503,N_3753,N_3742);
nor U6504 (N_6504,N_3552,N_4417);
or U6505 (N_6505,N_3390,N_3637);
or U6506 (N_6506,N_2960,N_4325);
nand U6507 (N_6507,N_2705,N_2589);
or U6508 (N_6508,N_2916,N_4275);
nor U6509 (N_6509,N_2510,N_2911);
and U6510 (N_6510,N_3220,N_4916);
nand U6511 (N_6511,N_2536,N_3334);
or U6512 (N_6512,N_4796,N_3752);
or U6513 (N_6513,N_4670,N_3357);
and U6514 (N_6514,N_4021,N_2833);
nor U6515 (N_6515,N_4301,N_3669);
and U6516 (N_6516,N_4331,N_2912);
nand U6517 (N_6517,N_3310,N_3315);
or U6518 (N_6518,N_3223,N_3713);
nand U6519 (N_6519,N_4877,N_3188);
and U6520 (N_6520,N_4344,N_2955);
and U6521 (N_6521,N_3594,N_2800);
or U6522 (N_6522,N_4633,N_3787);
nor U6523 (N_6523,N_2609,N_4815);
nor U6524 (N_6524,N_4699,N_4314);
and U6525 (N_6525,N_4409,N_4652);
nand U6526 (N_6526,N_4516,N_3923);
or U6527 (N_6527,N_4083,N_4529);
nor U6528 (N_6528,N_3118,N_4670);
or U6529 (N_6529,N_4463,N_4021);
or U6530 (N_6530,N_3705,N_2826);
nand U6531 (N_6531,N_2697,N_4904);
nor U6532 (N_6532,N_2538,N_4363);
nand U6533 (N_6533,N_3830,N_3642);
nor U6534 (N_6534,N_2921,N_3141);
and U6535 (N_6535,N_3567,N_3058);
nor U6536 (N_6536,N_4930,N_4759);
and U6537 (N_6537,N_2547,N_3631);
nand U6538 (N_6538,N_2905,N_3395);
nand U6539 (N_6539,N_4537,N_3031);
or U6540 (N_6540,N_4818,N_4482);
or U6541 (N_6541,N_3785,N_4435);
nand U6542 (N_6542,N_3202,N_4926);
nand U6543 (N_6543,N_3040,N_2571);
nand U6544 (N_6544,N_2571,N_3831);
or U6545 (N_6545,N_3542,N_4193);
and U6546 (N_6546,N_2972,N_4945);
and U6547 (N_6547,N_4685,N_4427);
nand U6548 (N_6548,N_4569,N_2905);
nand U6549 (N_6549,N_3335,N_3910);
and U6550 (N_6550,N_4322,N_4142);
nand U6551 (N_6551,N_4082,N_4619);
and U6552 (N_6552,N_4244,N_3157);
and U6553 (N_6553,N_3257,N_3688);
nor U6554 (N_6554,N_3702,N_3276);
nor U6555 (N_6555,N_3616,N_2511);
or U6556 (N_6556,N_2929,N_2971);
and U6557 (N_6557,N_4339,N_3704);
or U6558 (N_6558,N_2640,N_4629);
nand U6559 (N_6559,N_3404,N_2730);
nand U6560 (N_6560,N_3456,N_4864);
nand U6561 (N_6561,N_4807,N_4912);
nand U6562 (N_6562,N_3106,N_2732);
nor U6563 (N_6563,N_4074,N_3460);
or U6564 (N_6564,N_2644,N_3206);
or U6565 (N_6565,N_4525,N_4251);
nand U6566 (N_6566,N_4991,N_4493);
nand U6567 (N_6567,N_2879,N_3052);
and U6568 (N_6568,N_2738,N_4335);
nor U6569 (N_6569,N_2532,N_4125);
and U6570 (N_6570,N_2951,N_4890);
or U6571 (N_6571,N_4033,N_4501);
nand U6572 (N_6572,N_4653,N_2844);
nand U6573 (N_6573,N_3870,N_4050);
or U6574 (N_6574,N_4728,N_3455);
nand U6575 (N_6575,N_3335,N_4156);
nand U6576 (N_6576,N_3717,N_4250);
and U6577 (N_6577,N_3726,N_3434);
or U6578 (N_6578,N_2863,N_2604);
or U6579 (N_6579,N_3691,N_4647);
nor U6580 (N_6580,N_3545,N_4903);
nor U6581 (N_6581,N_4819,N_4334);
and U6582 (N_6582,N_3246,N_3093);
nor U6583 (N_6583,N_4535,N_3178);
or U6584 (N_6584,N_4946,N_3015);
nand U6585 (N_6585,N_2934,N_4861);
and U6586 (N_6586,N_4632,N_4621);
or U6587 (N_6587,N_4277,N_2714);
and U6588 (N_6588,N_2624,N_4048);
nand U6589 (N_6589,N_4835,N_3208);
nor U6590 (N_6590,N_2651,N_4786);
nand U6591 (N_6591,N_3682,N_4704);
nand U6592 (N_6592,N_3563,N_2721);
nor U6593 (N_6593,N_4039,N_3336);
nand U6594 (N_6594,N_2768,N_3541);
or U6595 (N_6595,N_3431,N_3193);
nand U6596 (N_6596,N_4067,N_2727);
xnor U6597 (N_6597,N_2633,N_3777);
and U6598 (N_6598,N_4816,N_3435);
or U6599 (N_6599,N_2963,N_4328);
or U6600 (N_6600,N_2652,N_3457);
and U6601 (N_6601,N_4034,N_2854);
or U6602 (N_6602,N_4688,N_3511);
nor U6603 (N_6603,N_2713,N_2698);
and U6604 (N_6604,N_3243,N_4639);
and U6605 (N_6605,N_3819,N_4693);
and U6606 (N_6606,N_4562,N_4829);
nor U6607 (N_6607,N_3266,N_4864);
nor U6608 (N_6608,N_3057,N_2558);
or U6609 (N_6609,N_2941,N_3672);
and U6610 (N_6610,N_4556,N_3849);
or U6611 (N_6611,N_2849,N_2966);
or U6612 (N_6612,N_4406,N_2958);
nand U6613 (N_6613,N_4647,N_2606);
nand U6614 (N_6614,N_3579,N_3815);
and U6615 (N_6615,N_3893,N_4911);
and U6616 (N_6616,N_4196,N_2920);
nor U6617 (N_6617,N_2551,N_3218);
nor U6618 (N_6618,N_3582,N_3209);
or U6619 (N_6619,N_4374,N_4606);
nand U6620 (N_6620,N_4798,N_3465);
nand U6621 (N_6621,N_4530,N_4717);
or U6622 (N_6622,N_4652,N_2654);
or U6623 (N_6623,N_3777,N_4220);
and U6624 (N_6624,N_4384,N_3976);
or U6625 (N_6625,N_4419,N_2543);
and U6626 (N_6626,N_4243,N_3494);
or U6627 (N_6627,N_4514,N_3130);
nand U6628 (N_6628,N_3234,N_4874);
nand U6629 (N_6629,N_4963,N_4378);
or U6630 (N_6630,N_4752,N_4356);
nand U6631 (N_6631,N_3692,N_4869);
nand U6632 (N_6632,N_3935,N_2970);
xor U6633 (N_6633,N_2815,N_4091);
nor U6634 (N_6634,N_3663,N_3582);
nor U6635 (N_6635,N_4921,N_3656);
or U6636 (N_6636,N_4004,N_3494);
nand U6637 (N_6637,N_2912,N_4535);
nor U6638 (N_6638,N_4407,N_2807);
and U6639 (N_6639,N_3724,N_2663);
nor U6640 (N_6640,N_3985,N_3440);
nand U6641 (N_6641,N_3604,N_4102);
and U6642 (N_6642,N_3626,N_4380);
nor U6643 (N_6643,N_3612,N_2843);
xnor U6644 (N_6644,N_3515,N_2911);
or U6645 (N_6645,N_4002,N_4292);
nor U6646 (N_6646,N_2764,N_2854);
nand U6647 (N_6647,N_4132,N_3929);
or U6648 (N_6648,N_2998,N_3294);
and U6649 (N_6649,N_4458,N_4345);
nand U6650 (N_6650,N_3553,N_4065);
or U6651 (N_6651,N_2606,N_3254);
or U6652 (N_6652,N_3172,N_3736);
or U6653 (N_6653,N_3614,N_4265);
nand U6654 (N_6654,N_2653,N_3928);
nand U6655 (N_6655,N_4002,N_3058);
or U6656 (N_6656,N_4760,N_2999);
or U6657 (N_6657,N_3050,N_4393);
or U6658 (N_6658,N_3526,N_3720);
and U6659 (N_6659,N_4441,N_2614);
or U6660 (N_6660,N_4647,N_4101);
and U6661 (N_6661,N_3115,N_3524);
nand U6662 (N_6662,N_3937,N_3602);
or U6663 (N_6663,N_4722,N_2878);
and U6664 (N_6664,N_4675,N_4782);
nand U6665 (N_6665,N_3418,N_4775);
and U6666 (N_6666,N_4341,N_4535);
nand U6667 (N_6667,N_4024,N_4643);
and U6668 (N_6668,N_3874,N_3248);
and U6669 (N_6669,N_4827,N_4274);
or U6670 (N_6670,N_2928,N_3020);
nor U6671 (N_6671,N_2952,N_4141);
nand U6672 (N_6672,N_3569,N_3454);
or U6673 (N_6673,N_3825,N_2583);
nand U6674 (N_6674,N_3336,N_4900);
nand U6675 (N_6675,N_3288,N_4247);
nor U6676 (N_6676,N_3720,N_3015);
and U6677 (N_6677,N_4645,N_4328);
or U6678 (N_6678,N_3500,N_4359);
nor U6679 (N_6679,N_3612,N_3324);
or U6680 (N_6680,N_4285,N_4040);
or U6681 (N_6681,N_3820,N_4602);
nor U6682 (N_6682,N_2632,N_3526);
or U6683 (N_6683,N_4807,N_4940);
nor U6684 (N_6684,N_4437,N_4656);
nor U6685 (N_6685,N_2698,N_2899);
nor U6686 (N_6686,N_4151,N_4544);
or U6687 (N_6687,N_3088,N_4172);
nand U6688 (N_6688,N_3285,N_4741);
nor U6689 (N_6689,N_2936,N_4916);
or U6690 (N_6690,N_4971,N_4080);
nor U6691 (N_6691,N_4358,N_3576);
nand U6692 (N_6692,N_4015,N_4461);
and U6693 (N_6693,N_3399,N_3654);
nand U6694 (N_6694,N_3270,N_3874);
nor U6695 (N_6695,N_3319,N_3317);
nor U6696 (N_6696,N_4334,N_4580);
nor U6697 (N_6697,N_2790,N_3171);
nand U6698 (N_6698,N_2611,N_3575);
and U6699 (N_6699,N_3729,N_4699);
and U6700 (N_6700,N_2592,N_2559);
nor U6701 (N_6701,N_2650,N_4782);
nand U6702 (N_6702,N_4949,N_4109);
and U6703 (N_6703,N_2571,N_3542);
or U6704 (N_6704,N_3815,N_2717);
nand U6705 (N_6705,N_4319,N_4573);
nand U6706 (N_6706,N_2569,N_4358);
and U6707 (N_6707,N_3749,N_4080);
nand U6708 (N_6708,N_4122,N_4575);
xor U6709 (N_6709,N_4776,N_2794);
or U6710 (N_6710,N_4204,N_2813);
or U6711 (N_6711,N_3007,N_2864);
or U6712 (N_6712,N_3169,N_4769);
and U6713 (N_6713,N_3648,N_4042);
nand U6714 (N_6714,N_4155,N_3689);
and U6715 (N_6715,N_4243,N_4398);
nand U6716 (N_6716,N_4285,N_3210);
or U6717 (N_6717,N_4558,N_3901);
nand U6718 (N_6718,N_2942,N_4477);
or U6719 (N_6719,N_3361,N_2747);
and U6720 (N_6720,N_4092,N_4171);
nand U6721 (N_6721,N_3246,N_4076);
and U6722 (N_6722,N_4352,N_4086);
nor U6723 (N_6723,N_4669,N_3510);
nor U6724 (N_6724,N_4395,N_3219);
and U6725 (N_6725,N_4313,N_2939);
and U6726 (N_6726,N_3918,N_3437);
nor U6727 (N_6727,N_3928,N_3915);
nand U6728 (N_6728,N_3692,N_4818);
and U6729 (N_6729,N_3484,N_3412);
and U6730 (N_6730,N_3950,N_4146);
nand U6731 (N_6731,N_4588,N_3337);
nor U6732 (N_6732,N_3258,N_4721);
nor U6733 (N_6733,N_2641,N_3825);
nand U6734 (N_6734,N_2603,N_2664);
and U6735 (N_6735,N_3302,N_3229);
and U6736 (N_6736,N_3693,N_4687);
nor U6737 (N_6737,N_3880,N_3955);
nor U6738 (N_6738,N_3988,N_4905);
or U6739 (N_6739,N_3737,N_4221);
or U6740 (N_6740,N_4488,N_4244);
and U6741 (N_6741,N_4090,N_4348);
nand U6742 (N_6742,N_4248,N_3844);
nand U6743 (N_6743,N_2787,N_2935);
nand U6744 (N_6744,N_2829,N_3975);
nor U6745 (N_6745,N_4188,N_2998);
and U6746 (N_6746,N_4201,N_2748);
and U6747 (N_6747,N_4861,N_3832);
or U6748 (N_6748,N_3406,N_3554);
nand U6749 (N_6749,N_3958,N_3201);
or U6750 (N_6750,N_4507,N_3025);
or U6751 (N_6751,N_3912,N_2805);
or U6752 (N_6752,N_4471,N_4237);
nand U6753 (N_6753,N_3262,N_2761);
and U6754 (N_6754,N_4373,N_4832);
nand U6755 (N_6755,N_3099,N_3000);
xor U6756 (N_6756,N_3256,N_3617);
or U6757 (N_6757,N_4386,N_4427);
nand U6758 (N_6758,N_4826,N_3488);
or U6759 (N_6759,N_3218,N_4718);
nor U6760 (N_6760,N_4754,N_3206);
or U6761 (N_6761,N_4529,N_3182);
or U6762 (N_6762,N_4026,N_3345);
nor U6763 (N_6763,N_4490,N_3791);
nor U6764 (N_6764,N_4036,N_3068);
nor U6765 (N_6765,N_3903,N_3298);
or U6766 (N_6766,N_4964,N_3876);
and U6767 (N_6767,N_4675,N_3976);
nor U6768 (N_6768,N_2898,N_4846);
nor U6769 (N_6769,N_2509,N_3194);
and U6770 (N_6770,N_4856,N_2669);
nand U6771 (N_6771,N_3938,N_4299);
nand U6772 (N_6772,N_3796,N_4346);
nor U6773 (N_6773,N_3082,N_4142);
nand U6774 (N_6774,N_2620,N_2530);
nand U6775 (N_6775,N_3578,N_4875);
nand U6776 (N_6776,N_2942,N_4299);
nor U6777 (N_6777,N_3693,N_4095);
and U6778 (N_6778,N_3280,N_4927);
nor U6779 (N_6779,N_4724,N_3236);
or U6780 (N_6780,N_4231,N_3439);
or U6781 (N_6781,N_3396,N_4849);
or U6782 (N_6782,N_4558,N_3125);
or U6783 (N_6783,N_4066,N_2540);
and U6784 (N_6784,N_3553,N_3675);
and U6785 (N_6785,N_4573,N_4417);
and U6786 (N_6786,N_2751,N_4025);
or U6787 (N_6787,N_4839,N_2573);
or U6788 (N_6788,N_3715,N_4775);
nor U6789 (N_6789,N_2627,N_3924);
and U6790 (N_6790,N_2713,N_2805);
nand U6791 (N_6791,N_4979,N_4981);
and U6792 (N_6792,N_3642,N_4839);
nand U6793 (N_6793,N_3238,N_2585);
nand U6794 (N_6794,N_3013,N_3763);
and U6795 (N_6795,N_3089,N_3952);
nor U6796 (N_6796,N_4001,N_4118);
or U6797 (N_6797,N_3813,N_3752);
nand U6798 (N_6798,N_2949,N_3128);
nand U6799 (N_6799,N_4861,N_2718);
nand U6800 (N_6800,N_4110,N_2785);
nor U6801 (N_6801,N_2932,N_3789);
nor U6802 (N_6802,N_3317,N_2721);
nand U6803 (N_6803,N_4768,N_2927);
nand U6804 (N_6804,N_3152,N_3196);
nand U6805 (N_6805,N_4938,N_3837);
nor U6806 (N_6806,N_4561,N_4886);
and U6807 (N_6807,N_2588,N_4587);
nor U6808 (N_6808,N_2855,N_3280);
nor U6809 (N_6809,N_2748,N_2732);
and U6810 (N_6810,N_2739,N_3341);
and U6811 (N_6811,N_4279,N_4620);
nor U6812 (N_6812,N_4131,N_3897);
nor U6813 (N_6813,N_4235,N_3749);
nand U6814 (N_6814,N_4483,N_4120);
and U6815 (N_6815,N_4654,N_2789);
nand U6816 (N_6816,N_3688,N_4826);
and U6817 (N_6817,N_4905,N_3818);
or U6818 (N_6818,N_4287,N_4158);
or U6819 (N_6819,N_3606,N_3279);
and U6820 (N_6820,N_3463,N_3884);
nand U6821 (N_6821,N_4590,N_4257);
or U6822 (N_6822,N_3765,N_2914);
nor U6823 (N_6823,N_3941,N_3733);
nand U6824 (N_6824,N_2507,N_3114);
or U6825 (N_6825,N_4136,N_4198);
nand U6826 (N_6826,N_4015,N_4119);
nand U6827 (N_6827,N_3281,N_4370);
nor U6828 (N_6828,N_3878,N_3156);
and U6829 (N_6829,N_4009,N_3155);
nor U6830 (N_6830,N_4644,N_4154);
or U6831 (N_6831,N_3282,N_3009);
and U6832 (N_6832,N_4437,N_4356);
or U6833 (N_6833,N_4638,N_3130);
and U6834 (N_6834,N_3189,N_4620);
or U6835 (N_6835,N_2894,N_3710);
nor U6836 (N_6836,N_4705,N_2982);
nand U6837 (N_6837,N_2527,N_4185);
or U6838 (N_6838,N_4011,N_4731);
or U6839 (N_6839,N_3365,N_2855);
and U6840 (N_6840,N_3414,N_2594);
nand U6841 (N_6841,N_4858,N_4295);
or U6842 (N_6842,N_4838,N_4371);
nand U6843 (N_6843,N_3263,N_3152);
and U6844 (N_6844,N_2761,N_2621);
or U6845 (N_6845,N_3501,N_4255);
or U6846 (N_6846,N_4710,N_4351);
nor U6847 (N_6847,N_3133,N_4672);
and U6848 (N_6848,N_4010,N_2713);
or U6849 (N_6849,N_3601,N_2700);
and U6850 (N_6850,N_4575,N_2541);
nor U6851 (N_6851,N_3167,N_4909);
or U6852 (N_6852,N_4180,N_3336);
or U6853 (N_6853,N_3622,N_2543);
nand U6854 (N_6854,N_3882,N_4521);
nor U6855 (N_6855,N_2694,N_2644);
nand U6856 (N_6856,N_4336,N_4350);
and U6857 (N_6857,N_3987,N_3821);
nand U6858 (N_6858,N_3849,N_3301);
and U6859 (N_6859,N_4038,N_3594);
and U6860 (N_6860,N_4976,N_2888);
nand U6861 (N_6861,N_3408,N_4626);
nand U6862 (N_6862,N_4458,N_2592);
nand U6863 (N_6863,N_3421,N_4947);
nand U6864 (N_6864,N_2691,N_2733);
nand U6865 (N_6865,N_2697,N_4632);
or U6866 (N_6866,N_3018,N_3653);
and U6867 (N_6867,N_4846,N_4717);
or U6868 (N_6868,N_4601,N_2599);
nand U6869 (N_6869,N_2907,N_4221);
and U6870 (N_6870,N_3515,N_4657);
and U6871 (N_6871,N_3651,N_3275);
or U6872 (N_6872,N_4498,N_3241);
nor U6873 (N_6873,N_3046,N_3565);
nor U6874 (N_6874,N_3903,N_4962);
nand U6875 (N_6875,N_3907,N_4313);
nor U6876 (N_6876,N_4883,N_4043);
or U6877 (N_6877,N_4289,N_3773);
or U6878 (N_6878,N_2689,N_4909);
nand U6879 (N_6879,N_2690,N_3884);
or U6880 (N_6880,N_4364,N_4355);
nand U6881 (N_6881,N_3860,N_3758);
xnor U6882 (N_6882,N_4062,N_3421);
nor U6883 (N_6883,N_3713,N_4207);
or U6884 (N_6884,N_4087,N_4235);
or U6885 (N_6885,N_2884,N_4192);
nor U6886 (N_6886,N_2879,N_3896);
nand U6887 (N_6887,N_3708,N_4740);
nor U6888 (N_6888,N_3071,N_4457);
or U6889 (N_6889,N_2825,N_4380);
or U6890 (N_6890,N_4677,N_3235);
and U6891 (N_6891,N_4274,N_4957);
or U6892 (N_6892,N_4098,N_4686);
and U6893 (N_6893,N_4856,N_4456);
or U6894 (N_6894,N_2618,N_4039);
and U6895 (N_6895,N_4228,N_3988);
or U6896 (N_6896,N_4891,N_4844);
or U6897 (N_6897,N_2909,N_4371);
nor U6898 (N_6898,N_4343,N_3737);
nand U6899 (N_6899,N_2631,N_3763);
nand U6900 (N_6900,N_4667,N_2913);
and U6901 (N_6901,N_4813,N_4773);
nor U6902 (N_6902,N_4323,N_4774);
or U6903 (N_6903,N_3404,N_4182);
or U6904 (N_6904,N_3314,N_4548);
and U6905 (N_6905,N_2500,N_4977);
nand U6906 (N_6906,N_4408,N_4590);
or U6907 (N_6907,N_3359,N_3607);
and U6908 (N_6908,N_4107,N_3279);
nand U6909 (N_6909,N_4322,N_3971);
nand U6910 (N_6910,N_4383,N_3861);
and U6911 (N_6911,N_2866,N_3813);
and U6912 (N_6912,N_3121,N_4939);
and U6913 (N_6913,N_4907,N_2700);
nand U6914 (N_6914,N_2559,N_4567);
and U6915 (N_6915,N_2994,N_3299);
nand U6916 (N_6916,N_4284,N_4885);
and U6917 (N_6917,N_3859,N_4099);
and U6918 (N_6918,N_4909,N_2824);
or U6919 (N_6919,N_3309,N_2823);
xor U6920 (N_6920,N_3976,N_2552);
nor U6921 (N_6921,N_4670,N_3543);
nor U6922 (N_6922,N_3279,N_4254);
or U6923 (N_6923,N_2547,N_3430);
or U6924 (N_6924,N_4396,N_3907);
or U6925 (N_6925,N_2970,N_3899);
and U6926 (N_6926,N_4964,N_4042);
and U6927 (N_6927,N_3486,N_4694);
nor U6928 (N_6928,N_4419,N_3652);
and U6929 (N_6929,N_4880,N_4582);
nand U6930 (N_6930,N_4100,N_4883);
nor U6931 (N_6931,N_4844,N_2855);
or U6932 (N_6932,N_4920,N_4591);
or U6933 (N_6933,N_3054,N_4313);
nand U6934 (N_6934,N_4077,N_2600);
nor U6935 (N_6935,N_3158,N_2825);
nand U6936 (N_6936,N_3630,N_2796);
and U6937 (N_6937,N_4528,N_3162);
nand U6938 (N_6938,N_4910,N_4267);
nor U6939 (N_6939,N_4496,N_3320);
and U6940 (N_6940,N_2630,N_3998);
nor U6941 (N_6941,N_3192,N_3683);
nor U6942 (N_6942,N_2538,N_4807);
and U6943 (N_6943,N_3813,N_4140);
and U6944 (N_6944,N_3263,N_4168);
nor U6945 (N_6945,N_4975,N_2866);
and U6946 (N_6946,N_4573,N_4472);
nor U6947 (N_6947,N_2502,N_4674);
nor U6948 (N_6948,N_3187,N_2671);
and U6949 (N_6949,N_2741,N_2763);
nand U6950 (N_6950,N_2528,N_4578);
and U6951 (N_6951,N_2846,N_3569);
nand U6952 (N_6952,N_4966,N_2941);
nand U6953 (N_6953,N_4143,N_3060);
nand U6954 (N_6954,N_4594,N_4308);
nor U6955 (N_6955,N_4757,N_2746);
nor U6956 (N_6956,N_4938,N_4829);
and U6957 (N_6957,N_4773,N_3400);
and U6958 (N_6958,N_3853,N_4471);
or U6959 (N_6959,N_3279,N_2942);
or U6960 (N_6960,N_2802,N_3204);
nor U6961 (N_6961,N_2994,N_4259);
and U6962 (N_6962,N_3319,N_4900);
nor U6963 (N_6963,N_2805,N_2947);
or U6964 (N_6964,N_4686,N_2822);
and U6965 (N_6965,N_2983,N_4303);
nand U6966 (N_6966,N_4662,N_3541);
and U6967 (N_6967,N_4967,N_4345);
or U6968 (N_6968,N_4704,N_4200);
and U6969 (N_6969,N_2679,N_4942);
or U6970 (N_6970,N_4650,N_3980);
nor U6971 (N_6971,N_3448,N_4644);
or U6972 (N_6972,N_4102,N_2710);
nor U6973 (N_6973,N_4998,N_3499);
nor U6974 (N_6974,N_4530,N_4460);
nand U6975 (N_6975,N_4821,N_4917);
nand U6976 (N_6976,N_2558,N_4502);
nand U6977 (N_6977,N_3169,N_4990);
or U6978 (N_6978,N_4303,N_2772);
or U6979 (N_6979,N_2995,N_4476);
or U6980 (N_6980,N_2659,N_3523);
or U6981 (N_6981,N_3230,N_3724);
nand U6982 (N_6982,N_4258,N_2928);
and U6983 (N_6983,N_4071,N_3962);
or U6984 (N_6984,N_4625,N_4614);
nand U6985 (N_6985,N_4953,N_4901);
nor U6986 (N_6986,N_2677,N_2685);
nand U6987 (N_6987,N_3128,N_2560);
nand U6988 (N_6988,N_4171,N_3844);
nand U6989 (N_6989,N_4714,N_3127);
and U6990 (N_6990,N_2711,N_3653);
nor U6991 (N_6991,N_3488,N_4135);
and U6992 (N_6992,N_4948,N_2621);
nand U6993 (N_6993,N_4909,N_4543);
and U6994 (N_6994,N_3420,N_3677);
nand U6995 (N_6995,N_4036,N_3876);
and U6996 (N_6996,N_4896,N_4608);
or U6997 (N_6997,N_2936,N_2990);
nand U6998 (N_6998,N_4836,N_4277);
nand U6999 (N_6999,N_4200,N_4360);
nand U7000 (N_7000,N_4581,N_4543);
nor U7001 (N_7001,N_3979,N_2527);
nand U7002 (N_7002,N_3709,N_3154);
nand U7003 (N_7003,N_2806,N_3001);
and U7004 (N_7004,N_4394,N_3655);
nor U7005 (N_7005,N_3055,N_3116);
nor U7006 (N_7006,N_4308,N_4528);
and U7007 (N_7007,N_4030,N_3812);
or U7008 (N_7008,N_2994,N_2646);
or U7009 (N_7009,N_4888,N_4893);
nor U7010 (N_7010,N_3099,N_3622);
nand U7011 (N_7011,N_2973,N_4044);
or U7012 (N_7012,N_3477,N_3997);
nand U7013 (N_7013,N_3006,N_4881);
and U7014 (N_7014,N_4518,N_4377);
or U7015 (N_7015,N_4737,N_4783);
or U7016 (N_7016,N_3822,N_4349);
nand U7017 (N_7017,N_3912,N_4411);
nand U7018 (N_7018,N_3358,N_3591);
and U7019 (N_7019,N_4021,N_4426);
nand U7020 (N_7020,N_3215,N_4894);
nand U7021 (N_7021,N_3905,N_4252);
nor U7022 (N_7022,N_3555,N_4172);
or U7023 (N_7023,N_4235,N_2517);
nor U7024 (N_7024,N_4132,N_3203);
nor U7025 (N_7025,N_4112,N_2683);
and U7026 (N_7026,N_3548,N_3331);
nor U7027 (N_7027,N_3284,N_2728);
nor U7028 (N_7028,N_4939,N_3120);
and U7029 (N_7029,N_4949,N_3726);
and U7030 (N_7030,N_4471,N_4789);
and U7031 (N_7031,N_3662,N_4804);
or U7032 (N_7032,N_2947,N_3519);
nand U7033 (N_7033,N_4034,N_4905);
nor U7034 (N_7034,N_3842,N_4392);
and U7035 (N_7035,N_3544,N_3213);
nor U7036 (N_7036,N_4636,N_2978);
or U7037 (N_7037,N_3955,N_2702);
and U7038 (N_7038,N_3032,N_4080);
nor U7039 (N_7039,N_3269,N_4078);
nand U7040 (N_7040,N_4941,N_4940);
or U7041 (N_7041,N_3897,N_4620);
or U7042 (N_7042,N_2971,N_4434);
nand U7043 (N_7043,N_3832,N_3145);
nor U7044 (N_7044,N_3819,N_4896);
nand U7045 (N_7045,N_4739,N_3232);
and U7046 (N_7046,N_4455,N_4486);
nor U7047 (N_7047,N_2773,N_2831);
or U7048 (N_7048,N_3538,N_2985);
nand U7049 (N_7049,N_4285,N_4809);
and U7050 (N_7050,N_2913,N_4409);
or U7051 (N_7051,N_3506,N_3405);
or U7052 (N_7052,N_2737,N_4429);
nand U7053 (N_7053,N_4589,N_2549);
nor U7054 (N_7054,N_4222,N_3729);
nand U7055 (N_7055,N_4091,N_2641);
nand U7056 (N_7056,N_3778,N_2946);
nand U7057 (N_7057,N_4294,N_4083);
nand U7058 (N_7058,N_4203,N_4217);
or U7059 (N_7059,N_3688,N_4495);
nand U7060 (N_7060,N_3804,N_4625);
nand U7061 (N_7061,N_4448,N_3708);
nor U7062 (N_7062,N_4742,N_3161);
or U7063 (N_7063,N_2897,N_3690);
nand U7064 (N_7064,N_3922,N_2988);
or U7065 (N_7065,N_4309,N_3568);
nor U7066 (N_7066,N_3366,N_2930);
nand U7067 (N_7067,N_2984,N_2783);
nand U7068 (N_7068,N_4996,N_4859);
or U7069 (N_7069,N_3336,N_2553);
nand U7070 (N_7070,N_3026,N_4567);
or U7071 (N_7071,N_2634,N_3434);
nor U7072 (N_7072,N_4045,N_2922);
nor U7073 (N_7073,N_3283,N_4037);
or U7074 (N_7074,N_3381,N_4373);
or U7075 (N_7075,N_3561,N_4310);
nand U7076 (N_7076,N_3314,N_3371);
and U7077 (N_7077,N_4499,N_4872);
and U7078 (N_7078,N_4956,N_3029);
nand U7079 (N_7079,N_4034,N_4562);
nor U7080 (N_7080,N_4289,N_3547);
or U7081 (N_7081,N_4225,N_3294);
nor U7082 (N_7082,N_2888,N_2700);
nand U7083 (N_7083,N_4464,N_3589);
nor U7084 (N_7084,N_4909,N_4855);
and U7085 (N_7085,N_3533,N_4003);
nor U7086 (N_7086,N_4372,N_2763);
nand U7087 (N_7087,N_4067,N_3264);
and U7088 (N_7088,N_3812,N_3967);
nor U7089 (N_7089,N_2540,N_3850);
or U7090 (N_7090,N_4419,N_3045);
nand U7091 (N_7091,N_4267,N_4398);
nor U7092 (N_7092,N_3580,N_4428);
nor U7093 (N_7093,N_4230,N_4314);
nor U7094 (N_7094,N_3075,N_4172);
or U7095 (N_7095,N_3913,N_3692);
nand U7096 (N_7096,N_4712,N_2696);
and U7097 (N_7097,N_4903,N_3473);
and U7098 (N_7098,N_3052,N_4355);
nor U7099 (N_7099,N_3035,N_2676);
or U7100 (N_7100,N_3462,N_4712);
or U7101 (N_7101,N_3712,N_2709);
nand U7102 (N_7102,N_2777,N_4506);
or U7103 (N_7103,N_3274,N_2672);
nor U7104 (N_7104,N_4248,N_2755);
or U7105 (N_7105,N_3287,N_3582);
and U7106 (N_7106,N_3090,N_4669);
and U7107 (N_7107,N_4455,N_4249);
nor U7108 (N_7108,N_3116,N_3275);
nand U7109 (N_7109,N_3713,N_4776);
nand U7110 (N_7110,N_4286,N_3017);
and U7111 (N_7111,N_2770,N_3398);
and U7112 (N_7112,N_3958,N_3672);
nand U7113 (N_7113,N_2644,N_4964);
nand U7114 (N_7114,N_3896,N_3617);
nand U7115 (N_7115,N_4859,N_3557);
nor U7116 (N_7116,N_2858,N_2997);
and U7117 (N_7117,N_2664,N_3507);
or U7118 (N_7118,N_4799,N_4844);
nor U7119 (N_7119,N_2859,N_3172);
xnor U7120 (N_7120,N_2786,N_3083);
nand U7121 (N_7121,N_3950,N_2890);
or U7122 (N_7122,N_4596,N_2762);
and U7123 (N_7123,N_3867,N_3445);
and U7124 (N_7124,N_4764,N_4817);
or U7125 (N_7125,N_3359,N_4643);
and U7126 (N_7126,N_4725,N_3088);
and U7127 (N_7127,N_3318,N_3081);
and U7128 (N_7128,N_4741,N_4131);
nand U7129 (N_7129,N_4876,N_2572);
or U7130 (N_7130,N_3451,N_2934);
and U7131 (N_7131,N_3627,N_3445);
nor U7132 (N_7132,N_3942,N_3100);
and U7133 (N_7133,N_3923,N_4948);
nor U7134 (N_7134,N_4492,N_3412);
and U7135 (N_7135,N_3004,N_2595);
nor U7136 (N_7136,N_4882,N_4975);
or U7137 (N_7137,N_3902,N_3155);
or U7138 (N_7138,N_4502,N_3346);
or U7139 (N_7139,N_3676,N_4894);
or U7140 (N_7140,N_3585,N_4588);
nor U7141 (N_7141,N_2527,N_4411);
and U7142 (N_7142,N_3393,N_3283);
nand U7143 (N_7143,N_2955,N_4143);
or U7144 (N_7144,N_3617,N_3897);
nand U7145 (N_7145,N_3884,N_3738);
and U7146 (N_7146,N_3294,N_3531);
nand U7147 (N_7147,N_4093,N_4325);
or U7148 (N_7148,N_3020,N_2600);
or U7149 (N_7149,N_4603,N_2663);
nand U7150 (N_7150,N_4374,N_3510);
and U7151 (N_7151,N_2609,N_4502);
or U7152 (N_7152,N_3161,N_4649);
nand U7153 (N_7153,N_4015,N_2813);
nand U7154 (N_7154,N_2935,N_2851);
nor U7155 (N_7155,N_4268,N_2585);
nand U7156 (N_7156,N_4510,N_4305);
nand U7157 (N_7157,N_2858,N_2534);
nand U7158 (N_7158,N_4400,N_4395);
nand U7159 (N_7159,N_3621,N_3029);
or U7160 (N_7160,N_3336,N_3762);
and U7161 (N_7161,N_3680,N_4253);
and U7162 (N_7162,N_2845,N_3606);
nor U7163 (N_7163,N_4774,N_4882);
nand U7164 (N_7164,N_4298,N_4850);
nand U7165 (N_7165,N_3735,N_4884);
nand U7166 (N_7166,N_4184,N_2745);
and U7167 (N_7167,N_3373,N_4283);
and U7168 (N_7168,N_2633,N_4762);
nor U7169 (N_7169,N_2743,N_4033);
nand U7170 (N_7170,N_2598,N_4129);
nor U7171 (N_7171,N_4192,N_3271);
nor U7172 (N_7172,N_4208,N_2528);
nor U7173 (N_7173,N_2649,N_3330);
and U7174 (N_7174,N_3938,N_2774);
and U7175 (N_7175,N_4672,N_4587);
and U7176 (N_7176,N_4328,N_4331);
nand U7177 (N_7177,N_3773,N_4942);
nand U7178 (N_7178,N_4374,N_2745);
nand U7179 (N_7179,N_3466,N_4807);
and U7180 (N_7180,N_4580,N_4249);
nor U7181 (N_7181,N_4159,N_2872);
or U7182 (N_7182,N_3408,N_3294);
or U7183 (N_7183,N_4523,N_4531);
or U7184 (N_7184,N_2787,N_2849);
nor U7185 (N_7185,N_3504,N_4245);
or U7186 (N_7186,N_4032,N_4706);
or U7187 (N_7187,N_4290,N_4684);
or U7188 (N_7188,N_4467,N_4681);
or U7189 (N_7189,N_4583,N_4712);
and U7190 (N_7190,N_3650,N_3023);
or U7191 (N_7191,N_4496,N_4622);
nand U7192 (N_7192,N_2650,N_4622);
nand U7193 (N_7193,N_4117,N_4601);
or U7194 (N_7194,N_4871,N_3750);
and U7195 (N_7195,N_4042,N_3696);
or U7196 (N_7196,N_4567,N_3131);
nand U7197 (N_7197,N_4295,N_2888);
or U7198 (N_7198,N_4791,N_3093);
nor U7199 (N_7199,N_2960,N_3587);
nand U7200 (N_7200,N_4326,N_3863);
or U7201 (N_7201,N_3406,N_2979);
nand U7202 (N_7202,N_3146,N_3077);
or U7203 (N_7203,N_2955,N_4876);
nor U7204 (N_7204,N_3312,N_3187);
nor U7205 (N_7205,N_4692,N_4350);
nand U7206 (N_7206,N_4858,N_4707);
or U7207 (N_7207,N_3787,N_3010);
nand U7208 (N_7208,N_4617,N_4319);
nand U7209 (N_7209,N_2562,N_2729);
nor U7210 (N_7210,N_4025,N_4421);
nor U7211 (N_7211,N_4233,N_2537);
nor U7212 (N_7212,N_3088,N_2829);
nor U7213 (N_7213,N_4100,N_4719);
xnor U7214 (N_7214,N_4548,N_3164);
and U7215 (N_7215,N_4250,N_4175);
or U7216 (N_7216,N_4790,N_3338);
nand U7217 (N_7217,N_4759,N_2685);
or U7218 (N_7218,N_4193,N_4624);
and U7219 (N_7219,N_4934,N_4709);
xnor U7220 (N_7220,N_3231,N_3562);
or U7221 (N_7221,N_4791,N_4869);
and U7222 (N_7222,N_3236,N_4449);
and U7223 (N_7223,N_2857,N_4553);
nand U7224 (N_7224,N_3495,N_2656);
nand U7225 (N_7225,N_4764,N_3444);
or U7226 (N_7226,N_3331,N_4226);
and U7227 (N_7227,N_4196,N_2753);
nand U7228 (N_7228,N_2638,N_2525);
or U7229 (N_7229,N_2730,N_3960);
nand U7230 (N_7230,N_3606,N_4715);
nor U7231 (N_7231,N_3221,N_4965);
or U7232 (N_7232,N_3653,N_4745);
nand U7233 (N_7233,N_3684,N_2888);
and U7234 (N_7234,N_3489,N_3273);
or U7235 (N_7235,N_4025,N_3198);
nand U7236 (N_7236,N_3541,N_3330);
or U7237 (N_7237,N_3291,N_2514);
nand U7238 (N_7238,N_4336,N_2725);
nor U7239 (N_7239,N_3073,N_2537);
and U7240 (N_7240,N_4488,N_3059);
or U7241 (N_7241,N_2899,N_3983);
nor U7242 (N_7242,N_4510,N_4527);
or U7243 (N_7243,N_2545,N_4186);
or U7244 (N_7244,N_4457,N_3115);
nand U7245 (N_7245,N_4436,N_3799);
and U7246 (N_7246,N_4588,N_4863);
and U7247 (N_7247,N_2850,N_4555);
nand U7248 (N_7248,N_3758,N_2770);
and U7249 (N_7249,N_4366,N_3936);
nor U7250 (N_7250,N_3765,N_3209);
nand U7251 (N_7251,N_3406,N_3377);
nor U7252 (N_7252,N_2561,N_3630);
and U7253 (N_7253,N_4033,N_4625);
nor U7254 (N_7254,N_3314,N_4256);
or U7255 (N_7255,N_4711,N_3477);
or U7256 (N_7256,N_3292,N_4036);
or U7257 (N_7257,N_4064,N_2938);
nor U7258 (N_7258,N_3978,N_3078);
nand U7259 (N_7259,N_4009,N_3171);
or U7260 (N_7260,N_3946,N_3109);
nor U7261 (N_7261,N_3306,N_2636);
nor U7262 (N_7262,N_4477,N_3210);
or U7263 (N_7263,N_2790,N_3903);
and U7264 (N_7264,N_4043,N_4878);
and U7265 (N_7265,N_4292,N_3334);
nand U7266 (N_7266,N_3639,N_3967);
and U7267 (N_7267,N_3404,N_3031);
or U7268 (N_7268,N_3328,N_4532);
and U7269 (N_7269,N_2866,N_3113);
and U7270 (N_7270,N_2678,N_4729);
and U7271 (N_7271,N_3201,N_3522);
or U7272 (N_7272,N_4859,N_3964);
and U7273 (N_7273,N_4666,N_4125);
nor U7274 (N_7274,N_3003,N_3019);
and U7275 (N_7275,N_3344,N_2817);
nor U7276 (N_7276,N_2787,N_3211);
and U7277 (N_7277,N_4037,N_2984);
and U7278 (N_7278,N_3458,N_3243);
nand U7279 (N_7279,N_4461,N_4371);
and U7280 (N_7280,N_4627,N_3101);
or U7281 (N_7281,N_3603,N_4494);
nand U7282 (N_7282,N_4440,N_2658);
and U7283 (N_7283,N_3991,N_3672);
nand U7284 (N_7284,N_4347,N_3885);
and U7285 (N_7285,N_3162,N_4125);
nand U7286 (N_7286,N_3628,N_3033);
and U7287 (N_7287,N_4903,N_3327);
nand U7288 (N_7288,N_2702,N_4472);
nand U7289 (N_7289,N_3694,N_4108);
or U7290 (N_7290,N_2873,N_3836);
nor U7291 (N_7291,N_3103,N_4943);
nand U7292 (N_7292,N_3821,N_4766);
nand U7293 (N_7293,N_4563,N_4790);
nor U7294 (N_7294,N_3969,N_2731);
and U7295 (N_7295,N_4634,N_3793);
and U7296 (N_7296,N_4856,N_3472);
nand U7297 (N_7297,N_3004,N_3738);
nor U7298 (N_7298,N_3323,N_2826);
nor U7299 (N_7299,N_4684,N_3139);
and U7300 (N_7300,N_2566,N_4605);
and U7301 (N_7301,N_4646,N_2649);
nand U7302 (N_7302,N_3984,N_3687);
or U7303 (N_7303,N_4617,N_4141);
and U7304 (N_7304,N_4632,N_4171);
and U7305 (N_7305,N_2803,N_3611);
nand U7306 (N_7306,N_3167,N_4839);
nor U7307 (N_7307,N_2860,N_4948);
nand U7308 (N_7308,N_4811,N_3873);
and U7309 (N_7309,N_3910,N_2884);
nor U7310 (N_7310,N_4821,N_3066);
nand U7311 (N_7311,N_3474,N_4548);
and U7312 (N_7312,N_4493,N_3371);
nor U7313 (N_7313,N_4611,N_4517);
or U7314 (N_7314,N_4591,N_2896);
nor U7315 (N_7315,N_4408,N_3332);
and U7316 (N_7316,N_4867,N_3100);
nand U7317 (N_7317,N_4404,N_2808);
nor U7318 (N_7318,N_3631,N_2579);
and U7319 (N_7319,N_2789,N_4966);
nand U7320 (N_7320,N_3887,N_4645);
nor U7321 (N_7321,N_3899,N_3300);
nor U7322 (N_7322,N_4331,N_2934);
nor U7323 (N_7323,N_3235,N_2960);
and U7324 (N_7324,N_3634,N_2626);
and U7325 (N_7325,N_4105,N_3485);
nand U7326 (N_7326,N_4997,N_4229);
and U7327 (N_7327,N_3154,N_4792);
and U7328 (N_7328,N_2871,N_3966);
and U7329 (N_7329,N_3790,N_4973);
and U7330 (N_7330,N_2765,N_4819);
nor U7331 (N_7331,N_4628,N_4382);
nor U7332 (N_7332,N_4570,N_3748);
nand U7333 (N_7333,N_4388,N_3084);
nand U7334 (N_7334,N_3330,N_2575);
and U7335 (N_7335,N_4614,N_4181);
or U7336 (N_7336,N_4068,N_4221);
nand U7337 (N_7337,N_2724,N_4851);
nor U7338 (N_7338,N_3488,N_3969);
or U7339 (N_7339,N_3800,N_3985);
nor U7340 (N_7340,N_3680,N_3269);
nand U7341 (N_7341,N_4855,N_4293);
nor U7342 (N_7342,N_2515,N_4140);
nand U7343 (N_7343,N_3564,N_3914);
and U7344 (N_7344,N_2677,N_3576);
and U7345 (N_7345,N_4648,N_2929);
nor U7346 (N_7346,N_3048,N_4894);
nand U7347 (N_7347,N_4520,N_4957);
and U7348 (N_7348,N_3533,N_4638);
nor U7349 (N_7349,N_4521,N_4979);
nand U7350 (N_7350,N_3083,N_2895);
and U7351 (N_7351,N_4714,N_2691);
nand U7352 (N_7352,N_4971,N_3205);
or U7353 (N_7353,N_3850,N_3616);
nor U7354 (N_7354,N_3061,N_3408);
and U7355 (N_7355,N_2623,N_3189);
or U7356 (N_7356,N_3674,N_4119);
nor U7357 (N_7357,N_4816,N_3300);
nor U7358 (N_7358,N_4099,N_4748);
or U7359 (N_7359,N_4518,N_4841);
nor U7360 (N_7360,N_2672,N_2928);
and U7361 (N_7361,N_3746,N_4105);
and U7362 (N_7362,N_4758,N_4515);
or U7363 (N_7363,N_2932,N_4271);
nor U7364 (N_7364,N_4173,N_3754);
nand U7365 (N_7365,N_4568,N_2694);
nand U7366 (N_7366,N_4645,N_3018);
or U7367 (N_7367,N_4505,N_4002);
and U7368 (N_7368,N_3032,N_3479);
nand U7369 (N_7369,N_4699,N_3488);
nand U7370 (N_7370,N_4528,N_2891);
or U7371 (N_7371,N_2574,N_4981);
nor U7372 (N_7372,N_4887,N_4834);
nand U7373 (N_7373,N_3661,N_3493);
and U7374 (N_7374,N_4732,N_2739);
nand U7375 (N_7375,N_4149,N_4688);
and U7376 (N_7376,N_4111,N_4614);
nand U7377 (N_7377,N_3389,N_3589);
nand U7378 (N_7378,N_4178,N_3884);
nor U7379 (N_7379,N_3904,N_4205);
nor U7380 (N_7380,N_3721,N_3783);
or U7381 (N_7381,N_4048,N_4907);
and U7382 (N_7382,N_4011,N_4296);
nor U7383 (N_7383,N_4089,N_2684);
nand U7384 (N_7384,N_3055,N_3387);
or U7385 (N_7385,N_2538,N_3905);
and U7386 (N_7386,N_3203,N_2666);
nand U7387 (N_7387,N_3904,N_4845);
or U7388 (N_7388,N_4033,N_3350);
nor U7389 (N_7389,N_4519,N_4765);
and U7390 (N_7390,N_4737,N_3135);
nor U7391 (N_7391,N_3009,N_3513);
and U7392 (N_7392,N_3073,N_3022);
or U7393 (N_7393,N_3224,N_3992);
nand U7394 (N_7394,N_4936,N_3499);
and U7395 (N_7395,N_2542,N_2744);
or U7396 (N_7396,N_3133,N_4395);
nor U7397 (N_7397,N_2644,N_2566);
nor U7398 (N_7398,N_4933,N_3406);
and U7399 (N_7399,N_2995,N_3452);
nand U7400 (N_7400,N_3661,N_4084);
xor U7401 (N_7401,N_4654,N_3717);
nand U7402 (N_7402,N_3771,N_3738);
or U7403 (N_7403,N_2974,N_2857);
or U7404 (N_7404,N_4480,N_3534);
or U7405 (N_7405,N_3647,N_3861);
and U7406 (N_7406,N_3759,N_2566);
nand U7407 (N_7407,N_2700,N_3376);
and U7408 (N_7408,N_3393,N_3113);
nor U7409 (N_7409,N_4195,N_4741);
and U7410 (N_7410,N_3890,N_3945);
nor U7411 (N_7411,N_4000,N_3208);
nand U7412 (N_7412,N_3766,N_3250);
nor U7413 (N_7413,N_3679,N_4285);
or U7414 (N_7414,N_3119,N_3510);
and U7415 (N_7415,N_3146,N_3724);
and U7416 (N_7416,N_3997,N_3801);
nand U7417 (N_7417,N_2677,N_2865);
nor U7418 (N_7418,N_4703,N_3602);
and U7419 (N_7419,N_3550,N_2708);
or U7420 (N_7420,N_4519,N_2794);
or U7421 (N_7421,N_3851,N_3706);
or U7422 (N_7422,N_4671,N_3771);
xor U7423 (N_7423,N_4888,N_3561);
and U7424 (N_7424,N_4160,N_2940);
nand U7425 (N_7425,N_4293,N_2716);
and U7426 (N_7426,N_4311,N_3434);
and U7427 (N_7427,N_2887,N_2916);
nand U7428 (N_7428,N_3103,N_2638);
or U7429 (N_7429,N_3690,N_2886);
nor U7430 (N_7430,N_4882,N_3108);
and U7431 (N_7431,N_3794,N_3318);
or U7432 (N_7432,N_3405,N_2593);
or U7433 (N_7433,N_4069,N_3394);
and U7434 (N_7434,N_3407,N_3144);
nor U7435 (N_7435,N_2908,N_4452);
nand U7436 (N_7436,N_3344,N_3908);
or U7437 (N_7437,N_4064,N_2992);
or U7438 (N_7438,N_4548,N_3058);
and U7439 (N_7439,N_4162,N_3582);
or U7440 (N_7440,N_3179,N_3344);
or U7441 (N_7441,N_4946,N_4224);
nand U7442 (N_7442,N_4416,N_2593);
or U7443 (N_7443,N_3190,N_4943);
or U7444 (N_7444,N_4112,N_3766);
nand U7445 (N_7445,N_2821,N_3144);
and U7446 (N_7446,N_2922,N_2586);
nor U7447 (N_7447,N_3105,N_3992);
or U7448 (N_7448,N_2903,N_3772);
nor U7449 (N_7449,N_2581,N_3931);
nor U7450 (N_7450,N_3997,N_3436);
nand U7451 (N_7451,N_4934,N_3094);
and U7452 (N_7452,N_3893,N_4487);
and U7453 (N_7453,N_4114,N_4183);
nand U7454 (N_7454,N_4540,N_4592);
nor U7455 (N_7455,N_4425,N_4710);
nand U7456 (N_7456,N_3536,N_4767);
nor U7457 (N_7457,N_3072,N_3369);
nor U7458 (N_7458,N_2934,N_4096);
and U7459 (N_7459,N_4512,N_4521);
nor U7460 (N_7460,N_3140,N_4908);
or U7461 (N_7461,N_3342,N_4902);
nand U7462 (N_7462,N_3733,N_3463);
nor U7463 (N_7463,N_3887,N_3270);
xor U7464 (N_7464,N_4033,N_3929);
nor U7465 (N_7465,N_3803,N_4670);
or U7466 (N_7466,N_3430,N_4279);
or U7467 (N_7467,N_3946,N_3497);
nand U7468 (N_7468,N_4734,N_3699);
and U7469 (N_7469,N_2736,N_4573);
nand U7470 (N_7470,N_4722,N_4299);
nor U7471 (N_7471,N_4842,N_3035);
nand U7472 (N_7472,N_4843,N_2807);
nand U7473 (N_7473,N_3332,N_2627);
nand U7474 (N_7474,N_4551,N_2765);
nand U7475 (N_7475,N_4490,N_3814);
nand U7476 (N_7476,N_2949,N_2587);
nor U7477 (N_7477,N_3183,N_4572);
or U7478 (N_7478,N_3542,N_3807);
nand U7479 (N_7479,N_4381,N_3374);
and U7480 (N_7480,N_4658,N_3711);
or U7481 (N_7481,N_2915,N_3847);
and U7482 (N_7482,N_2622,N_3021);
and U7483 (N_7483,N_3029,N_4864);
or U7484 (N_7484,N_4099,N_4813);
and U7485 (N_7485,N_2787,N_4402);
or U7486 (N_7486,N_4375,N_3046);
nand U7487 (N_7487,N_2894,N_4996);
or U7488 (N_7488,N_3324,N_4225);
nor U7489 (N_7489,N_4771,N_2529);
and U7490 (N_7490,N_3872,N_4064);
or U7491 (N_7491,N_4282,N_4272);
and U7492 (N_7492,N_4262,N_4893);
nand U7493 (N_7493,N_4006,N_2517);
or U7494 (N_7494,N_3498,N_4345);
or U7495 (N_7495,N_3555,N_3333);
or U7496 (N_7496,N_3997,N_4955);
and U7497 (N_7497,N_2960,N_3104);
nand U7498 (N_7498,N_4797,N_3156);
and U7499 (N_7499,N_4474,N_4849);
and U7500 (N_7500,N_6145,N_5343);
nand U7501 (N_7501,N_7002,N_6358);
and U7502 (N_7502,N_7160,N_5661);
nand U7503 (N_7503,N_7386,N_5688);
nand U7504 (N_7504,N_5142,N_6940);
or U7505 (N_7505,N_6737,N_6905);
nor U7506 (N_7506,N_7154,N_7390);
or U7507 (N_7507,N_5791,N_6198);
nor U7508 (N_7508,N_5497,N_6763);
nand U7509 (N_7509,N_6000,N_6510);
and U7510 (N_7510,N_6027,N_6294);
xnor U7511 (N_7511,N_5905,N_6394);
nand U7512 (N_7512,N_5761,N_6893);
or U7513 (N_7513,N_5704,N_6982);
nor U7514 (N_7514,N_7023,N_6711);
or U7515 (N_7515,N_7289,N_6659);
nand U7516 (N_7516,N_6962,N_5233);
nand U7517 (N_7517,N_6330,N_6877);
and U7518 (N_7518,N_5380,N_5296);
and U7519 (N_7519,N_7279,N_6464);
nand U7520 (N_7520,N_7372,N_5702);
and U7521 (N_7521,N_5340,N_5718);
nand U7522 (N_7522,N_6752,N_6726);
nor U7523 (N_7523,N_5051,N_6835);
nand U7524 (N_7524,N_6170,N_6578);
or U7525 (N_7525,N_6319,N_5720);
nor U7526 (N_7526,N_6239,N_5395);
nor U7527 (N_7527,N_5848,N_5262);
and U7528 (N_7528,N_7064,N_5199);
or U7529 (N_7529,N_6479,N_6998);
nand U7530 (N_7530,N_7342,N_5279);
xnor U7531 (N_7531,N_6790,N_6252);
and U7532 (N_7532,N_5064,N_5630);
nand U7533 (N_7533,N_7183,N_5636);
nor U7534 (N_7534,N_5339,N_5842);
nor U7535 (N_7535,N_6825,N_5959);
and U7536 (N_7536,N_7124,N_5878);
or U7537 (N_7537,N_5290,N_7441);
nand U7538 (N_7538,N_7428,N_5972);
nand U7539 (N_7539,N_6341,N_6728);
and U7540 (N_7540,N_7267,N_7405);
and U7541 (N_7541,N_5113,N_5446);
nand U7542 (N_7542,N_6587,N_6543);
and U7543 (N_7543,N_5460,N_7226);
or U7544 (N_7544,N_5091,N_5531);
or U7545 (N_7545,N_5190,N_5278);
or U7546 (N_7546,N_6303,N_6591);
or U7547 (N_7547,N_5696,N_5889);
nand U7548 (N_7548,N_5969,N_6794);
nand U7549 (N_7549,N_5373,N_5714);
nor U7550 (N_7550,N_6514,N_6563);
nor U7551 (N_7551,N_7102,N_7085);
nand U7552 (N_7552,N_6759,N_6118);
nor U7553 (N_7553,N_6805,N_6097);
xnor U7554 (N_7554,N_5646,N_7337);
and U7555 (N_7555,N_6882,N_6971);
and U7556 (N_7556,N_7158,N_6574);
and U7557 (N_7557,N_6683,N_5964);
nor U7558 (N_7558,N_5161,N_5455);
and U7559 (N_7559,N_6180,N_5287);
or U7560 (N_7560,N_7254,N_5214);
nand U7561 (N_7561,N_7317,N_5856);
or U7562 (N_7562,N_5949,N_5479);
nor U7563 (N_7563,N_6934,N_6916);
nand U7564 (N_7564,N_6743,N_5028);
nor U7565 (N_7565,N_5013,N_6401);
nor U7566 (N_7566,N_5633,N_5082);
nand U7567 (N_7567,N_7482,N_6979);
or U7568 (N_7568,N_5819,N_6436);
nor U7569 (N_7569,N_5937,N_6349);
nand U7570 (N_7570,N_6645,N_5726);
and U7571 (N_7571,N_6379,N_5100);
or U7572 (N_7572,N_5931,N_5077);
nand U7573 (N_7573,N_7392,N_6206);
and U7574 (N_7574,N_5768,N_6875);
nor U7575 (N_7575,N_6070,N_7086);
nor U7576 (N_7576,N_7403,N_6526);
nor U7577 (N_7577,N_6710,N_6599);
or U7578 (N_7578,N_6700,N_6864);
or U7579 (N_7579,N_6692,N_6681);
or U7580 (N_7580,N_6884,N_7437);
or U7581 (N_7581,N_7103,N_6985);
nand U7582 (N_7582,N_7224,N_6111);
nor U7583 (N_7583,N_6634,N_7370);
nand U7584 (N_7584,N_6192,N_6693);
nor U7585 (N_7585,N_5269,N_7000);
nand U7586 (N_7586,N_5315,N_5534);
or U7587 (N_7587,N_5106,N_7299);
and U7588 (N_7588,N_6222,N_6656);
nor U7589 (N_7589,N_6902,N_6872);
and U7590 (N_7590,N_7033,N_6623);
nor U7591 (N_7591,N_6562,N_6449);
and U7592 (N_7592,N_6997,N_5514);
and U7593 (N_7593,N_5505,N_5140);
nand U7594 (N_7594,N_6371,N_6477);
nand U7595 (N_7595,N_5752,N_5435);
or U7596 (N_7596,N_7179,N_6175);
nor U7597 (N_7597,N_5176,N_7368);
or U7598 (N_7598,N_7380,N_7166);
nor U7599 (N_7599,N_7399,N_5986);
or U7600 (N_7600,N_7051,N_6618);
nor U7601 (N_7601,N_5466,N_5488);
nand U7602 (N_7602,N_6775,N_5162);
nand U7603 (N_7603,N_5489,N_5298);
nor U7604 (N_7604,N_7088,N_5256);
nand U7605 (N_7605,N_5102,N_5118);
nand U7606 (N_7606,N_5332,N_6461);
nor U7607 (N_7607,N_5863,N_7150);
and U7608 (N_7608,N_6367,N_7151);
nand U7609 (N_7609,N_5763,N_6582);
nor U7610 (N_7610,N_5486,N_6124);
and U7611 (N_7611,N_6523,N_5306);
nor U7612 (N_7612,N_7209,N_6856);
nand U7613 (N_7613,N_6983,N_6189);
or U7614 (N_7614,N_5825,N_7436);
or U7615 (N_7615,N_6253,N_5253);
or U7616 (N_7616,N_5745,N_5780);
nand U7617 (N_7617,N_5400,N_6363);
or U7618 (N_7618,N_5483,N_7439);
or U7619 (N_7619,N_5284,N_5494);
or U7620 (N_7620,N_7291,N_7340);
and U7621 (N_7621,N_5731,N_6501);
or U7622 (N_7622,N_5853,N_5172);
and U7623 (N_7623,N_7463,N_7449);
or U7624 (N_7624,N_5653,N_5007);
and U7625 (N_7625,N_7475,N_6063);
nand U7626 (N_7626,N_7229,N_6376);
nor U7627 (N_7627,N_7255,N_5705);
nor U7628 (N_7628,N_6791,N_6020);
nand U7629 (N_7629,N_5174,N_5979);
nand U7630 (N_7630,N_7050,N_6719);
and U7631 (N_7631,N_6762,N_6570);
nor U7632 (N_7632,N_6758,N_5195);
nor U7633 (N_7633,N_6018,N_5620);
nand U7634 (N_7634,N_6107,N_5366);
and U7635 (N_7635,N_5708,N_5880);
and U7636 (N_7636,N_7235,N_5834);
and U7637 (N_7637,N_7132,N_5010);
or U7638 (N_7638,N_6411,N_5442);
or U7639 (N_7639,N_6955,N_6249);
nor U7640 (N_7640,N_5755,N_5440);
nand U7641 (N_7641,N_6845,N_7334);
nor U7642 (N_7642,N_5178,N_5042);
and U7643 (N_7643,N_5907,N_6141);
nor U7644 (N_7644,N_7264,N_5612);
nor U7645 (N_7645,N_5533,N_5684);
and U7646 (N_7646,N_7323,N_7478);
nor U7647 (N_7647,N_7492,N_5350);
and U7648 (N_7648,N_6136,N_6876);
or U7649 (N_7649,N_5131,N_5980);
nand U7650 (N_7650,N_6002,N_7363);
nand U7651 (N_7651,N_7397,N_6725);
nand U7652 (N_7652,N_6478,N_7316);
or U7653 (N_7653,N_6053,N_5790);
and U7654 (N_7654,N_7141,N_7322);
and U7655 (N_7655,N_6888,N_5736);
nor U7656 (N_7656,N_7073,N_5618);
nor U7657 (N_7657,N_5918,N_6324);
and U7658 (N_7658,N_6515,N_6355);
nor U7659 (N_7659,N_6615,N_5313);
and U7660 (N_7660,N_6680,N_7353);
xor U7661 (N_7661,N_5286,N_6544);
or U7662 (N_7662,N_5149,N_6891);
and U7663 (N_7663,N_5751,N_6148);
nor U7664 (N_7664,N_6142,N_6316);
or U7665 (N_7665,N_5583,N_5798);
nor U7666 (N_7666,N_5194,N_5732);
and U7667 (N_7667,N_5982,N_5811);
and U7668 (N_7668,N_6270,N_6497);
and U7669 (N_7669,N_5554,N_5881);
nor U7670 (N_7670,N_5629,N_7230);
nor U7671 (N_7671,N_5717,N_5478);
or U7672 (N_7672,N_5643,N_5966);
nor U7673 (N_7673,N_6164,N_5060);
or U7674 (N_7674,N_5401,N_5901);
nand U7675 (N_7675,N_6325,N_6240);
nor U7676 (N_7676,N_5295,N_7159);
and U7677 (N_7677,N_7280,N_5860);
nor U7678 (N_7678,N_6250,N_6028);
and U7679 (N_7679,N_6244,N_6248);
and U7680 (N_7680,N_7349,N_7007);
or U7681 (N_7681,N_7129,N_6128);
nand U7682 (N_7682,N_7225,N_5125);
or U7683 (N_7683,N_5816,N_7288);
nor U7684 (N_7684,N_5083,N_5965);
and U7685 (N_7685,N_6345,N_5338);
nand U7686 (N_7686,N_5536,N_6936);
and U7687 (N_7687,N_5275,N_5764);
and U7688 (N_7688,N_5086,N_6978);
nand U7689 (N_7689,N_6718,N_7243);
nand U7690 (N_7690,N_5715,N_6846);
or U7691 (N_7691,N_5826,N_5428);
or U7692 (N_7692,N_6412,N_7341);
and U7693 (N_7693,N_5151,N_5387);
nor U7694 (N_7694,N_5379,N_5258);
and U7695 (N_7695,N_6369,N_6406);
and U7696 (N_7696,N_5852,N_6465);
nor U7697 (N_7697,N_6799,N_5706);
and U7698 (N_7698,N_5270,N_6105);
nor U7699 (N_7699,N_7027,N_6057);
and U7700 (N_7700,N_7458,N_7336);
and U7701 (N_7701,N_7090,N_5989);
and U7702 (N_7702,N_7447,N_6911);
and U7703 (N_7703,N_6652,N_6422);
and U7704 (N_7704,N_5650,N_6443);
and U7705 (N_7705,N_6722,N_5575);
xor U7706 (N_7706,N_5666,N_6704);
nand U7707 (N_7707,N_6397,N_6427);
nand U7708 (N_7708,N_6382,N_6573);
nor U7709 (N_7709,N_7101,N_7057);
nand U7710 (N_7710,N_5915,N_6387);
and U7711 (N_7711,N_6372,N_6096);
nor U7712 (N_7712,N_6944,N_7009);
nand U7713 (N_7713,N_6460,N_6662);
nand U7714 (N_7714,N_5364,N_7443);
and U7715 (N_7715,N_5875,N_5866);
nand U7716 (N_7716,N_6641,N_6739);
or U7717 (N_7717,N_5375,N_6467);
or U7718 (N_7718,N_6988,N_7055);
and U7719 (N_7719,N_5261,N_5529);
or U7720 (N_7720,N_5458,N_7419);
or U7721 (N_7721,N_5712,N_6429);
nor U7722 (N_7722,N_6259,N_6607);
nand U7723 (N_7723,N_6228,N_5838);
nand U7724 (N_7724,N_6043,N_5527);
nor U7725 (N_7725,N_6409,N_6616);
and U7726 (N_7726,N_7261,N_7082);
or U7727 (N_7727,N_6104,N_6407);
or U7728 (N_7728,N_5030,N_6328);
nand U7729 (N_7729,N_5724,N_6741);
nand U7730 (N_7730,N_5570,N_7219);
nor U7731 (N_7731,N_5021,N_7016);
nand U7732 (N_7732,N_6859,N_7048);
or U7733 (N_7733,N_5242,N_7022);
or U7734 (N_7734,N_6229,N_6207);
or U7735 (N_7735,N_7417,N_6132);
or U7736 (N_7736,N_6871,N_6702);
nor U7737 (N_7737,N_7237,N_5119);
or U7738 (N_7738,N_5464,N_5044);
nand U7739 (N_7739,N_7369,N_6356);
and U7740 (N_7740,N_7177,N_6542);
or U7741 (N_7741,N_5203,N_6258);
and U7742 (N_7742,N_6194,N_6052);
or U7743 (N_7743,N_5652,N_5039);
or U7744 (N_7744,N_7497,N_6046);
nor U7745 (N_7745,N_5234,N_6143);
nor U7746 (N_7746,N_6486,N_6083);
and U7747 (N_7747,N_5208,N_7496);
or U7748 (N_7748,N_7347,N_6747);
or U7749 (N_7749,N_5941,N_5268);
or U7750 (N_7750,N_7355,N_5823);
and U7751 (N_7751,N_6770,N_6205);
nor U7752 (N_7752,N_6802,N_5674);
or U7753 (N_7753,N_7295,N_5267);
nor U7754 (N_7754,N_7400,N_6195);
nand U7755 (N_7755,N_5308,N_6246);
or U7756 (N_7756,N_7139,N_6772);
nor U7757 (N_7757,N_6773,N_6651);
or U7758 (N_7758,N_7311,N_5774);
nand U7759 (N_7759,N_5422,N_7494);
and U7760 (N_7760,N_6441,N_5182);
nor U7761 (N_7761,N_6423,N_6660);
nand U7762 (N_7762,N_5777,N_6342);
nand U7763 (N_7763,N_6211,N_6044);
and U7764 (N_7764,N_6226,N_6473);
and U7765 (N_7765,N_6224,N_5563);
xor U7766 (N_7766,N_7402,N_5681);
nand U7767 (N_7767,N_6072,N_5632);
or U7768 (N_7768,N_6927,N_6099);
nand U7769 (N_7769,N_7100,N_6903);
or U7770 (N_7770,N_7123,N_7327);
nand U7771 (N_7771,N_5266,N_7412);
nor U7772 (N_7772,N_6992,N_5782);
nand U7773 (N_7773,N_5624,N_6314);
nand U7774 (N_7774,N_6863,N_7253);
nor U7775 (N_7775,N_5024,N_6865);
or U7776 (N_7776,N_6391,N_7360);
nor U7777 (N_7777,N_5382,N_6067);
nor U7778 (N_7778,N_5167,N_6162);
and U7779 (N_7779,N_6504,N_6381);
nor U7780 (N_7780,N_7221,N_7283);
or U7781 (N_7781,N_5961,N_5457);
and U7782 (N_7782,N_6450,N_5225);
or U7783 (N_7783,N_6167,N_5904);
or U7784 (N_7784,N_7152,N_5733);
or U7785 (N_7785,N_6405,N_5574);
and U7786 (N_7786,N_7157,N_6041);
or U7787 (N_7787,N_5381,N_6939);
nor U7788 (N_7788,N_6622,N_6631);
or U7789 (N_7789,N_5076,N_6291);
nand U7790 (N_7790,N_5254,N_7074);
nand U7791 (N_7791,N_6675,N_7115);
nor U7792 (N_7792,N_5232,N_7217);
nor U7793 (N_7793,N_6188,N_7053);
nand U7794 (N_7794,N_5509,N_6352);
and U7795 (N_7795,N_6673,N_5245);
nand U7796 (N_7796,N_5515,N_6075);
nor U7797 (N_7797,N_7364,N_7054);
and U7798 (N_7798,N_5074,N_5571);
or U7799 (N_7799,N_7144,N_5065);
nor U7800 (N_7800,N_5283,N_6370);
nor U7801 (N_7801,N_6416,N_6365);
and U7802 (N_7802,N_7131,N_5827);
nand U7803 (N_7803,N_6343,N_6779);
and U7804 (N_7804,N_7005,N_6781);
nor U7805 (N_7805,N_5396,N_5410);
nor U7806 (N_7806,N_5050,N_7306);
nor U7807 (N_7807,N_5601,N_6163);
nand U7808 (N_7808,N_7444,N_6899);
nor U7809 (N_7809,N_6947,N_5311);
and U7810 (N_7810,N_7361,N_6265);
nand U7811 (N_7811,N_5333,N_6446);
and U7812 (N_7812,N_5744,N_5522);
or U7813 (N_7813,N_6843,N_6418);
nor U7814 (N_7814,N_5716,N_5792);
and U7815 (N_7815,N_6468,N_6932);
or U7816 (N_7816,N_6953,N_6881);
nand U7817 (N_7817,N_6442,N_6968);
and U7818 (N_7818,N_7003,N_6530);
and U7819 (N_7819,N_5196,N_5588);
nor U7820 (N_7820,N_6952,N_6642);
or U7821 (N_7821,N_5784,N_7108);
and U7822 (N_7822,N_6281,N_7236);
or U7823 (N_7823,N_5282,N_7499);
or U7824 (N_7824,N_5540,N_6009);
nand U7825 (N_7825,N_7195,N_6855);
nand U7826 (N_7826,N_5775,N_5679);
or U7827 (N_7827,N_5205,N_7382);
and U7828 (N_7828,N_5222,N_5080);
or U7829 (N_7829,N_5274,N_6995);
or U7830 (N_7830,N_7422,N_5459);
and U7831 (N_7831,N_7287,N_7142);
nand U7832 (N_7832,N_5993,N_5445);
nor U7833 (N_7833,N_6546,N_5701);
or U7834 (N_7834,N_7099,N_5526);
nor U7835 (N_7835,N_6402,N_7191);
nand U7836 (N_7836,N_5465,N_6392);
nor U7837 (N_7837,N_7296,N_5351);
or U7838 (N_7838,N_7378,N_5146);
and U7839 (N_7839,N_6077,N_7168);
and U7840 (N_7840,N_6059,N_5448);
or U7841 (N_7841,N_6216,N_6948);
nand U7842 (N_7842,N_6339,N_5691);
or U7843 (N_7843,N_6679,N_6254);
nor U7844 (N_7844,N_6567,N_6453);
nor U7845 (N_7845,N_5741,N_6961);
nor U7846 (N_7846,N_5215,N_5589);
xnor U7847 (N_7847,N_5319,N_7211);
and U7848 (N_7848,N_5155,N_6912);
or U7849 (N_7849,N_5911,N_7414);
and U7850 (N_7850,N_6808,N_5424);
nor U7851 (N_7851,N_5957,N_7024);
nand U7852 (N_7852,N_5061,N_7331);
and U7853 (N_7853,N_6147,N_5300);
nand U7854 (N_7854,N_5638,N_7259);
and U7855 (N_7855,N_6215,N_6428);
nor U7856 (N_7856,N_5198,N_7117);
nand U7857 (N_7857,N_6388,N_6946);
nand U7858 (N_7858,N_6081,N_5595);
and U7859 (N_7859,N_6271,N_6586);
nand U7860 (N_7860,N_7174,N_5663);
and U7861 (N_7861,N_6437,N_6016);
or U7862 (N_7862,N_7476,N_6089);
xor U7863 (N_7863,N_5939,N_7187);
nor U7864 (N_7864,N_5089,N_6774);
and U7865 (N_7865,N_5327,N_7484);
and U7866 (N_7866,N_5743,N_5619);
and U7867 (N_7867,N_5265,N_7469);
or U7868 (N_7868,N_5850,N_5425);
nor U7869 (N_7869,N_6021,N_7376);
nand U7870 (N_7870,N_6158,N_5090);
nor U7871 (N_7871,N_5081,N_5864);
nor U7872 (N_7872,N_6156,N_5492);
and U7873 (N_7873,N_7242,N_6151);
nor U7874 (N_7874,N_6347,N_6595);
nand U7875 (N_7875,N_6448,N_5328);
nor U7876 (N_7876,N_6285,N_6293);
or U7877 (N_7877,N_5239,N_5822);
or U7878 (N_7878,N_5138,N_6986);
nand U7879 (N_7879,N_5591,N_5087);
nand U7880 (N_7880,N_5305,N_7208);
nand U7881 (N_7881,N_6060,N_5431);
and U7882 (N_7882,N_6191,N_6015);
and U7883 (N_7883,N_5136,N_7346);
nand U7884 (N_7884,N_6237,N_6590);
nand U7885 (N_7885,N_6594,N_5748);
nor U7886 (N_7886,N_6333,N_7453);
nor U7887 (N_7887,N_5257,N_5555);
nand U7888 (N_7888,N_5271,N_6640);
nand U7889 (N_7889,N_5071,N_5452);
nor U7890 (N_7890,N_6307,N_5675);
or U7891 (N_7891,N_6236,N_5451);
nand U7892 (N_7892,N_6545,N_7391);
nor U7893 (N_7893,N_5603,N_7284);
nor U7894 (N_7894,N_5677,N_6247);
xor U7895 (N_7895,N_5159,N_7351);
and U7896 (N_7896,N_5924,N_6695);
or U7897 (N_7897,N_6208,N_7058);
nor U7898 (N_7898,N_7089,N_5615);
nand U7899 (N_7899,N_6832,N_6034);
nand U7900 (N_7900,N_6276,N_6470);
and U7901 (N_7901,N_5654,N_6055);
or U7902 (N_7902,N_7450,N_7461);
nand U7903 (N_7903,N_6621,N_7176);
and U7904 (N_7904,N_6264,N_6095);
nor U7905 (N_7905,N_7029,N_5046);
nand U7906 (N_7906,N_5128,N_5625);
nor U7907 (N_7907,N_5836,N_7328);
or U7908 (N_7908,N_5481,N_5635);
nand U7909 (N_7909,N_6928,N_6529);
nand U7910 (N_7910,N_5970,N_5829);
nor U7911 (N_7911,N_5157,N_7122);
and U7912 (N_7912,N_5892,N_5659);
nand U7913 (N_7913,N_5596,N_7012);
and U7914 (N_7914,N_6897,N_6697);
or U7915 (N_7915,N_6637,N_5525);
or U7916 (N_7916,N_5272,N_6575);
nor U7917 (N_7917,N_6223,N_6687);
or U7918 (N_7918,N_5600,N_5873);
and U7919 (N_7919,N_6149,N_6456);
nand U7920 (N_7920,N_6506,N_5568);
or U7921 (N_7921,N_7095,N_5660);
and U7922 (N_7922,N_6218,N_5248);
or U7923 (N_7923,N_7480,N_5499);
or U7924 (N_7924,N_5491,N_5068);
nand U7925 (N_7925,N_5839,N_6197);
nand U7926 (N_7926,N_5056,N_6821);
nand U7927 (N_7927,N_6909,N_5349);
or U7928 (N_7928,N_6108,N_5587);
xnor U7929 (N_7929,N_7020,N_7119);
nand U7930 (N_7930,N_6812,N_7344);
nand U7931 (N_7931,N_6671,N_5228);
and U7932 (N_7932,N_5797,N_5477);
or U7933 (N_7933,N_5043,N_7169);
and U7934 (N_7934,N_6001,N_6026);
nor U7935 (N_7935,N_5399,N_6404);
or U7936 (N_7936,N_5032,N_7348);
or U7937 (N_7937,N_5407,N_5160);
nor U7938 (N_7938,N_5981,N_5219);
nor U7939 (N_7939,N_6445,N_7145);
or U7940 (N_7940,N_7199,N_5285);
or U7941 (N_7941,N_7113,N_7079);
or U7942 (N_7942,N_6666,N_6256);
or U7943 (N_7943,N_7314,N_5882);
nor U7944 (N_7944,N_6649,N_5651);
nand U7945 (N_7945,N_5847,N_6549);
nand U7946 (N_7946,N_7134,N_5148);
nand U7947 (N_7947,N_7013,N_5134);
or U7948 (N_7948,N_5210,N_5132);
and U7949 (N_7949,N_6701,N_7147);
or U7950 (N_7950,N_7472,N_6630);
and U7951 (N_7951,N_6789,N_5067);
and U7952 (N_7952,N_5078,N_7362);
and U7953 (N_7953,N_6740,N_5055);
or U7954 (N_7954,N_6713,N_7366);
and U7955 (N_7955,N_5700,N_6929);
nand U7956 (N_7956,N_5259,N_5211);
nor U7957 (N_7957,N_6426,N_6869);
nor U7958 (N_7958,N_6155,N_5184);
nor U7959 (N_7959,N_5206,N_6362);
nand U7960 (N_7960,N_5001,N_6179);
and U7961 (N_7961,N_5897,N_6166);
nor U7962 (N_7962,N_7215,N_6359);
nand U7963 (N_7963,N_6949,N_5687);
nor U7964 (N_7964,N_7034,N_5057);
nand U7965 (N_7965,N_6287,N_5095);
and U7966 (N_7966,N_5331,N_6699);
or U7967 (N_7967,N_7214,N_7474);
or U7968 (N_7968,N_7321,N_7423);
or U7969 (N_7969,N_5019,N_6963);
nand U7970 (N_7970,N_6977,N_5231);
nand U7971 (N_7971,N_5378,N_6487);
or U7972 (N_7972,N_5389,N_6677);
or U7973 (N_7973,N_5862,N_7047);
nor U7974 (N_7974,N_7276,N_5419);
nand U7975 (N_7975,N_5154,N_5070);
nand U7976 (N_7976,N_6357,N_5324);
nand U7977 (N_7977,N_7239,N_5000);
or U7978 (N_7978,N_5416,N_5686);
nor U7979 (N_7979,N_5747,N_5721);
nand U7980 (N_7980,N_5519,N_7257);
xnor U7981 (N_7981,N_6079,N_6727);
nand U7982 (N_7982,N_7452,N_5927);
nor U7983 (N_7983,N_5289,N_5197);
nand U7984 (N_7984,N_6811,N_5742);
or U7985 (N_7985,N_6323,N_5449);
and U7986 (N_7986,N_5634,N_6554);
nand U7987 (N_7987,N_6037,N_5512);
nor U7988 (N_7988,N_7354,N_5746);
and U7989 (N_7989,N_6661,N_5441);
nor U7990 (N_7990,N_6455,N_6798);
and U7991 (N_7991,N_6930,N_7008);
or U7992 (N_7992,N_6064,N_5830);
and U7993 (N_7993,N_6847,N_5213);
or U7994 (N_7994,N_5122,N_5226);
xor U7995 (N_7995,N_6308,N_6255);
and U7996 (N_7996,N_6724,N_6138);
or U7997 (N_7997,N_6190,N_5586);
or U7998 (N_7998,N_7080,N_5063);
nand U7999 (N_7999,N_6756,N_6769);
nand U8000 (N_8000,N_7190,N_6159);
nor U8001 (N_8001,N_6459,N_5402);
nand U8002 (N_8002,N_6560,N_7281);
nand U8003 (N_8003,N_6600,N_5942);
nor U8004 (N_8004,N_6503,N_6417);
nand U8005 (N_8005,N_5936,N_7332);
nor U8006 (N_8006,N_6196,N_7359);
xnor U8007 (N_8007,N_7120,N_6498);
nor U8008 (N_8008,N_5928,N_6913);
nand U8009 (N_8009,N_6419,N_5240);
nand U8010 (N_8010,N_6827,N_5599);
nor U8011 (N_8011,N_7192,N_6536);
and U8012 (N_8012,N_5454,N_6140);
or U8013 (N_8013,N_6901,N_6605);
nor U8014 (N_8014,N_7062,N_6251);
nor U8015 (N_8015,N_6750,N_5566);
and U8016 (N_8016,N_5357,N_7293);
nor U8017 (N_8017,N_7188,N_5580);
or U8018 (N_8018,N_5695,N_6466);
nor U8019 (N_8019,N_6221,N_6655);
and U8020 (N_8020,N_6767,N_6139);
and U8021 (N_8021,N_6433,N_7164);
nor U8022 (N_8022,N_5246,N_6261);
nor U8023 (N_8023,N_7127,N_6822);
and U8024 (N_8024,N_6326,N_6174);
nand U8025 (N_8025,N_6654,N_5758);
nand U8026 (N_8026,N_5318,N_5840);
or U8027 (N_8027,N_6608,N_7307);
and U8028 (N_8028,N_5163,N_6113);
nand U8029 (N_8029,N_6220,N_7075);
nor U8030 (N_8030,N_7451,N_5079);
nor U8031 (N_8031,N_5408,N_7133);
and U8032 (N_8032,N_7308,N_6518);
or U8033 (N_8033,N_5785,N_5141);
and U8034 (N_8034,N_5938,N_6547);
nor U8035 (N_8035,N_7410,N_6959);
nand U8036 (N_8036,N_5807,N_7087);
and U8037 (N_8037,N_5053,N_6795);
xnor U8038 (N_8038,N_5516,N_5556);
or U8039 (N_8039,N_5922,N_5414);
or U8040 (N_8040,N_6296,N_6302);
nand U8041 (N_8041,N_5096,N_7069);
and U8042 (N_8042,N_6217,N_6993);
and U8043 (N_8043,N_5577,N_6736);
or U8044 (N_8044,N_7434,N_6807);
or U8045 (N_8045,N_5301,N_6625);
or U8046 (N_8046,N_7250,N_6100);
xor U8047 (N_8047,N_5126,N_6183);
nand U8048 (N_8048,N_5069,N_6996);
or U8049 (N_8049,N_5626,N_5690);
and U8050 (N_8050,N_6908,N_5365);
nand U8051 (N_8051,N_5362,N_5598);
nand U8052 (N_8052,N_6049,N_6047);
and U8053 (N_8053,N_6494,N_6824);
or U8054 (N_8054,N_7271,N_7248);
and U8055 (N_8055,N_5770,N_6786);
or U8056 (N_8056,N_6120,N_5845);
nand U8057 (N_8057,N_7184,N_5562);
nand U8058 (N_8058,N_7042,N_6242);
and U8059 (N_8059,N_6335,N_7438);
and U8060 (N_8060,N_7305,N_6245);
nand U8061 (N_8061,N_6490,N_5417);
nor U8062 (N_8062,N_5956,N_6213);
nor U8063 (N_8063,N_5361,N_6629);
nor U8064 (N_8064,N_6234,N_6941);
or U8065 (N_8065,N_5179,N_6492);
or U8066 (N_8066,N_6130,N_6212);
or U8067 (N_8067,N_6716,N_6885);
nor U8068 (N_8068,N_5776,N_5247);
and U8069 (N_8069,N_7333,N_5009);
or U8070 (N_8070,N_6088,N_6676);
nor U8071 (N_8071,N_7375,N_6814);
or U8072 (N_8072,N_5244,N_6386);
and U8073 (N_8073,N_7228,N_6068);
nand U8074 (N_8074,N_5766,N_6819);
nand U8075 (N_8075,N_5934,N_5664);
or U8076 (N_8076,N_5910,N_6969);
nor U8077 (N_8077,N_6628,N_7040);
nand U8078 (N_8078,N_6867,N_6069);
and U8079 (N_8079,N_5342,N_5252);
nand U8080 (N_8080,N_6023,N_6493);
nor U8081 (N_8081,N_5806,N_5217);
and U8082 (N_8082,N_5075,N_7483);
nor U8083 (N_8083,N_5218,N_6286);
nand U8084 (N_8084,N_7223,N_5114);
nor U8085 (N_8085,N_6257,N_5369);
or U8086 (N_8086,N_5251,N_5461);
nor U8087 (N_8087,N_6525,N_7477);
or U8088 (N_8088,N_6375,N_7345);
nor U8089 (N_8089,N_5049,N_5180);
nand U8090 (N_8090,N_5846,N_5548);
nor U8091 (N_8091,N_6839,N_6395);
nand U8092 (N_8092,N_5487,N_6238);
and U8093 (N_8093,N_6277,N_5031);
or U8094 (N_8094,N_7206,N_6742);
and U8095 (N_8095,N_5299,N_5530);
nor U8096 (N_8096,N_6592,N_5757);
and U8097 (N_8097,N_6505,N_6288);
or U8098 (N_8098,N_5614,N_5730);
and U8099 (N_8099,N_5330,N_5953);
or U8100 (N_8100,N_7300,N_6974);
or U8101 (N_8101,N_6917,N_5902);
nand U8102 (N_8102,N_6564,N_7457);
nand U8103 (N_8103,N_5413,N_6298);
or U8104 (N_8104,N_5954,N_6850);
or U8105 (N_8105,N_7011,N_5018);
nand U8106 (N_8106,N_7357,N_7421);
or U8107 (N_8107,N_6366,N_5528);
or U8108 (N_8108,N_6569,N_5760);
or U8109 (N_8109,N_5320,N_5191);
or U8110 (N_8110,N_5971,N_6792);
or U8111 (N_8111,N_6678,N_6033);
and U8112 (N_8112,N_6636,N_6818);
nor U8113 (N_8113,N_5443,N_7470);
or U8114 (N_8114,N_5781,N_5621);
or U8115 (N_8115,N_5667,N_5789);
nand U8116 (N_8116,N_6894,N_7106);
nand U8117 (N_8117,N_5310,N_5805);
and U8118 (N_8118,N_5647,N_5040);
or U8119 (N_8119,N_7146,N_6066);
nand U8120 (N_8120,N_6091,N_5473);
and U8121 (N_8121,N_5861,N_6396);
nor U8122 (N_8122,N_5314,N_5994);
and U8123 (N_8123,N_5552,N_7456);
or U8124 (N_8124,N_7093,N_5277);
or U8125 (N_8125,N_5609,N_5950);
or U8126 (N_8126,N_5759,N_6619);
nor U8127 (N_8127,N_7493,N_6331);
nor U8128 (N_8128,N_6280,N_5325);
nand U8129 (N_8129,N_6474,N_5987);
nor U8130 (N_8130,N_7227,N_6421);
xor U8131 (N_8131,N_7467,N_6219);
and U8132 (N_8132,N_6810,N_5352);
nor U8133 (N_8133,N_5983,N_5337);
or U8134 (N_8134,N_5249,N_6266);
or U8135 (N_8135,N_7097,N_7339);
nand U8136 (N_8136,N_6481,N_5345);
or U8137 (N_8137,N_5243,N_5359);
or U8138 (N_8138,N_6793,N_6146);
nor U8139 (N_8139,N_6413,N_6535);
nor U8140 (N_8140,N_6844,N_5500);
and U8141 (N_8141,N_6160,N_6058);
xor U8142 (N_8142,N_5561,N_6836);
nand U8143 (N_8143,N_5393,N_5037);
and U8144 (N_8144,N_5511,N_6109);
nor U8145 (N_8145,N_5482,N_5344);
xor U8146 (N_8146,N_5029,N_7035);
nor U8147 (N_8147,N_6061,N_6585);
or U8148 (N_8148,N_6444,N_6757);
or U8149 (N_8149,N_5573,N_7460);
nand U8150 (N_8150,N_6588,N_7116);
and U8151 (N_8151,N_7010,N_5426);
and U8152 (N_8152,N_5753,N_6707);
nor U8153 (N_8153,N_6670,N_6937);
or U8154 (N_8154,N_7379,N_6933);
nand U8155 (N_8155,N_5849,N_6597);
nand U8156 (N_8156,N_5940,N_7063);
or U8157 (N_8157,N_5576,N_5909);
nand U8158 (N_8158,N_7032,N_7153);
and U8159 (N_8159,N_7388,N_5164);
and U8160 (N_8160,N_5973,N_5041);
nor U8161 (N_8161,N_5117,N_7350);
nor U8162 (N_8162,N_7049,N_6074);
or U8163 (N_8163,N_5912,N_5868);
nand U8164 (N_8164,N_6613,N_5409);
or U8165 (N_8165,N_7274,N_5220);
and U8166 (N_8166,N_5434,N_6112);
or U8167 (N_8167,N_7290,N_6768);
and U8168 (N_8168,N_7408,N_5648);
or U8169 (N_8169,N_6682,N_5523);
and U8170 (N_8170,N_7171,N_7433);
and U8171 (N_8171,N_6976,N_7473);
nand U8172 (N_8172,N_7046,N_6880);
nand U8173 (N_8173,N_5991,N_5017);
or U8174 (N_8174,N_6471,N_7495);
or U8175 (N_8175,N_5984,N_6951);
nand U8176 (N_8176,N_6972,N_5558);
nand U8177 (N_8177,N_5469,N_5925);
or U8178 (N_8178,N_6451,N_5996);
or U8179 (N_8179,N_6321,N_6831);
and U8180 (N_8180,N_5346,N_7377);
or U8181 (N_8181,N_5368,N_5147);
nand U8182 (N_8182,N_5038,N_6185);
or U8183 (N_8183,N_6565,N_5133);
nor U8184 (N_8184,N_7216,N_6874);
nand U8185 (N_8185,N_5628,N_6694);
nor U8186 (N_8186,N_5565,N_7310);
and U8187 (N_8187,N_7256,N_5224);
xnor U8188 (N_8188,N_5392,N_5772);
or U8189 (N_8189,N_5348,N_6516);
nand U8190 (N_8190,N_5877,N_7067);
nand U8191 (N_8191,N_6476,N_6313);
nor U8192 (N_8192,N_6182,N_5144);
nor U8193 (N_8193,N_5238,N_7491);
nor U8194 (N_8194,N_5824,N_6119);
or U8195 (N_8195,N_6895,N_7427);
nand U8196 (N_8196,N_7136,N_6489);
or U8197 (N_8197,N_6131,N_5356);
or U8198 (N_8198,N_7425,N_5404);
and U8199 (N_8199,N_7137,N_7409);
and U8200 (N_8200,N_6778,N_5608);
nor U8201 (N_8201,N_5470,N_6290);
nor U8202 (N_8202,N_7149,N_5294);
nor U8203 (N_8203,N_5828,N_5116);
or U8204 (N_8204,N_5740,N_5223);
or U8205 (N_8205,N_6472,N_6233);
nand U8206 (N_8206,N_5003,N_5175);
nor U8207 (N_8207,N_6931,N_5188);
nand U8208 (N_8208,N_7084,N_5590);
nor U8209 (N_8209,N_5859,N_5463);
nand U8210 (N_8210,N_6878,N_7109);
nor U8211 (N_8211,N_7172,N_5900);
nand U8212 (N_8212,N_6051,N_5787);
nand U8213 (N_8213,N_5689,N_5398);
nor U8214 (N_8214,N_5358,N_5207);
nor U8215 (N_8215,N_5995,N_5412);
or U8216 (N_8216,N_6715,N_6320);
nor U8217 (N_8217,N_6005,N_6106);
or U8218 (N_8218,N_6915,N_6135);
nand U8219 (N_8219,N_6488,N_6689);
nor U8220 (N_8220,N_5411,N_6116);
nand U8221 (N_8221,N_6870,N_6771);
or U8222 (N_8222,N_5495,N_6943);
nand U8223 (N_8223,N_7249,N_6553);
nand U8224 (N_8224,N_7320,N_6861);
nor U8225 (N_8225,N_7258,N_6611);
nand U8226 (N_8226,N_5771,N_7037);
and U8227 (N_8227,N_7393,N_7266);
or U8228 (N_8228,N_5496,N_5678);
nand U8229 (N_8229,N_6048,N_7180);
nand U8230 (N_8230,N_5011,N_5480);
nor U8231 (N_8231,N_5112,N_6420);
nand U8232 (N_8232,N_5168,N_6776);
nand U8233 (N_8233,N_5120,N_6604);
or U8234 (N_8234,N_7148,N_6981);
nor U8235 (N_8235,N_6583,N_5560);
and U8236 (N_8236,N_6065,N_6273);
nor U8237 (N_8237,N_7381,N_7181);
and U8238 (N_8238,N_6262,N_6491);
or U8239 (N_8239,N_6646,N_5723);
nand U8240 (N_8240,N_5923,N_6432);
nand U8241 (N_8241,N_6663,N_5988);
nor U8242 (N_8242,N_5546,N_5645);
or U8243 (N_8243,N_6964,N_5818);
nor U8244 (N_8244,N_5788,N_7045);
nand U8245 (N_8245,N_6966,N_5475);
nand U8246 (N_8246,N_6424,N_6950);
and U8247 (N_8247,N_6841,N_7459);
or U8248 (N_8248,N_6624,N_5669);
or U8249 (N_8249,N_7189,N_6938);
nor U8250 (N_8250,N_5707,N_5066);
or U8251 (N_8251,N_5671,N_5769);
or U8252 (N_8252,N_5453,N_7365);
nand U8253 (N_8253,N_6019,N_5385);
or U8254 (N_8254,N_7077,N_6551);
or U8255 (N_8255,N_7270,N_7110);
nand U8256 (N_8256,N_5564,N_7383);
nor U8257 (N_8257,N_7041,N_7260);
and U8258 (N_8258,N_6561,N_7275);
nand U8259 (N_8259,N_5551,N_6868);
and U8260 (N_8260,N_5975,N_5150);
and U8261 (N_8261,N_6054,N_6708);
nor U8262 (N_8262,N_5115,N_7465);
nor U8263 (N_8263,N_7038,N_6309);
or U8264 (N_8264,N_7065,N_5883);
nand U8265 (N_8265,N_7424,N_7173);
and U8266 (N_8266,N_5508,N_6337);
nor U8267 (N_8267,N_7396,N_5809);
or U8268 (N_8268,N_6110,N_5935);
or U8269 (N_8269,N_6760,N_5383);
nand U8270 (N_8270,N_6093,N_5189);
nor U8271 (N_8271,N_5812,N_5288);
nand U8272 (N_8272,N_5430,N_6509);
and U8273 (N_8273,N_5682,N_7092);
and U8274 (N_8274,N_5193,N_5204);
nand U8275 (N_8275,N_5105,N_7335);
nor U8276 (N_8276,N_5820,N_6165);
nor U8277 (N_8277,N_6748,N_7329);
and U8278 (N_8278,N_6889,N_5644);
nor U8279 (N_8279,N_7140,N_6360);
nor U8280 (N_8280,N_6965,N_6834);
nand U8281 (N_8281,N_5810,N_6383);
or U8282 (N_8282,N_6780,N_7170);
nand U8283 (N_8283,N_5186,N_5498);
nand U8284 (N_8284,N_6826,N_6890);
and U8285 (N_8285,N_5280,N_6803);
or U8286 (N_8286,N_6733,N_7302);
nand U8287 (N_8287,N_5185,N_7246);
nand U8288 (N_8288,N_5209,N_6853);
and U8289 (N_8289,N_5438,N_5665);
or U8290 (N_8290,N_5794,N_7315);
nand U8291 (N_8291,N_7481,N_7429);
nor U8292 (N_8292,N_6186,N_5355);
nand U8293 (N_8293,N_7430,N_5023);
nor U8294 (N_8294,N_5592,N_6840);
nand U8295 (N_8295,N_6521,N_6647);
nor U8296 (N_8296,N_5773,N_6210);
or U8297 (N_8297,N_6080,N_6577);
nand U8298 (N_8298,N_5597,N_7389);
and U8299 (N_8299,N_5004,N_5229);
or U8300 (N_8300,N_6508,N_7252);
or U8301 (N_8301,N_6272,N_5898);
and U8302 (N_8302,N_6633,N_5153);
and U8303 (N_8303,N_6975,N_7416);
and U8304 (N_8304,N_7471,N_5921);
nand U8305 (N_8305,N_6076,N_5870);
or U8306 (N_8306,N_6800,N_6664);
nor U8307 (N_8307,N_5722,N_6924);
nand U8308 (N_8308,N_5418,N_5553);
or U8309 (N_8309,N_6452,N_5367);
and U8310 (N_8310,N_5370,N_6062);
or U8311 (N_8311,N_7442,N_5025);
nand U8312 (N_8312,N_5607,N_5778);
nand U8313 (N_8313,N_7207,N_6085);
nand U8314 (N_8314,N_5680,N_5073);
and U8315 (N_8315,N_6187,N_7021);
nor U8316 (N_8316,N_6910,N_5673);
nand U8317 (N_8317,N_5012,N_6973);
nor U8318 (N_8318,N_5572,N_6230);
nor U8319 (N_8319,N_5749,N_5616);
and U8320 (N_8320,N_7107,N_5316);
and U8321 (N_8321,N_6685,N_6193);
and U8322 (N_8322,N_5710,N_5594);
nand U8323 (N_8323,N_7234,N_6267);
and U8324 (N_8324,N_5433,N_5559);
nand U8325 (N_8325,N_6475,N_7241);
nand U8326 (N_8326,N_6094,N_5906);
nor U8327 (N_8327,N_5544,N_6300);
or U8328 (N_8328,N_6384,N_7039);
or U8329 (N_8329,N_5436,N_7490);
or U8330 (N_8330,N_5699,N_7487);
nor U8331 (N_8331,N_5978,N_5177);
and U8332 (N_8332,N_6517,N_5047);
nand U8333 (N_8333,N_6614,N_6374);
or U8334 (N_8334,N_7185,N_6435);
nor U8335 (N_8335,N_6483,N_5951);
and U8336 (N_8336,N_6361,N_5985);
or U8337 (N_8337,N_5672,N_6350);
and U8338 (N_8338,N_5293,N_6809);
and U8339 (N_8339,N_5123,N_5384);
or U8340 (N_8340,N_5127,N_6038);
nor U8341 (N_8341,N_7205,N_5471);
or U8342 (N_8342,N_5297,N_7418);
or U8343 (N_8343,N_6306,N_7387);
nor U8344 (N_8344,N_7330,N_5513);
nor U8345 (N_8345,N_6598,N_7019);
nor U8346 (N_8346,N_7298,N_6507);
nand U8347 (N_8347,N_6169,N_5072);
or U8348 (N_8348,N_7231,N_6480);
nor U8349 (N_8349,N_5088,N_6045);
nor U8350 (N_8350,N_7078,N_6945);
or U8351 (N_8351,N_5567,N_7401);
nand U8352 (N_8352,N_5990,N_7251);
nor U8353 (N_8353,N_5052,N_6301);
nand U8354 (N_8354,N_7036,N_6200);
nand U8355 (N_8355,N_7384,N_7031);
nand U8356 (N_8356,N_5035,N_7356);
and U8357 (N_8357,N_6603,N_6705);
nor U8358 (N_8358,N_7468,N_7446);
or U8359 (N_8359,N_6990,N_5312);
nand U8360 (N_8360,N_6398,N_7394);
nor U8361 (N_8361,N_6334,N_6235);
and U8362 (N_8362,N_5027,N_6987);
nor U8363 (N_8363,N_5727,N_6278);
nor U8364 (N_8364,N_6765,N_5524);
xnor U8365 (N_8365,N_6815,N_6866);
and U8366 (N_8366,N_6279,N_5711);
and U8367 (N_8367,N_5237,N_6820);
nor U8368 (N_8368,N_5837,N_5698);
nor U8369 (N_8369,N_5520,N_7178);
nor U8370 (N_8370,N_6292,N_7198);
or U8371 (N_8371,N_5948,N_6862);
nor U8372 (N_8372,N_5322,N_5347);
nand U8373 (N_8373,N_6580,N_6648);
and U8374 (N_8374,N_5579,N_6571);
nor U8375 (N_8375,N_5016,N_6686);
nor U8376 (N_8376,N_5578,N_5097);
xor U8377 (N_8377,N_7121,N_5143);
and U8378 (N_8378,N_6227,N_5181);
or U8379 (N_8379,N_6056,N_6295);
nand U8380 (N_8380,N_5946,N_6539);
and U8381 (N_8381,N_5832,N_7081);
and U8382 (N_8382,N_6698,N_6754);
and U8383 (N_8383,N_6415,N_5493);
nor U8384 (N_8384,N_7326,N_6084);
nand U8385 (N_8385,N_5917,N_5374);
or U8386 (N_8386,N_5444,N_5765);
nor U8387 (N_8387,N_6202,N_5098);
nand U8388 (N_8388,N_5476,N_6954);
nand U8389 (N_8389,N_6559,N_6712);
and U8390 (N_8390,N_5821,N_5386);
nand U8391 (N_8391,N_6532,N_5371);
and U8392 (N_8392,N_5998,N_5899);
nor U8393 (N_8393,N_5450,N_5737);
nor U8394 (N_8394,N_6674,N_5541);
nor U8395 (N_8395,N_5627,N_5872);
or U8396 (N_8396,N_6653,N_7406);
nor U8397 (N_8397,N_6204,N_6761);
or U8398 (N_8398,N_5896,N_5919);
or U8399 (N_8399,N_6556,N_5649);
or U8400 (N_8400,N_6907,N_6639);
or U8401 (N_8401,N_6340,N_5854);
nand U8402 (N_8402,N_6838,N_6035);
or U8403 (N_8403,N_7435,N_6351);
nor U8404 (N_8404,N_5212,N_5631);
and U8405 (N_8405,N_5992,N_5192);
or U8406 (N_8406,N_5887,N_5623);
or U8407 (N_8407,N_7068,N_5813);
or U8408 (N_8408,N_5876,N_5884);
nor U8409 (N_8409,N_6006,N_5890);
nor U8410 (N_8410,N_6709,N_6117);
or U8411 (N_8411,N_5703,N_5545);
and U8412 (N_8412,N_5165,N_5685);
nand U8413 (N_8413,N_5094,N_6385);
or U8414 (N_8414,N_6887,N_5439);
nand U8415 (N_8415,N_7464,N_5394);
nand U8416 (N_8416,N_5532,N_7407);
nor U8417 (N_8417,N_5391,N_7373);
or U8418 (N_8418,N_6610,N_7071);
nand U8419 (N_8419,N_7265,N_5697);
nand U8420 (N_8420,N_5604,N_6746);
and U8421 (N_8421,N_5767,N_6102);
and U8422 (N_8422,N_6121,N_6289);
xnor U8423 (N_8423,N_6390,N_6425);
or U8424 (N_8424,N_6123,N_5403);
nand U8425 (N_8425,N_6462,N_5273);
nand U8426 (N_8426,N_7059,N_6626);
and U8427 (N_8427,N_5506,N_7294);
nand U8428 (N_8428,N_6942,N_6284);
or U8429 (N_8429,N_5518,N_6353);
nor U8430 (N_8430,N_5639,N_6103);
or U8431 (N_8431,N_7278,N_6438);
nor U8432 (N_8432,N_7303,N_7194);
and U8433 (N_8433,N_6958,N_5920);
nand U8434 (N_8434,N_7203,N_6596);
nor U8435 (N_8435,N_7126,N_7324);
nor U8436 (N_8436,N_7056,N_6644);
nor U8437 (N_8437,N_6534,N_5640);
nand U8438 (N_8438,N_5793,N_5020);
nor U8439 (N_8439,N_5933,N_7319);
and U8440 (N_8440,N_7292,N_5642);
nor U8441 (N_8441,N_7263,N_7201);
nand U8442 (N_8442,N_7130,N_7238);
and U8443 (N_8443,N_7338,N_6617);
nand U8444 (N_8444,N_6528,N_6364);
or U8445 (N_8445,N_6311,N_6269);
or U8446 (N_8446,N_7202,N_7269);
or U8447 (N_8447,N_6011,N_5504);
or U8448 (N_8448,N_5045,N_5786);
or U8449 (N_8449,N_5255,N_7218);
or U8450 (N_8450,N_6282,N_7143);
nor U8451 (N_8451,N_6032,N_6082);
or U8452 (N_8452,N_7212,N_7325);
or U8453 (N_8453,N_5354,N_7028);
nand U8454 (N_8454,N_7222,N_6851);
nand U8455 (N_8455,N_6469,N_6378);
and U8456 (N_8456,N_5729,N_6785);
nor U8457 (N_8457,N_6522,N_7070);
nor U8458 (N_8458,N_5303,N_6007);
and U8459 (N_8459,N_5662,N_5582);
and U8460 (N_8460,N_6797,N_6755);
nand U8461 (N_8461,N_6857,N_7210);
nor U8462 (N_8462,N_6344,N_6804);
nor U8463 (N_8463,N_6181,N_6732);
xnor U8464 (N_8464,N_5610,N_7489);
and U8465 (N_8465,N_5326,N_6541);
or U8466 (N_8466,N_6317,N_5656);
nor U8467 (N_8467,N_6373,N_5015);
nand U8468 (N_8468,N_7114,N_6879);
and U8469 (N_8469,N_7498,N_6087);
or U8470 (N_8470,N_6013,N_5107);
nor U8471 (N_8471,N_6014,N_5952);
nand U8472 (N_8472,N_6454,N_5655);
or U8473 (N_8473,N_7415,N_5750);
nand U8474 (N_8474,N_7431,N_6837);
and U8475 (N_8475,N_5363,N_6620);
and U8476 (N_8476,N_6691,N_6399);
nor U8477 (N_8477,N_5034,N_6040);
nor U8478 (N_8478,N_7309,N_6601);
and U8479 (N_8479,N_7286,N_5171);
and U8480 (N_8480,N_5719,N_6440);
and U8481 (N_8481,N_6150,N_6346);
nand U8482 (N_8482,N_6241,N_6209);
nand U8483 (N_8483,N_6801,N_6263);
nor U8484 (N_8484,N_5510,N_6989);
nor U8485 (N_8485,N_7282,N_5858);
nand U8486 (N_8486,N_5406,N_7196);
nor U8487 (N_8487,N_5997,N_6137);
and U8488 (N_8488,N_6690,N_5865);
nand U8489 (N_8489,N_5713,N_5397);
and U8490 (N_8490,N_6696,N_7448);
and U8491 (N_8491,N_5474,N_6900);
nor U8492 (N_8492,N_7486,N_6268);
nand U8493 (N_8493,N_5539,N_5955);
nor U8494 (N_8494,N_6650,N_6134);
nor U8495 (N_8495,N_5485,N_6177);
or U8496 (N_8496,N_7466,N_5944);
nand U8497 (N_8497,N_5913,N_6499);
and U8498 (N_8498,N_6753,N_7245);
and U8499 (N_8499,N_5084,N_6231);
and U8500 (N_8500,N_5693,N_5547);
nand U8501 (N_8501,N_5606,N_5947);
and U8502 (N_8502,N_5874,N_6558);
or U8503 (N_8503,N_6858,N_5779);
nand U8504 (N_8504,N_6612,N_5535);
and U8505 (N_8505,N_6572,N_5152);
nand U8506 (N_8506,N_6994,N_7455);
or U8507 (N_8507,N_5804,N_7161);
nand U8508 (N_8508,N_6531,N_7232);
or U8509 (N_8509,N_5291,N_5871);
nand U8510 (N_8510,N_6557,N_6667);
nor U8511 (N_8511,N_5613,N_6152);
nor U8512 (N_8512,N_5835,N_6527);
nor U8513 (N_8513,N_6720,N_6519);
nor U8514 (N_8514,N_6657,N_5054);
nor U8515 (N_8515,N_6717,N_5605);
or U8516 (N_8516,N_5569,N_5187);
nand U8517 (N_8517,N_5895,N_6457);
nor U8518 (N_8518,N_5307,N_6744);
and U8519 (N_8519,N_5967,N_5227);
nand U8520 (N_8520,N_5725,N_7268);
or U8521 (N_8521,N_5099,N_5085);
nor U8522 (N_8522,N_6706,N_6957);
or U8523 (N_8523,N_5962,N_5808);
and U8524 (N_8524,N_5885,N_5093);
nor U8525 (N_8525,N_5976,N_6327);
nand U8526 (N_8526,N_5958,N_6243);
or U8527 (N_8527,N_6550,N_7162);
and U8528 (N_8528,N_6749,N_6777);
or U8529 (N_8529,N_5538,N_5893);
nand U8530 (N_8530,N_6991,N_6606);
nor U8531 (N_8531,N_5456,N_6078);
nand U8532 (N_8532,N_5415,N_6304);
nand U8533 (N_8533,N_7352,N_6389);
nor U8534 (N_8534,N_7213,N_5831);
and U8535 (N_8535,N_7432,N_7104);
or U8536 (N_8536,N_5264,N_6782);
nand U8537 (N_8537,N_5423,N_5336);
or U8538 (N_8538,N_5390,N_6090);
nand U8539 (N_8539,N_7244,N_6297);
nand U8540 (N_8540,N_7312,N_6447);
and U8541 (N_8541,N_7304,N_6999);
nor U8542 (N_8542,N_6734,N_5334);
nor U8543 (N_8543,N_7404,N_6042);
and U8544 (N_8544,N_6368,N_6576);
xor U8545 (N_8545,N_5008,N_5101);
nor U8546 (N_8546,N_6031,N_5062);
nor U8547 (N_8547,N_7052,N_7135);
nand U8548 (N_8548,N_6312,N_6923);
nand U8549 (N_8549,N_5783,N_6848);
nor U8550 (N_8550,N_6003,N_6830);
or U8551 (N_8551,N_6400,N_5170);
or U8552 (N_8552,N_6703,N_6906);
nand U8553 (N_8553,N_6668,N_6566);
or U8554 (N_8554,N_6322,N_6672);
nor U8555 (N_8555,N_6852,N_5999);
nand U8556 (N_8556,N_5903,N_6318);
or U8557 (N_8557,N_5914,N_5467);
nand U8558 (N_8558,N_5109,N_6823);
or U8559 (N_8559,N_5129,N_7462);
or U8560 (N_8560,N_5894,N_6173);
nor U8561 (N_8561,N_5963,N_6788);
nand U8562 (N_8562,N_5641,N_6548);
or U8563 (N_8563,N_5059,N_5945);
nand U8564 (N_8564,N_6458,N_7233);
or U8565 (N_8565,N_7182,N_6030);
nor U8566 (N_8566,N_5472,N_7272);
and U8567 (N_8567,N_6926,N_5602);
nand U8568 (N_8568,N_5542,N_5033);
nor U8569 (N_8569,N_6833,N_6935);
or U8570 (N_8570,N_7060,N_5103);
nand U8571 (N_8571,N_6114,N_5026);
nor U8572 (N_8572,N_5802,N_6883);
xnor U8573 (N_8573,N_7440,N_6495);
nor U8574 (N_8574,N_7204,N_7358);
or U8575 (N_8575,N_7072,N_6496);
and U8576 (N_8576,N_6751,N_6984);
nor U8577 (N_8577,N_7111,N_5139);
or U8578 (N_8578,N_7395,N_5014);
and U8579 (N_8579,N_5036,N_5376);
and U8580 (N_8580,N_7083,N_6581);
and U8581 (N_8581,N_5388,N_6589);
nand U8582 (N_8582,N_5420,N_7112);
and U8583 (N_8583,N_5124,N_5796);
xor U8584 (N_8584,N_7273,N_7167);
and U8585 (N_8585,N_5490,N_5158);
and U8586 (N_8586,N_5694,N_6176);
nor U8587 (N_8587,N_6168,N_7165);
nor U8588 (N_8588,N_5833,N_6126);
nor U8589 (N_8589,N_5005,N_7096);
nor U8590 (N_8590,N_6348,N_6329);
nor U8591 (N_8591,N_5879,N_5676);
nor U8592 (N_8592,N_6766,N_6153);
nor U8593 (N_8593,N_5800,N_7175);
and U8594 (N_8594,N_6980,N_5593);
or U8595 (N_8595,N_6178,N_6012);
and U8596 (N_8596,N_5891,N_6408);
and U8597 (N_8597,N_5236,N_6730);
or U8598 (N_8598,N_6627,N_5263);
nand U8599 (N_8599,N_5728,N_6764);
nor U8600 (N_8600,N_6854,N_5584);
or U8601 (N_8601,N_6638,N_5173);
or U8602 (N_8602,N_6658,N_6584);
nor U8603 (N_8603,N_5437,N_7262);
and U8604 (N_8604,N_5549,N_5581);
or U8605 (N_8605,N_5341,N_5908);
nor U8606 (N_8606,N_5622,N_6214);
and U8607 (N_8607,N_5250,N_6533);
and U8608 (N_8608,N_7371,N_6555);
or U8609 (N_8609,N_6723,N_5657);
nor U8610 (N_8610,N_6925,N_6914);
and U8611 (N_8611,N_7426,N_5427);
nor U8612 (N_8612,N_7001,N_5843);
nand U8613 (N_8613,N_6232,N_5335);
or U8614 (N_8614,N_6513,N_5851);
nor U8615 (N_8615,N_7061,N_5201);
nand U8616 (N_8616,N_6004,N_6918);
and U8617 (N_8617,N_7318,N_7367);
and U8618 (N_8618,N_6071,N_7125);
or U8619 (N_8619,N_7006,N_6922);
or U8620 (N_8620,N_5857,N_7193);
or U8621 (N_8621,N_7025,N_6017);
nand U8622 (N_8622,N_7479,N_7018);
and U8623 (N_8623,N_7445,N_5137);
nand U8624 (N_8624,N_5200,N_5468);
nand U8625 (N_8625,N_5135,N_5762);
nand U8626 (N_8626,N_6609,N_6816);
nand U8627 (N_8627,N_5795,N_5557);
or U8628 (N_8628,N_6122,N_6842);
nor U8629 (N_8629,N_5817,N_5974);
nor U8630 (N_8630,N_6310,N_5429);
nand U8631 (N_8631,N_5670,N_6904);
nand U8632 (N_8632,N_6502,N_6919);
or U8633 (N_8633,N_7098,N_6787);
nor U8634 (N_8634,N_6632,N_5932);
nor U8635 (N_8635,N_5658,N_5668);
or U8636 (N_8636,N_6784,N_5537);
and U8637 (N_8637,N_5421,N_5260);
and U8638 (N_8638,N_5867,N_5735);
nand U8639 (N_8639,N_5353,N_6101);
and U8640 (N_8640,N_7014,N_6796);
xnor U8641 (N_8641,N_6552,N_6593);
nand U8642 (N_8642,N_6050,N_6520);
and U8643 (N_8643,N_5799,N_6133);
nand U8644 (N_8644,N_6439,N_7200);
nor U8645 (N_8645,N_7030,N_6500);
nand U8646 (N_8646,N_7094,N_5611);
nand U8647 (N_8647,N_6688,N_5977);
nor U8648 (N_8648,N_7118,N_5683);
nand U8649 (N_8649,N_6956,N_5108);
nand U8650 (N_8650,N_6025,N_6010);
nand U8651 (N_8651,N_5221,N_5230);
or U8652 (N_8652,N_6154,N_6886);
or U8653 (N_8653,N_5304,N_5916);
nand U8654 (N_8654,N_5501,N_5104);
or U8655 (N_8655,N_6579,N_5329);
and U8656 (N_8656,N_6665,N_6896);
nand U8657 (N_8657,N_6225,N_7398);
nand U8658 (N_8658,N_7301,N_5169);
nor U8659 (N_8659,N_5617,N_7105);
nand U8660 (N_8660,N_7313,N_6738);
nor U8661 (N_8661,N_6144,N_7015);
nor U8662 (N_8662,N_6203,N_6022);
nor U8663 (N_8663,N_5462,N_5156);
nand U8664 (N_8664,N_5092,N_7091);
nor U8665 (N_8665,N_7285,N_6538);
nand U8666 (N_8666,N_7156,N_6898);
or U8667 (N_8667,N_5447,N_5692);
nand U8668 (N_8668,N_6115,N_6414);
and U8669 (N_8669,N_5503,N_6721);
nand U8670 (N_8670,N_5869,N_5377);
nor U8671 (N_8671,N_5145,N_6377);
nand U8672 (N_8672,N_6463,N_6873);
nor U8673 (N_8673,N_5022,N_7043);
or U8674 (N_8674,N_6092,N_5739);
nand U8675 (N_8675,N_5815,N_5803);
nor U8676 (N_8676,N_5756,N_6336);
and U8677 (N_8677,N_7220,N_5292);
or U8678 (N_8678,N_7197,N_5372);
nor U8679 (N_8679,N_6849,N_5276);
and U8680 (N_8680,N_6008,N_7485);
and U8681 (N_8681,N_6684,N_5507);
or U8682 (N_8682,N_6967,N_7297);
nand U8683 (N_8683,N_6029,N_6828);
nand U8684 (N_8684,N_5888,N_5321);
and U8685 (N_8685,N_6332,N_6184);
nand U8686 (N_8686,N_5521,N_6430);
and U8687 (N_8687,N_7004,N_5637);
or U8688 (N_8688,N_5235,N_5960);
and U8689 (N_8689,N_6482,N_6157);
or U8690 (N_8690,N_5734,N_6393);
nor U8691 (N_8691,N_6283,N_6338);
nor U8692 (N_8692,N_6540,N_5121);
or U8693 (N_8693,N_7017,N_5484);
nor U8694 (N_8694,N_6129,N_7026);
xor U8695 (N_8695,N_6410,N_5929);
nand U8696 (N_8696,N_5738,N_5968);
nor U8697 (N_8697,N_6511,N_7186);
or U8698 (N_8698,N_6568,N_7343);
nand U8699 (N_8699,N_6201,N_7488);
nand U8700 (N_8700,N_7240,N_5841);
nor U8701 (N_8701,N_5110,N_6970);
nor U8702 (N_8702,N_6161,N_6669);
nand U8703 (N_8703,N_6039,N_6860);
nand U8704 (N_8704,N_5048,N_7128);
and U8705 (N_8705,N_5886,N_5405);
nand U8706 (N_8706,N_7044,N_5814);
or U8707 (N_8707,N_6729,N_7454);
nor U8708 (N_8708,N_6125,N_6434);
nand U8709 (N_8709,N_7374,N_6745);
nor U8710 (N_8710,N_7247,N_6431);
nor U8711 (N_8711,N_5709,N_5926);
nand U8712 (N_8712,N_6921,N_6602);
nor U8713 (N_8713,N_7411,N_5432);
and U8714 (N_8714,N_5281,N_5502);
nand U8715 (N_8715,N_6813,N_6960);
or U8716 (N_8716,N_6714,N_5930);
or U8717 (N_8717,N_6086,N_5166);
or U8718 (N_8718,N_7420,N_6299);
nor U8719 (N_8719,N_6260,N_6643);
or U8720 (N_8720,N_6275,N_6635);
nand U8721 (N_8721,N_5317,N_6731);
nand U8722 (N_8722,N_5058,N_5801);
nand U8723 (N_8723,N_5241,N_5302);
nand U8724 (N_8724,N_6484,N_6512);
and U8725 (N_8725,N_6537,N_7155);
nand U8726 (N_8726,N_6315,N_7138);
nor U8727 (N_8727,N_7277,N_7163);
or U8728 (N_8728,N_6892,N_5130);
nand U8729 (N_8729,N_6172,N_5216);
or U8730 (N_8730,N_6354,N_6380);
or U8731 (N_8731,N_5943,N_6305);
and U8732 (N_8732,N_5309,N_6783);
and U8733 (N_8733,N_6920,N_5543);
nand U8734 (N_8734,N_6817,N_7076);
and U8735 (N_8735,N_6171,N_6036);
and U8736 (N_8736,N_5517,N_6127);
and U8737 (N_8737,N_5002,N_5111);
nand U8738 (N_8738,N_6073,N_6199);
or U8739 (N_8739,N_5585,N_5183);
or U8740 (N_8740,N_7413,N_6485);
or U8741 (N_8741,N_5844,N_6524);
and U8742 (N_8742,N_6403,N_7385);
nor U8743 (N_8743,N_6098,N_5202);
nand U8744 (N_8744,N_5323,N_6829);
and U8745 (N_8745,N_6735,N_5855);
or U8746 (N_8746,N_5754,N_6024);
nand U8747 (N_8747,N_7066,N_6274);
or U8748 (N_8748,N_6806,N_5550);
nand U8749 (N_8749,N_5360,N_5006);
nand U8750 (N_8750,N_5747,N_6473);
and U8751 (N_8751,N_7348,N_7257);
or U8752 (N_8752,N_6228,N_5841);
or U8753 (N_8753,N_6992,N_6220);
or U8754 (N_8754,N_5577,N_6230);
nand U8755 (N_8755,N_7415,N_5319);
nor U8756 (N_8756,N_5980,N_6476);
nor U8757 (N_8757,N_6030,N_5652);
nand U8758 (N_8758,N_7264,N_6230);
and U8759 (N_8759,N_6035,N_6759);
and U8760 (N_8760,N_6175,N_6768);
nand U8761 (N_8761,N_6660,N_7320);
or U8762 (N_8762,N_6117,N_5495);
or U8763 (N_8763,N_6893,N_5717);
or U8764 (N_8764,N_6089,N_5764);
xnor U8765 (N_8765,N_6641,N_6721);
and U8766 (N_8766,N_6341,N_6900);
nand U8767 (N_8767,N_5279,N_6857);
nor U8768 (N_8768,N_5338,N_5082);
and U8769 (N_8769,N_5970,N_7281);
nand U8770 (N_8770,N_5590,N_5437);
nor U8771 (N_8771,N_7003,N_7314);
nor U8772 (N_8772,N_6926,N_5429);
and U8773 (N_8773,N_5645,N_7037);
or U8774 (N_8774,N_5325,N_5868);
or U8775 (N_8775,N_5349,N_5736);
nand U8776 (N_8776,N_5291,N_6412);
nor U8777 (N_8777,N_5793,N_5609);
and U8778 (N_8778,N_6519,N_7346);
nor U8779 (N_8779,N_6436,N_6424);
nor U8780 (N_8780,N_6404,N_5770);
or U8781 (N_8781,N_5280,N_5517);
or U8782 (N_8782,N_5586,N_5464);
nor U8783 (N_8783,N_7081,N_7379);
and U8784 (N_8784,N_6984,N_6799);
and U8785 (N_8785,N_6955,N_5888);
nand U8786 (N_8786,N_7414,N_5799);
and U8787 (N_8787,N_5798,N_6024);
nor U8788 (N_8788,N_6700,N_7282);
or U8789 (N_8789,N_7127,N_6063);
and U8790 (N_8790,N_5224,N_6692);
nand U8791 (N_8791,N_7117,N_6996);
nor U8792 (N_8792,N_6129,N_7427);
nand U8793 (N_8793,N_5588,N_7271);
or U8794 (N_8794,N_6467,N_6952);
nor U8795 (N_8795,N_7443,N_6734);
or U8796 (N_8796,N_7380,N_5025);
or U8797 (N_8797,N_6276,N_6944);
nor U8798 (N_8798,N_5342,N_5756);
nand U8799 (N_8799,N_6580,N_7382);
or U8800 (N_8800,N_5485,N_6957);
and U8801 (N_8801,N_5884,N_6558);
and U8802 (N_8802,N_6228,N_6363);
or U8803 (N_8803,N_5014,N_5695);
nor U8804 (N_8804,N_6443,N_5661);
and U8805 (N_8805,N_7206,N_5497);
or U8806 (N_8806,N_6714,N_7438);
nor U8807 (N_8807,N_6601,N_5791);
nand U8808 (N_8808,N_6987,N_5017);
nor U8809 (N_8809,N_6150,N_5800);
and U8810 (N_8810,N_6218,N_6824);
nor U8811 (N_8811,N_5816,N_6432);
or U8812 (N_8812,N_6064,N_7307);
nand U8813 (N_8813,N_6057,N_5199);
or U8814 (N_8814,N_7205,N_5304);
nor U8815 (N_8815,N_5574,N_5939);
and U8816 (N_8816,N_7252,N_7185);
and U8817 (N_8817,N_5559,N_5011);
or U8818 (N_8818,N_5736,N_7184);
nor U8819 (N_8819,N_7154,N_6735);
nand U8820 (N_8820,N_5673,N_7290);
or U8821 (N_8821,N_7223,N_5053);
nand U8822 (N_8822,N_6342,N_7470);
or U8823 (N_8823,N_5834,N_6218);
nand U8824 (N_8824,N_6612,N_6804);
and U8825 (N_8825,N_6807,N_7080);
xnor U8826 (N_8826,N_5550,N_5651);
and U8827 (N_8827,N_6939,N_6109);
nor U8828 (N_8828,N_5878,N_5009);
or U8829 (N_8829,N_7009,N_7192);
and U8830 (N_8830,N_6419,N_6917);
nor U8831 (N_8831,N_6637,N_6710);
nand U8832 (N_8832,N_5458,N_5390);
and U8833 (N_8833,N_6920,N_6282);
nand U8834 (N_8834,N_5288,N_6513);
or U8835 (N_8835,N_6986,N_5296);
nand U8836 (N_8836,N_6831,N_7186);
nor U8837 (N_8837,N_6966,N_6186);
or U8838 (N_8838,N_6317,N_7091);
or U8839 (N_8839,N_5075,N_6349);
and U8840 (N_8840,N_6104,N_5806);
nor U8841 (N_8841,N_5051,N_6749);
nand U8842 (N_8842,N_5431,N_6576);
and U8843 (N_8843,N_5716,N_5621);
nand U8844 (N_8844,N_7053,N_7446);
nand U8845 (N_8845,N_7023,N_5605);
nor U8846 (N_8846,N_6816,N_6697);
and U8847 (N_8847,N_6781,N_5453);
or U8848 (N_8848,N_5484,N_5578);
or U8849 (N_8849,N_5565,N_6344);
nor U8850 (N_8850,N_6086,N_6398);
and U8851 (N_8851,N_5054,N_5646);
or U8852 (N_8852,N_6329,N_5161);
nand U8853 (N_8853,N_7336,N_5313);
nor U8854 (N_8854,N_7411,N_5705);
or U8855 (N_8855,N_6304,N_5585);
and U8856 (N_8856,N_7339,N_7203);
nor U8857 (N_8857,N_5538,N_5757);
or U8858 (N_8858,N_5115,N_6449);
and U8859 (N_8859,N_5345,N_5966);
nand U8860 (N_8860,N_5094,N_6677);
nand U8861 (N_8861,N_6580,N_5307);
nand U8862 (N_8862,N_5777,N_6115);
nand U8863 (N_8863,N_7043,N_6085);
and U8864 (N_8864,N_6002,N_6237);
nor U8865 (N_8865,N_7497,N_6039);
nor U8866 (N_8866,N_6724,N_5492);
and U8867 (N_8867,N_6350,N_6351);
nor U8868 (N_8868,N_5751,N_6266);
nand U8869 (N_8869,N_6593,N_7066);
or U8870 (N_8870,N_7463,N_5994);
nand U8871 (N_8871,N_6924,N_5273);
and U8872 (N_8872,N_5602,N_5324);
or U8873 (N_8873,N_7273,N_6598);
and U8874 (N_8874,N_6743,N_5055);
and U8875 (N_8875,N_5625,N_7416);
or U8876 (N_8876,N_7378,N_6778);
nor U8877 (N_8877,N_6483,N_5220);
nor U8878 (N_8878,N_6474,N_6632);
or U8879 (N_8879,N_7047,N_6384);
and U8880 (N_8880,N_5481,N_6198);
nand U8881 (N_8881,N_6470,N_6245);
and U8882 (N_8882,N_5206,N_5494);
nor U8883 (N_8883,N_7215,N_6379);
and U8884 (N_8884,N_6048,N_5398);
and U8885 (N_8885,N_5917,N_6837);
nor U8886 (N_8886,N_5367,N_5259);
nand U8887 (N_8887,N_7168,N_7039);
or U8888 (N_8888,N_5423,N_6953);
and U8889 (N_8889,N_6175,N_6999);
and U8890 (N_8890,N_5721,N_7170);
and U8891 (N_8891,N_5045,N_6643);
nand U8892 (N_8892,N_7031,N_5370);
nand U8893 (N_8893,N_6192,N_6411);
nand U8894 (N_8894,N_6418,N_5489);
nand U8895 (N_8895,N_7334,N_7237);
or U8896 (N_8896,N_7310,N_6404);
nand U8897 (N_8897,N_6842,N_5996);
nor U8898 (N_8898,N_6078,N_5810);
nand U8899 (N_8899,N_7310,N_6072);
or U8900 (N_8900,N_5383,N_5400);
nor U8901 (N_8901,N_6366,N_7210);
nor U8902 (N_8902,N_7104,N_5464);
or U8903 (N_8903,N_5090,N_7457);
and U8904 (N_8904,N_6882,N_5523);
nor U8905 (N_8905,N_7030,N_6936);
and U8906 (N_8906,N_6985,N_7046);
or U8907 (N_8907,N_5479,N_7049);
or U8908 (N_8908,N_7223,N_7228);
or U8909 (N_8909,N_5985,N_5658);
nor U8910 (N_8910,N_5939,N_6460);
nand U8911 (N_8911,N_6960,N_6703);
or U8912 (N_8912,N_5008,N_6936);
nor U8913 (N_8913,N_5238,N_6437);
and U8914 (N_8914,N_5895,N_6777);
and U8915 (N_8915,N_5611,N_6802);
and U8916 (N_8916,N_5821,N_6142);
nand U8917 (N_8917,N_6031,N_6656);
or U8918 (N_8918,N_5771,N_7157);
nor U8919 (N_8919,N_6805,N_7083);
or U8920 (N_8920,N_5336,N_6438);
nor U8921 (N_8921,N_5527,N_6383);
nand U8922 (N_8922,N_5955,N_6417);
or U8923 (N_8923,N_6002,N_6583);
nand U8924 (N_8924,N_5393,N_6438);
and U8925 (N_8925,N_5769,N_5105);
and U8926 (N_8926,N_7467,N_6367);
or U8927 (N_8927,N_6385,N_6241);
and U8928 (N_8928,N_6414,N_6450);
and U8929 (N_8929,N_7431,N_5505);
nand U8930 (N_8930,N_7269,N_7374);
nand U8931 (N_8931,N_6659,N_6406);
nor U8932 (N_8932,N_5683,N_6083);
nor U8933 (N_8933,N_6569,N_6742);
nor U8934 (N_8934,N_5750,N_5486);
and U8935 (N_8935,N_6075,N_5080);
and U8936 (N_8936,N_6648,N_6292);
and U8937 (N_8937,N_6415,N_6356);
nor U8938 (N_8938,N_6594,N_7061);
nor U8939 (N_8939,N_5436,N_5275);
nand U8940 (N_8940,N_7414,N_6745);
nor U8941 (N_8941,N_5834,N_6821);
nor U8942 (N_8942,N_5204,N_7170);
or U8943 (N_8943,N_5694,N_5160);
and U8944 (N_8944,N_6593,N_6737);
nor U8945 (N_8945,N_5016,N_6271);
or U8946 (N_8946,N_5405,N_5369);
or U8947 (N_8947,N_6468,N_5877);
nor U8948 (N_8948,N_5683,N_7027);
nand U8949 (N_8949,N_5530,N_6676);
nor U8950 (N_8950,N_7095,N_6229);
and U8951 (N_8951,N_7221,N_6309);
or U8952 (N_8952,N_5319,N_6288);
nand U8953 (N_8953,N_7084,N_6881);
nand U8954 (N_8954,N_5702,N_5174);
nand U8955 (N_8955,N_7441,N_6209);
or U8956 (N_8956,N_7131,N_7349);
or U8957 (N_8957,N_6106,N_7172);
or U8958 (N_8958,N_5176,N_5828);
nor U8959 (N_8959,N_7180,N_7355);
or U8960 (N_8960,N_5552,N_6663);
or U8961 (N_8961,N_7272,N_6455);
nand U8962 (N_8962,N_6587,N_7471);
or U8963 (N_8963,N_7336,N_5617);
or U8964 (N_8964,N_6776,N_6171);
or U8965 (N_8965,N_5178,N_5716);
and U8966 (N_8966,N_7232,N_6481);
or U8967 (N_8967,N_5479,N_5441);
xor U8968 (N_8968,N_6601,N_5741);
nand U8969 (N_8969,N_5399,N_6131);
nor U8970 (N_8970,N_5031,N_5509);
and U8971 (N_8971,N_6423,N_5824);
nand U8972 (N_8972,N_6185,N_5461);
nor U8973 (N_8973,N_6091,N_6204);
or U8974 (N_8974,N_6316,N_6319);
or U8975 (N_8975,N_7426,N_5497);
and U8976 (N_8976,N_6900,N_7147);
and U8977 (N_8977,N_5785,N_5451);
and U8978 (N_8978,N_5819,N_6962);
nor U8979 (N_8979,N_5592,N_5506);
nand U8980 (N_8980,N_5725,N_7481);
nand U8981 (N_8981,N_5594,N_6193);
nor U8982 (N_8982,N_6682,N_5117);
nand U8983 (N_8983,N_7232,N_6930);
or U8984 (N_8984,N_6410,N_5215);
nor U8985 (N_8985,N_6968,N_6480);
nor U8986 (N_8986,N_7330,N_6106);
and U8987 (N_8987,N_6460,N_5146);
and U8988 (N_8988,N_5757,N_6830);
or U8989 (N_8989,N_7352,N_5990);
or U8990 (N_8990,N_6267,N_5188);
nor U8991 (N_8991,N_5812,N_5041);
nand U8992 (N_8992,N_5167,N_5928);
nor U8993 (N_8993,N_5060,N_7078);
or U8994 (N_8994,N_6122,N_6070);
or U8995 (N_8995,N_6620,N_6285);
nor U8996 (N_8996,N_6621,N_6537);
nor U8997 (N_8997,N_5796,N_5531);
or U8998 (N_8998,N_7466,N_6843);
nor U8999 (N_8999,N_6956,N_5341);
or U9000 (N_9000,N_7496,N_5596);
xnor U9001 (N_9001,N_6110,N_6876);
and U9002 (N_9002,N_6218,N_7338);
and U9003 (N_9003,N_5555,N_6230);
xnor U9004 (N_9004,N_6572,N_7459);
nor U9005 (N_9005,N_6960,N_5876);
or U9006 (N_9006,N_6868,N_5801);
and U9007 (N_9007,N_7070,N_6937);
nand U9008 (N_9008,N_5768,N_5880);
and U9009 (N_9009,N_5149,N_6459);
nor U9010 (N_9010,N_6108,N_7135);
nand U9011 (N_9011,N_5946,N_6088);
nor U9012 (N_9012,N_5724,N_5355);
nor U9013 (N_9013,N_5367,N_5570);
and U9014 (N_9014,N_6274,N_5597);
and U9015 (N_9015,N_5399,N_5970);
and U9016 (N_9016,N_5256,N_7260);
and U9017 (N_9017,N_6148,N_6265);
or U9018 (N_9018,N_5713,N_5576);
nor U9019 (N_9019,N_7089,N_5224);
or U9020 (N_9020,N_6815,N_5115);
nor U9021 (N_9021,N_5799,N_6298);
nand U9022 (N_9022,N_7342,N_6356);
or U9023 (N_9023,N_5194,N_6980);
nand U9024 (N_9024,N_6441,N_5921);
and U9025 (N_9025,N_5863,N_6234);
nor U9026 (N_9026,N_6672,N_6909);
nand U9027 (N_9027,N_6045,N_5356);
and U9028 (N_9028,N_6906,N_5510);
and U9029 (N_9029,N_5694,N_6524);
nor U9030 (N_9030,N_7310,N_7019);
nor U9031 (N_9031,N_6223,N_5234);
nand U9032 (N_9032,N_5862,N_6752);
nor U9033 (N_9033,N_5384,N_6396);
and U9034 (N_9034,N_6801,N_5339);
nor U9035 (N_9035,N_6291,N_7489);
and U9036 (N_9036,N_6115,N_5191);
nand U9037 (N_9037,N_7077,N_6727);
and U9038 (N_9038,N_6622,N_5617);
nor U9039 (N_9039,N_5070,N_6687);
or U9040 (N_9040,N_6444,N_6636);
or U9041 (N_9041,N_7251,N_7472);
xnor U9042 (N_9042,N_5649,N_6080);
nor U9043 (N_9043,N_5176,N_6373);
nor U9044 (N_9044,N_7432,N_7023);
or U9045 (N_9045,N_5355,N_6263);
nor U9046 (N_9046,N_6516,N_7197);
nand U9047 (N_9047,N_6767,N_7130);
nor U9048 (N_9048,N_5159,N_6718);
nor U9049 (N_9049,N_5163,N_6749);
and U9050 (N_9050,N_6799,N_5352);
xor U9051 (N_9051,N_6113,N_5826);
or U9052 (N_9052,N_5806,N_7147);
or U9053 (N_9053,N_6721,N_7255);
nor U9054 (N_9054,N_5196,N_5447);
or U9055 (N_9055,N_6046,N_5429);
or U9056 (N_9056,N_7069,N_6511);
and U9057 (N_9057,N_5047,N_5876);
and U9058 (N_9058,N_5103,N_7027);
and U9059 (N_9059,N_7262,N_7346);
or U9060 (N_9060,N_6387,N_7107);
nand U9061 (N_9061,N_6948,N_7215);
and U9062 (N_9062,N_5382,N_5596);
or U9063 (N_9063,N_6424,N_6681);
nand U9064 (N_9064,N_6746,N_6127);
and U9065 (N_9065,N_5879,N_7488);
or U9066 (N_9066,N_5358,N_5067);
nand U9067 (N_9067,N_5880,N_5478);
nand U9068 (N_9068,N_5200,N_5533);
nand U9069 (N_9069,N_7186,N_5398);
or U9070 (N_9070,N_6550,N_6947);
nor U9071 (N_9071,N_5074,N_6054);
and U9072 (N_9072,N_5627,N_5365);
nand U9073 (N_9073,N_5279,N_6619);
nor U9074 (N_9074,N_5629,N_6521);
nor U9075 (N_9075,N_6570,N_7461);
xnor U9076 (N_9076,N_6072,N_7069);
nand U9077 (N_9077,N_5014,N_5086);
or U9078 (N_9078,N_7311,N_6629);
and U9079 (N_9079,N_6946,N_5535);
or U9080 (N_9080,N_5704,N_7367);
and U9081 (N_9081,N_5622,N_6654);
nand U9082 (N_9082,N_6779,N_6586);
nor U9083 (N_9083,N_7115,N_6074);
nand U9084 (N_9084,N_5232,N_6491);
and U9085 (N_9085,N_5555,N_5720);
nand U9086 (N_9086,N_5707,N_5220);
and U9087 (N_9087,N_5131,N_6463);
and U9088 (N_9088,N_6297,N_6994);
or U9089 (N_9089,N_5641,N_7424);
nand U9090 (N_9090,N_7276,N_7185);
nand U9091 (N_9091,N_6239,N_6857);
or U9092 (N_9092,N_6272,N_7104);
and U9093 (N_9093,N_5370,N_5267);
or U9094 (N_9094,N_6783,N_6174);
nor U9095 (N_9095,N_5602,N_5747);
nor U9096 (N_9096,N_5148,N_6250);
or U9097 (N_9097,N_6688,N_7344);
nand U9098 (N_9098,N_7431,N_5356);
nand U9099 (N_9099,N_5637,N_5623);
and U9100 (N_9100,N_5348,N_7379);
nand U9101 (N_9101,N_6937,N_6921);
nor U9102 (N_9102,N_6004,N_6353);
nand U9103 (N_9103,N_7043,N_5208);
and U9104 (N_9104,N_6540,N_6610);
nor U9105 (N_9105,N_6470,N_5695);
or U9106 (N_9106,N_5765,N_6996);
nand U9107 (N_9107,N_6955,N_6732);
nand U9108 (N_9108,N_5178,N_7311);
and U9109 (N_9109,N_6485,N_7265);
nand U9110 (N_9110,N_5052,N_6090);
or U9111 (N_9111,N_7335,N_6231);
or U9112 (N_9112,N_5325,N_6619);
xnor U9113 (N_9113,N_5162,N_6697);
or U9114 (N_9114,N_5316,N_6237);
or U9115 (N_9115,N_6870,N_5931);
and U9116 (N_9116,N_7379,N_6419);
and U9117 (N_9117,N_5499,N_7297);
nand U9118 (N_9118,N_5926,N_6263);
or U9119 (N_9119,N_5159,N_5214);
nor U9120 (N_9120,N_6647,N_5213);
and U9121 (N_9121,N_7426,N_6332);
and U9122 (N_9122,N_5966,N_7221);
nor U9123 (N_9123,N_5516,N_6005);
nand U9124 (N_9124,N_6542,N_6629);
or U9125 (N_9125,N_6932,N_5251);
and U9126 (N_9126,N_5538,N_6733);
or U9127 (N_9127,N_5746,N_6317);
or U9128 (N_9128,N_6999,N_5873);
and U9129 (N_9129,N_5974,N_6635);
and U9130 (N_9130,N_6728,N_7277);
nand U9131 (N_9131,N_6773,N_7498);
nand U9132 (N_9132,N_5709,N_7117);
nand U9133 (N_9133,N_6488,N_5941);
nor U9134 (N_9134,N_5063,N_6492);
nand U9135 (N_9135,N_5157,N_6886);
nand U9136 (N_9136,N_5702,N_5626);
nor U9137 (N_9137,N_5023,N_7309);
nand U9138 (N_9138,N_6998,N_5161);
nand U9139 (N_9139,N_6084,N_6655);
or U9140 (N_9140,N_6045,N_5428);
or U9141 (N_9141,N_7061,N_5699);
nor U9142 (N_9142,N_6212,N_7227);
and U9143 (N_9143,N_6375,N_5807);
nor U9144 (N_9144,N_6136,N_6487);
or U9145 (N_9145,N_5515,N_5863);
nand U9146 (N_9146,N_6018,N_5899);
or U9147 (N_9147,N_6080,N_6596);
and U9148 (N_9148,N_6160,N_5411);
nor U9149 (N_9149,N_5752,N_6353);
and U9150 (N_9150,N_6793,N_7310);
and U9151 (N_9151,N_7311,N_5236);
nor U9152 (N_9152,N_5131,N_6406);
nor U9153 (N_9153,N_5421,N_6094);
and U9154 (N_9154,N_5462,N_5803);
or U9155 (N_9155,N_5661,N_5863);
and U9156 (N_9156,N_5991,N_5023);
and U9157 (N_9157,N_6738,N_6270);
and U9158 (N_9158,N_6400,N_6091);
nor U9159 (N_9159,N_6914,N_5879);
nand U9160 (N_9160,N_6923,N_6448);
nand U9161 (N_9161,N_6152,N_7252);
nor U9162 (N_9162,N_5846,N_6769);
nor U9163 (N_9163,N_6444,N_6476);
or U9164 (N_9164,N_6019,N_6989);
nor U9165 (N_9165,N_6288,N_5303);
nor U9166 (N_9166,N_6705,N_7215);
nand U9167 (N_9167,N_6083,N_6141);
nor U9168 (N_9168,N_7250,N_5172);
nand U9169 (N_9169,N_6916,N_7477);
nor U9170 (N_9170,N_6739,N_5968);
or U9171 (N_9171,N_6356,N_6346);
nor U9172 (N_9172,N_6715,N_7488);
nand U9173 (N_9173,N_5475,N_7379);
and U9174 (N_9174,N_6375,N_5722);
nor U9175 (N_9175,N_6682,N_6114);
nor U9176 (N_9176,N_7398,N_5147);
or U9177 (N_9177,N_6694,N_6827);
nand U9178 (N_9178,N_5039,N_6794);
nor U9179 (N_9179,N_6844,N_6896);
and U9180 (N_9180,N_6503,N_7153);
or U9181 (N_9181,N_5538,N_6866);
nand U9182 (N_9182,N_5985,N_5816);
or U9183 (N_9183,N_5205,N_5820);
and U9184 (N_9184,N_6908,N_5770);
xnor U9185 (N_9185,N_5864,N_6108);
nor U9186 (N_9186,N_5865,N_5261);
nor U9187 (N_9187,N_5760,N_6082);
or U9188 (N_9188,N_6700,N_6348);
and U9189 (N_9189,N_5106,N_5832);
nand U9190 (N_9190,N_6070,N_6393);
nand U9191 (N_9191,N_5461,N_5478);
nor U9192 (N_9192,N_6536,N_5891);
and U9193 (N_9193,N_5665,N_7092);
and U9194 (N_9194,N_5731,N_6035);
or U9195 (N_9195,N_7337,N_5532);
and U9196 (N_9196,N_7453,N_5306);
nor U9197 (N_9197,N_7279,N_6440);
or U9198 (N_9198,N_5362,N_6837);
or U9199 (N_9199,N_7401,N_5268);
nor U9200 (N_9200,N_6050,N_5524);
and U9201 (N_9201,N_5935,N_5203);
nand U9202 (N_9202,N_5867,N_6737);
nor U9203 (N_9203,N_5118,N_7259);
or U9204 (N_9204,N_6903,N_5460);
or U9205 (N_9205,N_6031,N_6194);
and U9206 (N_9206,N_5294,N_7018);
or U9207 (N_9207,N_5032,N_7367);
or U9208 (N_9208,N_6812,N_6781);
nor U9209 (N_9209,N_7257,N_6303);
nor U9210 (N_9210,N_5471,N_5492);
nand U9211 (N_9211,N_7445,N_6372);
or U9212 (N_9212,N_5746,N_6541);
and U9213 (N_9213,N_6931,N_5740);
nor U9214 (N_9214,N_6293,N_5993);
and U9215 (N_9215,N_7184,N_6303);
nand U9216 (N_9216,N_6695,N_7113);
and U9217 (N_9217,N_6514,N_5714);
nand U9218 (N_9218,N_6730,N_6449);
or U9219 (N_9219,N_6422,N_6768);
nor U9220 (N_9220,N_6038,N_6980);
nand U9221 (N_9221,N_5542,N_7117);
nand U9222 (N_9222,N_6711,N_7416);
or U9223 (N_9223,N_6061,N_6845);
or U9224 (N_9224,N_5269,N_7208);
nor U9225 (N_9225,N_5071,N_5583);
or U9226 (N_9226,N_6577,N_6163);
and U9227 (N_9227,N_5784,N_5455);
or U9228 (N_9228,N_7159,N_6907);
or U9229 (N_9229,N_6491,N_7029);
nand U9230 (N_9230,N_6531,N_5794);
nor U9231 (N_9231,N_6085,N_5145);
xnor U9232 (N_9232,N_7037,N_7171);
and U9233 (N_9233,N_7059,N_5076);
and U9234 (N_9234,N_6134,N_7484);
and U9235 (N_9235,N_5758,N_5015);
nor U9236 (N_9236,N_7263,N_7210);
nor U9237 (N_9237,N_5923,N_7242);
nand U9238 (N_9238,N_7428,N_6403);
nand U9239 (N_9239,N_5373,N_6399);
or U9240 (N_9240,N_5731,N_6263);
and U9241 (N_9241,N_6747,N_6844);
or U9242 (N_9242,N_5286,N_5657);
nor U9243 (N_9243,N_5102,N_6392);
nand U9244 (N_9244,N_7476,N_5154);
nand U9245 (N_9245,N_6530,N_5512);
or U9246 (N_9246,N_6471,N_6127);
and U9247 (N_9247,N_5134,N_7220);
nand U9248 (N_9248,N_6697,N_6609);
nand U9249 (N_9249,N_5791,N_6173);
or U9250 (N_9250,N_5604,N_5243);
and U9251 (N_9251,N_7143,N_6097);
or U9252 (N_9252,N_5799,N_6363);
nand U9253 (N_9253,N_5527,N_5591);
nand U9254 (N_9254,N_6865,N_7104);
nand U9255 (N_9255,N_6005,N_5240);
nand U9256 (N_9256,N_5673,N_7022);
nor U9257 (N_9257,N_5748,N_7131);
nor U9258 (N_9258,N_5791,N_7322);
nor U9259 (N_9259,N_5781,N_6994);
and U9260 (N_9260,N_6404,N_5570);
nand U9261 (N_9261,N_6536,N_5587);
and U9262 (N_9262,N_7234,N_5603);
and U9263 (N_9263,N_7214,N_7158);
or U9264 (N_9264,N_5076,N_5609);
nand U9265 (N_9265,N_5000,N_5871);
or U9266 (N_9266,N_6581,N_5762);
nor U9267 (N_9267,N_5698,N_6679);
nor U9268 (N_9268,N_6843,N_5698);
and U9269 (N_9269,N_5492,N_6856);
or U9270 (N_9270,N_6959,N_7031);
nand U9271 (N_9271,N_7257,N_7081);
nand U9272 (N_9272,N_5463,N_6340);
or U9273 (N_9273,N_6336,N_5268);
and U9274 (N_9274,N_5849,N_5121);
and U9275 (N_9275,N_6579,N_7463);
or U9276 (N_9276,N_5209,N_7113);
nor U9277 (N_9277,N_6460,N_5836);
nand U9278 (N_9278,N_6552,N_7114);
nor U9279 (N_9279,N_5270,N_7367);
nand U9280 (N_9280,N_5506,N_7258);
nor U9281 (N_9281,N_7254,N_6868);
or U9282 (N_9282,N_6030,N_5432);
and U9283 (N_9283,N_5554,N_6017);
or U9284 (N_9284,N_6023,N_7252);
or U9285 (N_9285,N_6965,N_7061);
nand U9286 (N_9286,N_6284,N_5011);
nand U9287 (N_9287,N_6790,N_7490);
nand U9288 (N_9288,N_5350,N_6038);
and U9289 (N_9289,N_6929,N_7269);
or U9290 (N_9290,N_5948,N_5413);
or U9291 (N_9291,N_6177,N_5544);
and U9292 (N_9292,N_7232,N_5000);
nand U9293 (N_9293,N_7359,N_5651);
and U9294 (N_9294,N_6574,N_6679);
nor U9295 (N_9295,N_5530,N_7280);
or U9296 (N_9296,N_6944,N_7441);
and U9297 (N_9297,N_5122,N_5021);
and U9298 (N_9298,N_5412,N_6056);
and U9299 (N_9299,N_6527,N_5227);
and U9300 (N_9300,N_7356,N_6027);
and U9301 (N_9301,N_7291,N_5262);
or U9302 (N_9302,N_5712,N_5327);
nand U9303 (N_9303,N_5197,N_5121);
or U9304 (N_9304,N_6372,N_6427);
and U9305 (N_9305,N_6724,N_5295);
or U9306 (N_9306,N_7446,N_5366);
nand U9307 (N_9307,N_6067,N_6002);
nand U9308 (N_9308,N_5210,N_5896);
nor U9309 (N_9309,N_6084,N_7467);
nor U9310 (N_9310,N_6512,N_7198);
or U9311 (N_9311,N_6588,N_6533);
nor U9312 (N_9312,N_5297,N_5045);
and U9313 (N_9313,N_7442,N_5776);
nor U9314 (N_9314,N_5670,N_5133);
and U9315 (N_9315,N_6068,N_6128);
nand U9316 (N_9316,N_6037,N_6374);
or U9317 (N_9317,N_6481,N_7438);
nor U9318 (N_9318,N_5470,N_5205);
or U9319 (N_9319,N_6048,N_6111);
nand U9320 (N_9320,N_5519,N_5780);
nand U9321 (N_9321,N_5596,N_6512);
nor U9322 (N_9322,N_5129,N_7089);
nand U9323 (N_9323,N_6680,N_5515);
nand U9324 (N_9324,N_5241,N_7387);
and U9325 (N_9325,N_5722,N_5056);
nor U9326 (N_9326,N_7491,N_6897);
nand U9327 (N_9327,N_5903,N_7001);
xor U9328 (N_9328,N_5256,N_6944);
or U9329 (N_9329,N_6769,N_6508);
nand U9330 (N_9330,N_5603,N_5956);
and U9331 (N_9331,N_6845,N_6518);
and U9332 (N_9332,N_6709,N_5765);
or U9333 (N_9333,N_7486,N_5483);
nor U9334 (N_9334,N_5326,N_7082);
nand U9335 (N_9335,N_5893,N_5235);
nor U9336 (N_9336,N_6998,N_5486);
nand U9337 (N_9337,N_5481,N_7312);
or U9338 (N_9338,N_5998,N_6787);
nor U9339 (N_9339,N_5934,N_5323);
nor U9340 (N_9340,N_6552,N_6588);
nor U9341 (N_9341,N_5204,N_7168);
nor U9342 (N_9342,N_6462,N_5066);
nor U9343 (N_9343,N_6416,N_7083);
nor U9344 (N_9344,N_5312,N_5644);
nor U9345 (N_9345,N_5943,N_6269);
nor U9346 (N_9346,N_7039,N_5350);
or U9347 (N_9347,N_5908,N_5208);
nor U9348 (N_9348,N_5388,N_5071);
nand U9349 (N_9349,N_6979,N_6736);
and U9350 (N_9350,N_5100,N_5149);
or U9351 (N_9351,N_6458,N_5526);
or U9352 (N_9352,N_5983,N_6006);
and U9353 (N_9353,N_5412,N_6519);
nor U9354 (N_9354,N_5964,N_6470);
and U9355 (N_9355,N_7050,N_5487);
or U9356 (N_9356,N_5563,N_5236);
nand U9357 (N_9357,N_5284,N_6655);
and U9358 (N_9358,N_5466,N_7239);
or U9359 (N_9359,N_7262,N_6228);
nor U9360 (N_9360,N_6748,N_6340);
xnor U9361 (N_9361,N_5660,N_6972);
or U9362 (N_9362,N_6462,N_6799);
and U9363 (N_9363,N_6436,N_6322);
and U9364 (N_9364,N_6725,N_5821);
nor U9365 (N_9365,N_6845,N_6129);
and U9366 (N_9366,N_5420,N_6933);
or U9367 (N_9367,N_5144,N_5299);
nand U9368 (N_9368,N_5745,N_6497);
nand U9369 (N_9369,N_6780,N_6336);
or U9370 (N_9370,N_5290,N_5956);
nor U9371 (N_9371,N_6481,N_5512);
nand U9372 (N_9372,N_6944,N_6826);
nand U9373 (N_9373,N_6737,N_6293);
and U9374 (N_9374,N_6125,N_5840);
or U9375 (N_9375,N_5731,N_7379);
nor U9376 (N_9376,N_6664,N_6984);
or U9377 (N_9377,N_5233,N_5123);
nand U9378 (N_9378,N_6928,N_6979);
or U9379 (N_9379,N_6268,N_6645);
nor U9380 (N_9380,N_6329,N_6832);
nor U9381 (N_9381,N_6207,N_5213);
and U9382 (N_9382,N_7437,N_5643);
nor U9383 (N_9383,N_5002,N_5609);
nand U9384 (N_9384,N_5720,N_5831);
or U9385 (N_9385,N_5862,N_5660);
nand U9386 (N_9386,N_6971,N_5650);
nand U9387 (N_9387,N_5474,N_7305);
nand U9388 (N_9388,N_6920,N_5761);
nor U9389 (N_9389,N_5956,N_5087);
nor U9390 (N_9390,N_6963,N_6632);
nor U9391 (N_9391,N_5800,N_7157);
nand U9392 (N_9392,N_6889,N_5062);
xor U9393 (N_9393,N_5172,N_5626);
or U9394 (N_9394,N_7121,N_5553);
and U9395 (N_9395,N_5459,N_5655);
or U9396 (N_9396,N_6856,N_5923);
nor U9397 (N_9397,N_6684,N_7443);
or U9398 (N_9398,N_7177,N_6140);
nor U9399 (N_9399,N_6574,N_5465);
nand U9400 (N_9400,N_6697,N_6909);
nor U9401 (N_9401,N_5260,N_6375);
nor U9402 (N_9402,N_7037,N_5154);
and U9403 (N_9403,N_5888,N_7107);
and U9404 (N_9404,N_6234,N_6831);
or U9405 (N_9405,N_7183,N_5244);
nand U9406 (N_9406,N_5552,N_5110);
and U9407 (N_9407,N_6001,N_6787);
and U9408 (N_9408,N_6467,N_7377);
nand U9409 (N_9409,N_6779,N_6819);
and U9410 (N_9410,N_7447,N_7245);
nand U9411 (N_9411,N_5066,N_7157);
nor U9412 (N_9412,N_5206,N_7275);
and U9413 (N_9413,N_5811,N_6975);
and U9414 (N_9414,N_6562,N_7225);
nand U9415 (N_9415,N_6756,N_6469);
and U9416 (N_9416,N_5277,N_6127);
or U9417 (N_9417,N_6511,N_5910);
and U9418 (N_9418,N_5717,N_6067);
nand U9419 (N_9419,N_7089,N_5780);
and U9420 (N_9420,N_5312,N_6902);
nand U9421 (N_9421,N_6015,N_6349);
or U9422 (N_9422,N_7229,N_5813);
nand U9423 (N_9423,N_5024,N_5705);
nand U9424 (N_9424,N_6830,N_5550);
nor U9425 (N_9425,N_5442,N_6117);
nor U9426 (N_9426,N_5370,N_6260);
and U9427 (N_9427,N_6845,N_5714);
nor U9428 (N_9428,N_5096,N_7212);
or U9429 (N_9429,N_5410,N_6677);
nand U9430 (N_9430,N_5273,N_5827);
nand U9431 (N_9431,N_5379,N_6385);
or U9432 (N_9432,N_6941,N_7299);
and U9433 (N_9433,N_5815,N_7232);
or U9434 (N_9434,N_6546,N_6631);
nand U9435 (N_9435,N_5238,N_5141);
xnor U9436 (N_9436,N_6589,N_6542);
nor U9437 (N_9437,N_6691,N_5488);
or U9438 (N_9438,N_6395,N_5302);
nand U9439 (N_9439,N_5021,N_6314);
nand U9440 (N_9440,N_5360,N_5732);
and U9441 (N_9441,N_5839,N_5082);
nand U9442 (N_9442,N_5883,N_6674);
and U9443 (N_9443,N_6781,N_5147);
xor U9444 (N_9444,N_7303,N_6832);
and U9445 (N_9445,N_5969,N_6059);
or U9446 (N_9446,N_6239,N_5040);
and U9447 (N_9447,N_6879,N_7133);
or U9448 (N_9448,N_6517,N_6939);
or U9449 (N_9449,N_5970,N_6750);
nand U9450 (N_9450,N_5935,N_6834);
or U9451 (N_9451,N_5086,N_5092);
nor U9452 (N_9452,N_6555,N_5340);
nand U9453 (N_9453,N_7026,N_7271);
nor U9454 (N_9454,N_7488,N_6740);
nand U9455 (N_9455,N_6515,N_5961);
nand U9456 (N_9456,N_6314,N_6763);
nor U9457 (N_9457,N_6333,N_6707);
or U9458 (N_9458,N_5477,N_7471);
nand U9459 (N_9459,N_5150,N_5348);
and U9460 (N_9460,N_6524,N_5471);
or U9461 (N_9461,N_6384,N_6191);
or U9462 (N_9462,N_7311,N_7284);
and U9463 (N_9463,N_7374,N_5615);
or U9464 (N_9464,N_6126,N_5885);
nor U9465 (N_9465,N_6673,N_6217);
or U9466 (N_9466,N_6581,N_7463);
nand U9467 (N_9467,N_6677,N_6508);
or U9468 (N_9468,N_5101,N_5809);
nor U9469 (N_9469,N_6050,N_6144);
nand U9470 (N_9470,N_6028,N_5754);
or U9471 (N_9471,N_5253,N_5965);
and U9472 (N_9472,N_5256,N_7137);
nand U9473 (N_9473,N_5403,N_7205);
nand U9474 (N_9474,N_5236,N_5312);
and U9475 (N_9475,N_7478,N_5417);
or U9476 (N_9476,N_6556,N_7120);
nand U9477 (N_9477,N_7244,N_5909);
nand U9478 (N_9478,N_5811,N_7383);
nand U9479 (N_9479,N_6650,N_5047);
xor U9480 (N_9480,N_7344,N_6074);
or U9481 (N_9481,N_6041,N_6937);
nand U9482 (N_9482,N_6873,N_5975);
and U9483 (N_9483,N_7291,N_5706);
or U9484 (N_9484,N_5576,N_5983);
or U9485 (N_9485,N_5458,N_7101);
nand U9486 (N_9486,N_6318,N_6106);
or U9487 (N_9487,N_5107,N_5598);
or U9488 (N_9488,N_5536,N_6268);
and U9489 (N_9489,N_5006,N_5202);
nor U9490 (N_9490,N_5265,N_7047);
or U9491 (N_9491,N_7049,N_5096);
nand U9492 (N_9492,N_5598,N_5405);
nor U9493 (N_9493,N_6058,N_5014);
nor U9494 (N_9494,N_7374,N_5727);
nand U9495 (N_9495,N_6227,N_7474);
nand U9496 (N_9496,N_5777,N_5588);
nand U9497 (N_9497,N_7222,N_5079);
and U9498 (N_9498,N_6249,N_6017);
and U9499 (N_9499,N_6468,N_6099);
nand U9500 (N_9500,N_6495,N_5873);
or U9501 (N_9501,N_6245,N_5501);
or U9502 (N_9502,N_5680,N_7381);
nor U9503 (N_9503,N_6175,N_6111);
or U9504 (N_9504,N_6792,N_7433);
nor U9505 (N_9505,N_6768,N_6083);
nand U9506 (N_9506,N_6673,N_6414);
and U9507 (N_9507,N_7210,N_7108);
nand U9508 (N_9508,N_5473,N_7060);
nor U9509 (N_9509,N_6204,N_5763);
or U9510 (N_9510,N_5763,N_5549);
nor U9511 (N_9511,N_5987,N_7023);
nor U9512 (N_9512,N_6832,N_6857);
nor U9513 (N_9513,N_6569,N_6050);
and U9514 (N_9514,N_7339,N_5430);
or U9515 (N_9515,N_6347,N_7469);
or U9516 (N_9516,N_5960,N_6343);
or U9517 (N_9517,N_7001,N_6045);
and U9518 (N_9518,N_6424,N_6655);
nor U9519 (N_9519,N_5564,N_6020);
nand U9520 (N_9520,N_5657,N_6248);
and U9521 (N_9521,N_6916,N_6529);
xor U9522 (N_9522,N_6894,N_7163);
nor U9523 (N_9523,N_6768,N_5636);
and U9524 (N_9524,N_6644,N_5742);
and U9525 (N_9525,N_5736,N_6646);
or U9526 (N_9526,N_5648,N_7332);
or U9527 (N_9527,N_6879,N_7249);
nand U9528 (N_9528,N_5269,N_6823);
nor U9529 (N_9529,N_5047,N_7410);
or U9530 (N_9530,N_5959,N_5901);
and U9531 (N_9531,N_5986,N_7263);
nand U9532 (N_9532,N_6903,N_6098);
nor U9533 (N_9533,N_6496,N_6289);
and U9534 (N_9534,N_6970,N_6428);
and U9535 (N_9535,N_6584,N_7221);
nor U9536 (N_9536,N_5425,N_5431);
and U9537 (N_9537,N_5519,N_6552);
or U9538 (N_9538,N_5361,N_7008);
nand U9539 (N_9539,N_5469,N_7494);
nand U9540 (N_9540,N_6815,N_6391);
nand U9541 (N_9541,N_7495,N_6019);
nor U9542 (N_9542,N_6218,N_6978);
nor U9543 (N_9543,N_5377,N_6484);
and U9544 (N_9544,N_5311,N_6726);
nor U9545 (N_9545,N_6606,N_5601);
nand U9546 (N_9546,N_6356,N_7182);
nand U9547 (N_9547,N_5258,N_6429);
and U9548 (N_9548,N_6451,N_5496);
nand U9549 (N_9549,N_7064,N_6765);
nand U9550 (N_9550,N_5442,N_5566);
nor U9551 (N_9551,N_6158,N_5623);
nand U9552 (N_9552,N_7492,N_5126);
nand U9553 (N_9553,N_5469,N_6445);
or U9554 (N_9554,N_5016,N_7475);
nand U9555 (N_9555,N_5322,N_5072);
nor U9556 (N_9556,N_7183,N_6900);
nor U9557 (N_9557,N_7082,N_5465);
nand U9558 (N_9558,N_7187,N_7499);
or U9559 (N_9559,N_5645,N_5122);
nor U9560 (N_9560,N_5910,N_5896);
nor U9561 (N_9561,N_6383,N_5482);
nor U9562 (N_9562,N_6376,N_6322);
nor U9563 (N_9563,N_5536,N_6946);
or U9564 (N_9564,N_6229,N_5929);
and U9565 (N_9565,N_6595,N_6707);
nand U9566 (N_9566,N_5307,N_6147);
nand U9567 (N_9567,N_5126,N_7018);
nand U9568 (N_9568,N_6533,N_6659);
and U9569 (N_9569,N_6858,N_5254);
and U9570 (N_9570,N_5863,N_5658);
nand U9571 (N_9571,N_6350,N_5884);
or U9572 (N_9572,N_6968,N_6885);
nand U9573 (N_9573,N_6452,N_6837);
and U9574 (N_9574,N_6610,N_6088);
nand U9575 (N_9575,N_5525,N_5068);
and U9576 (N_9576,N_6261,N_6982);
or U9577 (N_9577,N_6745,N_6871);
nand U9578 (N_9578,N_6615,N_6935);
and U9579 (N_9579,N_6182,N_6542);
and U9580 (N_9580,N_5672,N_6609);
nand U9581 (N_9581,N_5036,N_7350);
and U9582 (N_9582,N_5412,N_7337);
and U9583 (N_9583,N_6339,N_6983);
or U9584 (N_9584,N_6991,N_6476);
or U9585 (N_9585,N_7154,N_5993);
or U9586 (N_9586,N_6337,N_5734);
nand U9587 (N_9587,N_5715,N_6347);
or U9588 (N_9588,N_5920,N_7492);
nand U9589 (N_9589,N_7297,N_6089);
and U9590 (N_9590,N_5191,N_5846);
and U9591 (N_9591,N_7234,N_6848);
and U9592 (N_9592,N_6542,N_7469);
and U9593 (N_9593,N_6343,N_6240);
nand U9594 (N_9594,N_7350,N_6533);
nor U9595 (N_9595,N_6430,N_6758);
or U9596 (N_9596,N_5393,N_6746);
nor U9597 (N_9597,N_7180,N_7131);
nor U9598 (N_9598,N_5054,N_6387);
and U9599 (N_9599,N_6999,N_5404);
or U9600 (N_9600,N_6407,N_6487);
nand U9601 (N_9601,N_7158,N_5747);
and U9602 (N_9602,N_6910,N_5754);
and U9603 (N_9603,N_5477,N_6524);
nor U9604 (N_9604,N_5693,N_5107);
nor U9605 (N_9605,N_5771,N_5201);
nand U9606 (N_9606,N_5171,N_6573);
and U9607 (N_9607,N_6641,N_6113);
and U9608 (N_9608,N_6804,N_6772);
nand U9609 (N_9609,N_7465,N_7412);
or U9610 (N_9610,N_6795,N_6244);
and U9611 (N_9611,N_6329,N_7278);
nand U9612 (N_9612,N_5448,N_7051);
nor U9613 (N_9613,N_7017,N_7319);
and U9614 (N_9614,N_6662,N_6113);
and U9615 (N_9615,N_6777,N_6912);
or U9616 (N_9616,N_6796,N_5535);
nand U9617 (N_9617,N_6564,N_7389);
or U9618 (N_9618,N_5474,N_6088);
nand U9619 (N_9619,N_7239,N_5602);
nor U9620 (N_9620,N_7030,N_7043);
nor U9621 (N_9621,N_7228,N_6900);
or U9622 (N_9622,N_7386,N_7007);
nor U9623 (N_9623,N_5517,N_6775);
nor U9624 (N_9624,N_5583,N_5649);
and U9625 (N_9625,N_5971,N_6843);
and U9626 (N_9626,N_5024,N_6927);
or U9627 (N_9627,N_5693,N_7118);
or U9628 (N_9628,N_6500,N_5478);
nand U9629 (N_9629,N_6999,N_7478);
and U9630 (N_9630,N_6175,N_6470);
nand U9631 (N_9631,N_5792,N_5527);
nor U9632 (N_9632,N_5728,N_5311);
nand U9633 (N_9633,N_7352,N_6992);
nand U9634 (N_9634,N_5804,N_7156);
nand U9635 (N_9635,N_5841,N_7105);
nand U9636 (N_9636,N_7024,N_7398);
or U9637 (N_9637,N_6617,N_7421);
nor U9638 (N_9638,N_6372,N_5847);
and U9639 (N_9639,N_7299,N_5532);
or U9640 (N_9640,N_5706,N_5848);
or U9641 (N_9641,N_5577,N_6731);
or U9642 (N_9642,N_5908,N_6121);
nor U9643 (N_9643,N_5681,N_7328);
nor U9644 (N_9644,N_6286,N_7275);
nand U9645 (N_9645,N_5349,N_5005);
nor U9646 (N_9646,N_5300,N_6036);
or U9647 (N_9647,N_6663,N_5733);
nor U9648 (N_9648,N_5007,N_5935);
or U9649 (N_9649,N_7012,N_7139);
or U9650 (N_9650,N_5837,N_7266);
or U9651 (N_9651,N_6736,N_5164);
or U9652 (N_9652,N_6973,N_7085);
and U9653 (N_9653,N_5430,N_6328);
nand U9654 (N_9654,N_6119,N_7362);
nor U9655 (N_9655,N_5703,N_5619);
nand U9656 (N_9656,N_6799,N_7213);
nor U9657 (N_9657,N_7128,N_6473);
nor U9658 (N_9658,N_5001,N_5622);
or U9659 (N_9659,N_7241,N_6129);
or U9660 (N_9660,N_5556,N_6634);
or U9661 (N_9661,N_7223,N_7111);
or U9662 (N_9662,N_6943,N_5968);
or U9663 (N_9663,N_7392,N_5052);
or U9664 (N_9664,N_5836,N_6963);
nor U9665 (N_9665,N_6093,N_5804);
nor U9666 (N_9666,N_6757,N_6141);
and U9667 (N_9667,N_6829,N_6244);
nand U9668 (N_9668,N_7039,N_6142);
nand U9669 (N_9669,N_5654,N_5136);
nor U9670 (N_9670,N_5049,N_5681);
nor U9671 (N_9671,N_5122,N_6374);
nor U9672 (N_9672,N_5224,N_6078);
nand U9673 (N_9673,N_5091,N_5533);
or U9674 (N_9674,N_7315,N_6903);
xnor U9675 (N_9675,N_7188,N_6265);
nor U9676 (N_9676,N_5675,N_5026);
or U9677 (N_9677,N_6644,N_5633);
and U9678 (N_9678,N_6095,N_5022);
and U9679 (N_9679,N_5099,N_6144);
xor U9680 (N_9680,N_7136,N_5363);
nand U9681 (N_9681,N_7093,N_7381);
nor U9682 (N_9682,N_6124,N_7236);
nor U9683 (N_9683,N_5062,N_5610);
and U9684 (N_9684,N_7198,N_6950);
nand U9685 (N_9685,N_5458,N_5685);
nand U9686 (N_9686,N_7487,N_5305);
or U9687 (N_9687,N_5941,N_6347);
or U9688 (N_9688,N_6621,N_7496);
and U9689 (N_9689,N_6693,N_6398);
nand U9690 (N_9690,N_6417,N_6937);
and U9691 (N_9691,N_6243,N_6097);
and U9692 (N_9692,N_5879,N_5304);
and U9693 (N_9693,N_5690,N_7011);
or U9694 (N_9694,N_6932,N_7339);
and U9695 (N_9695,N_6586,N_5555);
or U9696 (N_9696,N_5346,N_6178);
nand U9697 (N_9697,N_5641,N_6760);
and U9698 (N_9698,N_5712,N_6097);
nor U9699 (N_9699,N_6250,N_7145);
nor U9700 (N_9700,N_5498,N_7335);
and U9701 (N_9701,N_5020,N_5717);
and U9702 (N_9702,N_5212,N_5681);
nor U9703 (N_9703,N_6602,N_6643);
and U9704 (N_9704,N_6117,N_5119);
or U9705 (N_9705,N_6696,N_5904);
and U9706 (N_9706,N_6063,N_7007);
nand U9707 (N_9707,N_5463,N_5492);
nor U9708 (N_9708,N_5659,N_5949);
nor U9709 (N_9709,N_7236,N_5238);
or U9710 (N_9710,N_6698,N_5595);
xnor U9711 (N_9711,N_7456,N_6999);
and U9712 (N_9712,N_5118,N_6900);
or U9713 (N_9713,N_6387,N_6080);
nand U9714 (N_9714,N_6479,N_5703);
nand U9715 (N_9715,N_6328,N_5733);
xor U9716 (N_9716,N_5155,N_7165);
nand U9717 (N_9717,N_6911,N_6682);
and U9718 (N_9718,N_7282,N_5048);
and U9719 (N_9719,N_5780,N_7261);
nor U9720 (N_9720,N_7360,N_7265);
nand U9721 (N_9721,N_5410,N_6169);
and U9722 (N_9722,N_5079,N_6953);
and U9723 (N_9723,N_5239,N_7443);
or U9724 (N_9724,N_7014,N_5953);
nor U9725 (N_9725,N_7272,N_5097);
and U9726 (N_9726,N_5818,N_5798);
nand U9727 (N_9727,N_6007,N_6459);
nand U9728 (N_9728,N_5905,N_6829);
nand U9729 (N_9729,N_6201,N_6910);
nand U9730 (N_9730,N_6257,N_6664);
nand U9731 (N_9731,N_7217,N_5996);
or U9732 (N_9732,N_5607,N_5700);
or U9733 (N_9733,N_5075,N_6932);
nand U9734 (N_9734,N_5654,N_5032);
or U9735 (N_9735,N_7177,N_6532);
xnor U9736 (N_9736,N_7468,N_5884);
nor U9737 (N_9737,N_7378,N_5692);
nand U9738 (N_9738,N_7420,N_7165);
and U9739 (N_9739,N_5120,N_5867);
nor U9740 (N_9740,N_6873,N_7416);
or U9741 (N_9741,N_7372,N_6793);
nand U9742 (N_9742,N_5014,N_5718);
and U9743 (N_9743,N_5580,N_5251);
or U9744 (N_9744,N_5276,N_6544);
and U9745 (N_9745,N_6459,N_5467);
nand U9746 (N_9746,N_5444,N_5973);
nor U9747 (N_9747,N_5777,N_6295);
or U9748 (N_9748,N_6063,N_5928);
or U9749 (N_9749,N_5122,N_5395);
or U9750 (N_9750,N_5360,N_5436);
nor U9751 (N_9751,N_5301,N_5383);
xor U9752 (N_9752,N_6147,N_7253);
and U9753 (N_9753,N_7343,N_6604);
nor U9754 (N_9754,N_5306,N_7194);
or U9755 (N_9755,N_7394,N_7197);
nand U9756 (N_9756,N_5288,N_5281);
or U9757 (N_9757,N_6719,N_5739);
and U9758 (N_9758,N_6695,N_5010);
nor U9759 (N_9759,N_6864,N_6159);
or U9760 (N_9760,N_7235,N_5284);
xor U9761 (N_9761,N_6011,N_6091);
or U9762 (N_9762,N_5340,N_5314);
nor U9763 (N_9763,N_6382,N_7455);
or U9764 (N_9764,N_6275,N_5749);
nand U9765 (N_9765,N_6319,N_5974);
and U9766 (N_9766,N_7348,N_7019);
nand U9767 (N_9767,N_6579,N_5442);
xnor U9768 (N_9768,N_5937,N_6334);
or U9769 (N_9769,N_6180,N_6654);
nor U9770 (N_9770,N_6638,N_7040);
xnor U9771 (N_9771,N_5100,N_5554);
and U9772 (N_9772,N_5318,N_5835);
or U9773 (N_9773,N_6202,N_6093);
nand U9774 (N_9774,N_6545,N_5680);
or U9775 (N_9775,N_6211,N_5795);
nand U9776 (N_9776,N_5991,N_6945);
and U9777 (N_9777,N_5945,N_5298);
and U9778 (N_9778,N_7332,N_6505);
nor U9779 (N_9779,N_6118,N_5582);
nor U9780 (N_9780,N_5989,N_6905);
nor U9781 (N_9781,N_5488,N_6122);
and U9782 (N_9782,N_6784,N_6146);
or U9783 (N_9783,N_6268,N_6034);
nor U9784 (N_9784,N_5396,N_5108);
or U9785 (N_9785,N_5819,N_5328);
and U9786 (N_9786,N_6541,N_5271);
nand U9787 (N_9787,N_7300,N_7030);
nor U9788 (N_9788,N_6984,N_6659);
or U9789 (N_9789,N_5021,N_7359);
or U9790 (N_9790,N_5467,N_6184);
or U9791 (N_9791,N_7251,N_6425);
or U9792 (N_9792,N_6906,N_6224);
nor U9793 (N_9793,N_6495,N_6134);
nand U9794 (N_9794,N_7236,N_6471);
or U9795 (N_9795,N_5780,N_6028);
nor U9796 (N_9796,N_7381,N_5996);
nor U9797 (N_9797,N_7075,N_6664);
nand U9798 (N_9798,N_6525,N_6986);
or U9799 (N_9799,N_6495,N_5564);
nand U9800 (N_9800,N_6283,N_5210);
nand U9801 (N_9801,N_5450,N_5972);
or U9802 (N_9802,N_5779,N_5715);
nand U9803 (N_9803,N_6443,N_6293);
and U9804 (N_9804,N_5986,N_6097);
nand U9805 (N_9805,N_6184,N_5766);
and U9806 (N_9806,N_5948,N_6019);
nand U9807 (N_9807,N_5961,N_5010);
and U9808 (N_9808,N_6250,N_7298);
nand U9809 (N_9809,N_7006,N_5034);
or U9810 (N_9810,N_5407,N_6565);
and U9811 (N_9811,N_5553,N_5752);
nand U9812 (N_9812,N_7197,N_5097);
or U9813 (N_9813,N_7073,N_5092);
nor U9814 (N_9814,N_7257,N_5934);
nor U9815 (N_9815,N_5212,N_6023);
or U9816 (N_9816,N_6990,N_6142);
and U9817 (N_9817,N_5264,N_6513);
nand U9818 (N_9818,N_6464,N_7444);
nor U9819 (N_9819,N_7337,N_5521);
or U9820 (N_9820,N_5887,N_6122);
and U9821 (N_9821,N_5073,N_7251);
or U9822 (N_9822,N_5524,N_6333);
or U9823 (N_9823,N_5507,N_6167);
or U9824 (N_9824,N_7141,N_5274);
or U9825 (N_9825,N_6693,N_5620);
nand U9826 (N_9826,N_6192,N_5297);
and U9827 (N_9827,N_5957,N_6529);
and U9828 (N_9828,N_7279,N_6152);
and U9829 (N_9829,N_6649,N_5799);
nor U9830 (N_9830,N_6542,N_6048);
nand U9831 (N_9831,N_6506,N_7038);
nor U9832 (N_9832,N_7347,N_6587);
nand U9833 (N_9833,N_6202,N_7126);
nand U9834 (N_9834,N_6849,N_6898);
and U9835 (N_9835,N_6064,N_6686);
nand U9836 (N_9836,N_7266,N_6463);
or U9837 (N_9837,N_6361,N_6438);
and U9838 (N_9838,N_6058,N_6164);
or U9839 (N_9839,N_5385,N_5839);
and U9840 (N_9840,N_6314,N_5755);
nand U9841 (N_9841,N_6707,N_5174);
and U9842 (N_9842,N_6547,N_6155);
nor U9843 (N_9843,N_7304,N_5349);
nand U9844 (N_9844,N_6117,N_5534);
or U9845 (N_9845,N_5484,N_5630);
nand U9846 (N_9846,N_7106,N_7497);
or U9847 (N_9847,N_5900,N_6731);
or U9848 (N_9848,N_5307,N_7370);
or U9849 (N_9849,N_5715,N_6804);
nor U9850 (N_9850,N_5214,N_6747);
nand U9851 (N_9851,N_7250,N_5076);
nor U9852 (N_9852,N_7221,N_5267);
nor U9853 (N_9853,N_6865,N_5297);
nand U9854 (N_9854,N_5923,N_5060);
nand U9855 (N_9855,N_6202,N_7128);
or U9856 (N_9856,N_6739,N_5840);
or U9857 (N_9857,N_7126,N_5154);
or U9858 (N_9858,N_5576,N_5750);
nand U9859 (N_9859,N_5685,N_6124);
nand U9860 (N_9860,N_5377,N_5292);
and U9861 (N_9861,N_6463,N_6991);
and U9862 (N_9862,N_5632,N_6038);
or U9863 (N_9863,N_6144,N_5280);
nor U9864 (N_9864,N_5895,N_5426);
xor U9865 (N_9865,N_5821,N_6326);
and U9866 (N_9866,N_6254,N_5983);
nor U9867 (N_9867,N_7018,N_5037);
nand U9868 (N_9868,N_6313,N_5882);
and U9869 (N_9869,N_7414,N_6078);
and U9870 (N_9870,N_6171,N_5815);
and U9871 (N_9871,N_7469,N_5549);
nand U9872 (N_9872,N_7155,N_5739);
nor U9873 (N_9873,N_5273,N_6463);
nor U9874 (N_9874,N_6229,N_7181);
nand U9875 (N_9875,N_5346,N_5567);
and U9876 (N_9876,N_5354,N_5912);
and U9877 (N_9877,N_7385,N_5818);
and U9878 (N_9878,N_5701,N_5498);
or U9879 (N_9879,N_7233,N_5527);
nand U9880 (N_9880,N_6825,N_7321);
nand U9881 (N_9881,N_5893,N_6626);
or U9882 (N_9882,N_5540,N_6742);
xor U9883 (N_9883,N_5182,N_7339);
nor U9884 (N_9884,N_5673,N_6928);
and U9885 (N_9885,N_7129,N_6448);
nor U9886 (N_9886,N_6894,N_6168);
or U9887 (N_9887,N_5610,N_6636);
nand U9888 (N_9888,N_5642,N_7192);
or U9889 (N_9889,N_6431,N_6238);
and U9890 (N_9890,N_6985,N_6982);
nor U9891 (N_9891,N_5347,N_5036);
nor U9892 (N_9892,N_7022,N_7096);
nor U9893 (N_9893,N_7469,N_5705);
and U9894 (N_9894,N_5913,N_7347);
or U9895 (N_9895,N_6712,N_7079);
and U9896 (N_9896,N_6116,N_6226);
nor U9897 (N_9897,N_5980,N_6436);
and U9898 (N_9898,N_7404,N_5161);
or U9899 (N_9899,N_7186,N_5269);
and U9900 (N_9900,N_6086,N_5292);
nand U9901 (N_9901,N_6044,N_6577);
or U9902 (N_9902,N_5761,N_5500);
nor U9903 (N_9903,N_6128,N_7368);
or U9904 (N_9904,N_6926,N_5655);
and U9905 (N_9905,N_6796,N_5172);
and U9906 (N_9906,N_6702,N_5241);
and U9907 (N_9907,N_5102,N_5483);
or U9908 (N_9908,N_5010,N_7457);
or U9909 (N_9909,N_5967,N_6654);
and U9910 (N_9910,N_5013,N_6074);
nor U9911 (N_9911,N_6977,N_7120);
nand U9912 (N_9912,N_5383,N_7373);
or U9913 (N_9913,N_5219,N_5261);
or U9914 (N_9914,N_6007,N_5954);
nor U9915 (N_9915,N_6716,N_6163);
or U9916 (N_9916,N_5423,N_6164);
and U9917 (N_9917,N_5717,N_5655);
and U9918 (N_9918,N_5276,N_5558);
and U9919 (N_9919,N_6799,N_5040);
nor U9920 (N_9920,N_6824,N_7264);
or U9921 (N_9921,N_6250,N_7278);
and U9922 (N_9922,N_5395,N_6935);
and U9923 (N_9923,N_5195,N_7202);
nor U9924 (N_9924,N_5256,N_5593);
nor U9925 (N_9925,N_6963,N_6544);
nand U9926 (N_9926,N_5974,N_6961);
nand U9927 (N_9927,N_5581,N_5984);
and U9928 (N_9928,N_5318,N_7108);
and U9929 (N_9929,N_5958,N_6384);
nand U9930 (N_9930,N_6580,N_6311);
and U9931 (N_9931,N_7346,N_6112);
or U9932 (N_9932,N_5992,N_5408);
or U9933 (N_9933,N_7034,N_5595);
or U9934 (N_9934,N_6667,N_6584);
nand U9935 (N_9935,N_6404,N_5329);
nor U9936 (N_9936,N_5594,N_5054);
and U9937 (N_9937,N_7257,N_6705);
or U9938 (N_9938,N_6344,N_5995);
nand U9939 (N_9939,N_7302,N_7038);
and U9940 (N_9940,N_5522,N_7054);
nand U9941 (N_9941,N_6792,N_6343);
nand U9942 (N_9942,N_6636,N_6293);
and U9943 (N_9943,N_5502,N_6078);
nor U9944 (N_9944,N_7222,N_6236);
and U9945 (N_9945,N_5317,N_5415);
or U9946 (N_9946,N_7357,N_7381);
nand U9947 (N_9947,N_6301,N_6913);
or U9948 (N_9948,N_7279,N_7278);
nand U9949 (N_9949,N_5239,N_7388);
nor U9950 (N_9950,N_7452,N_7394);
nor U9951 (N_9951,N_6376,N_5982);
nand U9952 (N_9952,N_6348,N_5359);
nand U9953 (N_9953,N_7253,N_5535);
nand U9954 (N_9954,N_6410,N_5131);
xnor U9955 (N_9955,N_7278,N_5417);
and U9956 (N_9956,N_6077,N_5733);
nor U9957 (N_9957,N_7146,N_7214);
nand U9958 (N_9958,N_5203,N_5350);
nor U9959 (N_9959,N_5582,N_6455);
and U9960 (N_9960,N_5992,N_6655);
nand U9961 (N_9961,N_5674,N_6230);
and U9962 (N_9962,N_5315,N_5299);
and U9963 (N_9963,N_7179,N_7020);
or U9964 (N_9964,N_5664,N_7487);
nand U9965 (N_9965,N_6330,N_7071);
nand U9966 (N_9966,N_5782,N_6769);
nand U9967 (N_9967,N_7042,N_6980);
and U9968 (N_9968,N_7427,N_5934);
nor U9969 (N_9969,N_5191,N_7168);
or U9970 (N_9970,N_6200,N_6202);
nand U9971 (N_9971,N_6995,N_6558);
nor U9972 (N_9972,N_6487,N_6262);
nor U9973 (N_9973,N_5274,N_6859);
nor U9974 (N_9974,N_7239,N_6298);
nor U9975 (N_9975,N_6403,N_6161);
nor U9976 (N_9976,N_6648,N_6287);
and U9977 (N_9977,N_5180,N_5466);
or U9978 (N_9978,N_5743,N_5305);
and U9979 (N_9979,N_5923,N_6343);
nor U9980 (N_9980,N_7161,N_6880);
nor U9981 (N_9981,N_7216,N_7296);
nand U9982 (N_9982,N_6399,N_5908);
nand U9983 (N_9983,N_6598,N_6082);
nand U9984 (N_9984,N_5718,N_5464);
nand U9985 (N_9985,N_6439,N_6224);
and U9986 (N_9986,N_6398,N_5998);
nand U9987 (N_9987,N_5502,N_5843);
or U9988 (N_9988,N_5761,N_7279);
or U9989 (N_9989,N_6235,N_5530);
nor U9990 (N_9990,N_5604,N_6903);
and U9991 (N_9991,N_7222,N_5625);
nand U9992 (N_9992,N_6664,N_6063);
nand U9993 (N_9993,N_6928,N_5237);
and U9994 (N_9994,N_7437,N_5740);
nand U9995 (N_9995,N_6500,N_7274);
nor U9996 (N_9996,N_5668,N_6899);
nor U9997 (N_9997,N_7026,N_5454);
nor U9998 (N_9998,N_6468,N_5288);
nor U9999 (N_9999,N_6675,N_6358);
and U10000 (N_10000,N_9479,N_9856);
and U10001 (N_10001,N_7997,N_8264);
nand U10002 (N_10002,N_8626,N_9114);
and U10003 (N_10003,N_8006,N_9616);
or U10004 (N_10004,N_9739,N_9065);
or U10005 (N_10005,N_8598,N_8368);
or U10006 (N_10006,N_9555,N_8194);
nor U10007 (N_10007,N_7936,N_8787);
or U10008 (N_10008,N_9144,N_8523);
nand U10009 (N_10009,N_8268,N_9539);
and U10010 (N_10010,N_8360,N_9228);
nor U10011 (N_10011,N_8242,N_9897);
and U10012 (N_10012,N_9116,N_7914);
and U10013 (N_10013,N_9466,N_7577);
and U10014 (N_10014,N_8563,N_9870);
or U10015 (N_10015,N_8485,N_8997);
nand U10016 (N_10016,N_7855,N_8344);
nor U10017 (N_10017,N_7580,N_9060);
or U10018 (N_10018,N_8929,N_9854);
nor U10019 (N_10019,N_7835,N_9209);
and U10020 (N_10020,N_9269,N_8202);
and U10021 (N_10021,N_7651,N_8298);
nor U10022 (N_10022,N_7711,N_9980);
nor U10023 (N_10023,N_9247,N_9160);
or U10024 (N_10024,N_9796,N_8966);
nand U10025 (N_10025,N_8948,N_9750);
nor U10026 (N_10026,N_8822,N_8043);
nor U10027 (N_10027,N_9632,N_8795);
nor U10028 (N_10028,N_9890,N_8687);
nand U10029 (N_10029,N_9028,N_8471);
nand U10030 (N_10030,N_8001,N_8486);
nor U10031 (N_10031,N_7660,N_9241);
nand U10032 (N_10032,N_8784,N_9418);
nand U10033 (N_10033,N_7766,N_8155);
nor U10034 (N_10034,N_8064,N_8529);
nor U10035 (N_10035,N_8976,N_9839);
nor U10036 (N_10036,N_8509,N_7776);
or U10037 (N_10037,N_7941,N_9438);
or U10038 (N_10038,N_7630,N_8540);
or U10039 (N_10039,N_7884,N_8084);
xor U10040 (N_10040,N_8203,N_8371);
or U10041 (N_10041,N_9793,N_9042);
nand U10042 (N_10042,N_9199,N_8534);
nand U10043 (N_10043,N_9688,N_7638);
and U10044 (N_10044,N_8317,N_7569);
xnor U10045 (N_10045,N_8081,N_9930);
and U10046 (N_10046,N_9267,N_9665);
nand U10047 (N_10047,N_9359,N_9195);
nor U10048 (N_10048,N_7597,N_9159);
and U10049 (N_10049,N_7998,N_9718);
and U10050 (N_10050,N_9562,N_8234);
nor U10051 (N_10051,N_7684,N_8335);
nor U10052 (N_10052,N_9553,N_8530);
and U10053 (N_10053,N_9902,N_9458);
or U10054 (N_10054,N_8710,N_9168);
nor U10055 (N_10055,N_7818,N_8852);
nor U10056 (N_10056,N_7792,N_9163);
or U10057 (N_10057,N_8220,N_8040);
nand U10058 (N_10058,N_7975,N_8481);
and U10059 (N_10059,N_8960,N_8536);
nor U10060 (N_10060,N_9222,N_8857);
nor U10061 (N_10061,N_8926,N_9573);
nor U10062 (N_10062,N_7947,N_7523);
nand U10063 (N_10063,N_7952,N_7524);
nor U10064 (N_10064,N_9327,N_8136);
and U10065 (N_10065,N_9243,N_9432);
nand U10066 (N_10066,N_8849,N_9231);
and U10067 (N_10067,N_7848,N_9900);
and U10068 (N_10068,N_8649,N_8621);
and U10069 (N_10069,N_9627,N_8083);
or U10070 (N_10070,N_7772,N_8694);
and U10071 (N_10071,N_8810,N_8443);
nor U10072 (N_10072,N_7655,N_7666);
nor U10073 (N_10073,N_9309,N_7511);
and U10074 (N_10074,N_8989,N_8178);
and U10075 (N_10075,N_9943,N_9957);
or U10076 (N_10076,N_9284,N_7981);
nor U10077 (N_10077,N_7592,N_8060);
nor U10078 (N_10078,N_8950,N_8867);
and U10079 (N_10079,N_7957,N_9026);
nand U10080 (N_10080,N_8856,N_9178);
nand U10081 (N_10081,N_9423,N_9310);
xnor U10082 (N_10082,N_9841,N_8881);
and U10083 (N_10083,N_7858,N_9487);
nor U10084 (N_10084,N_8351,N_9440);
nor U10085 (N_10085,N_9477,N_7650);
or U10086 (N_10086,N_9837,N_9869);
nand U10087 (N_10087,N_9765,N_7632);
or U10088 (N_10088,N_8745,N_8158);
nand U10089 (N_10089,N_9707,N_7877);
and U10090 (N_10090,N_9713,N_8514);
or U10091 (N_10091,N_9364,N_8827);
nor U10092 (N_10092,N_8601,N_9568);
and U10093 (N_10093,N_7538,N_7609);
nor U10094 (N_10094,N_8569,N_9365);
nand U10095 (N_10095,N_8454,N_9374);
and U10096 (N_10096,N_8915,N_9758);
nor U10097 (N_10097,N_7620,N_9536);
nand U10098 (N_10098,N_8968,N_7903);
nor U10099 (N_10099,N_8754,N_9133);
and U10100 (N_10100,N_9912,N_7752);
nor U10101 (N_10101,N_9524,N_9814);
and U10102 (N_10102,N_8640,N_7814);
and U10103 (N_10103,N_8975,N_7764);
nand U10104 (N_10104,N_8251,N_9817);
and U10105 (N_10105,N_7951,N_8904);
and U10106 (N_10106,N_8899,N_7929);
and U10107 (N_10107,N_9219,N_9139);
and U10108 (N_10108,N_9731,N_8100);
and U10109 (N_10109,N_8386,N_9409);
nor U10110 (N_10110,N_7992,N_8134);
and U10111 (N_10111,N_7823,N_9981);
and U10112 (N_10112,N_8165,N_8786);
nor U10113 (N_10113,N_9608,N_9610);
or U10114 (N_10114,N_9300,N_8357);
xnor U10115 (N_10115,N_9229,N_8492);
nand U10116 (N_10116,N_8753,N_9389);
nor U10117 (N_10117,N_7587,N_8637);
nand U10118 (N_10118,N_7810,N_9007);
or U10119 (N_10119,N_7667,N_8613);
and U10120 (N_10120,N_8225,N_7867);
and U10121 (N_10121,N_8107,N_8027);
nor U10122 (N_10122,N_8507,N_8126);
or U10123 (N_10123,N_8348,N_7549);
or U10124 (N_10124,N_9532,N_9911);
or U10125 (N_10125,N_9768,N_8253);
nand U10126 (N_10126,N_9344,N_9112);
or U10127 (N_10127,N_8572,N_7924);
or U10128 (N_10128,N_9755,N_9188);
or U10129 (N_10129,N_8157,N_9150);
nand U10130 (N_10130,N_8431,N_9887);
or U10131 (N_10131,N_8943,N_7505);
nor U10132 (N_10132,N_9262,N_7850);
and U10133 (N_10133,N_9771,N_9170);
nand U10134 (N_10134,N_8416,N_8110);
nor U10135 (N_10135,N_9121,N_8010);
nand U10136 (N_10136,N_9506,N_8893);
nor U10137 (N_10137,N_9543,N_8266);
and U10138 (N_10138,N_8248,N_9778);
or U10139 (N_10139,N_8362,N_8697);
and U10140 (N_10140,N_8952,N_9507);
or U10141 (N_10141,N_8617,N_8581);
and U10142 (N_10142,N_8538,N_9097);
nor U10143 (N_10143,N_9021,N_8630);
xnor U10144 (N_10144,N_9516,N_9772);
or U10145 (N_10145,N_9513,N_9586);
nand U10146 (N_10146,N_8680,N_9455);
and U10147 (N_10147,N_9431,N_7500);
nor U10148 (N_10148,N_7898,N_7748);
nor U10149 (N_10149,N_7842,N_9411);
or U10150 (N_10150,N_9034,N_7985);
or U10151 (N_10151,N_9719,N_9860);
or U10152 (N_10152,N_9711,N_8373);
nand U10153 (N_10153,N_7829,N_7782);
and U10154 (N_10154,N_8879,N_9214);
and U10155 (N_10155,N_9629,N_8295);
or U10156 (N_10156,N_9434,N_8669);
nand U10157 (N_10157,N_8823,N_9518);
nor U10158 (N_10158,N_9106,N_9978);
nand U10159 (N_10159,N_7537,N_8252);
and U10160 (N_10160,N_7532,N_9154);
or U10161 (N_10161,N_8546,N_9350);
xnor U10162 (N_10162,N_9538,N_8654);
and U10163 (N_10163,N_7624,N_9552);
nand U10164 (N_10164,N_8876,N_9279);
and U10165 (N_10165,N_8472,N_9955);
nand U10166 (N_10166,N_8781,N_9853);
or U10167 (N_10167,N_9250,N_8489);
and U10168 (N_10168,N_9172,N_7796);
and U10169 (N_10169,N_9657,N_8327);
and U10170 (N_10170,N_8661,N_8848);
and U10171 (N_10171,N_9313,N_8861);
nand U10172 (N_10172,N_9041,N_8378);
nor U10173 (N_10173,N_8618,N_9166);
nor U10174 (N_10174,N_7746,N_8686);
and U10175 (N_10175,N_9481,N_8185);
or U10176 (N_10176,N_8478,N_7674);
and U10177 (N_10177,N_9879,N_9500);
nor U10178 (N_10178,N_9966,N_8620);
and U10179 (N_10179,N_8183,N_7771);
nand U10180 (N_10180,N_8983,N_9009);
nor U10181 (N_10181,N_9642,N_9478);
nand U10182 (N_10182,N_8015,N_9035);
nor U10183 (N_10183,N_8095,N_8473);
nand U10184 (N_10184,N_8738,N_9910);
nor U10185 (N_10185,N_8636,N_8981);
nand U10186 (N_10186,N_8219,N_8945);
and U10187 (N_10187,N_9167,N_9877);
or U10188 (N_10188,N_9015,N_9847);
nor U10189 (N_10189,N_8312,N_7610);
and U10190 (N_10190,N_8839,N_9623);
nor U10191 (N_10191,N_8227,N_9463);
and U10192 (N_10192,N_8168,N_9985);
and U10193 (N_10193,N_8773,N_7988);
nand U10194 (N_10194,N_9488,N_9174);
nand U10195 (N_10195,N_7544,N_9357);
nand U10196 (N_10196,N_9164,N_9117);
or U10197 (N_10197,N_8097,N_9210);
or U10198 (N_10198,N_9726,N_9614);
nor U10199 (N_10199,N_7800,N_9000);
or U10200 (N_10200,N_7598,N_7557);
or U10201 (N_10201,N_7560,N_9609);
nor U10202 (N_10202,N_7989,N_9131);
nand U10203 (N_10203,N_8777,N_8265);
nor U10204 (N_10204,N_7959,N_8858);
or U10205 (N_10205,N_9446,N_7837);
nor U10206 (N_10206,N_9052,N_9384);
or U10207 (N_10207,N_8307,N_8476);
nand U10208 (N_10208,N_9027,N_8676);
nor U10209 (N_10209,N_8998,N_9343);
nor U10210 (N_10210,N_9550,N_7503);
nor U10211 (N_10211,N_8763,N_7590);
or U10212 (N_10212,N_9073,N_9227);
nand U10213 (N_10213,N_8591,N_8086);
and U10214 (N_10214,N_9119,N_8840);
nor U10215 (N_10215,N_9883,N_8955);
and U10216 (N_10216,N_8646,N_9085);
and U10217 (N_10217,N_8462,N_8016);
and U10218 (N_10218,N_8608,N_8908);
and U10219 (N_10219,N_9053,N_9485);
or U10220 (N_10220,N_8728,N_7912);
and U10221 (N_10221,N_9456,N_9744);
and U10222 (N_10222,N_7728,N_9014);
nor U10223 (N_10223,N_8761,N_8008);
nand U10224 (N_10224,N_8048,N_8042);
nor U10225 (N_10225,N_9889,N_8369);
nor U10226 (N_10226,N_8275,N_9412);
nor U10227 (N_10227,N_9512,N_8632);
nand U10228 (N_10228,N_7819,N_8731);
nor U10229 (N_10229,N_9931,N_9740);
nand U10230 (N_10230,N_7967,N_8394);
nand U10231 (N_10231,N_7956,N_9273);
or U10232 (N_10232,N_9305,N_8512);
nor U10233 (N_10233,N_9829,N_9450);
or U10234 (N_10234,N_9659,N_7716);
nor U10235 (N_10235,N_8841,N_7866);
or U10236 (N_10236,N_9563,N_8237);
and U10237 (N_10237,N_9406,N_8971);
or U10238 (N_10238,N_8885,N_8580);
nand U10239 (N_10239,N_9795,N_8583);
nor U10240 (N_10240,N_8869,N_8663);
nor U10241 (N_10241,N_7636,N_7955);
xnor U10242 (N_10242,N_8390,N_7890);
nor U10243 (N_10243,N_7901,N_8515);
or U10244 (N_10244,N_7953,N_9179);
or U10245 (N_10245,N_9748,N_8117);
nor U10246 (N_10246,N_9878,N_8482);
or U10247 (N_10247,N_8940,N_9358);
or U10248 (N_10248,N_8291,N_7554);
and U10249 (N_10249,N_7775,N_7783);
nand U10250 (N_10250,N_9193,N_8678);
nor U10251 (N_10251,N_8333,N_9521);
and U10252 (N_10252,N_7822,N_9819);
or U10253 (N_10253,N_9625,N_7589);
nand U10254 (N_10254,N_9903,N_8720);
or U10255 (N_10255,N_9048,N_7812);
nor U10256 (N_10256,N_8429,N_9529);
nor U10257 (N_10257,N_9451,N_7994);
nand U10258 (N_10258,N_8210,N_8779);
and U10259 (N_10259,N_8593,N_9782);
or U10260 (N_10260,N_9098,N_8576);
or U10261 (N_10261,N_9844,N_8764);
nand U10262 (N_10262,N_8077,N_9396);
and U10263 (N_10263,N_9898,N_9064);
or U10264 (N_10264,N_8316,N_8588);
or U10265 (N_10265,N_9324,N_7558);
nor U10266 (N_10266,N_8901,N_8545);
nand U10267 (N_10267,N_9548,N_9452);
nand U10268 (N_10268,N_9695,N_9323);
nor U10269 (N_10269,N_9025,N_8717);
and U10270 (N_10270,N_9245,N_9443);
nor U10271 (N_10271,N_8011,N_8766);
and U10272 (N_10272,N_9843,N_9528);
nand U10273 (N_10273,N_7767,N_9437);
and U10274 (N_10274,N_8294,N_8343);
or U10275 (N_10275,N_8657,N_8667);
or U10276 (N_10276,N_7540,N_9636);
nand U10277 (N_10277,N_8883,N_7599);
or U10278 (N_10278,N_7564,N_8332);
nor U10279 (N_10279,N_9630,N_9095);
and U10280 (N_10280,N_8181,N_7991);
xor U10281 (N_10281,N_9476,N_8286);
and U10282 (N_10282,N_9770,N_9546);
nand U10283 (N_10283,N_9801,N_8148);
nand U10284 (N_10284,N_9958,N_9331);
xnor U10285 (N_10285,N_8129,N_9611);
nor U10286 (N_10286,N_9705,N_8760);
and U10287 (N_10287,N_7679,N_9348);
or U10288 (N_10288,N_8282,N_7567);
or U10289 (N_10289,N_7622,N_9033);
xor U10290 (N_10290,N_8411,N_9111);
nand U10291 (N_10291,N_8555,N_8192);
nor U10292 (N_10292,N_8401,N_8897);
nor U10293 (N_10293,N_9427,N_9866);
or U10294 (N_10294,N_8740,N_9909);
and U10295 (N_10295,N_8956,N_7713);
nand U10296 (N_10296,N_8263,N_8603);
and U10297 (N_10297,N_9482,N_9729);
nand U10298 (N_10298,N_9896,N_8552);
and U10299 (N_10299,N_9678,N_9289);
and U10300 (N_10300,N_9387,N_8169);
and U10301 (N_10301,N_7826,N_7509);
nand U10302 (N_10302,N_9263,N_7768);
or U10303 (N_10303,N_8022,N_7677);
and U10304 (N_10304,N_9551,N_9276);
and U10305 (N_10305,N_8979,N_9804);
nand U10306 (N_10306,N_7779,N_9652);
or U10307 (N_10307,N_8375,N_9850);
and U10308 (N_10308,N_8393,N_7830);
nor U10309 (N_10309,N_7832,N_9992);
or U10310 (N_10310,N_8428,N_9975);
nand U10311 (N_10311,N_9846,N_8109);
and U10312 (N_10312,N_9401,N_8914);
and U10313 (N_10313,N_7714,N_8793);
nand U10314 (N_10314,N_9558,N_8715);
nand U10315 (N_10315,N_8870,N_9071);
nand U10316 (N_10316,N_9619,N_8522);
or U10317 (N_10317,N_9311,N_8108);
and U10318 (N_10318,N_9047,N_8074);
or U10319 (N_10319,N_9249,N_7659);
or U10320 (N_10320,N_8171,N_7904);
or U10321 (N_10321,N_8909,N_8681);
and U10322 (N_10322,N_9306,N_8487);
nor U10323 (N_10323,N_8382,N_7707);
nor U10324 (N_10324,N_9236,N_7581);
nand U10325 (N_10325,N_8341,N_9445);
nor U10326 (N_10326,N_9288,N_7512);
or U10327 (N_10327,N_8366,N_8293);
nor U10328 (N_10328,N_9338,N_9658);
nor U10329 (N_10329,N_7999,N_8161);
nor U10330 (N_10330,N_8318,N_9886);
or U10331 (N_10331,N_7908,N_8934);
nor U10332 (N_10332,N_8118,N_9928);
and U10333 (N_10333,N_8775,N_8067);
nand U10334 (N_10334,N_8888,N_9205);
or U10335 (N_10335,N_9607,N_8651);
or U10336 (N_10336,N_9907,N_9848);
nand U10337 (N_10337,N_8385,N_9371);
or U10338 (N_10338,N_9895,N_9134);
and U10339 (N_10339,N_7552,N_7520);
nor U10340 (N_10340,N_7911,N_8440);
or U10341 (N_10341,N_8695,N_7586);
nand U10342 (N_10342,N_7945,N_8093);
nand U10343 (N_10343,N_9746,N_8614);
and U10344 (N_10344,N_8223,N_8647);
nor U10345 (N_10345,N_8553,N_9029);
and U10346 (N_10346,N_9667,N_7611);
or U10347 (N_10347,N_8031,N_9986);
nand U10348 (N_10348,N_9380,N_9326);
nand U10349 (N_10349,N_9058,N_8882);
or U10350 (N_10350,N_8656,N_8211);
nor U10351 (N_10351,N_8400,N_7717);
and U10352 (N_10352,N_8682,N_8708);
or U10353 (N_10353,N_8337,N_8907);
nand U10354 (N_10354,N_9840,N_7652);
nor U10355 (N_10355,N_9915,N_8533);
and U10356 (N_10356,N_8670,N_9303);
nor U10357 (N_10357,N_7778,N_8246);
or U10358 (N_10358,N_9526,N_8550);
and U10359 (N_10359,N_9835,N_9424);
nor U10360 (N_10360,N_9838,N_9537);
nand U10361 (N_10361,N_8034,N_9504);
or U10362 (N_10362,N_9467,N_7614);
nand U10363 (N_10363,N_9135,N_7750);
and U10364 (N_10364,N_9290,N_9360);
nor U10365 (N_10365,N_9472,N_7799);
nand U10366 (N_10366,N_9349,N_8551);
xnor U10367 (N_10367,N_8494,N_9062);
nand U10368 (N_10368,N_8424,N_9011);
or U10369 (N_10369,N_8674,N_9091);
nand U10370 (N_10370,N_7661,N_8224);
and U10371 (N_10371,N_7977,N_7879);
nand U10372 (N_10372,N_7853,N_9519);
nand U10373 (N_10373,N_8056,N_9618);
nor U10374 (N_10374,N_8582,N_8499);
or U10375 (N_10375,N_8842,N_8936);
nor U10376 (N_10376,N_9641,N_9132);
or U10377 (N_10377,N_9691,N_9102);
nor U10378 (N_10378,N_7789,N_9833);
and U10379 (N_10379,N_8741,N_9407);
nand U10380 (N_10380,N_8430,N_8752);
nand U10381 (N_10381,N_9670,N_9716);
nand U10382 (N_10382,N_8402,N_9644);
or U10383 (N_10383,N_8387,N_8349);
and U10384 (N_10384,N_9924,N_9920);
and U10385 (N_10385,N_7543,N_9702);
nor U10386 (N_10386,N_7504,N_7887);
and U10387 (N_10387,N_9717,N_9834);
or U10388 (N_10388,N_8174,N_8313);
or U10389 (N_10389,N_9394,N_7920);
nand U10390 (N_10390,N_9312,N_9023);
xor U10391 (N_10391,N_7574,N_8491);
or U10392 (N_10392,N_8277,N_7980);
nand U10393 (N_10393,N_7939,N_7653);
nor U10394 (N_10394,N_9584,N_8379);
and U10395 (N_10395,N_7896,N_7600);
nor U10396 (N_10396,N_8041,N_9733);
nand U10397 (N_10397,N_9668,N_8150);
and U10398 (N_10398,N_9540,N_8190);
nor U10399 (N_10399,N_8450,N_9341);
and U10400 (N_10400,N_8999,N_9080);
nor U10401 (N_10401,N_9480,N_7712);
or U10402 (N_10402,N_7563,N_9317);
and U10403 (N_10403,N_8619,N_7935);
nor U10404 (N_10404,N_7798,N_9010);
or U10405 (N_10405,N_9974,N_8751);
or U10406 (N_10406,N_8123,N_7733);
nand U10407 (N_10407,N_8012,N_7897);
and U10408 (N_10408,N_9322,N_9325);
and U10409 (N_10409,N_8921,N_9603);
or U10410 (N_10410,N_9185,N_7629);
nand U10411 (N_10411,N_9191,N_8624);
nand U10412 (N_10412,N_8771,N_9926);
nor U10413 (N_10413,N_9809,N_9818);
nand U10414 (N_10414,N_9462,N_9950);
and U10415 (N_10415,N_8359,N_9218);
nor U10416 (N_10416,N_9684,N_9580);
nand U10417 (N_10417,N_9656,N_8575);
and U10418 (N_10418,N_9496,N_8742);
nand U10419 (N_10419,N_8249,N_7665);
or U10420 (N_10420,N_8834,N_8684);
nand U10421 (N_10421,N_9318,N_9781);
and U10422 (N_10422,N_8244,N_9275);
nor U10423 (N_10423,N_9587,N_8377);
nand U10424 (N_10424,N_7777,N_9631);
or U10425 (N_10425,N_9646,N_8791);
and U10426 (N_10426,N_9560,N_8496);
nand U10427 (N_10427,N_9031,N_9395);
or U10428 (N_10428,N_8510,N_9938);
nand U10429 (N_10429,N_7669,N_8007);
or U10430 (N_10430,N_8232,N_8207);
and U10431 (N_10431,N_9392,N_8917);
and U10432 (N_10432,N_9280,N_8954);
and U10433 (N_10433,N_8447,N_9808);
and U10434 (N_10434,N_8701,N_8325);
or U10435 (N_10435,N_9328,N_8420);
and U10436 (N_10436,N_8625,N_8096);
or U10437 (N_10437,N_8564,N_8306);
nand U10438 (N_10438,N_8898,N_9489);
nor U10439 (N_10439,N_7657,N_8951);
or U10440 (N_10440,N_8653,N_8596);
or U10441 (N_10441,N_9066,N_8149);
nor U10442 (N_10442,N_8860,N_9484);
nand U10443 (N_10443,N_9334,N_9595);
nand U10444 (N_10444,N_9505,N_7555);
or U10445 (N_10445,N_8816,N_9416);
and U10446 (N_10446,N_8895,N_8941);
and U10447 (N_10447,N_8991,N_8292);
nand U10448 (N_10448,N_9137,N_9292);
and U10449 (N_10449,N_8438,N_9791);
or U10450 (N_10450,N_8115,N_7693);
nor U10451 (N_10451,N_7513,N_8570);
and U10452 (N_10452,N_8836,N_9192);
nand U10453 (N_10453,N_9961,N_8389);
nor U10454 (N_10454,N_7781,N_8116);
nand U10455 (N_10455,N_7708,N_8970);
and U10456 (N_10456,N_7770,N_8597);
or U10457 (N_10457,N_7795,N_7742);
and U10458 (N_10458,N_7978,N_7900);
and U10459 (N_10459,N_9430,N_8837);
nand U10460 (N_10460,N_9346,N_9240);
and U10461 (N_10461,N_8578,N_8783);
and U10462 (N_10462,N_8047,N_8415);
and U10463 (N_10463,N_8833,N_9068);
and U10464 (N_10464,N_8103,N_8739);
nand U10465 (N_10465,N_9547,N_9723);
nand U10466 (N_10466,N_8498,N_8470);
and U10467 (N_10467,N_7642,N_7575);
nand U10468 (N_10468,N_9599,N_9594);
nand U10469 (N_10469,N_7883,N_9494);
or U10470 (N_10470,N_8247,N_8910);
and U10471 (N_10471,N_8151,N_9200);
or U10472 (N_10472,N_8974,N_8635);
nand U10473 (N_10473,N_7595,N_7919);
nand U10474 (N_10474,N_7612,N_9802);
nand U10475 (N_10475,N_9622,N_8121);
xnor U10476 (N_10476,N_8304,N_7545);
and U10477 (N_10477,N_9696,N_9320);
and U10478 (N_10478,N_9643,N_9579);
nor U10479 (N_10479,N_8437,N_8274);
or U10480 (N_10480,N_8830,N_9891);
nor U10481 (N_10481,N_9149,N_8843);
or U10482 (N_10482,N_8090,N_8612);
nor U10483 (N_10483,N_8537,N_7931);
and U10484 (N_10484,N_8054,N_8557);
and U10485 (N_10485,N_7553,N_7601);
and U10486 (N_10486,N_9790,N_9979);
nand U10487 (N_10487,N_9464,N_8631);
and U10488 (N_10488,N_9822,N_8407);
nand U10489 (N_10489,N_7976,N_9248);
or U10490 (N_10490,N_9677,N_9118);
or U10491 (N_10491,N_8864,N_8388);
nor U10492 (N_10492,N_9525,N_7573);
and U10493 (N_10493,N_9983,N_9984);
nor U10494 (N_10494,N_7670,N_9486);
or U10495 (N_10495,N_9465,N_9626);
or U10496 (N_10496,N_9302,N_8014);
or U10497 (N_10497,N_9020,N_7803);
nor U10498 (N_10498,N_9473,N_8502);
and U10499 (N_10499,N_8505,N_7582);
nor U10500 (N_10500,N_7649,N_8668);
and U10501 (N_10501,N_8147,N_9849);
or U10502 (N_10502,N_8949,N_7940);
or U10503 (N_10503,N_8854,N_8850);
or U10504 (N_10504,N_9260,N_9259);
and U10505 (N_10505,N_7725,N_8243);
or U10506 (N_10506,N_9354,N_8214);
or U10507 (N_10507,N_8285,N_8642);
nor U10508 (N_10508,N_9655,N_7643);
and U10509 (N_10509,N_9803,N_9405);
and U10510 (N_10510,N_7510,N_9422);
or U10511 (N_10511,N_9198,N_8182);
and U10512 (N_10512,N_9018,N_9736);
nand U10513 (N_10513,N_9105,N_8193);
or U10514 (N_10514,N_7730,N_9712);
nor U10515 (N_10515,N_9710,N_7790);
or U10516 (N_10516,N_9087,N_9760);
nand U10517 (N_10517,N_8794,N_9251);
or U10518 (N_10518,N_8871,N_9812);
nand U10519 (N_10519,N_8690,N_9184);
or U10520 (N_10520,N_8567,N_8946);
and U10521 (N_10521,N_7846,N_7747);
nor U10522 (N_10522,N_9730,N_9171);
nor U10523 (N_10523,N_8930,N_8939);
nor U10524 (N_10524,N_7514,N_9686);
nor U10525 (N_10525,N_8566,N_8330);
nand U10526 (N_10526,N_8127,N_8521);
and U10527 (N_10527,N_8868,N_9737);
nand U10528 (N_10528,N_9220,N_9460);
nor U10529 (N_10529,N_9202,N_8206);
nor U10530 (N_10530,N_8425,N_7983);
nor U10531 (N_10531,N_9542,N_7838);
and U10532 (N_10532,N_8130,N_9293);
nor U10533 (N_10533,N_9510,N_8577);
nor U10534 (N_10534,N_8920,N_7993);
or U10535 (N_10535,N_9330,N_7698);
nor U10536 (N_10536,N_7882,N_9086);
nand U10537 (N_10537,N_8495,N_8942);
or U10538 (N_10538,N_9238,N_8104);
or U10539 (N_10539,N_9763,N_9304);
or U10540 (N_10540,N_7880,N_8911);
and U10541 (N_10541,N_8352,N_8547);
nand U10542 (N_10542,N_8044,N_9811);
nand U10543 (N_10543,N_9008,N_7971);
and U10544 (N_10544,N_7815,N_8135);
nor U10545 (N_10545,N_9012,N_8560);
and U10546 (N_10546,N_7561,N_9875);
nand U10547 (N_10547,N_7909,N_9299);
nor U10548 (N_10548,N_8666,N_8452);
and U10549 (N_10549,N_7596,N_8785);
or U10550 (N_10550,N_8455,N_9232);
and U10551 (N_10551,N_8336,N_8200);
or U10552 (N_10552,N_9935,N_9013);
nand U10553 (N_10553,N_7943,N_9633);
nor U10554 (N_10554,N_8638,N_9217);
or U10555 (N_10555,N_8314,N_8627);
nor U10556 (N_10556,N_8988,N_9127);
nand U10557 (N_10557,N_8805,N_7949);
nand U10558 (N_10558,N_9993,N_9593);
or U10559 (N_10559,N_9408,N_9351);
and U10560 (N_10560,N_8984,N_8436);
nand U10561 (N_10561,N_8659,N_7892);
or U10562 (N_10562,N_9270,N_7825);
nor U10563 (N_10563,N_9367,N_7547);
or U10564 (N_10564,N_7979,N_8391);
nand U10565 (N_10565,N_8338,N_9382);
and U10566 (N_10566,N_9805,N_8933);
and U10567 (N_10567,N_8800,N_7787);
nor U10568 (N_10568,N_8776,N_8925);
nand U10569 (N_10569,N_7518,N_7671);
and U10570 (N_10570,N_7902,N_9180);
nand U10571 (N_10571,N_8723,N_8209);
nor U10572 (N_10572,N_9828,N_8633);
nand U10573 (N_10573,N_9520,N_9206);
nor U10574 (N_10574,N_8213,N_9821);
nor U10575 (N_10575,N_7811,N_7735);
nand U10576 (N_10576,N_9597,N_9393);
nor U10577 (N_10577,N_7710,N_8713);
nor U10578 (N_10578,N_9258,N_8721);
or U10579 (N_10579,N_7806,N_9882);
and U10580 (N_10580,N_8906,N_8039);
nor U10581 (N_10581,N_8579,N_9997);
or U10582 (N_10582,N_7678,N_9088);
nor U10583 (N_10583,N_8735,N_8821);
nand U10584 (N_10584,N_8480,N_8606);
nand U10585 (N_10585,N_7996,N_9441);
and U10586 (N_10586,N_8924,N_9099);
and U10587 (N_10587,N_7604,N_9352);
nor U10588 (N_10588,N_9442,N_8217);
nor U10589 (N_10589,N_8257,N_7786);
nor U10590 (N_10590,N_9973,N_8091);
or U10591 (N_10591,N_9541,N_9651);
or U10592 (N_10592,N_9138,N_7753);
nand U10593 (N_10593,N_9868,N_7893);
nor U10594 (N_10594,N_9161,N_9428);
nand U10595 (N_10595,N_8900,N_8334);
nand U10596 (N_10596,N_8356,N_9307);
nand U10597 (N_10597,N_7761,N_7541);
or U10598 (N_10598,N_8140,N_7579);
or U10599 (N_10599,N_7916,N_8700);
and U10600 (N_10600,N_9932,N_9383);
or U10601 (N_10601,N_7905,N_7954);
nand U10602 (N_10602,N_9905,N_7757);
nand U10603 (N_10603,N_8819,N_9561);
nand U10604 (N_10604,N_8590,N_8395);
nor U10605 (N_10605,N_7588,N_8872);
or U10606 (N_10606,N_8665,N_8996);
nor U10607 (N_10607,N_9283,N_8434);
nor U10608 (N_10608,N_7841,N_9146);
nor U10609 (N_10609,N_9495,N_9815);
or U10610 (N_10610,N_9294,N_7950);
and U10611 (N_10611,N_7862,N_8392);
nand U10612 (N_10612,N_9436,N_7802);
or U10613 (N_10613,N_8702,N_9904);
nor U10614 (N_10614,N_9151,N_7527);
nor U10615 (N_10615,N_7501,N_7721);
or U10616 (N_10616,N_9533,N_9761);
or U10617 (N_10617,N_8978,N_9749);
nand U10618 (N_10618,N_9559,N_9453);
nor U10619 (N_10619,N_9234,N_9335);
or U10620 (N_10620,N_7700,N_9454);
or U10621 (N_10621,N_8520,N_8111);
nor U10622 (N_10622,N_8051,N_9084);
nor U10623 (N_10623,N_8221,N_8463);
or U10624 (N_10624,N_8170,N_7664);
or U10625 (N_10625,N_9939,N_7754);
or U10626 (N_10626,N_7616,N_9693);
or U10627 (N_10627,N_8071,N_7606);
or U10628 (N_10628,N_8287,N_8714);
and U10629 (N_10629,N_7565,N_7517);
or U10630 (N_10630,N_9582,N_9576);
nand U10631 (N_10631,N_8574,N_8229);
nand U10632 (N_10632,N_8049,N_9372);
nor U10633 (N_10633,N_9660,N_8238);
or U10634 (N_10634,N_8299,N_9089);
nand U10635 (N_10635,N_8704,N_8053);
and U10636 (N_10636,N_8500,N_8609);
nand U10637 (N_10637,N_9994,N_7921);
xnor U10638 (N_10638,N_8743,N_8166);
and U10639 (N_10639,N_9929,N_9954);
or U10640 (N_10640,N_9720,N_7548);
nor U10641 (N_10641,N_8281,N_8085);
nor U10642 (N_10642,N_8812,N_9650);
nor U10643 (N_10643,N_8446,N_8384);
or U10644 (N_10644,N_9531,N_8802);
xor U10645 (N_10645,N_8855,N_9375);
or U10646 (N_10646,N_8113,N_8033);
nand U10647 (N_10647,N_7656,N_8623);
nand U10648 (N_10648,N_8412,N_8535);
nor U10649 (N_10649,N_8995,N_8722);
or U10650 (N_10650,N_9753,N_7762);
nand U10651 (N_10651,N_8878,N_9577);
or U10652 (N_10652,N_9591,N_7515);
or U10653 (N_10653,N_8815,N_8350);
or U10654 (N_10654,N_9556,N_8009);
and U10655 (N_10655,N_8231,N_8549);
xor U10656 (N_10656,N_8101,N_7986);
or U10657 (N_10657,N_7704,N_8397);
nor U10658 (N_10658,N_8453,N_7645);
nor U10659 (N_10659,N_8605,N_8442);
nand U10660 (N_10660,N_8208,N_7968);
nand U10661 (N_10661,N_8464,N_8189);
or U10662 (N_10662,N_9715,N_8762);
and U10663 (N_10663,N_8340,N_7922);
nand U10664 (N_10664,N_9735,N_9301);
nand U10665 (N_10665,N_9413,N_8187);
nor U10666 (N_10666,N_7619,N_7727);
nand U10667 (N_10667,N_7736,N_7519);
and U10668 (N_10668,N_8270,N_7720);
and U10669 (N_10669,N_8972,N_9982);
nand U10670 (N_10670,N_9329,N_9005);
nor U10671 (N_10671,N_7965,N_9662);
or U10672 (N_10672,N_7637,N_8218);
nor U10673 (N_10673,N_7780,N_9789);
nor U10674 (N_10674,N_8279,N_9377);
nor U10675 (N_10675,N_7572,N_9820);
or U10676 (N_10676,N_9004,N_9754);
nor U10677 (N_10677,N_8548,N_8005);
or U10678 (N_10678,N_7613,N_9224);
nand U10679 (N_10679,N_9638,N_8832);
or U10680 (N_10680,N_9752,N_8982);
or U10681 (N_10681,N_8036,N_9321);
nand U10682 (N_10682,N_9128,N_7937);
or U10683 (N_10683,N_7691,N_9922);
or U10684 (N_10684,N_9140,N_8028);
and U10685 (N_10685,N_8772,N_8828);
nand U10686 (N_10686,N_9063,N_7530);
nand U10687 (N_10687,N_8021,N_9046);
nor U10688 (N_10688,N_8128,N_9862);
and U10689 (N_10689,N_9810,N_7763);
or U10690 (N_10690,N_8571,N_9743);
nand U10691 (N_10691,N_9333,N_8912);
or U10692 (N_10692,N_7640,N_8250);
and U10693 (N_10693,N_9421,N_7556);
nor U10694 (N_10694,N_7641,N_9873);
and U10695 (N_10695,N_8894,N_9037);
nor U10696 (N_10696,N_8331,N_9773);
or U10697 (N_10697,N_7627,N_8880);
or U10698 (N_10698,N_8156,N_9876);
or U10699 (N_10699,N_9203,N_9277);
nand U10700 (N_10700,N_8584,N_9523);
nor U10701 (N_10701,N_9634,N_8874);
or U10702 (N_10702,N_9419,N_8080);
nor U10703 (N_10703,N_7918,N_8068);
nor U10704 (N_10704,N_8354,N_9295);
and U10705 (N_10705,N_9530,N_9965);
nand U10706 (N_10706,N_7773,N_7857);
xnor U10707 (N_10707,N_8891,N_8561);
nand U10708 (N_10708,N_8018,N_9798);
nand U10709 (N_10709,N_9757,N_9498);
nor U10710 (N_10710,N_9470,N_7942);
and U10711 (N_10711,N_9162,N_8241);
nor U10712 (N_10712,N_8256,N_9399);
and U10713 (N_10713,N_9177,N_9970);
nand U10714 (N_10714,N_8376,N_7621);
nor U10715 (N_10715,N_9388,N_7570);
or U10716 (N_10716,N_8105,N_9575);
nor U10717 (N_10717,N_9687,N_9635);
or U10718 (N_10718,N_7774,N_9971);
nor U10719 (N_10719,N_8835,N_8922);
nor U10720 (N_10720,N_9110,N_8652);
nor U10721 (N_10721,N_7690,N_9700);
nor U10722 (N_10722,N_8846,N_7602);
or U10723 (N_10723,N_7689,N_9792);
xor U10724 (N_10724,N_8019,N_7594);
or U10725 (N_10725,N_8037,N_9617);
or U10726 (N_10726,N_7966,N_9892);
nand U10727 (N_10727,N_9942,N_9226);
and U10728 (N_10728,N_9213,N_8967);
nor U10729 (N_10729,N_9257,N_8516);
nand U10730 (N_10730,N_8228,N_9081);
or U10731 (N_10731,N_9692,N_9515);
and U10732 (N_10732,N_9823,N_7987);
or U10733 (N_10733,N_9271,N_7964);
nor U10734 (N_10734,N_7646,N_9884);
nor U10735 (N_10735,N_9457,N_9208);
nor U10736 (N_10736,N_8662,N_8877);
nor U10737 (N_10737,N_9654,N_7765);
nor U10738 (N_10738,N_8239,N_8346);
and U10739 (N_10739,N_9756,N_7508);
or U10740 (N_10740,N_9129,N_9917);
nand U10741 (N_10741,N_8973,N_7930);
nand U10742 (N_10742,N_7963,N_7584);
nor U10743 (N_10743,N_8319,N_8639);
nor U10744 (N_10744,N_8504,N_9867);
nand U10745 (N_10745,N_9925,N_9706);
or U10746 (N_10746,N_7734,N_8131);
or U10747 (N_10747,N_8094,N_8532);
nor U10748 (N_10748,N_9680,N_9787);
nor U10749 (N_10749,N_8903,N_8986);
or U10750 (N_10750,N_9369,N_9264);
and U10751 (N_10751,N_9433,N_8527);
nand U10752 (N_10752,N_9522,N_9079);
nor U10753 (N_10753,N_8847,N_9893);
and U10754 (N_10754,N_7658,N_9246);
nor U10755 (N_10755,N_7843,N_8322);
nor U10756 (N_10756,N_9858,N_8778);
nand U10757 (N_10757,N_8448,N_9449);
nor U10758 (N_10758,N_8947,N_8004);
or U10759 (N_10759,N_7681,N_8517);
or U10760 (N_10760,N_7705,N_9585);
nor U10761 (N_10761,N_7723,N_8916);
and U10762 (N_10762,N_9953,N_9602);
xnor U10763 (N_10763,N_7851,N_8918);
and U10764 (N_10764,N_9061,N_8075);
nor U10765 (N_10765,N_8458,N_8052);
xor U10766 (N_10766,N_9336,N_7926);
or U10767 (N_10767,N_8405,N_8280);
and U10768 (N_10768,N_8699,N_8353);
nor U10769 (N_10769,N_9885,N_8276);
and U10770 (N_10770,N_9824,N_9002);
and U10771 (N_10771,N_7961,N_7809);
nand U10772 (N_10772,N_7793,N_7578);
nand U10773 (N_10773,N_9674,N_9130);
and U10774 (N_10774,N_9666,N_8825);
or U10775 (N_10775,N_8730,N_7969);
nand U10776 (N_10776,N_9747,N_9492);
and U10777 (N_10777,N_9420,N_8089);
and U10778 (N_10778,N_9447,N_7635);
and U10779 (N_10779,N_9759,N_9738);
nand U10780 (N_10780,N_9148,N_9989);
and U10781 (N_10781,N_9709,N_9152);
and U10782 (N_10782,N_9339,N_8254);
or U10783 (N_10783,N_7917,N_9050);
nand U10784 (N_10784,N_7876,N_9016);
nor U10785 (N_10785,N_8935,N_8062);
or U10786 (N_10786,N_8114,N_8607);
or U10787 (N_10787,N_8477,N_9239);
nor U10788 (N_10788,N_9113,N_7888);
nor U10789 (N_10789,N_8380,N_8261);
or U10790 (N_10790,N_8641,N_7872);
or U10791 (N_10791,N_8406,N_7934);
or U10792 (N_10792,N_8604,N_8413);
or U10793 (N_10793,N_9122,N_7889);
nor U10794 (N_10794,N_8092,N_7932);
or U10795 (N_10795,N_8796,N_9055);
nand U10796 (N_10796,N_9583,N_9775);
nand U10797 (N_10797,N_8398,N_8600);
or U10798 (N_10798,N_8746,N_7840);
nand U10799 (N_10799,N_9197,N_8602);
nand U10800 (N_10800,N_7706,N_8159);
or U10801 (N_10801,N_8737,N_8175);
and U10802 (N_10802,N_9386,N_8418);
or U10803 (N_10803,N_8539,N_7683);
nor U10804 (N_10804,N_9751,N_8383);
and U10805 (N_10805,N_8501,N_9664);
nand U10806 (N_10806,N_7794,N_9265);
nand U10807 (N_10807,N_7662,N_7854);
and U10808 (N_10808,N_9836,N_7536);
nand U10809 (N_10809,N_9813,N_9673);
or U10810 (N_10810,N_8315,N_9851);
or U10811 (N_10811,N_7928,N_9800);
and U10812 (N_10812,N_8152,N_7970);
or U10813 (N_10813,N_9285,N_8483);
or U10814 (N_10814,N_9908,N_9036);
or U10815 (N_10815,N_9483,N_9698);
nand U10816 (N_10816,N_9059,N_9572);
and U10817 (N_10817,N_8829,N_9825);
nor U10818 (N_10818,N_8003,N_8993);
nor U10819 (N_10819,N_8050,N_8977);
nor U10820 (N_10820,N_8519,N_9070);
or U10821 (N_10821,N_7871,N_7828);
nand U10822 (N_10822,N_9379,N_9832);
nor U10823 (N_10823,N_9972,N_9956);
nand U10824 (N_10824,N_7885,N_9566);
or U10825 (N_10825,N_8798,N_9780);
and U10826 (N_10826,N_8233,N_9762);
and U10827 (N_10827,N_8414,N_8139);
and U10828 (N_10828,N_9233,N_8141);
and U10829 (N_10829,N_9355,N_9962);
or U10830 (N_10830,N_9187,N_7938);
and U10831 (N_10831,N_8475,N_8544);
or U10832 (N_10832,N_8423,N_8137);
or U10833 (N_10833,N_7695,N_8179);
or U10834 (N_10834,N_8059,N_7680);
nand U10835 (N_10835,N_9968,N_8363);
or U10836 (N_10836,N_8289,N_9923);
and U10837 (N_10837,N_8045,N_9370);
nand U10838 (N_10838,N_8484,N_8057);
and U10839 (N_10839,N_9806,N_9914);
and U10840 (N_10840,N_9211,N_9067);
or U10841 (N_10841,N_8184,N_9946);
xor U10842 (N_10842,N_9779,N_7566);
or U10843 (N_10843,N_9176,N_7583);
and U10844 (N_10844,N_9244,N_7863);
nor U10845 (N_10845,N_7626,N_9298);
nand U10846 (N_10846,N_9143,N_7944);
and U10847 (N_10847,N_8066,N_8026);
and U10848 (N_10848,N_9136,N_8809);
nand U10849 (N_10849,N_9906,N_9256);
nor U10850 (N_10850,N_9921,N_9499);
nor U10851 (N_10851,N_8962,N_8622);
nor U10852 (N_10852,N_9769,N_8177);
and U10853 (N_10853,N_8524,N_8518);
or U10854 (N_10854,N_8980,N_7948);
nand U10855 (N_10855,N_8167,N_9024);
or U10856 (N_10856,N_8919,N_8706);
nand U10857 (N_10857,N_8245,N_8073);
or U10858 (N_10858,N_7542,N_8863);
nand U10859 (N_10859,N_9831,N_8873);
nand U10860 (N_10860,N_8734,N_8188);
nor U10861 (N_10861,N_9049,N_9278);
nand U10862 (N_10862,N_9827,N_7741);
nand U10863 (N_10863,N_8195,N_8079);
or U10864 (N_10864,N_8326,N_9308);
nand U10865 (N_10865,N_8303,N_7827);
nor U10866 (N_10866,N_9090,N_8427);
and U10867 (N_10867,N_8599,N_8799);
or U10868 (N_10868,N_9296,N_9030);
xnor U10869 (N_10869,N_9469,N_9268);
or U10870 (N_10870,N_8865,N_9281);
nor U10871 (N_10871,N_8000,N_8461);
or U10872 (N_10872,N_9254,N_9727);
nor U10873 (N_10873,N_9581,N_8323);
or U10874 (N_10874,N_8269,N_7817);
and U10875 (N_10875,N_8284,N_9991);
xor U10876 (N_10876,N_9045,N_9663);
and U10877 (N_10877,N_9072,N_9934);
nor U10878 (N_10878,N_8573,N_8660);
and U10879 (N_10879,N_8445,N_8162);
or U10880 (N_10880,N_8931,N_8204);
nand U10881 (N_10881,N_8409,N_7699);
and U10882 (N_10882,N_9342,N_9852);
nand U10883 (N_10883,N_7703,N_8419);
nand U10884 (N_10884,N_8272,N_8164);
and U10885 (N_10885,N_9040,N_8197);
nor U10886 (N_10886,N_8768,N_8435);
nor U10887 (N_10887,N_8146,N_9511);
nand U10888 (N_10888,N_9032,N_8927);
or U10889 (N_10889,N_7647,N_9728);
or U10890 (N_10890,N_8744,N_9165);
and U10891 (N_10891,N_9894,N_9977);
and U10892 (N_10892,N_9676,N_8689);
nor U10893 (N_10893,N_8508,N_8705);
nor U10894 (N_10894,N_9941,N_9842);
nand U10895 (N_10895,N_9816,N_8692);
xnor U10896 (N_10896,N_7894,N_8106);
or U10897 (N_10897,N_7927,N_9545);
xor U10898 (N_10898,N_8176,N_7839);
or U10899 (N_10899,N_9003,N_7933);
or U10900 (N_10900,N_9527,N_7718);
and U10901 (N_10901,N_9661,N_7831);
or U10902 (N_10902,N_8240,N_7833);
nor U10903 (N_10903,N_9940,N_8562);
nand U10904 (N_10904,N_9077,N_8506);
nand U10905 (N_10905,N_8311,N_8082);
and U10906 (N_10906,N_9429,N_9685);
or U10907 (N_10907,N_7824,N_9865);
or U10908 (N_10908,N_9742,N_9038);
nor U10909 (N_10909,N_8258,N_8339);
nand U10910 (N_10910,N_9252,N_9390);
and U10911 (N_10911,N_9807,N_9459);
nor U10912 (N_10912,N_7682,N_9286);
nand U10913 (N_10913,N_9044,N_8719);
nand U10914 (N_10914,N_8173,N_7522);
and U10915 (N_10915,N_9874,N_9400);
nor U10916 (N_10916,N_9175,N_9776);
nor U10917 (N_10917,N_7571,N_9291);
or U10918 (N_10918,N_8862,N_8216);
nand U10919 (N_10919,N_9589,N_8585);
nand U10920 (N_10920,N_7805,N_9094);
or U10921 (N_10921,N_8320,N_9588);
and U10922 (N_10922,N_8525,N_9403);
and U10923 (N_10923,N_8457,N_7516);
and U10924 (N_10924,N_7603,N_9682);
nand U10925 (N_10925,N_7808,N_8408);
nor U10926 (N_10926,N_7692,N_9212);
and U10927 (N_10927,N_9361,N_9398);
nor U10928 (N_10928,N_9444,N_9056);
nand U10929 (N_10929,N_7958,N_8154);
or U10930 (N_10930,N_7644,N_9919);
nor U10931 (N_10931,N_8801,N_9142);
nand U10932 (N_10932,N_8467,N_8098);
nand U10933 (N_10933,N_7697,N_9969);
nand U10934 (N_10934,N_9624,N_9987);
nor U10935 (N_10935,N_8142,N_8886);
or U10936 (N_10936,N_7535,N_9502);
and U10937 (N_10937,N_8138,N_7605);
nand U10938 (N_10938,N_9948,N_8814);
and U10939 (N_10939,N_8361,N_7673);
nand U10940 (N_10940,N_7531,N_8163);
nor U10941 (N_10941,N_7550,N_7506);
nor U10942 (N_10942,N_9314,N_9859);
and U10943 (N_10943,N_9414,N_9201);
nor U10944 (N_10944,N_8466,N_9671);
nor U10945 (N_10945,N_7849,N_9613);
xor U10946 (N_10946,N_8212,N_8818);
and U10947 (N_10947,N_7559,N_9057);
nor U10948 (N_10948,N_9082,N_9888);
nand U10949 (N_10949,N_7861,N_8513);
or U10950 (N_10950,N_9741,N_9937);
nand U10951 (N_10951,N_7801,N_8449);
or U10952 (N_10952,N_8774,N_8770);
nand U10953 (N_10953,N_8594,N_8677);
nor U10954 (N_10954,N_8568,N_8887);
and U10955 (N_10955,N_9725,N_8889);
xor U10956 (N_10956,N_8310,N_8712);
or U10957 (N_10957,N_8643,N_9628);
or U10958 (N_10958,N_9951,N_8201);
or U10959 (N_10959,N_8087,N_9315);
and U10960 (N_10960,N_9612,N_9871);
and U10961 (N_10961,N_7820,N_8905);
or U10962 (N_10962,N_8020,N_7568);
nor U10963 (N_10963,N_7607,N_9783);
nor U10964 (N_10964,N_9356,N_9714);
and U10965 (N_10965,N_7756,N_8267);
nor U10966 (N_10966,N_8683,N_8693);
nand U10967 (N_10967,N_9169,N_8300);
and U10968 (N_10968,N_9799,N_8417);
and U10969 (N_10969,N_7740,N_9100);
nor U10970 (N_10970,N_9147,N_7676);
or U10971 (N_10971,N_8866,N_8076);
nand U10972 (N_10972,N_9215,N_9266);
nand U10973 (N_10973,N_8072,N_9125);
nor U10974 (N_10974,N_9120,N_9703);
nor U10975 (N_10975,N_9381,N_7751);
and U10976 (N_10976,N_8358,N_9508);
nor U10977 (N_10977,N_7608,N_8365);
nor U10978 (N_10978,N_8987,N_8938);
and U10979 (N_10979,N_9237,N_9123);
or U10980 (N_10980,N_9439,N_8990);
or U10981 (N_10981,N_8273,N_9565);
or U10982 (N_10982,N_9497,N_8884);
and U10983 (N_10983,N_8490,N_8372);
and U10984 (N_10984,N_9933,N_8965);
and U10985 (N_10985,N_8592,N_9415);
and U10986 (N_10986,N_8892,N_7533);
or U10987 (N_10987,N_7821,N_9857);
nand U10988 (N_10988,N_9669,N_7910);
nand U10989 (N_10989,N_8589,N_8817);
or U10990 (N_10990,N_8961,N_8707);
nand U10991 (N_10991,N_9694,N_7685);
nand U10992 (N_10992,N_9093,N_9640);
nand U10993 (N_10993,N_7886,N_9108);
nor U10994 (N_10994,N_9391,N_7984);
nor U10995 (N_10995,N_8797,N_9944);
or U10996 (N_10996,N_8748,N_8444);
nor U10997 (N_10997,N_8556,N_8433);
nand U10998 (N_10998,N_8790,N_9207);
nor U10999 (N_10999,N_9282,N_9722);
and U11000 (N_11000,N_9101,N_9615);
nand U11001 (N_11001,N_7915,N_9990);
or U11002 (N_11002,N_9764,N_9039);
xnor U11003 (N_11003,N_7732,N_7648);
nand U11004 (N_11004,N_9272,N_8497);
or U11005 (N_11005,N_8679,N_9096);
or U11006 (N_11006,N_7816,N_9777);
nand U11007 (N_11007,N_8404,N_7576);
or U11008 (N_11008,N_7663,N_8629);
nand U11009 (N_11009,N_9845,N_8664);
nor U11010 (N_11010,N_8644,N_8994);
or U11011 (N_11011,N_8558,N_9104);
nand U11012 (N_11012,N_8469,N_8932);
and U11013 (N_11013,N_9503,N_7726);
and U11014 (N_11014,N_7585,N_7797);
nand U11015 (N_11015,N_7591,N_7722);
and U11016 (N_11016,N_8610,N_7834);
or U11017 (N_11017,N_7715,N_9242);
nand U11018 (N_11018,N_7634,N_9373);
nor U11019 (N_11019,N_7631,N_8441);
nand U11020 (N_11020,N_8696,N_9766);
nor U11021 (N_11021,N_8283,N_7895);
nand U11022 (N_11022,N_9679,N_8260);
or U11023 (N_11023,N_8859,N_8543);
and U11024 (N_11024,N_8724,N_9181);
nor U11025 (N_11025,N_9967,N_8046);
or U11026 (N_11026,N_8838,N_7878);
and U11027 (N_11027,N_8381,N_9794);
or U11028 (N_11028,N_7639,N_7759);
and U11029 (N_11029,N_7749,N_9362);
and U11030 (N_11030,N_8088,N_9952);
nand U11031 (N_11031,N_9590,N_9567);
nand U11032 (N_11032,N_8969,N_9999);
nor U11033 (N_11033,N_7675,N_8650);
and U11034 (N_11034,N_8186,N_8716);
nand U11035 (N_11035,N_8811,N_9216);
nor U11036 (N_11036,N_8456,N_7785);
nand U11037 (N_11037,N_9606,N_9156);
nand U11038 (N_11038,N_8985,N_9601);
nor U11039 (N_11039,N_9404,N_7760);
and U11040 (N_11040,N_8025,N_8459);
or U11041 (N_11041,N_8439,N_8732);
and U11042 (N_11042,N_7623,N_8586);
and U11043 (N_11043,N_9721,N_8308);
and U11044 (N_11044,N_8826,N_7528);
and U11045 (N_11045,N_8122,N_9683);
and U11046 (N_11046,N_8528,N_9689);
and U11047 (N_11047,N_9115,N_7847);
xnor U11048 (N_11048,N_8759,N_9767);
nand U11049 (N_11049,N_7534,N_8017);
nor U11050 (N_11050,N_8259,N_8645);
or U11051 (N_11051,N_9043,N_8554);
nor U11052 (N_11052,N_7521,N_9949);
nand U11053 (N_11053,N_7899,N_7856);
nor U11054 (N_11054,N_8964,N_9076);
nand U11055 (N_11055,N_7873,N_8526);
and U11056 (N_11056,N_8426,N_9785);
and U11057 (N_11057,N_9493,N_8230);
nor U11058 (N_11058,N_9855,N_8711);
nor U11059 (N_11059,N_8937,N_9899);
and U11060 (N_11060,N_9544,N_7864);
and U11061 (N_11061,N_7870,N_9880);
or U11062 (N_11062,N_9319,N_7907);
nor U11063 (N_11063,N_8875,N_9425);
and U11064 (N_11064,N_8465,N_9960);
and U11065 (N_11065,N_7551,N_8718);
or U11066 (N_11066,N_8070,N_8963);
nand U11067 (N_11067,N_7974,N_9620);
nor U11068 (N_11068,N_8112,N_7852);
nand U11069 (N_11069,N_9998,N_8672);
and U11070 (N_11070,N_7719,N_7724);
or U11071 (N_11071,N_9019,N_7807);
or U11072 (N_11072,N_9261,N_8288);
nor U11073 (N_11073,N_8703,N_7731);
and U11074 (N_11074,N_8769,N_9598);
or U11075 (N_11075,N_8957,N_8144);
and U11076 (N_11076,N_9491,N_8328);
and U11077 (N_11077,N_8460,N_7709);
and U11078 (N_11078,N_7923,N_9368);
and U11079 (N_11079,N_8671,N_7694);
nor U11080 (N_11080,N_9155,N_8749);
and U11081 (N_11081,N_8844,N_7784);
and U11082 (N_11082,N_7995,N_8180);
nor U11083 (N_11083,N_9690,N_7972);
nor U11084 (N_11084,N_9708,N_7529);
and U11085 (N_11085,N_9189,N_8944);
and U11086 (N_11086,N_9448,N_8831);
or U11087 (N_11087,N_9103,N_7769);
and U11088 (N_11088,N_9332,N_8758);
or U11089 (N_11089,N_8367,N_7744);
and U11090 (N_11090,N_8851,N_8078);
nor U11091 (N_11091,N_9704,N_9183);
nor U11092 (N_11092,N_8616,N_8410);
nor U11093 (N_11093,N_8262,N_8255);
or U11094 (N_11094,N_9517,N_8347);
nor U11095 (N_11095,N_8813,N_8132);
and U11096 (N_11096,N_7836,N_9645);
nand U11097 (N_11097,N_8145,N_8055);
or U11098 (N_11098,N_8587,N_9069);
and U11099 (N_11099,N_9426,N_9916);
and U11100 (N_11100,N_9230,N_8913);
or U11101 (N_11101,N_7960,N_9074);
and U11102 (N_11102,N_9959,N_9235);
nor U11103 (N_11103,N_8023,N_8757);
nand U11104 (N_11104,N_8172,N_9158);
nor U11105 (N_11105,N_9605,N_8205);
or U11106 (N_11106,N_9596,N_9927);
nand U11107 (N_11107,N_7617,N_8119);
nor U11108 (N_11108,N_8301,N_8493);
nor U11109 (N_11109,N_8729,N_7859);
nand U11110 (N_11110,N_8780,N_9054);
nand U11111 (N_11111,N_8782,N_8824);
and U11112 (N_11112,N_7788,N_9490);
and U11113 (N_11113,N_9774,N_8364);
and U11114 (N_11114,N_7739,N_9410);
and U11115 (N_11115,N_8198,N_8309);
nor U11116 (N_11116,N_8024,N_8923);
and U11117 (N_11117,N_7593,N_8160);
or U11118 (N_11118,N_8226,N_8675);
nand U11119 (N_11119,N_9006,N_8733);
and U11120 (N_11120,N_8215,N_9647);
or U11121 (N_11121,N_7874,N_8542);
nand U11122 (N_11122,N_9126,N_7844);
nand U11123 (N_11123,N_9826,N_9639);
nor U11124 (N_11124,N_9734,N_9083);
nand U11125 (N_11125,N_8658,N_9964);
nand U11126 (N_11126,N_7875,N_8342);
or U11127 (N_11127,N_7906,N_9675);
and U11128 (N_11128,N_8727,N_8673);
or U11129 (N_11129,N_8133,N_8890);
or U11130 (N_11130,N_9182,N_9988);
and U11131 (N_11131,N_9699,N_9863);
nor U11132 (N_11132,N_9397,N_7743);
nor U11133 (N_11133,N_7755,N_7804);
or U11134 (N_11134,N_9287,N_9881);
nand U11135 (N_11135,N_8736,N_9363);
nand U11136 (N_11136,N_9468,N_8709);
nor U11137 (N_11137,N_9534,N_7615);
and U11138 (N_11138,N_8222,N_7962);
or U11139 (N_11139,N_9996,N_8191);
nand U11140 (N_11140,N_8541,N_8958);
and U11141 (N_11141,N_8565,N_8806);
nand U11142 (N_11142,N_8820,N_8807);
or U11143 (N_11143,N_9022,N_7686);
nand U11144 (N_11144,N_8305,N_9402);
or U11145 (N_11145,N_8474,N_9637);
nor U11146 (N_11146,N_8655,N_8069);
nand U11147 (N_11147,N_9701,N_7973);
nand U11148 (N_11148,N_8726,N_8345);
nor U11149 (N_11149,N_9075,N_9578);
and U11150 (N_11150,N_7845,N_9366);
nor U11151 (N_11151,N_8302,N_9078);
nand U11152 (N_11152,N_8403,N_7654);
or U11153 (N_11153,N_8928,N_8953);
and U11154 (N_11154,N_9417,N_8767);
nand U11155 (N_11155,N_9435,N_8559);
or U11156 (N_11156,N_9223,N_7869);
or U11157 (N_11157,N_7737,N_9337);
nand U11158 (N_11158,N_9697,N_7502);
nand U11159 (N_11159,N_8611,N_8628);
or U11160 (N_11160,N_8065,N_9976);
nor U11161 (N_11161,N_9092,N_9509);
nand U11162 (N_11162,N_9501,N_8511);
nor U11163 (N_11163,N_8688,N_8685);
and U11164 (N_11164,N_9378,N_9124);
nand U11165 (N_11165,N_8747,N_7865);
and U11166 (N_11166,N_8278,N_9107);
nor U11167 (N_11167,N_8765,N_9901);
and U11168 (N_11168,N_8235,N_9514);
nor U11169 (N_11169,N_7925,N_9621);
nor U11170 (N_11170,N_8013,N_9173);
and U11171 (N_11171,N_9145,N_7625);
and U11172 (N_11172,N_9745,N_9274);
nand U11173 (N_11173,N_8099,N_9672);
and U11174 (N_11174,N_8329,N_7738);
or U11175 (N_11175,N_8648,N_8959);
nand U11176 (N_11176,N_8531,N_9297);
nand U11177 (N_11177,N_8789,N_8755);
or U11178 (N_11178,N_8853,N_8002);
and U11179 (N_11179,N_9221,N_8422);
or U11180 (N_11180,N_8061,N_9475);
or U11181 (N_11181,N_7758,N_7618);
nor U11182 (N_11182,N_7628,N_9569);
or U11183 (N_11183,N_8032,N_8451);
nor U11184 (N_11184,N_9648,N_9864);
or U11185 (N_11185,N_9347,N_9600);
nand U11186 (N_11186,N_9190,N_9017);
nor U11187 (N_11187,N_9253,N_8750);
nand U11188 (N_11188,N_9194,N_9786);
or U11189 (N_11189,N_9947,N_8396);
and U11190 (N_11190,N_7860,N_8029);
and U11191 (N_11191,N_8479,N_7688);
or U11192 (N_11192,N_8035,N_9157);
nor U11193 (N_11193,N_8421,N_7982);
or U11194 (N_11194,N_8845,N_8143);
nand U11195 (N_11195,N_8788,N_9861);
or U11196 (N_11196,N_7913,N_7701);
or U11197 (N_11197,N_9557,N_9345);
and U11198 (N_11198,N_7633,N_7729);
and U11199 (N_11199,N_8374,N_8803);
nor U11200 (N_11200,N_7745,N_9945);
nor U11201 (N_11201,N_9196,N_7546);
nand U11202 (N_11202,N_7791,N_9963);
and U11203 (N_11203,N_8153,N_9554);
or U11204 (N_11204,N_8804,N_8399);
xor U11205 (N_11205,N_9204,N_9549);
or U11206 (N_11206,N_9797,N_9141);
nor U11207 (N_11207,N_9724,N_8792);
nor U11208 (N_11208,N_8503,N_9995);
nor U11209 (N_11209,N_9830,N_8698);
and U11210 (N_11210,N_8355,N_8432);
nor U11211 (N_11211,N_7696,N_7525);
or U11212 (N_11212,N_8290,N_8992);
xor U11213 (N_11213,N_8595,N_7813);
nand U11214 (N_11214,N_9255,N_8199);
and U11215 (N_11215,N_7539,N_9653);
nand U11216 (N_11216,N_8808,N_9913);
and U11217 (N_11217,N_8321,N_9570);
nand U11218 (N_11218,N_9574,N_9376);
and U11219 (N_11219,N_8725,N_8324);
nor U11220 (N_11220,N_8124,N_9571);
nand U11221 (N_11221,N_8120,N_7526);
and U11222 (N_11222,N_9788,N_8756);
nor U11223 (N_11223,N_8468,N_8488);
nand U11224 (N_11224,N_7946,N_9604);
nor U11225 (N_11225,N_9649,N_9732);
nor U11226 (N_11226,N_7702,N_7990);
and U11227 (N_11227,N_8125,N_8297);
nor U11228 (N_11228,N_9474,N_9535);
nor U11229 (N_11229,N_7562,N_8896);
and U11230 (N_11230,N_9385,N_8063);
nor U11231 (N_11231,N_8902,N_9872);
nand U11232 (N_11232,N_7507,N_9186);
and U11233 (N_11233,N_8370,N_9316);
nand U11234 (N_11234,N_9936,N_9340);
or U11235 (N_11235,N_8296,N_9225);
nand U11236 (N_11236,N_8271,N_9109);
nor U11237 (N_11237,N_7868,N_7672);
and U11238 (N_11238,N_8236,N_8102);
nand U11239 (N_11239,N_9592,N_8615);
nor U11240 (N_11240,N_8038,N_8691);
nor U11241 (N_11241,N_9353,N_7687);
and U11242 (N_11242,N_9681,N_9784);
nand U11243 (N_11243,N_9471,N_8196);
nor U11244 (N_11244,N_9001,N_8058);
or U11245 (N_11245,N_9564,N_8030);
nor U11246 (N_11246,N_9051,N_7891);
or U11247 (N_11247,N_9153,N_8634);
or U11248 (N_11248,N_9918,N_7668);
nand U11249 (N_11249,N_7881,N_9461);
nand U11250 (N_11250,N_7779,N_9885);
xor U11251 (N_11251,N_8118,N_7786);
nor U11252 (N_11252,N_8742,N_9585);
nand U11253 (N_11253,N_8938,N_9352);
or U11254 (N_11254,N_9556,N_7885);
and U11255 (N_11255,N_9562,N_9270);
and U11256 (N_11256,N_9178,N_8478);
and U11257 (N_11257,N_9652,N_9517);
nor U11258 (N_11258,N_8869,N_9492);
nor U11259 (N_11259,N_9871,N_8052);
and U11260 (N_11260,N_8270,N_9943);
nand U11261 (N_11261,N_8132,N_8268);
or U11262 (N_11262,N_8166,N_8850);
nand U11263 (N_11263,N_9428,N_8493);
nor U11264 (N_11264,N_9838,N_7754);
or U11265 (N_11265,N_9326,N_8874);
nand U11266 (N_11266,N_8081,N_9206);
and U11267 (N_11267,N_9731,N_8872);
nand U11268 (N_11268,N_8250,N_9399);
and U11269 (N_11269,N_8528,N_9300);
nor U11270 (N_11270,N_8229,N_9189);
or U11271 (N_11271,N_7821,N_8503);
nor U11272 (N_11272,N_8369,N_8218);
and U11273 (N_11273,N_9454,N_8454);
nor U11274 (N_11274,N_8850,N_9635);
or U11275 (N_11275,N_8199,N_8242);
xnor U11276 (N_11276,N_8713,N_9590);
nand U11277 (N_11277,N_9460,N_8511);
nand U11278 (N_11278,N_8743,N_9122);
or U11279 (N_11279,N_9720,N_7927);
and U11280 (N_11280,N_8442,N_9641);
nor U11281 (N_11281,N_7599,N_7551);
and U11282 (N_11282,N_8802,N_8405);
and U11283 (N_11283,N_8023,N_8958);
nand U11284 (N_11284,N_8384,N_8940);
and U11285 (N_11285,N_9524,N_7561);
or U11286 (N_11286,N_9387,N_9986);
or U11287 (N_11287,N_7668,N_9709);
and U11288 (N_11288,N_9280,N_7507);
nor U11289 (N_11289,N_9833,N_8342);
nand U11290 (N_11290,N_8811,N_9492);
and U11291 (N_11291,N_8371,N_9479);
and U11292 (N_11292,N_8688,N_9531);
and U11293 (N_11293,N_7785,N_7983);
and U11294 (N_11294,N_8108,N_8444);
nor U11295 (N_11295,N_8149,N_9171);
nand U11296 (N_11296,N_8251,N_9636);
nor U11297 (N_11297,N_9797,N_9422);
and U11298 (N_11298,N_8973,N_8448);
and U11299 (N_11299,N_9580,N_8671);
and U11300 (N_11300,N_9891,N_8465);
nor U11301 (N_11301,N_9467,N_8713);
and U11302 (N_11302,N_8652,N_7620);
or U11303 (N_11303,N_7719,N_9682);
or U11304 (N_11304,N_7565,N_9936);
or U11305 (N_11305,N_7665,N_9554);
and U11306 (N_11306,N_9349,N_9674);
and U11307 (N_11307,N_9905,N_8198);
and U11308 (N_11308,N_8452,N_8936);
or U11309 (N_11309,N_9661,N_8040);
nor U11310 (N_11310,N_8811,N_9354);
and U11311 (N_11311,N_7840,N_9195);
nand U11312 (N_11312,N_9918,N_9506);
nand U11313 (N_11313,N_8215,N_8625);
and U11314 (N_11314,N_9721,N_7586);
or U11315 (N_11315,N_8358,N_7623);
nor U11316 (N_11316,N_9619,N_8480);
nor U11317 (N_11317,N_7688,N_8957);
nand U11318 (N_11318,N_8421,N_8034);
or U11319 (N_11319,N_8292,N_7904);
nand U11320 (N_11320,N_7528,N_9990);
and U11321 (N_11321,N_9255,N_9669);
nand U11322 (N_11322,N_9165,N_9017);
nand U11323 (N_11323,N_9206,N_8355);
xor U11324 (N_11324,N_7839,N_9731);
nor U11325 (N_11325,N_7811,N_9357);
or U11326 (N_11326,N_8317,N_9817);
and U11327 (N_11327,N_7800,N_8251);
nor U11328 (N_11328,N_7533,N_9077);
nand U11329 (N_11329,N_9678,N_9186);
and U11330 (N_11330,N_9689,N_8104);
nand U11331 (N_11331,N_8278,N_8589);
nor U11332 (N_11332,N_9218,N_8001);
nand U11333 (N_11333,N_8736,N_9978);
or U11334 (N_11334,N_8260,N_8900);
or U11335 (N_11335,N_8977,N_9412);
or U11336 (N_11336,N_8640,N_8652);
nand U11337 (N_11337,N_8890,N_8928);
and U11338 (N_11338,N_7671,N_8157);
nand U11339 (N_11339,N_8556,N_8352);
or U11340 (N_11340,N_8248,N_9596);
nor U11341 (N_11341,N_7979,N_9249);
nor U11342 (N_11342,N_9368,N_9246);
nand U11343 (N_11343,N_9748,N_9224);
and U11344 (N_11344,N_8749,N_8977);
or U11345 (N_11345,N_9847,N_8772);
nor U11346 (N_11346,N_8089,N_7852);
or U11347 (N_11347,N_9034,N_8047);
or U11348 (N_11348,N_9053,N_8808);
nand U11349 (N_11349,N_7501,N_9027);
or U11350 (N_11350,N_9570,N_9296);
nor U11351 (N_11351,N_8378,N_9052);
or U11352 (N_11352,N_7634,N_9854);
nand U11353 (N_11353,N_9183,N_7533);
nor U11354 (N_11354,N_7641,N_7538);
nand U11355 (N_11355,N_8749,N_7735);
nand U11356 (N_11356,N_8179,N_7676);
nand U11357 (N_11357,N_8504,N_7777);
nor U11358 (N_11358,N_9807,N_8720);
or U11359 (N_11359,N_9004,N_7903);
nor U11360 (N_11360,N_9746,N_8499);
or U11361 (N_11361,N_7676,N_9731);
or U11362 (N_11362,N_7848,N_8833);
or U11363 (N_11363,N_9075,N_8377);
and U11364 (N_11364,N_9134,N_8213);
nand U11365 (N_11365,N_9356,N_9681);
or U11366 (N_11366,N_9421,N_9357);
and U11367 (N_11367,N_8345,N_7536);
or U11368 (N_11368,N_9671,N_7829);
nor U11369 (N_11369,N_8545,N_8636);
nor U11370 (N_11370,N_9205,N_7630);
nand U11371 (N_11371,N_8597,N_7669);
or U11372 (N_11372,N_8131,N_9902);
and U11373 (N_11373,N_8704,N_9590);
xnor U11374 (N_11374,N_9676,N_8107);
nand U11375 (N_11375,N_8309,N_7537);
nor U11376 (N_11376,N_8401,N_7614);
nand U11377 (N_11377,N_7774,N_7970);
and U11378 (N_11378,N_7938,N_9851);
or U11379 (N_11379,N_8212,N_8705);
nand U11380 (N_11380,N_7919,N_8263);
and U11381 (N_11381,N_8503,N_7653);
nor U11382 (N_11382,N_9162,N_9114);
nand U11383 (N_11383,N_8513,N_7622);
or U11384 (N_11384,N_8253,N_7831);
nand U11385 (N_11385,N_8917,N_7864);
nor U11386 (N_11386,N_7525,N_9837);
and U11387 (N_11387,N_8480,N_8286);
and U11388 (N_11388,N_9695,N_9265);
nor U11389 (N_11389,N_7604,N_9262);
and U11390 (N_11390,N_8347,N_8652);
nand U11391 (N_11391,N_9878,N_9534);
nand U11392 (N_11392,N_8552,N_9233);
xor U11393 (N_11393,N_9704,N_7783);
and U11394 (N_11394,N_8457,N_8096);
and U11395 (N_11395,N_9081,N_9260);
nand U11396 (N_11396,N_9829,N_7757);
nand U11397 (N_11397,N_9566,N_9829);
or U11398 (N_11398,N_9266,N_9755);
nand U11399 (N_11399,N_8690,N_8049);
nand U11400 (N_11400,N_9262,N_8594);
nand U11401 (N_11401,N_9015,N_8492);
nor U11402 (N_11402,N_7688,N_7908);
or U11403 (N_11403,N_8911,N_8945);
nand U11404 (N_11404,N_8571,N_9258);
nand U11405 (N_11405,N_8341,N_8745);
and U11406 (N_11406,N_9825,N_9604);
nand U11407 (N_11407,N_9440,N_9320);
nor U11408 (N_11408,N_9636,N_9642);
nand U11409 (N_11409,N_9013,N_9059);
nor U11410 (N_11410,N_8793,N_9460);
and U11411 (N_11411,N_8144,N_8906);
or U11412 (N_11412,N_9895,N_7524);
nor U11413 (N_11413,N_8798,N_8458);
xnor U11414 (N_11414,N_9173,N_9908);
xor U11415 (N_11415,N_7546,N_7822);
nand U11416 (N_11416,N_7748,N_9266);
nor U11417 (N_11417,N_9960,N_8414);
and U11418 (N_11418,N_8678,N_8697);
nand U11419 (N_11419,N_8796,N_9517);
and U11420 (N_11420,N_8800,N_8604);
or U11421 (N_11421,N_9854,N_7992);
or U11422 (N_11422,N_7878,N_9753);
or U11423 (N_11423,N_9167,N_9299);
and U11424 (N_11424,N_8877,N_9020);
and U11425 (N_11425,N_7554,N_7867);
and U11426 (N_11426,N_7809,N_9204);
nor U11427 (N_11427,N_7803,N_9945);
or U11428 (N_11428,N_8077,N_8047);
nand U11429 (N_11429,N_8046,N_9746);
and U11430 (N_11430,N_9442,N_9140);
and U11431 (N_11431,N_8915,N_8860);
nor U11432 (N_11432,N_8572,N_8851);
nand U11433 (N_11433,N_8128,N_9532);
or U11434 (N_11434,N_8277,N_9394);
and U11435 (N_11435,N_9701,N_8037);
nand U11436 (N_11436,N_9661,N_9222);
and U11437 (N_11437,N_9463,N_8434);
and U11438 (N_11438,N_7756,N_8563);
or U11439 (N_11439,N_8365,N_8783);
nand U11440 (N_11440,N_8062,N_8709);
nand U11441 (N_11441,N_7947,N_8451);
nand U11442 (N_11442,N_8919,N_9594);
nand U11443 (N_11443,N_8871,N_9674);
or U11444 (N_11444,N_9641,N_9048);
nor U11445 (N_11445,N_9064,N_9312);
or U11446 (N_11446,N_8535,N_7992);
nand U11447 (N_11447,N_7516,N_9533);
or U11448 (N_11448,N_8812,N_8258);
nand U11449 (N_11449,N_7718,N_9948);
or U11450 (N_11450,N_8804,N_9316);
and U11451 (N_11451,N_9269,N_7881);
or U11452 (N_11452,N_8405,N_7775);
and U11453 (N_11453,N_7830,N_9593);
nor U11454 (N_11454,N_7907,N_9243);
nor U11455 (N_11455,N_7967,N_8187);
and U11456 (N_11456,N_7761,N_9254);
or U11457 (N_11457,N_8044,N_9377);
nand U11458 (N_11458,N_7582,N_7752);
and U11459 (N_11459,N_9660,N_9223);
or U11460 (N_11460,N_8544,N_9687);
nand U11461 (N_11461,N_8099,N_8172);
and U11462 (N_11462,N_8989,N_8008);
nand U11463 (N_11463,N_8595,N_8133);
nand U11464 (N_11464,N_9241,N_8014);
and U11465 (N_11465,N_9263,N_7648);
nor U11466 (N_11466,N_9728,N_8713);
and U11467 (N_11467,N_8539,N_8674);
nor U11468 (N_11468,N_8760,N_7716);
and U11469 (N_11469,N_8435,N_8118);
nor U11470 (N_11470,N_9081,N_9174);
and U11471 (N_11471,N_9416,N_9195);
or U11472 (N_11472,N_9869,N_9191);
nand U11473 (N_11473,N_8897,N_7704);
nand U11474 (N_11474,N_9970,N_9540);
or U11475 (N_11475,N_8216,N_7775);
nor U11476 (N_11476,N_8017,N_9154);
or U11477 (N_11477,N_9487,N_9276);
nand U11478 (N_11478,N_8071,N_9373);
or U11479 (N_11479,N_9518,N_8782);
or U11480 (N_11480,N_8385,N_8021);
nand U11481 (N_11481,N_9025,N_8359);
nand U11482 (N_11482,N_8605,N_9354);
nand U11483 (N_11483,N_7902,N_9848);
nor U11484 (N_11484,N_9827,N_9948);
and U11485 (N_11485,N_8050,N_7676);
or U11486 (N_11486,N_7793,N_7695);
nand U11487 (N_11487,N_7977,N_8560);
and U11488 (N_11488,N_8915,N_9888);
nor U11489 (N_11489,N_9558,N_8119);
nand U11490 (N_11490,N_9797,N_8630);
nor U11491 (N_11491,N_9115,N_8011);
nand U11492 (N_11492,N_9706,N_8647);
or U11493 (N_11493,N_7779,N_9903);
nand U11494 (N_11494,N_8468,N_7893);
or U11495 (N_11495,N_7534,N_8693);
nand U11496 (N_11496,N_8700,N_8997);
nand U11497 (N_11497,N_8310,N_8361);
nand U11498 (N_11498,N_8067,N_9065);
or U11499 (N_11499,N_7794,N_8267);
or U11500 (N_11500,N_9878,N_9069);
or U11501 (N_11501,N_8850,N_9004);
nand U11502 (N_11502,N_8729,N_8794);
nor U11503 (N_11503,N_7659,N_9425);
and U11504 (N_11504,N_8798,N_7575);
nand U11505 (N_11505,N_9317,N_7790);
nor U11506 (N_11506,N_9415,N_8119);
and U11507 (N_11507,N_9424,N_8776);
or U11508 (N_11508,N_8530,N_7589);
nand U11509 (N_11509,N_8200,N_9604);
or U11510 (N_11510,N_7932,N_7877);
and U11511 (N_11511,N_8954,N_9533);
and U11512 (N_11512,N_9145,N_8789);
xnor U11513 (N_11513,N_8710,N_9790);
or U11514 (N_11514,N_7543,N_9400);
nand U11515 (N_11515,N_8772,N_7647);
nand U11516 (N_11516,N_8194,N_9886);
nand U11517 (N_11517,N_9413,N_8619);
nor U11518 (N_11518,N_8622,N_8592);
nand U11519 (N_11519,N_7857,N_9137);
nand U11520 (N_11520,N_7773,N_9386);
or U11521 (N_11521,N_7759,N_9281);
or U11522 (N_11522,N_8232,N_8928);
nor U11523 (N_11523,N_8792,N_8755);
nor U11524 (N_11524,N_8532,N_9210);
nand U11525 (N_11525,N_9375,N_9953);
or U11526 (N_11526,N_9537,N_7654);
and U11527 (N_11527,N_9659,N_7770);
or U11528 (N_11528,N_8342,N_9605);
nand U11529 (N_11529,N_9627,N_9361);
nor U11530 (N_11530,N_8651,N_9415);
or U11531 (N_11531,N_9992,N_9917);
nand U11532 (N_11532,N_8811,N_9814);
nor U11533 (N_11533,N_8990,N_8852);
or U11534 (N_11534,N_7648,N_7576);
or U11535 (N_11535,N_8191,N_9229);
nand U11536 (N_11536,N_8488,N_8843);
nand U11537 (N_11537,N_7892,N_9031);
nand U11538 (N_11538,N_9643,N_9242);
and U11539 (N_11539,N_8745,N_9121);
nor U11540 (N_11540,N_7985,N_8515);
and U11541 (N_11541,N_9850,N_9888);
nor U11542 (N_11542,N_9630,N_9632);
or U11543 (N_11543,N_8644,N_7713);
nor U11544 (N_11544,N_8039,N_7714);
and U11545 (N_11545,N_7706,N_8196);
or U11546 (N_11546,N_9554,N_8225);
and U11547 (N_11547,N_8148,N_7974);
nor U11548 (N_11548,N_9355,N_7858);
or U11549 (N_11549,N_9966,N_9911);
and U11550 (N_11550,N_7944,N_8299);
nand U11551 (N_11551,N_8783,N_9986);
and U11552 (N_11552,N_7576,N_9369);
and U11553 (N_11553,N_9072,N_7541);
nor U11554 (N_11554,N_8254,N_8791);
and U11555 (N_11555,N_9692,N_9595);
nor U11556 (N_11556,N_9993,N_9682);
and U11557 (N_11557,N_8359,N_9958);
and U11558 (N_11558,N_8417,N_7622);
nand U11559 (N_11559,N_8938,N_9118);
nand U11560 (N_11560,N_7902,N_9114);
nor U11561 (N_11561,N_9618,N_9852);
or U11562 (N_11562,N_9280,N_7674);
or U11563 (N_11563,N_9031,N_7699);
nand U11564 (N_11564,N_9896,N_8576);
nor U11565 (N_11565,N_8827,N_8134);
nand U11566 (N_11566,N_9493,N_9247);
or U11567 (N_11567,N_8753,N_8215);
nor U11568 (N_11568,N_9396,N_9758);
nor U11569 (N_11569,N_8721,N_8184);
and U11570 (N_11570,N_9722,N_8854);
or U11571 (N_11571,N_7808,N_7986);
xnor U11572 (N_11572,N_8928,N_9788);
nor U11573 (N_11573,N_8518,N_9025);
nor U11574 (N_11574,N_9199,N_8236);
and U11575 (N_11575,N_8956,N_8988);
or U11576 (N_11576,N_9590,N_8659);
nand U11577 (N_11577,N_9592,N_9645);
or U11578 (N_11578,N_9239,N_8452);
nand U11579 (N_11579,N_9327,N_8114);
nor U11580 (N_11580,N_8007,N_8746);
nor U11581 (N_11581,N_8023,N_8557);
and U11582 (N_11582,N_9180,N_9714);
nor U11583 (N_11583,N_8089,N_9155);
nor U11584 (N_11584,N_9724,N_9069);
nand U11585 (N_11585,N_8303,N_8641);
and U11586 (N_11586,N_7801,N_8874);
and U11587 (N_11587,N_9818,N_8123);
and U11588 (N_11588,N_9192,N_7678);
nor U11589 (N_11589,N_9966,N_7573);
and U11590 (N_11590,N_8242,N_8077);
and U11591 (N_11591,N_9694,N_8331);
nor U11592 (N_11592,N_9012,N_7989);
or U11593 (N_11593,N_9600,N_9955);
nor U11594 (N_11594,N_8994,N_8959);
and U11595 (N_11595,N_7586,N_9551);
or U11596 (N_11596,N_8199,N_8682);
nor U11597 (N_11597,N_7569,N_9270);
nand U11598 (N_11598,N_7976,N_9746);
nand U11599 (N_11599,N_7607,N_9305);
or U11600 (N_11600,N_8066,N_8881);
nand U11601 (N_11601,N_8311,N_9522);
nand U11602 (N_11602,N_9845,N_8209);
nand U11603 (N_11603,N_8093,N_9547);
nor U11604 (N_11604,N_9798,N_8754);
and U11605 (N_11605,N_8090,N_8048);
nand U11606 (N_11606,N_7897,N_8244);
and U11607 (N_11607,N_8381,N_8092);
and U11608 (N_11608,N_7642,N_7930);
and U11609 (N_11609,N_9342,N_8705);
nand U11610 (N_11610,N_7881,N_9301);
nor U11611 (N_11611,N_8472,N_9833);
and U11612 (N_11612,N_9505,N_7777);
nand U11613 (N_11613,N_9504,N_8189);
and U11614 (N_11614,N_8989,N_8770);
and U11615 (N_11615,N_8666,N_8354);
and U11616 (N_11616,N_7615,N_7886);
nand U11617 (N_11617,N_8067,N_8520);
nand U11618 (N_11618,N_8813,N_8851);
nand U11619 (N_11619,N_9354,N_8769);
nor U11620 (N_11620,N_9759,N_9918);
nand U11621 (N_11621,N_8701,N_7997);
nand U11622 (N_11622,N_7640,N_8310);
or U11623 (N_11623,N_9127,N_9239);
nand U11624 (N_11624,N_9253,N_9277);
nor U11625 (N_11625,N_9708,N_7634);
and U11626 (N_11626,N_9029,N_8364);
or U11627 (N_11627,N_9971,N_9699);
and U11628 (N_11628,N_8953,N_7754);
and U11629 (N_11629,N_8310,N_8540);
nand U11630 (N_11630,N_8217,N_9818);
or U11631 (N_11631,N_8216,N_7624);
xnor U11632 (N_11632,N_8861,N_9841);
or U11633 (N_11633,N_7559,N_9455);
nand U11634 (N_11634,N_7645,N_7918);
nor U11635 (N_11635,N_9103,N_9466);
or U11636 (N_11636,N_8470,N_8920);
nand U11637 (N_11637,N_7786,N_8415);
nand U11638 (N_11638,N_7750,N_8279);
and U11639 (N_11639,N_9808,N_8602);
or U11640 (N_11640,N_8632,N_9509);
nand U11641 (N_11641,N_8454,N_9666);
nor U11642 (N_11642,N_9168,N_8764);
or U11643 (N_11643,N_9520,N_8931);
and U11644 (N_11644,N_7889,N_9047);
nand U11645 (N_11645,N_9282,N_9968);
nor U11646 (N_11646,N_7996,N_8385);
nand U11647 (N_11647,N_8453,N_8352);
nor U11648 (N_11648,N_9060,N_8115);
nand U11649 (N_11649,N_8278,N_9552);
nand U11650 (N_11650,N_9842,N_9475);
nand U11651 (N_11651,N_7798,N_9197);
and U11652 (N_11652,N_8987,N_8427);
or U11653 (N_11653,N_9740,N_8309);
and U11654 (N_11654,N_9906,N_8551);
and U11655 (N_11655,N_8953,N_9746);
and U11656 (N_11656,N_8421,N_7644);
nor U11657 (N_11657,N_7579,N_7998);
and U11658 (N_11658,N_7816,N_9319);
nand U11659 (N_11659,N_7715,N_8541);
or U11660 (N_11660,N_8714,N_8207);
nor U11661 (N_11661,N_8511,N_7876);
nand U11662 (N_11662,N_9477,N_8921);
or U11663 (N_11663,N_9261,N_8101);
nor U11664 (N_11664,N_8763,N_7955);
or U11665 (N_11665,N_8012,N_9407);
nor U11666 (N_11666,N_9452,N_7809);
nor U11667 (N_11667,N_9135,N_9052);
and U11668 (N_11668,N_8397,N_9212);
and U11669 (N_11669,N_9109,N_9119);
and U11670 (N_11670,N_9811,N_9806);
and U11671 (N_11671,N_8964,N_7937);
and U11672 (N_11672,N_8990,N_8089);
or U11673 (N_11673,N_8365,N_8449);
and U11674 (N_11674,N_9549,N_9611);
nor U11675 (N_11675,N_8976,N_8153);
and U11676 (N_11676,N_8925,N_8127);
or U11677 (N_11677,N_9417,N_8042);
or U11678 (N_11678,N_7872,N_9588);
or U11679 (N_11679,N_8117,N_9063);
or U11680 (N_11680,N_9217,N_8089);
nor U11681 (N_11681,N_9445,N_8406);
nor U11682 (N_11682,N_7621,N_9143);
and U11683 (N_11683,N_8296,N_8319);
or U11684 (N_11684,N_9210,N_9374);
nand U11685 (N_11685,N_9225,N_9977);
nand U11686 (N_11686,N_8802,N_7937);
nor U11687 (N_11687,N_9670,N_9184);
nand U11688 (N_11688,N_9879,N_9174);
and U11689 (N_11689,N_8804,N_9789);
nor U11690 (N_11690,N_8084,N_9024);
and U11691 (N_11691,N_7741,N_8434);
xor U11692 (N_11692,N_9250,N_9596);
nor U11693 (N_11693,N_8571,N_7603);
and U11694 (N_11694,N_7964,N_8163);
nand U11695 (N_11695,N_8783,N_8814);
and U11696 (N_11696,N_8941,N_8370);
nor U11697 (N_11697,N_9017,N_9752);
or U11698 (N_11698,N_9961,N_9179);
nor U11699 (N_11699,N_9959,N_8543);
and U11700 (N_11700,N_8743,N_8936);
nor U11701 (N_11701,N_9405,N_7769);
nor U11702 (N_11702,N_9288,N_7881);
and U11703 (N_11703,N_8065,N_7651);
or U11704 (N_11704,N_8516,N_8571);
or U11705 (N_11705,N_8268,N_9008);
and U11706 (N_11706,N_7882,N_8793);
nor U11707 (N_11707,N_7563,N_9888);
and U11708 (N_11708,N_9991,N_9910);
or U11709 (N_11709,N_8288,N_9235);
nor U11710 (N_11710,N_8423,N_9119);
xor U11711 (N_11711,N_8037,N_9773);
nand U11712 (N_11712,N_8006,N_8626);
nor U11713 (N_11713,N_8237,N_8338);
nand U11714 (N_11714,N_9554,N_9975);
and U11715 (N_11715,N_9039,N_8223);
nand U11716 (N_11716,N_9126,N_7613);
or U11717 (N_11717,N_7790,N_9657);
and U11718 (N_11718,N_9035,N_8606);
nand U11719 (N_11719,N_9640,N_9665);
nand U11720 (N_11720,N_9641,N_9772);
nor U11721 (N_11721,N_9205,N_7982);
nor U11722 (N_11722,N_8163,N_9008);
and U11723 (N_11723,N_7805,N_9622);
and U11724 (N_11724,N_8364,N_9967);
or U11725 (N_11725,N_8480,N_9220);
and U11726 (N_11726,N_9373,N_7928);
and U11727 (N_11727,N_9141,N_7937);
nand U11728 (N_11728,N_9988,N_9632);
and U11729 (N_11729,N_7903,N_9537);
nor U11730 (N_11730,N_9818,N_9311);
nor U11731 (N_11731,N_8847,N_9361);
or U11732 (N_11732,N_8064,N_7876);
or U11733 (N_11733,N_9061,N_8069);
nand U11734 (N_11734,N_9288,N_8218);
nand U11735 (N_11735,N_8060,N_8404);
nand U11736 (N_11736,N_8563,N_9969);
nand U11737 (N_11737,N_8726,N_8670);
nor U11738 (N_11738,N_7907,N_8501);
nand U11739 (N_11739,N_8219,N_9185);
nand U11740 (N_11740,N_9325,N_7573);
nand U11741 (N_11741,N_8187,N_8918);
and U11742 (N_11742,N_9384,N_9538);
and U11743 (N_11743,N_8630,N_8659);
or U11744 (N_11744,N_8752,N_8370);
or U11745 (N_11745,N_8439,N_7986);
nand U11746 (N_11746,N_9557,N_8167);
and U11747 (N_11747,N_9560,N_7707);
nand U11748 (N_11748,N_7531,N_9962);
or U11749 (N_11749,N_8890,N_8643);
and U11750 (N_11750,N_9518,N_9063);
and U11751 (N_11751,N_9180,N_8393);
xor U11752 (N_11752,N_7776,N_9782);
nor U11753 (N_11753,N_9553,N_9449);
nor U11754 (N_11754,N_9061,N_7560);
nand U11755 (N_11755,N_8035,N_9830);
and U11756 (N_11756,N_8212,N_9753);
nor U11757 (N_11757,N_9913,N_7848);
nor U11758 (N_11758,N_7648,N_9342);
and U11759 (N_11759,N_8386,N_7791);
nor U11760 (N_11760,N_8452,N_9979);
nand U11761 (N_11761,N_9218,N_9451);
nand U11762 (N_11762,N_9079,N_8274);
or U11763 (N_11763,N_9975,N_8119);
nor U11764 (N_11764,N_9199,N_9042);
nand U11765 (N_11765,N_8887,N_7809);
or U11766 (N_11766,N_8379,N_7802);
nand U11767 (N_11767,N_8485,N_8459);
nand U11768 (N_11768,N_9880,N_8743);
and U11769 (N_11769,N_9271,N_9289);
or U11770 (N_11770,N_9746,N_9065);
nand U11771 (N_11771,N_9252,N_8251);
nand U11772 (N_11772,N_8964,N_9825);
or U11773 (N_11773,N_8780,N_9926);
nand U11774 (N_11774,N_8037,N_9247);
nor U11775 (N_11775,N_9024,N_8531);
nor U11776 (N_11776,N_7911,N_9449);
or U11777 (N_11777,N_9926,N_8858);
and U11778 (N_11778,N_7785,N_9680);
or U11779 (N_11779,N_8488,N_7963);
or U11780 (N_11780,N_8502,N_8725);
nand U11781 (N_11781,N_8239,N_9426);
nor U11782 (N_11782,N_8623,N_9640);
or U11783 (N_11783,N_7866,N_8741);
and U11784 (N_11784,N_8905,N_8392);
or U11785 (N_11785,N_9375,N_7733);
nand U11786 (N_11786,N_8540,N_8631);
nor U11787 (N_11787,N_9461,N_7952);
nor U11788 (N_11788,N_9308,N_7819);
nand U11789 (N_11789,N_8819,N_9558);
and U11790 (N_11790,N_9904,N_8930);
nand U11791 (N_11791,N_9287,N_8567);
nor U11792 (N_11792,N_8003,N_9941);
and U11793 (N_11793,N_8707,N_8889);
nor U11794 (N_11794,N_9072,N_9317);
and U11795 (N_11795,N_9385,N_8750);
or U11796 (N_11796,N_7605,N_9365);
or U11797 (N_11797,N_8670,N_8086);
nand U11798 (N_11798,N_9179,N_9892);
or U11799 (N_11799,N_9859,N_7539);
nor U11800 (N_11800,N_7592,N_8562);
or U11801 (N_11801,N_9212,N_8641);
nor U11802 (N_11802,N_8767,N_9826);
and U11803 (N_11803,N_9596,N_9689);
and U11804 (N_11804,N_8335,N_9188);
or U11805 (N_11805,N_9292,N_9330);
or U11806 (N_11806,N_9760,N_8949);
and U11807 (N_11807,N_8332,N_9842);
or U11808 (N_11808,N_7651,N_8453);
nand U11809 (N_11809,N_9521,N_9939);
nand U11810 (N_11810,N_8399,N_9811);
nand U11811 (N_11811,N_9195,N_9267);
nand U11812 (N_11812,N_9231,N_9325);
nor U11813 (N_11813,N_7778,N_9502);
nor U11814 (N_11814,N_7955,N_8073);
and U11815 (N_11815,N_7709,N_8650);
or U11816 (N_11816,N_9822,N_9649);
and U11817 (N_11817,N_9690,N_9661);
nor U11818 (N_11818,N_8643,N_9214);
nor U11819 (N_11819,N_8648,N_8294);
nor U11820 (N_11820,N_9037,N_8367);
or U11821 (N_11821,N_9700,N_8063);
nand U11822 (N_11822,N_9565,N_7588);
or U11823 (N_11823,N_8391,N_9873);
nand U11824 (N_11824,N_9238,N_9297);
nor U11825 (N_11825,N_7598,N_9099);
nand U11826 (N_11826,N_9736,N_8155);
nand U11827 (N_11827,N_7964,N_7699);
or U11828 (N_11828,N_9365,N_9776);
xor U11829 (N_11829,N_8020,N_8331);
nor U11830 (N_11830,N_9933,N_8646);
nor U11831 (N_11831,N_9256,N_9300);
and U11832 (N_11832,N_7745,N_7819);
nor U11833 (N_11833,N_8768,N_8419);
nand U11834 (N_11834,N_9548,N_9111);
and U11835 (N_11835,N_8473,N_8477);
nor U11836 (N_11836,N_8926,N_9105);
nor U11837 (N_11837,N_9792,N_9299);
and U11838 (N_11838,N_7852,N_9267);
or U11839 (N_11839,N_9496,N_8218);
and U11840 (N_11840,N_9625,N_9364);
nand U11841 (N_11841,N_8318,N_7611);
nand U11842 (N_11842,N_8009,N_8441);
and U11843 (N_11843,N_8872,N_9473);
and U11844 (N_11844,N_9424,N_8264);
nand U11845 (N_11845,N_7634,N_7975);
and U11846 (N_11846,N_8406,N_8423);
and U11847 (N_11847,N_8082,N_7527);
nor U11848 (N_11848,N_7953,N_8808);
nor U11849 (N_11849,N_8057,N_8300);
nand U11850 (N_11850,N_9615,N_7648);
nand U11851 (N_11851,N_8404,N_8361);
nand U11852 (N_11852,N_8045,N_8769);
and U11853 (N_11853,N_9527,N_7771);
nand U11854 (N_11854,N_8856,N_8408);
and U11855 (N_11855,N_7886,N_8548);
or U11856 (N_11856,N_7709,N_8810);
or U11857 (N_11857,N_9477,N_9180);
nand U11858 (N_11858,N_7875,N_9675);
nand U11859 (N_11859,N_7660,N_9106);
xor U11860 (N_11860,N_9357,N_8354);
nor U11861 (N_11861,N_8562,N_8146);
nand U11862 (N_11862,N_7849,N_8538);
nand U11863 (N_11863,N_9958,N_8932);
and U11864 (N_11864,N_8366,N_9658);
or U11865 (N_11865,N_7875,N_8136);
or U11866 (N_11866,N_8850,N_8046);
nor U11867 (N_11867,N_9905,N_9475);
nand U11868 (N_11868,N_8023,N_7772);
and U11869 (N_11869,N_7685,N_7513);
or U11870 (N_11870,N_8440,N_9683);
and U11871 (N_11871,N_7885,N_9736);
or U11872 (N_11872,N_8781,N_8828);
nand U11873 (N_11873,N_7507,N_8147);
or U11874 (N_11874,N_9350,N_7791);
nand U11875 (N_11875,N_9743,N_8682);
or U11876 (N_11876,N_7608,N_8249);
nand U11877 (N_11877,N_8124,N_8740);
or U11878 (N_11878,N_9462,N_9565);
nor U11879 (N_11879,N_7659,N_9128);
nand U11880 (N_11880,N_9065,N_9624);
or U11881 (N_11881,N_8185,N_9276);
nand U11882 (N_11882,N_7569,N_9752);
or U11883 (N_11883,N_8091,N_7796);
or U11884 (N_11884,N_8813,N_7723);
nor U11885 (N_11885,N_9799,N_7896);
and U11886 (N_11886,N_7661,N_7786);
nand U11887 (N_11887,N_9964,N_8956);
nand U11888 (N_11888,N_8455,N_9227);
nor U11889 (N_11889,N_8387,N_8377);
or U11890 (N_11890,N_8987,N_9030);
nand U11891 (N_11891,N_7710,N_9177);
nand U11892 (N_11892,N_9160,N_7823);
and U11893 (N_11893,N_9519,N_7894);
and U11894 (N_11894,N_8946,N_9762);
and U11895 (N_11895,N_9674,N_8748);
or U11896 (N_11896,N_7962,N_8810);
nand U11897 (N_11897,N_9387,N_8611);
and U11898 (N_11898,N_8735,N_8034);
or U11899 (N_11899,N_9469,N_7927);
and U11900 (N_11900,N_8529,N_7839);
or U11901 (N_11901,N_9907,N_9333);
nand U11902 (N_11902,N_8592,N_8956);
and U11903 (N_11903,N_9473,N_8387);
and U11904 (N_11904,N_9766,N_8210);
nand U11905 (N_11905,N_8636,N_9858);
or U11906 (N_11906,N_9929,N_8463);
nand U11907 (N_11907,N_9684,N_7996);
or U11908 (N_11908,N_9633,N_9609);
or U11909 (N_11909,N_7922,N_8145);
or U11910 (N_11910,N_8903,N_8840);
or U11911 (N_11911,N_8024,N_8016);
or U11912 (N_11912,N_8962,N_7928);
or U11913 (N_11913,N_9379,N_9311);
and U11914 (N_11914,N_9034,N_8231);
or U11915 (N_11915,N_9449,N_8439);
nand U11916 (N_11916,N_8510,N_8981);
nor U11917 (N_11917,N_9829,N_7828);
and U11918 (N_11918,N_9819,N_9178);
or U11919 (N_11919,N_9699,N_7513);
nor U11920 (N_11920,N_7853,N_9873);
or U11921 (N_11921,N_7817,N_8368);
nand U11922 (N_11922,N_9879,N_8652);
nor U11923 (N_11923,N_9974,N_7621);
or U11924 (N_11924,N_9277,N_8330);
nand U11925 (N_11925,N_9490,N_9983);
nand U11926 (N_11926,N_8312,N_9294);
or U11927 (N_11927,N_7763,N_9695);
and U11928 (N_11928,N_7646,N_9512);
or U11929 (N_11929,N_8551,N_8583);
nor U11930 (N_11930,N_8565,N_8148);
nand U11931 (N_11931,N_9751,N_8012);
and U11932 (N_11932,N_8007,N_8489);
nor U11933 (N_11933,N_8977,N_9830);
and U11934 (N_11934,N_9383,N_8686);
or U11935 (N_11935,N_9361,N_8793);
nand U11936 (N_11936,N_8463,N_9175);
nand U11937 (N_11937,N_7904,N_7788);
nand U11938 (N_11938,N_9265,N_7883);
or U11939 (N_11939,N_8057,N_8336);
or U11940 (N_11940,N_8776,N_9651);
or U11941 (N_11941,N_9562,N_9312);
nor U11942 (N_11942,N_9416,N_8623);
or U11943 (N_11943,N_9653,N_9278);
nor U11944 (N_11944,N_8362,N_8150);
nor U11945 (N_11945,N_9918,N_8056);
nor U11946 (N_11946,N_9704,N_9590);
nor U11947 (N_11947,N_9542,N_9120);
or U11948 (N_11948,N_7968,N_8489);
nor U11949 (N_11949,N_8714,N_9239);
nor U11950 (N_11950,N_8224,N_9283);
nor U11951 (N_11951,N_8089,N_8760);
or U11952 (N_11952,N_8898,N_9773);
and U11953 (N_11953,N_8884,N_8591);
and U11954 (N_11954,N_8259,N_9625);
or U11955 (N_11955,N_9422,N_9538);
and U11956 (N_11956,N_9475,N_8283);
and U11957 (N_11957,N_8613,N_8884);
nor U11958 (N_11958,N_8604,N_9712);
and U11959 (N_11959,N_9351,N_8948);
nand U11960 (N_11960,N_9880,N_8861);
nor U11961 (N_11961,N_8143,N_9757);
and U11962 (N_11962,N_8108,N_7943);
or U11963 (N_11963,N_9083,N_7757);
nor U11964 (N_11964,N_9932,N_7856);
nand U11965 (N_11965,N_9486,N_8759);
or U11966 (N_11966,N_7591,N_7737);
nand U11967 (N_11967,N_9923,N_7631);
nor U11968 (N_11968,N_9728,N_8332);
or U11969 (N_11969,N_9263,N_9330);
nand U11970 (N_11970,N_9993,N_9605);
nand U11971 (N_11971,N_8866,N_8421);
nand U11972 (N_11972,N_7853,N_9903);
nand U11973 (N_11973,N_9272,N_8542);
and U11974 (N_11974,N_8679,N_9066);
and U11975 (N_11975,N_8246,N_7531);
or U11976 (N_11976,N_9775,N_8570);
or U11977 (N_11977,N_9402,N_9766);
or U11978 (N_11978,N_7623,N_9436);
and U11979 (N_11979,N_8184,N_9530);
nor U11980 (N_11980,N_9454,N_8119);
nand U11981 (N_11981,N_8076,N_9541);
nor U11982 (N_11982,N_7698,N_9036);
or U11983 (N_11983,N_8535,N_8138);
and U11984 (N_11984,N_9727,N_8675);
nor U11985 (N_11985,N_8247,N_7546);
nand U11986 (N_11986,N_7772,N_8792);
nand U11987 (N_11987,N_9616,N_7719);
or U11988 (N_11988,N_9387,N_9562);
nor U11989 (N_11989,N_8900,N_8076);
and U11990 (N_11990,N_9156,N_8527);
or U11991 (N_11991,N_8737,N_9366);
nor U11992 (N_11992,N_9423,N_8625);
or U11993 (N_11993,N_9620,N_8188);
nand U11994 (N_11994,N_8462,N_9650);
and U11995 (N_11995,N_8238,N_7821);
or U11996 (N_11996,N_9411,N_9908);
nand U11997 (N_11997,N_9442,N_9700);
nand U11998 (N_11998,N_8907,N_9773);
nand U11999 (N_11999,N_8099,N_8483);
nand U12000 (N_12000,N_8595,N_7683);
or U12001 (N_12001,N_9990,N_9819);
and U12002 (N_12002,N_8424,N_7681);
or U12003 (N_12003,N_8270,N_9433);
or U12004 (N_12004,N_8376,N_7956);
nand U12005 (N_12005,N_9686,N_7985);
nor U12006 (N_12006,N_9630,N_8747);
and U12007 (N_12007,N_8846,N_9144);
nor U12008 (N_12008,N_7655,N_9225);
or U12009 (N_12009,N_9917,N_7719);
nand U12010 (N_12010,N_8801,N_8204);
xor U12011 (N_12011,N_8590,N_8322);
and U12012 (N_12012,N_8593,N_7727);
nand U12013 (N_12013,N_9712,N_8096);
and U12014 (N_12014,N_8103,N_9612);
and U12015 (N_12015,N_9528,N_8253);
or U12016 (N_12016,N_8606,N_8142);
nor U12017 (N_12017,N_8228,N_8489);
nand U12018 (N_12018,N_8245,N_7890);
nor U12019 (N_12019,N_9407,N_8088);
or U12020 (N_12020,N_8276,N_7605);
or U12021 (N_12021,N_8941,N_7889);
and U12022 (N_12022,N_8665,N_8256);
nor U12023 (N_12023,N_9151,N_8390);
or U12024 (N_12024,N_8302,N_8436);
and U12025 (N_12025,N_8440,N_8789);
nand U12026 (N_12026,N_8110,N_9187);
nor U12027 (N_12027,N_9476,N_8345);
or U12028 (N_12028,N_7809,N_8745);
nor U12029 (N_12029,N_8670,N_9596);
nor U12030 (N_12030,N_8438,N_8106);
nand U12031 (N_12031,N_8641,N_7596);
or U12032 (N_12032,N_9020,N_9355);
nor U12033 (N_12033,N_8834,N_9918);
nand U12034 (N_12034,N_7770,N_7709);
nand U12035 (N_12035,N_9796,N_9880);
nor U12036 (N_12036,N_9044,N_9582);
or U12037 (N_12037,N_8136,N_9900);
and U12038 (N_12038,N_7939,N_8188);
nor U12039 (N_12039,N_8610,N_7806);
nor U12040 (N_12040,N_8585,N_9082);
nand U12041 (N_12041,N_8289,N_9441);
or U12042 (N_12042,N_9809,N_8754);
or U12043 (N_12043,N_9704,N_8593);
nor U12044 (N_12044,N_9968,N_8579);
and U12045 (N_12045,N_9634,N_9081);
and U12046 (N_12046,N_9144,N_9801);
nand U12047 (N_12047,N_9443,N_7615);
nand U12048 (N_12048,N_9960,N_9751);
or U12049 (N_12049,N_9401,N_8936);
nand U12050 (N_12050,N_8184,N_7695);
nor U12051 (N_12051,N_9631,N_8044);
nor U12052 (N_12052,N_7845,N_7995);
or U12053 (N_12053,N_8709,N_8296);
or U12054 (N_12054,N_8564,N_9323);
nor U12055 (N_12055,N_7766,N_9451);
or U12056 (N_12056,N_9368,N_7707);
xor U12057 (N_12057,N_8836,N_9150);
nor U12058 (N_12058,N_7960,N_9828);
and U12059 (N_12059,N_9037,N_9475);
and U12060 (N_12060,N_9398,N_8945);
or U12061 (N_12061,N_9783,N_8101);
nor U12062 (N_12062,N_7782,N_8782);
or U12063 (N_12063,N_8462,N_9141);
nand U12064 (N_12064,N_9207,N_9616);
nor U12065 (N_12065,N_8956,N_7542);
and U12066 (N_12066,N_9662,N_7679);
nor U12067 (N_12067,N_7887,N_7765);
or U12068 (N_12068,N_9288,N_7758);
and U12069 (N_12069,N_8734,N_7609);
nor U12070 (N_12070,N_9331,N_8266);
nand U12071 (N_12071,N_8342,N_9100);
nor U12072 (N_12072,N_8636,N_8471);
and U12073 (N_12073,N_9730,N_7809);
and U12074 (N_12074,N_7951,N_8402);
nand U12075 (N_12075,N_9898,N_8752);
and U12076 (N_12076,N_8670,N_9378);
and U12077 (N_12077,N_8384,N_8183);
nor U12078 (N_12078,N_9022,N_9766);
and U12079 (N_12079,N_9448,N_9377);
nor U12080 (N_12080,N_8922,N_7863);
nand U12081 (N_12081,N_7998,N_8274);
nor U12082 (N_12082,N_7617,N_8963);
or U12083 (N_12083,N_7741,N_8133);
or U12084 (N_12084,N_8392,N_9875);
and U12085 (N_12085,N_9483,N_8009);
or U12086 (N_12086,N_9647,N_7645);
xnor U12087 (N_12087,N_8694,N_9604);
nor U12088 (N_12088,N_8749,N_7752);
nand U12089 (N_12089,N_8981,N_8982);
nor U12090 (N_12090,N_8068,N_7726);
nand U12091 (N_12091,N_7956,N_8095);
nor U12092 (N_12092,N_9590,N_9759);
nor U12093 (N_12093,N_9663,N_9116);
nand U12094 (N_12094,N_8953,N_9463);
or U12095 (N_12095,N_7787,N_8324);
or U12096 (N_12096,N_8951,N_7885);
xnor U12097 (N_12097,N_7859,N_8497);
nand U12098 (N_12098,N_8534,N_7888);
nand U12099 (N_12099,N_8025,N_8592);
nor U12100 (N_12100,N_9495,N_9576);
nand U12101 (N_12101,N_8627,N_8779);
or U12102 (N_12102,N_9332,N_9437);
nand U12103 (N_12103,N_9536,N_7847);
or U12104 (N_12104,N_9944,N_8308);
or U12105 (N_12105,N_9537,N_9346);
and U12106 (N_12106,N_7714,N_9774);
nand U12107 (N_12107,N_7578,N_9677);
or U12108 (N_12108,N_9586,N_8453);
and U12109 (N_12109,N_7564,N_9778);
and U12110 (N_12110,N_8692,N_8541);
and U12111 (N_12111,N_8458,N_7701);
nand U12112 (N_12112,N_9079,N_9033);
or U12113 (N_12113,N_8868,N_7767);
nor U12114 (N_12114,N_9827,N_7510);
nand U12115 (N_12115,N_9719,N_9706);
nor U12116 (N_12116,N_9093,N_7992);
and U12117 (N_12117,N_8245,N_8438);
or U12118 (N_12118,N_8383,N_8237);
and U12119 (N_12119,N_8836,N_8626);
nand U12120 (N_12120,N_9691,N_7762);
nand U12121 (N_12121,N_9475,N_7942);
or U12122 (N_12122,N_8808,N_8717);
and U12123 (N_12123,N_9004,N_9024);
and U12124 (N_12124,N_8635,N_7571);
nor U12125 (N_12125,N_9239,N_7786);
and U12126 (N_12126,N_9204,N_8543);
and U12127 (N_12127,N_9311,N_7990);
or U12128 (N_12128,N_8587,N_9446);
or U12129 (N_12129,N_9043,N_9134);
or U12130 (N_12130,N_7743,N_9003);
nand U12131 (N_12131,N_9741,N_8959);
or U12132 (N_12132,N_8455,N_9715);
nor U12133 (N_12133,N_8049,N_8520);
nand U12134 (N_12134,N_7600,N_9993);
nand U12135 (N_12135,N_8172,N_7508);
or U12136 (N_12136,N_9191,N_7788);
nor U12137 (N_12137,N_7922,N_9453);
nor U12138 (N_12138,N_8463,N_8592);
or U12139 (N_12139,N_8880,N_9653);
or U12140 (N_12140,N_9789,N_7768);
nand U12141 (N_12141,N_8569,N_9216);
nor U12142 (N_12142,N_9804,N_8965);
and U12143 (N_12143,N_9792,N_9060);
nand U12144 (N_12144,N_7625,N_7812);
and U12145 (N_12145,N_8719,N_8306);
nor U12146 (N_12146,N_7669,N_9682);
and U12147 (N_12147,N_7980,N_8411);
nor U12148 (N_12148,N_9211,N_7646);
nor U12149 (N_12149,N_9000,N_8258);
or U12150 (N_12150,N_9434,N_7934);
nor U12151 (N_12151,N_7810,N_7858);
or U12152 (N_12152,N_7837,N_7758);
or U12153 (N_12153,N_7527,N_9627);
xnor U12154 (N_12154,N_8796,N_9190);
or U12155 (N_12155,N_8015,N_7642);
nor U12156 (N_12156,N_9666,N_9253);
nand U12157 (N_12157,N_9348,N_9860);
nor U12158 (N_12158,N_9071,N_9872);
nand U12159 (N_12159,N_8748,N_7981);
nand U12160 (N_12160,N_9427,N_8230);
and U12161 (N_12161,N_8199,N_8054);
or U12162 (N_12162,N_8561,N_9197);
nor U12163 (N_12163,N_8975,N_9215);
and U12164 (N_12164,N_8352,N_9154);
or U12165 (N_12165,N_8817,N_8475);
nor U12166 (N_12166,N_7700,N_9161);
and U12167 (N_12167,N_8197,N_7954);
or U12168 (N_12168,N_8821,N_7899);
nand U12169 (N_12169,N_9763,N_8150);
and U12170 (N_12170,N_9157,N_7593);
or U12171 (N_12171,N_9116,N_8379);
and U12172 (N_12172,N_7943,N_8624);
and U12173 (N_12173,N_9969,N_9796);
and U12174 (N_12174,N_8026,N_7979);
nand U12175 (N_12175,N_9704,N_8355);
nand U12176 (N_12176,N_9972,N_9971);
nor U12177 (N_12177,N_9671,N_9568);
or U12178 (N_12178,N_9212,N_8542);
or U12179 (N_12179,N_7546,N_9655);
and U12180 (N_12180,N_8814,N_9679);
and U12181 (N_12181,N_8334,N_9359);
and U12182 (N_12182,N_7986,N_9398);
and U12183 (N_12183,N_8087,N_7996);
nand U12184 (N_12184,N_9448,N_7664);
nand U12185 (N_12185,N_9678,N_8896);
nor U12186 (N_12186,N_9596,N_7969);
or U12187 (N_12187,N_7775,N_8081);
and U12188 (N_12188,N_7550,N_8830);
nand U12189 (N_12189,N_8995,N_8143);
or U12190 (N_12190,N_8055,N_9779);
and U12191 (N_12191,N_7898,N_8072);
or U12192 (N_12192,N_8993,N_9621);
nand U12193 (N_12193,N_8095,N_7693);
and U12194 (N_12194,N_7940,N_8911);
and U12195 (N_12195,N_8504,N_9896);
nand U12196 (N_12196,N_8139,N_9076);
and U12197 (N_12197,N_9513,N_9744);
or U12198 (N_12198,N_9925,N_9884);
or U12199 (N_12199,N_8623,N_9392);
nor U12200 (N_12200,N_8095,N_7690);
nor U12201 (N_12201,N_9522,N_8865);
nand U12202 (N_12202,N_9129,N_8049);
nand U12203 (N_12203,N_8701,N_9984);
nor U12204 (N_12204,N_8732,N_8418);
or U12205 (N_12205,N_8076,N_9442);
and U12206 (N_12206,N_9873,N_9984);
or U12207 (N_12207,N_8114,N_8102);
and U12208 (N_12208,N_8476,N_9930);
nor U12209 (N_12209,N_9533,N_8503);
nor U12210 (N_12210,N_9559,N_8791);
nor U12211 (N_12211,N_9049,N_9906);
nor U12212 (N_12212,N_8147,N_7749);
and U12213 (N_12213,N_7764,N_7622);
and U12214 (N_12214,N_8194,N_8727);
nor U12215 (N_12215,N_7737,N_9381);
and U12216 (N_12216,N_7741,N_8363);
nand U12217 (N_12217,N_8643,N_7756);
and U12218 (N_12218,N_7902,N_7934);
or U12219 (N_12219,N_9291,N_9732);
nand U12220 (N_12220,N_9999,N_7717);
and U12221 (N_12221,N_8887,N_9442);
nor U12222 (N_12222,N_9726,N_9470);
and U12223 (N_12223,N_9315,N_9711);
nand U12224 (N_12224,N_8231,N_7928);
nor U12225 (N_12225,N_9949,N_9764);
xor U12226 (N_12226,N_9611,N_8264);
nand U12227 (N_12227,N_8973,N_9103);
nor U12228 (N_12228,N_9640,N_9047);
or U12229 (N_12229,N_9638,N_9352);
nor U12230 (N_12230,N_8337,N_9298);
and U12231 (N_12231,N_9052,N_9232);
nor U12232 (N_12232,N_7681,N_9117);
nor U12233 (N_12233,N_8187,N_9214);
and U12234 (N_12234,N_8280,N_8200);
xor U12235 (N_12235,N_9516,N_7829);
or U12236 (N_12236,N_8334,N_7988);
nand U12237 (N_12237,N_8605,N_8770);
nor U12238 (N_12238,N_9049,N_8842);
nor U12239 (N_12239,N_9815,N_9605);
nand U12240 (N_12240,N_9101,N_7800);
or U12241 (N_12241,N_9574,N_8296);
nand U12242 (N_12242,N_7877,N_8311);
nor U12243 (N_12243,N_9670,N_9364);
nand U12244 (N_12244,N_8271,N_7880);
nor U12245 (N_12245,N_9421,N_9427);
nand U12246 (N_12246,N_8078,N_8536);
nor U12247 (N_12247,N_8223,N_9379);
or U12248 (N_12248,N_9524,N_8970);
and U12249 (N_12249,N_8879,N_9663);
and U12250 (N_12250,N_9978,N_9476);
nor U12251 (N_12251,N_8271,N_7576);
and U12252 (N_12252,N_8320,N_8631);
nor U12253 (N_12253,N_7773,N_8146);
nor U12254 (N_12254,N_7585,N_9418);
nand U12255 (N_12255,N_8439,N_9495);
and U12256 (N_12256,N_7661,N_8135);
and U12257 (N_12257,N_8454,N_8343);
or U12258 (N_12258,N_9072,N_9957);
or U12259 (N_12259,N_9560,N_9714);
or U12260 (N_12260,N_9310,N_9126);
nand U12261 (N_12261,N_7837,N_9899);
nor U12262 (N_12262,N_8546,N_9469);
and U12263 (N_12263,N_7986,N_9065);
and U12264 (N_12264,N_9518,N_8708);
and U12265 (N_12265,N_9468,N_7595);
nand U12266 (N_12266,N_7640,N_9792);
nand U12267 (N_12267,N_9410,N_8061);
or U12268 (N_12268,N_9168,N_8975);
nand U12269 (N_12269,N_9275,N_9506);
or U12270 (N_12270,N_7822,N_8887);
nor U12271 (N_12271,N_9126,N_8857);
and U12272 (N_12272,N_7548,N_9199);
nor U12273 (N_12273,N_8541,N_9662);
or U12274 (N_12274,N_9553,N_8708);
nor U12275 (N_12275,N_8328,N_8953);
or U12276 (N_12276,N_7785,N_8031);
nor U12277 (N_12277,N_9332,N_7981);
and U12278 (N_12278,N_7586,N_9844);
and U12279 (N_12279,N_8559,N_9503);
or U12280 (N_12280,N_8500,N_8803);
or U12281 (N_12281,N_8704,N_7534);
nor U12282 (N_12282,N_8145,N_9380);
or U12283 (N_12283,N_8062,N_8349);
or U12284 (N_12284,N_7780,N_7948);
or U12285 (N_12285,N_9027,N_9594);
and U12286 (N_12286,N_7687,N_9751);
or U12287 (N_12287,N_9983,N_9873);
and U12288 (N_12288,N_9743,N_8944);
or U12289 (N_12289,N_8611,N_8019);
or U12290 (N_12290,N_8667,N_9520);
or U12291 (N_12291,N_8503,N_8693);
nand U12292 (N_12292,N_7706,N_8263);
and U12293 (N_12293,N_8222,N_7621);
and U12294 (N_12294,N_9302,N_7902);
nor U12295 (N_12295,N_9666,N_7629);
and U12296 (N_12296,N_9013,N_8941);
nor U12297 (N_12297,N_8083,N_9427);
nand U12298 (N_12298,N_7993,N_7774);
and U12299 (N_12299,N_9228,N_8030);
nand U12300 (N_12300,N_9497,N_8549);
nand U12301 (N_12301,N_9806,N_8150);
nand U12302 (N_12302,N_7661,N_9059);
nand U12303 (N_12303,N_7581,N_9457);
or U12304 (N_12304,N_9726,N_9166);
nor U12305 (N_12305,N_8448,N_9084);
or U12306 (N_12306,N_7500,N_9461);
nand U12307 (N_12307,N_9646,N_7569);
nand U12308 (N_12308,N_8369,N_8309);
and U12309 (N_12309,N_8821,N_8640);
xor U12310 (N_12310,N_9880,N_9922);
nand U12311 (N_12311,N_9277,N_8848);
or U12312 (N_12312,N_7815,N_8999);
nor U12313 (N_12313,N_9789,N_7634);
and U12314 (N_12314,N_9121,N_8858);
nand U12315 (N_12315,N_8057,N_9564);
nand U12316 (N_12316,N_9048,N_9743);
or U12317 (N_12317,N_7512,N_8521);
nor U12318 (N_12318,N_8085,N_7948);
nand U12319 (N_12319,N_9010,N_9663);
or U12320 (N_12320,N_9330,N_8887);
or U12321 (N_12321,N_9116,N_8824);
nand U12322 (N_12322,N_9086,N_8919);
nor U12323 (N_12323,N_9319,N_8710);
and U12324 (N_12324,N_9449,N_8604);
nand U12325 (N_12325,N_9336,N_8086);
nand U12326 (N_12326,N_7874,N_8558);
nand U12327 (N_12327,N_7926,N_8893);
and U12328 (N_12328,N_8515,N_8711);
xnor U12329 (N_12329,N_8759,N_9636);
and U12330 (N_12330,N_7564,N_8207);
nor U12331 (N_12331,N_9887,N_7545);
nand U12332 (N_12332,N_9446,N_9989);
nand U12333 (N_12333,N_8549,N_9823);
or U12334 (N_12334,N_9594,N_7773);
nor U12335 (N_12335,N_8836,N_9197);
and U12336 (N_12336,N_8052,N_8387);
nand U12337 (N_12337,N_8591,N_8519);
and U12338 (N_12338,N_7669,N_8703);
nor U12339 (N_12339,N_8387,N_8969);
nor U12340 (N_12340,N_8606,N_9280);
nand U12341 (N_12341,N_9590,N_9575);
nand U12342 (N_12342,N_8330,N_8687);
and U12343 (N_12343,N_9253,N_8583);
or U12344 (N_12344,N_9262,N_9500);
and U12345 (N_12345,N_8305,N_8917);
or U12346 (N_12346,N_8169,N_9028);
and U12347 (N_12347,N_8879,N_7664);
nand U12348 (N_12348,N_8777,N_9022);
nand U12349 (N_12349,N_8962,N_9114);
nor U12350 (N_12350,N_7774,N_9414);
nor U12351 (N_12351,N_7514,N_8668);
and U12352 (N_12352,N_9064,N_9084);
nor U12353 (N_12353,N_9979,N_9222);
or U12354 (N_12354,N_9831,N_8842);
and U12355 (N_12355,N_8906,N_8111);
nand U12356 (N_12356,N_8543,N_8072);
and U12357 (N_12357,N_9116,N_7912);
and U12358 (N_12358,N_7743,N_9104);
nor U12359 (N_12359,N_9191,N_9425);
and U12360 (N_12360,N_8508,N_9260);
and U12361 (N_12361,N_9130,N_9693);
or U12362 (N_12362,N_7584,N_8978);
nor U12363 (N_12363,N_7933,N_8453);
nor U12364 (N_12364,N_8353,N_9379);
and U12365 (N_12365,N_8502,N_8303);
and U12366 (N_12366,N_9587,N_8295);
nor U12367 (N_12367,N_9049,N_7657);
and U12368 (N_12368,N_7640,N_8380);
nand U12369 (N_12369,N_8195,N_9404);
nand U12370 (N_12370,N_8538,N_9352);
and U12371 (N_12371,N_7775,N_8124);
and U12372 (N_12372,N_7952,N_9679);
or U12373 (N_12373,N_9448,N_9571);
and U12374 (N_12374,N_9174,N_8297);
or U12375 (N_12375,N_9263,N_8807);
and U12376 (N_12376,N_9234,N_8050);
or U12377 (N_12377,N_9207,N_9727);
and U12378 (N_12378,N_7906,N_9985);
or U12379 (N_12379,N_8039,N_8324);
or U12380 (N_12380,N_8105,N_9404);
nand U12381 (N_12381,N_9578,N_9485);
or U12382 (N_12382,N_8779,N_7853);
and U12383 (N_12383,N_8801,N_8137);
and U12384 (N_12384,N_9091,N_9703);
or U12385 (N_12385,N_9115,N_8380);
nand U12386 (N_12386,N_8891,N_9524);
nor U12387 (N_12387,N_8797,N_9523);
or U12388 (N_12388,N_9038,N_7967);
nor U12389 (N_12389,N_9922,N_8862);
or U12390 (N_12390,N_9731,N_9006);
and U12391 (N_12391,N_8274,N_7808);
nor U12392 (N_12392,N_9384,N_8469);
nor U12393 (N_12393,N_7567,N_8431);
nand U12394 (N_12394,N_9981,N_9880);
nor U12395 (N_12395,N_9368,N_9917);
nor U12396 (N_12396,N_8142,N_9322);
nand U12397 (N_12397,N_8253,N_8418);
and U12398 (N_12398,N_8476,N_9213);
nor U12399 (N_12399,N_7779,N_7630);
nor U12400 (N_12400,N_8963,N_8871);
nand U12401 (N_12401,N_7722,N_8832);
and U12402 (N_12402,N_7555,N_8403);
or U12403 (N_12403,N_8743,N_9138);
nand U12404 (N_12404,N_9845,N_9513);
or U12405 (N_12405,N_8970,N_9458);
nor U12406 (N_12406,N_9576,N_7723);
and U12407 (N_12407,N_9548,N_9619);
and U12408 (N_12408,N_9405,N_9312);
nand U12409 (N_12409,N_7747,N_9332);
or U12410 (N_12410,N_7959,N_8580);
or U12411 (N_12411,N_7711,N_8325);
and U12412 (N_12412,N_8961,N_7893);
nor U12413 (N_12413,N_9971,N_9213);
nand U12414 (N_12414,N_7854,N_9383);
nor U12415 (N_12415,N_9891,N_8582);
and U12416 (N_12416,N_8449,N_9447);
nor U12417 (N_12417,N_7631,N_8840);
and U12418 (N_12418,N_8892,N_8093);
nor U12419 (N_12419,N_8406,N_8925);
or U12420 (N_12420,N_8037,N_8260);
or U12421 (N_12421,N_8517,N_9752);
nand U12422 (N_12422,N_9819,N_8014);
nand U12423 (N_12423,N_9364,N_7579);
or U12424 (N_12424,N_9248,N_9325);
nor U12425 (N_12425,N_9681,N_8494);
nor U12426 (N_12426,N_9297,N_8511);
and U12427 (N_12427,N_8752,N_9825);
or U12428 (N_12428,N_8030,N_8590);
and U12429 (N_12429,N_7616,N_9049);
and U12430 (N_12430,N_7571,N_9619);
nor U12431 (N_12431,N_8505,N_9555);
and U12432 (N_12432,N_8952,N_8664);
nand U12433 (N_12433,N_9499,N_7817);
and U12434 (N_12434,N_8359,N_8007);
or U12435 (N_12435,N_7992,N_8226);
and U12436 (N_12436,N_8654,N_7882);
and U12437 (N_12437,N_9746,N_9558);
nand U12438 (N_12438,N_7785,N_7609);
or U12439 (N_12439,N_8349,N_9170);
or U12440 (N_12440,N_9012,N_9679);
nand U12441 (N_12441,N_8467,N_9219);
nand U12442 (N_12442,N_8375,N_7604);
and U12443 (N_12443,N_9442,N_7871);
nor U12444 (N_12444,N_8506,N_8504);
or U12445 (N_12445,N_9659,N_7842);
or U12446 (N_12446,N_8011,N_7930);
nand U12447 (N_12447,N_8575,N_8025);
or U12448 (N_12448,N_8900,N_7598);
or U12449 (N_12449,N_8580,N_8010);
nor U12450 (N_12450,N_8156,N_9102);
nand U12451 (N_12451,N_8760,N_9276);
and U12452 (N_12452,N_9218,N_8670);
or U12453 (N_12453,N_9886,N_9109);
or U12454 (N_12454,N_8531,N_7763);
nor U12455 (N_12455,N_8888,N_8510);
nor U12456 (N_12456,N_7885,N_7644);
nand U12457 (N_12457,N_9538,N_8371);
xor U12458 (N_12458,N_9229,N_8246);
or U12459 (N_12459,N_9399,N_9417);
or U12460 (N_12460,N_8636,N_9237);
or U12461 (N_12461,N_7525,N_8397);
and U12462 (N_12462,N_8913,N_8703);
nand U12463 (N_12463,N_8637,N_9044);
or U12464 (N_12464,N_7689,N_8967);
and U12465 (N_12465,N_9851,N_9920);
or U12466 (N_12466,N_9753,N_7882);
nor U12467 (N_12467,N_9013,N_9654);
nor U12468 (N_12468,N_8731,N_8670);
nor U12469 (N_12469,N_9575,N_9980);
and U12470 (N_12470,N_8634,N_9436);
nor U12471 (N_12471,N_8171,N_8506);
and U12472 (N_12472,N_8063,N_9939);
nor U12473 (N_12473,N_9934,N_8056);
nand U12474 (N_12474,N_7678,N_9863);
nor U12475 (N_12475,N_8490,N_7870);
nand U12476 (N_12476,N_8695,N_8360);
and U12477 (N_12477,N_8443,N_8410);
nand U12478 (N_12478,N_8248,N_9519);
nand U12479 (N_12479,N_9149,N_8400);
and U12480 (N_12480,N_7938,N_9134);
nor U12481 (N_12481,N_7668,N_7717);
nand U12482 (N_12482,N_7753,N_9715);
or U12483 (N_12483,N_8254,N_8833);
and U12484 (N_12484,N_8934,N_9018);
nor U12485 (N_12485,N_9974,N_8007);
or U12486 (N_12486,N_8154,N_9187);
nor U12487 (N_12487,N_7765,N_7685);
nand U12488 (N_12488,N_9347,N_8396);
nor U12489 (N_12489,N_8887,N_8841);
nor U12490 (N_12490,N_9849,N_8951);
nand U12491 (N_12491,N_8146,N_9202);
and U12492 (N_12492,N_9260,N_8786);
or U12493 (N_12493,N_9483,N_8495);
nor U12494 (N_12494,N_9669,N_8161);
nand U12495 (N_12495,N_7728,N_8133);
and U12496 (N_12496,N_9705,N_9246);
and U12497 (N_12497,N_9326,N_9922);
and U12498 (N_12498,N_8900,N_9015);
nand U12499 (N_12499,N_9573,N_8551);
nand U12500 (N_12500,N_10475,N_10902);
nor U12501 (N_12501,N_12283,N_11425);
or U12502 (N_12502,N_10380,N_11165);
nand U12503 (N_12503,N_10495,N_10656);
or U12504 (N_12504,N_10825,N_10006);
nand U12505 (N_12505,N_10402,N_11399);
xnor U12506 (N_12506,N_12118,N_12474);
or U12507 (N_12507,N_10239,N_10878);
nor U12508 (N_12508,N_10839,N_11078);
or U12509 (N_12509,N_11680,N_10954);
nand U12510 (N_12510,N_12137,N_11777);
or U12511 (N_12511,N_10057,N_11660);
or U12512 (N_12512,N_11297,N_12237);
and U12513 (N_12513,N_11008,N_11267);
nand U12514 (N_12514,N_12451,N_12444);
nand U12515 (N_12515,N_10214,N_11772);
nor U12516 (N_12516,N_11367,N_11100);
and U12517 (N_12517,N_10225,N_10833);
nand U12518 (N_12518,N_10769,N_10453);
nor U12519 (N_12519,N_11606,N_11403);
xnor U12520 (N_12520,N_10981,N_12420);
or U12521 (N_12521,N_10976,N_12262);
and U12522 (N_12522,N_10900,N_12472);
nand U12523 (N_12523,N_10032,N_11433);
and U12524 (N_12524,N_10562,N_12167);
and U12525 (N_12525,N_10428,N_11511);
nor U12526 (N_12526,N_10369,N_10560);
or U12527 (N_12527,N_10873,N_10767);
nor U12528 (N_12528,N_11191,N_10235);
nor U12529 (N_12529,N_11327,N_11101);
nor U12530 (N_12530,N_10025,N_10664);
or U12531 (N_12531,N_11280,N_11380);
nand U12532 (N_12532,N_12402,N_11373);
or U12533 (N_12533,N_12315,N_10060);
nand U12534 (N_12534,N_11994,N_12067);
nor U12535 (N_12535,N_11933,N_12495);
and U12536 (N_12536,N_12486,N_12412);
and U12537 (N_12537,N_11821,N_12117);
and U12538 (N_12538,N_12440,N_10172);
nor U12539 (N_12539,N_11796,N_10359);
nand U12540 (N_12540,N_11113,N_12348);
nor U12541 (N_12541,N_10663,N_11362);
or U12542 (N_12542,N_11109,N_12467);
and U12543 (N_12543,N_10383,N_11354);
nand U12544 (N_12544,N_10166,N_10881);
or U12545 (N_12545,N_11455,N_11833);
and U12546 (N_12546,N_10207,N_10228);
and U12547 (N_12547,N_11937,N_12105);
nor U12548 (N_12548,N_11807,N_10675);
or U12549 (N_12549,N_11181,N_11454);
nand U12550 (N_12550,N_10922,N_10851);
nor U12551 (N_12551,N_10665,N_11147);
and U12552 (N_12552,N_11934,N_10119);
and U12553 (N_12553,N_11914,N_10582);
nor U12554 (N_12554,N_12497,N_10846);
and U12555 (N_12555,N_10290,N_12260);
nand U12556 (N_12556,N_10363,N_11621);
nand U12557 (N_12557,N_12265,N_12312);
nand U12558 (N_12558,N_10892,N_10611);
nor U12559 (N_12559,N_10474,N_10563);
nand U12560 (N_12560,N_12211,N_10432);
nand U12561 (N_12561,N_11315,N_11537);
and U12562 (N_12562,N_12430,N_11528);
and U12563 (N_12563,N_10101,N_11941);
nor U12564 (N_12564,N_10821,N_11577);
or U12565 (N_12565,N_11750,N_11457);
nand U12566 (N_12566,N_11339,N_12101);
xnor U12567 (N_12567,N_11017,N_10038);
nor U12568 (N_12568,N_10926,N_11224);
or U12569 (N_12569,N_11086,N_10764);
or U12570 (N_12570,N_10606,N_10061);
and U12571 (N_12571,N_11659,N_10492);
or U12572 (N_12572,N_11963,N_10883);
and U12573 (N_12573,N_10638,N_12295);
nand U12574 (N_12574,N_12383,N_11910);
nor U12575 (N_12575,N_10350,N_10173);
and U12576 (N_12576,N_10418,N_10260);
nand U12577 (N_12577,N_10800,N_12016);
or U12578 (N_12578,N_11095,N_11903);
and U12579 (N_12579,N_10730,N_11820);
nor U12580 (N_12580,N_12041,N_10882);
nand U12581 (N_12581,N_10157,N_12243);
or U12582 (N_12582,N_12465,N_11350);
or U12583 (N_12583,N_10862,N_10646);
or U12584 (N_12584,N_10915,N_10738);
or U12585 (N_12585,N_12446,N_12064);
nor U12586 (N_12586,N_11954,N_10278);
or U12587 (N_12587,N_10681,N_10340);
nand U12588 (N_12588,N_11895,N_12112);
and U12589 (N_12589,N_10558,N_12212);
or U12590 (N_12590,N_12036,N_11250);
or U12591 (N_12591,N_12287,N_10128);
or U12592 (N_12592,N_10106,N_11762);
or U12593 (N_12593,N_10921,N_10852);
nand U12594 (N_12594,N_10850,N_10238);
or U12595 (N_12595,N_11790,N_11310);
nand U12596 (N_12596,N_11429,N_11091);
nand U12597 (N_12597,N_12019,N_10812);
nor U12598 (N_12598,N_11203,N_10206);
and U12599 (N_12599,N_11948,N_11460);
nor U12600 (N_12600,N_10412,N_12086);
or U12601 (N_12601,N_12475,N_10975);
and U12602 (N_12602,N_11004,N_11335);
nand U12603 (N_12603,N_12106,N_10494);
and U12604 (N_12604,N_11111,N_10010);
and U12605 (N_12605,N_11502,N_10470);
nand U12606 (N_12606,N_11170,N_10572);
xor U12607 (N_12607,N_12460,N_10771);
nor U12608 (N_12608,N_11139,N_11013);
or U12609 (N_12609,N_12289,N_10395);
nand U12610 (N_12610,N_11296,N_10991);
nand U12611 (N_12611,N_12352,N_10605);
or U12612 (N_12612,N_10045,N_10911);
or U12613 (N_12613,N_11931,N_10810);
nor U12614 (N_12614,N_11506,N_10068);
nand U12615 (N_12615,N_12405,N_11898);
nand U12616 (N_12616,N_11396,N_11079);
or U12617 (N_12617,N_12489,N_10160);
and U12618 (N_12618,N_11241,N_10874);
and U12619 (N_12619,N_10177,N_11843);
or U12620 (N_12620,N_10818,N_11329);
nand U12621 (N_12621,N_11318,N_11791);
nor U12622 (N_12622,N_10592,N_11251);
and U12623 (N_12623,N_10216,N_10078);
and U12624 (N_12624,N_10808,N_10472);
nand U12625 (N_12625,N_12411,N_12194);
or U12626 (N_12626,N_12452,N_12135);
nand U12627 (N_12627,N_10398,N_11355);
nand U12628 (N_12628,N_12234,N_10224);
or U12629 (N_12629,N_11787,N_11152);
or U12630 (N_12630,N_12206,N_12363);
or U12631 (N_12631,N_10209,N_12132);
nand U12632 (N_12632,N_12425,N_12242);
and U12633 (N_12633,N_11048,N_10493);
or U12634 (N_12634,N_10924,N_10385);
nor U12635 (N_12635,N_10880,N_10967);
nand U12636 (N_12636,N_12169,N_10707);
or U12637 (N_12637,N_11923,N_10132);
and U12638 (N_12638,N_10074,N_11627);
and U12639 (N_12639,N_11240,N_11021);
nor U12640 (N_12640,N_12360,N_10763);
or U12641 (N_12641,N_11904,N_10030);
and U12642 (N_12642,N_11944,N_10628);
and U12643 (N_12643,N_10055,N_12025);
nor U12644 (N_12644,N_10896,N_12048);
nor U12645 (N_12645,N_11317,N_11379);
and U12646 (N_12646,N_12170,N_10002);
nor U12647 (N_12647,N_12291,N_11908);
nand U12648 (N_12648,N_10727,N_11563);
and U12649 (N_12649,N_10854,N_11749);
and U12650 (N_12650,N_11920,N_11440);
and U12651 (N_12651,N_12192,N_10033);
nor U12652 (N_12652,N_10781,N_11445);
nand U12653 (N_12653,N_10410,N_10249);
nor U12654 (N_12654,N_10276,N_12040);
or U12655 (N_12655,N_12244,N_11564);
nand U12656 (N_12656,N_12031,N_11729);
nand U12657 (N_12657,N_11603,N_11880);
nor U12658 (N_12658,N_10661,N_11047);
nand U12659 (N_12659,N_10263,N_11375);
or U12660 (N_12660,N_11515,N_10670);
nor U12661 (N_12661,N_10872,N_10169);
or U12662 (N_12662,N_11344,N_10136);
nand U12663 (N_12663,N_11299,N_11084);
or U12664 (N_12664,N_11995,N_12091);
and U12665 (N_12665,N_10639,N_12447);
and U12666 (N_12666,N_11847,N_10017);
nand U12667 (N_12667,N_11716,N_12078);
or U12668 (N_12668,N_10481,N_11166);
or U12669 (N_12669,N_10761,N_10579);
xor U12670 (N_12670,N_10886,N_10258);
and U12671 (N_12671,N_11651,N_10325);
and U12672 (N_12672,N_10236,N_10840);
or U12673 (N_12673,N_10012,N_11629);
and U12674 (N_12674,N_12252,N_10159);
or U12675 (N_12675,N_11149,N_11632);
or U12676 (N_12676,N_11658,N_10645);
or U12677 (N_12677,N_12274,N_11492);
nand U12678 (N_12678,N_11822,N_10411);
and U12679 (N_12679,N_12341,N_11523);
nor U12680 (N_12680,N_12056,N_11089);
nand U12681 (N_12681,N_11337,N_10015);
nor U12682 (N_12682,N_10845,N_12417);
nor U12683 (N_12683,N_12351,N_12026);
and U12684 (N_12684,N_12225,N_12410);
and U12685 (N_12685,N_10403,N_11067);
or U12686 (N_12686,N_11090,N_10754);
nor U12687 (N_12687,N_10425,N_12487);
nand U12688 (N_12688,N_10875,N_11728);
and U12689 (N_12689,N_11643,N_11487);
nand U12690 (N_12690,N_10460,N_10511);
or U12691 (N_12691,N_10163,N_10677);
nand U12692 (N_12692,N_11901,N_12218);
nand U12693 (N_12693,N_11692,N_11256);
and U12694 (N_12694,N_10589,N_10770);
or U12695 (N_12695,N_12346,N_10253);
and U12696 (N_12696,N_11174,N_10360);
and U12697 (N_12697,N_10778,N_11589);
nor U12698 (N_12698,N_12095,N_10051);
nand U12699 (N_12699,N_10552,N_11947);
nand U12700 (N_12700,N_12380,N_10586);
or U12701 (N_12701,N_11612,N_11190);
nand U12702 (N_12702,N_11075,N_11962);
nand U12703 (N_12703,N_11424,N_11129);
and U12704 (N_12704,N_10629,N_12071);
nor U12705 (N_12705,N_10441,N_11925);
nand U12706 (N_12706,N_10145,N_10614);
xor U12707 (N_12707,N_12272,N_11974);
and U12708 (N_12708,N_12496,N_12202);
and U12709 (N_12709,N_11894,N_11881);
nand U12710 (N_12710,N_10540,N_11185);
or U12711 (N_12711,N_10435,N_11292);
and U12712 (N_12712,N_10903,N_10690);
nand U12713 (N_12713,N_10528,N_10804);
nor U12714 (N_12714,N_10264,N_11080);
nand U12715 (N_12715,N_12266,N_10518);
or U12716 (N_12716,N_12069,N_10721);
and U12717 (N_12717,N_10052,N_11382);
nand U12718 (N_12718,N_10523,N_11939);
or U12719 (N_12719,N_10148,N_10534);
and U12720 (N_12720,N_10514,N_12092);
and U12721 (N_12721,N_11574,N_11193);
or U12722 (N_12722,N_11779,N_11970);
or U12723 (N_12723,N_12150,N_11630);
nand U12724 (N_12724,N_12152,N_10631);
or U12725 (N_12725,N_10233,N_12473);
or U12726 (N_12726,N_12462,N_12396);
nor U12727 (N_12727,N_12024,N_10442);
nor U12728 (N_12728,N_12392,N_11746);
or U12729 (N_12729,N_10925,N_12379);
and U12730 (N_12730,N_11110,N_10280);
nand U12731 (N_12731,N_10465,N_11488);
and U12732 (N_12732,N_12052,N_11102);
or U12733 (N_12733,N_11037,N_10698);
or U12734 (N_12734,N_11795,N_10019);
nand U12735 (N_12735,N_10246,N_12373);
or U12736 (N_12736,N_11419,N_12196);
and U12737 (N_12737,N_12314,N_10640);
nand U12738 (N_12738,N_12399,N_10667);
nand U12739 (N_12739,N_10554,N_11381);
nand U12740 (N_12740,N_11818,N_12388);
nor U12741 (N_12741,N_10368,N_10901);
nor U12742 (N_12742,N_10848,N_11215);
nor U12743 (N_12743,N_10088,N_11205);
nor U12744 (N_12744,N_10099,N_11919);
and U12745 (N_12745,N_12061,N_11398);
and U12746 (N_12746,N_11252,N_11176);
nand U12747 (N_12747,N_10682,N_10516);
and U12748 (N_12748,N_12131,N_11156);
and U12749 (N_12749,N_11525,N_11366);
and U12750 (N_12750,N_10498,N_10861);
and U12751 (N_12751,N_11592,N_11439);
nand U12752 (N_12752,N_11063,N_11049);
or U12753 (N_12753,N_11413,N_12469);
nand U12754 (N_12754,N_12357,N_12442);
nand U12755 (N_12755,N_11199,N_11167);
and U12756 (N_12756,N_12459,N_12426);
nand U12757 (N_12757,N_12200,N_10809);
or U12758 (N_12758,N_11300,N_11059);
nor U12759 (N_12759,N_12271,N_12386);
and U12760 (N_12760,N_10244,N_10351);
and U12761 (N_12761,N_10179,N_12207);
and U12762 (N_12762,N_10745,N_12264);
or U12763 (N_12763,N_10919,N_11119);
nor U12764 (N_12764,N_10488,N_11549);
or U12765 (N_12765,N_10584,N_10650);
or U12766 (N_12766,N_10195,N_10390);
nand U12767 (N_12767,N_10701,N_11596);
xor U12768 (N_12768,N_12393,N_11858);
nor U12769 (N_12769,N_10381,N_10227);
or U12770 (N_12770,N_11495,N_11340);
and U12771 (N_12771,N_11801,N_12156);
nor U12772 (N_12772,N_11260,N_10868);
or U12773 (N_12773,N_11108,N_11666);
and U12774 (N_12774,N_10413,N_11276);
nor U12775 (N_12775,N_12190,N_11093);
or U12776 (N_12776,N_12171,N_11529);
nor U12777 (N_12777,N_10815,N_11846);
or U12778 (N_12778,N_10034,N_10610);
nor U12779 (N_12779,N_11107,N_10737);
or U12780 (N_12780,N_12498,N_10344);
or U12781 (N_12781,N_11640,N_10705);
nor U12782 (N_12782,N_10741,N_11099);
nand U12783 (N_12783,N_11896,N_11493);
nor U12784 (N_12784,N_10277,N_12468);
nor U12785 (N_12785,N_12075,N_11283);
nor U12786 (N_12786,N_11733,N_11972);
nor U12787 (N_12787,N_10619,N_10097);
and U12788 (N_12788,N_10699,N_11432);
or U12789 (N_12789,N_12466,N_11784);
or U12790 (N_12790,N_10142,N_11872);
nor U12791 (N_12791,N_11561,N_11231);
nand U12792 (N_12792,N_11575,N_11799);
nor U12793 (N_12793,N_12356,N_10603);
and U12794 (N_12794,N_11540,N_12147);
nor U12795 (N_12795,N_10053,N_12185);
or U12796 (N_12796,N_10816,N_10288);
nor U12797 (N_12797,N_11652,N_10792);
nor U12798 (N_12798,N_12236,N_11352);
and U12799 (N_12799,N_10083,N_10086);
and U12800 (N_12800,N_11590,N_12209);
and U12801 (N_12801,N_11556,N_10312);
nor U12802 (N_12802,N_11247,N_11552);
or U12803 (N_12803,N_11501,N_11177);
or U12804 (N_12804,N_10303,N_10537);
nand U12805 (N_12805,N_12285,N_10805);
nand U12806 (N_12806,N_11142,N_10930);
or U12807 (N_12807,N_11553,N_12333);
and U12808 (N_12808,N_10555,N_10292);
nand U12809 (N_12809,N_10354,N_12324);
or U12810 (N_12810,N_12197,N_10170);
or U12811 (N_12811,N_11187,N_10152);
nand U12812 (N_12812,N_12414,N_11298);
and U12813 (N_12813,N_10267,N_11324);
and U12814 (N_12814,N_11731,N_10501);
nand U12815 (N_12815,N_11125,N_11538);
or U12816 (N_12816,N_11263,N_10377);
nor U12817 (N_12817,N_10668,N_10593);
or U12818 (N_12818,N_12336,N_11869);
xor U12819 (N_12819,N_11326,N_12240);
nand U12820 (N_12820,N_11245,N_10294);
nor U12821 (N_12821,N_10662,N_11226);
nand U12822 (N_12822,N_11124,N_10400);
nand U12823 (N_12823,N_10201,N_11158);
nor U12824 (N_12824,N_11971,N_10115);
or U12825 (N_12825,N_10433,N_10081);
or U12826 (N_12826,N_10073,N_11991);
and U12827 (N_12827,N_11855,N_10026);
or U12828 (N_12828,N_11464,N_10040);
nor U12829 (N_12829,N_11206,N_11076);
and U12830 (N_12830,N_11244,N_12002);
nand U12831 (N_12831,N_12110,N_10256);
nand U12832 (N_12832,N_11611,N_10210);
nand U12833 (N_12833,N_11507,N_11294);
xor U12834 (N_12834,N_10348,N_12251);
and U12835 (N_12835,N_11854,N_11421);
nor U12836 (N_12836,N_10291,N_10215);
nand U12837 (N_12837,N_10625,N_11544);
nor U12838 (N_12838,N_11988,N_11926);
or U12839 (N_12839,N_11953,N_10329);
nor U12840 (N_12840,N_10574,N_10255);
or U12841 (N_12841,N_10564,N_10069);
nor U12842 (N_12842,N_11491,N_12001);
or U12843 (N_12843,N_12104,N_10482);
nor U12844 (N_12844,N_12404,N_11718);
nand U12845 (N_12845,N_10849,N_10229);
nand U12846 (N_12846,N_11810,N_11647);
or U12847 (N_12847,N_11234,N_12406);
and U12848 (N_12848,N_11532,N_12088);
or U12849 (N_12849,N_10013,N_12005);
nand U12850 (N_12850,N_10916,N_11325);
nand U12851 (N_12851,N_10884,N_11351);
and U12852 (N_12852,N_11661,N_12491);
and U12853 (N_12853,N_11946,N_11936);
and U12854 (N_12854,N_10687,N_11547);
nand U12855 (N_12855,N_11850,N_10232);
xor U12856 (N_12856,N_10020,N_10304);
nand U12857 (N_12857,N_10118,N_11376);
nor U12858 (N_12858,N_11745,N_10343);
nand U12859 (N_12859,N_10143,N_11435);
or U12860 (N_12860,N_12176,N_11586);
or U12861 (N_12861,N_12142,N_12070);
nand U12862 (N_12862,N_10694,N_10895);
and U12863 (N_12863,N_11968,N_11684);
and U12864 (N_12864,N_11580,N_11703);
nor U12865 (N_12865,N_11571,N_11709);
nand U12866 (N_12866,N_11357,N_10612);
or U12867 (N_12867,N_12120,N_11437);
nand U12868 (N_12868,N_10752,N_10813);
or U12869 (N_12869,N_10478,N_10120);
and U12870 (N_12870,N_12318,N_11565);
nand U12871 (N_12871,N_11530,N_12046);
nand U12872 (N_12872,N_11816,N_12121);
or U12873 (N_12873,N_10655,N_10336);
nor U12874 (N_12874,N_10525,N_10462);
nand U12875 (N_12875,N_10702,N_12178);
and U12876 (N_12876,N_10134,N_11035);
nand U12877 (N_12877,N_10247,N_12445);
nor U12878 (N_12878,N_11415,N_10212);
and U12879 (N_12879,N_11906,N_11578);
or U12880 (N_12880,N_10957,N_10447);
nand U12881 (N_12881,N_11092,N_10176);
nand U12882 (N_12882,N_10155,N_11932);
or U12883 (N_12883,N_11469,N_10379);
nand U12884 (N_12884,N_10445,N_12258);
nand U12885 (N_12885,N_10185,N_10287);
and U12886 (N_12886,N_12384,N_10768);
nor U12887 (N_12887,N_12302,N_11978);
nand U12888 (N_12888,N_10955,N_11277);
or U12889 (N_12889,N_10674,N_10859);
nand U12890 (N_12890,N_11334,N_12327);
nand U12891 (N_12891,N_11653,N_11074);
or U12892 (N_12892,N_11907,N_11442);
and U12893 (N_12893,N_10855,N_11020);
nor U12894 (N_12894,N_11773,N_12480);
nor U12895 (N_12895,N_11572,N_12011);
nand U12896 (N_12896,N_11293,N_12073);
and U12897 (N_12897,N_11077,N_12372);
nor U12898 (N_12898,N_10414,N_10141);
nand U12899 (N_12899,N_11738,N_10806);
or U12900 (N_12900,N_10964,N_10984);
nand U12901 (N_12901,N_10347,N_11874);
nor U12902 (N_12902,N_10865,N_12173);
nor U12903 (N_12903,N_10717,N_10198);
and U12904 (N_12904,N_11751,N_10417);
and U12905 (N_12905,N_11761,N_11401);
or U12906 (N_12906,N_11559,N_11998);
and U12907 (N_12907,N_11056,N_10993);
nor U12908 (N_12908,N_11451,N_12248);
nor U12909 (N_12909,N_12035,N_11723);
and U12910 (N_12910,N_10685,N_10936);
nand U12911 (N_12911,N_12074,N_11527);
nor U12912 (N_12912,N_11747,N_12208);
or U12913 (N_12913,N_12353,N_11184);
or U12914 (N_12914,N_11007,N_11830);
or U12915 (N_12915,N_11051,N_11900);
nand U12916 (N_12916,N_11225,N_10602);
nand U12917 (N_12917,N_12102,N_11394);
and U12918 (N_12918,N_11585,N_12432);
or U12919 (N_12919,N_11774,N_10736);
nand U12920 (N_12920,N_10999,N_10434);
nor U12921 (N_12921,N_11985,N_11624);
nand U12922 (N_12922,N_11342,N_11393);
nand U12923 (N_12923,N_11160,N_12115);
and U12924 (N_12924,N_11060,N_12037);
nand U12925 (N_12925,N_12449,N_10509);
xor U12926 (N_12926,N_12081,N_11849);
nor U12927 (N_12927,N_11689,N_11212);
or U12928 (N_12928,N_10608,N_11441);
nand U12929 (N_12929,N_12317,N_10407);
and U12930 (N_12930,N_11369,N_10718);
nor U12931 (N_12931,N_11227,N_10457);
nand U12932 (N_12932,N_11798,N_11600);
and U12933 (N_12933,N_11182,N_10723);
nand U12934 (N_12934,N_11094,N_11752);
nand U12935 (N_12935,N_10811,N_10652);
and U12936 (N_12936,N_11311,N_10489);
or U12937 (N_12937,N_12345,N_11710);
or U12938 (N_12938,N_12470,N_10080);
or U12939 (N_12939,N_11246,N_10609);
nand U12940 (N_12940,N_11960,N_10647);
nor U12941 (N_12941,N_10302,N_11949);
or U12942 (N_12942,N_11669,N_10814);
and U12943 (N_12943,N_11172,N_11304);
nor U12944 (N_12944,N_10673,N_11786);
nor U12945 (N_12945,N_10150,N_11794);
and U12946 (N_12946,N_11253,N_11546);
and U12947 (N_12947,N_12155,N_10422);
nand U12948 (N_12948,N_10133,N_10144);
or U12949 (N_12949,N_11967,N_11628);
nor U12950 (N_12950,N_11186,N_11368);
nor U12951 (N_12951,N_11857,N_10456);
and U12952 (N_12952,N_10468,N_10765);
nor U12953 (N_12953,N_10949,N_12483);
or U12954 (N_12954,N_11599,N_11068);
or U12955 (N_12955,N_10683,N_10042);
and U12956 (N_12956,N_10372,N_10879);
nand U12957 (N_12957,N_10636,N_12136);
and U12958 (N_12958,N_10746,N_12205);
nand U12959 (N_12959,N_10194,N_12492);
nand U12960 (N_12960,N_11155,N_10987);
or U12961 (N_12961,N_11679,N_12422);
nand U12962 (N_12962,N_11959,N_10947);
nand U12963 (N_12963,N_10918,N_12490);
and U12964 (N_12964,N_11918,N_12476);
nor U12965 (N_12965,N_10654,N_11804);
nor U12966 (N_12966,N_11588,N_11498);
or U12967 (N_12967,N_11593,N_11775);
nand U12968 (N_12968,N_11028,N_12198);
and U12969 (N_12969,N_10419,N_11126);
nand U12970 (N_12970,N_10458,N_11922);
nor U12971 (N_12971,N_10421,N_10706);
nor U12972 (N_12972,N_12099,N_11913);
nor U12973 (N_12973,N_11386,N_11265);
and U12974 (N_12974,N_10823,N_11870);
nand U12975 (N_12975,N_10213,N_11204);
and U12976 (N_12976,N_10679,N_10766);
nor U12977 (N_12977,N_10842,N_10463);
nor U12978 (N_12978,N_10618,N_11496);
nor U12979 (N_12979,N_11064,N_11414);
and U12980 (N_12980,N_12481,N_10406);
and U12981 (N_12981,N_11510,N_10459);
or U12982 (N_12982,N_10500,N_10952);
nor U12983 (N_12983,N_10512,N_11213);
or U12984 (N_12984,N_12204,N_10440);
nor U12985 (N_12985,N_10945,N_12416);
nor U12986 (N_12986,N_11197,N_10904);
or U12987 (N_12987,N_12113,N_11598);
and U12988 (N_12988,N_12066,N_10063);
nand U12989 (N_12989,N_11130,N_10491);
and U12990 (N_12990,N_10082,N_11040);
or U12991 (N_12991,N_11837,N_10031);
or U12992 (N_12992,N_10098,N_10786);
and U12993 (N_12993,N_11404,N_10062);
nand U12994 (N_12994,N_11584,N_10322);
or U12995 (N_12995,N_12219,N_11178);
and U12996 (N_12996,N_11287,N_10835);
or U12997 (N_12997,N_10838,N_12122);
or U12998 (N_12998,N_10864,N_12096);
nand U12999 (N_12999,N_11838,N_10029);
or U13000 (N_13000,N_10275,N_10743);
or U13001 (N_13001,N_10230,N_11168);
nand U13002 (N_13002,N_11248,N_10977);
nand U13003 (N_13003,N_10268,N_11302);
nor U13004 (N_13004,N_10091,N_12288);
nand U13005 (N_13005,N_12221,N_10583);
and U13006 (N_13006,N_12164,N_10910);
nand U13007 (N_13007,N_12034,N_11144);
or U13008 (N_13008,N_11741,N_10378);
nor U13009 (N_13009,N_11452,N_11468);
nand U13010 (N_13010,N_11476,N_11148);
or U13011 (N_13011,N_11743,N_10265);
nor U13012 (N_13012,N_10963,N_10750);
or U13013 (N_13013,N_11238,N_10490);
and U13014 (N_13014,N_10054,N_10696);
or U13015 (N_13015,N_10121,N_12453);
or U13016 (N_13016,N_11470,N_11817);
and U13017 (N_13017,N_10154,N_11462);
nor U13018 (N_13018,N_10067,N_10757);
nand U13019 (N_13019,N_12390,N_11286);
and U13020 (N_13020,N_10797,N_11066);
nand U13021 (N_13021,N_12129,N_11873);
nor U13022 (N_13022,N_10357,N_10594);
nor U13023 (N_13023,N_12292,N_11388);
nor U13024 (N_13024,N_10416,N_10871);
or U13025 (N_13025,N_12323,N_11072);
or U13026 (N_13026,N_10789,N_10906);
nor U13027 (N_13027,N_11607,N_10587);
nor U13028 (N_13028,N_11509,N_11522);
nand U13029 (N_13029,N_10345,N_11730);
or U13030 (N_13030,N_11430,N_12397);
nand U13031 (N_13031,N_11882,N_10775);
nand U13032 (N_13032,N_11494,N_12456);
nor U13033 (N_13033,N_11453,N_10960);
nor U13034 (N_13034,N_10124,N_11322);
or U13035 (N_13035,N_11853,N_10917);
nor U13036 (N_13036,N_10355,N_12350);
nand U13037 (N_13037,N_10866,N_11997);
nor U13038 (N_13038,N_11217,N_10335);
nand U13039 (N_13039,N_11416,N_12213);
and U13040 (N_13040,N_10521,N_11301);
and U13041 (N_13041,N_12340,N_10342);
or U13042 (N_13042,N_10556,N_12220);
and U13043 (N_13043,N_11050,N_10373);
and U13044 (N_13044,N_10158,N_10744);
or U13045 (N_13045,N_11569,N_10467);
or U13046 (N_13046,N_11961,N_10932);
nor U13047 (N_13047,N_11306,N_12280);
nand U13048 (N_13048,N_11279,N_12343);
nor U13049 (N_13049,N_11361,N_10632);
nand U13050 (N_13050,N_10847,N_11417);
nand U13051 (N_13051,N_11521,N_10200);
nand U13052 (N_13052,N_10734,N_10935);
nor U13053 (N_13053,N_11765,N_10496);
and U13054 (N_13054,N_10680,N_11157);
and U13055 (N_13055,N_10095,N_11255);
nor U13056 (N_13056,N_10146,N_11977);
nor U13057 (N_13057,N_11374,N_11022);
nand U13058 (N_13058,N_10349,N_11018);
or U13059 (N_13059,N_10190,N_11132);
nor U13060 (N_13060,N_11668,N_11587);
or U13061 (N_13061,N_12233,N_10392);
nor U13062 (N_13062,N_11305,N_11636);
nand U13063 (N_13063,N_10486,N_12123);
nand U13064 (N_13064,N_12427,N_11019);
nand U13065 (N_13065,N_11045,N_11364);
and U13066 (N_13066,N_11842,N_11863);
and U13067 (N_13067,N_12421,N_11428);
and U13068 (N_13068,N_10751,N_10223);
or U13069 (N_13069,N_10666,N_11291);
and U13070 (N_13070,N_10001,N_10837);
nor U13071 (N_13071,N_10795,N_10382);
nand U13072 (N_13072,N_11281,N_10161);
or U13073 (N_13073,N_10505,N_12134);
nor U13074 (N_13074,N_12273,N_10131);
nand U13075 (N_13075,N_10566,N_10497);
or U13076 (N_13076,N_10762,N_11641);
or U13077 (N_13077,N_12349,N_10836);
nand U13078 (N_13078,N_10988,N_11519);
or U13079 (N_13079,N_12143,N_10365);
nand U13080 (N_13080,N_10990,N_12424);
or U13081 (N_13081,N_10044,N_11054);
or U13082 (N_13082,N_10968,N_10245);
or U13083 (N_13083,N_10827,N_12413);
and U13084 (N_13084,N_10909,N_10188);
nand U13085 (N_13085,N_11303,N_11637);
nor U13086 (N_13086,N_12013,N_10022);
nand U13087 (N_13087,N_10595,N_11688);
and U13088 (N_13088,N_11753,N_11087);
and U13089 (N_13089,N_11475,N_10164);
and U13090 (N_13090,N_11697,N_10484);
and U13091 (N_13091,N_10995,N_10139);
nand U13092 (N_13092,N_10424,N_10598);
or U13093 (N_13093,N_10064,N_11195);
nor U13094 (N_13094,N_10396,N_12371);
or U13095 (N_13095,N_10222,N_10621);
nor U13096 (N_13096,N_11812,N_11883);
nand U13097 (N_13097,N_11536,N_12189);
nand U13098 (N_13098,N_12133,N_11082);
and U13099 (N_13099,N_11824,N_10193);
or U13100 (N_13100,N_10832,N_12215);
and U13101 (N_13101,N_11924,N_10897);
nor U13102 (N_13102,N_12083,N_10076);
nand U13103 (N_13103,N_11105,N_10072);
or U13104 (N_13104,N_11793,N_11987);
and U13105 (N_13105,N_11031,N_12477);
and U13106 (N_13106,N_10105,N_11721);
or U13107 (N_13107,N_10626,N_10783);
nor U13108 (N_13108,N_11323,N_10408);
nand U13109 (N_13109,N_10807,N_11626);
nor U13110 (N_13110,N_10844,N_12418);
or U13111 (N_13111,N_11138,N_10234);
or U13112 (N_13112,N_10471,N_12347);
nor U13113 (N_13113,N_12439,N_12181);
nor U13114 (N_13114,N_10449,N_10642);
or U13115 (N_13115,N_12094,N_10079);
nor U13116 (N_13116,N_10671,N_10251);
and U13117 (N_13117,N_12151,N_11979);
and U13118 (N_13118,N_11268,N_11346);
nor U13119 (N_13119,N_11038,N_10798);
and U13120 (N_13120,N_11006,N_12305);
or U13121 (N_13121,N_11363,N_10996);
and U13122 (N_13122,N_10499,N_10863);
and U13123 (N_13123,N_12033,N_10483);
nand U13124 (N_13124,N_10109,N_11992);
nor U13125 (N_13125,N_10711,N_12389);
nor U13126 (N_13126,N_10300,N_10777);
or U13127 (N_13127,N_11555,N_10204);
or U13128 (N_13128,N_12114,N_11497);
nor U13129 (N_13129,N_12253,N_11980);
nand U13130 (N_13130,N_11755,N_11010);
and U13131 (N_13131,N_10826,N_11249);
nand U13132 (N_13132,N_11663,N_12245);
nand U13133 (N_13133,N_11313,N_11690);
nor U13134 (N_13134,N_12458,N_11272);
nand U13135 (N_13135,N_11594,N_11356);
or U13136 (N_13136,N_11909,N_11566);
or U13137 (N_13137,N_11614,N_11264);
nand U13138 (N_13138,N_11208,N_11826);
or U13139 (N_13139,N_12119,N_10959);
or U13140 (N_13140,N_11736,N_12051);
nand U13141 (N_13141,N_10000,N_11560);
nand U13142 (N_13142,N_11675,N_12325);
or U13143 (N_13143,N_11886,N_11449);
nor U13144 (N_13144,N_10970,N_11719);
nor U13145 (N_13145,N_11825,N_10782);
nor U13146 (N_13146,N_12039,N_10332);
or U13147 (N_13147,N_11805,N_12408);
nand U13148 (N_13148,N_11180,N_12282);
and U13149 (N_13149,N_12227,N_11030);
or U13150 (N_13150,N_11955,N_11695);
nand U13151 (N_13151,N_11678,N_10567);
and U13152 (N_13152,N_10125,N_10530);
and U13153 (N_13153,N_11143,N_11196);
nor U13154 (N_13154,N_11349,N_11484);
or U13155 (N_13155,N_10502,N_10732);
or U13156 (N_13156,N_12222,N_11073);
nor U13157 (N_13157,N_10093,N_10018);
nor U13158 (N_13158,N_12079,N_11889);
nand U13159 (N_13159,N_10542,N_11656);
or U13160 (N_13160,N_12298,N_11154);
nand U13161 (N_13161,N_11258,N_10049);
nand U13162 (N_13162,N_10905,N_11214);
or U13163 (N_13163,N_11671,N_11693);
nand U13164 (N_13164,N_11211,N_10376);
nor U13165 (N_13165,N_11085,N_10196);
nor U13166 (N_13166,N_10653,N_10182);
nor U13167 (N_13167,N_12398,N_10992);
or U13168 (N_13168,N_11290,N_12277);
nand U13169 (N_13169,N_10731,N_10041);
nand U13170 (N_13170,N_11975,N_10710);
xor U13171 (N_13171,N_10568,N_11771);
and U13172 (N_13172,N_10140,N_10257);
or U13173 (N_13173,N_10713,N_11179);
and U13174 (N_13174,N_11456,N_11616);
or U13175 (N_13175,N_11892,N_10785);
and U13176 (N_13176,N_10538,N_11389);
nor U13177 (N_13177,N_11032,N_12161);
nand U13178 (N_13178,N_10046,N_11969);
nand U13179 (N_13179,N_11732,N_10520);
or U13180 (N_13180,N_11687,N_10966);
nor U13181 (N_13181,N_10028,N_10600);
or U13182 (N_13182,N_10565,N_12090);
and U13183 (N_13183,N_11016,N_10221);
or U13184 (N_13184,N_12203,N_11921);
nor U13185 (N_13185,N_11707,N_12300);
and U13186 (N_13186,N_10973,N_12044);
nand U13187 (N_13187,N_11400,N_12140);
nand U13188 (N_13188,N_12058,N_11711);
nor U13189 (N_13189,N_10888,N_10108);
and U13190 (N_13190,N_11034,N_10065);
nand U13191 (N_13191,N_12281,N_11288);
or U13192 (N_13192,N_12157,N_10824);
nand U13193 (N_13193,N_10087,N_11489);
and U13194 (N_13194,N_12030,N_11405);
or U13195 (N_13195,N_10858,N_11864);
and U13196 (N_13196,N_10285,N_11467);
nand U13197 (N_13197,N_12269,N_11778);
nor U13198 (N_13198,N_10452,N_11024);
nand U13199 (N_13199,N_11121,N_10519);
nor U13200 (N_13200,N_10830,N_11043);
nand U13201 (N_13201,N_11320,N_10508);
and U13202 (N_13202,N_11966,N_10371);
and U13203 (N_13203,N_10299,N_12177);
nor U13204 (N_13204,N_11543,N_12223);
and U13205 (N_13205,N_11216,N_10283);
and U13206 (N_13206,N_10444,N_12391);
or U13207 (N_13207,N_11070,N_12362);
and U13208 (N_13208,N_11957,N_10700);
xnor U13209 (N_13209,N_12354,N_10709);
nor U13210 (N_13210,N_11159,N_12448);
or U13211 (N_13211,N_12464,N_11811);
or U13212 (N_13212,N_11912,N_11674);
nand U13213 (N_13213,N_12344,N_10423);
nor U13214 (N_13214,N_11295,N_11759);
or U13215 (N_13215,N_10024,N_10703);
or U13216 (N_13216,N_10479,N_10420);
nor U13217 (N_13217,N_12216,N_10330);
and U13218 (N_13218,N_11232,N_12008);
and U13219 (N_13219,N_10735,N_11631);
nor U13220 (N_13220,N_10834,N_10448);
nand U13221 (N_13221,N_10570,N_11237);
nand U13222 (N_13222,N_11735,N_10107);
nand U13223 (N_13223,N_12250,N_12268);
and U13224 (N_13224,N_12438,N_10760);
and U13225 (N_13225,N_11742,N_10931);
or U13226 (N_13226,N_11989,N_10780);
and U13227 (N_13227,N_11878,N_12313);
nor U13228 (N_13228,N_12010,N_12231);
nor U13229 (N_13229,N_12254,N_10541);
and U13230 (N_13230,N_12457,N_11657);
nor U13231 (N_13231,N_10953,N_12055);
nand U13232 (N_13232,N_10323,N_11789);
nor U13233 (N_13233,N_10279,N_12478);
nand U13234 (N_13234,N_12097,N_11649);
nor U13235 (N_13235,N_10337,N_10352);
nor U13236 (N_13236,N_10720,N_10651);
nand U13237 (N_13237,N_11840,N_12138);
and U13238 (N_13238,N_11567,N_10096);
nand U13239 (N_13239,N_10370,N_12415);
or U13240 (N_13240,N_10929,N_11754);
xor U13241 (N_13241,N_10747,N_10191);
nand U13242 (N_13242,N_10704,N_10615);
nor U13243 (N_13243,N_11229,N_10793);
nor U13244 (N_13244,N_11052,N_10090);
nor U13245 (N_13245,N_11672,N_10867);
or U13246 (N_13246,N_10515,N_10311);
nand U13247 (N_13247,N_10982,N_10887);
nand U13248 (N_13248,N_10333,N_12235);
or U13249 (N_13249,N_10167,N_12382);
or U13250 (N_13250,N_10480,N_10553);
nor U13251 (N_13251,N_10367,N_12293);
or U13252 (N_13252,N_10016,N_10270);
nor U13253 (N_13253,N_11542,N_10998);
nor U13254 (N_13254,N_11145,N_10114);
nor U13255 (N_13255,N_10199,N_10241);
and U13256 (N_13256,N_12331,N_11336);
nor U13257 (N_13257,N_11461,N_10712);
nand U13258 (N_13258,N_11055,N_10617);
or U13259 (N_13259,N_10237,N_11866);
and U13260 (N_13260,N_10733,N_10779);
or U13261 (N_13261,N_12299,N_10550);
nor U13262 (N_13262,N_10314,N_10790);
nor U13263 (N_13263,N_12179,N_11545);
or U13264 (N_13264,N_11372,N_11450);
nor U13265 (N_13265,N_10117,N_10728);
nand U13266 (N_13266,N_11383,N_12241);
and U13267 (N_13267,N_10772,N_10856);
and U13268 (N_13268,N_12111,N_10788);
nand U13269 (N_13269,N_11411,N_11667);
nand U13270 (N_13270,N_11887,N_11734);
and U13271 (N_13271,N_12259,N_11230);
or U13272 (N_13272,N_12419,N_10532);
nor U13273 (N_13273,N_11444,N_11477);
or U13274 (N_13274,N_11482,N_12077);
nor U13275 (N_13275,N_10689,N_11333);
nor U13276 (N_13276,N_10506,N_11783);
or U13277 (N_13277,N_10175,N_11312);
or U13278 (N_13278,N_12159,N_10684);
or U13279 (N_13279,N_12308,N_11984);
nand U13280 (N_13280,N_10362,N_11151);
nand U13281 (N_13281,N_10171,N_11557);
or U13282 (N_13282,N_11860,N_10749);
and U13283 (N_13283,N_10755,N_10817);
or U13284 (N_13284,N_11005,N_10974);
nand U13285 (N_13285,N_10591,N_12355);
nor U13286 (N_13286,N_11254,N_10401);
or U13287 (N_13287,N_11427,N_11410);
nor U13288 (N_13288,N_10688,N_11797);
nand U13289 (N_13289,N_11257,N_10889);
nor U13290 (N_13290,N_11696,N_11478);
nor U13291 (N_13291,N_11128,N_12038);
and U13292 (N_13292,N_11504,N_10252);
nand U13293 (N_13293,N_12158,N_10575);
nor U13294 (N_13294,N_11262,N_12141);
or U13295 (N_13295,N_12021,N_11026);
or U13296 (N_13296,N_12023,N_10739);
nor U13297 (N_13297,N_11014,N_12482);
nor U13298 (N_13298,N_11459,N_10487);
nand U13299 (N_13299,N_12316,N_10476);
or U13300 (N_13300,N_10364,N_10820);
or U13301 (N_13301,N_12276,N_11958);
nand U13302 (N_13302,N_12076,N_12004);
or U13303 (N_13303,N_10588,N_11235);
or U13304 (N_13304,N_11137,N_11813);
nor U13305 (N_13305,N_12082,N_12029);
and U13306 (N_13306,N_10934,N_12322);
and U13307 (N_13307,N_11513,N_11233);
nor U13308 (N_13308,N_10526,N_11802);
nor U13309 (N_13309,N_10321,N_12116);
nor U13310 (N_13310,N_10389,N_10784);
nor U13311 (N_13311,N_10569,N_11986);
or U13312 (N_13312,N_11646,N_10043);
nand U13313 (N_13313,N_10439,N_10983);
nor U13314 (N_13314,N_12165,N_12230);
or U13315 (N_13315,N_10356,N_11387);
and U13316 (N_13316,N_10309,N_11447);
or U13317 (N_13317,N_10898,N_10269);
nand U13318 (N_13318,N_12130,N_11029);
and U13319 (N_13319,N_12499,N_10104);
or U13320 (N_13320,N_10697,N_11164);
nand U13321 (N_13321,N_12407,N_11620);
and U13322 (N_13322,N_10281,N_12270);
nand U13323 (N_13323,N_11071,N_10129);
or U13324 (N_13324,N_11608,N_10008);
nand U13325 (N_13325,N_11514,N_11472);
nand U13326 (N_13326,N_11644,N_11814);
nor U13327 (N_13327,N_11141,N_11950);
or U13328 (N_13328,N_10219,N_11655);
nor U13329 (N_13329,N_10011,N_11473);
nor U13330 (N_13330,N_11665,N_11391);
nor U13331 (N_13331,N_11065,N_12228);
nand U13332 (N_13332,N_11884,N_10271);
and U13333 (N_13333,N_10248,N_10084);
or U13334 (N_13334,N_11479,N_12145);
nand U13335 (N_13335,N_10409,N_12366);
and U13336 (N_13336,N_11061,N_12068);
and U13337 (N_13337,N_10986,N_11331);
and U13338 (N_13338,N_11964,N_10429);
or U13339 (N_13339,N_11505,N_10184);
nor U13340 (N_13340,N_10218,N_10923);
and U13341 (N_13341,N_11650,N_10686);
and U13342 (N_13342,N_10920,N_11377);
and U13343 (N_13343,N_12434,N_11171);
or U13344 (N_13344,N_11384,N_10669);
or U13345 (N_13345,N_11766,N_10450);
or U13346 (N_13346,N_11831,N_10828);
nand U13347 (N_13347,N_10841,N_11106);
nand U13348 (N_13348,N_11201,N_11591);
nor U13349 (N_13349,N_11638,N_12153);
nor U13350 (N_13350,N_12182,N_11083);
or U13351 (N_13351,N_11219,N_10576);
nand U13352 (N_13352,N_10071,N_11426);
and U13353 (N_13353,N_10796,N_10633);
nor U13354 (N_13354,N_11876,N_11782);
and U13355 (N_13355,N_10604,N_11041);
and U13356 (N_13356,N_10869,N_11271);
or U13357 (N_13357,N_11981,N_12367);
nand U13358 (N_13358,N_11033,N_11436);
and U13359 (N_13359,N_11691,N_11942);
nor U13360 (N_13360,N_12054,N_12429);
nand U13361 (N_13361,N_11717,N_10539);
and U13362 (N_13362,N_11161,N_12232);
and U13363 (N_13363,N_11897,N_10259);
and U13364 (N_13364,N_12149,N_11929);
nor U13365 (N_13365,N_12275,N_11792);
nand U13366 (N_13366,N_11408,N_12377);
nor U13367 (N_13367,N_12217,N_10843);
and U13368 (N_13368,N_11027,N_12378);
and U13369 (N_13369,N_10165,N_10137);
nand U13370 (N_13370,N_10438,N_10578);
and U13371 (N_13371,N_10980,N_11785);
and U13372 (N_13372,N_10014,N_11117);
and U13373 (N_13373,N_12256,N_10386);
or U13374 (N_13374,N_11088,N_11943);
nand U13375 (N_13375,N_10913,N_11316);
and U13376 (N_13376,N_11945,N_11518);
or U13377 (N_13377,N_11698,N_11409);
or U13378 (N_13378,N_10994,N_12278);
nor U13379 (N_13379,N_11823,N_10004);
or U13380 (N_13380,N_11744,N_11524);
and U13381 (N_13381,N_10135,N_10944);
nand U13382 (N_13382,N_12000,N_10529);
or U13383 (N_13383,N_10361,N_11371);
and U13384 (N_13384,N_10313,N_10577);
and U13385 (N_13385,N_11579,N_10822);
xnor U13386 (N_13386,N_10860,N_11173);
or U13387 (N_13387,N_11044,N_11535);
nand U13388 (N_13388,N_11202,N_10958);
nor U13389 (N_13389,N_10585,N_10168);
nand U13390 (N_13390,N_11701,N_11617);
and U13391 (N_13391,N_10791,N_11261);
nand U13392 (N_13392,N_11713,N_12284);
or U13393 (N_13393,N_11000,N_10358);
or U13394 (N_13394,N_12290,N_12463);
or U13395 (N_13395,N_11239,N_10599);
nor U13396 (N_13396,N_10597,N_10485);
nand U13397 (N_13397,N_10469,N_12065);
or U13398 (N_13398,N_10641,N_11856);
and U13399 (N_13399,N_12326,N_12267);
or U13400 (N_13400,N_10056,N_10243);
nor U13401 (N_13401,N_11118,N_10544);
nor U13402 (N_13402,N_12339,N_11917);
nor U13403 (N_13403,N_12226,N_10938);
or U13404 (N_13404,N_12261,N_10985);
nand U13405 (N_13405,N_11554,N_11466);
nor U13406 (N_13406,N_11639,N_11757);
or U13407 (N_13407,N_11756,N_12249);
nand U13408 (N_13408,N_10503,N_12214);
nand U13409 (N_13409,N_10774,N_10058);
and U13410 (N_13410,N_10802,N_10978);
nand U13411 (N_13411,N_10231,N_11122);
or U13412 (N_13412,N_11677,N_12229);
and U13413 (N_13413,N_10630,N_12160);
and U13414 (N_13414,N_11726,N_10643);
and U13415 (N_13415,N_10310,N_10388);
nand U13416 (N_13416,N_10316,N_11581);
and U13417 (N_13417,N_11915,N_11618);
nand U13418 (N_13418,N_12087,N_10187);
nor U13419 (N_13419,N_11699,N_12125);
xnor U13420 (N_13420,N_10543,N_12423);
nand U13421 (N_13421,N_11576,N_12124);
or U13422 (N_13422,N_10426,N_11123);
nand U13423 (N_13423,N_10927,N_10306);
and U13424 (N_13424,N_12435,N_11550);
nor U13425 (N_13425,N_11332,N_10581);
and U13426 (N_13426,N_10138,N_12246);
and U13427 (N_13427,N_10627,N_10716);
nor U13428 (N_13428,N_11976,N_10773);
or U13429 (N_13429,N_12304,N_10548);
nor U13430 (N_13430,N_12328,N_12337);
nand U13431 (N_13431,N_11407,N_11633);
and U13432 (N_13432,N_10205,N_10110);
nand U13433 (N_13433,N_10353,N_11769);
and U13434 (N_13434,N_10876,N_11402);
nand U13435 (N_13435,N_10339,N_10513);
and U13436 (N_13436,N_11446,N_10549);
nand U13437 (N_13437,N_11645,N_12338);
nor U13438 (N_13438,N_11474,N_12062);
nor U13439 (N_13439,N_10436,N_11764);
nor U13440 (N_13440,N_11911,N_10658);
nor U13441 (N_13441,N_11228,N_11069);
nand U13442 (N_13442,N_12428,N_12370);
nand U13443 (N_13443,N_10111,N_11194);
nand U13444 (N_13444,N_11508,N_11002);
nand U13445 (N_13445,N_11861,N_10437);
nor U13446 (N_13446,N_10384,N_11116);
nand U13447 (N_13447,N_10753,N_11714);
nor U13448 (N_13448,N_11480,N_11865);
nand U13449 (N_13449,N_10261,N_12263);
or U13450 (N_13450,N_12224,N_10853);
nor U13451 (N_13451,N_12247,N_10186);
and U13452 (N_13452,N_11192,N_11573);
nor U13453 (N_13453,N_11702,N_11036);
and U13454 (N_13454,N_12400,N_11890);
and U13455 (N_13455,N_11605,N_11112);
nand U13456 (N_13456,N_11685,N_10695);
or U13457 (N_13457,N_11788,N_12049);
xor U13458 (N_13458,N_10391,N_10634);
nand U13459 (N_13459,N_10103,N_12193);
and U13460 (N_13460,N_11358,N_10893);
nand U13461 (N_13461,N_11406,N_10242);
nor U13462 (N_13462,N_12126,N_10130);
nor U13463 (N_13463,N_11443,N_10151);
nand U13464 (N_13464,N_11725,N_11438);
or U13465 (N_13465,N_10305,N_10559);
nand U13466 (N_13466,N_10622,N_11058);
nand U13467 (N_13467,N_11708,N_10477);
nor U13468 (N_13468,N_12401,N_11808);
or U13469 (N_13469,N_11965,N_10127);
or U13470 (N_13470,N_10580,N_11673);
nor U13471 (N_13471,N_12493,N_11819);
and U13472 (N_13472,N_11526,N_11583);
nand U13473 (N_13473,N_12375,N_11500);
nand U13474 (N_13474,N_10510,N_11623);
nand U13475 (N_13475,N_10907,N_10147);
nor U13476 (N_13476,N_11270,N_11015);
nor U13477 (N_13477,N_10308,N_10250);
and U13478 (N_13478,N_10116,N_12403);
or U13479 (N_13479,N_12433,N_11531);
and U13480 (N_13480,N_11284,N_11223);
nand U13481 (N_13481,N_10007,N_11120);
or U13482 (N_13482,N_11930,N_12342);
nand U13483 (N_13483,N_11720,N_11664);
and U13484 (N_13484,N_11803,N_11654);
or U13485 (N_13485,N_10660,N_10203);
nor U13486 (N_13486,N_10284,N_11499);
nand U13487 (N_13487,N_12127,N_11285);
and U13488 (N_13488,N_11648,N_10535);
or U13489 (N_13489,N_10740,N_10551);
nor U13490 (N_13490,N_11236,N_10338);
nand U13491 (N_13491,N_10415,N_10524);
and U13492 (N_13492,N_12239,N_10404);
nor U13493 (N_13493,N_10939,N_11360);
nor U13494 (N_13494,N_11613,N_11431);
and U13495 (N_13495,N_10573,N_12320);
nand U13496 (N_13496,N_10950,N_11935);
and U13497 (N_13497,N_12047,N_10431);
nand U13498 (N_13498,N_12461,N_10274);
nand U13499 (N_13499,N_11815,N_10961);
nand U13500 (N_13500,N_11727,N_10341);
nor U13501 (N_13501,N_11634,N_11057);
or U13502 (N_13502,N_10693,N_10003);
nand U13503 (N_13503,N_11338,N_10942);
nand U13504 (N_13504,N_10113,N_10546);
and U13505 (N_13505,N_11737,N_11996);
nand U13506 (N_13506,N_12450,N_11023);
and U13507 (N_13507,N_10298,N_12162);
nand U13508 (N_13508,N_11982,N_10036);
nor U13509 (N_13509,N_12394,N_11562);
and U13510 (N_13510,N_12437,N_11539);
nor U13511 (N_13511,N_12319,N_10273);
or U13512 (N_13512,N_12009,N_10620);
nor U13513 (N_13513,N_11307,N_12455);
nand U13514 (N_13514,N_11458,N_11222);
and U13515 (N_13515,N_11341,N_12172);
nand U13516 (N_13516,N_10180,N_12080);
nor U13517 (N_13517,N_11845,N_10644);
nor U13518 (N_13518,N_11127,N_10531);
nor U13519 (N_13519,N_10678,N_11952);
nor U13520 (N_13520,N_11169,N_10517);
or U13521 (N_13521,N_10149,N_11131);
and U13522 (N_13522,N_10297,N_10315);
and U13523 (N_13523,N_11520,N_11282);
nor U13524 (N_13524,N_11039,N_11893);
or U13525 (N_13525,N_11534,N_11486);
or U13526 (N_13526,N_10894,N_10153);
nand U13527 (N_13527,N_11150,N_10857);
nor U13528 (N_13528,N_12168,N_12297);
nand U13529 (N_13529,N_11308,N_10399);
or U13530 (N_13530,N_11175,N_12012);
nand U13531 (N_13531,N_10758,N_10870);
nor U13532 (N_13532,N_10226,N_12210);
nor U13533 (N_13533,N_11888,N_11042);
or U13534 (N_13534,N_12184,N_10616);
or U13535 (N_13535,N_11809,N_10307);
nand U13536 (N_13536,N_10374,N_10676);
nand U13537 (N_13537,N_10296,N_10211);
or U13538 (N_13538,N_10799,N_11739);
nor U13539 (N_13539,N_10039,N_12365);
nand U13540 (N_13540,N_12310,N_11533);
xnor U13541 (N_13541,N_10005,N_11483);
or U13542 (N_13542,N_11776,N_12027);
nand U13543 (N_13543,N_11905,N_10192);
or U13544 (N_13544,N_11162,N_11700);
and U13545 (N_13545,N_11604,N_12154);
nand U13546 (N_13546,N_12146,N_10181);
xor U13547 (N_13547,N_12306,N_10748);
nor U13548 (N_13548,N_10969,N_11153);
nor U13549 (N_13549,N_11448,N_10397);
and U13550 (N_13550,N_12166,N_11780);
nand U13551 (N_13551,N_10443,N_12103);
or U13552 (N_13552,N_11715,N_11243);
or U13553 (N_13553,N_10262,N_10220);
nand U13554 (N_13554,N_12238,N_12286);
and U13555 (N_13555,N_10466,N_11642);
nand U13556 (N_13556,N_10545,N_10366);
and U13557 (N_13557,N_11397,N_12100);
and U13558 (N_13558,N_11763,N_11218);
or U13559 (N_13559,N_11834,N_11582);
or U13560 (N_13560,N_12072,N_11378);
nand U13561 (N_13561,N_10504,N_10943);
nand U13562 (N_13562,N_11670,N_11683);
nor U13563 (N_13563,N_10979,N_10596);
nor U13564 (N_13564,N_10446,N_11289);
nor U13565 (N_13565,N_11423,N_10324);
nor U13566 (N_13566,N_11481,N_11365);
nor U13567 (N_13567,N_10972,N_11829);
nor U13568 (N_13568,N_12139,N_11274);
or U13569 (N_13569,N_12369,N_10899);
nand U13570 (N_13570,N_11003,N_11601);
nand U13571 (N_13571,N_10048,N_11420);
and U13572 (N_13572,N_11770,N_10208);
and U13573 (N_13573,N_11848,N_11740);
nand U13574 (N_13574,N_11053,N_12334);
and U13575 (N_13575,N_10971,N_11135);
and U13576 (N_13576,N_12108,N_11852);
nand U13577 (N_13577,N_10561,N_11973);
and U13578 (N_13578,N_11956,N_11682);
nand U13579 (N_13579,N_10346,N_10326);
nor U13580 (N_13580,N_10059,N_11859);
nand U13581 (N_13581,N_12032,N_11851);
or U13582 (N_13582,N_12484,N_10393);
xor U13583 (N_13583,N_10427,N_12381);
nand U13584 (N_13584,N_12007,N_12436);
or U13585 (N_13585,N_10089,N_10183);
or U13586 (N_13586,N_12186,N_10454);
nor U13587 (N_13587,N_10989,N_10473);
and U13588 (N_13588,N_10877,N_11485);
and U13589 (N_13589,N_11828,N_11597);
and U13590 (N_13590,N_12303,N_10461);
nor U13591 (N_13591,N_11146,N_12180);
and U13592 (N_13592,N_11418,N_12084);
nand U13593 (N_13593,N_12309,N_10331);
and U13594 (N_13594,N_12053,N_10320);
and U13595 (N_13595,N_10112,N_12059);
nor U13596 (N_13596,N_10715,N_10319);
nand U13597 (N_13597,N_10607,N_12311);
and U13598 (N_13598,N_12014,N_10794);
nand U13599 (N_13599,N_11412,N_11347);
nor U13600 (N_13600,N_12109,N_10197);
and U13601 (N_13601,N_11676,N_10908);
and U13602 (N_13602,N_12485,N_12089);
nand U13603 (N_13603,N_11999,N_10571);
nor U13604 (N_13604,N_12301,N_11343);
or U13605 (N_13605,N_12199,N_10430);
nand U13606 (N_13606,N_11348,N_11844);
nand U13607 (N_13607,N_10122,N_10266);
or U13608 (N_13608,N_12335,N_10956);
and U13609 (N_13609,N_12085,N_12494);
and U13610 (N_13610,N_12174,N_10729);
nand U13611 (N_13611,N_10289,N_12020);
or U13612 (N_13612,N_11704,N_10672);
nand U13613 (N_13613,N_11951,N_10659);
and U13614 (N_13614,N_11609,N_10405);
and U13615 (N_13615,N_12431,N_11983);
nand U13616 (N_13616,N_11885,N_12329);
or U13617 (N_13617,N_11114,N_11927);
nor U13618 (N_13618,N_12479,N_11207);
nor U13619 (N_13619,N_10891,N_11189);
and U13620 (N_13620,N_12454,N_10507);
nor U13621 (N_13621,N_10648,N_11722);
nor U13622 (N_13622,N_11622,N_10557);
nand U13623 (N_13623,N_11097,N_12257);
and U13624 (N_13624,N_12374,N_11748);
or U13625 (N_13625,N_11841,N_10387);
or U13626 (N_13626,N_10102,N_12279);
or U13627 (N_13627,N_10601,N_10070);
xnor U13628 (N_13628,N_10037,N_12488);
nor U13629 (N_13629,N_12443,N_10085);
nor U13630 (N_13630,N_10724,N_11871);
nand U13631 (N_13631,N_12191,N_12128);
and U13632 (N_13632,N_12296,N_11463);
nand U13633 (N_13633,N_11862,N_10174);
nor U13634 (N_13634,N_10066,N_12060);
nor U13635 (N_13635,N_11096,N_12332);
nor U13636 (N_13636,N_11705,N_11104);
nor U13637 (N_13637,N_12175,N_11938);
nand U13638 (N_13638,N_12017,N_10217);
nor U13639 (N_13639,N_10536,N_12255);
nor U13640 (N_13640,N_12321,N_11098);
or U13641 (N_13641,N_11390,N_12006);
xor U13642 (N_13642,N_10885,N_10948);
and U13643 (N_13643,N_11465,N_10692);
or U13644 (N_13644,N_10455,N_11133);
or U13645 (N_13645,N_10725,N_11615);
and U13646 (N_13646,N_11011,N_11009);
nand U13647 (N_13647,N_11662,N_12045);
and U13648 (N_13648,N_11273,N_10756);
nand U13649 (N_13649,N_11879,N_10759);
and U13650 (N_13650,N_10318,N_10094);
nand U13651 (N_13651,N_10522,N_11993);
nor U13652 (N_13652,N_11570,N_11220);
or U13653 (N_13653,N_11610,N_11395);
nor U13654 (N_13654,N_10464,N_10965);
nor U13655 (N_13655,N_11940,N_11760);
nor U13656 (N_13656,N_11359,N_10050);
and U13657 (N_13657,N_11163,N_11899);
nand U13658 (N_13658,N_11242,N_11183);
nor U13659 (N_13659,N_11602,N_11025);
or U13660 (N_13660,N_12015,N_11471);
nand U13661 (N_13661,N_11517,N_11314);
or U13662 (N_13662,N_11012,N_11209);
nor U13663 (N_13663,N_12359,N_12409);
or U13664 (N_13664,N_10328,N_10962);
or U13665 (N_13665,N_11827,N_10451);
nand U13666 (N_13666,N_10928,N_10100);
nor U13667 (N_13667,N_12195,N_10776);
or U13668 (N_13668,N_11319,N_11259);
or U13669 (N_13669,N_11328,N_10282);
or U13670 (N_13670,N_11275,N_10047);
nand U13671 (N_13671,N_11200,N_11800);
or U13672 (N_13672,N_10254,N_11619);
nor U13673 (N_13673,N_11541,N_11877);
nor U13674 (N_13674,N_10719,N_12187);
and U13675 (N_13675,N_12107,N_10156);
nand U13676 (N_13676,N_10742,N_11832);
and U13677 (N_13677,N_12307,N_10997);
nand U13678 (N_13678,N_12361,N_12188);
and U13679 (N_13679,N_10035,N_10286);
or U13680 (N_13680,N_11839,N_10831);
nand U13681 (N_13681,N_11768,N_11134);
nand U13682 (N_13682,N_11558,N_12022);
or U13683 (N_13683,N_12043,N_11635);
and U13684 (N_13684,N_11140,N_10317);
or U13685 (N_13685,N_12163,N_10590);
nor U13686 (N_13686,N_11503,N_11568);
and U13687 (N_13687,N_11902,N_10941);
and U13688 (N_13688,N_12028,N_12294);
nand U13689 (N_13689,N_11928,N_10272);
or U13690 (N_13690,N_12376,N_10951);
nand U13691 (N_13691,N_11706,N_11758);
nor U13692 (N_13692,N_11916,N_12364);
nor U13693 (N_13693,N_10375,N_11891);
or U13694 (N_13694,N_11046,N_12387);
nand U13695 (N_13695,N_10819,N_11321);
nand U13696 (N_13696,N_10940,N_11516);
nor U13697 (N_13697,N_11115,N_10657);
or U13698 (N_13698,N_10162,N_11867);
nand U13699 (N_13699,N_11686,N_12148);
and U13700 (N_13700,N_10009,N_11836);
nor U13701 (N_13701,N_12018,N_11781);
nor U13702 (N_13702,N_10295,N_11221);
or U13703 (N_13703,N_10077,N_11269);
nor U13704 (N_13704,N_12098,N_11370);
or U13705 (N_13705,N_11345,N_10293);
and U13706 (N_13706,N_11392,N_11062);
and U13707 (N_13707,N_12093,N_12471);
nand U13708 (N_13708,N_11278,N_12201);
or U13709 (N_13709,N_10021,N_10027);
nor U13710 (N_13710,N_10801,N_10202);
or U13711 (N_13711,N_10092,N_10946);
nor U13712 (N_13712,N_10075,N_11001);
nand U13713 (N_13713,N_12441,N_10914);
nand U13714 (N_13714,N_11990,N_10803);
and U13715 (N_13715,N_10624,N_11595);
xor U13716 (N_13716,N_12063,N_10334);
and U13717 (N_13717,N_10178,N_10635);
nor U13718 (N_13718,N_10123,N_12144);
nand U13719 (N_13719,N_11490,N_11875);
nor U13720 (N_13720,N_11548,N_10023);
or U13721 (N_13721,N_11081,N_11210);
and U13722 (N_13722,N_12395,N_12330);
nand U13723 (N_13723,N_10327,N_11681);
or U13724 (N_13724,N_10890,N_10708);
or U13725 (N_13725,N_10637,N_10787);
nor U13726 (N_13726,N_10933,N_11625);
or U13727 (N_13727,N_11136,N_10726);
nor U13728 (N_13728,N_11694,N_12057);
and U13729 (N_13729,N_11353,N_10691);
or U13730 (N_13730,N_12183,N_11385);
or U13731 (N_13731,N_11806,N_10829);
and U13732 (N_13732,N_10623,N_10613);
and U13733 (N_13733,N_11724,N_11188);
and U13734 (N_13734,N_10722,N_10937);
nor U13735 (N_13735,N_11330,N_10301);
nor U13736 (N_13736,N_11309,N_10126);
and U13737 (N_13737,N_10649,N_12368);
and U13738 (N_13738,N_12003,N_11266);
nor U13739 (N_13739,N_10189,N_10240);
nor U13740 (N_13740,N_12385,N_10533);
and U13741 (N_13741,N_11198,N_10912);
nand U13742 (N_13742,N_11422,N_10714);
nand U13743 (N_13743,N_11868,N_11434);
and U13744 (N_13744,N_12042,N_11712);
nor U13745 (N_13745,N_10394,N_11835);
and U13746 (N_13746,N_11551,N_11512);
or U13747 (N_13747,N_10547,N_10527);
nor U13748 (N_13748,N_11767,N_12050);
nand U13749 (N_13749,N_12358,N_11103);
and U13750 (N_13750,N_10066,N_11492);
nor U13751 (N_13751,N_10788,N_12308);
nor U13752 (N_13752,N_11260,N_11072);
or U13753 (N_13753,N_11510,N_10588);
and U13754 (N_13754,N_12353,N_12082);
or U13755 (N_13755,N_10451,N_11550);
and U13756 (N_13756,N_11302,N_10128);
or U13757 (N_13757,N_10222,N_12253);
nand U13758 (N_13758,N_10200,N_11182);
nand U13759 (N_13759,N_10634,N_12297);
nand U13760 (N_13760,N_11763,N_11715);
nor U13761 (N_13761,N_11715,N_11382);
or U13762 (N_13762,N_10416,N_11630);
and U13763 (N_13763,N_10884,N_10110);
and U13764 (N_13764,N_10054,N_11621);
and U13765 (N_13765,N_11702,N_10930);
and U13766 (N_13766,N_11511,N_10835);
and U13767 (N_13767,N_10807,N_10151);
nand U13768 (N_13768,N_10402,N_11267);
and U13769 (N_13769,N_12246,N_10386);
nor U13770 (N_13770,N_11730,N_11935);
and U13771 (N_13771,N_12155,N_12002);
and U13772 (N_13772,N_11196,N_11734);
nor U13773 (N_13773,N_10407,N_10870);
nor U13774 (N_13774,N_11220,N_12308);
and U13775 (N_13775,N_10397,N_11111);
nand U13776 (N_13776,N_11796,N_10250);
nor U13777 (N_13777,N_10222,N_11609);
nor U13778 (N_13778,N_10212,N_11161);
or U13779 (N_13779,N_11546,N_10991);
or U13780 (N_13780,N_12366,N_12304);
nor U13781 (N_13781,N_10233,N_10671);
nand U13782 (N_13782,N_11805,N_10094);
nor U13783 (N_13783,N_12491,N_11433);
nor U13784 (N_13784,N_10007,N_12416);
or U13785 (N_13785,N_10823,N_11881);
or U13786 (N_13786,N_11839,N_11716);
nor U13787 (N_13787,N_11768,N_10939);
nor U13788 (N_13788,N_11246,N_10598);
xnor U13789 (N_13789,N_12049,N_11965);
nand U13790 (N_13790,N_11678,N_11647);
nor U13791 (N_13791,N_12028,N_10827);
nor U13792 (N_13792,N_12470,N_10888);
and U13793 (N_13793,N_10393,N_10697);
nor U13794 (N_13794,N_11880,N_12290);
nor U13795 (N_13795,N_11255,N_12068);
nand U13796 (N_13796,N_12315,N_11942);
nor U13797 (N_13797,N_12264,N_11432);
nand U13798 (N_13798,N_10422,N_10074);
or U13799 (N_13799,N_10978,N_11172);
nand U13800 (N_13800,N_10421,N_10923);
nand U13801 (N_13801,N_12053,N_10342);
nand U13802 (N_13802,N_11974,N_11939);
nor U13803 (N_13803,N_10982,N_11471);
xnor U13804 (N_13804,N_12274,N_12395);
nor U13805 (N_13805,N_11011,N_12053);
or U13806 (N_13806,N_11604,N_11924);
nor U13807 (N_13807,N_12058,N_11209);
nand U13808 (N_13808,N_11176,N_12481);
or U13809 (N_13809,N_12163,N_10462);
or U13810 (N_13810,N_10513,N_11042);
nand U13811 (N_13811,N_10078,N_11088);
and U13812 (N_13812,N_10684,N_12060);
nor U13813 (N_13813,N_11827,N_11293);
and U13814 (N_13814,N_10875,N_12071);
or U13815 (N_13815,N_12297,N_12321);
nand U13816 (N_13816,N_11062,N_11941);
nor U13817 (N_13817,N_12064,N_11132);
and U13818 (N_13818,N_10202,N_12144);
nor U13819 (N_13819,N_10543,N_12280);
nor U13820 (N_13820,N_12466,N_11939);
nor U13821 (N_13821,N_12450,N_12328);
and U13822 (N_13822,N_11306,N_11483);
and U13823 (N_13823,N_10159,N_10598);
or U13824 (N_13824,N_12394,N_10800);
or U13825 (N_13825,N_10640,N_12280);
or U13826 (N_13826,N_12376,N_10038);
nor U13827 (N_13827,N_11453,N_10017);
nor U13828 (N_13828,N_11785,N_11833);
nor U13829 (N_13829,N_10917,N_12161);
or U13830 (N_13830,N_10416,N_10865);
nand U13831 (N_13831,N_11244,N_10061);
or U13832 (N_13832,N_11772,N_10874);
nor U13833 (N_13833,N_11965,N_12354);
nand U13834 (N_13834,N_10135,N_10643);
and U13835 (N_13835,N_11071,N_11716);
nor U13836 (N_13836,N_11129,N_10669);
nor U13837 (N_13837,N_10094,N_11831);
nor U13838 (N_13838,N_10449,N_10811);
or U13839 (N_13839,N_12120,N_10425);
nor U13840 (N_13840,N_11478,N_10186);
or U13841 (N_13841,N_10851,N_12199);
nor U13842 (N_13842,N_11441,N_10634);
nand U13843 (N_13843,N_11216,N_11479);
or U13844 (N_13844,N_12116,N_11367);
or U13845 (N_13845,N_10485,N_12036);
or U13846 (N_13846,N_10356,N_11103);
nor U13847 (N_13847,N_12374,N_10469);
and U13848 (N_13848,N_11459,N_10502);
nand U13849 (N_13849,N_11259,N_11708);
nor U13850 (N_13850,N_11664,N_10116);
and U13851 (N_13851,N_10661,N_10246);
and U13852 (N_13852,N_10057,N_10849);
nand U13853 (N_13853,N_12497,N_10910);
nor U13854 (N_13854,N_11003,N_11730);
and U13855 (N_13855,N_11492,N_12243);
nor U13856 (N_13856,N_10621,N_10740);
and U13857 (N_13857,N_12021,N_10250);
nand U13858 (N_13858,N_11477,N_10689);
nand U13859 (N_13859,N_11138,N_11502);
or U13860 (N_13860,N_10800,N_10554);
or U13861 (N_13861,N_11005,N_11798);
or U13862 (N_13862,N_12147,N_11718);
or U13863 (N_13863,N_11653,N_12091);
or U13864 (N_13864,N_11191,N_11918);
or U13865 (N_13865,N_12162,N_11376);
or U13866 (N_13866,N_11683,N_10929);
nor U13867 (N_13867,N_10155,N_11455);
nor U13868 (N_13868,N_11500,N_11286);
and U13869 (N_13869,N_12361,N_11023);
nor U13870 (N_13870,N_12455,N_10838);
nor U13871 (N_13871,N_10374,N_10390);
or U13872 (N_13872,N_10157,N_12472);
nor U13873 (N_13873,N_11061,N_10624);
or U13874 (N_13874,N_11094,N_10850);
and U13875 (N_13875,N_11173,N_11725);
or U13876 (N_13876,N_11082,N_11561);
or U13877 (N_13877,N_10433,N_10318);
and U13878 (N_13878,N_10907,N_11930);
or U13879 (N_13879,N_11148,N_12034);
and U13880 (N_13880,N_10704,N_10358);
nand U13881 (N_13881,N_11400,N_10998);
or U13882 (N_13882,N_12355,N_12476);
nor U13883 (N_13883,N_10632,N_11856);
nand U13884 (N_13884,N_11025,N_11850);
nor U13885 (N_13885,N_12415,N_10936);
and U13886 (N_13886,N_10493,N_10175);
and U13887 (N_13887,N_10757,N_11982);
nor U13888 (N_13888,N_11606,N_12277);
nor U13889 (N_13889,N_11398,N_10566);
nor U13890 (N_13890,N_12075,N_10716);
and U13891 (N_13891,N_11836,N_10003);
nand U13892 (N_13892,N_10918,N_11439);
nand U13893 (N_13893,N_10452,N_12462);
nor U13894 (N_13894,N_11389,N_11562);
nand U13895 (N_13895,N_12308,N_11699);
nand U13896 (N_13896,N_12246,N_11455);
or U13897 (N_13897,N_11472,N_11205);
or U13898 (N_13898,N_11844,N_11103);
nor U13899 (N_13899,N_11530,N_11240);
and U13900 (N_13900,N_11625,N_11918);
nor U13901 (N_13901,N_11405,N_11498);
or U13902 (N_13902,N_10922,N_11947);
or U13903 (N_13903,N_12100,N_12013);
nor U13904 (N_13904,N_10797,N_10697);
and U13905 (N_13905,N_11635,N_10264);
and U13906 (N_13906,N_10745,N_11102);
nand U13907 (N_13907,N_10353,N_12476);
nor U13908 (N_13908,N_12309,N_11672);
nor U13909 (N_13909,N_11358,N_11721);
or U13910 (N_13910,N_12092,N_11014);
or U13911 (N_13911,N_11661,N_11248);
and U13912 (N_13912,N_10481,N_10741);
and U13913 (N_13913,N_11128,N_10190);
or U13914 (N_13914,N_11918,N_10640);
nand U13915 (N_13915,N_12457,N_11883);
and U13916 (N_13916,N_12002,N_10693);
nand U13917 (N_13917,N_10624,N_12105);
nand U13918 (N_13918,N_11514,N_12390);
nand U13919 (N_13919,N_11581,N_11844);
nor U13920 (N_13920,N_10764,N_11798);
or U13921 (N_13921,N_12214,N_11590);
nand U13922 (N_13922,N_10129,N_10433);
or U13923 (N_13923,N_11524,N_10970);
or U13924 (N_13924,N_10349,N_11302);
nor U13925 (N_13925,N_11841,N_11854);
nor U13926 (N_13926,N_11641,N_10128);
or U13927 (N_13927,N_11471,N_10114);
and U13928 (N_13928,N_12185,N_12472);
or U13929 (N_13929,N_11237,N_11303);
nor U13930 (N_13930,N_10056,N_12109);
and U13931 (N_13931,N_10191,N_11107);
nand U13932 (N_13932,N_11835,N_11717);
or U13933 (N_13933,N_12148,N_11887);
or U13934 (N_13934,N_11005,N_10254);
nor U13935 (N_13935,N_11308,N_11687);
nand U13936 (N_13936,N_11231,N_11278);
xor U13937 (N_13937,N_10989,N_11129);
or U13938 (N_13938,N_11584,N_10324);
nand U13939 (N_13939,N_11167,N_12164);
or U13940 (N_13940,N_10901,N_12224);
nor U13941 (N_13941,N_10025,N_10806);
or U13942 (N_13942,N_11664,N_10005);
or U13943 (N_13943,N_11570,N_11723);
or U13944 (N_13944,N_10103,N_11471);
or U13945 (N_13945,N_10573,N_11995);
and U13946 (N_13946,N_10609,N_10144);
or U13947 (N_13947,N_10410,N_12377);
and U13948 (N_13948,N_10349,N_10548);
or U13949 (N_13949,N_11221,N_10799);
and U13950 (N_13950,N_11047,N_10172);
and U13951 (N_13951,N_10466,N_10932);
nand U13952 (N_13952,N_12050,N_11695);
nand U13953 (N_13953,N_10872,N_11872);
and U13954 (N_13954,N_12296,N_11832);
nor U13955 (N_13955,N_11875,N_10826);
nor U13956 (N_13956,N_11440,N_10507);
nor U13957 (N_13957,N_11616,N_12125);
nand U13958 (N_13958,N_11837,N_10768);
nor U13959 (N_13959,N_11559,N_11012);
and U13960 (N_13960,N_12044,N_11145);
or U13961 (N_13961,N_10168,N_12317);
nand U13962 (N_13962,N_10250,N_12051);
nand U13963 (N_13963,N_11721,N_10790);
nor U13964 (N_13964,N_11418,N_12354);
or U13965 (N_13965,N_10751,N_11349);
and U13966 (N_13966,N_12309,N_11406);
and U13967 (N_13967,N_10622,N_11776);
nor U13968 (N_13968,N_11294,N_12153);
and U13969 (N_13969,N_10331,N_12499);
or U13970 (N_13970,N_12219,N_11594);
and U13971 (N_13971,N_11656,N_10558);
nand U13972 (N_13972,N_10934,N_11109);
and U13973 (N_13973,N_12339,N_12452);
nor U13974 (N_13974,N_11442,N_10616);
nor U13975 (N_13975,N_11060,N_11237);
and U13976 (N_13976,N_11766,N_11332);
nor U13977 (N_13977,N_10639,N_11185);
and U13978 (N_13978,N_12092,N_10618);
nand U13979 (N_13979,N_11171,N_10264);
or U13980 (N_13980,N_10205,N_12096);
or U13981 (N_13981,N_10598,N_12388);
or U13982 (N_13982,N_12180,N_11082);
nor U13983 (N_13983,N_11500,N_10840);
nand U13984 (N_13984,N_11029,N_12034);
and U13985 (N_13985,N_11386,N_11069);
and U13986 (N_13986,N_11662,N_10516);
and U13987 (N_13987,N_12187,N_10051);
nand U13988 (N_13988,N_10071,N_10136);
nand U13989 (N_13989,N_10455,N_11707);
or U13990 (N_13990,N_10521,N_10292);
or U13991 (N_13991,N_11808,N_11751);
and U13992 (N_13992,N_10502,N_12333);
nor U13993 (N_13993,N_12333,N_11230);
and U13994 (N_13994,N_11684,N_12275);
nand U13995 (N_13995,N_10372,N_10135);
or U13996 (N_13996,N_10434,N_11769);
or U13997 (N_13997,N_11204,N_11722);
nand U13998 (N_13998,N_12221,N_10165);
nand U13999 (N_13999,N_12231,N_11485);
nand U14000 (N_14000,N_11307,N_10304);
or U14001 (N_14001,N_11278,N_10142);
and U14002 (N_14002,N_10699,N_11871);
nor U14003 (N_14003,N_11848,N_10808);
nor U14004 (N_14004,N_11121,N_10580);
and U14005 (N_14005,N_11792,N_12244);
nand U14006 (N_14006,N_11482,N_12378);
or U14007 (N_14007,N_10111,N_11131);
and U14008 (N_14008,N_11672,N_11888);
nand U14009 (N_14009,N_10379,N_12086);
nor U14010 (N_14010,N_11885,N_11062);
or U14011 (N_14011,N_11394,N_10387);
and U14012 (N_14012,N_10584,N_11296);
or U14013 (N_14013,N_10858,N_10370);
nor U14014 (N_14014,N_12208,N_11708);
or U14015 (N_14015,N_12354,N_11789);
nor U14016 (N_14016,N_12395,N_10124);
and U14017 (N_14017,N_10273,N_11757);
and U14018 (N_14018,N_11655,N_11230);
nand U14019 (N_14019,N_11778,N_11554);
nand U14020 (N_14020,N_12107,N_11706);
and U14021 (N_14021,N_11868,N_10953);
xor U14022 (N_14022,N_11184,N_11312);
nor U14023 (N_14023,N_11722,N_11775);
nor U14024 (N_14024,N_10255,N_11354);
nor U14025 (N_14025,N_11780,N_10588);
or U14026 (N_14026,N_10351,N_10015);
nand U14027 (N_14027,N_12178,N_10468);
or U14028 (N_14028,N_10525,N_11705);
or U14029 (N_14029,N_12345,N_10737);
nor U14030 (N_14030,N_11248,N_10454);
or U14031 (N_14031,N_10988,N_12257);
and U14032 (N_14032,N_10304,N_11542);
or U14033 (N_14033,N_11606,N_11894);
nand U14034 (N_14034,N_11203,N_10359);
nand U14035 (N_14035,N_12452,N_10952);
nand U14036 (N_14036,N_10762,N_11017);
nor U14037 (N_14037,N_11436,N_12367);
or U14038 (N_14038,N_10895,N_11976);
or U14039 (N_14039,N_11512,N_10157);
nand U14040 (N_14040,N_11084,N_10006);
nand U14041 (N_14041,N_10484,N_11748);
and U14042 (N_14042,N_10843,N_11829);
or U14043 (N_14043,N_10187,N_10155);
nor U14044 (N_14044,N_11008,N_10527);
nor U14045 (N_14045,N_10506,N_11333);
nand U14046 (N_14046,N_11257,N_10948);
nor U14047 (N_14047,N_11245,N_11205);
nor U14048 (N_14048,N_10253,N_11725);
nor U14049 (N_14049,N_12113,N_10566);
nand U14050 (N_14050,N_11113,N_12151);
or U14051 (N_14051,N_10500,N_12219);
nand U14052 (N_14052,N_11018,N_10626);
nor U14053 (N_14053,N_10773,N_10215);
nand U14054 (N_14054,N_11048,N_11772);
nand U14055 (N_14055,N_11547,N_11251);
or U14056 (N_14056,N_12483,N_10428);
and U14057 (N_14057,N_11413,N_11755);
nand U14058 (N_14058,N_10991,N_11410);
and U14059 (N_14059,N_12309,N_10396);
and U14060 (N_14060,N_10476,N_11636);
nand U14061 (N_14061,N_10373,N_11801);
nand U14062 (N_14062,N_11484,N_11382);
or U14063 (N_14063,N_10564,N_11425);
nor U14064 (N_14064,N_10909,N_12413);
and U14065 (N_14065,N_10922,N_11860);
nand U14066 (N_14066,N_12087,N_12402);
or U14067 (N_14067,N_11919,N_10651);
nor U14068 (N_14068,N_11167,N_10884);
nor U14069 (N_14069,N_11525,N_10107);
and U14070 (N_14070,N_12305,N_11721);
and U14071 (N_14071,N_10834,N_10310);
nand U14072 (N_14072,N_11337,N_11551);
nand U14073 (N_14073,N_11088,N_10270);
nor U14074 (N_14074,N_10672,N_11559);
and U14075 (N_14075,N_11659,N_10198);
nor U14076 (N_14076,N_12428,N_12454);
nor U14077 (N_14077,N_10522,N_11245);
or U14078 (N_14078,N_10149,N_12192);
and U14079 (N_14079,N_12140,N_12376);
nand U14080 (N_14080,N_11627,N_11639);
or U14081 (N_14081,N_11690,N_10225);
or U14082 (N_14082,N_12289,N_11312);
nor U14083 (N_14083,N_11112,N_11160);
or U14084 (N_14084,N_10269,N_11823);
nand U14085 (N_14085,N_10638,N_11356);
nand U14086 (N_14086,N_11603,N_11630);
nor U14087 (N_14087,N_10054,N_11270);
and U14088 (N_14088,N_10084,N_11096);
nand U14089 (N_14089,N_12111,N_11882);
nand U14090 (N_14090,N_11526,N_11946);
or U14091 (N_14091,N_12337,N_11555);
nand U14092 (N_14092,N_12092,N_11275);
or U14093 (N_14093,N_11860,N_10609);
and U14094 (N_14094,N_11888,N_12251);
and U14095 (N_14095,N_11329,N_12103);
nor U14096 (N_14096,N_11987,N_10692);
or U14097 (N_14097,N_10585,N_10544);
and U14098 (N_14098,N_10821,N_10189);
or U14099 (N_14099,N_11571,N_10909);
and U14100 (N_14100,N_10893,N_10734);
and U14101 (N_14101,N_11365,N_11495);
and U14102 (N_14102,N_11088,N_12037);
and U14103 (N_14103,N_10825,N_11346);
and U14104 (N_14104,N_10294,N_12474);
or U14105 (N_14105,N_10759,N_10590);
and U14106 (N_14106,N_10409,N_10926);
and U14107 (N_14107,N_10553,N_11642);
nand U14108 (N_14108,N_11826,N_12389);
or U14109 (N_14109,N_12212,N_12411);
and U14110 (N_14110,N_10135,N_10360);
nand U14111 (N_14111,N_12411,N_10146);
or U14112 (N_14112,N_10535,N_11973);
nor U14113 (N_14113,N_11995,N_12090);
or U14114 (N_14114,N_10590,N_11005);
or U14115 (N_14115,N_12425,N_10427);
and U14116 (N_14116,N_11617,N_10887);
nor U14117 (N_14117,N_10669,N_11447);
nand U14118 (N_14118,N_11073,N_10337);
nand U14119 (N_14119,N_10213,N_10327);
nor U14120 (N_14120,N_11848,N_11359);
or U14121 (N_14121,N_11248,N_12238);
nor U14122 (N_14122,N_10687,N_11005);
nand U14123 (N_14123,N_12371,N_12184);
and U14124 (N_14124,N_10318,N_11260);
or U14125 (N_14125,N_10390,N_11712);
and U14126 (N_14126,N_11100,N_11893);
or U14127 (N_14127,N_10775,N_11090);
or U14128 (N_14128,N_11864,N_10668);
and U14129 (N_14129,N_11939,N_10929);
nor U14130 (N_14130,N_10066,N_10949);
and U14131 (N_14131,N_10425,N_10874);
and U14132 (N_14132,N_12367,N_11124);
nand U14133 (N_14133,N_11457,N_10201);
nand U14134 (N_14134,N_10770,N_10100);
or U14135 (N_14135,N_10409,N_12304);
or U14136 (N_14136,N_12050,N_12234);
and U14137 (N_14137,N_11487,N_10177);
nand U14138 (N_14138,N_12394,N_11176);
nor U14139 (N_14139,N_11209,N_11502);
and U14140 (N_14140,N_11189,N_10858);
and U14141 (N_14141,N_10356,N_10036);
or U14142 (N_14142,N_10000,N_11650);
nand U14143 (N_14143,N_11924,N_11309);
nor U14144 (N_14144,N_11669,N_11083);
and U14145 (N_14145,N_11920,N_10450);
and U14146 (N_14146,N_11114,N_10083);
and U14147 (N_14147,N_11482,N_10955);
nor U14148 (N_14148,N_10051,N_10736);
or U14149 (N_14149,N_10643,N_10398);
or U14150 (N_14150,N_11506,N_10015);
nor U14151 (N_14151,N_10898,N_12224);
nor U14152 (N_14152,N_10998,N_11137);
nor U14153 (N_14153,N_10481,N_12016);
and U14154 (N_14154,N_10929,N_11841);
nand U14155 (N_14155,N_11393,N_10224);
and U14156 (N_14156,N_12197,N_12247);
nand U14157 (N_14157,N_11957,N_10805);
nand U14158 (N_14158,N_11978,N_10945);
nor U14159 (N_14159,N_12231,N_12122);
and U14160 (N_14160,N_10333,N_10374);
and U14161 (N_14161,N_11273,N_11772);
and U14162 (N_14162,N_11509,N_11680);
nand U14163 (N_14163,N_10165,N_11108);
nor U14164 (N_14164,N_10504,N_10693);
nor U14165 (N_14165,N_12225,N_10970);
nand U14166 (N_14166,N_12032,N_11941);
and U14167 (N_14167,N_11256,N_11550);
or U14168 (N_14168,N_11100,N_12475);
nand U14169 (N_14169,N_11826,N_11550);
nand U14170 (N_14170,N_12005,N_10497);
and U14171 (N_14171,N_10396,N_11866);
or U14172 (N_14172,N_10242,N_12431);
nand U14173 (N_14173,N_12176,N_10011);
and U14174 (N_14174,N_11862,N_11282);
nand U14175 (N_14175,N_11922,N_12167);
nor U14176 (N_14176,N_12181,N_11087);
nor U14177 (N_14177,N_10588,N_12242);
or U14178 (N_14178,N_10421,N_12101);
or U14179 (N_14179,N_11623,N_12250);
nor U14180 (N_14180,N_12051,N_10545);
nor U14181 (N_14181,N_11224,N_10800);
nand U14182 (N_14182,N_11771,N_12484);
and U14183 (N_14183,N_10681,N_10552);
and U14184 (N_14184,N_10221,N_11409);
and U14185 (N_14185,N_12108,N_11481);
and U14186 (N_14186,N_12059,N_11436);
or U14187 (N_14187,N_11801,N_11122);
and U14188 (N_14188,N_12149,N_11820);
nor U14189 (N_14189,N_10640,N_11264);
or U14190 (N_14190,N_11100,N_10783);
nand U14191 (N_14191,N_10982,N_11723);
nor U14192 (N_14192,N_12245,N_10167);
nand U14193 (N_14193,N_10551,N_12459);
or U14194 (N_14194,N_12088,N_12022);
and U14195 (N_14195,N_10647,N_11964);
or U14196 (N_14196,N_11304,N_12179);
or U14197 (N_14197,N_11153,N_11405);
or U14198 (N_14198,N_11562,N_11460);
nor U14199 (N_14199,N_10908,N_11618);
and U14200 (N_14200,N_11568,N_12419);
and U14201 (N_14201,N_11546,N_11083);
or U14202 (N_14202,N_12099,N_10971);
nand U14203 (N_14203,N_12042,N_10700);
or U14204 (N_14204,N_10833,N_11291);
nand U14205 (N_14205,N_12432,N_11721);
and U14206 (N_14206,N_11616,N_10868);
nor U14207 (N_14207,N_11992,N_10654);
and U14208 (N_14208,N_12115,N_11671);
nor U14209 (N_14209,N_12434,N_10155);
and U14210 (N_14210,N_10451,N_11688);
nor U14211 (N_14211,N_12267,N_10941);
or U14212 (N_14212,N_11495,N_10654);
or U14213 (N_14213,N_11340,N_10526);
xor U14214 (N_14214,N_11834,N_10472);
or U14215 (N_14215,N_12167,N_12107);
and U14216 (N_14216,N_11091,N_11737);
nor U14217 (N_14217,N_10415,N_12009);
xnor U14218 (N_14218,N_10776,N_11936);
and U14219 (N_14219,N_10947,N_12258);
nand U14220 (N_14220,N_10723,N_10618);
and U14221 (N_14221,N_10523,N_12468);
or U14222 (N_14222,N_10289,N_11392);
or U14223 (N_14223,N_10453,N_10359);
nor U14224 (N_14224,N_11162,N_10340);
nand U14225 (N_14225,N_11881,N_11945);
nor U14226 (N_14226,N_12147,N_10985);
or U14227 (N_14227,N_12481,N_12088);
nand U14228 (N_14228,N_11190,N_10029);
nand U14229 (N_14229,N_11785,N_12264);
nor U14230 (N_14230,N_12358,N_11294);
or U14231 (N_14231,N_11327,N_11220);
nor U14232 (N_14232,N_11500,N_10097);
or U14233 (N_14233,N_10930,N_10407);
nand U14234 (N_14234,N_10489,N_12339);
and U14235 (N_14235,N_10394,N_10206);
nor U14236 (N_14236,N_10644,N_10659);
nand U14237 (N_14237,N_11569,N_12466);
nand U14238 (N_14238,N_11801,N_12358);
nor U14239 (N_14239,N_11149,N_12152);
nor U14240 (N_14240,N_11896,N_10906);
and U14241 (N_14241,N_10981,N_11624);
nor U14242 (N_14242,N_12388,N_10583);
and U14243 (N_14243,N_11378,N_11161);
and U14244 (N_14244,N_11221,N_10485);
and U14245 (N_14245,N_11244,N_11263);
nor U14246 (N_14246,N_12208,N_11737);
nand U14247 (N_14247,N_11377,N_11679);
or U14248 (N_14248,N_10784,N_11755);
xnor U14249 (N_14249,N_11376,N_11036);
or U14250 (N_14250,N_11309,N_10819);
or U14251 (N_14251,N_11882,N_11588);
or U14252 (N_14252,N_12165,N_11159);
nand U14253 (N_14253,N_10745,N_10010);
nor U14254 (N_14254,N_10940,N_11573);
or U14255 (N_14255,N_11550,N_11096);
nand U14256 (N_14256,N_10327,N_12359);
nand U14257 (N_14257,N_12370,N_10002);
xnor U14258 (N_14258,N_10024,N_10386);
and U14259 (N_14259,N_10153,N_10713);
nand U14260 (N_14260,N_11955,N_10557);
nor U14261 (N_14261,N_10939,N_12078);
nor U14262 (N_14262,N_12357,N_11667);
nor U14263 (N_14263,N_10388,N_10672);
nor U14264 (N_14264,N_11493,N_10003);
nand U14265 (N_14265,N_11083,N_11304);
nor U14266 (N_14266,N_10542,N_10805);
nand U14267 (N_14267,N_12128,N_11917);
and U14268 (N_14268,N_10394,N_10498);
and U14269 (N_14269,N_12391,N_11820);
and U14270 (N_14270,N_10743,N_12015);
or U14271 (N_14271,N_11895,N_11538);
nor U14272 (N_14272,N_10883,N_12223);
and U14273 (N_14273,N_11263,N_11582);
nor U14274 (N_14274,N_10590,N_12373);
nor U14275 (N_14275,N_10194,N_10061);
nor U14276 (N_14276,N_11937,N_10440);
nand U14277 (N_14277,N_11903,N_11402);
nor U14278 (N_14278,N_10843,N_12458);
nand U14279 (N_14279,N_10545,N_10073);
nor U14280 (N_14280,N_12443,N_10426);
or U14281 (N_14281,N_12287,N_10402);
xnor U14282 (N_14282,N_11689,N_12487);
nand U14283 (N_14283,N_11858,N_12171);
nand U14284 (N_14284,N_12045,N_11126);
and U14285 (N_14285,N_10885,N_10738);
nand U14286 (N_14286,N_10962,N_11047);
nand U14287 (N_14287,N_12324,N_10599);
or U14288 (N_14288,N_11282,N_10961);
and U14289 (N_14289,N_11466,N_11497);
or U14290 (N_14290,N_11351,N_11414);
nand U14291 (N_14291,N_11519,N_10011);
or U14292 (N_14292,N_12112,N_11108);
or U14293 (N_14293,N_12082,N_10024);
nor U14294 (N_14294,N_11428,N_12416);
or U14295 (N_14295,N_11973,N_11210);
or U14296 (N_14296,N_11607,N_12389);
or U14297 (N_14297,N_10679,N_10184);
or U14298 (N_14298,N_12099,N_12018);
and U14299 (N_14299,N_10344,N_12016);
nor U14300 (N_14300,N_10383,N_10250);
nor U14301 (N_14301,N_10496,N_12280);
nand U14302 (N_14302,N_12412,N_10479);
nand U14303 (N_14303,N_12000,N_11735);
and U14304 (N_14304,N_10819,N_10791);
or U14305 (N_14305,N_10952,N_10343);
and U14306 (N_14306,N_10093,N_11042);
or U14307 (N_14307,N_11907,N_12193);
and U14308 (N_14308,N_11238,N_11621);
or U14309 (N_14309,N_10752,N_10445);
and U14310 (N_14310,N_12234,N_11490);
and U14311 (N_14311,N_11600,N_11449);
nor U14312 (N_14312,N_12052,N_11004);
and U14313 (N_14313,N_11371,N_11319);
nor U14314 (N_14314,N_10709,N_10279);
nor U14315 (N_14315,N_10607,N_11071);
nor U14316 (N_14316,N_11979,N_11288);
and U14317 (N_14317,N_12492,N_12167);
and U14318 (N_14318,N_11911,N_10891);
or U14319 (N_14319,N_11445,N_10483);
or U14320 (N_14320,N_10048,N_10390);
or U14321 (N_14321,N_11723,N_11607);
nor U14322 (N_14322,N_10102,N_10983);
nor U14323 (N_14323,N_12363,N_11107);
nor U14324 (N_14324,N_12386,N_12383);
nor U14325 (N_14325,N_10927,N_11201);
or U14326 (N_14326,N_12227,N_11076);
nor U14327 (N_14327,N_12138,N_10386);
nand U14328 (N_14328,N_10761,N_11925);
nor U14329 (N_14329,N_11537,N_10038);
and U14330 (N_14330,N_10327,N_11342);
nor U14331 (N_14331,N_12229,N_11822);
nand U14332 (N_14332,N_11270,N_11157);
and U14333 (N_14333,N_10570,N_10222);
nand U14334 (N_14334,N_11943,N_11892);
or U14335 (N_14335,N_11801,N_12244);
nand U14336 (N_14336,N_10862,N_12147);
or U14337 (N_14337,N_11931,N_11234);
nand U14338 (N_14338,N_12427,N_12400);
and U14339 (N_14339,N_10944,N_10655);
and U14340 (N_14340,N_12248,N_11760);
and U14341 (N_14341,N_10832,N_11200);
nor U14342 (N_14342,N_10114,N_11060);
nor U14343 (N_14343,N_11289,N_11014);
nor U14344 (N_14344,N_10351,N_12161);
nor U14345 (N_14345,N_10351,N_11863);
nand U14346 (N_14346,N_11856,N_11089);
or U14347 (N_14347,N_11220,N_10308);
or U14348 (N_14348,N_12170,N_10076);
nor U14349 (N_14349,N_10231,N_10182);
xor U14350 (N_14350,N_12223,N_10312);
or U14351 (N_14351,N_10793,N_10716);
nor U14352 (N_14352,N_12005,N_11171);
xor U14353 (N_14353,N_11773,N_11028);
nand U14354 (N_14354,N_11905,N_12374);
nand U14355 (N_14355,N_10354,N_11596);
nor U14356 (N_14356,N_12246,N_11291);
and U14357 (N_14357,N_10040,N_10860);
nand U14358 (N_14358,N_10129,N_10720);
nor U14359 (N_14359,N_10083,N_10262);
or U14360 (N_14360,N_10535,N_10237);
and U14361 (N_14361,N_11556,N_11869);
and U14362 (N_14362,N_11371,N_10733);
nand U14363 (N_14363,N_10072,N_11559);
nor U14364 (N_14364,N_10223,N_11506);
and U14365 (N_14365,N_10895,N_11074);
or U14366 (N_14366,N_11685,N_11729);
or U14367 (N_14367,N_12014,N_11785);
and U14368 (N_14368,N_10947,N_10103);
nand U14369 (N_14369,N_10753,N_11603);
or U14370 (N_14370,N_11865,N_12408);
and U14371 (N_14371,N_10038,N_11064);
nand U14372 (N_14372,N_11378,N_10321);
nor U14373 (N_14373,N_11526,N_11166);
nor U14374 (N_14374,N_12446,N_12061);
or U14375 (N_14375,N_11455,N_10509);
nand U14376 (N_14376,N_10201,N_12204);
or U14377 (N_14377,N_11346,N_10882);
or U14378 (N_14378,N_11952,N_10334);
or U14379 (N_14379,N_10837,N_10827);
and U14380 (N_14380,N_10275,N_10481);
nand U14381 (N_14381,N_10192,N_12002);
or U14382 (N_14382,N_12006,N_10761);
or U14383 (N_14383,N_10455,N_10186);
nor U14384 (N_14384,N_10196,N_11164);
and U14385 (N_14385,N_10664,N_12316);
or U14386 (N_14386,N_10046,N_10217);
and U14387 (N_14387,N_11226,N_10521);
nand U14388 (N_14388,N_12260,N_10775);
nand U14389 (N_14389,N_10169,N_11345);
and U14390 (N_14390,N_11983,N_12030);
or U14391 (N_14391,N_11579,N_11120);
nor U14392 (N_14392,N_10977,N_11153);
and U14393 (N_14393,N_10937,N_12475);
nand U14394 (N_14394,N_10504,N_11927);
and U14395 (N_14395,N_10070,N_10255);
nand U14396 (N_14396,N_11128,N_10177);
and U14397 (N_14397,N_10561,N_10508);
and U14398 (N_14398,N_11941,N_11738);
or U14399 (N_14399,N_12432,N_11131);
nor U14400 (N_14400,N_10509,N_10038);
nor U14401 (N_14401,N_10826,N_10224);
nor U14402 (N_14402,N_11201,N_12224);
or U14403 (N_14403,N_11330,N_11791);
nor U14404 (N_14404,N_11096,N_11136);
or U14405 (N_14405,N_10310,N_10380);
and U14406 (N_14406,N_11300,N_10223);
or U14407 (N_14407,N_10113,N_12062);
or U14408 (N_14408,N_10578,N_11433);
and U14409 (N_14409,N_12313,N_11674);
or U14410 (N_14410,N_10052,N_12429);
nor U14411 (N_14411,N_10164,N_11990);
nor U14412 (N_14412,N_10612,N_11059);
and U14413 (N_14413,N_11885,N_10146);
and U14414 (N_14414,N_10028,N_10723);
xor U14415 (N_14415,N_10859,N_11817);
and U14416 (N_14416,N_10951,N_10469);
or U14417 (N_14417,N_11375,N_10503);
nand U14418 (N_14418,N_10424,N_11098);
and U14419 (N_14419,N_12392,N_11711);
and U14420 (N_14420,N_11554,N_10807);
and U14421 (N_14421,N_11422,N_11919);
nand U14422 (N_14422,N_10666,N_11932);
nor U14423 (N_14423,N_11244,N_11073);
nor U14424 (N_14424,N_11964,N_11332);
and U14425 (N_14425,N_10705,N_10820);
nand U14426 (N_14426,N_12060,N_11441);
nor U14427 (N_14427,N_11308,N_10735);
and U14428 (N_14428,N_10567,N_11416);
and U14429 (N_14429,N_10765,N_12456);
or U14430 (N_14430,N_10921,N_12214);
nand U14431 (N_14431,N_12419,N_10739);
or U14432 (N_14432,N_10495,N_11032);
and U14433 (N_14433,N_11842,N_10117);
or U14434 (N_14434,N_10791,N_10041);
and U14435 (N_14435,N_11628,N_11476);
and U14436 (N_14436,N_10635,N_10954);
nor U14437 (N_14437,N_11445,N_10148);
nor U14438 (N_14438,N_10394,N_12362);
nor U14439 (N_14439,N_12138,N_10671);
nor U14440 (N_14440,N_11576,N_12315);
nand U14441 (N_14441,N_10539,N_10602);
and U14442 (N_14442,N_10024,N_10675);
nand U14443 (N_14443,N_10464,N_12028);
and U14444 (N_14444,N_10411,N_11982);
and U14445 (N_14445,N_11925,N_10481);
nor U14446 (N_14446,N_10407,N_12390);
and U14447 (N_14447,N_10476,N_10906);
or U14448 (N_14448,N_10701,N_10581);
nand U14449 (N_14449,N_10026,N_10358);
nand U14450 (N_14450,N_11522,N_11625);
or U14451 (N_14451,N_10440,N_11722);
nand U14452 (N_14452,N_10253,N_12497);
nand U14453 (N_14453,N_11241,N_12188);
nand U14454 (N_14454,N_10710,N_10175);
nor U14455 (N_14455,N_11006,N_12330);
and U14456 (N_14456,N_12206,N_10566);
nor U14457 (N_14457,N_11062,N_10542);
nor U14458 (N_14458,N_10969,N_10798);
and U14459 (N_14459,N_11056,N_11355);
or U14460 (N_14460,N_11018,N_10909);
nand U14461 (N_14461,N_10712,N_11109);
or U14462 (N_14462,N_12357,N_12387);
nand U14463 (N_14463,N_10586,N_12219);
or U14464 (N_14464,N_10647,N_11345);
nor U14465 (N_14465,N_11853,N_10651);
or U14466 (N_14466,N_10940,N_11494);
nand U14467 (N_14467,N_12236,N_12026);
xnor U14468 (N_14468,N_10052,N_12338);
nor U14469 (N_14469,N_12002,N_12172);
nor U14470 (N_14470,N_11027,N_10145);
and U14471 (N_14471,N_10449,N_10612);
nor U14472 (N_14472,N_10584,N_11206);
nor U14473 (N_14473,N_12068,N_12026);
or U14474 (N_14474,N_10182,N_10226);
or U14475 (N_14475,N_11912,N_11571);
and U14476 (N_14476,N_10751,N_11740);
nor U14477 (N_14477,N_11320,N_11457);
nor U14478 (N_14478,N_12344,N_11599);
nand U14479 (N_14479,N_10634,N_10666);
nand U14480 (N_14480,N_11394,N_12194);
or U14481 (N_14481,N_11830,N_11586);
and U14482 (N_14482,N_10380,N_12151);
nor U14483 (N_14483,N_12116,N_10054);
nand U14484 (N_14484,N_12273,N_11390);
nor U14485 (N_14485,N_11244,N_11433);
or U14486 (N_14486,N_11807,N_10640);
nor U14487 (N_14487,N_10836,N_10785);
or U14488 (N_14488,N_11540,N_11584);
and U14489 (N_14489,N_12260,N_11179);
nor U14490 (N_14490,N_10485,N_11648);
or U14491 (N_14491,N_12461,N_10123);
or U14492 (N_14492,N_10196,N_10238);
or U14493 (N_14493,N_10698,N_10199);
nor U14494 (N_14494,N_11872,N_12004);
nor U14495 (N_14495,N_10278,N_12307);
or U14496 (N_14496,N_10558,N_10577);
nor U14497 (N_14497,N_10135,N_10578);
or U14498 (N_14498,N_10789,N_11058);
and U14499 (N_14499,N_11060,N_11668);
xor U14500 (N_14500,N_11172,N_12335);
and U14501 (N_14501,N_11366,N_10660);
nand U14502 (N_14502,N_10739,N_10559);
nor U14503 (N_14503,N_11417,N_11882);
or U14504 (N_14504,N_11486,N_12138);
nand U14505 (N_14505,N_10742,N_10120);
nor U14506 (N_14506,N_10117,N_10082);
nor U14507 (N_14507,N_12311,N_12411);
nor U14508 (N_14508,N_10684,N_10600);
nor U14509 (N_14509,N_11739,N_11268);
and U14510 (N_14510,N_11247,N_10019);
and U14511 (N_14511,N_10276,N_12224);
nand U14512 (N_14512,N_10660,N_10530);
or U14513 (N_14513,N_11694,N_11586);
and U14514 (N_14514,N_10044,N_10234);
nor U14515 (N_14515,N_10125,N_10311);
and U14516 (N_14516,N_12152,N_12374);
xnor U14517 (N_14517,N_11720,N_10360);
or U14518 (N_14518,N_12441,N_11036);
and U14519 (N_14519,N_11376,N_10201);
nand U14520 (N_14520,N_10523,N_10999);
and U14521 (N_14521,N_11267,N_11224);
nand U14522 (N_14522,N_10232,N_11048);
and U14523 (N_14523,N_11950,N_11603);
or U14524 (N_14524,N_11030,N_10827);
nand U14525 (N_14525,N_10473,N_10240);
nand U14526 (N_14526,N_11718,N_11286);
or U14527 (N_14527,N_10921,N_11483);
and U14528 (N_14528,N_12230,N_12074);
nor U14529 (N_14529,N_10895,N_11938);
nor U14530 (N_14530,N_12345,N_10651);
or U14531 (N_14531,N_12082,N_11672);
and U14532 (N_14532,N_11037,N_10410);
nor U14533 (N_14533,N_10545,N_11802);
nand U14534 (N_14534,N_11896,N_11012);
nand U14535 (N_14535,N_12164,N_11197);
nor U14536 (N_14536,N_10335,N_12145);
or U14537 (N_14537,N_11493,N_11554);
or U14538 (N_14538,N_11396,N_11807);
nor U14539 (N_14539,N_11367,N_11413);
nor U14540 (N_14540,N_10715,N_10474);
or U14541 (N_14541,N_12431,N_12009);
nor U14542 (N_14542,N_10549,N_12086);
nand U14543 (N_14543,N_11240,N_11799);
or U14544 (N_14544,N_10439,N_11583);
and U14545 (N_14545,N_11843,N_11930);
and U14546 (N_14546,N_10799,N_10851);
and U14547 (N_14547,N_10366,N_10183);
or U14548 (N_14548,N_11064,N_10875);
and U14549 (N_14549,N_12159,N_11554);
nand U14550 (N_14550,N_11547,N_10934);
nor U14551 (N_14551,N_11491,N_10647);
nor U14552 (N_14552,N_11718,N_11651);
and U14553 (N_14553,N_12234,N_11587);
nand U14554 (N_14554,N_11341,N_12265);
nand U14555 (N_14555,N_11781,N_11204);
or U14556 (N_14556,N_11739,N_10580);
or U14557 (N_14557,N_11474,N_10402);
nor U14558 (N_14558,N_11408,N_10627);
or U14559 (N_14559,N_12216,N_10435);
or U14560 (N_14560,N_11159,N_12261);
and U14561 (N_14561,N_12059,N_10981);
xnor U14562 (N_14562,N_10844,N_11893);
nand U14563 (N_14563,N_11810,N_10477);
nand U14564 (N_14564,N_12254,N_11389);
nor U14565 (N_14565,N_11058,N_10854);
nand U14566 (N_14566,N_10891,N_12427);
and U14567 (N_14567,N_12163,N_11370);
nor U14568 (N_14568,N_12283,N_12248);
nand U14569 (N_14569,N_12391,N_12227);
or U14570 (N_14570,N_10533,N_12441);
and U14571 (N_14571,N_11209,N_11330);
nor U14572 (N_14572,N_10312,N_10365);
or U14573 (N_14573,N_12239,N_12361);
or U14574 (N_14574,N_12210,N_10786);
and U14575 (N_14575,N_11556,N_10717);
nand U14576 (N_14576,N_10854,N_10603);
or U14577 (N_14577,N_11738,N_11007);
xor U14578 (N_14578,N_12081,N_10637);
nor U14579 (N_14579,N_11190,N_10275);
nand U14580 (N_14580,N_11766,N_11015);
or U14581 (N_14581,N_11090,N_10898);
nand U14582 (N_14582,N_11615,N_11356);
and U14583 (N_14583,N_11243,N_10641);
nor U14584 (N_14584,N_11839,N_11398);
and U14585 (N_14585,N_12484,N_12173);
and U14586 (N_14586,N_11553,N_10576);
nand U14587 (N_14587,N_10719,N_11391);
and U14588 (N_14588,N_10773,N_10338);
nand U14589 (N_14589,N_12191,N_10631);
or U14590 (N_14590,N_10007,N_11599);
or U14591 (N_14591,N_12226,N_11544);
or U14592 (N_14592,N_10855,N_11351);
nand U14593 (N_14593,N_10473,N_10008);
nor U14594 (N_14594,N_12145,N_10709);
and U14595 (N_14595,N_11052,N_11188);
and U14596 (N_14596,N_11357,N_12321);
nor U14597 (N_14597,N_12243,N_11327);
and U14598 (N_14598,N_11088,N_11179);
nand U14599 (N_14599,N_11299,N_12493);
nand U14600 (N_14600,N_10291,N_10455);
nor U14601 (N_14601,N_10797,N_11464);
nor U14602 (N_14602,N_10605,N_12453);
and U14603 (N_14603,N_11846,N_10104);
nand U14604 (N_14604,N_10466,N_11615);
nor U14605 (N_14605,N_11969,N_10383);
nand U14606 (N_14606,N_10281,N_10377);
or U14607 (N_14607,N_10624,N_12366);
nor U14608 (N_14608,N_10200,N_12240);
or U14609 (N_14609,N_11648,N_11241);
nor U14610 (N_14610,N_11338,N_12220);
nor U14611 (N_14611,N_10440,N_10568);
nor U14612 (N_14612,N_11333,N_10278);
nand U14613 (N_14613,N_10879,N_11409);
or U14614 (N_14614,N_11549,N_12316);
and U14615 (N_14615,N_11635,N_11230);
and U14616 (N_14616,N_11152,N_11303);
nor U14617 (N_14617,N_11063,N_11986);
nor U14618 (N_14618,N_10385,N_12356);
nand U14619 (N_14619,N_10756,N_10650);
nor U14620 (N_14620,N_11138,N_12458);
or U14621 (N_14621,N_12120,N_10888);
nor U14622 (N_14622,N_11615,N_10346);
and U14623 (N_14623,N_12120,N_10014);
and U14624 (N_14624,N_10161,N_11423);
and U14625 (N_14625,N_10634,N_10744);
or U14626 (N_14626,N_11052,N_11903);
nor U14627 (N_14627,N_10252,N_10508);
xnor U14628 (N_14628,N_10342,N_12459);
and U14629 (N_14629,N_12252,N_12320);
or U14630 (N_14630,N_12189,N_11130);
or U14631 (N_14631,N_11534,N_11152);
and U14632 (N_14632,N_10243,N_10086);
nand U14633 (N_14633,N_11299,N_12469);
nand U14634 (N_14634,N_11039,N_11638);
nor U14635 (N_14635,N_11316,N_10890);
or U14636 (N_14636,N_11174,N_12373);
or U14637 (N_14637,N_11005,N_11202);
nor U14638 (N_14638,N_11863,N_11992);
and U14639 (N_14639,N_10531,N_10092);
nand U14640 (N_14640,N_11559,N_11530);
nor U14641 (N_14641,N_11598,N_11430);
nor U14642 (N_14642,N_11504,N_11372);
nand U14643 (N_14643,N_10448,N_11418);
nand U14644 (N_14644,N_11334,N_11513);
or U14645 (N_14645,N_10215,N_11536);
or U14646 (N_14646,N_11346,N_12462);
nor U14647 (N_14647,N_10252,N_10957);
nand U14648 (N_14648,N_10491,N_10485);
nand U14649 (N_14649,N_12382,N_11135);
nor U14650 (N_14650,N_11142,N_11073);
nor U14651 (N_14651,N_10633,N_11892);
and U14652 (N_14652,N_11920,N_10949);
nand U14653 (N_14653,N_10009,N_10123);
and U14654 (N_14654,N_11857,N_10701);
nor U14655 (N_14655,N_10030,N_10209);
or U14656 (N_14656,N_10503,N_11832);
and U14657 (N_14657,N_10381,N_12154);
and U14658 (N_14658,N_10391,N_12016);
and U14659 (N_14659,N_10175,N_12192);
nand U14660 (N_14660,N_12475,N_12264);
and U14661 (N_14661,N_10983,N_11688);
nor U14662 (N_14662,N_12380,N_10925);
nand U14663 (N_14663,N_10326,N_10898);
nand U14664 (N_14664,N_12021,N_10662);
and U14665 (N_14665,N_10315,N_11569);
or U14666 (N_14666,N_11046,N_10704);
and U14667 (N_14667,N_10700,N_10385);
nor U14668 (N_14668,N_10366,N_10642);
and U14669 (N_14669,N_11933,N_10860);
nor U14670 (N_14670,N_12165,N_11063);
and U14671 (N_14671,N_12311,N_10411);
nor U14672 (N_14672,N_10018,N_11920);
nor U14673 (N_14673,N_11064,N_12401);
nand U14674 (N_14674,N_11471,N_11229);
or U14675 (N_14675,N_10526,N_11697);
nor U14676 (N_14676,N_10337,N_11524);
or U14677 (N_14677,N_10381,N_10605);
nor U14678 (N_14678,N_11817,N_11639);
and U14679 (N_14679,N_10693,N_11508);
and U14680 (N_14680,N_11821,N_11607);
and U14681 (N_14681,N_11248,N_12296);
nor U14682 (N_14682,N_11896,N_12100);
nor U14683 (N_14683,N_11139,N_10050);
and U14684 (N_14684,N_10411,N_12187);
xnor U14685 (N_14685,N_10572,N_10343);
nand U14686 (N_14686,N_10959,N_10095);
and U14687 (N_14687,N_10400,N_11529);
nand U14688 (N_14688,N_10227,N_11378);
nor U14689 (N_14689,N_10512,N_11306);
nand U14690 (N_14690,N_11870,N_12002);
or U14691 (N_14691,N_11552,N_11975);
and U14692 (N_14692,N_12015,N_11708);
nand U14693 (N_14693,N_11035,N_12477);
nand U14694 (N_14694,N_10165,N_12357);
xor U14695 (N_14695,N_12087,N_12308);
nor U14696 (N_14696,N_11950,N_12234);
nand U14697 (N_14697,N_10090,N_11780);
nor U14698 (N_14698,N_11027,N_10319);
and U14699 (N_14699,N_11790,N_11419);
nand U14700 (N_14700,N_12277,N_12339);
or U14701 (N_14701,N_11006,N_10624);
nand U14702 (N_14702,N_11923,N_11527);
nor U14703 (N_14703,N_10255,N_10792);
xor U14704 (N_14704,N_10760,N_11261);
and U14705 (N_14705,N_11580,N_11682);
nand U14706 (N_14706,N_10734,N_11762);
nor U14707 (N_14707,N_10871,N_11478);
or U14708 (N_14708,N_11625,N_11925);
and U14709 (N_14709,N_10003,N_11334);
and U14710 (N_14710,N_11192,N_11495);
nor U14711 (N_14711,N_10371,N_11174);
nand U14712 (N_14712,N_10255,N_11290);
nor U14713 (N_14713,N_11389,N_11139);
or U14714 (N_14714,N_10810,N_11016);
nor U14715 (N_14715,N_12182,N_11196);
nand U14716 (N_14716,N_11662,N_12496);
nor U14717 (N_14717,N_11294,N_12116);
nor U14718 (N_14718,N_11727,N_10464);
or U14719 (N_14719,N_11859,N_11847);
nand U14720 (N_14720,N_10279,N_11087);
nand U14721 (N_14721,N_10533,N_11872);
nand U14722 (N_14722,N_10953,N_11687);
nand U14723 (N_14723,N_12423,N_11161);
and U14724 (N_14724,N_11343,N_11481);
or U14725 (N_14725,N_10974,N_11236);
or U14726 (N_14726,N_11712,N_10317);
nand U14727 (N_14727,N_11616,N_10410);
nor U14728 (N_14728,N_11076,N_11934);
nor U14729 (N_14729,N_11894,N_10153);
or U14730 (N_14730,N_12376,N_10633);
nor U14731 (N_14731,N_11154,N_12213);
nand U14732 (N_14732,N_10948,N_10660);
nand U14733 (N_14733,N_11536,N_10835);
and U14734 (N_14734,N_11568,N_11950);
nand U14735 (N_14735,N_12343,N_12266);
nand U14736 (N_14736,N_10075,N_12230);
nand U14737 (N_14737,N_10268,N_11098);
nor U14738 (N_14738,N_11625,N_12157);
or U14739 (N_14739,N_10467,N_12268);
nor U14740 (N_14740,N_11535,N_10223);
xor U14741 (N_14741,N_11597,N_10369);
nand U14742 (N_14742,N_12491,N_12052);
or U14743 (N_14743,N_11223,N_12321);
nor U14744 (N_14744,N_10369,N_11829);
or U14745 (N_14745,N_12163,N_10711);
nor U14746 (N_14746,N_12488,N_11351);
nor U14747 (N_14747,N_11224,N_10411);
nand U14748 (N_14748,N_12313,N_10812);
nand U14749 (N_14749,N_10316,N_10970);
and U14750 (N_14750,N_10267,N_10849);
or U14751 (N_14751,N_11607,N_11744);
or U14752 (N_14752,N_12054,N_10044);
and U14753 (N_14753,N_12316,N_11872);
nand U14754 (N_14754,N_11038,N_10992);
or U14755 (N_14755,N_12177,N_10685);
nand U14756 (N_14756,N_12366,N_11578);
and U14757 (N_14757,N_12062,N_11344);
and U14758 (N_14758,N_10845,N_11403);
and U14759 (N_14759,N_12192,N_10664);
nor U14760 (N_14760,N_10440,N_11487);
nor U14761 (N_14761,N_11853,N_10590);
or U14762 (N_14762,N_11821,N_12166);
nand U14763 (N_14763,N_11122,N_12067);
nor U14764 (N_14764,N_12155,N_11620);
and U14765 (N_14765,N_12020,N_11028);
nand U14766 (N_14766,N_10709,N_10048);
nand U14767 (N_14767,N_11790,N_11432);
or U14768 (N_14768,N_10707,N_10378);
nand U14769 (N_14769,N_10157,N_10602);
nand U14770 (N_14770,N_10828,N_11438);
nor U14771 (N_14771,N_11962,N_10098);
and U14772 (N_14772,N_12325,N_12285);
and U14773 (N_14773,N_10699,N_10133);
nand U14774 (N_14774,N_11852,N_12403);
and U14775 (N_14775,N_12356,N_12260);
or U14776 (N_14776,N_11547,N_11495);
xnor U14777 (N_14777,N_11073,N_11736);
nor U14778 (N_14778,N_11352,N_11509);
and U14779 (N_14779,N_10437,N_10284);
nor U14780 (N_14780,N_11733,N_10198);
nand U14781 (N_14781,N_11091,N_10921);
nor U14782 (N_14782,N_11346,N_12096);
nor U14783 (N_14783,N_10279,N_12219);
and U14784 (N_14784,N_12416,N_10322);
or U14785 (N_14785,N_11370,N_11085);
nor U14786 (N_14786,N_11284,N_12205);
nand U14787 (N_14787,N_10676,N_11492);
nor U14788 (N_14788,N_12048,N_10385);
and U14789 (N_14789,N_11003,N_11733);
nand U14790 (N_14790,N_10362,N_11342);
nand U14791 (N_14791,N_12398,N_11862);
nor U14792 (N_14792,N_10732,N_12490);
and U14793 (N_14793,N_11717,N_10733);
and U14794 (N_14794,N_12205,N_11575);
or U14795 (N_14795,N_12032,N_10236);
xnor U14796 (N_14796,N_11143,N_12107);
and U14797 (N_14797,N_10998,N_11406);
and U14798 (N_14798,N_11366,N_10287);
and U14799 (N_14799,N_12403,N_11466);
nand U14800 (N_14800,N_12104,N_11633);
nand U14801 (N_14801,N_12133,N_11704);
or U14802 (N_14802,N_10694,N_10553);
and U14803 (N_14803,N_11874,N_10180);
or U14804 (N_14804,N_10603,N_12367);
or U14805 (N_14805,N_10560,N_11125);
or U14806 (N_14806,N_11855,N_12320);
or U14807 (N_14807,N_12190,N_11603);
nor U14808 (N_14808,N_12326,N_11821);
or U14809 (N_14809,N_10477,N_11203);
and U14810 (N_14810,N_12267,N_11717);
and U14811 (N_14811,N_10752,N_12457);
nand U14812 (N_14812,N_11016,N_11450);
and U14813 (N_14813,N_12423,N_10739);
or U14814 (N_14814,N_11027,N_10618);
or U14815 (N_14815,N_11931,N_10043);
or U14816 (N_14816,N_10192,N_12105);
or U14817 (N_14817,N_11748,N_12234);
nand U14818 (N_14818,N_10768,N_12246);
nor U14819 (N_14819,N_11726,N_10273);
and U14820 (N_14820,N_12019,N_12374);
nor U14821 (N_14821,N_12310,N_10875);
or U14822 (N_14822,N_11514,N_11527);
nand U14823 (N_14823,N_11613,N_12351);
nand U14824 (N_14824,N_11002,N_11565);
or U14825 (N_14825,N_10297,N_12457);
nand U14826 (N_14826,N_11441,N_10856);
or U14827 (N_14827,N_10814,N_10848);
and U14828 (N_14828,N_10130,N_10795);
or U14829 (N_14829,N_11241,N_11129);
xor U14830 (N_14830,N_10028,N_10418);
nor U14831 (N_14831,N_11784,N_10865);
nor U14832 (N_14832,N_12264,N_11604);
or U14833 (N_14833,N_10361,N_10108);
nand U14834 (N_14834,N_10957,N_11354);
nor U14835 (N_14835,N_11407,N_11527);
nor U14836 (N_14836,N_11103,N_10901);
nor U14837 (N_14837,N_10334,N_10408);
and U14838 (N_14838,N_11439,N_10110);
nor U14839 (N_14839,N_11086,N_11441);
nor U14840 (N_14840,N_11965,N_10916);
nor U14841 (N_14841,N_11370,N_11333);
and U14842 (N_14842,N_11074,N_11495);
nand U14843 (N_14843,N_12491,N_10778);
and U14844 (N_14844,N_10127,N_11172);
or U14845 (N_14845,N_12423,N_11543);
or U14846 (N_14846,N_11419,N_11254);
and U14847 (N_14847,N_10289,N_11406);
and U14848 (N_14848,N_10710,N_12305);
nand U14849 (N_14849,N_11013,N_11772);
or U14850 (N_14850,N_12045,N_10850);
or U14851 (N_14851,N_10795,N_11532);
nor U14852 (N_14852,N_11600,N_10659);
or U14853 (N_14853,N_11660,N_11053);
nor U14854 (N_14854,N_10647,N_11680);
nand U14855 (N_14855,N_10895,N_10754);
nor U14856 (N_14856,N_11219,N_12020);
nand U14857 (N_14857,N_10301,N_11587);
or U14858 (N_14858,N_12311,N_11488);
or U14859 (N_14859,N_12030,N_11219);
and U14860 (N_14860,N_10870,N_11747);
nor U14861 (N_14861,N_12189,N_11541);
and U14862 (N_14862,N_12308,N_12442);
or U14863 (N_14863,N_11309,N_10998);
nor U14864 (N_14864,N_12134,N_10422);
nor U14865 (N_14865,N_11890,N_11493);
and U14866 (N_14866,N_10937,N_10805);
and U14867 (N_14867,N_10808,N_10550);
nor U14868 (N_14868,N_11067,N_11261);
nand U14869 (N_14869,N_11987,N_10100);
nand U14870 (N_14870,N_12237,N_10464);
nand U14871 (N_14871,N_10768,N_10823);
or U14872 (N_14872,N_11515,N_12459);
nor U14873 (N_14873,N_12459,N_10194);
nor U14874 (N_14874,N_12470,N_11123);
and U14875 (N_14875,N_10666,N_11404);
and U14876 (N_14876,N_10286,N_11036);
or U14877 (N_14877,N_11932,N_10506);
or U14878 (N_14878,N_11775,N_12040);
nor U14879 (N_14879,N_11893,N_10113);
and U14880 (N_14880,N_10465,N_11542);
and U14881 (N_14881,N_11802,N_11774);
and U14882 (N_14882,N_10850,N_11324);
nor U14883 (N_14883,N_10067,N_12085);
nand U14884 (N_14884,N_10409,N_11968);
nand U14885 (N_14885,N_11918,N_11490);
nor U14886 (N_14886,N_10362,N_10255);
or U14887 (N_14887,N_12224,N_11698);
nand U14888 (N_14888,N_10198,N_12240);
xor U14889 (N_14889,N_10291,N_11262);
nand U14890 (N_14890,N_10022,N_12218);
nand U14891 (N_14891,N_11965,N_10355);
and U14892 (N_14892,N_11611,N_11572);
or U14893 (N_14893,N_10714,N_12405);
nand U14894 (N_14894,N_11114,N_11966);
and U14895 (N_14895,N_11253,N_10424);
or U14896 (N_14896,N_11469,N_10869);
nor U14897 (N_14897,N_10001,N_11776);
nand U14898 (N_14898,N_12287,N_10829);
and U14899 (N_14899,N_11436,N_12116);
and U14900 (N_14900,N_10114,N_10582);
nand U14901 (N_14901,N_10843,N_12257);
nand U14902 (N_14902,N_11217,N_12433);
nor U14903 (N_14903,N_12229,N_11825);
and U14904 (N_14904,N_11865,N_10677);
nand U14905 (N_14905,N_11959,N_10184);
nor U14906 (N_14906,N_11124,N_10522);
nand U14907 (N_14907,N_10433,N_11453);
nand U14908 (N_14908,N_12126,N_12024);
nor U14909 (N_14909,N_10604,N_12337);
nand U14910 (N_14910,N_10654,N_12242);
nand U14911 (N_14911,N_11040,N_10674);
nor U14912 (N_14912,N_10102,N_11175);
nor U14913 (N_14913,N_10466,N_11968);
and U14914 (N_14914,N_12017,N_11949);
nand U14915 (N_14915,N_11343,N_10438);
and U14916 (N_14916,N_12128,N_10165);
and U14917 (N_14917,N_12496,N_10132);
and U14918 (N_14918,N_11185,N_10657);
nor U14919 (N_14919,N_10482,N_10079);
or U14920 (N_14920,N_10132,N_10409);
nand U14921 (N_14921,N_11611,N_11170);
or U14922 (N_14922,N_12165,N_11749);
nand U14923 (N_14923,N_11841,N_12159);
nand U14924 (N_14924,N_11581,N_12067);
and U14925 (N_14925,N_10446,N_10846);
or U14926 (N_14926,N_11423,N_11242);
nor U14927 (N_14927,N_11235,N_12340);
nor U14928 (N_14928,N_11419,N_12291);
nor U14929 (N_14929,N_11439,N_12351);
or U14930 (N_14930,N_11330,N_11351);
or U14931 (N_14931,N_11356,N_11149);
nand U14932 (N_14932,N_11563,N_11529);
or U14933 (N_14933,N_10270,N_11198);
nand U14934 (N_14934,N_12452,N_10380);
nand U14935 (N_14935,N_11076,N_11155);
nor U14936 (N_14936,N_10206,N_11443);
or U14937 (N_14937,N_11720,N_11232);
or U14938 (N_14938,N_10762,N_10356);
nand U14939 (N_14939,N_11726,N_11067);
and U14940 (N_14940,N_11594,N_10171);
or U14941 (N_14941,N_10580,N_11913);
or U14942 (N_14942,N_10928,N_11587);
nor U14943 (N_14943,N_12415,N_12322);
and U14944 (N_14944,N_11783,N_12388);
nor U14945 (N_14945,N_11907,N_10849);
and U14946 (N_14946,N_10827,N_10331);
nand U14947 (N_14947,N_10786,N_11149);
nand U14948 (N_14948,N_10641,N_11084);
and U14949 (N_14949,N_11697,N_10516);
or U14950 (N_14950,N_11561,N_11194);
or U14951 (N_14951,N_12078,N_10282);
nand U14952 (N_14952,N_10646,N_11397);
or U14953 (N_14953,N_12102,N_11897);
nand U14954 (N_14954,N_10440,N_10187);
and U14955 (N_14955,N_10956,N_11715);
or U14956 (N_14956,N_10000,N_10227);
nor U14957 (N_14957,N_12047,N_10537);
and U14958 (N_14958,N_11619,N_10480);
nor U14959 (N_14959,N_11722,N_10022);
or U14960 (N_14960,N_11827,N_11634);
nor U14961 (N_14961,N_10145,N_10108);
nor U14962 (N_14962,N_11499,N_11755);
nor U14963 (N_14963,N_12161,N_11812);
and U14964 (N_14964,N_10704,N_11878);
nand U14965 (N_14965,N_11053,N_11826);
nor U14966 (N_14966,N_12403,N_12397);
nand U14967 (N_14967,N_10572,N_11578);
nor U14968 (N_14968,N_11226,N_10239);
or U14969 (N_14969,N_10011,N_12103);
and U14970 (N_14970,N_11085,N_11967);
or U14971 (N_14971,N_11313,N_11578);
nand U14972 (N_14972,N_11774,N_11092);
and U14973 (N_14973,N_11641,N_11940);
nand U14974 (N_14974,N_12409,N_11836);
xor U14975 (N_14975,N_11477,N_10112);
or U14976 (N_14976,N_10287,N_12157);
and U14977 (N_14977,N_12273,N_11863);
and U14978 (N_14978,N_10202,N_11139);
and U14979 (N_14979,N_10824,N_12051);
or U14980 (N_14980,N_11269,N_10321);
or U14981 (N_14981,N_11532,N_10924);
nor U14982 (N_14982,N_12352,N_10195);
nor U14983 (N_14983,N_12428,N_10296);
or U14984 (N_14984,N_10803,N_11835);
nor U14985 (N_14985,N_10770,N_11392);
or U14986 (N_14986,N_10303,N_10353);
nand U14987 (N_14987,N_11127,N_11104);
or U14988 (N_14988,N_10261,N_11174);
and U14989 (N_14989,N_12223,N_10096);
and U14990 (N_14990,N_12252,N_10177);
nand U14991 (N_14991,N_10524,N_11839);
nor U14992 (N_14992,N_11488,N_11506);
or U14993 (N_14993,N_12012,N_11279);
nand U14994 (N_14994,N_12016,N_10088);
or U14995 (N_14995,N_12164,N_12460);
and U14996 (N_14996,N_11335,N_10213);
and U14997 (N_14997,N_10250,N_10655);
nor U14998 (N_14998,N_10352,N_10161);
nand U14999 (N_14999,N_11768,N_11067);
and U15000 (N_15000,N_13254,N_14140);
or U15001 (N_15001,N_12532,N_13459);
nor U15002 (N_15002,N_13187,N_14629);
nand U15003 (N_15003,N_14390,N_14931);
and U15004 (N_15004,N_14979,N_14290);
or U15005 (N_15005,N_13753,N_14442);
and U15006 (N_15006,N_12860,N_13184);
and U15007 (N_15007,N_13932,N_14714);
xor U15008 (N_15008,N_13587,N_14652);
and U15009 (N_15009,N_14309,N_13629);
nand U15010 (N_15010,N_13831,N_14493);
and U15011 (N_15011,N_12562,N_14919);
and U15012 (N_15012,N_14000,N_12872);
or U15013 (N_15013,N_12653,N_14159);
or U15014 (N_15014,N_12730,N_12985);
nand U15015 (N_15015,N_14544,N_13675);
and U15016 (N_15016,N_13097,N_13899);
or U15017 (N_15017,N_14437,N_13827);
and U15018 (N_15018,N_14752,N_12571);
and U15019 (N_15019,N_13394,N_14877);
or U15020 (N_15020,N_14021,N_14126);
and U15021 (N_15021,N_13940,N_14732);
nand U15022 (N_15022,N_14529,N_13712);
and U15023 (N_15023,N_14247,N_12839);
nand U15024 (N_15024,N_14808,N_13944);
nand U15025 (N_15025,N_14993,N_14900);
and U15026 (N_15026,N_13590,N_12752);
nand U15027 (N_15027,N_13724,N_13444);
nor U15028 (N_15028,N_14851,N_14588);
or U15029 (N_15029,N_13664,N_13242);
nor U15030 (N_15030,N_14013,N_14199);
or U15031 (N_15031,N_12593,N_14858);
nor U15032 (N_15032,N_12501,N_13741);
or U15033 (N_15033,N_14826,N_14232);
and U15034 (N_15034,N_14091,N_14246);
nor U15035 (N_15035,N_13967,N_14139);
or U15036 (N_15036,N_12699,N_13199);
or U15037 (N_15037,N_14121,N_12785);
or U15038 (N_15038,N_13466,N_13418);
nor U15039 (N_15039,N_14372,N_12568);
or U15040 (N_15040,N_14947,N_13258);
or U15041 (N_15041,N_12645,N_14878);
and U15042 (N_15042,N_13045,N_13739);
nor U15043 (N_15043,N_14743,N_13111);
nor U15044 (N_15044,N_14517,N_14870);
xnor U15045 (N_15045,N_14884,N_12605);
and U15046 (N_15046,N_14347,N_14936);
nor U15047 (N_15047,N_13439,N_14830);
nor U15048 (N_15048,N_14114,N_12831);
nand U15049 (N_15049,N_13130,N_14671);
nand U15050 (N_15050,N_13088,N_14319);
nand U15051 (N_15051,N_14036,N_13002);
nor U15052 (N_15052,N_14577,N_12707);
nand U15053 (N_15053,N_13680,N_12865);
nor U15054 (N_15054,N_14105,N_12959);
nor U15055 (N_15055,N_14343,N_14145);
nor U15056 (N_15056,N_12914,N_14181);
or U15057 (N_15057,N_14917,N_14736);
and U15058 (N_15058,N_14062,N_13257);
and U15059 (N_15059,N_13970,N_12517);
and U15060 (N_15060,N_12512,N_14429);
nor U15061 (N_15061,N_13244,N_14642);
nor U15062 (N_15062,N_14408,N_13938);
and U15063 (N_15063,N_12869,N_13329);
or U15064 (N_15064,N_13151,N_14829);
nand U15065 (N_15065,N_14607,N_12725);
or U15066 (N_15066,N_13089,N_12680);
and U15067 (N_15067,N_13843,N_12989);
nand U15068 (N_15068,N_14983,N_13505);
nand U15069 (N_15069,N_13272,N_13732);
nand U15070 (N_15070,N_14700,N_14797);
or U15071 (N_15071,N_14565,N_14701);
nand U15072 (N_15072,N_12846,N_13772);
or U15073 (N_15073,N_13322,N_13348);
nor U15074 (N_15074,N_12650,N_13145);
nand U15075 (N_15075,N_14560,N_13536);
nor U15076 (N_15076,N_13457,N_14321);
or U15077 (N_15077,N_14217,N_14951);
nand U15078 (N_15078,N_12669,N_14253);
nor U15079 (N_15079,N_14401,N_14001);
nor U15080 (N_15080,N_12954,N_13610);
and U15081 (N_15081,N_12743,N_13583);
nand U15082 (N_15082,N_13478,N_13033);
nor U15083 (N_15083,N_12889,N_14399);
and U15084 (N_15084,N_13029,N_14019);
or U15085 (N_15085,N_13341,N_14859);
nand U15086 (N_15086,N_13204,N_14035);
nor U15087 (N_15087,N_12878,N_12681);
nand U15088 (N_15088,N_13174,N_13308);
or U15089 (N_15089,N_13708,N_13992);
nand U15090 (N_15090,N_13074,N_14890);
and U15091 (N_15091,N_12587,N_13818);
nor U15092 (N_15092,N_14778,N_13851);
nand U15093 (N_15093,N_12996,N_13847);
nand U15094 (N_15094,N_14152,N_14513);
nor U15095 (N_15095,N_13364,N_14194);
nand U15096 (N_15096,N_14627,N_14078);
nand U15097 (N_15097,N_14967,N_13054);
nand U15098 (N_15098,N_12871,N_12777);
nor U15099 (N_15099,N_13490,N_14481);
or U15100 (N_15100,N_13568,N_13744);
nand U15101 (N_15101,N_12746,N_13201);
and U15102 (N_15102,N_14280,N_12736);
nand U15103 (N_15103,N_12897,N_13621);
nor U15104 (N_15104,N_12599,N_13372);
nand U15105 (N_15105,N_13396,N_12504);
nor U15106 (N_15106,N_12634,N_14382);
nand U15107 (N_15107,N_12659,N_14193);
or U15108 (N_15108,N_14227,N_13259);
or U15109 (N_15109,N_12670,N_13848);
and U15110 (N_15110,N_14759,N_14075);
or U15111 (N_15111,N_13353,N_13981);
nand U15112 (N_15112,N_13278,N_13090);
and U15113 (N_15113,N_14596,N_14862);
nand U15114 (N_15114,N_13662,N_14080);
and U15115 (N_15115,N_13585,N_14601);
or U15116 (N_15116,N_14123,N_13541);
nor U15117 (N_15117,N_13248,N_13942);
or U15118 (N_15118,N_13286,N_13876);
nand U15119 (N_15119,N_14383,N_12993);
or U15120 (N_15120,N_14089,N_13865);
nor U15121 (N_15121,N_14605,N_14179);
nand U15122 (N_15122,N_14471,N_13246);
and U15123 (N_15123,N_13344,N_14675);
and U15124 (N_15124,N_14052,N_14317);
or U15125 (N_15125,N_13626,N_13497);
and U15126 (N_15126,N_13691,N_13704);
nand U15127 (N_15127,N_12738,N_13104);
nand U15128 (N_15128,N_13212,N_13224);
and U15129 (N_15129,N_14106,N_13702);
nand U15130 (N_15130,N_14010,N_12810);
nor U15131 (N_15131,N_14932,N_13220);
or U15132 (N_15132,N_13654,N_14856);
nand U15133 (N_15133,N_13358,N_14248);
or U15134 (N_15134,N_12945,N_14341);
or U15135 (N_15135,N_13953,N_14180);
or U15136 (N_15136,N_13751,N_14874);
or U15137 (N_15137,N_13122,N_14754);
and U15138 (N_15138,N_13207,N_13429);
and U15139 (N_15139,N_14817,N_14772);
nor U15140 (N_15140,N_14130,N_13565);
nand U15141 (N_15141,N_14998,N_14537);
or U15142 (N_15142,N_13208,N_13183);
nor U15143 (N_15143,N_12661,N_13602);
nand U15144 (N_15144,N_13909,N_13113);
nand U15145 (N_15145,N_13126,N_14679);
and U15146 (N_15146,N_13862,N_13376);
nor U15147 (N_15147,N_14503,N_12982);
nor U15148 (N_15148,N_13034,N_14370);
nand U15149 (N_15149,N_14421,N_14452);
or U15150 (N_15150,N_12908,N_14526);
nor U15151 (N_15151,N_13889,N_13345);
or U15152 (N_15152,N_14040,N_13219);
nor U15153 (N_15153,N_14475,N_12665);
nand U15154 (N_15154,N_12980,N_13973);
or U15155 (N_15155,N_14305,N_12566);
and U15156 (N_15156,N_14655,N_12994);
or U15157 (N_15157,N_13530,N_13337);
or U15158 (N_15158,N_12613,N_14992);
nand U15159 (N_15159,N_12692,N_12862);
or U15160 (N_15160,N_14511,N_14834);
and U15161 (N_15161,N_12974,N_14753);
and U15162 (N_15162,N_13488,N_13014);
nor U15163 (N_15163,N_12886,N_14125);
nor U15164 (N_15164,N_14205,N_12523);
nor U15165 (N_15165,N_14359,N_14901);
or U15166 (N_15166,N_13399,N_14231);
nand U15167 (N_15167,N_14470,N_12554);
nor U15168 (N_15168,N_14581,N_13816);
or U15169 (N_15169,N_14320,N_14624);
nor U15170 (N_15170,N_14004,N_13213);
or U15171 (N_15171,N_13920,N_14164);
and U15172 (N_15172,N_13161,N_13579);
nand U15173 (N_15173,N_14924,N_13300);
and U15174 (N_15174,N_12833,N_14096);
and U15175 (N_15175,N_12882,N_13028);
nand U15176 (N_15176,N_14820,N_12911);
and U15177 (N_15177,N_14354,N_14651);
and U15178 (N_15178,N_13716,N_13262);
nor U15179 (N_15179,N_12917,N_14069);
or U15180 (N_15180,N_14413,N_14965);
and U15181 (N_15181,N_13817,N_13471);
nor U15182 (N_15182,N_12899,N_14852);
nor U15183 (N_15183,N_13555,N_12697);
nor U15184 (N_15184,N_12840,N_12711);
or U15185 (N_15185,N_13327,N_14974);
nor U15186 (N_15186,N_14682,N_14095);
nor U15187 (N_15187,N_13863,N_13449);
and U15188 (N_15188,N_12935,N_14240);
or U15189 (N_15189,N_14891,N_14886);
and U15190 (N_15190,N_14045,N_14697);
or U15191 (N_15191,N_12766,N_14433);
nor U15192 (N_15192,N_13401,N_13163);
or U15193 (N_15193,N_14746,N_13160);
nor U15194 (N_15194,N_13634,N_14144);
and U15195 (N_15195,N_14047,N_13321);
nand U15196 (N_15196,N_13050,N_12879);
or U15197 (N_15197,N_14358,N_14079);
and U15198 (N_15198,N_12767,N_12552);
and U15199 (N_15199,N_14518,N_13616);
nand U15200 (N_15200,N_13519,N_14550);
and U15201 (N_15201,N_14060,N_12696);
nand U15202 (N_15202,N_14574,N_14132);
or U15203 (N_15203,N_14249,N_14585);
or U15204 (N_15204,N_13374,N_13234);
and U15205 (N_15205,N_12693,N_14446);
or U15206 (N_15206,N_14773,N_14988);
nand U15207 (N_15207,N_12850,N_13975);
nand U15208 (N_15208,N_13727,N_12544);
nor U15209 (N_15209,N_13378,N_13446);
or U15210 (N_15210,N_13336,N_14533);
or U15211 (N_15211,N_13375,N_12798);
nor U15212 (N_15212,N_14717,N_14610);
nand U15213 (N_15213,N_12758,N_14448);
and U15214 (N_15214,N_13470,N_14122);
and U15215 (N_15215,N_13092,N_14216);
and U15216 (N_15216,N_13983,N_14757);
or U15217 (N_15217,N_12818,N_13604);
or U15218 (N_15218,N_13682,N_12888);
nor U15219 (N_15219,N_14135,N_13767);
or U15220 (N_15220,N_13195,N_12928);
nand U15221 (N_15221,N_12652,N_13011);
and U15222 (N_15222,N_14483,N_14861);
or U15223 (N_15223,N_13804,N_14920);
or U15224 (N_15224,N_13227,N_13454);
or U15225 (N_15225,N_13526,N_14573);
or U15226 (N_15226,N_12960,N_12856);
nand U15227 (N_15227,N_13007,N_14907);
or U15228 (N_15228,N_12944,N_14670);
and U15229 (N_15229,N_14278,N_12976);
and U15230 (N_15230,N_14074,N_12557);
nor U15231 (N_15231,N_14938,N_14895);
nor U15232 (N_15232,N_12760,N_13821);
or U15233 (N_15233,N_12816,N_13858);
and U15234 (N_15234,N_13543,N_13022);
nand U15235 (N_15235,N_13283,N_12970);
and U15236 (N_15236,N_13020,N_14767);
and U15237 (N_15237,N_12870,N_13295);
nand U15238 (N_15238,N_13575,N_13241);
or U15239 (N_15239,N_14669,N_14527);
and U15240 (N_15240,N_14188,N_14602);
nor U15241 (N_15241,N_12967,N_13968);
or U15242 (N_15242,N_14724,N_14785);
nor U15243 (N_15243,N_14349,N_14510);
and U15244 (N_15244,N_13696,N_14620);
nand U15245 (N_15245,N_14257,N_13748);
and U15246 (N_15246,N_12607,N_14136);
nand U15247 (N_15247,N_14559,N_13016);
and U15248 (N_15248,N_13546,N_12648);
nor U15249 (N_15249,N_14944,N_14970);
nand U15250 (N_15250,N_14948,N_13946);
nor U15251 (N_15251,N_13389,N_13733);
and U15252 (N_15252,N_12780,N_14011);
or U15253 (N_15253,N_13124,N_13788);
and U15254 (N_15254,N_12931,N_12761);
nand U15255 (N_15255,N_12988,N_14831);
or U15256 (N_15256,N_12529,N_14594);
nor U15257 (N_15257,N_14222,N_14889);
and U15258 (N_15258,N_13492,N_14101);
nor U15259 (N_15259,N_13841,N_13084);
or U15260 (N_15260,N_14569,N_12705);
nand U15261 (N_15261,N_13082,N_13203);
and U15262 (N_15262,N_14727,N_14532);
nor U15263 (N_15263,N_14688,N_13169);
nand U15264 (N_15264,N_12877,N_14650);
nor U15265 (N_15265,N_13971,N_14049);
nor U15266 (N_15266,N_13655,N_14038);
nand U15267 (N_15267,N_14171,N_14364);
nor U15268 (N_15268,N_12597,N_14281);
nand U15269 (N_15269,N_12809,N_14996);
and U15270 (N_15270,N_13857,N_14561);
nor U15271 (N_15271,N_12811,N_12749);
or U15272 (N_15272,N_14906,N_14668);
nand U15273 (N_15273,N_14638,N_12875);
nor U15274 (N_15274,N_13026,N_13943);
nor U15275 (N_15275,N_13917,N_13365);
nand U15276 (N_15276,N_14915,N_13989);
and U15277 (N_15277,N_13578,N_12732);
nand U15278 (N_15278,N_13522,N_13040);
nor U15279 (N_15279,N_13310,N_13738);
nand U15280 (N_15280,N_13003,N_14064);
or U15281 (N_15281,N_14183,N_12937);
nor U15282 (N_15282,N_14275,N_12550);
nand U15283 (N_15283,N_13021,N_14213);
nand U15284 (N_15284,N_14326,N_14362);
nand U15285 (N_15285,N_13529,N_14392);
and U15286 (N_15286,N_14952,N_14003);
nand U15287 (N_15287,N_13162,N_14684);
and U15288 (N_15288,N_14720,N_14903);
nand U15289 (N_15289,N_14905,N_14755);
and U15290 (N_15290,N_14960,N_12995);
nand U15291 (N_15291,N_13980,N_12703);
nand U15292 (N_15292,N_13379,N_14299);
and U15293 (N_15293,N_14498,N_13233);
nand U15294 (N_15294,N_13605,N_14735);
and U15295 (N_15295,N_13066,N_13468);
nand U15296 (N_15296,N_13722,N_13041);
nor U15297 (N_15297,N_14792,N_13377);
and U15298 (N_15298,N_14657,N_13994);
nand U15299 (N_15299,N_12756,N_12903);
and U15300 (N_15300,N_12644,N_12943);
nand U15301 (N_15301,N_14490,N_13370);
and U15302 (N_15302,N_14150,N_14315);
nor U15303 (N_15303,N_12519,N_14053);
nand U15304 (N_15304,N_13701,N_13839);
or U15305 (N_15305,N_12987,N_14634);
nand U15306 (N_15306,N_13990,N_14378);
nor U15307 (N_15307,N_13229,N_14625);
xnor U15308 (N_15308,N_13690,N_12812);
nor U15309 (N_15309,N_12606,N_14107);
or U15310 (N_15310,N_13672,N_13812);
and U15311 (N_15311,N_14953,N_14980);
nand U15312 (N_15312,N_14568,N_13633);
and U15313 (N_15313,N_14048,N_14268);
or U15314 (N_15314,N_14954,N_13436);
or U15315 (N_15315,N_14853,N_13914);
xor U15316 (N_15316,N_13349,N_13385);
nand U15317 (N_15317,N_14595,N_13540);
or U15318 (N_15318,N_13661,N_13271);
and U15319 (N_15319,N_13746,N_14474);
nand U15320 (N_15320,N_12867,N_14530);
or U15321 (N_15321,N_13576,N_14263);
nor U15322 (N_15322,N_13637,N_13235);
nand U15323 (N_15323,N_12969,N_12841);
nand U15324 (N_15324,N_14881,N_13673);
or U15325 (N_15325,N_14043,N_13534);
and U15326 (N_15326,N_14578,N_14643);
or U15327 (N_15327,N_12941,N_12984);
or U15328 (N_15328,N_13031,N_14946);
and U15329 (N_15329,N_14266,N_13928);
and U15330 (N_15330,N_13784,N_13191);
nand U15331 (N_15331,N_14940,N_14549);
nand U15332 (N_15332,N_12880,N_13451);
nor U15333 (N_15333,N_13307,N_14329);
and U15334 (N_15334,N_14613,N_13511);
and U15335 (N_15335,N_14459,N_12503);
nor U15336 (N_15336,N_12721,N_13877);
and U15337 (N_15337,N_13500,N_14719);
and U15338 (N_15338,N_14387,N_13935);
or U15339 (N_15339,N_13595,N_14796);
and U15340 (N_15340,N_13077,N_13562);
nor U15341 (N_15341,N_14499,N_13987);
or U15342 (N_15342,N_13678,N_13391);
nor U15343 (N_15343,N_13745,N_13240);
nor U15344 (N_15344,N_12589,N_14207);
and U15345 (N_15345,N_13347,N_14288);
or U15346 (N_15346,N_14371,N_14187);
or U15347 (N_15347,N_13431,N_13086);
nor U15348 (N_15348,N_13116,N_13493);
nor U15349 (N_15349,N_14108,N_14854);
nand U15350 (N_15350,N_12775,N_12894);
nand U15351 (N_15351,N_12893,N_14495);
nor U15352 (N_15352,N_13660,N_14109);
and U15353 (N_15353,N_12772,N_12895);
or U15354 (N_15354,N_14633,N_13171);
or U15355 (N_15355,N_12973,N_12962);
nor U15356 (N_15356,N_14764,N_13893);
nand U15357 (N_15357,N_13190,N_13969);
nand U15358 (N_15358,N_14212,N_14848);
nor U15359 (N_15359,N_13730,N_14704);
or U15360 (N_15360,N_14520,N_13480);
nor U15361 (N_15361,N_14681,N_13132);
or U15362 (N_15362,N_12977,N_14251);
nor U15363 (N_15363,N_12814,N_13273);
or U15364 (N_15364,N_13383,N_13405);
or U15365 (N_15365,N_14611,N_13102);
nand U15366 (N_15366,N_14178,N_14663);
nand U15367 (N_15367,N_14564,N_12508);
or U15368 (N_15368,N_13479,N_13790);
nor U15369 (N_15369,N_12958,N_12639);
nor U15370 (N_15370,N_12778,N_13589);
or U15371 (N_15371,N_12592,N_13101);
and U15372 (N_15372,N_12972,N_13434);
and U15373 (N_15373,N_13866,N_14070);
or U15374 (N_15374,N_14570,N_14496);
and U15375 (N_15375,N_13384,N_14492);
and U15376 (N_15376,N_14331,N_12535);
or U15377 (N_15377,N_13416,N_12804);
or U15378 (N_15378,N_14203,N_13905);
nand U15379 (N_15379,N_14056,N_12750);
nand U15380 (N_15380,N_12660,N_13736);
or U15381 (N_15381,N_13571,N_14406);
or U15382 (N_15382,N_13901,N_13409);
nor U15383 (N_15383,N_12531,N_13718);
or U15384 (N_15384,N_13950,N_14985);
and U15385 (N_15385,N_13648,N_14076);
and U15386 (N_15386,N_14142,N_13129);
and U15387 (N_15387,N_13181,N_14925);
and U15388 (N_15388,N_12631,N_12637);
nor U15389 (N_15389,N_12649,N_14738);
and U15390 (N_15390,N_14360,N_12666);
and U15391 (N_15391,N_13957,N_13873);
nand U15392 (N_15392,N_14864,N_13447);
or U15393 (N_15393,N_13411,N_14184);
nor U15394 (N_15394,N_14664,N_14762);
and U15395 (N_15395,N_14444,N_13228);
nand U15396 (N_15396,N_14812,N_14748);
or U15397 (N_15397,N_12755,N_14761);
nor U15398 (N_15398,N_13598,N_14350);
and U15399 (N_15399,N_14017,N_13710);
and U15400 (N_15400,N_14779,N_13995);
and U15401 (N_15401,N_14943,N_14312);
and U15402 (N_15402,N_14380,N_13609);
and U15403 (N_15403,N_14020,N_12788);
and U15404 (N_15404,N_13964,N_12510);
or U15405 (N_15405,N_13757,N_13252);
and U15406 (N_15406,N_14297,N_12786);
and U15407 (N_15407,N_13754,N_12898);
nor U15408 (N_15408,N_13027,N_12539);
xor U15409 (N_15409,N_12857,N_13810);
and U15410 (N_15410,N_13908,N_13046);
nor U15411 (N_15411,N_13561,N_14644);
nand U15412 (N_15412,N_13063,N_14733);
nor U15413 (N_15413,N_13632,N_13627);
or U15414 (N_15414,N_13548,N_13527);
nor U15415 (N_15415,N_14435,N_12578);
or U15416 (N_15416,N_14863,N_13175);
xor U15417 (N_15417,N_13249,N_13421);
nand U15418 (N_15418,N_13549,N_12731);
nand U15419 (N_15419,N_13338,N_13062);
nand U15420 (N_15420,N_12609,N_13216);
nor U15421 (N_15421,N_13453,N_12997);
or U15422 (N_15422,N_13842,N_12845);
and U15423 (N_15423,N_14647,N_13387);
nor U15424 (N_15424,N_13887,N_14381);
or U15425 (N_15425,N_13870,N_13933);
or U15426 (N_15426,N_14612,N_14072);
nor U15427 (N_15427,N_14333,N_13335);
or U15428 (N_15428,N_14723,N_13666);
nor U15429 (N_15429,N_12754,N_13972);
nor U15430 (N_15430,N_13093,N_13138);
or U15431 (N_15431,N_14803,N_14186);
nand U15432 (N_15432,N_13837,N_13267);
nand U15433 (N_15433,N_14237,N_13282);
and U15434 (N_15434,N_12858,N_13628);
nor U15435 (N_15435,N_13306,N_13649);
nand U15436 (N_15436,N_13049,N_12983);
and U15437 (N_15437,N_14054,N_13406);
nor U15438 (N_15438,N_14990,N_12570);
or U15439 (N_15439,N_14200,N_14587);
or U15440 (N_15440,N_13440,N_14637);
nor U15441 (N_15441,N_12751,N_14986);
or U15442 (N_15442,N_13872,N_12663);
nor U15443 (N_15443,N_13095,N_14391);
nor U15444 (N_15444,N_13781,N_14810);
xnor U15445 (N_15445,N_13528,N_14818);
nor U15446 (N_15446,N_12540,N_13679);
or U15447 (N_15447,N_12689,N_13787);
nand U15448 (N_15448,N_14747,N_13830);
or U15449 (N_15449,N_12506,N_13395);
nor U15450 (N_15450,N_14141,N_13400);
and U15451 (N_15451,N_14417,N_14695);
nor U15452 (N_15452,N_12619,N_13709);
and U15453 (N_15453,N_13402,N_13897);
nand U15454 (N_15454,N_12549,N_13539);
and U15455 (N_15455,N_13556,N_14847);
and U15456 (N_15456,N_14806,N_12791);
or U15457 (N_15457,N_12724,N_14226);
nand U15458 (N_15458,N_13956,N_13765);
nand U15459 (N_15459,N_13715,N_13988);
and U15460 (N_15460,N_13991,N_14500);
or U15461 (N_15461,N_12849,N_14712);
and U15462 (N_15462,N_14718,N_14165);
nand U15463 (N_15463,N_14287,N_13508);
nor U15464 (N_15464,N_12511,N_14340);
nor U15465 (N_15465,N_12803,N_13978);
nor U15466 (N_15466,N_14082,N_13339);
nand U15467 (N_15467,N_13210,N_12939);
or U15468 (N_15468,N_12773,N_14814);
nand U15469 (N_15469,N_12543,N_13474);
nand U15470 (N_15470,N_13371,N_13276);
nor U15471 (N_15471,N_12741,N_12559);
or U15472 (N_15472,N_13776,N_12674);
and U15473 (N_15473,N_14509,N_13168);
nand U15474 (N_15474,N_12842,N_13018);
or U15475 (N_15475,N_13965,N_13923);
and U15476 (N_15476,N_14137,N_13001);
nand U15477 (N_15477,N_12564,N_13828);
or U15478 (N_15478,N_13071,N_13042);
or U15479 (N_15479,N_13159,N_13363);
or U15480 (N_15480,N_14426,N_13105);
or U15481 (N_15481,N_14937,N_12968);
or U15482 (N_15482,N_14768,N_13800);
nand U15483 (N_15483,N_14014,N_13334);
and U15484 (N_15484,N_14172,N_13211);
and U15485 (N_15485,N_13180,N_14478);
nor U15486 (N_15486,N_14094,N_13017);
and U15487 (N_15487,N_12646,N_14677);
and U15488 (N_15488,N_14269,N_14691);
nor U15489 (N_15489,N_13836,N_14161);
or U15490 (N_15490,N_13918,N_13361);
nand U15491 (N_15491,N_12709,N_13560);
nand U15492 (N_15492,N_14086,N_12579);
and U15493 (N_15493,N_12602,N_13326);
and U15494 (N_15494,N_13714,N_13886);
nand U15495 (N_15495,N_13277,N_13198);
nand U15496 (N_15496,N_12971,N_14555);
or U15497 (N_15497,N_14781,N_12753);
and U15498 (N_15498,N_13805,N_13217);
and U15499 (N_15499,N_14745,N_13134);
or U15500 (N_15500,N_13798,N_13551);
nand U15501 (N_15501,N_13960,N_13778);
nand U15502 (N_15502,N_14788,N_13535);
nand U15503 (N_15503,N_13318,N_12558);
and U15504 (N_15504,N_13773,N_14844);
and U15505 (N_15505,N_13728,N_14440);
nand U15506 (N_15506,N_12658,N_13237);
or U15507 (N_15507,N_14335,N_14210);
xor U15508 (N_15508,N_14962,N_13346);
and U15509 (N_15509,N_13427,N_13596);
nor U15510 (N_15510,N_14973,N_14477);
nor U15511 (N_15511,N_13255,N_13850);
nor U15512 (N_15512,N_13705,N_13215);
or U15513 (N_15513,N_14129,N_14262);
and U15514 (N_15514,N_12942,N_12542);
and U15515 (N_15515,N_13896,N_13777);
and U15516 (N_15516,N_14073,N_14394);
and U15517 (N_15517,N_12545,N_14398);
or U15518 (N_15518,N_13251,N_13076);
nand U15519 (N_15519,N_14909,N_13067);
and U15520 (N_15520,N_13513,N_12500);
and U15521 (N_15521,N_12887,N_12583);
and U15522 (N_15522,N_13100,N_13867);
nor U15523 (N_15523,N_12627,N_14291);
nor U15524 (N_15524,N_13775,N_14639);
nand U15525 (N_15525,N_14685,N_14431);
nor U15526 (N_15526,N_14598,N_14507);
nor U15527 (N_15527,N_14175,N_14097);
nor U15528 (N_15528,N_13055,N_14005);
nand U15529 (N_15529,N_12915,N_13636);
or U15530 (N_15530,N_14786,N_14308);
or U15531 (N_15531,N_14327,N_13331);
or U15532 (N_15532,N_12826,N_14201);
or U15533 (N_15533,N_14843,N_14153);
nor U15534 (N_15534,N_13080,N_12956);
nand U15535 (N_15535,N_12923,N_14282);
nand U15536 (N_15536,N_13121,N_14794);
and U15537 (N_15537,N_13895,N_14361);
or U15538 (N_15538,N_12774,N_12726);
or U15539 (N_15539,N_13463,N_14857);
nor U15540 (N_15540,N_14316,N_13435);
nand U15541 (N_15541,N_12533,N_14473);
or U15542 (N_15542,N_13167,N_12683);
and U15543 (N_15543,N_12733,N_12690);
or U15544 (N_15544,N_13315,N_14964);
nand U15545 (N_15545,N_13683,N_13860);
and U15546 (N_15546,N_14591,N_14683);
nor U15547 (N_15547,N_14479,N_14032);
or U15548 (N_15548,N_13424,N_12628);
and U15549 (N_15549,N_12802,N_13445);
xor U15550 (N_15550,N_13239,N_13352);
nand U15551 (N_15551,N_14157,N_14363);
nor U15552 (N_15552,N_13231,N_14271);
nand U15553 (N_15553,N_12626,N_13412);
and U15554 (N_15554,N_12975,N_13652);
and U15555 (N_15555,N_12896,N_13222);
nand U15556 (N_15556,N_14787,N_14547);
and U15557 (N_15557,N_14336,N_14115);
nor U15558 (N_15558,N_12916,N_14419);
nand U15559 (N_15559,N_12520,N_13142);
nand U15560 (N_15560,N_12902,N_13265);
nand U15561 (N_15561,N_14100,N_13750);
and U15562 (N_15562,N_14058,N_14375);
nor U15563 (N_15563,N_14068,N_14636);
nor U15564 (N_15564,N_14868,N_13189);
nor U15565 (N_15565,N_14751,N_12866);
or U15566 (N_15566,N_13807,N_14265);
nand U15567 (N_15567,N_13927,N_13663);
or U15568 (N_15568,N_14916,N_12832);
or U15569 (N_15569,N_13958,N_13506);
and U15570 (N_15570,N_13109,N_14516);
nor U15571 (N_15571,N_13977,N_14580);
nand U15572 (N_15572,N_13849,N_14339);
nand U15573 (N_15573,N_14286,N_14730);
and U15574 (N_15574,N_13763,N_14197);
nor U15575 (N_15575,N_12591,N_12614);
and U15576 (N_15576,N_14635,N_14807);
or U15577 (N_15577,N_13279,N_13961);
nor U15578 (N_15578,N_14386,N_14763);
nor U15579 (N_15579,N_14384,N_13755);
or U15580 (N_15580,N_14104,N_13829);
and U15581 (N_15581,N_14012,N_12695);
nand U15582 (N_15582,N_13756,N_12582);
or U15583 (N_15583,N_12817,N_14770);
or U15584 (N_15584,N_13465,N_12717);
nand U15585 (N_15585,N_12672,N_14008);
or U15586 (N_15586,N_13432,N_13202);
nand U15587 (N_15587,N_14323,N_14777);
or U15588 (N_15588,N_13880,N_12808);
and U15589 (N_15589,N_14221,N_13015);
nor U15590 (N_15590,N_13611,N_14456);
nand U15591 (N_15591,N_14427,N_14666);
and U15592 (N_15592,N_14978,N_14220);
and U15593 (N_15593,N_14991,N_12979);
and U15594 (N_15594,N_12518,N_14855);
nor U15595 (N_15595,N_13623,N_13515);
or U15596 (N_15596,N_14041,N_14959);
and U15597 (N_15597,N_14346,N_13462);
nor U15598 (N_15598,N_14223,N_12538);
nand U15599 (N_15599,N_14177,N_13013);
nor U15600 (N_15600,N_13883,N_14337);
nor U15601 (N_15601,N_12828,N_12978);
or U15602 (N_15602,N_12799,N_14835);
and U15603 (N_15603,N_13482,N_12623);
and U15604 (N_15604,N_13761,N_12522);
nor U15605 (N_15605,N_12502,N_14402);
nor U15606 (N_15606,N_13036,N_14775);
nor U15607 (N_15607,N_14063,N_14273);
nand U15608 (N_15608,N_14345,N_14805);
nand U15609 (N_15609,N_13024,N_14092);
nand U15610 (N_15610,N_12938,N_12636);
nor U15611 (N_15611,N_14024,N_14128);
and U15612 (N_15612,N_14673,N_13408);
and U15613 (N_15613,N_12596,N_14630);
nand U15614 (N_15614,N_13438,N_13035);
or U15615 (N_15615,N_14558,N_13051);
nor U15616 (N_15616,N_14576,N_13966);
and U15617 (N_15617,N_14703,N_14825);
or U15618 (N_15618,N_13099,N_14646);
nor U15619 (N_15619,N_12734,N_12561);
nor U15620 (N_15620,N_13247,N_13783);
nor U15621 (N_15621,N_14608,N_14057);
nand U15622 (N_15622,N_14883,N_13532);
and U15623 (N_15623,N_14002,N_12604);
nor U15624 (N_15624,N_12864,N_13081);
or U15625 (N_15625,N_13137,N_13123);
and U15626 (N_15626,N_12918,N_14676);
or U15627 (N_15627,N_14648,N_14994);
nor U15628 (N_15628,N_12556,N_13106);
nand U15629 (N_15629,N_13000,N_14229);
nor U15630 (N_15630,N_13808,N_12961);
nand U15631 (N_15631,N_13250,N_14618);
and U15632 (N_15632,N_13502,N_12509);
or U15633 (N_15633,N_13150,N_13456);
or U15634 (N_15634,N_14482,N_13593);
nand U15635 (N_15635,N_14224,N_13687);
or U15636 (N_15636,N_14311,N_12712);
nand U15637 (N_15637,N_14711,N_14113);
nor U15638 (N_15638,N_12615,N_13152);
and U15639 (N_15639,N_13906,N_12560);
and U15640 (N_15640,N_13726,N_13261);
or U15641 (N_15641,N_14815,N_14833);
nand U15642 (N_15642,N_14832,N_14415);
or U15643 (N_15643,N_12925,N_14077);
or U15644 (N_15644,N_13390,N_14007);
nor U15645 (N_15645,N_14649,N_12685);
or U15646 (N_15646,N_14887,N_12546);
and U15647 (N_15647,N_14480,N_13826);
or U15648 (N_15648,N_14457,N_13524);
xnor U15649 (N_15649,N_14950,N_14531);
or U15650 (N_15650,N_14776,N_14615);
nand U15651 (N_15651,N_13644,N_13407);
nor U15652 (N_15652,N_14124,N_13430);
and U15653 (N_15653,N_14409,N_14298);
nand U15654 (N_15654,N_14230,N_14882);
nand U15655 (N_15655,N_13061,N_12584);
nor U15656 (N_15656,N_13510,N_14127);
or U15657 (N_15657,N_14913,N_14111);
and U15658 (N_15658,N_14869,N_13780);
and U15659 (N_15659,N_13925,N_13342);
or U15660 (N_15660,N_12527,N_13949);
and U15661 (N_15661,N_12742,N_13794);
and U15662 (N_15662,N_12909,N_13945);
or U15663 (N_15663,N_14765,N_12824);
nand U15664 (N_15664,N_13178,N_14836);
nor U15665 (N_15665,N_14252,N_14971);
nor U15666 (N_15666,N_12706,N_12763);
nand U15667 (N_15667,N_13999,N_14219);
nand U15668 (N_15668,N_13473,N_14450);
nand U15669 (N_15669,N_13179,N_13297);
or U15670 (N_15670,N_13083,N_14672);
and U15671 (N_15671,N_14374,N_12719);
nand U15672 (N_15672,N_14295,N_13303);
and U15673 (N_15673,N_12838,N_13911);
or U15674 (N_15674,N_14083,N_13937);
nand U15675 (N_15675,N_14102,N_13139);
or U15676 (N_15676,N_14894,N_14860);
nand U15677 (N_15677,N_13809,N_12676);
nand U15678 (N_15678,N_12534,N_13314);
nand U15679 (N_15679,N_12955,N_14572);
nand U15680 (N_15680,N_13356,N_13302);
and U15681 (N_15681,N_13760,N_12795);
nor U15682 (N_15682,N_12565,N_14488);
nand U15683 (N_15683,N_13245,N_13143);
or U15684 (N_15684,N_13369,N_12610);
or U15685 (N_15685,N_14904,N_14930);
and U15686 (N_15686,N_14928,N_14543);
nor U15687 (N_15687,N_12748,N_14472);
nand U15688 (N_15688,N_13119,N_13624);
nor U15689 (N_15689,N_14154,N_13214);
or U15690 (N_15690,N_12668,N_14567);
and U15691 (N_15691,N_13328,N_14018);
nand U15692 (N_15692,N_14713,N_13658);
nand U15693 (N_15693,N_14158,N_12823);
and U15694 (N_15694,N_14667,N_12675);
nand U15695 (N_15695,N_14405,N_13362);
and U15696 (N_15696,N_12727,N_14170);
or U15697 (N_15697,N_12555,N_14031);
or U15698 (N_15698,N_14512,N_13993);
nor U15699 (N_15699,N_12853,N_14379);
and U15700 (N_15700,N_13165,N_12553);
or U15701 (N_15701,N_13699,N_14554);
and U15702 (N_15702,N_14438,N_14769);
nand U15703 (N_15703,N_13912,N_14811);
nand U15704 (N_15704,N_13127,N_13795);
and U15705 (N_15705,N_14865,N_13128);
or U15706 (N_15706,N_14423,N_13172);
nand U15707 (N_15707,N_12735,N_13620);
nand U15708 (N_15708,N_13544,N_13789);
nand U15709 (N_15709,N_13915,N_13603);
or U15710 (N_15710,N_14088,N_14424);
nor U15711 (N_15711,N_13537,N_14628);
and U15712 (N_15712,N_12595,N_12952);
nand U15713 (N_15713,N_13052,N_14593);
or U15714 (N_15714,N_14542,N_12863);
nor U15715 (N_15715,N_14303,N_13646);
nor U15716 (N_15716,N_13005,N_12797);
nand U15717 (N_15717,N_13268,N_14356);
nor U15718 (N_15718,N_14793,N_14918);
and U15719 (N_15719,N_14501,N_13864);
nand U15720 (N_15720,N_12629,N_14981);
or U15721 (N_15721,N_13019,N_14722);
and U15722 (N_15722,N_13366,N_14888);
or U15723 (N_15723,N_14353,N_13786);
and U15724 (N_15724,N_13025,N_13835);
nor U15725 (N_15725,N_13811,N_13381);
and U15726 (N_15726,N_12825,N_14502);
nor U15727 (N_15727,N_14274,N_13641);
nand U15728 (N_15728,N_12716,N_14439);
or U15729 (N_15729,N_13770,N_13592);
and U15730 (N_15730,N_13443,N_13588);
xnor U15731 (N_15731,N_14464,N_12505);
nor U15732 (N_15732,N_14556,N_13700);
or U15733 (N_15733,N_12855,N_13902);
nor U15734 (N_15734,N_13317,N_14294);
nor U15735 (N_15735,N_13197,N_14388);
and U15736 (N_15736,N_12940,N_14897);
nor U15737 (N_15737,N_14085,N_14600);
nand U15738 (N_15738,N_14956,N_13657);
or U15739 (N_15739,N_14715,N_12829);
nor U15740 (N_15740,N_14352,N_13298);
nand U15741 (N_15741,N_13221,N_13512);
nor U15742 (N_15742,N_14489,N_13460);
xor U15743 (N_15743,N_14819,N_14911);
and U15744 (N_15744,N_14324,N_13963);
nor U15745 (N_15745,N_12684,N_13861);
nand U15746 (N_15746,N_14828,N_13685);
nand U15747 (N_15747,N_12625,N_13521);
or U15748 (N_15748,N_13688,N_14801);
and U15749 (N_15749,N_14461,N_14051);
and U15750 (N_15750,N_14837,N_14133);
or U15751 (N_15751,N_13853,N_14243);
and U15752 (N_15752,N_13289,N_13574);
and U15753 (N_15753,N_13591,N_13939);
nor U15754 (N_15754,N_12513,N_14270);
and U15755 (N_15755,N_13846,N_12927);
or U15756 (N_15756,N_14015,N_13330);
nor U15757 (N_15757,N_14705,N_13639);
nand U15758 (N_15758,N_14789,N_12548);
or U15759 (N_15759,N_14716,N_12641);
or U15760 (N_15760,N_12913,N_14975);
nor U15761 (N_15761,N_14443,N_13423);
nand U15762 (N_15762,N_14702,N_14800);
nand U15763 (N_15763,N_13367,N_14899);
and U15764 (N_15764,N_14497,N_12776);
or U15765 (N_15765,N_14680,N_14313);
nor U15766 (N_15766,N_14506,N_14385);
and U15767 (N_15767,N_13774,N_13892);
and U15768 (N_15768,N_14942,N_12981);
nor U15769 (N_15769,N_13650,N_12792);
or U15770 (N_15770,N_13832,N_14945);
and U15771 (N_15771,N_14148,N_13458);
nor U15772 (N_15772,N_12922,N_13206);
and U15773 (N_15773,N_12787,N_12764);
nor U15774 (N_15774,N_12783,N_14515);
or U15775 (N_15775,N_13313,N_13825);
and U15776 (N_15776,N_12590,N_13677);
or U15777 (N_15777,N_13731,N_13158);
and U15778 (N_15778,N_14146,N_12620);
nand U15779 (N_15779,N_13030,N_14289);
or U15780 (N_15780,N_12933,N_12905);
nor U15781 (N_15781,N_12612,N_12635);
nor U15782 (N_15782,N_13393,N_14867);
nand U15783 (N_15783,N_13155,N_14044);
and U15784 (N_15784,N_14455,N_12822);
and U15785 (N_15785,N_12514,N_12745);
or U15786 (N_15786,N_13485,N_13351);
and U15787 (N_15787,N_12530,N_14822);
or U15788 (N_15788,N_13058,N_13612);
nor U15789 (N_15789,N_14631,N_13428);
and U15790 (N_15790,N_13838,N_13904);
and U15791 (N_15791,N_13494,N_13467);
or U15792 (N_15792,N_13617,N_13009);
or U15793 (N_15793,N_14771,N_14357);
nor U15794 (N_15794,N_14425,N_14283);
and U15795 (N_15795,N_13785,N_13547);
nand U15796 (N_15796,N_14099,N_12999);
and U15797 (N_15797,N_13869,N_13997);
or U15798 (N_15798,N_14659,N_13669);
or U15799 (N_15799,N_13743,N_13762);
nand U15800 (N_15800,N_14118,N_12819);
nand U15801 (N_15801,N_14606,N_14276);
nand U15802 (N_15802,N_12848,N_14454);
or U15803 (N_15803,N_14307,N_12594);
nor U15804 (N_15804,N_14261,N_12563);
and U15805 (N_15805,N_13599,N_13671);
nand U15806 (N_15806,N_13433,N_13096);
and U15807 (N_15807,N_12528,N_14491);
nor U15808 (N_15808,N_13618,N_12964);
nor U15809 (N_15809,N_13448,N_14376);
nor U15810 (N_15810,N_14081,N_13373);
nand U15811 (N_15811,N_13703,N_13504);
and U15812 (N_15812,N_13157,N_14009);
or U15813 (N_15813,N_12651,N_13926);
and U15814 (N_15814,N_14093,N_14710);
nand U15815 (N_15815,N_12580,N_12947);
or U15816 (N_15816,N_13580,N_12852);
nand U15817 (N_15817,N_14414,N_13114);
nand U15818 (N_15818,N_12581,N_13284);
and U15819 (N_15819,N_14709,N_14022);
nor U15820 (N_15820,N_14692,N_13243);
or U15821 (N_15821,N_13954,N_13148);
and U15822 (N_15822,N_14120,N_13929);
and U15823 (N_15823,N_14367,N_13840);
and U15824 (N_15824,N_13900,N_12643);
or U15825 (N_15825,N_12801,N_13010);
nand U15826 (N_15826,N_13359,N_13834);
nor U15827 (N_15827,N_13694,N_14239);
nand U15828 (N_15828,N_13647,N_13475);
or U15829 (N_15829,N_14255,N_12873);
nor U15830 (N_15830,N_13450,N_13290);
nor U15831 (N_15831,N_14037,N_12992);
nand U15832 (N_15832,N_14557,N_14678);
nor U15833 (N_15833,N_12541,N_12874);
or U15834 (N_15834,N_13766,N_13006);
nand U15835 (N_15835,N_13023,N_14302);
and U15836 (N_15836,N_14840,N_13878);
nor U15837 (N_15837,N_12793,N_14228);
or U15838 (N_15838,N_13056,N_14999);
nor U15839 (N_15839,N_13559,N_13670);
and U15840 (N_15840,N_13656,N_14742);
nand U15841 (N_15841,N_13684,N_14055);
nand U15842 (N_15842,N_13280,N_14766);
nand U15843 (N_15843,N_12524,N_14293);
nor U15844 (N_15844,N_13903,N_13188);
nand U15845 (N_15845,N_13797,N_14505);
nand U15846 (N_15846,N_13764,N_13226);
nand U15847 (N_15847,N_14447,N_12701);
or U15848 (N_15848,N_14599,N_14850);
nor U15849 (N_15849,N_13441,N_14804);
xor U15850 (N_15850,N_13645,N_13170);
nor U15851 (N_15851,N_12946,N_14466);
or U15852 (N_15852,N_13414,N_13292);
nand U15853 (N_15853,N_14741,N_13720);
and U15854 (N_15854,N_14902,N_12537);
nor U15855 (N_15855,N_14050,N_13577);
and U15856 (N_15856,N_13793,N_14783);
nand U15857 (N_15857,N_14654,N_13296);
and U15858 (N_15858,N_13455,N_13288);
nand U15859 (N_15859,N_13380,N_14662);
xnor U15860 (N_15860,N_12667,N_14866);
or U15861 (N_15861,N_12633,N_12617);
and U15862 (N_15862,N_13098,N_12737);
or U15863 (N_15863,N_14355,N_13072);
nand U15864 (N_15864,N_12521,N_13814);
nand U15865 (N_15865,N_13442,N_14658);
nand U15866 (N_15866,N_14661,N_12662);
or U15867 (N_15867,N_13425,N_14369);
and U15868 (N_15868,N_14465,N_13998);
or U15869 (N_15869,N_12536,N_13824);
or U15870 (N_15870,N_12747,N_12924);
nand U15871 (N_15871,N_14338,N_14995);
and U15872 (N_15872,N_13631,N_14071);
or U15873 (N_15873,N_13931,N_14103);
nand U15874 (N_15874,N_14264,N_14389);
nor U15875 (N_15875,N_13936,N_14586);
nand U15876 (N_15876,N_12948,N_14539);
nand U15877 (N_15877,N_13185,N_13472);
nor U15878 (N_15878,N_14729,N_14185);
nor U15879 (N_15879,N_12813,N_13489);
and U15880 (N_15880,N_13464,N_12700);
or U15881 (N_15881,N_12679,N_13354);
nand U15882 (N_15882,N_14332,N_14131);
nand U15883 (N_15883,N_12779,N_14460);
nor U15884 (N_15884,N_14156,N_14579);
nor U15885 (N_15885,N_14259,N_13230);
nand U15886 (N_15886,N_13043,N_14067);
or U15887 (N_15887,N_14416,N_14432);
or U15888 (N_15888,N_12907,N_14622);
nand U15889 (N_15889,N_13223,N_14285);
and U15890 (N_15890,N_14196,N_13469);
nand U15891 (N_15891,N_13498,N_13822);
or U15892 (N_15892,N_14059,N_13934);
or U15893 (N_15893,N_14245,N_14614);
nand U15894 (N_15894,N_13586,N_12790);
nand U15895 (N_15895,N_13110,N_14065);
nor U15896 (N_15896,N_14873,N_13320);
nor U15897 (N_15897,N_13452,N_13768);
nand U15898 (N_15898,N_13156,N_13004);
or U15899 (N_15899,N_13270,N_14214);
nor U15900 (N_15900,N_14926,N_12654);
nand U15901 (N_15901,N_13196,N_14235);
or U15902 (N_15902,N_12820,N_14653);
nor U15903 (N_15903,N_13919,N_14523);
nand U15904 (N_15904,N_14025,N_12708);
nand U15905 (N_15905,N_14522,N_13065);
nor U15906 (N_15906,N_12698,N_14422);
nor U15907 (N_15907,N_13205,N_14134);
and U15908 (N_15908,N_13117,N_14689);
nor U15909 (N_15909,N_13461,N_13868);
nor U15910 (N_15910,N_14519,N_14029);
or U15911 (N_15911,N_14656,N_13312);
nand U15912 (N_15912,N_14566,N_12720);
nor U15913 (N_15913,N_13625,N_13360);
and U15914 (N_15914,N_12525,N_12837);
nand U15915 (N_15915,N_13749,N_14562);
and U15916 (N_15916,N_14451,N_14373);
and U15917 (N_15917,N_14827,N_14744);
nor U15918 (N_15918,N_14528,N_12744);
and U15919 (N_15919,N_14626,N_13115);
or U15920 (N_15920,N_13426,N_13107);
or U15921 (N_15921,N_14342,N_13523);
and U15922 (N_15922,N_13894,N_12729);
nor U15923 (N_15923,N_13048,N_13552);
nor U15924 (N_15924,N_12574,N_14445);
xor U15925 (N_15925,N_13108,N_14254);
or U15926 (N_15926,N_13038,N_13594);
and U15927 (N_15927,N_13667,N_14485);
nor U15928 (N_15928,N_13087,N_13146);
nor U15929 (N_15929,N_13260,N_12806);
and U15930 (N_15930,N_14155,N_13884);
nand U15931 (N_15931,N_14784,N_13735);
nor U15932 (N_15932,N_14468,N_13069);
or U15933 (N_15933,N_14434,N_13717);
nand U15934 (N_15934,N_13538,N_14514);
and U15935 (N_15935,N_12815,N_12926);
nand U15936 (N_15936,N_12851,N_13806);
or U15937 (N_15937,N_14571,N_13801);
nand U15938 (N_15938,N_13550,N_13135);
or U15939 (N_15939,N_12762,N_14234);
nor U15940 (N_15940,N_13542,N_12910);
nand U15941 (N_15941,N_14540,N_13659);
nand U15942 (N_15942,N_14721,N_14969);
nor U15943 (N_15943,N_12687,N_12618);
and U15944 (N_15944,N_14876,N_14292);
or U15945 (N_15945,N_14318,N_13410);
nor U15946 (N_15946,N_14244,N_12884);
or U15947 (N_15947,N_12759,N_12603);
nor U15948 (N_15948,N_13734,N_12765);
nor U15949 (N_15949,N_13332,N_12547);
and U15950 (N_15950,N_14524,N_14504);
and U15951 (N_15951,N_13304,N_14816);
or U15952 (N_15952,N_14116,N_14430);
nor U15953 (N_15953,N_14166,N_13802);
and U15954 (N_15954,N_14645,N_14824);
and U15955 (N_15955,N_12740,N_14404);
nand U15956 (N_15956,N_13852,N_14366);
nor U15957 (N_15957,N_12757,N_14242);
or U15958 (N_15958,N_12836,N_14174);
and U15959 (N_15959,N_13959,N_13301);
and U15960 (N_15960,N_14026,N_13477);
or U15961 (N_15961,N_14149,N_14538);
nand U15962 (N_15962,N_13293,N_13885);
nand U15963 (N_15963,N_12682,N_12789);
or U15964 (N_15964,N_14304,N_14163);
or U15965 (N_15965,N_13073,N_13813);
or U15966 (N_15966,N_13044,N_13698);
and U15967 (N_15967,N_12575,N_14279);
and U15968 (N_15968,N_13653,N_14192);
nand U15969 (N_15969,N_13729,N_13144);
or U15970 (N_15970,N_14674,N_13759);
nor U15971 (N_15971,N_14453,N_14739);
nand U15972 (N_15972,N_14147,N_13979);
xor U15973 (N_15973,N_13386,N_12691);
nand U15974 (N_15974,N_13350,N_13676);
nand U15975 (N_15975,N_13200,N_13642);
or U15976 (N_15976,N_12821,N_13253);
nor U15977 (N_15977,N_14972,N_13343);
or U15978 (N_15978,N_13638,N_12963);
nand U15979 (N_15979,N_14551,N_14912);
nor U15980 (N_15980,N_12919,N_12647);
nand U15981 (N_15981,N_13269,N_13882);
nor U15982 (N_15982,N_14204,N_13681);
nand U15983 (N_15983,N_12621,N_13264);
and U15984 (N_15984,N_12966,N_14660);
and U15985 (N_15985,N_13012,N_12678);
nor U15986 (N_15986,N_14176,N_13615);
xor U15987 (N_15987,N_14300,N_13907);
nor U15988 (N_15988,N_14173,N_13517);
and U15989 (N_15989,N_12912,N_14823);
nor U15990 (N_15990,N_14621,N_12671);
nand U15991 (N_15991,N_12936,N_14241);
and U15992 (N_15992,N_14167,N_12807);
nand U15993 (N_15993,N_12718,N_12805);
nor U15994 (N_15994,N_14699,N_14536);
or U15995 (N_15995,N_14272,N_14325);
nor U15996 (N_15996,N_14028,N_12616);
nand U15997 (N_15997,N_14690,N_12990);
nand U15998 (N_15998,N_14728,N_13141);
and U15999 (N_15999,N_14583,N_13913);
or U16000 (N_16000,N_14922,N_13948);
or U16001 (N_16001,N_14541,N_13799);
and U16002 (N_16002,N_13103,N_13706);
and U16003 (N_16003,N_14330,N_14845);
nor U16004 (N_16004,N_13737,N_14494);
nor U16005 (N_16005,N_12950,N_13582);
and U16006 (N_16006,N_13951,N_13112);
or U16007 (N_16007,N_14420,N_13420);
nand U16008 (N_16008,N_12770,N_14225);
or U16009 (N_16009,N_12573,N_12771);
and U16010 (N_16010,N_12953,N_13483);
nor U16011 (N_16011,N_14790,N_14546);
nand U16012 (N_16012,N_13419,N_13316);
and U16013 (N_16013,N_13803,N_13819);
nor U16014 (N_16014,N_13325,N_12722);
and U16015 (N_16015,N_14284,N_12551);
nand U16016 (N_16016,N_14590,N_12957);
xnor U16017 (N_16017,N_12854,N_14921);
nor U16018 (N_16018,N_14640,N_12932);
nor U16019 (N_16019,N_14582,N_14958);
and U16020 (N_16020,N_13859,N_14487);
xnor U16021 (N_16021,N_14795,N_13779);
nor U16022 (N_16022,N_13068,N_14314);
nor U16023 (N_16023,N_14821,N_13397);
nand U16024 (N_16024,N_14872,N_14813);
and U16025 (N_16025,N_14604,N_14034);
nand U16026 (N_16026,N_12830,N_12713);
nand U16027 (N_16027,N_14545,N_14258);
nand U16028 (N_16028,N_13758,N_12904);
nor U16029 (N_16029,N_14842,N_13133);
and U16030 (N_16030,N_12642,N_12906);
and U16031 (N_16031,N_14160,N_14597);
nand U16032 (N_16032,N_12630,N_14976);
nand U16033 (N_16033,N_14623,N_13771);
nand U16034 (N_16034,N_13281,N_14933);
nand U16035 (N_16035,N_14849,N_14734);
or U16036 (N_16036,N_13355,N_14006);
or U16037 (N_16037,N_14963,N_14791);
nor U16038 (N_16038,N_14112,N_13299);
nor U16039 (N_16039,N_12611,N_13782);
nor U16040 (N_16040,N_13533,N_14707);
and U16041 (N_16041,N_14760,N_13357);
nor U16042 (N_16042,N_13635,N_12694);
nand U16043 (N_16043,N_12847,N_13569);
and U16044 (N_16044,N_14046,N_13723);
nor U16045 (N_16045,N_12710,N_13572);
nor U16046 (N_16046,N_13875,N_12715);
and U16047 (N_16047,N_13140,N_14838);
or U16048 (N_16048,N_14033,N_12890);
nor U16049 (N_16049,N_13518,N_13545);
or U16050 (N_16050,N_14809,N_13403);
nor U16051 (N_16051,N_14260,N_14238);
or U16052 (N_16052,N_14344,N_12608);
nor U16053 (N_16053,N_13070,N_14484);
or U16054 (N_16054,N_13319,N_13037);
nor U16055 (N_16055,N_14774,N_14740);
nand U16056 (N_16056,N_13392,N_13075);
nand U16057 (N_16057,N_13060,N_12624);
nand U16058 (N_16058,N_13294,N_14143);
and U16059 (N_16059,N_14984,N_12572);
or U16060 (N_16060,N_13324,N_12526);
nand U16061 (N_16061,N_13566,N_13274);
or U16062 (N_16062,N_14871,N_13120);
nor U16063 (N_16063,N_13608,N_12515);
and U16064 (N_16064,N_12859,N_14525);
nor U16065 (N_16065,N_13844,N_13719);
nand U16066 (N_16066,N_12784,N_13601);
nand U16067 (N_16067,N_14467,N_13125);
or U16068 (N_16068,N_14351,N_13340);
or U16069 (N_16069,N_12891,N_13854);
or U16070 (N_16070,N_14462,N_13651);
nor U16071 (N_16071,N_13597,N_14449);
and U16072 (N_16072,N_14190,N_13833);
nor U16073 (N_16073,N_13291,N_13855);
or U16074 (N_16074,N_14949,N_14934);
nor U16075 (N_16075,N_14211,N_13845);
and U16076 (N_16076,N_13186,N_13496);
and U16077 (N_16077,N_14407,N_12892);
and U16078 (N_16078,N_12569,N_14400);
nor U16079 (N_16079,N_12640,N_12781);
nand U16080 (N_16080,N_13501,N_12769);
and U16081 (N_16081,N_12920,N_13747);
and U16082 (N_16082,N_13078,N_13606);
nand U16083 (N_16083,N_13607,N_12782);
and U16084 (N_16084,N_13791,N_12883);
or U16085 (N_16085,N_12686,N_12585);
nor U16086 (N_16086,N_13713,N_14084);
nor U16087 (N_16087,N_14694,N_13820);
and U16088 (N_16088,N_14328,N_13236);
nor U16089 (N_16089,N_13525,N_13955);
and U16090 (N_16090,N_13514,N_14412);
or U16091 (N_16091,N_12638,N_13064);
and U16092 (N_16092,N_13823,N_13567);
nand U16093 (N_16093,N_13856,N_14087);
and U16094 (N_16094,N_13581,N_13404);
or U16095 (N_16095,N_14463,N_13476);
or U16096 (N_16096,N_14030,N_13173);
nand U16097 (N_16097,N_13952,N_14534);
nand U16098 (N_16098,N_12794,N_13881);
or U16099 (N_16099,N_12881,N_14898);
nand U16100 (N_16100,N_14117,N_13890);
or U16101 (N_16101,N_13622,N_13520);
nor U16102 (N_16102,N_12702,N_14395);
nor U16103 (N_16103,N_13792,N_13147);
or U16104 (N_16104,N_14798,N_14841);
or U16105 (N_16105,N_13697,N_13287);
xor U16106 (N_16106,N_12843,N_13499);
and U16107 (N_16107,N_13008,N_14039);
and U16108 (N_16108,N_13182,N_13668);
or U16109 (N_16109,N_13614,N_13573);
or U16110 (N_16110,N_14411,N_13149);
and U16111 (N_16111,N_14377,N_14896);
and U16112 (N_16112,N_12739,N_14592);
nor U16113 (N_16113,N_13564,N_14023);
nor U16114 (N_16114,N_13563,N_13898);
nor U16115 (N_16115,N_13570,N_14616);
nand U16116 (N_16116,N_13094,N_13285);
nand U16117 (N_16117,N_13815,N_12600);
or U16118 (N_16118,N_14322,N_14189);
or U16119 (N_16119,N_14749,N_14708);
nor U16120 (N_16120,N_12949,N_13643);
or U16121 (N_16121,N_13874,N_14202);
nand U16122 (N_16122,N_14393,N_13194);
and U16123 (N_16123,N_13118,N_14725);
nor U16124 (N_16124,N_14267,N_14365);
nor U16125 (N_16125,N_13164,N_13619);
nor U16126 (N_16126,N_14687,N_14923);
and U16127 (N_16127,N_14589,N_14119);
or U16128 (N_16128,N_14885,N_13557);
nor U16129 (N_16129,N_14696,N_14310);
nand U16130 (N_16130,N_14782,N_14151);
or U16131 (N_16131,N_14737,N_13382);
nand U16132 (N_16132,N_12901,N_12844);
nor U16133 (N_16133,N_13415,N_12921);
nand U16134 (N_16134,N_14110,N_13153);
and U16135 (N_16135,N_14458,N_13871);
and U16136 (N_16136,N_14508,N_13686);
nor U16137 (N_16137,N_14403,N_14535);
nor U16138 (N_16138,N_14966,N_13947);
or U16139 (N_16139,N_13584,N_13238);
nor U16140 (N_16140,N_12632,N_13692);
or U16141 (N_16141,N_13368,N_13695);
and U16142 (N_16142,N_14997,N_12586);
or U16143 (N_16143,N_12601,N_13398);
and U16144 (N_16144,N_13941,N_12728);
or U16145 (N_16145,N_14756,N_13422);
nand U16146 (N_16146,N_14968,N_13930);
or U16147 (N_16147,N_12930,N_14521);
nand U16148 (N_16148,N_14731,N_14846);
nand U16149 (N_16149,N_13437,N_14206);
or U16150 (N_16150,N_12656,N_14641);
nor U16151 (N_16151,N_12876,N_14090);
nor U16152 (N_16152,N_13032,N_14168);
nand U16153 (N_16153,N_13554,N_14368);
and U16154 (N_16154,N_12567,N_13910);
nor U16155 (N_16155,N_14875,N_13263);
nor U16156 (N_16156,N_14880,N_14397);
xor U16157 (N_16157,N_12834,N_14632);
or U16158 (N_16158,N_14839,N_14334);
or U16159 (N_16159,N_13154,N_13333);
nand U16160 (N_16160,N_14665,N_14066);
nor U16161 (N_16161,N_13481,N_14277);
and U16162 (N_16162,N_12598,N_14441);
nand U16163 (N_16163,N_13982,N_13674);
and U16164 (N_16164,N_13613,N_13323);
and U16165 (N_16165,N_13693,N_13924);
xnor U16166 (N_16166,N_13177,N_12714);
nand U16167 (N_16167,N_13487,N_12507);
and U16168 (N_16168,N_13059,N_14042);
nand U16169 (N_16169,N_14548,N_14686);
nor U16170 (N_16170,N_13131,N_14619);
nand U16171 (N_16171,N_13091,N_13689);
nand U16172 (N_16172,N_13640,N_14195);
and U16173 (N_16173,N_13984,N_13079);
nor U16174 (N_16174,N_13256,N_14486);
or U16175 (N_16175,N_14617,N_13742);
and U16176 (N_16176,N_13752,N_14016);
or U16177 (N_16177,N_12677,N_14182);
and U16178 (N_16178,N_13986,N_14584);
xnor U16179 (N_16179,N_13721,N_12704);
or U16180 (N_16180,N_14469,N_14910);
and U16181 (N_16181,N_14758,N_12796);
and U16182 (N_16182,N_13136,N_14799);
nor U16183 (N_16183,N_14802,N_14162);
and U16184 (N_16184,N_13707,N_14296);
nor U16185 (N_16185,N_14603,N_13053);
nor U16186 (N_16186,N_13507,N_14209);
nand U16187 (N_16187,N_13711,N_14957);
nand U16188 (N_16188,N_12657,N_12723);
nor U16189 (N_16189,N_14609,N_13976);
nand U16190 (N_16190,N_12577,N_13891);
nor U16191 (N_16191,N_12868,N_14941);
nor U16192 (N_16192,N_14410,N_14698);
nand U16193 (N_16193,N_12800,N_14396);
nand U16194 (N_16194,N_14476,N_14250);
nor U16195 (N_16195,N_12835,N_12934);
nand U16196 (N_16196,N_14138,N_13193);
and U16197 (N_16197,N_12885,N_14892);
nor U16198 (N_16198,N_14256,N_14563);
and U16199 (N_16199,N_12965,N_14098);
nand U16200 (N_16200,N_13166,N_13665);
nand U16201 (N_16201,N_14191,N_13769);
or U16202 (N_16202,N_14436,N_13558);
nand U16203 (N_16203,N_13600,N_13275);
or U16204 (N_16204,N_14879,N_12827);
nand U16205 (N_16205,N_14750,N_13047);
or U16206 (N_16206,N_14575,N_14306);
nor U16207 (N_16207,N_12622,N_12655);
and U16208 (N_16208,N_14236,N_13311);
and U16209 (N_16209,N_12991,N_12576);
or U16210 (N_16210,N_12588,N_14233);
nor U16211 (N_16211,N_13495,N_14693);
or U16212 (N_16212,N_13305,N_12673);
or U16213 (N_16213,N_13985,N_13740);
or U16214 (N_16214,N_14027,N_13879);
or U16215 (N_16215,N_13996,N_14929);
nand U16216 (N_16216,N_14061,N_13413);
or U16217 (N_16217,N_14893,N_14908);
and U16218 (N_16218,N_13176,N_14927);
or U16219 (N_16219,N_12664,N_13192);
or U16220 (N_16220,N_12768,N_13309);
nand U16221 (N_16221,N_13484,N_13974);
or U16222 (N_16222,N_12516,N_14169);
and U16223 (N_16223,N_14553,N_13516);
nand U16224 (N_16224,N_12986,N_13503);
and U16225 (N_16225,N_13725,N_14987);
and U16226 (N_16226,N_14955,N_13531);
nor U16227 (N_16227,N_13916,N_13232);
or U16228 (N_16228,N_14218,N_13218);
nor U16229 (N_16229,N_14418,N_12998);
and U16230 (N_16230,N_12929,N_12900);
nand U16231 (N_16231,N_14706,N_13057);
nor U16232 (N_16232,N_13796,N_14552);
nor U16233 (N_16233,N_14198,N_13491);
nor U16234 (N_16234,N_13417,N_14989);
or U16235 (N_16235,N_14428,N_14780);
and U16236 (N_16236,N_13039,N_14982);
nor U16237 (N_16237,N_14961,N_14977);
or U16238 (N_16238,N_14348,N_14301);
and U16239 (N_16239,N_14939,N_13553);
or U16240 (N_16240,N_14215,N_12951);
or U16241 (N_16241,N_14914,N_12861);
or U16242 (N_16242,N_13921,N_12688);
nand U16243 (N_16243,N_13962,N_13225);
nor U16244 (N_16244,N_13888,N_13388);
nand U16245 (N_16245,N_14935,N_13209);
nand U16246 (N_16246,N_13922,N_13486);
nor U16247 (N_16247,N_13266,N_13509);
and U16248 (N_16248,N_13630,N_14208);
or U16249 (N_16249,N_13085,N_14726);
and U16250 (N_16250,N_14367,N_14943);
and U16251 (N_16251,N_13475,N_13087);
and U16252 (N_16252,N_13508,N_14180);
and U16253 (N_16253,N_13899,N_14935);
or U16254 (N_16254,N_13256,N_13455);
and U16255 (N_16255,N_14982,N_12711);
and U16256 (N_16256,N_12671,N_14308);
or U16257 (N_16257,N_14554,N_13306);
nand U16258 (N_16258,N_13202,N_14893);
or U16259 (N_16259,N_14130,N_14227);
and U16260 (N_16260,N_12916,N_14324);
or U16261 (N_16261,N_13873,N_14284);
or U16262 (N_16262,N_14137,N_13435);
nand U16263 (N_16263,N_13114,N_12754);
nand U16264 (N_16264,N_14091,N_13756);
or U16265 (N_16265,N_14666,N_14019);
nand U16266 (N_16266,N_14045,N_14653);
and U16267 (N_16267,N_12614,N_14479);
or U16268 (N_16268,N_12843,N_12559);
nor U16269 (N_16269,N_13414,N_14161);
and U16270 (N_16270,N_12715,N_14729);
nor U16271 (N_16271,N_14528,N_13389);
or U16272 (N_16272,N_13069,N_14027);
nor U16273 (N_16273,N_13231,N_13723);
or U16274 (N_16274,N_13464,N_12957);
xor U16275 (N_16275,N_14349,N_13353);
nand U16276 (N_16276,N_12687,N_14640);
and U16277 (N_16277,N_14437,N_14014);
and U16278 (N_16278,N_13951,N_14674);
and U16279 (N_16279,N_13375,N_12674);
and U16280 (N_16280,N_14080,N_13466);
nand U16281 (N_16281,N_12619,N_13204);
and U16282 (N_16282,N_13128,N_14416);
nand U16283 (N_16283,N_14547,N_14373);
and U16284 (N_16284,N_14107,N_14450);
nor U16285 (N_16285,N_14824,N_13065);
nor U16286 (N_16286,N_14313,N_14895);
nor U16287 (N_16287,N_14956,N_14884);
or U16288 (N_16288,N_14715,N_13750);
and U16289 (N_16289,N_13125,N_12640);
and U16290 (N_16290,N_13159,N_13906);
and U16291 (N_16291,N_13813,N_13747);
nand U16292 (N_16292,N_14712,N_12866);
nor U16293 (N_16293,N_12791,N_13998);
and U16294 (N_16294,N_14087,N_12688);
and U16295 (N_16295,N_12963,N_12575);
or U16296 (N_16296,N_14690,N_12690);
xor U16297 (N_16297,N_13393,N_13004);
or U16298 (N_16298,N_13488,N_14166);
and U16299 (N_16299,N_14600,N_13519);
or U16300 (N_16300,N_14107,N_14596);
and U16301 (N_16301,N_12701,N_14690);
and U16302 (N_16302,N_13257,N_13943);
and U16303 (N_16303,N_12857,N_14123);
nand U16304 (N_16304,N_12750,N_14444);
nand U16305 (N_16305,N_14351,N_14274);
nor U16306 (N_16306,N_13216,N_14267);
nand U16307 (N_16307,N_14372,N_12818);
nor U16308 (N_16308,N_13072,N_12874);
nor U16309 (N_16309,N_13471,N_14247);
nor U16310 (N_16310,N_14832,N_13799);
nand U16311 (N_16311,N_13655,N_13831);
nor U16312 (N_16312,N_14935,N_14491);
nor U16313 (N_16313,N_12864,N_13141);
nand U16314 (N_16314,N_14356,N_12828);
or U16315 (N_16315,N_13724,N_14438);
nor U16316 (N_16316,N_13255,N_14403);
and U16317 (N_16317,N_13388,N_14124);
nor U16318 (N_16318,N_13711,N_12750);
or U16319 (N_16319,N_14845,N_14564);
nand U16320 (N_16320,N_14609,N_14725);
and U16321 (N_16321,N_12608,N_13694);
and U16322 (N_16322,N_14342,N_12609);
nand U16323 (N_16323,N_13288,N_14132);
and U16324 (N_16324,N_13125,N_14930);
nor U16325 (N_16325,N_12564,N_14385);
nor U16326 (N_16326,N_13032,N_13744);
nand U16327 (N_16327,N_12569,N_14871);
or U16328 (N_16328,N_13827,N_12906);
and U16329 (N_16329,N_14957,N_13961);
nor U16330 (N_16330,N_13959,N_14672);
or U16331 (N_16331,N_13767,N_13046);
nand U16332 (N_16332,N_13625,N_13281);
xnor U16333 (N_16333,N_14569,N_14383);
nor U16334 (N_16334,N_13676,N_13241);
nand U16335 (N_16335,N_13156,N_14793);
nor U16336 (N_16336,N_12689,N_14337);
nor U16337 (N_16337,N_12862,N_14909);
and U16338 (N_16338,N_13302,N_12712);
and U16339 (N_16339,N_13700,N_13492);
nor U16340 (N_16340,N_12622,N_14338);
nand U16341 (N_16341,N_12584,N_13967);
nor U16342 (N_16342,N_13584,N_14903);
and U16343 (N_16343,N_12978,N_14812);
or U16344 (N_16344,N_14181,N_14842);
or U16345 (N_16345,N_13695,N_13575);
and U16346 (N_16346,N_14136,N_13177);
and U16347 (N_16347,N_12582,N_13592);
and U16348 (N_16348,N_14403,N_13770);
or U16349 (N_16349,N_14582,N_12686);
nor U16350 (N_16350,N_13458,N_14556);
nor U16351 (N_16351,N_14379,N_13442);
and U16352 (N_16352,N_13248,N_12880);
nor U16353 (N_16353,N_14212,N_12629);
nand U16354 (N_16354,N_12787,N_12832);
or U16355 (N_16355,N_13737,N_13681);
nand U16356 (N_16356,N_13708,N_12966);
nor U16357 (N_16357,N_14580,N_13617);
nor U16358 (N_16358,N_14664,N_13420);
nor U16359 (N_16359,N_13312,N_13347);
or U16360 (N_16360,N_13581,N_12811);
nor U16361 (N_16361,N_14452,N_12824);
xnor U16362 (N_16362,N_13675,N_13553);
nor U16363 (N_16363,N_13775,N_14184);
nand U16364 (N_16364,N_14532,N_14792);
nor U16365 (N_16365,N_14793,N_13682);
and U16366 (N_16366,N_13993,N_13465);
nand U16367 (N_16367,N_13443,N_14427);
and U16368 (N_16368,N_13320,N_14830);
and U16369 (N_16369,N_14132,N_13852);
nand U16370 (N_16370,N_14819,N_13252);
and U16371 (N_16371,N_14885,N_13428);
or U16372 (N_16372,N_13275,N_14398);
nand U16373 (N_16373,N_13203,N_13139);
or U16374 (N_16374,N_14982,N_12825);
and U16375 (N_16375,N_14372,N_13008);
nor U16376 (N_16376,N_14874,N_13260);
and U16377 (N_16377,N_12978,N_14975);
nand U16378 (N_16378,N_12518,N_14910);
and U16379 (N_16379,N_14433,N_12625);
and U16380 (N_16380,N_14106,N_14744);
nor U16381 (N_16381,N_13158,N_13678);
nand U16382 (N_16382,N_13475,N_12939);
nand U16383 (N_16383,N_14887,N_14826);
nor U16384 (N_16384,N_14167,N_12841);
nor U16385 (N_16385,N_12874,N_14774);
or U16386 (N_16386,N_14147,N_14544);
nand U16387 (N_16387,N_14003,N_14482);
nand U16388 (N_16388,N_13990,N_14319);
xnor U16389 (N_16389,N_13102,N_14270);
nor U16390 (N_16390,N_13119,N_14732);
nand U16391 (N_16391,N_13916,N_12831);
nor U16392 (N_16392,N_14400,N_13102);
nand U16393 (N_16393,N_13339,N_13793);
xnor U16394 (N_16394,N_12890,N_12882);
xnor U16395 (N_16395,N_13185,N_12881);
and U16396 (N_16396,N_14700,N_12711);
nor U16397 (N_16397,N_14276,N_12655);
nor U16398 (N_16398,N_13388,N_13826);
xor U16399 (N_16399,N_13199,N_13015);
and U16400 (N_16400,N_14879,N_14198);
and U16401 (N_16401,N_14462,N_13312);
nor U16402 (N_16402,N_14435,N_14966);
nand U16403 (N_16403,N_13909,N_12846);
or U16404 (N_16404,N_12944,N_14111);
nor U16405 (N_16405,N_13072,N_14713);
or U16406 (N_16406,N_13647,N_13075);
and U16407 (N_16407,N_13030,N_13781);
nand U16408 (N_16408,N_14409,N_13464);
nor U16409 (N_16409,N_13704,N_14882);
nand U16410 (N_16410,N_14444,N_14660);
or U16411 (N_16411,N_12827,N_13401);
or U16412 (N_16412,N_13332,N_14113);
nand U16413 (N_16413,N_14368,N_14550);
nand U16414 (N_16414,N_12847,N_14762);
nand U16415 (N_16415,N_14189,N_14556);
and U16416 (N_16416,N_13650,N_14217);
and U16417 (N_16417,N_12697,N_14707);
nand U16418 (N_16418,N_13461,N_13846);
nand U16419 (N_16419,N_14373,N_14458);
nand U16420 (N_16420,N_13805,N_13971);
or U16421 (N_16421,N_14777,N_14356);
and U16422 (N_16422,N_14622,N_13487);
and U16423 (N_16423,N_12524,N_13931);
and U16424 (N_16424,N_13152,N_14345);
and U16425 (N_16425,N_13585,N_14654);
nand U16426 (N_16426,N_13568,N_14440);
and U16427 (N_16427,N_14780,N_14321);
or U16428 (N_16428,N_14896,N_13159);
and U16429 (N_16429,N_13749,N_12674);
and U16430 (N_16430,N_14533,N_13331);
nor U16431 (N_16431,N_14599,N_12963);
xnor U16432 (N_16432,N_14416,N_14692);
or U16433 (N_16433,N_13980,N_12645);
or U16434 (N_16434,N_13461,N_14704);
or U16435 (N_16435,N_14722,N_13291);
nand U16436 (N_16436,N_13359,N_12758);
nor U16437 (N_16437,N_13314,N_14819);
or U16438 (N_16438,N_13210,N_12827);
and U16439 (N_16439,N_14400,N_13057);
or U16440 (N_16440,N_14589,N_14962);
and U16441 (N_16441,N_14758,N_14243);
nand U16442 (N_16442,N_14924,N_14528);
nor U16443 (N_16443,N_13214,N_14576);
nand U16444 (N_16444,N_12669,N_13487);
nand U16445 (N_16445,N_12976,N_12941);
and U16446 (N_16446,N_14598,N_13255);
nand U16447 (N_16447,N_14857,N_12718);
nand U16448 (N_16448,N_14170,N_14903);
nor U16449 (N_16449,N_13558,N_13608);
nand U16450 (N_16450,N_14972,N_13316);
nand U16451 (N_16451,N_12666,N_14690);
nand U16452 (N_16452,N_14074,N_12812);
or U16453 (N_16453,N_13674,N_13233);
or U16454 (N_16454,N_14911,N_14593);
nor U16455 (N_16455,N_14221,N_14363);
nand U16456 (N_16456,N_12828,N_12647);
xor U16457 (N_16457,N_13863,N_13417);
or U16458 (N_16458,N_12899,N_14573);
or U16459 (N_16459,N_14833,N_12723);
nand U16460 (N_16460,N_14596,N_13587);
nor U16461 (N_16461,N_13888,N_14222);
nand U16462 (N_16462,N_13616,N_13843);
or U16463 (N_16463,N_13593,N_13556);
nor U16464 (N_16464,N_13601,N_12761);
or U16465 (N_16465,N_14275,N_12977);
xor U16466 (N_16466,N_14319,N_12501);
and U16467 (N_16467,N_13752,N_14894);
nand U16468 (N_16468,N_13671,N_14994);
nor U16469 (N_16469,N_14911,N_12518);
or U16470 (N_16470,N_14035,N_13809);
nor U16471 (N_16471,N_14792,N_13871);
nor U16472 (N_16472,N_12999,N_14510);
and U16473 (N_16473,N_13891,N_14254);
nand U16474 (N_16474,N_13116,N_13423);
nand U16475 (N_16475,N_13193,N_13800);
nor U16476 (N_16476,N_14595,N_13565);
nand U16477 (N_16477,N_12680,N_14625);
or U16478 (N_16478,N_14582,N_14189);
nor U16479 (N_16479,N_14249,N_13497);
nand U16480 (N_16480,N_13721,N_14351);
nor U16481 (N_16481,N_14059,N_14751);
nor U16482 (N_16482,N_12795,N_12693);
or U16483 (N_16483,N_13179,N_13309);
nand U16484 (N_16484,N_14097,N_13449);
or U16485 (N_16485,N_14888,N_14231);
and U16486 (N_16486,N_14569,N_12631);
nor U16487 (N_16487,N_14569,N_12827);
nor U16488 (N_16488,N_13907,N_14586);
and U16489 (N_16489,N_12827,N_13799);
or U16490 (N_16490,N_14884,N_14784);
nand U16491 (N_16491,N_14088,N_13752);
nor U16492 (N_16492,N_14899,N_13155);
and U16493 (N_16493,N_13779,N_13729);
nand U16494 (N_16494,N_14783,N_13315);
or U16495 (N_16495,N_13466,N_12561);
or U16496 (N_16496,N_13599,N_12841);
nand U16497 (N_16497,N_12749,N_14109);
and U16498 (N_16498,N_13110,N_13345);
and U16499 (N_16499,N_12692,N_14318);
or U16500 (N_16500,N_12779,N_13683);
nor U16501 (N_16501,N_14643,N_12606);
and U16502 (N_16502,N_13060,N_13074);
nand U16503 (N_16503,N_14026,N_14556);
and U16504 (N_16504,N_13006,N_14527);
or U16505 (N_16505,N_13375,N_14774);
nand U16506 (N_16506,N_13094,N_13831);
nor U16507 (N_16507,N_12740,N_14295);
or U16508 (N_16508,N_13211,N_14704);
and U16509 (N_16509,N_13644,N_13298);
nand U16510 (N_16510,N_14680,N_13192);
or U16511 (N_16511,N_14428,N_14253);
nand U16512 (N_16512,N_13312,N_12959);
nand U16513 (N_16513,N_13196,N_14370);
nand U16514 (N_16514,N_13639,N_13808);
nor U16515 (N_16515,N_14300,N_12571);
or U16516 (N_16516,N_12999,N_13823);
nand U16517 (N_16517,N_13398,N_14524);
and U16518 (N_16518,N_13308,N_14814);
nand U16519 (N_16519,N_13277,N_13135);
and U16520 (N_16520,N_13219,N_14841);
nor U16521 (N_16521,N_12745,N_13599);
or U16522 (N_16522,N_14002,N_14703);
or U16523 (N_16523,N_12710,N_12791);
or U16524 (N_16524,N_14271,N_12913);
nand U16525 (N_16525,N_14652,N_12538);
nor U16526 (N_16526,N_14403,N_14834);
or U16527 (N_16527,N_14992,N_12506);
nand U16528 (N_16528,N_12511,N_12941);
or U16529 (N_16529,N_14562,N_14400);
and U16530 (N_16530,N_13764,N_12757);
and U16531 (N_16531,N_13961,N_13908);
or U16532 (N_16532,N_14416,N_14459);
nand U16533 (N_16533,N_13350,N_12988);
or U16534 (N_16534,N_14685,N_13246);
and U16535 (N_16535,N_13168,N_14681);
nand U16536 (N_16536,N_13922,N_13333);
and U16537 (N_16537,N_14713,N_14969);
nor U16538 (N_16538,N_13257,N_13427);
and U16539 (N_16539,N_12693,N_14794);
nor U16540 (N_16540,N_13544,N_14424);
and U16541 (N_16541,N_13129,N_13010);
nor U16542 (N_16542,N_14990,N_14410);
and U16543 (N_16543,N_13916,N_13715);
and U16544 (N_16544,N_14247,N_14497);
or U16545 (N_16545,N_13531,N_13721);
nor U16546 (N_16546,N_14384,N_13718);
nand U16547 (N_16547,N_14559,N_14201);
and U16548 (N_16548,N_14738,N_13592);
nand U16549 (N_16549,N_12615,N_14605);
or U16550 (N_16550,N_13065,N_14341);
or U16551 (N_16551,N_12804,N_14672);
and U16552 (N_16552,N_14455,N_13564);
or U16553 (N_16553,N_13305,N_14050);
and U16554 (N_16554,N_14223,N_12869);
nor U16555 (N_16555,N_14732,N_12905);
nor U16556 (N_16556,N_13424,N_14097);
or U16557 (N_16557,N_12924,N_13117);
and U16558 (N_16558,N_12783,N_14342);
nand U16559 (N_16559,N_12587,N_13433);
and U16560 (N_16560,N_14630,N_12697);
nor U16561 (N_16561,N_12872,N_13650);
nor U16562 (N_16562,N_12549,N_13504);
or U16563 (N_16563,N_13409,N_13467);
and U16564 (N_16564,N_13131,N_13676);
and U16565 (N_16565,N_14337,N_14718);
nand U16566 (N_16566,N_13409,N_13727);
and U16567 (N_16567,N_13769,N_14672);
nor U16568 (N_16568,N_13404,N_14146);
nor U16569 (N_16569,N_14956,N_12695);
or U16570 (N_16570,N_13552,N_13962);
nand U16571 (N_16571,N_12878,N_14698);
or U16572 (N_16572,N_12885,N_13369);
or U16573 (N_16573,N_12590,N_12940);
or U16574 (N_16574,N_13224,N_14909);
nor U16575 (N_16575,N_14840,N_14547);
nor U16576 (N_16576,N_13191,N_12772);
nand U16577 (N_16577,N_13310,N_13090);
or U16578 (N_16578,N_14329,N_14945);
nor U16579 (N_16579,N_14212,N_13195);
nor U16580 (N_16580,N_13406,N_12736);
and U16581 (N_16581,N_14636,N_13032);
or U16582 (N_16582,N_14521,N_12635);
or U16583 (N_16583,N_14733,N_14409);
xor U16584 (N_16584,N_14942,N_12650);
nor U16585 (N_16585,N_14184,N_14359);
and U16586 (N_16586,N_14275,N_14924);
nand U16587 (N_16587,N_14622,N_12818);
nand U16588 (N_16588,N_13093,N_14412);
nor U16589 (N_16589,N_13321,N_13271);
and U16590 (N_16590,N_14303,N_13626);
and U16591 (N_16591,N_13456,N_14093);
nor U16592 (N_16592,N_13902,N_13506);
or U16593 (N_16593,N_13313,N_14856);
nand U16594 (N_16594,N_13172,N_13475);
and U16595 (N_16595,N_13925,N_13950);
and U16596 (N_16596,N_13200,N_13249);
nor U16597 (N_16597,N_14643,N_14836);
nand U16598 (N_16598,N_14895,N_12581);
or U16599 (N_16599,N_14870,N_13138);
nand U16600 (N_16600,N_13716,N_12797);
and U16601 (N_16601,N_14429,N_14098);
nand U16602 (N_16602,N_13175,N_13383);
nand U16603 (N_16603,N_12656,N_13647);
nor U16604 (N_16604,N_13151,N_14356);
nand U16605 (N_16605,N_14435,N_14788);
and U16606 (N_16606,N_12596,N_13527);
nor U16607 (N_16607,N_14828,N_12744);
and U16608 (N_16608,N_12537,N_14470);
nor U16609 (N_16609,N_12681,N_14308);
nor U16610 (N_16610,N_14517,N_14600);
or U16611 (N_16611,N_14300,N_12874);
nand U16612 (N_16612,N_14378,N_13403);
or U16613 (N_16613,N_14686,N_13796);
and U16614 (N_16614,N_12895,N_13200);
and U16615 (N_16615,N_13912,N_13430);
or U16616 (N_16616,N_12940,N_14687);
nor U16617 (N_16617,N_14729,N_14541);
nor U16618 (N_16618,N_14226,N_13429);
nand U16619 (N_16619,N_14790,N_14980);
nor U16620 (N_16620,N_12681,N_14978);
or U16621 (N_16621,N_13027,N_12515);
nor U16622 (N_16622,N_14377,N_13697);
nand U16623 (N_16623,N_14903,N_14552);
and U16624 (N_16624,N_14629,N_13704);
and U16625 (N_16625,N_12516,N_14066);
and U16626 (N_16626,N_14155,N_13933);
nor U16627 (N_16627,N_13000,N_12526);
nand U16628 (N_16628,N_12839,N_13277);
or U16629 (N_16629,N_13044,N_14177);
or U16630 (N_16630,N_13136,N_14182);
nor U16631 (N_16631,N_14534,N_14962);
nand U16632 (N_16632,N_14310,N_13474);
and U16633 (N_16633,N_13898,N_13867);
or U16634 (N_16634,N_14514,N_12963);
xor U16635 (N_16635,N_12965,N_14901);
and U16636 (N_16636,N_14518,N_14968);
nor U16637 (N_16637,N_13020,N_14643);
and U16638 (N_16638,N_13364,N_12552);
nor U16639 (N_16639,N_13584,N_13411);
or U16640 (N_16640,N_12909,N_14746);
and U16641 (N_16641,N_14406,N_14115);
nor U16642 (N_16642,N_14887,N_13057);
nand U16643 (N_16643,N_13087,N_14481);
nand U16644 (N_16644,N_12539,N_12877);
or U16645 (N_16645,N_14991,N_13798);
and U16646 (N_16646,N_14238,N_14232);
or U16647 (N_16647,N_12848,N_14952);
or U16648 (N_16648,N_12599,N_13772);
nor U16649 (N_16649,N_13901,N_12560);
nand U16650 (N_16650,N_14911,N_14118);
and U16651 (N_16651,N_14604,N_13425);
and U16652 (N_16652,N_14178,N_13871);
or U16653 (N_16653,N_12638,N_12927);
and U16654 (N_16654,N_14205,N_13002);
nor U16655 (N_16655,N_14057,N_14194);
nor U16656 (N_16656,N_14174,N_12587);
nand U16657 (N_16657,N_12610,N_13697);
or U16658 (N_16658,N_14989,N_13865);
nor U16659 (N_16659,N_13870,N_14270);
nand U16660 (N_16660,N_12693,N_12993);
or U16661 (N_16661,N_14460,N_14933);
nor U16662 (N_16662,N_12517,N_13356);
nor U16663 (N_16663,N_14681,N_14499);
nor U16664 (N_16664,N_14413,N_13255);
nand U16665 (N_16665,N_13566,N_14463);
nand U16666 (N_16666,N_12884,N_12597);
and U16667 (N_16667,N_14277,N_12873);
and U16668 (N_16668,N_12766,N_13221);
nand U16669 (N_16669,N_14270,N_13519);
nand U16670 (N_16670,N_13979,N_13819);
nor U16671 (N_16671,N_14782,N_13588);
nor U16672 (N_16672,N_13284,N_13574);
and U16673 (N_16673,N_14066,N_13059);
and U16674 (N_16674,N_12705,N_12577);
or U16675 (N_16675,N_14436,N_12801);
or U16676 (N_16676,N_13957,N_13677);
and U16677 (N_16677,N_13154,N_13559);
or U16678 (N_16678,N_13195,N_13699);
or U16679 (N_16679,N_12694,N_14129);
and U16680 (N_16680,N_13500,N_13814);
and U16681 (N_16681,N_12853,N_13608);
or U16682 (N_16682,N_14679,N_13897);
and U16683 (N_16683,N_13956,N_12830);
or U16684 (N_16684,N_14326,N_14874);
or U16685 (N_16685,N_13427,N_12525);
or U16686 (N_16686,N_14796,N_14470);
and U16687 (N_16687,N_13322,N_13197);
and U16688 (N_16688,N_12788,N_12869);
nor U16689 (N_16689,N_13573,N_13670);
xor U16690 (N_16690,N_14863,N_13854);
nor U16691 (N_16691,N_13762,N_14896);
nor U16692 (N_16692,N_14929,N_14476);
and U16693 (N_16693,N_13255,N_14770);
xor U16694 (N_16694,N_13201,N_14884);
and U16695 (N_16695,N_13810,N_14163);
nand U16696 (N_16696,N_12976,N_14746);
nand U16697 (N_16697,N_14433,N_14977);
nand U16698 (N_16698,N_14547,N_13499);
and U16699 (N_16699,N_12827,N_13978);
and U16700 (N_16700,N_13470,N_14159);
nand U16701 (N_16701,N_13854,N_13587);
nand U16702 (N_16702,N_13755,N_13034);
nor U16703 (N_16703,N_14885,N_13097);
or U16704 (N_16704,N_13625,N_13666);
and U16705 (N_16705,N_14441,N_13550);
nand U16706 (N_16706,N_12914,N_13106);
or U16707 (N_16707,N_13471,N_14829);
nand U16708 (N_16708,N_13156,N_12980);
and U16709 (N_16709,N_13922,N_14277);
or U16710 (N_16710,N_13498,N_13990);
nor U16711 (N_16711,N_14915,N_14863);
or U16712 (N_16712,N_14576,N_13174);
and U16713 (N_16713,N_14991,N_12507);
nand U16714 (N_16714,N_14402,N_13852);
nor U16715 (N_16715,N_13094,N_13068);
nor U16716 (N_16716,N_14923,N_14978);
nor U16717 (N_16717,N_14877,N_12555);
nor U16718 (N_16718,N_13215,N_13333);
nand U16719 (N_16719,N_12518,N_14156);
nand U16720 (N_16720,N_13893,N_14882);
or U16721 (N_16721,N_13962,N_14774);
or U16722 (N_16722,N_14194,N_14378);
or U16723 (N_16723,N_14650,N_13594);
nand U16724 (N_16724,N_13513,N_14819);
nor U16725 (N_16725,N_14547,N_14179);
or U16726 (N_16726,N_12887,N_14378);
and U16727 (N_16727,N_12876,N_13158);
or U16728 (N_16728,N_13441,N_14215);
nor U16729 (N_16729,N_14255,N_14793);
nor U16730 (N_16730,N_14044,N_14610);
nor U16731 (N_16731,N_14733,N_13016);
nor U16732 (N_16732,N_12992,N_14493);
or U16733 (N_16733,N_14586,N_13329);
nand U16734 (N_16734,N_13610,N_12892);
nor U16735 (N_16735,N_14543,N_12883);
nand U16736 (N_16736,N_14426,N_12873);
nand U16737 (N_16737,N_13930,N_13319);
or U16738 (N_16738,N_13943,N_13010);
and U16739 (N_16739,N_12685,N_12769);
nand U16740 (N_16740,N_14515,N_13885);
nand U16741 (N_16741,N_13907,N_14747);
and U16742 (N_16742,N_14816,N_14590);
nor U16743 (N_16743,N_14216,N_14870);
or U16744 (N_16744,N_14924,N_14100);
nor U16745 (N_16745,N_13324,N_14698);
or U16746 (N_16746,N_14325,N_12905);
nor U16747 (N_16747,N_14656,N_13579);
nand U16748 (N_16748,N_13647,N_13167);
nand U16749 (N_16749,N_12809,N_14393);
and U16750 (N_16750,N_13902,N_12524);
nand U16751 (N_16751,N_13612,N_13986);
nor U16752 (N_16752,N_13750,N_13568);
nor U16753 (N_16753,N_13168,N_13086);
nor U16754 (N_16754,N_14551,N_13331);
nand U16755 (N_16755,N_12709,N_13479);
nor U16756 (N_16756,N_13615,N_14174);
and U16757 (N_16757,N_13922,N_12696);
nand U16758 (N_16758,N_13758,N_12602);
nand U16759 (N_16759,N_12970,N_13304);
or U16760 (N_16760,N_12699,N_12772);
nor U16761 (N_16761,N_12691,N_14782);
and U16762 (N_16762,N_14392,N_14563);
and U16763 (N_16763,N_13213,N_12990);
nand U16764 (N_16764,N_14156,N_12768);
nor U16765 (N_16765,N_14956,N_13887);
nand U16766 (N_16766,N_13374,N_12592);
or U16767 (N_16767,N_13514,N_12911);
or U16768 (N_16768,N_12659,N_13675);
nor U16769 (N_16769,N_14241,N_12970);
nor U16770 (N_16770,N_14843,N_14437);
or U16771 (N_16771,N_14627,N_12926);
nor U16772 (N_16772,N_13810,N_14472);
and U16773 (N_16773,N_14482,N_13391);
and U16774 (N_16774,N_13830,N_14994);
nor U16775 (N_16775,N_14312,N_13689);
nand U16776 (N_16776,N_14843,N_12526);
nand U16777 (N_16777,N_14499,N_13561);
or U16778 (N_16778,N_12848,N_12611);
or U16779 (N_16779,N_13788,N_13722);
or U16780 (N_16780,N_14578,N_14427);
nor U16781 (N_16781,N_13868,N_13917);
nand U16782 (N_16782,N_12646,N_14037);
nand U16783 (N_16783,N_14594,N_13547);
or U16784 (N_16784,N_12683,N_13298);
nor U16785 (N_16785,N_14415,N_14172);
nand U16786 (N_16786,N_12985,N_14080);
nor U16787 (N_16787,N_14169,N_12800);
nor U16788 (N_16788,N_14560,N_14872);
nor U16789 (N_16789,N_12886,N_14658);
and U16790 (N_16790,N_14605,N_13490);
or U16791 (N_16791,N_14117,N_13555);
nor U16792 (N_16792,N_14093,N_14867);
nor U16793 (N_16793,N_12940,N_13209);
or U16794 (N_16794,N_12957,N_13941);
and U16795 (N_16795,N_13623,N_13554);
nand U16796 (N_16796,N_13015,N_13557);
nor U16797 (N_16797,N_14416,N_13199);
and U16798 (N_16798,N_14756,N_14470);
and U16799 (N_16799,N_13826,N_13340);
or U16800 (N_16800,N_13024,N_12566);
or U16801 (N_16801,N_14090,N_13919);
or U16802 (N_16802,N_12942,N_14369);
nor U16803 (N_16803,N_14806,N_14186);
or U16804 (N_16804,N_14276,N_12804);
nor U16805 (N_16805,N_14963,N_14382);
nor U16806 (N_16806,N_14835,N_13311);
nor U16807 (N_16807,N_13717,N_14629);
nor U16808 (N_16808,N_13801,N_13381);
nand U16809 (N_16809,N_14407,N_12589);
or U16810 (N_16810,N_14351,N_13844);
nand U16811 (N_16811,N_14076,N_12762);
nor U16812 (N_16812,N_13807,N_14263);
nor U16813 (N_16813,N_14078,N_13775);
nor U16814 (N_16814,N_13116,N_14345);
and U16815 (N_16815,N_12769,N_12791);
and U16816 (N_16816,N_12833,N_13323);
nand U16817 (N_16817,N_13881,N_14732);
nand U16818 (N_16818,N_14624,N_12879);
nor U16819 (N_16819,N_12997,N_13328);
and U16820 (N_16820,N_13732,N_14433);
or U16821 (N_16821,N_14904,N_14162);
or U16822 (N_16822,N_13027,N_12860);
or U16823 (N_16823,N_12533,N_12570);
nand U16824 (N_16824,N_14453,N_13046);
nor U16825 (N_16825,N_14236,N_13521);
nand U16826 (N_16826,N_13914,N_13668);
or U16827 (N_16827,N_12542,N_13008);
nor U16828 (N_16828,N_12561,N_13938);
or U16829 (N_16829,N_14985,N_12557);
or U16830 (N_16830,N_13072,N_14552);
and U16831 (N_16831,N_12824,N_12555);
nor U16832 (N_16832,N_13800,N_14773);
and U16833 (N_16833,N_14597,N_13270);
and U16834 (N_16834,N_13422,N_13281);
nor U16835 (N_16835,N_14305,N_13351);
or U16836 (N_16836,N_13859,N_14190);
nor U16837 (N_16837,N_13507,N_13516);
and U16838 (N_16838,N_13662,N_13498);
and U16839 (N_16839,N_14527,N_12934);
or U16840 (N_16840,N_12611,N_14403);
and U16841 (N_16841,N_12700,N_13589);
nand U16842 (N_16842,N_12966,N_13898);
nor U16843 (N_16843,N_13479,N_13881);
or U16844 (N_16844,N_14557,N_13946);
nand U16845 (N_16845,N_14936,N_13807);
nor U16846 (N_16846,N_14588,N_14296);
nand U16847 (N_16847,N_12935,N_14321);
or U16848 (N_16848,N_14358,N_14153);
and U16849 (N_16849,N_14797,N_13159);
or U16850 (N_16850,N_12550,N_12613);
nand U16851 (N_16851,N_13229,N_12596);
or U16852 (N_16852,N_13103,N_12733);
nor U16853 (N_16853,N_13479,N_13801);
or U16854 (N_16854,N_14298,N_14551);
or U16855 (N_16855,N_14898,N_14495);
or U16856 (N_16856,N_14983,N_12891);
and U16857 (N_16857,N_13183,N_13341);
or U16858 (N_16858,N_13752,N_14920);
and U16859 (N_16859,N_14359,N_14663);
and U16860 (N_16860,N_13142,N_12674);
or U16861 (N_16861,N_14437,N_14121);
and U16862 (N_16862,N_12994,N_13052);
or U16863 (N_16863,N_14001,N_13663);
or U16864 (N_16864,N_12719,N_14465);
nor U16865 (N_16865,N_13271,N_14835);
and U16866 (N_16866,N_12502,N_13587);
and U16867 (N_16867,N_13887,N_14332);
nor U16868 (N_16868,N_14956,N_14541);
nor U16869 (N_16869,N_12885,N_13163);
nor U16870 (N_16870,N_12729,N_12623);
nand U16871 (N_16871,N_13968,N_14539);
nor U16872 (N_16872,N_14584,N_14226);
nand U16873 (N_16873,N_13110,N_13417);
and U16874 (N_16874,N_13615,N_12984);
nand U16875 (N_16875,N_14415,N_13967);
and U16876 (N_16876,N_13724,N_13091);
nor U16877 (N_16877,N_14448,N_13869);
nor U16878 (N_16878,N_14186,N_14779);
or U16879 (N_16879,N_14906,N_14859);
or U16880 (N_16880,N_14156,N_14327);
and U16881 (N_16881,N_12529,N_13770);
nand U16882 (N_16882,N_14376,N_13222);
nand U16883 (N_16883,N_14429,N_13913);
nor U16884 (N_16884,N_12681,N_12807);
or U16885 (N_16885,N_14645,N_13544);
and U16886 (N_16886,N_13917,N_14176);
or U16887 (N_16887,N_14788,N_14907);
and U16888 (N_16888,N_14333,N_14851);
or U16889 (N_16889,N_13523,N_14531);
nand U16890 (N_16890,N_14210,N_13303);
and U16891 (N_16891,N_12834,N_14506);
nor U16892 (N_16892,N_13120,N_12967);
nor U16893 (N_16893,N_14121,N_13310);
nand U16894 (N_16894,N_12510,N_13471);
or U16895 (N_16895,N_14066,N_14470);
nor U16896 (N_16896,N_13495,N_13606);
nand U16897 (N_16897,N_14497,N_12735);
nor U16898 (N_16898,N_14599,N_14498);
nand U16899 (N_16899,N_14897,N_13830);
nor U16900 (N_16900,N_14490,N_14579);
and U16901 (N_16901,N_13783,N_13636);
or U16902 (N_16902,N_13191,N_12605);
nor U16903 (N_16903,N_13667,N_14821);
nor U16904 (N_16904,N_12602,N_13648);
nor U16905 (N_16905,N_14535,N_14589);
or U16906 (N_16906,N_13637,N_12812);
and U16907 (N_16907,N_13252,N_12970);
nand U16908 (N_16908,N_12572,N_13863);
and U16909 (N_16909,N_14077,N_14806);
or U16910 (N_16910,N_14929,N_14510);
and U16911 (N_16911,N_12761,N_14972);
nand U16912 (N_16912,N_14624,N_14967);
and U16913 (N_16913,N_14819,N_13243);
or U16914 (N_16914,N_14810,N_13801);
nor U16915 (N_16915,N_13470,N_13044);
and U16916 (N_16916,N_14705,N_14392);
and U16917 (N_16917,N_14210,N_13315);
and U16918 (N_16918,N_12807,N_14863);
nand U16919 (N_16919,N_12712,N_12809);
and U16920 (N_16920,N_14827,N_13440);
nor U16921 (N_16921,N_12892,N_14738);
xor U16922 (N_16922,N_14595,N_13974);
nand U16923 (N_16923,N_14563,N_13113);
nand U16924 (N_16924,N_14576,N_13507);
and U16925 (N_16925,N_13253,N_12541);
nand U16926 (N_16926,N_12926,N_14991);
nor U16927 (N_16927,N_12583,N_13225);
and U16928 (N_16928,N_14689,N_13583);
nor U16929 (N_16929,N_13117,N_14059);
nand U16930 (N_16930,N_12638,N_12500);
or U16931 (N_16931,N_14996,N_14384);
and U16932 (N_16932,N_14728,N_14926);
or U16933 (N_16933,N_12977,N_14056);
or U16934 (N_16934,N_14874,N_14722);
and U16935 (N_16935,N_14409,N_12933);
nor U16936 (N_16936,N_14575,N_13899);
nand U16937 (N_16937,N_13962,N_13630);
or U16938 (N_16938,N_13558,N_12580);
and U16939 (N_16939,N_14961,N_13824);
and U16940 (N_16940,N_13083,N_14628);
nand U16941 (N_16941,N_14573,N_14028);
nor U16942 (N_16942,N_12890,N_13699);
and U16943 (N_16943,N_13002,N_13854);
or U16944 (N_16944,N_12777,N_14189);
nor U16945 (N_16945,N_14041,N_13564);
nor U16946 (N_16946,N_14300,N_13128);
or U16947 (N_16947,N_12755,N_13109);
nor U16948 (N_16948,N_14051,N_13149);
or U16949 (N_16949,N_13785,N_13271);
xnor U16950 (N_16950,N_13063,N_13662);
or U16951 (N_16951,N_13984,N_14304);
or U16952 (N_16952,N_14190,N_13089);
nor U16953 (N_16953,N_14215,N_13802);
nor U16954 (N_16954,N_12660,N_13635);
and U16955 (N_16955,N_12582,N_14249);
and U16956 (N_16956,N_14604,N_13258);
nand U16957 (N_16957,N_14868,N_13799);
and U16958 (N_16958,N_13061,N_13170);
nand U16959 (N_16959,N_14917,N_14407);
nand U16960 (N_16960,N_12601,N_12510);
nand U16961 (N_16961,N_12869,N_14383);
nor U16962 (N_16962,N_14031,N_12536);
and U16963 (N_16963,N_14913,N_14225);
and U16964 (N_16964,N_13962,N_12975);
nor U16965 (N_16965,N_14565,N_14166);
nor U16966 (N_16966,N_12637,N_14417);
nor U16967 (N_16967,N_14615,N_13910);
or U16968 (N_16968,N_14529,N_13024);
nor U16969 (N_16969,N_14191,N_14671);
and U16970 (N_16970,N_14192,N_14994);
or U16971 (N_16971,N_14594,N_12535);
nor U16972 (N_16972,N_13350,N_14944);
and U16973 (N_16973,N_14046,N_14399);
nor U16974 (N_16974,N_13245,N_14574);
nor U16975 (N_16975,N_13865,N_14034);
nor U16976 (N_16976,N_13272,N_14024);
nor U16977 (N_16977,N_13933,N_14943);
or U16978 (N_16978,N_13265,N_13911);
or U16979 (N_16979,N_12550,N_14926);
nor U16980 (N_16980,N_13410,N_13224);
nand U16981 (N_16981,N_14782,N_13611);
nor U16982 (N_16982,N_12794,N_14399);
or U16983 (N_16983,N_13326,N_13447);
nand U16984 (N_16984,N_14180,N_13718);
and U16985 (N_16985,N_13467,N_13679);
or U16986 (N_16986,N_14672,N_13652);
or U16987 (N_16987,N_13560,N_14937);
nor U16988 (N_16988,N_14817,N_13186);
and U16989 (N_16989,N_12767,N_13358);
or U16990 (N_16990,N_12738,N_13792);
nor U16991 (N_16991,N_13289,N_13014);
nand U16992 (N_16992,N_13956,N_14609);
nand U16993 (N_16993,N_14083,N_12832);
or U16994 (N_16994,N_13903,N_14738);
or U16995 (N_16995,N_13668,N_12976);
or U16996 (N_16996,N_14437,N_14732);
nor U16997 (N_16997,N_14219,N_14369);
and U16998 (N_16998,N_12777,N_13710);
and U16999 (N_16999,N_13656,N_14897);
nor U17000 (N_17000,N_13924,N_13059);
nand U17001 (N_17001,N_14355,N_12547);
or U17002 (N_17002,N_12784,N_14700);
nand U17003 (N_17003,N_14943,N_12567);
and U17004 (N_17004,N_14785,N_13682);
and U17005 (N_17005,N_14825,N_13267);
nand U17006 (N_17006,N_14687,N_14427);
nor U17007 (N_17007,N_12523,N_14051);
or U17008 (N_17008,N_12573,N_14308);
nor U17009 (N_17009,N_13622,N_12763);
or U17010 (N_17010,N_14621,N_14857);
nand U17011 (N_17011,N_13358,N_14524);
or U17012 (N_17012,N_13639,N_14916);
nand U17013 (N_17013,N_13765,N_13936);
nor U17014 (N_17014,N_13701,N_12713);
and U17015 (N_17015,N_13089,N_14627);
nand U17016 (N_17016,N_14442,N_14198);
nand U17017 (N_17017,N_14992,N_14797);
xnor U17018 (N_17018,N_12850,N_14402);
or U17019 (N_17019,N_13049,N_14384);
nor U17020 (N_17020,N_12710,N_13836);
or U17021 (N_17021,N_12630,N_14359);
or U17022 (N_17022,N_12641,N_14906);
nor U17023 (N_17023,N_12686,N_13261);
and U17024 (N_17024,N_13352,N_14253);
xor U17025 (N_17025,N_12862,N_12840);
nand U17026 (N_17026,N_14753,N_14037);
or U17027 (N_17027,N_12996,N_13892);
or U17028 (N_17028,N_14294,N_14586);
or U17029 (N_17029,N_14175,N_13883);
nand U17030 (N_17030,N_14071,N_14009);
nor U17031 (N_17031,N_14640,N_13906);
nand U17032 (N_17032,N_13007,N_14006);
and U17033 (N_17033,N_12790,N_13834);
nand U17034 (N_17034,N_14100,N_13561);
or U17035 (N_17035,N_13306,N_12970);
nand U17036 (N_17036,N_14226,N_12705);
nor U17037 (N_17037,N_14198,N_14047);
or U17038 (N_17038,N_14391,N_13572);
nand U17039 (N_17039,N_13758,N_12998);
and U17040 (N_17040,N_14413,N_14313);
nor U17041 (N_17041,N_14386,N_14663);
nor U17042 (N_17042,N_13439,N_13597);
nand U17043 (N_17043,N_13017,N_14670);
or U17044 (N_17044,N_14588,N_13208);
nor U17045 (N_17045,N_13326,N_12639);
or U17046 (N_17046,N_14120,N_13163);
nand U17047 (N_17047,N_13543,N_14525);
nand U17048 (N_17048,N_12918,N_14853);
or U17049 (N_17049,N_13859,N_12743);
nor U17050 (N_17050,N_14169,N_13836);
or U17051 (N_17051,N_13692,N_12502);
and U17052 (N_17052,N_14150,N_14478);
nor U17053 (N_17053,N_13093,N_12851);
and U17054 (N_17054,N_13747,N_12834);
or U17055 (N_17055,N_14008,N_14583);
or U17056 (N_17056,N_13986,N_13789);
and U17057 (N_17057,N_13538,N_12931);
and U17058 (N_17058,N_12688,N_12944);
or U17059 (N_17059,N_12601,N_14746);
and U17060 (N_17060,N_14064,N_14093);
nor U17061 (N_17061,N_13908,N_14933);
nand U17062 (N_17062,N_14175,N_14331);
nor U17063 (N_17063,N_13101,N_14752);
nand U17064 (N_17064,N_14260,N_14031);
and U17065 (N_17065,N_13474,N_14071);
and U17066 (N_17066,N_13101,N_13998);
nand U17067 (N_17067,N_14244,N_13179);
nand U17068 (N_17068,N_14984,N_13909);
and U17069 (N_17069,N_13221,N_13543);
or U17070 (N_17070,N_14264,N_14866);
and U17071 (N_17071,N_12864,N_12882);
or U17072 (N_17072,N_14620,N_14639);
and U17073 (N_17073,N_13466,N_12701);
nor U17074 (N_17074,N_14823,N_14034);
and U17075 (N_17075,N_14807,N_13023);
or U17076 (N_17076,N_13122,N_14385);
nor U17077 (N_17077,N_13878,N_14948);
nor U17078 (N_17078,N_12619,N_14017);
nor U17079 (N_17079,N_14394,N_12524);
nand U17080 (N_17080,N_13270,N_14078);
nand U17081 (N_17081,N_12506,N_14245);
nand U17082 (N_17082,N_14526,N_13920);
or U17083 (N_17083,N_12830,N_13114);
or U17084 (N_17084,N_13935,N_12723);
or U17085 (N_17085,N_12939,N_13451);
nor U17086 (N_17086,N_12847,N_13193);
and U17087 (N_17087,N_13776,N_14835);
nor U17088 (N_17088,N_14588,N_13963);
or U17089 (N_17089,N_12778,N_13959);
and U17090 (N_17090,N_14628,N_12620);
and U17091 (N_17091,N_13111,N_14507);
xnor U17092 (N_17092,N_14767,N_14762);
or U17093 (N_17093,N_13423,N_13970);
nor U17094 (N_17094,N_13651,N_13584);
nor U17095 (N_17095,N_13897,N_12905);
nand U17096 (N_17096,N_14327,N_14301);
and U17097 (N_17097,N_13493,N_12863);
nor U17098 (N_17098,N_13978,N_13594);
or U17099 (N_17099,N_13702,N_12634);
and U17100 (N_17100,N_12999,N_13231);
and U17101 (N_17101,N_14293,N_13173);
nor U17102 (N_17102,N_14206,N_14167);
or U17103 (N_17103,N_12733,N_14883);
nand U17104 (N_17104,N_13068,N_13747);
and U17105 (N_17105,N_14801,N_14975);
and U17106 (N_17106,N_14701,N_13414);
nand U17107 (N_17107,N_13585,N_12561);
and U17108 (N_17108,N_14948,N_13163);
nand U17109 (N_17109,N_14224,N_12999);
or U17110 (N_17110,N_13493,N_13376);
nor U17111 (N_17111,N_12940,N_14311);
nor U17112 (N_17112,N_14129,N_12778);
and U17113 (N_17113,N_13002,N_12791);
or U17114 (N_17114,N_14401,N_14527);
nor U17115 (N_17115,N_13426,N_14891);
nand U17116 (N_17116,N_12624,N_13758);
or U17117 (N_17117,N_12567,N_13433);
nor U17118 (N_17118,N_14269,N_13279);
nand U17119 (N_17119,N_12871,N_13354);
nand U17120 (N_17120,N_13245,N_13791);
and U17121 (N_17121,N_12695,N_13266);
or U17122 (N_17122,N_13400,N_13837);
nand U17123 (N_17123,N_12857,N_12509);
and U17124 (N_17124,N_13913,N_14093);
nand U17125 (N_17125,N_14267,N_13000);
nor U17126 (N_17126,N_14430,N_13972);
nand U17127 (N_17127,N_14645,N_13869);
nand U17128 (N_17128,N_14187,N_13689);
or U17129 (N_17129,N_13611,N_12807);
nor U17130 (N_17130,N_14039,N_13296);
or U17131 (N_17131,N_13138,N_13008);
nand U17132 (N_17132,N_14221,N_14718);
or U17133 (N_17133,N_13119,N_13772);
or U17134 (N_17134,N_14298,N_13529);
nand U17135 (N_17135,N_14806,N_14786);
nand U17136 (N_17136,N_13057,N_13757);
nor U17137 (N_17137,N_13701,N_12617);
nand U17138 (N_17138,N_14106,N_12619);
nor U17139 (N_17139,N_14333,N_13893);
or U17140 (N_17140,N_14990,N_14220);
nand U17141 (N_17141,N_13540,N_13498);
and U17142 (N_17142,N_13470,N_13881);
nor U17143 (N_17143,N_13198,N_13045);
nor U17144 (N_17144,N_12862,N_14721);
nor U17145 (N_17145,N_14519,N_14923);
or U17146 (N_17146,N_14982,N_14170);
or U17147 (N_17147,N_14361,N_14967);
nor U17148 (N_17148,N_14054,N_14502);
or U17149 (N_17149,N_13398,N_14170);
nand U17150 (N_17150,N_13054,N_14128);
nand U17151 (N_17151,N_14412,N_12607);
or U17152 (N_17152,N_14493,N_13201);
and U17153 (N_17153,N_14415,N_12866);
and U17154 (N_17154,N_14853,N_12667);
or U17155 (N_17155,N_13081,N_13543);
and U17156 (N_17156,N_13393,N_13581);
and U17157 (N_17157,N_13230,N_12671);
or U17158 (N_17158,N_13157,N_14147);
or U17159 (N_17159,N_14997,N_12776);
nor U17160 (N_17160,N_12757,N_13252);
nand U17161 (N_17161,N_14230,N_13019);
or U17162 (N_17162,N_14034,N_12799);
nand U17163 (N_17163,N_14555,N_13295);
nand U17164 (N_17164,N_13007,N_13829);
nor U17165 (N_17165,N_13878,N_12785);
nand U17166 (N_17166,N_14341,N_13337);
nand U17167 (N_17167,N_12654,N_14420);
nor U17168 (N_17168,N_12660,N_12801);
nand U17169 (N_17169,N_13144,N_12554);
or U17170 (N_17170,N_12873,N_13962);
or U17171 (N_17171,N_14038,N_14536);
nor U17172 (N_17172,N_14132,N_13757);
and U17173 (N_17173,N_14032,N_13463);
xor U17174 (N_17174,N_14438,N_13279);
or U17175 (N_17175,N_14296,N_14708);
nand U17176 (N_17176,N_13885,N_14720);
nor U17177 (N_17177,N_14372,N_13391);
nand U17178 (N_17178,N_14708,N_13367);
nor U17179 (N_17179,N_14711,N_13780);
nand U17180 (N_17180,N_13495,N_12904);
and U17181 (N_17181,N_12742,N_14298);
or U17182 (N_17182,N_14108,N_13757);
nor U17183 (N_17183,N_14423,N_14336);
nor U17184 (N_17184,N_13096,N_13163);
nand U17185 (N_17185,N_14093,N_14104);
nor U17186 (N_17186,N_14390,N_14186);
nand U17187 (N_17187,N_13191,N_13483);
or U17188 (N_17188,N_14130,N_14895);
and U17189 (N_17189,N_14544,N_14388);
nand U17190 (N_17190,N_14366,N_13483);
nor U17191 (N_17191,N_12963,N_13391);
or U17192 (N_17192,N_14363,N_12555);
nand U17193 (N_17193,N_14265,N_14396);
or U17194 (N_17194,N_13702,N_13140);
or U17195 (N_17195,N_13841,N_13601);
or U17196 (N_17196,N_14258,N_14886);
and U17197 (N_17197,N_13488,N_12558);
and U17198 (N_17198,N_14988,N_13732);
nand U17199 (N_17199,N_14902,N_14377);
or U17200 (N_17200,N_13733,N_13322);
nor U17201 (N_17201,N_13762,N_14472);
and U17202 (N_17202,N_14575,N_14905);
nand U17203 (N_17203,N_13674,N_14734);
nand U17204 (N_17204,N_13978,N_12949);
nor U17205 (N_17205,N_14135,N_14821);
or U17206 (N_17206,N_13893,N_13468);
nor U17207 (N_17207,N_12826,N_14981);
or U17208 (N_17208,N_14208,N_12834);
or U17209 (N_17209,N_13201,N_14013);
nor U17210 (N_17210,N_14705,N_12750);
or U17211 (N_17211,N_14715,N_13734);
nand U17212 (N_17212,N_13756,N_13358);
or U17213 (N_17213,N_13784,N_13115);
xnor U17214 (N_17214,N_12987,N_12960);
nand U17215 (N_17215,N_13888,N_14328);
nand U17216 (N_17216,N_14869,N_14230);
or U17217 (N_17217,N_12777,N_13039);
nor U17218 (N_17218,N_13559,N_14601);
nor U17219 (N_17219,N_14345,N_14254);
and U17220 (N_17220,N_14215,N_12675);
and U17221 (N_17221,N_14504,N_14973);
or U17222 (N_17222,N_12889,N_14143);
or U17223 (N_17223,N_14069,N_13010);
or U17224 (N_17224,N_14024,N_12810);
nand U17225 (N_17225,N_14818,N_13942);
nor U17226 (N_17226,N_14227,N_13502);
nor U17227 (N_17227,N_13972,N_14088);
or U17228 (N_17228,N_13958,N_12524);
nand U17229 (N_17229,N_14748,N_12854);
nor U17230 (N_17230,N_12893,N_13110);
or U17231 (N_17231,N_13090,N_14002);
and U17232 (N_17232,N_13296,N_12863);
nand U17233 (N_17233,N_12956,N_13769);
or U17234 (N_17234,N_13796,N_12755);
or U17235 (N_17235,N_13754,N_14080);
nand U17236 (N_17236,N_13916,N_14072);
nor U17237 (N_17237,N_12563,N_13943);
or U17238 (N_17238,N_13070,N_14194);
nand U17239 (N_17239,N_13038,N_14994);
nand U17240 (N_17240,N_12659,N_14310);
xor U17241 (N_17241,N_14738,N_13754);
or U17242 (N_17242,N_12969,N_14414);
or U17243 (N_17243,N_13708,N_13751);
nor U17244 (N_17244,N_13852,N_12525);
or U17245 (N_17245,N_13019,N_12630);
nand U17246 (N_17246,N_14813,N_12653);
or U17247 (N_17247,N_13238,N_12595);
and U17248 (N_17248,N_14822,N_13565);
nor U17249 (N_17249,N_14275,N_13463);
nor U17250 (N_17250,N_14765,N_14221);
and U17251 (N_17251,N_12549,N_14622);
and U17252 (N_17252,N_13273,N_14015);
or U17253 (N_17253,N_12707,N_12774);
nand U17254 (N_17254,N_14148,N_14397);
or U17255 (N_17255,N_14607,N_14496);
and U17256 (N_17256,N_14793,N_14477);
or U17257 (N_17257,N_13899,N_14310);
nand U17258 (N_17258,N_13536,N_14212);
nor U17259 (N_17259,N_13130,N_14378);
nand U17260 (N_17260,N_14012,N_14982);
nor U17261 (N_17261,N_14249,N_12740);
and U17262 (N_17262,N_14622,N_14758);
nand U17263 (N_17263,N_14750,N_14992);
nand U17264 (N_17264,N_13165,N_13540);
and U17265 (N_17265,N_13681,N_14184);
or U17266 (N_17266,N_12989,N_14478);
nand U17267 (N_17267,N_13596,N_14026);
and U17268 (N_17268,N_14651,N_12613);
and U17269 (N_17269,N_13529,N_13703);
nand U17270 (N_17270,N_12728,N_14818);
nand U17271 (N_17271,N_13169,N_13632);
and U17272 (N_17272,N_13564,N_14970);
or U17273 (N_17273,N_14427,N_14112);
nand U17274 (N_17274,N_13512,N_14818);
nor U17275 (N_17275,N_13070,N_12559);
or U17276 (N_17276,N_14912,N_13964);
nor U17277 (N_17277,N_13232,N_13131);
or U17278 (N_17278,N_13083,N_12854);
nor U17279 (N_17279,N_12852,N_14535);
nor U17280 (N_17280,N_14710,N_14103);
nand U17281 (N_17281,N_14609,N_13320);
and U17282 (N_17282,N_13309,N_14764);
or U17283 (N_17283,N_13153,N_13406);
nor U17284 (N_17284,N_13848,N_12725);
xor U17285 (N_17285,N_14247,N_14753);
or U17286 (N_17286,N_14519,N_13163);
or U17287 (N_17287,N_12900,N_12958);
nor U17288 (N_17288,N_13199,N_13291);
nor U17289 (N_17289,N_14936,N_12660);
nor U17290 (N_17290,N_13348,N_13587);
or U17291 (N_17291,N_13538,N_12587);
xnor U17292 (N_17292,N_14453,N_14108);
nand U17293 (N_17293,N_14217,N_14321);
and U17294 (N_17294,N_14431,N_14245);
or U17295 (N_17295,N_14166,N_13071);
nor U17296 (N_17296,N_12834,N_14441);
nand U17297 (N_17297,N_13839,N_13825);
and U17298 (N_17298,N_13527,N_13856);
or U17299 (N_17299,N_13191,N_12680);
and U17300 (N_17300,N_12597,N_14701);
or U17301 (N_17301,N_12602,N_13941);
nor U17302 (N_17302,N_13764,N_13799);
and U17303 (N_17303,N_13006,N_13787);
nand U17304 (N_17304,N_13239,N_12913);
and U17305 (N_17305,N_13160,N_14195);
nor U17306 (N_17306,N_13949,N_13222);
and U17307 (N_17307,N_14633,N_13645);
nor U17308 (N_17308,N_13877,N_14762);
and U17309 (N_17309,N_13237,N_12928);
or U17310 (N_17310,N_14103,N_14123);
nand U17311 (N_17311,N_13756,N_13013);
nor U17312 (N_17312,N_12538,N_14357);
nor U17313 (N_17313,N_12800,N_12916);
or U17314 (N_17314,N_12857,N_14831);
and U17315 (N_17315,N_12727,N_12533);
and U17316 (N_17316,N_13065,N_13280);
nand U17317 (N_17317,N_14255,N_13060);
nor U17318 (N_17318,N_14257,N_13836);
nor U17319 (N_17319,N_12972,N_14156);
nand U17320 (N_17320,N_13273,N_13419);
nand U17321 (N_17321,N_12695,N_13125);
and U17322 (N_17322,N_14641,N_14195);
and U17323 (N_17323,N_13728,N_13361);
xor U17324 (N_17324,N_13037,N_13652);
and U17325 (N_17325,N_12571,N_12632);
nand U17326 (N_17326,N_13493,N_14714);
nor U17327 (N_17327,N_14769,N_12937);
nand U17328 (N_17328,N_13179,N_14505);
nor U17329 (N_17329,N_14297,N_13677);
and U17330 (N_17330,N_14795,N_14307);
nor U17331 (N_17331,N_13613,N_14489);
nand U17332 (N_17332,N_14282,N_13750);
nand U17333 (N_17333,N_14710,N_13711);
or U17334 (N_17334,N_14919,N_14288);
and U17335 (N_17335,N_13513,N_13360);
or U17336 (N_17336,N_14305,N_14585);
nand U17337 (N_17337,N_13790,N_14722);
or U17338 (N_17338,N_13871,N_13990);
nor U17339 (N_17339,N_13178,N_13314);
and U17340 (N_17340,N_13600,N_14962);
nor U17341 (N_17341,N_13745,N_14930);
nand U17342 (N_17342,N_13771,N_14706);
nor U17343 (N_17343,N_12768,N_13549);
and U17344 (N_17344,N_13339,N_14015);
nand U17345 (N_17345,N_12635,N_12755);
and U17346 (N_17346,N_14801,N_12698);
and U17347 (N_17347,N_14228,N_12944);
and U17348 (N_17348,N_12705,N_14892);
nor U17349 (N_17349,N_14070,N_14459);
or U17350 (N_17350,N_13891,N_13759);
or U17351 (N_17351,N_12937,N_14143);
or U17352 (N_17352,N_12746,N_14263);
nand U17353 (N_17353,N_12791,N_14759);
nand U17354 (N_17354,N_13758,N_13188);
nor U17355 (N_17355,N_13831,N_13935);
or U17356 (N_17356,N_14101,N_14578);
or U17357 (N_17357,N_14220,N_14236);
nand U17358 (N_17358,N_12894,N_14179);
nor U17359 (N_17359,N_13393,N_14707);
and U17360 (N_17360,N_12781,N_14890);
or U17361 (N_17361,N_12501,N_14411);
or U17362 (N_17362,N_14266,N_14192);
nand U17363 (N_17363,N_12860,N_12761);
nor U17364 (N_17364,N_12608,N_14602);
nand U17365 (N_17365,N_13917,N_13883);
or U17366 (N_17366,N_13033,N_13659);
nand U17367 (N_17367,N_12919,N_13304);
and U17368 (N_17368,N_14062,N_13276);
or U17369 (N_17369,N_13967,N_12955);
and U17370 (N_17370,N_13723,N_14568);
and U17371 (N_17371,N_14570,N_14431);
or U17372 (N_17372,N_13810,N_14262);
or U17373 (N_17373,N_14093,N_14879);
nand U17374 (N_17374,N_13939,N_13953);
nor U17375 (N_17375,N_13165,N_14860);
or U17376 (N_17376,N_12707,N_14153);
and U17377 (N_17377,N_12932,N_13678);
nand U17378 (N_17378,N_13807,N_14023);
nand U17379 (N_17379,N_14156,N_13707);
and U17380 (N_17380,N_14799,N_12724);
nand U17381 (N_17381,N_13783,N_14486);
nor U17382 (N_17382,N_14281,N_14493);
nand U17383 (N_17383,N_14904,N_14972);
nor U17384 (N_17384,N_14589,N_14627);
and U17385 (N_17385,N_13832,N_14314);
and U17386 (N_17386,N_14330,N_14837);
or U17387 (N_17387,N_13454,N_13483);
nor U17388 (N_17388,N_13793,N_12953);
nor U17389 (N_17389,N_14063,N_14628);
or U17390 (N_17390,N_13190,N_13897);
nand U17391 (N_17391,N_13091,N_14715);
nand U17392 (N_17392,N_13112,N_14144);
and U17393 (N_17393,N_14180,N_12947);
and U17394 (N_17394,N_14624,N_14594);
nand U17395 (N_17395,N_14537,N_13739);
and U17396 (N_17396,N_13979,N_14391);
xor U17397 (N_17397,N_14280,N_14379);
and U17398 (N_17398,N_13538,N_12760);
and U17399 (N_17399,N_14488,N_13345);
and U17400 (N_17400,N_13463,N_13734);
nor U17401 (N_17401,N_12936,N_13486);
nor U17402 (N_17402,N_13984,N_14755);
nor U17403 (N_17403,N_14560,N_12951);
or U17404 (N_17404,N_14314,N_14596);
nor U17405 (N_17405,N_13398,N_14878);
or U17406 (N_17406,N_14010,N_14249);
nor U17407 (N_17407,N_12855,N_14720);
nor U17408 (N_17408,N_14287,N_13756);
nand U17409 (N_17409,N_13424,N_13009);
or U17410 (N_17410,N_13879,N_13790);
nand U17411 (N_17411,N_12802,N_13127);
and U17412 (N_17412,N_14631,N_13232);
and U17413 (N_17413,N_14982,N_14328);
nand U17414 (N_17414,N_14382,N_14298);
xor U17415 (N_17415,N_14028,N_14213);
or U17416 (N_17416,N_12988,N_14703);
nand U17417 (N_17417,N_14199,N_14812);
nand U17418 (N_17418,N_13134,N_13435);
nand U17419 (N_17419,N_14850,N_12725);
and U17420 (N_17420,N_14171,N_14685);
nor U17421 (N_17421,N_14971,N_14411);
and U17422 (N_17422,N_14985,N_13949);
nor U17423 (N_17423,N_14149,N_12844);
nand U17424 (N_17424,N_14496,N_12695);
nor U17425 (N_17425,N_14415,N_13183);
nor U17426 (N_17426,N_14131,N_13773);
nand U17427 (N_17427,N_12608,N_13314);
nor U17428 (N_17428,N_14591,N_12636);
or U17429 (N_17429,N_13340,N_14554);
or U17430 (N_17430,N_13458,N_14488);
and U17431 (N_17431,N_13634,N_14241);
or U17432 (N_17432,N_14290,N_13193);
and U17433 (N_17433,N_14353,N_14305);
nand U17434 (N_17434,N_14786,N_14468);
nor U17435 (N_17435,N_12771,N_12692);
nor U17436 (N_17436,N_14846,N_13179);
nand U17437 (N_17437,N_13547,N_13946);
and U17438 (N_17438,N_14510,N_13126);
and U17439 (N_17439,N_12934,N_12820);
and U17440 (N_17440,N_13257,N_14776);
and U17441 (N_17441,N_14706,N_14422);
and U17442 (N_17442,N_12554,N_13873);
or U17443 (N_17443,N_14668,N_12820);
or U17444 (N_17444,N_14643,N_13396);
nor U17445 (N_17445,N_12718,N_14781);
nor U17446 (N_17446,N_14034,N_12583);
nor U17447 (N_17447,N_13996,N_14027);
nand U17448 (N_17448,N_13815,N_12729);
nand U17449 (N_17449,N_14928,N_13659);
nand U17450 (N_17450,N_12608,N_14884);
and U17451 (N_17451,N_14208,N_13041);
xor U17452 (N_17452,N_12797,N_12762);
or U17453 (N_17453,N_14136,N_14686);
and U17454 (N_17454,N_13030,N_13225);
nand U17455 (N_17455,N_14743,N_13168);
xor U17456 (N_17456,N_12547,N_14335);
nand U17457 (N_17457,N_14267,N_13281);
and U17458 (N_17458,N_13952,N_14709);
and U17459 (N_17459,N_12952,N_14149);
nand U17460 (N_17460,N_14856,N_12736);
nor U17461 (N_17461,N_12657,N_13349);
nand U17462 (N_17462,N_12658,N_13010);
nor U17463 (N_17463,N_14644,N_14295);
or U17464 (N_17464,N_14961,N_14513);
nand U17465 (N_17465,N_13016,N_13031);
nand U17466 (N_17466,N_12611,N_13809);
or U17467 (N_17467,N_13900,N_14058);
nand U17468 (N_17468,N_14168,N_13582);
nand U17469 (N_17469,N_13902,N_14767);
or U17470 (N_17470,N_13920,N_14319);
nand U17471 (N_17471,N_14058,N_12557);
or U17472 (N_17472,N_12631,N_12773);
and U17473 (N_17473,N_13715,N_13635);
and U17474 (N_17474,N_14995,N_13449);
and U17475 (N_17475,N_13459,N_14938);
or U17476 (N_17476,N_14393,N_13374);
nand U17477 (N_17477,N_14495,N_14009);
nor U17478 (N_17478,N_13170,N_13889);
nor U17479 (N_17479,N_13426,N_14494);
nand U17480 (N_17480,N_13611,N_14415);
and U17481 (N_17481,N_13019,N_12844);
nand U17482 (N_17482,N_13315,N_13748);
nand U17483 (N_17483,N_12900,N_14135);
or U17484 (N_17484,N_12613,N_14464);
nor U17485 (N_17485,N_12649,N_12674);
and U17486 (N_17486,N_13487,N_14700);
or U17487 (N_17487,N_13777,N_14646);
or U17488 (N_17488,N_14201,N_12642);
nor U17489 (N_17489,N_12913,N_13686);
or U17490 (N_17490,N_14200,N_14391);
nand U17491 (N_17491,N_14243,N_14316);
nand U17492 (N_17492,N_13659,N_14589);
nor U17493 (N_17493,N_13256,N_13440);
nor U17494 (N_17494,N_13067,N_13852);
nor U17495 (N_17495,N_14198,N_13340);
nor U17496 (N_17496,N_14213,N_13345);
and U17497 (N_17497,N_14309,N_14625);
and U17498 (N_17498,N_13750,N_13277);
nand U17499 (N_17499,N_12727,N_12743);
nand U17500 (N_17500,N_16842,N_16623);
nand U17501 (N_17501,N_17304,N_16424);
and U17502 (N_17502,N_17382,N_17457);
and U17503 (N_17503,N_16044,N_16238);
nor U17504 (N_17504,N_15376,N_16193);
nand U17505 (N_17505,N_15882,N_15552);
nor U17506 (N_17506,N_15934,N_15128);
or U17507 (N_17507,N_16157,N_16363);
nand U17508 (N_17508,N_16107,N_17464);
nand U17509 (N_17509,N_15687,N_15024);
nor U17510 (N_17510,N_16932,N_15461);
or U17511 (N_17511,N_17431,N_16043);
nor U17512 (N_17512,N_17094,N_16805);
nand U17513 (N_17513,N_17143,N_16445);
nand U17514 (N_17514,N_17479,N_15937);
nor U17515 (N_17515,N_16941,N_17091);
or U17516 (N_17516,N_15519,N_17386);
and U17517 (N_17517,N_16979,N_17490);
nor U17518 (N_17518,N_15413,N_17090);
nand U17519 (N_17519,N_15885,N_15133);
and U17520 (N_17520,N_15849,N_15699);
nor U17521 (N_17521,N_15135,N_15073);
nand U17522 (N_17522,N_15695,N_15455);
or U17523 (N_17523,N_16297,N_15223);
nand U17524 (N_17524,N_16456,N_16715);
nor U17525 (N_17525,N_16006,N_15613);
and U17526 (N_17526,N_15478,N_15603);
nor U17527 (N_17527,N_16147,N_17009);
and U17528 (N_17528,N_16796,N_15174);
nor U17529 (N_17529,N_16637,N_16959);
or U17530 (N_17530,N_17021,N_15653);
nor U17531 (N_17531,N_16684,N_17338);
or U17532 (N_17532,N_17290,N_15783);
nor U17533 (N_17533,N_16722,N_17132);
nor U17534 (N_17534,N_17354,N_15311);
and U17535 (N_17535,N_16426,N_15053);
xor U17536 (N_17536,N_15348,N_16574);
or U17537 (N_17537,N_15308,N_15343);
nand U17538 (N_17538,N_17327,N_16412);
or U17539 (N_17539,N_15522,N_16446);
nor U17540 (N_17540,N_15957,N_15987);
nand U17541 (N_17541,N_15458,N_15365);
nor U17542 (N_17542,N_16054,N_16306);
or U17543 (N_17543,N_16653,N_15044);
nand U17544 (N_17544,N_15755,N_15278);
and U17545 (N_17545,N_15319,N_16775);
nor U17546 (N_17546,N_16906,N_16443);
nand U17547 (N_17547,N_17230,N_17366);
or U17548 (N_17548,N_15147,N_16065);
and U17549 (N_17549,N_16196,N_15930);
or U17550 (N_17550,N_17289,N_15070);
or U17551 (N_17551,N_16388,N_16933);
and U17552 (N_17552,N_15842,N_15822);
nand U17553 (N_17553,N_16129,N_15642);
nand U17554 (N_17554,N_15107,N_16525);
nand U17555 (N_17555,N_15356,N_15960);
nor U17556 (N_17556,N_16516,N_17356);
nor U17557 (N_17557,N_15351,N_15471);
nor U17558 (N_17558,N_17022,N_17039);
nor U17559 (N_17559,N_15046,N_15355);
nand U17560 (N_17560,N_17153,N_17081);
and U17561 (N_17561,N_15159,N_16301);
and U17562 (N_17562,N_15679,N_16831);
or U17563 (N_17563,N_16307,N_16211);
and U17564 (N_17564,N_15340,N_16897);
nand U17565 (N_17565,N_15577,N_17387);
or U17566 (N_17566,N_15899,N_17195);
nand U17567 (N_17567,N_15948,N_15124);
or U17568 (N_17568,N_16045,N_16096);
nor U17569 (N_17569,N_17206,N_17053);
nand U17570 (N_17570,N_16850,N_16635);
nor U17571 (N_17571,N_16570,N_16340);
or U17572 (N_17572,N_17474,N_15908);
and U17573 (N_17573,N_16697,N_16540);
or U17574 (N_17574,N_15647,N_15417);
or U17575 (N_17575,N_16326,N_15239);
nand U17576 (N_17576,N_17309,N_16993);
and U17577 (N_17577,N_15267,N_17026);
or U17578 (N_17578,N_17446,N_16749);
or U17579 (N_17579,N_16234,N_16759);
nor U17580 (N_17580,N_15708,N_15538);
nor U17581 (N_17581,N_15148,N_15315);
nand U17582 (N_17582,N_15169,N_16122);
and U17583 (N_17583,N_17460,N_15126);
nand U17584 (N_17584,N_15359,N_17317);
and U17585 (N_17585,N_16547,N_15336);
or U17586 (N_17586,N_15254,N_16723);
and U17587 (N_17587,N_17003,N_16551);
or U17588 (N_17588,N_16575,N_16103);
or U17589 (N_17589,N_15399,N_15121);
xor U17590 (N_17590,N_15521,N_15415);
and U17591 (N_17591,N_15694,N_15122);
nor U17592 (N_17592,N_16506,N_17211);
and U17593 (N_17593,N_16144,N_16853);
or U17594 (N_17594,N_16510,N_17359);
and U17595 (N_17595,N_16199,N_15588);
nor U17596 (N_17596,N_15326,N_15219);
nand U17597 (N_17597,N_15207,N_16934);
or U17598 (N_17598,N_15890,N_16962);
nor U17599 (N_17599,N_16645,N_16581);
and U17600 (N_17600,N_16729,N_16800);
and U17601 (N_17601,N_15054,N_17286);
nor U17602 (N_17602,N_17133,N_15933);
nor U17603 (N_17603,N_15076,N_16185);
and U17604 (N_17604,N_16752,N_17448);
nand U17605 (N_17605,N_17277,N_15322);
nand U17606 (N_17606,N_16086,N_16782);
nand U17607 (N_17607,N_15697,N_16886);
and U17608 (N_17608,N_15596,N_15607);
or U17609 (N_17609,N_17067,N_15556);
and U17610 (N_17610,N_17451,N_16721);
nor U17611 (N_17611,N_16423,N_16849);
nand U17612 (N_17612,N_16847,N_17057);
or U17613 (N_17613,N_15196,N_15913);
and U17614 (N_17614,N_15422,N_15646);
or U17615 (N_17615,N_15508,N_15144);
nand U17616 (N_17616,N_15535,N_15759);
xnor U17617 (N_17617,N_15985,N_16779);
or U17618 (N_17618,N_17390,N_15280);
nand U17619 (N_17619,N_16611,N_15592);
nor U17620 (N_17620,N_15562,N_15495);
or U17621 (N_17621,N_15001,N_16826);
and U17622 (N_17622,N_15366,N_15705);
nor U17623 (N_17623,N_16056,N_16400);
and U17624 (N_17624,N_17353,N_15247);
nand U17625 (N_17625,N_15447,N_15850);
nand U17626 (N_17626,N_16174,N_17035);
nand U17627 (N_17627,N_16878,N_17433);
and U17628 (N_17628,N_16638,N_17496);
or U17629 (N_17629,N_15981,N_15450);
or U17630 (N_17630,N_16453,N_15777);
and U17631 (N_17631,N_15745,N_15578);
nand U17632 (N_17632,N_15680,N_15132);
or U17633 (N_17633,N_16596,N_15211);
or U17634 (N_17634,N_16376,N_17380);
or U17635 (N_17635,N_15035,N_16728);
nor U17636 (N_17636,N_17238,N_16736);
or U17637 (N_17637,N_16055,N_15640);
and U17638 (N_17638,N_15332,N_16434);
nand U17639 (N_17639,N_15905,N_17325);
nand U17640 (N_17640,N_15180,N_16594);
or U17641 (N_17641,N_17453,N_17241);
or U17642 (N_17642,N_16953,N_16682);
or U17643 (N_17643,N_16300,N_16288);
nand U17644 (N_17644,N_16040,N_16997);
and U17645 (N_17645,N_15955,N_16937);
and U17646 (N_17646,N_17258,N_16405);
or U17647 (N_17647,N_15733,N_17328);
or U17648 (N_17648,N_16656,N_16232);
and U17649 (N_17649,N_16472,N_15880);
and U17650 (N_17650,N_17093,N_16918);
nand U17651 (N_17651,N_16958,N_16244);
nor U17652 (N_17652,N_16414,N_15031);
nand U17653 (N_17653,N_17498,N_15995);
or U17654 (N_17654,N_15674,N_15164);
and U17655 (N_17655,N_15956,N_16140);
and U17656 (N_17656,N_16825,N_17414);
nor U17657 (N_17657,N_16974,N_15528);
and U17658 (N_17658,N_15958,N_17367);
and U17659 (N_17659,N_15190,N_15372);
nor U17660 (N_17660,N_15000,N_15090);
nand U17661 (N_17661,N_15566,N_17429);
nand U17662 (N_17662,N_16860,N_15406);
or U17663 (N_17663,N_15858,N_16823);
nor U17664 (N_17664,N_16145,N_16643);
or U17665 (N_17665,N_17183,N_17342);
nand U17666 (N_17666,N_15623,N_17476);
and U17667 (N_17667,N_16124,N_15205);
nand U17668 (N_17668,N_16318,N_16471);
or U17669 (N_17669,N_16685,N_15421);
and U17670 (N_17670,N_16245,N_16837);
nor U17671 (N_17671,N_15251,N_15184);
nand U17672 (N_17672,N_17240,N_16753);
and U17673 (N_17673,N_17017,N_16275);
or U17674 (N_17674,N_15630,N_15769);
and U17675 (N_17675,N_15770,N_16485);
and U17676 (N_17676,N_15405,N_17472);
nor U17677 (N_17677,N_17307,N_17377);
nor U17678 (N_17678,N_16907,N_17112);
or U17679 (N_17679,N_16520,N_15568);
nor U17680 (N_17680,N_16839,N_15496);
and U17681 (N_17681,N_16672,N_15860);
nand U17682 (N_17682,N_16406,N_15275);
nor U17683 (N_17683,N_15454,N_15884);
or U17684 (N_17684,N_17179,N_16696);
or U17685 (N_17685,N_16008,N_17182);
nor U17686 (N_17686,N_17301,N_15572);
or U17687 (N_17687,N_16755,N_15218);
or U17688 (N_17688,N_15230,N_17218);
xnor U17689 (N_17689,N_16207,N_15602);
nor U17690 (N_17690,N_16222,N_15906);
and U17691 (N_17691,N_15206,N_17260);
or U17692 (N_17692,N_15464,N_15056);
nand U17693 (N_17693,N_15241,N_15195);
and U17694 (N_17694,N_16130,N_17156);
or U17695 (N_17695,N_15507,N_15095);
or U17696 (N_17696,N_16619,N_17308);
or U17697 (N_17697,N_15651,N_16888);
nor U17698 (N_17698,N_16994,N_16950);
nand U17699 (N_17699,N_16532,N_15862);
and U17700 (N_17700,N_16135,N_15766);
and U17701 (N_17701,N_15537,N_15567);
nor U17702 (N_17702,N_15618,N_17397);
nor U17703 (N_17703,N_15487,N_16925);
nand U17704 (N_17704,N_15711,N_16502);
nand U17705 (N_17705,N_17122,N_15990);
nor U17706 (N_17706,N_16127,N_17121);
or U17707 (N_17707,N_15531,N_15814);
nor U17708 (N_17708,N_16731,N_17306);
nor U17709 (N_17709,N_15067,N_16865);
nand U17710 (N_17710,N_16957,N_16692);
or U17711 (N_17711,N_16660,N_16375);
nand U17712 (N_17712,N_16531,N_16571);
and U17713 (N_17713,N_16707,N_15720);
nor U17714 (N_17714,N_17494,N_17312);
nand U17715 (N_17715,N_17269,N_16902);
and U17716 (N_17716,N_17095,N_16354);
and U17717 (N_17717,N_16605,N_16968);
nor U17718 (N_17718,N_15941,N_17170);
or U17719 (N_17719,N_15010,N_16242);
or U17720 (N_17720,N_15545,N_16074);
and U17721 (N_17721,N_15456,N_15030);
nand U17722 (N_17722,N_15083,N_15624);
or U17723 (N_17723,N_16891,N_17219);
nand U17724 (N_17724,N_15982,N_16025);
or U17725 (N_17725,N_15292,N_17436);
nand U17726 (N_17726,N_15082,N_15220);
or U17727 (N_17727,N_15025,N_16746);
nor U17728 (N_17728,N_16970,N_17492);
nand U17729 (N_17729,N_15883,N_16708);
nor U17730 (N_17730,N_15373,N_15228);
and U17731 (N_17731,N_16789,N_15459);
nand U17732 (N_17732,N_16793,N_16599);
and U17733 (N_17733,N_15313,N_17008);
and U17734 (N_17734,N_17409,N_17172);
or U17735 (N_17735,N_16425,N_17271);
and U17736 (N_17736,N_15709,N_15810);
nand U17737 (N_17737,N_15377,N_15703);
or U17738 (N_17738,N_15418,N_15214);
nor U17739 (N_17739,N_16073,N_17276);
nand U17740 (N_17740,N_17344,N_15068);
or U17741 (N_17741,N_15523,N_16386);
nand U17742 (N_17742,N_15657,N_17295);
and U17743 (N_17743,N_16780,N_17469);
nor U17744 (N_17744,N_15802,N_15724);
nor U17745 (N_17745,N_16007,N_16740);
nor U17746 (N_17746,N_15162,N_17080);
or U17747 (N_17747,N_16119,N_15019);
nand U17748 (N_17748,N_16283,N_17234);
and U17749 (N_17749,N_17202,N_16360);
and U17750 (N_17750,N_16355,N_17049);
nor U17751 (N_17751,N_17161,N_16322);
nor U17752 (N_17752,N_15741,N_15172);
or U17753 (N_17753,N_15993,N_17399);
nor U17754 (N_17754,N_16900,N_15892);
nor U17755 (N_17755,N_17097,N_16109);
nor U17756 (N_17756,N_17044,N_17058);
or U17757 (N_17757,N_17106,N_17488);
nor U17758 (N_17758,N_15752,N_16572);
and U17759 (N_17759,N_16584,N_15084);
or U17760 (N_17760,N_16128,N_15998);
nor U17761 (N_17761,N_16545,N_16335);
nor U17762 (N_17762,N_16420,N_16105);
or U17763 (N_17763,N_16845,N_15361);
or U17764 (N_17764,N_15183,N_17125);
and U17765 (N_17765,N_15142,N_15331);
nor U17766 (N_17766,N_15500,N_15050);
nor U17767 (N_17767,N_15550,N_17071);
nor U17768 (N_17768,N_17020,N_16331);
or U17769 (N_17769,N_16436,N_16662);
nor U17770 (N_17770,N_15307,N_15115);
and U17771 (N_17771,N_15846,N_16015);
xnor U17772 (N_17772,N_15344,N_15660);
or U17773 (N_17773,N_17189,N_16181);
or U17774 (N_17774,N_16343,N_16260);
xnor U17775 (N_17775,N_16948,N_15160);
nor U17776 (N_17776,N_16451,N_16150);
nand U17777 (N_17777,N_15779,N_17096);
or U17778 (N_17778,N_15309,N_16352);
nor U17779 (N_17779,N_17216,N_17191);
nor U17780 (N_17780,N_17423,N_15134);
or U17781 (N_17781,N_15789,N_17173);
nor U17782 (N_17782,N_16734,N_16204);
nor U17783 (N_17783,N_15014,N_16587);
or U17784 (N_17784,N_15298,N_17030);
and U17785 (N_17785,N_15776,N_15499);
nor U17786 (N_17786,N_16665,N_15689);
nand U17787 (N_17787,N_15276,N_15834);
nor U17788 (N_17788,N_17484,N_17468);
and U17789 (N_17789,N_15514,N_16158);
or U17790 (N_17790,N_16912,N_16161);
or U17791 (N_17791,N_17394,N_15798);
or U17792 (N_17792,N_15028,N_16562);
and U17793 (N_17793,N_16390,N_16295);
or U17794 (N_17794,N_15598,N_17027);
or U17795 (N_17795,N_17131,N_16497);
xor U17796 (N_17796,N_15758,N_15645);
or U17797 (N_17797,N_15843,N_15966);
nor U17798 (N_17798,N_15467,N_17201);
and U17799 (N_17799,N_17034,N_16776);
or U17800 (N_17800,N_16050,N_16180);
nor U17801 (N_17801,N_15153,N_15775);
or U17802 (N_17802,N_16262,N_15631);
nor U17803 (N_17803,N_17224,N_16601);
nor U17804 (N_17804,N_16866,N_15612);
or U17805 (N_17805,N_17154,N_17120);
nand U17806 (N_17806,N_16975,N_16395);
and U17807 (N_17807,N_15668,N_17365);
or U17808 (N_17808,N_16982,N_16392);
and U17809 (N_17809,N_15715,N_15796);
nor U17810 (N_17810,N_15685,N_16088);
nand U17811 (N_17811,N_15064,N_16302);
and U17812 (N_17812,N_15018,N_15936);
or U17813 (N_17813,N_15226,N_15790);
or U17814 (N_17814,N_16818,N_15504);
nor U17815 (N_17815,N_15593,N_15087);
and U17816 (N_17816,N_16913,N_15480);
or U17817 (N_17817,N_16688,N_15609);
nor U17818 (N_17818,N_17486,N_17480);
nor U17819 (N_17819,N_15113,N_17198);
nand U17820 (N_17820,N_17016,N_17203);
and U17821 (N_17821,N_15388,N_17487);
and U17822 (N_17822,N_15836,N_15333);
or U17823 (N_17823,N_15327,N_15969);
nand U17824 (N_17824,N_16240,N_16976);
or U17825 (N_17825,N_16706,N_15542);
or U17826 (N_17826,N_17391,N_17054);
nor U17827 (N_17827,N_16654,N_16361);
nand U17828 (N_17828,N_17116,N_17250);
and U17829 (N_17829,N_15633,N_17231);
nand U17830 (N_17830,N_15093,N_16291);
or U17831 (N_17831,N_17171,N_15100);
nor U17832 (N_17832,N_16770,N_17443);
nand U17833 (N_17833,N_16998,N_15272);
and U17834 (N_17834,N_16021,N_15738);
and U17835 (N_17835,N_16589,N_15089);
nor U17836 (N_17836,N_16210,N_15546);
and U17837 (N_17837,N_16636,N_15864);
nor U17838 (N_17838,N_15787,N_16965);
or U17839 (N_17839,N_15563,N_16464);
nor U17840 (N_17840,N_17368,N_16440);
nand U17841 (N_17841,N_17184,N_15605);
nand U17842 (N_17842,N_16026,N_17302);
or U17843 (N_17843,N_15345,N_15608);
or U17844 (N_17844,N_16100,N_16033);
nor U17845 (N_17845,N_17422,N_17401);
nand U17846 (N_17846,N_15178,N_15739);
nor U17847 (N_17847,N_16000,N_15003);
nand U17848 (N_17848,N_15060,N_16926);
and U17849 (N_17849,N_15585,N_16338);
and U17850 (N_17850,N_17437,N_17149);
or U17851 (N_17851,N_17175,N_15510);
nor U17852 (N_17852,N_15101,N_15664);
nand U17853 (N_17853,N_17194,N_17174);
and U17854 (N_17854,N_15094,N_17188);
nand U17855 (N_17855,N_15774,N_15390);
nor U17856 (N_17856,N_15484,N_15938);
nor U17857 (N_17857,N_15501,N_15684);
and U17858 (N_17858,N_15785,N_16677);
and U17859 (N_17859,N_15973,N_16265);
nor U17860 (N_17860,N_15179,N_17018);
nor U17861 (N_17861,N_17385,N_15051);
nor U17862 (N_17862,N_17275,N_15554);
and U17863 (N_17863,N_16514,N_16252);
nor U17864 (N_17864,N_15648,N_16840);
nor U17865 (N_17865,N_16649,N_15394);
and U17866 (N_17866,N_15678,N_17345);
and U17867 (N_17867,N_15118,N_15509);
or U17868 (N_17868,N_15290,N_15482);
and U17869 (N_17869,N_16856,N_15518);
and U17870 (N_17870,N_15270,N_16059);
and U17871 (N_17871,N_15075,N_15740);
and U17872 (N_17872,N_17190,N_17374);
nor U17873 (N_17873,N_15665,N_16243);
and U17874 (N_17874,N_15271,N_15844);
nand U17875 (N_17875,N_16342,N_16841);
nand U17876 (N_17876,N_16387,N_16120);
or U17877 (N_17877,N_16590,N_16679);
nand U17878 (N_17878,N_16013,N_16577);
or U17879 (N_17879,N_15264,N_15114);
or U17880 (N_17880,N_15189,N_16330);
and U17881 (N_17881,N_15961,N_16247);
or U17882 (N_17882,N_16765,N_15475);
and U17883 (N_17883,N_16239,N_16750);
nor U17884 (N_17884,N_15666,N_15123);
nor U17885 (N_17885,N_16396,N_16737);
nor U17886 (N_17886,N_15731,N_15579);
nand U17887 (N_17887,N_16117,N_15116);
nor U17888 (N_17888,N_17483,N_15707);
or U17889 (N_17889,N_17226,N_16980);
nand U17890 (N_17890,N_16566,N_16334);
or U17891 (N_17891,N_15571,N_16168);
nand U17892 (N_17892,N_15236,N_16341);
nand U17893 (N_17893,N_16614,N_15168);
nand U17894 (N_17894,N_16220,N_15301);
nor U17895 (N_17895,N_15986,N_17105);
and U17896 (N_17896,N_16366,N_15152);
or U17897 (N_17897,N_16175,N_16588);
or U17898 (N_17898,N_17163,N_16089);
and U17899 (N_17899,N_15006,N_15329);
nor U17900 (N_17900,N_15291,N_16744);
nand U17901 (N_17901,N_16367,N_15763);
and U17902 (N_17902,N_15099,N_16552);
nor U17903 (N_17903,N_16690,N_15718);
nand U17904 (N_17904,N_16651,N_16370);
and U17905 (N_17905,N_17145,N_17262);
nand U17906 (N_17906,N_15516,N_16747);
nor U17907 (N_17907,N_16398,N_15419);
or U17908 (N_17908,N_15334,N_16910);
or U17909 (N_17909,N_16383,N_16814);
nor U17910 (N_17910,N_16467,N_15871);
or U17911 (N_17911,N_15526,N_16791);
or U17912 (N_17912,N_17418,N_16717);
nand U17913 (N_17913,N_17305,N_16009);
and U17914 (N_17914,N_17372,N_15176);
nand U17915 (N_17915,N_17334,N_15294);
nor U17916 (N_17916,N_15932,N_17235);
nand U17917 (N_17917,N_16591,N_16030);
nor U17918 (N_17918,N_16674,N_17413);
and U17919 (N_17919,N_15208,N_15661);
and U17920 (N_17920,N_15801,N_16364);
and U17921 (N_17921,N_16613,N_16309);
nor U17922 (N_17922,N_15245,N_16633);
nor U17923 (N_17923,N_16819,N_17274);
nor U17924 (N_17924,N_17192,N_15616);
xor U17925 (N_17925,N_15944,N_15873);
xor U17926 (N_17926,N_17257,N_15293);
nor U17927 (N_17927,N_15636,N_16689);
nor U17928 (N_17928,N_15644,N_17347);
nand U17929 (N_17929,N_15063,N_15202);
or U17930 (N_17930,N_15221,N_15716);
nor U17931 (N_17931,N_16267,N_16149);
and U17932 (N_17932,N_15852,N_15943);
and U17933 (N_17933,N_17396,N_17032);
nor U17934 (N_17934,N_17069,N_16176);
nor U17935 (N_17935,N_15491,N_16903);
or U17936 (N_17936,N_15011,N_15912);
nand U17937 (N_17937,N_15129,N_17352);
and U17938 (N_17938,N_16217,N_17270);
nor U17939 (N_17939,N_17314,N_15170);
nand U17940 (N_17940,N_17322,N_16031);
or U17941 (N_17941,N_15448,N_15547);
nor U17942 (N_17942,N_15358,N_15463);
nor U17943 (N_17943,N_15146,N_17421);
or U17944 (N_17944,N_17279,N_15881);
nand U17945 (N_17945,N_15753,N_16305);
nand U17946 (N_17946,N_15954,N_16246);
nor U17947 (N_17947,N_16087,N_15105);
xor U17948 (N_17948,N_15536,N_16431);
nor U17949 (N_17949,N_15988,N_16683);
or U17950 (N_17950,N_16554,N_15234);
and U17951 (N_17951,N_17313,N_16716);
nor U17952 (N_17952,N_15284,N_15061);
or U17953 (N_17953,N_16495,N_15493);
nand U17954 (N_17954,N_15553,N_16742);
or U17955 (N_17955,N_16099,N_17025);
and U17956 (N_17956,N_16905,N_17147);
nand U17957 (N_17957,N_17378,N_16206);
nand U17958 (N_17958,N_16983,N_17461);
nand U17959 (N_17959,N_15866,N_17348);
or U17960 (N_17960,N_15364,N_16678);
nand U17961 (N_17961,N_17495,N_16652);
nor U17962 (N_17962,N_15193,N_15041);
nor U17963 (N_17963,N_16470,N_16848);
and U17964 (N_17964,N_16359,N_15012);
nand U17965 (N_17965,N_16714,N_15112);
nand U17966 (N_17966,N_15444,N_16536);
and U17967 (N_17967,N_15964,N_16517);
nand U17968 (N_17968,N_16018,N_16137);
nor U17969 (N_17969,N_17477,N_17169);
nand U17970 (N_17970,N_16209,N_15201);
and U17971 (N_17971,N_15362,N_15224);
or U17972 (N_17972,N_17463,N_16593);
and U17973 (N_17973,N_15983,N_16719);
or U17974 (N_17974,N_16820,N_15439);
nor U17975 (N_17975,N_15681,N_17404);
or U17976 (N_17976,N_16754,N_17491);
nor U17977 (N_17977,N_16017,N_16304);
nor U17978 (N_17978,N_17259,N_16225);
nand U17979 (N_17979,N_17167,N_16313);
and U17980 (N_17980,N_17330,N_16650);
and U17981 (N_17981,N_16964,N_16922);
and U17982 (N_17982,N_16811,N_17245);
and U17983 (N_17983,N_15795,N_15723);
or U17984 (N_17984,N_15404,N_16557);
or U17985 (N_17985,N_15979,N_16830);
nand U17986 (N_17986,N_16930,N_16868);
or U17987 (N_17987,N_16067,N_15977);
and U17988 (N_17988,N_15791,N_17410);
and U17989 (N_17989,N_16399,N_15235);
or U17990 (N_17990,N_15274,N_16155);
nand U17991 (N_17991,N_15229,N_15649);
nor U17992 (N_17992,N_16720,N_16644);
nand U17993 (N_17993,N_15346,N_15296);
or U17994 (N_17994,N_16081,N_16080);
nor U17995 (N_17995,N_15347,N_16138);
or U17996 (N_17996,N_16756,N_15140);
and U17997 (N_17997,N_15845,N_15825);
or U17998 (N_17998,N_16430,N_16996);
nand U17999 (N_17999,N_17015,N_16563);
and U18000 (N_18000,N_15036,N_16567);
or U18001 (N_18001,N_17158,N_16310);
nand U18002 (N_18002,N_15071,N_15204);
and U18003 (N_18003,N_15859,N_15497);
nor U18004 (N_18004,N_16256,N_15768);
and U18005 (N_18005,N_16476,N_16862);
nor U18006 (N_18006,N_17362,N_16403);
nand U18007 (N_18007,N_17239,N_15869);
or U18008 (N_18008,N_15091,N_16439);
nor U18009 (N_18009,N_16325,N_15706);
or U18010 (N_18010,N_15772,N_15416);
or U18011 (N_18011,N_15942,N_15217);
or U18012 (N_18012,N_16846,N_17110);
nand U18013 (N_18013,N_15033,N_16854);
and U18014 (N_18014,N_16528,N_15260);
nand U18015 (N_18015,N_17331,N_15503);
nand U18016 (N_18016,N_17303,N_16876);
nand U18017 (N_18017,N_15200,N_15910);
nand U18018 (N_18018,N_17236,N_16833);
nor U18019 (N_18019,N_15506,N_16491);
nor U18020 (N_18020,N_16810,N_16870);
and U18021 (N_18021,N_15939,N_16486);
nand U18022 (N_18022,N_17168,N_16901);
nand U18023 (N_18023,N_15244,N_15318);
or U18024 (N_18024,N_17319,N_17134);
and U18025 (N_18025,N_16822,N_15805);
or U18026 (N_18026,N_17337,N_15137);
nand U18027 (N_18027,N_15875,N_15433);
and U18028 (N_18028,N_15688,N_15520);
or U18029 (N_18029,N_15565,N_16947);
nor U18030 (N_18030,N_15252,N_16449);
or U18031 (N_18031,N_16493,N_16328);
nor U18032 (N_18032,N_17292,N_16014);
and U18033 (N_18033,N_17459,N_15149);
and U18034 (N_18034,N_17223,N_16909);
or U18035 (N_18035,N_16938,N_15804);
and U18036 (N_18036,N_16208,N_15671);
nand U18037 (N_18037,N_16943,N_17400);
or U18038 (N_18038,N_15717,N_15306);
or U18039 (N_18039,N_16573,N_16187);
xnor U18040 (N_18040,N_15383,N_15305);
nor U18041 (N_18041,N_16991,N_16098);
nor U18042 (N_18042,N_15736,N_16835);
nor U18043 (N_18043,N_15161,N_16869);
or U18044 (N_18044,N_15898,N_15632);
or U18045 (N_18045,N_15992,N_16797);
or U18046 (N_18046,N_15316,N_17265);
nand U18047 (N_18047,N_16458,N_15436);
nand U18048 (N_18048,N_16829,N_16097);
or U18049 (N_18049,N_16249,N_16861);
nor U18050 (N_18050,N_16002,N_15916);
and U18051 (N_18051,N_16164,N_16289);
and U18052 (N_18052,N_16695,N_16290);
or U18053 (N_18053,N_16713,N_15601);
nand U18054 (N_18054,N_17229,N_17291);
nand U18055 (N_18055,N_17281,N_15074);
or U18056 (N_18056,N_15713,N_16492);
or U18057 (N_18057,N_16442,N_16299);
and U18058 (N_18058,N_17108,N_17146);
nor U18059 (N_18059,N_16494,N_15677);
and U18060 (N_18060,N_17389,N_15625);
and U18061 (N_18061,N_17082,N_15812);
nand U18062 (N_18062,N_15156,N_15452);
nand U18063 (N_18063,N_16374,N_16046);
nand U18064 (N_18064,N_15492,N_16751);
and U18065 (N_18065,N_16076,N_16203);
nand U18066 (N_18066,N_17298,N_15742);
and U18067 (N_18067,N_15569,N_15886);
nand U18068 (N_18068,N_15185,N_16710);
and U18069 (N_18069,N_16987,N_17037);
or U18070 (N_18070,N_16774,N_15265);
nor U18071 (N_18071,N_17031,N_16156);
nor U18072 (N_18072,N_17076,N_16264);
or U18073 (N_18073,N_15548,N_15861);
or U18074 (N_18074,N_17011,N_16999);
nor U18075 (N_18075,N_17242,N_16786);
nand U18076 (N_18076,N_15048,N_16788);
and U18077 (N_18077,N_16466,N_16227);
nor U18078 (N_18078,N_16487,N_15911);
nor U18079 (N_18079,N_16954,N_17176);
nor U18080 (N_18080,N_17023,N_16034);
and U18081 (N_18081,N_15971,N_16807);
nor U18082 (N_18082,N_17092,N_15412);
and U18083 (N_18083,N_16618,N_16610);
nor U18084 (N_18084,N_15473,N_15323);
nand U18085 (N_18085,N_17285,N_15980);
nor U18086 (N_18086,N_17126,N_16915);
nor U18087 (N_18087,N_16763,N_17014);
or U18088 (N_18088,N_15749,N_16268);
and U18089 (N_18089,N_16160,N_16236);
and U18090 (N_18090,N_17129,N_15026);
or U18091 (N_18091,N_16681,N_15266);
and U18092 (N_18092,N_16942,N_15434);
nand U18093 (N_18093,N_15778,N_16544);
nand U18094 (N_18094,N_17412,N_16693);
nor U18095 (N_18095,N_16864,N_15925);
and U18096 (N_18096,N_16278,N_16027);
nor U18097 (N_18097,N_16447,N_16162);
nor U18098 (N_18098,N_16365,N_15803);
xor U18099 (N_18099,N_16981,N_17228);
nand U18100 (N_18100,N_15029,N_16556);
or U18101 (N_18101,N_15544,N_17178);
or U18102 (N_18102,N_16687,N_17107);
and U18103 (N_18103,N_17072,N_16069);
nor U18104 (N_18104,N_17329,N_17357);
or U18105 (N_18105,N_15839,N_15079);
nor U18106 (N_18106,N_16042,N_16413);
or U18107 (N_18107,N_16172,N_16371);
or U18108 (N_18108,N_15693,N_16480);
nor U18109 (N_18109,N_15233,N_16029);
nand U18110 (N_18110,N_15767,N_15472);
and U18111 (N_18111,N_17458,N_15370);
and U18112 (N_18112,N_16308,N_16523);
and U18113 (N_18113,N_15575,N_17462);
or U18114 (N_18114,N_16131,N_15652);
or U18115 (N_18115,N_16255,N_16529);
or U18116 (N_18116,N_17253,N_17221);
or U18117 (N_18117,N_15287,N_17185);
nor U18118 (N_18118,N_15387,N_15922);
or U18119 (N_18119,N_17089,N_15215);
nand U18120 (N_18120,N_15756,N_15670);
or U18121 (N_18121,N_17045,N_15654);
nor U18122 (N_18122,N_15950,N_16657);
nand U18123 (N_18123,N_16576,N_16205);
or U18124 (N_18124,N_17209,N_16382);
and U18125 (N_18125,N_15854,N_17002);
nor U18126 (N_18126,N_15438,N_15761);
or U18127 (N_18127,N_15381,N_15069);
or U18128 (N_18128,N_16995,N_16726);
nand U18129 (N_18129,N_17056,N_17136);
nor U18130 (N_18130,N_17038,N_16141);
or U18131 (N_18131,N_15261,N_16024);
and U18132 (N_18132,N_16631,N_15401);
and U18133 (N_18133,N_17041,N_17442);
or U18134 (N_18134,N_16956,N_16767);
nor U18135 (N_18135,N_15232,N_15532);
nor U18136 (N_18136,N_16539,N_17197);
nor U18137 (N_18137,N_16004,N_15445);
or U18138 (N_18138,N_15295,N_16213);
nor U18139 (N_18139,N_15328,N_16266);
or U18140 (N_18140,N_16020,N_15258);
or U18141 (N_18141,N_16292,N_15929);
nor U18142 (N_18142,N_15828,N_15962);
or U18143 (N_18143,N_16022,N_16419);
and U18144 (N_18144,N_15641,N_15963);
nand U18145 (N_18145,N_15897,N_16923);
or U18146 (N_18146,N_16459,N_16852);
nand U18147 (N_18147,N_16808,N_17428);
nor U18148 (N_18148,N_17243,N_15324);
or U18149 (N_18149,N_15901,N_16385);
nand U18150 (N_18150,N_17225,N_16874);
nand U18151 (N_18151,N_15062,N_15700);
and U18152 (N_18152,N_16990,N_15835);
or U18153 (N_18153,N_17077,N_16011);
or U18154 (N_18154,N_15104,N_17475);
nand U18155 (N_18155,N_16163,N_15907);
and U18156 (N_18156,N_16189,N_16658);
nor U18157 (N_18157,N_15469,N_16879);
nor U18158 (N_18158,N_17293,N_16151);
and U18159 (N_18159,N_15800,N_15619);
nor U18160 (N_18160,N_15302,N_15020);
and U18161 (N_18161,N_17335,N_15468);
and U18162 (N_18162,N_15430,N_16667);
nand U18163 (N_18163,N_15728,N_15557);
nand U18164 (N_18164,N_16285,N_16899);
nor U18165 (N_18165,N_17111,N_15395);
nor U18166 (N_18166,N_16049,N_16603);
and U18167 (N_18167,N_15034,N_17333);
and U18168 (N_18168,N_16123,N_15304);
or U18169 (N_18169,N_17296,N_16315);
nor U18170 (N_18170,N_15017,N_17193);
or U18171 (N_18171,N_15177,N_16748);
and U18172 (N_18172,N_15638,N_16104);
and U18173 (N_18173,N_15167,N_15692);
or U18174 (N_18174,N_17162,N_16960);
and U18175 (N_18175,N_15494,N_16542);
or U18176 (N_18176,N_15746,N_16634);
or U18177 (N_18177,N_15868,N_16787);
and U18178 (N_18178,N_15829,N_15096);
or U18179 (N_18179,N_15999,N_15407);
nor U18180 (N_18180,N_17127,N_15154);
nand U18181 (N_18181,N_15673,N_16475);
nor U18182 (N_18182,N_15837,N_16524);
or U18183 (N_18183,N_16216,N_16978);
or U18184 (N_18184,N_16263,N_17232);
nor U18185 (N_18185,N_16478,N_16973);
nor U18186 (N_18186,N_16329,N_16051);
nor U18187 (N_18187,N_15946,N_15889);
or U18188 (N_18188,N_16802,N_16815);
or U18189 (N_18189,N_17249,N_16384);
nand U18190 (N_18190,N_16795,N_17024);
nor U18191 (N_18191,N_16812,N_16550);
nor U18192 (N_18192,N_15582,N_17441);
nand U18193 (N_18193,N_15512,N_17100);
nand U18194 (N_18194,N_15411,N_16877);
nor U18195 (N_18195,N_16287,N_16102);
nand U18196 (N_18196,N_15610,N_17434);
nand U18197 (N_18197,N_15838,N_16377);
or U18198 (N_18198,N_15476,N_16621);
or U18199 (N_18199,N_17248,N_15511);
and U18200 (N_18200,N_15502,N_16988);
or U18201 (N_18201,N_17444,N_16134);
nand U18202 (N_18202,N_16858,N_16518);
or U18203 (N_18203,N_15021,N_15683);
nand U18204 (N_18204,N_16257,N_16411);
nand U18205 (N_18205,N_16333,N_15710);
and U18206 (N_18206,N_17326,N_15970);
nand U18207 (N_18207,N_17361,N_15479);
and U18208 (N_18208,N_15634,N_16416);
and U18209 (N_18209,N_15909,N_16666);
nand U18210 (N_18210,N_17118,N_17310);
and U18211 (N_18211,N_17315,N_17419);
nor U18212 (N_18212,N_15924,N_16356);
and U18213 (N_18213,N_16178,N_16703);
nor U18214 (N_18214,N_16704,N_15682);
and U18215 (N_18215,N_15066,N_17376);
or U18216 (N_18216,N_15077,N_15996);
or U18217 (N_18217,N_15369,N_16896);
nand U18218 (N_18218,N_17255,N_15876);
nand U18219 (N_18219,N_16963,N_16409);
nor U18220 (N_18220,N_17164,N_15400);
and U18221 (N_18221,N_15606,N_16664);
nand U18222 (N_18222,N_17181,N_16700);
nand U18223 (N_18223,N_16694,N_15968);
nor U18224 (N_18224,N_15055,N_17237);
and U18225 (N_18225,N_15446,N_15363);
or U18226 (N_18226,N_17426,N_17355);
and U18227 (N_18227,N_15449,N_15915);
nor U18228 (N_18228,N_17300,N_16277);
nor U18229 (N_18229,N_16125,N_16012);
nand U18230 (N_18230,N_15517,N_17392);
nand U18231 (N_18231,N_16512,N_15097);
nand U18232 (N_18232,N_17316,N_15227);
nand U18233 (N_18233,N_17200,N_16111);
nor U18234 (N_18234,N_17166,N_17152);
or U18235 (N_18235,N_16270,N_15940);
or U18236 (N_18236,N_15902,N_16461);
or U18237 (N_18237,N_15675,N_17233);
or U18238 (N_18238,N_16345,N_17294);
and U18239 (N_18239,N_15032,N_15893);
or U18240 (N_18240,N_15959,N_15923);
nor U18241 (N_18241,N_16455,N_15549);
nand U18242 (N_18242,N_17288,N_15253);
and U18243 (N_18243,N_16961,N_16920);
nand U18244 (N_18244,N_17088,N_16939);
or U18245 (N_18245,N_16640,N_15457);
or U18246 (N_18246,N_16101,N_15597);
and U18247 (N_18247,N_16799,N_16437);
and U18248 (N_18248,N_17078,N_15587);
nor U18249 (N_18249,N_16781,N_15342);
nor U18250 (N_18250,N_16188,N_16062);
or U18251 (N_18251,N_17151,N_15863);
and U18252 (N_18252,N_16339,N_15188);
nand U18253 (N_18253,N_16857,N_17320);
nor U18254 (N_18254,N_17000,N_17222);
nand U18255 (N_18255,N_15927,N_15481);
nand U18256 (N_18256,N_17123,N_16380);
and U18257 (N_18257,N_15397,N_17036);
nand U18258 (N_18258,N_17052,N_17407);
nor U18259 (N_18259,N_16757,N_15145);
nor U18260 (N_18260,N_16202,N_16488);
and U18261 (N_18261,N_16661,N_16010);
or U18262 (N_18262,N_17402,N_16762);
and U18263 (N_18263,N_16739,N_17485);
nand U18264 (N_18264,N_15181,N_17101);
nand U18265 (N_18265,N_16883,N_16070);
nand U18266 (N_18266,N_15110,N_16259);
xnor U18267 (N_18267,N_15559,N_15285);
or U18268 (N_18268,N_15428,N_15255);
nor U18269 (N_18269,N_15794,N_16121);
nor U18270 (N_18270,N_17363,N_17138);
nand U18271 (N_18271,N_15663,N_16183);
or U18272 (N_18272,N_16481,N_16945);
and U18273 (N_18273,N_16058,N_15426);
nor U18274 (N_18274,N_15555,N_15040);
and U18275 (N_18275,N_15187,N_15820);
nand U18276 (N_18276,N_16609,N_16454);
and U18277 (N_18277,N_16035,N_16873);
and U18278 (N_18278,N_16499,N_15690);
or U18279 (N_18279,N_15994,N_16816);
or U18280 (N_18280,N_16118,N_16967);
or U18281 (N_18281,N_16404,N_17416);
nand U18282 (N_18282,N_15106,N_16916);
xnor U18283 (N_18283,N_16659,N_16642);
nand U18284 (N_18284,N_17098,N_16555);
or U18285 (N_18285,N_16221,N_15008);
and U18286 (N_18286,N_16955,N_16732);
and U18287 (N_18287,N_17099,N_16324);
or U18288 (N_18288,N_16989,N_16323);
nand U18289 (N_18289,N_16813,N_15833);
and U18290 (N_18290,N_16632,N_15719);
or U18291 (N_18291,N_16827,N_16462);
nor U18292 (N_18292,N_17139,N_15525);
and U18293 (N_18293,N_16804,N_15175);
nand U18294 (N_18294,N_15007,N_17332);
or U18295 (N_18295,N_16711,N_15246);
or U18296 (N_18296,N_17213,N_15534);
and U18297 (N_18297,N_16773,N_15442);
nand U18298 (N_18298,N_17471,N_17177);
nor U18299 (N_18299,N_15622,N_16625);
nand U18300 (N_18300,N_16935,N_15762);
and U18301 (N_18301,N_15141,N_16273);
and U18302 (N_18302,N_16337,N_16389);
and U18303 (N_18303,N_16686,N_15815);
or U18304 (N_18304,N_16503,N_15453);
nand U18305 (N_18305,N_16269,N_15248);
nand U18306 (N_18306,N_16761,N_17051);
nand U18307 (N_18307,N_15393,N_16250);
or U18308 (N_18308,N_17349,N_16490);
and U18309 (N_18309,N_17408,N_17010);
nor U18310 (N_18310,N_15629,N_16919);
nor U18311 (N_18311,N_16349,N_15757);
or U18312 (N_18312,N_16559,N_15978);
xnor U18313 (N_18313,N_15824,N_15976);
or U18314 (N_18314,N_16401,N_16867);
nand U18315 (N_18315,N_16228,N_16535);
or U18316 (N_18316,N_16586,N_15409);
nor U18317 (N_18317,N_17432,N_16887);
and U18318 (N_18318,N_17215,N_15599);
nor U18319 (N_18319,N_16612,N_16075);
and U18320 (N_18320,N_15367,N_15658);
and U18321 (N_18321,N_15595,N_16639);
and U18322 (N_18322,N_15714,N_17466);
or U18323 (N_18323,N_17117,N_16053);
nor U18324 (N_18324,N_15460,N_16641);
and U18325 (N_18325,N_15991,N_16484);
or U18326 (N_18326,N_15806,N_16855);
or U18327 (N_18327,N_16241,N_17499);
and U18328 (N_18328,N_15250,N_15297);
nand U18329 (N_18329,N_17266,N_15935);
nand U18330 (N_18330,N_15764,N_15917);
nand U18331 (N_18331,N_15627,N_16253);
and U18332 (N_18332,N_16393,N_17046);
nand U18333 (N_18333,N_16068,N_16169);
and U18334 (N_18334,N_17244,N_16078);
nand U18335 (N_18335,N_15303,N_15576);
nor U18336 (N_18336,N_16489,N_17104);
nand U18337 (N_18337,N_16680,N_16357);
nand U18338 (N_18338,N_16548,N_16582);
and U18339 (N_18339,N_15043,N_17141);
nand U18340 (N_18340,N_15614,N_16090);
nor U18341 (N_18341,N_17430,N_16585);
or U18342 (N_18342,N_15799,N_15997);
nor U18343 (N_18343,N_15879,N_16602);
and U18344 (N_18344,N_16139,N_17375);
nor U18345 (N_18345,N_15403,N_15424);
nand U18346 (N_18346,N_15158,N_16921);
or U18347 (N_18347,N_17063,N_15088);
and U18348 (N_18348,N_16951,N_16894);
nand U18349 (N_18349,N_17001,N_16235);
and U18350 (N_18350,N_15039,N_15580);
and U18351 (N_18351,N_15797,N_15379);
nor U18352 (N_18352,N_17263,N_15727);
and U18353 (N_18353,N_17299,N_16186);
nor U18354 (N_18354,N_16448,N_17346);
and U18355 (N_18355,N_15268,N_17452);
nor U18356 (N_18356,N_16060,N_17424);
nand U18357 (N_18357,N_17283,N_16143);
and U18358 (N_18358,N_16477,N_15443);
nor U18359 (N_18359,N_15953,N_15330);
and U18360 (N_18360,N_15895,N_15465);
or U18361 (N_18361,N_16949,N_15440);
nor U18362 (N_18362,N_17383,N_17311);
nor U18363 (N_18363,N_15166,N_16092);
nand U18364 (N_18364,N_16875,N_15462);
or U18365 (N_18365,N_16832,N_16082);
nand U18366 (N_18366,N_16085,N_16607);
xnor U18367 (N_18367,N_16606,N_16880);
nand U18368 (N_18368,N_16182,N_17142);
and U18369 (N_18369,N_15437,N_15353);
or U18370 (N_18370,N_16133,N_16838);
or U18371 (N_18371,N_17373,N_16889);
nor U18372 (N_18372,N_15655,N_16223);
nand U18373 (N_18373,N_15378,N_16992);
xnor U18374 (N_18374,N_16108,N_15257);
and U18375 (N_18375,N_15038,N_15972);
nor U18376 (N_18376,N_15281,N_16166);
and U18377 (N_18377,N_15748,N_15808);
nand U18378 (N_18378,N_15754,N_17205);
nor U18379 (N_18379,N_16892,N_16595);
nor U18380 (N_18380,N_16167,N_15249);
nor U18381 (N_18381,N_16258,N_16699);
and U18382 (N_18382,N_15788,N_15865);
nand U18383 (N_18383,N_16444,N_15139);
nor U18384 (N_18384,N_17212,N_16546);
or U18385 (N_18385,N_16673,N_15635);
and U18386 (N_18386,N_15744,N_15841);
nand U18387 (N_18387,N_16792,N_15870);
and U18388 (N_18388,N_16159,N_17278);
or U18389 (N_18389,N_16469,N_15840);
nand U18390 (N_18390,N_16429,N_16197);
nor U18391 (N_18391,N_16373,N_15380);
and U18392 (N_18392,N_15904,N_16911);
and U18393 (N_18393,N_16537,N_17013);
or U18394 (N_18394,N_16298,N_15477);
nor U18395 (N_18395,N_16698,N_15615);
or U18396 (N_18396,N_16415,N_15022);
and U18397 (N_18397,N_17074,N_16583);
or U18398 (N_18398,N_16378,N_15676);
nor U18399 (N_18399,N_16146,N_16093);
nor U18400 (N_18400,N_15847,N_16408);
and U18401 (N_18401,N_17124,N_15721);
and U18402 (N_18402,N_16348,N_15931);
and U18403 (N_18403,N_15967,N_15765);
nand U18404 (N_18404,N_17109,N_17028);
and U18405 (N_18405,N_16741,N_16116);
nor U18406 (N_18406,N_16676,N_16760);
nor U18407 (N_18407,N_15429,N_15015);
nand U18408 (N_18408,N_15650,N_16115);
nor U18409 (N_18409,N_16834,N_16432);
nor U18410 (N_18410,N_15131,N_16091);
or U18411 (N_18411,N_15877,N_15743);
and U18412 (N_18412,N_16615,N_15005);
or U18413 (N_18413,N_15819,N_15891);
nand U18414 (N_18414,N_15354,N_15386);
nor U18415 (N_18415,N_17395,N_17297);
nor U18416 (N_18416,N_16016,N_15286);
or U18417 (N_18417,N_15098,N_16622);
or U18418 (N_18418,N_16312,N_15667);
and U18419 (N_18419,N_16895,N_16179);
or U18420 (N_18420,N_15357,N_15212);
nor U18421 (N_18421,N_17066,N_15466);
and U18422 (N_18422,N_17196,N_16479);
nor U18423 (N_18423,N_15600,N_16177);
and U18424 (N_18424,N_15626,N_17493);
xor U18425 (N_18425,N_16195,N_17159);
nor U18426 (N_18426,N_16280,N_16350);
and U18427 (N_18427,N_15591,N_16533);
and U18428 (N_18428,N_17042,N_15109);
or U18429 (N_18429,N_16561,N_16032);
and U18430 (N_18430,N_16038,N_17360);
nand U18431 (N_18431,N_17059,N_17135);
and U18432 (N_18432,N_17398,N_15527);
nor U18433 (N_18433,N_15384,N_16663);
nand U18434 (N_18434,N_15811,N_15818);
and U18435 (N_18435,N_15529,N_15541);
nor U18436 (N_18436,N_17160,N_16279);
and U18437 (N_18437,N_15659,N_15581);
or U18438 (N_18438,N_15878,N_16801);
and U18439 (N_18439,N_15823,N_17083);
nand U18440 (N_18440,N_15117,N_17454);
and U18441 (N_18441,N_16284,N_15751);
nand U18442 (N_18442,N_16904,N_15349);
and U18443 (N_18443,N_16526,N_17455);
or U18444 (N_18444,N_16039,N_16254);
and U18445 (N_18445,N_17130,N_17450);
or U18446 (N_18446,N_15058,N_17417);
nand U18447 (N_18447,N_15414,N_15887);
nor U18448 (N_18448,N_16597,N_15222);
and U18449 (N_18449,N_16314,N_15059);
nand U18450 (N_18450,N_17340,N_15945);
and U18451 (N_18451,N_17155,N_16417);
or U18452 (N_18452,N_15564,N_17068);
nor U18453 (N_18453,N_16438,N_15947);
and U18454 (N_18454,N_16114,N_17497);
and U18455 (N_18455,N_16712,N_16527);
nand U18456 (N_18456,N_16048,N_15052);
nand U18457 (N_18457,N_17006,N_16794);
or U18458 (N_18458,N_17087,N_15611);
or U18459 (N_18459,N_15150,N_15300);
or U18460 (N_18460,N_15851,N_15045);
nor U18461 (N_18461,N_16190,N_16036);
nor U18462 (N_18462,N_16001,N_16165);
or U18463 (N_18463,N_15283,N_17449);
or U18464 (N_18464,N_17128,N_15590);
nand U18465 (N_18465,N_17427,N_17252);
and U18466 (N_18466,N_16433,N_16332);
nor U18467 (N_18467,N_15560,N_15339);
or U18468 (N_18468,N_15299,N_17012);
nand U18469 (N_18469,N_16543,N_16931);
and U18470 (N_18470,N_15080,N_17482);
or U18471 (N_18471,N_16063,N_16110);
or U18472 (N_18472,N_15078,N_15490);
or U18473 (N_18473,N_15856,N_15583);
or U18474 (N_18474,N_16817,N_16944);
nor U18475 (N_18475,N_16984,N_16407);
nor U18476 (N_18476,N_17208,N_15341);
nand U18477 (N_18477,N_16316,N_16184);
or U18478 (N_18478,N_16061,N_15277);
nand U18479 (N_18479,N_15573,N_15198);
nor U18480 (N_18480,N_16450,N_16702);
or U18481 (N_18481,N_17150,N_16421);
nor U18482 (N_18482,N_16604,N_17318);
or U18483 (N_18483,N_15337,N_16274);
nand U18484 (N_18484,N_15734,N_17381);
nor U18485 (N_18485,N_15621,N_17336);
nand U18486 (N_18486,N_15874,N_16508);
nor U18487 (N_18487,N_15952,N_17439);
or U18488 (N_18488,N_15102,N_17473);
nand U18489 (N_18489,N_16626,N_15857);
or U18490 (N_18490,N_15561,N_15203);
and U18491 (N_18491,N_15240,N_16766);
or U18492 (N_18492,N_15350,N_15813);
nand U18493 (N_18493,N_15423,N_16237);
nor U18494 (N_18494,N_15784,N_15750);
and U18495 (N_18495,N_16072,N_16418);
nand U18496 (N_18496,N_16735,N_15262);
nor U18497 (N_18497,N_17282,N_16251);
and U18498 (N_18498,N_15669,N_17369);
nand U18499 (N_18499,N_17256,N_17435);
nand U18500 (N_18500,N_16885,N_15900);
nand U18501 (N_18501,N_15136,N_16758);
nor U18502 (N_18502,N_16463,N_15786);
and U18503 (N_18503,N_17119,N_15023);
nor U18504 (N_18504,N_15282,N_15974);
nor U18505 (N_18505,N_16917,N_17144);
nor U18506 (N_18506,N_16768,N_15488);
nand U18507 (N_18507,N_17079,N_17210);
nand U18508 (N_18508,N_15586,N_15325);
nand U18509 (N_18509,N_16872,N_17033);
or U18510 (N_18510,N_15210,N_17489);
and U18511 (N_18511,N_15108,N_15530);
nand U18512 (N_18512,N_15213,N_17379);
and U18513 (N_18513,N_16230,N_17114);
nand U18514 (N_18514,N_16113,N_15965);
and U18515 (N_18515,N_16972,N_15817);
or U18516 (N_18516,N_15639,N_15735);
or U18517 (N_18517,N_15543,N_16669);
nand U18518 (N_18518,N_15288,N_15049);
and U18519 (N_18519,N_16224,N_15773);
nand U18520 (N_18520,N_15004,N_16771);
nand U18521 (N_18521,N_16410,N_16569);
nor U18522 (N_18522,N_15451,N_17048);
nor U18523 (N_18523,N_16064,N_16457);
or U18524 (N_18524,N_16136,N_16231);
or U18525 (N_18525,N_16513,N_16041);
nand U18526 (N_18526,N_15013,N_15125);
or U18527 (N_18527,N_15317,N_17060);
nor U18528 (N_18528,N_15729,N_16522);
or U18529 (N_18529,N_15656,N_16986);
nor U18530 (N_18530,N_16005,N_16598);
nand U18531 (N_18531,N_15470,N_17254);
nor U18532 (N_18532,N_17227,N_17005);
and U18533 (N_18533,N_16381,N_15382);
nor U18534 (N_18534,N_15872,N_17478);
or U18535 (N_18535,N_16549,N_16624);
and U18536 (N_18536,N_15826,N_15072);
nand U18537 (N_18537,N_15231,N_17405);
and U18538 (N_18538,N_16047,N_16727);
and U18539 (N_18539,N_15398,N_15951);
and U18540 (N_18540,N_16066,N_16296);
nor U18541 (N_18541,N_15269,N_16003);
or U18542 (N_18542,N_16336,N_17113);
nand U18543 (N_18543,N_15392,N_16271);
nand U18544 (N_18544,N_16372,N_16629);
nor U18545 (N_18545,N_17115,N_17180);
nor U18546 (N_18546,N_16985,N_16670);
and U18547 (N_18547,N_16317,N_16785);
nand U18548 (N_18548,N_16353,N_16509);
nor U18549 (N_18549,N_15238,N_17070);
or U18550 (N_18550,N_16148,N_15360);
or U18551 (N_18551,N_16369,N_16394);
nand U18552 (N_18552,N_16465,N_16630);
or U18553 (N_18553,N_15984,N_16824);
or U18554 (N_18554,N_16028,N_16851);
or U18555 (N_18555,N_15888,N_16803);
or U18556 (N_18556,N_17007,N_16733);
and U18557 (N_18557,N_15165,N_16940);
nor U18558 (N_18558,N_15374,N_15410);
or U18559 (N_18559,N_16778,N_15186);
and U18560 (N_18560,N_15722,N_16908);
or U18561 (N_18561,N_15427,N_15505);
or U18562 (N_18562,N_15216,N_16600);
or U18563 (N_18563,N_17220,N_17370);
nand U18564 (N_18564,N_15780,N_15589);
nand U18565 (N_18565,N_17358,N_16627);
and U18566 (N_18566,N_16152,N_16655);
or U18567 (N_18567,N_17019,N_17350);
or U18568 (N_18568,N_15009,N_15092);
or U18569 (N_18569,N_17364,N_16884);
and U18570 (N_18570,N_15574,N_16294);
and U18571 (N_18571,N_16946,N_15919);
nand U18572 (N_18572,N_15896,N_17251);
or U18573 (N_18573,N_16173,N_15975);
nand U18574 (N_18574,N_17324,N_15686);
and U18575 (N_18575,N_15726,N_15848);
nand U18576 (N_18576,N_16863,N_15338);
and U18577 (N_18577,N_17341,N_17470);
and U18578 (N_18578,N_16379,N_17247);
or U18579 (N_18579,N_17420,N_16777);
and U18580 (N_18580,N_16608,N_16498);
nor U18581 (N_18581,N_17323,N_17199);
and U18582 (N_18582,N_15701,N_15737);
or U18583 (N_18583,N_16725,N_15524);
and U18584 (N_18584,N_16668,N_17343);
nor U18585 (N_18585,N_16519,N_17148);
and U18586 (N_18586,N_15173,N_16214);
or U18587 (N_18587,N_17047,N_15832);
or U18588 (N_18588,N_15119,N_15391);
and U18589 (N_18589,N_15243,N_16971);
and U18590 (N_18590,N_16212,N_16286);
or U18591 (N_18591,N_17102,N_15027);
nand U18592 (N_18592,N_16293,N_15402);
nand U18593 (N_18593,N_16079,N_15111);
nor U18594 (N_18594,N_17186,N_17137);
xor U18595 (N_18595,N_17064,N_17204);
or U18596 (N_18596,N_15263,N_16347);
or U18597 (N_18597,N_16215,N_17055);
nor U18598 (N_18598,N_15485,N_17085);
nand U18599 (N_18599,N_16422,N_17403);
and U18600 (N_18600,N_15730,N_16745);
or U18601 (N_18601,N_15042,N_16474);
or U18602 (N_18602,N_17351,N_17061);
and U18603 (N_18603,N_15127,N_15793);
and U18604 (N_18604,N_15368,N_16037);
and U18605 (N_18605,N_16718,N_15712);
and U18606 (N_18606,N_15065,N_16368);
nand U18607 (N_18607,N_16427,N_15259);
nand U18608 (N_18608,N_16927,N_15130);
or U18609 (N_18609,N_15103,N_15279);
nand U18610 (N_18610,N_16783,N_16358);
nor U18611 (N_18611,N_15435,N_17261);
nand U18612 (N_18612,N_16671,N_16568);
or U18613 (N_18613,N_16738,N_17043);
nand U18614 (N_18614,N_16311,N_15867);
nand U18615 (N_18615,N_16617,N_17445);
nor U18616 (N_18616,N_15335,N_15420);
nand U18617 (N_18617,N_17165,N_15515);
and U18618 (N_18618,N_15558,N_15389);
nand U18619 (N_18619,N_15321,N_16871);
and U18620 (N_18620,N_16928,N_16052);
nor U18621 (N_18621,N_15928,N_15441);
nor U18622 (N_18622,N_15989,N_16530);
nor U18623 (N_18623,N_17217,N_15037);
nor U18624 (N_18624,N_16790,N_16675);
and U18625 (N_18625,N_16460,N_16560);
or U18626 (N_18626,N_15086,N_16936);
and U18627 (N_18627,N_15242,N_17465);
or U18628 (N_18628,N_15620,N_16023);
nand U18629 (N_18629,N_16218,N_16500);
or U18630 (N_18630,N_15352,N_17467);
or U18631 (N_18631,N_16893,N_15894);
nor U18632 (N_18632,N_16809,N_15771);
or U18633 (N_18633,N_16057,N_15151);
xnor U18634 (N_18634,N_15747,N_15120);
xnor U18635 (N_18635,N_15171,N_15584);
or U18636 (N_18636,N_15138,N_15486);
or U18637 (N_18637,N_16435,N_15192);
and U18638 (N_18638,N_16628,N_15691);
nand U18639 (N_18639,N_15314,N_16881);
nand U18640 (N_18640,N_17440,N_15237);
and U18641 (N_18641,N_15732,N_15551);
nand U18642 (N_18642,N_16844,N_16402);
nand U18643 (N_18643,N_15081,N_16171);
or U18644 (N_18644,N_15760,N_17075);
and U18645 (N_18645,N_16142,N_15256);
nor U18646 (N_18646,N_16391,N_16320);
nand U18647 (N_18647,N_16616,N_16579);
nor U18648 (N_18648,N_15533,N_15672);
and U18649 (N_18649,N_16772,N_17411);
or U18650 (N_18650,N_16647,N_16898);
and U18651 (N_18651,N_17264,N_16724);
nor U18652 (N_18652,N_17207,N_16346);
and U18653 (N_18653,N_16798,N_15489);
and U18654 (N_18654,N_15057,N_16452);
nand U18655 (N_18655,N_16836,N_16321);
nor U18656 (N_18656,N_17280,N_16441);
nand U18657 (N_18657,N_16821,N_17103);
nand U18658 (N_18658,N_16153,N_15725);
and U18659 (N_18659,N_16969,N_15827);
nor U18660 (N_18660,N_15821,N_17157);
and U18661 (N_18661,N_17062,N_15809);
or U18662 (N_18662,N_16538,N_17273);
or U18663 (N_18663,N_16094,N_15782);
and U18664 (N_18664,N_16106,N_15816);
and U18665 (N_18665,N_15781,N_16929);
nor U18666 (N_18666,N_16282,N_15914);
or U18667 (N_18667,N_17086,N_16468);
nand U18668 (N_18668,N_16592,N_15163);
nor U18669 (N_18669,N_15016,N_15197);
nand U18670 (N_18670,N_15853,N_15498);
and U18671 (N_18671,N_16843,N_16504);
and U18672 (N_18672,N_15807,N_15604);
nand U18673 (N_18673,N_15949,N_15273);
and U18674 (N_18674,N_15831,N_15320);
nand U18675 (N_18675,N_16705,N_16558);
or U18676 (N_18676,N_15698,N_16397);
nor U18677 (N_18677,N_16730,N_16966);
nand U18678 (N_18678,N_17393,N_16154);
and U18679 (N_18679,N_16276,N_15182);
or U18680 (N_18680,N_16303,N_15483);
nor U18681 (N_18681,N_17456,N_15431);
nor U18682 (N_18682,N_15085,N_15225);
nand U18683 (N_18683,N_15594,N_17050);
and U18684 (N_18684,N_16701,N_16496);
nor U18685 (N_18685,N_16084,N_15312);
nor U18686 (N_18686,N_16882,N_16473);
and U18687 (N_18687,N_16483,N_16077);
or U18688 (N_18688,N_16192,N_16233);
or U18689 (N_18689,N_15855,N_16482);
and U18690 (N_18690,N_16272,N_16743);
nor U18691 (N_18691,N_16764,N_16515);
and U18692 (N_18692,N_16507,N_16691);
or U18693 (N_18693,N_15289,N_15540);
nor U18694 (N_18694,N_16112,N_16924);
nand U18695 (N_18695,N_16194,N_15474);
and U18696 (N_18696,N_15918,N_17073);
nor U18697 (N_18697,N_16784,N_17438);
nor U18698 (N_18698,N_16198,N_17272);
or U18699 (N_18699,N_17040,N_17214);
nor U18700 (N_18700,N_15662,N_15570);
or U18701 (N_18701,N_17321,N_15926);
nor U18702 (N_18702,N_17339,N_17384);
or U18703 (N_18703,N_17246,N_15513);
nor U18704 (N_18704,N_15375,N_17267);
nor U18705 (N_18705,N_16281,N_16327);
nand U18706 (N_18706,N_16521,N_16553);
or U18707 (N_18707,N_16019,N_17425);
nand U18708 (N_18708,N_16261,N_17084);
or U18709 (N_18709,N_16126,N_16580);
nor U18710 (N_18710,N_17406,N_17140);
nor U18711 (N_18711,N_17481,N_16191);
and U18712 (N_18712,N_15408,N_16620);
and U18713 (N_18713,N_16071,N_15157);
and U18714 (N_18714,N_16219,N_16351);
or U18715 (N_18715,N_17187,N_15143);
or U18716 (N_18716,N_15432,N_15702);
and U18717 (N_18717,N_17065,N_16344);
nand U18718 (N_18718,N_15155,N_15539);
nand U18719 (N_18719,N_16578,N_15371);
and U18720 (N_18720,N_15792,N_15903);
or U18721 (N_18721,N_15199,N_16511);
nand U18722 (N_18722,N_15002,N_15643);
or U18723 (N_18723,N_16769,N_17371);
nand U18724 (N_18724,N_17029,N_15696);
or U18725 (N_18725,N_16200,N_17388);
or U18726 (N_18726,N_16083,N_16132);
nor U18727 (N_18727,N_17268,N_16709);
or U18728 (N_18728,N_17415,N_16501);
and U18729 (N_18729,N_15425,N_15830);
or U18730 (N_18730,N_16229,N_16828);
nand U18731 (N_18731,N_16914,N_16362);
nor U18732 (N_18732,N_15921,N_15310);
and U18733 (N_18733,N_15704,N_15628);
or U18734 (N_18734,N_16095,N_16170);
xnor U18735 (N_18735,N_16646,N_16952);
or U18736 (N_18736,N_16648,N_16977);
or U18737 (N_18737,N_15637,N_17447);
nand U18738 (N_18738,N_15191,N_15920);
xnor U18739 (N_18739,N_17287,N_16564);
or U18740 (N_18740,N_16428,N_15385);
or U18741 (N_18741,N_15396,N_16226);
nor U18742 (N_18742,N_16890,N_16565);
or U18743 (N_18743,N_16534,N_16505);
and U18744 (N_18744,N_16248,N_16319);
and U18745 (N_18745,N_15617,N_17284);
nand U18746 (N_18746,N_15194,N_15209);
nor U18747 (N_18747,N_16859,N_16541);
nand U18748 (N_18748,N_16201,N_16806);
or U18749 (N_18749,N_17004,N_15047);
nor U18750 (N_18750,N_15570,N_16727);
nand U18751 (N_18751,N_17248,N_15620);
nor U18752 (N_18752,N_15763,N_16877);
nor U18753 (N_18753,N_16868,N_16286);
nand U18754 (N_18754,N_15368,N_16605);
xnor U18755 (N_18755,N_16177,N_16803);
and U18756 (N_18756,N_16054,N_16252);
xor U18757 (N_18757,N_17094,N_16664);
nor U18758 (N_18758,N_17482,N_15056);
nor U18759 (N_18759,N_16112,N_16947);
and U18760 (N_18760,N_16451,N_16233);
nor U18761 (N_18761,N_16354,N_16492);
nor U18762 (N_18762,N_17186,N_16773);
or U18763 (N_18763,N_17399,N_15591);
nand U18764 (N_18764,N_16886,N_17145);
nor U18765 (N_18765,N_15612,N_15322);
and U18766 (N_18766,N_16659,N_16807);
and U18767 (N_18767,N_16864,N_17316);
nor U18768 (N_18768,N_15946,N_15494);
and U18769 (N_18769,N_15733,N_15797);
nor U18770 (N_18770,N_15657,N_15209);
and U18771 (N_18771,N_16425,N_15845);
nor U18772 (N_18772,N_17202,N_16244);
nand U18773 (N_18773,N_16978,N_17205);
or U18774 (N_18774,N_16964,N_17102);
nand U18775 (N_18775,N_16552,N_15216);
nand U18776 (N_18776,N_16831,N_17209);
and U18777 (N_18777,N_17138,N_16300);
nor U18778 (N_18778,N_15178,N_16645);
and U18779 (N_18779,N_15217,N_15737);
nand U18780 (N_18780,N_15985,N_15781);
xor U18781 (N_18781,N_15229,N_17146);
and U18782 (N_18782,N_15114,N_15928);
or U18783 (N_18783,N_17193,N_16584);
or U18784 (N_18784,N_17204,N_15795);
and U18785 (N_18785,N_15062,N_16635);
or U18786 (N_18786,N_17233,N_16956);
nand U18787 (N_18787,N_15847,N_15707);
or U18788 (N_18788,N_17469,N_15633);
and U18789 (N_18789,N_17424,N_15845);
or U18790 (N_18790,N_15912,N_16331);
and U18791 (N_18791,N_17085,N_16828);
nor U18792 (N_18792,N_15067,N_16588);
or U18793 (N_18793,N_15644,N_15360);
nand U18794 (N_18794,N_16447,N_15535);
nand U18795 (N_18795,N_16404,N_15372);
or U18796 (N_18796,N_16082,N_16414);
nor U18797 (N_18797,N_17378,N_16882);
nor U18798 (N_18798,N_15474,N_17005);
nand U18799 (N_18799,N_15868,N_15049);
or U18800 (N_18800,N_16512,N_16858);
or U18801 (N_18801,N_17208,N_16833);
nand U18802 (N_18802,N_16159,N_16037);
and U18803 (N_18803,N_15683,N_15817);
nand U18804 (N_18804,N_15715,N_16674);
or U18805 (N_18805,N_17137,N_15150);
nor U18806 (N_18806,N_16873,N_15971);
nor U18807 (N_18807,N_15986,N_15012);
and U18808 (N_18808,N_15795,N_15083);
and U18809 (N_18809,N_17209,N_16705);
and U18810 (N_18810,N_17340,N_17013);
nand U18811 (N_18811,N_16357,N_16747);
or U18812 (N_18812,N_17258,N_17261);
nand U18813 (N_18813,N_17172,N_16165);
nand U18814 (N_18814,N_16631,N_17060);
nor U18815 (N_18815,N_16874,N_15124);
nand U18816 (N_18816,N_17250,N_17376);
and U18817 (N_18817,N_16885,N_16806);
or U18818 (N_18818,N_17141,N_16913);
xor U18819 (N_18819,N_16525,N_16490);
and U18820 (N_18820,N_16840,N_16559);
nand U18821 (N_18821,N_15855,N_15204);
or U18822 (N_18822,N_17189,N_15327);
xor U18823 (N_18823,N_16912,N_15297);
nand U18824 (N_18824,N_16743,N_15991);
nand U18825 (N_18825,N_15984,N_17383);
nor U18826 (N_18826,N_15903,N_15680);
nor U18827 (N_18827,N_16934,N_16679);
and U18828 (N_18828,N_17349,N_15624);
nand U18829 (N_18829,N_15828,N_15953);
and U18830 (N_18830,N_17095,N_17062);
nor U18831 (N_18831,N_17468,N_16430);
or U18832 (N_18832,N_17321,N_17265);
or U18833 (N_18833,N_16300,N_15188);
or U18834 (N_18834,N_17274,N_16528);
nor U18835 (N_18835,N_17086,N_16935);
nor U18836 (N_18836,N_15284,N_16849);
nand U18837 (N_18837,N_15013,N_17310);
or U18838 (N_18838,N_16245,N_16212);
nor U18839 (N_18839,N_17297,N_17221);
nand U18840 (N_18840,N_16142,N_17341);
nand U18841 (N_18841,N_17403,N_15148);
nand U18842 (N_18842,N_17119,N_15848);
nor U18843 (N_18843,N_15981,N_15162);
nand U18844 (N_18844,N_16160,N_17342);
nand U18845 (N_18845,N_15140,N_16638);
nand U18846 (N_18846,N_15134,N_15712);
nor U18847 (N_18847,N_16275,N_16140);
or U18848 (N_18848,N_15335,N_15318);
nand U18849 (N_18849,N_15948,N_17016);
nand U18850 (N_18850,N_15129,N_17061);
or U18851 (N_18851,N_17306,N_16405);
xnor U18852 (N_18852,N_15228,N_16456);
and U18853 (N_18853,N_15575,N_15872);
or U18854 (N_18854,N_16663,N_15988);
nor U18855 (N_18855,N_15728,N_16483);
nand U18856 (N_18856,N_16302,N_17485);
or U18857 (N_18857,N_16194,N_15107);
or U18858 (N_18858,N_17047,N_15091);
nor U18859 (N_18859,N_16066,N_15015);
nor U18860 (N_18860,N_15005,N_16385);
xor U18861 (N_18861,N_16253,N_16918);
or U18862 (N_18862,N_15617,N_15152);
and U18863 (N_18863,N_15654,N_17263);
nand U18864 (N_18864,N_16910,N_15317);
nand U18865 (N_18865,N_16173,N_17183);
nor U18866 (N_18866,N_16546,N_15233);
and U18867 (N_18867,N_16954,N_16977);
and U18868 (N_18868,N_17385,N_15811);
and U18869 (N_18869,N_16068,N_17014);
nor U18870 (N_18870,N_16731,N_16835);
or U18871 (N_18871,N_15616,N_17476);
nor U18872 (N_18872,N_15275,N_16886);
nand U18873 (N_18873,N_16421,N_16473);
or U18874 (N_18874,N_16270,N_15053);
nor U18875 (N_18875,N_16878,N_15686);
nor U18876 (N_18876,N_15836,N_16546);
nor U18877 (N_18877,N_15200,N_16668);
and U18878 (N_18878,N_15585,N_17145);
and U18879 (N_18879,N_17079,N_17161);
nand U18880 (N_18880,N_16761,N_15117);
nor U18881 (N_18881,N_16274,N_15160);
or U18882 (N_18882,N_15827,N_16293);
or U18883 (N_18883,N_16704,N_15821);
and U18884 (N_18884,N_16302,N_15701);
nand U18885 (N_18885,N_16916,N_16174);
or U18886 (N_18886,N_16349,N_15393);
or U18887 (N_18887,N_17037,N_17100);
or U18888 (N_18888,N_16726,N_17140);
or U18889 (N_18889,N_16293,N_16524);
nand U18890 (N_18890,N_15416,N_16828);
and U18891 (N_18891,N_16876,N_16727);
nand U18892 (N_18892,N_16048,N_15556);
nor U18893 (N_18893,N_16493,N_16095);
and U18894 (N_18894,N_16714,N_16098);
or U18895 (N_18895,N_15467,N_15762);
nand U18896 (N_18896,N_16015,N_15993);
nand U18897 (N_18897,N_16274,N_16051);
or U18898 (N_18898,N_16703,N_16240);
and U18899 (N_18899,N_17229,N_16152);
nand U18900 (N_18900,N_16667,N_15262);
and U18901 (N_18901,N_17248,N_15238);
nand U18902 (N_18902,N_16109,N_15363);
nand U18903 (N_18903,N_15059,N_15799);
or U18904 (N_18904,N_17342,N_15437);
nor U18905 (N_18905,N_17428,N_15370);
or U18906 (N_18906,N_17284,N_16197);
and U18907 (N_18907,N_16736,N_15023);
nor U18908 (N_18908,N_16647,N_16150);
or U18909 (N_18909,N_15399,N_17451);
and U18910 (N_18910,N_15695,N_16687);
nand U18911 (N_18911,N_17047,N_17090);
or U18912 (N_18912,N_16615,N_15446);
nand U18913 (N_18913,N_15793,N_16651);
or U18914 (N_18914,N_16477,N_16068);
and U18915 (N_18915,N_16658,N_16297);
or U18916 (N_18916,N_15130,N_17244);
and U18917 (N_18917,N_16055,N_15234);
and U18918 (N_18918,N_16364,N_16843);
and U18919 (N_18919,N_17392,N_17426);
and U18920 (N_18920,N_16581,N_17268);
or U18921 (N_18921,N_16570,N_15134);
nand U18922 (N_18922,N_15874,N_16144);
nor U18923 (N_18923,N_16454,N_15979);
or U18924 (N_18924,N_16445,N_16628);
nor U18925 (N_18925,N_16893,N_17272);
and U18926 (N_18926,N_15114,N_16582);
and U18927 (N_18927,N_15313,N_15378);
nand U18928 (N_18928,N_16344,N_17164);
and U18929 (N_18929,N_17038,N_16668);
and U18930 (N_18930,N_15395,N_16423);
nor U18931 (N_18931,N_15331,N_17178);
or U18932 (N_18932,N_17455,N_16576);
and U18933 (N_18933,N_15998,N_16853);
and U18934 (N_18934,N_15883,N_15723);
and U18935 (N_18935,N_15593,N_15686);
nand U18936 (N_18936,N_15876,N_16992);
nand U18937 (N_18937,N_16905,N_16318);
and U18938 (N_18938,N_17177,N_16844);
nand U18939 (N_18939,N_17141,N_17093);
nor U18940 (N_18940,N_17417,N_16696);
and U18941 (N_18941,N_15757,N_15277);
nand U18942 (N_18942,N_16806,N_17226);
or U18943 (N_18943,N_17307,N_15378);
nor U18944 (N_18944,N_15357,N_15966);
xor U18945 (N_18945,N_15197,N_15155);
nor U18946 (N_18946,N_16092,N_15005);
nor U18947 (N_18947,N_17012,N_15228);
xor U18948 (N_18948,N_16680,N_16142);
nand U18949 (N_18949,N_15819,N_15762);
and U18950 (N_18950,N_15014,N_15284);
nor U18951 (N_18951,N_16404,N_16247);
and U18952 (N_18952,N_16943,N_17357);
and U18953 (N_18953,N_16321,N_17101);
and U18954 (N_18954,N_17457,N_15637);
or U18955 (N_18955,N_15827,N_15269);
and U18956 (N_18956,N_15421,N_15549);
nand U18957 (N_18957,N_15522,N_16381);
nor U18958 (N_18958,N_16017,N_16803);
nand U18959 (N_18959,N_15368,N_17307);
and U18960 (N_18960,N_17304,N_15987);
nand U18961 (N_18961,N_16174,N_15148);
or U18962 (N_18962,N_16922,N_17235);
or U18963 (N_18963,N_16495,N_15095);
or U18964 (N_18964,N_16256,N_15928);
and U18965 (N_18965,N_16519,N_15598);
and U18966 (N_18966,N_16478,N_15973);
nor U18967 (N_18967,N_16530,N_16770);
and U18968 (N_18968,N_17303,N_15871);
nand U18969 (N_18969,N_15980,N_16013);
or U18970 (N_18970,N_17469,N_17228);
nor U18971 (N_18971,N_15405,N_15411);
and U18972 (N_18972,N_15960,N_16973);
nor U18973 (N_18973,N_16815,N_17339);
nand U18974 (N_18974,N_15291,N_16225);
or U18975 (N_18975,N_15011,N_15316);
or U18976 (N_18976,N_15984,N_15508);
and U18977 (N_18977,N_15716,N_17158);
or U18978 (N_18978,N_16656,N_15539);
nand U18979 (N_18979,N_17407,N_15508);
and U18980 (N_18980,N_16737,N_17376);
and U18981 (N_18981,N_15938,N_16507);
nand U18982 (N_18982,N_16754,N_15072);
or U18983 (N_18983,N_16699,N_15067);
and U18984 (N_18984,N_16722,N_15467);
nand U18985 (N_18985,N_16550,N_15144);
nand U18986 (N_18986,N_16847,N_15518);
nor U18987 (N_18987,N_16210,N_15138);
nand U18988 (N_18988,N_15313,N_15090);
and U18989 (N_18989,N_16214,N_16527);
nand U18990 (N_18990,N_17203,N_16698);
nor U18991 (N_18991,N_16302,N_15630);
nor U18992 (N_18992,N_16874,N_15021);
or U18993 (N_18993,N_15302,N_15282);
nor U18994 (N_18994,N_16126,N_15603);
nor U18995 (N_18995,N_15211,N_17327);
and U18996 (N_18996,N_15318,N_16846);
nor U18997 (N_18997,N_15322,N_16644);
and U18998 (N_18998,N_16809,N_16138);
and U18999 (N_18999,N_16300,N_16291);
and U19000 (N_19000,N_15851,N_17206);
nor U19001 (N_19001,N_16224,N_16703);
or U19002 (N_19002,N_16923,N_15433);
and U19003 (N_19003,N_16351,N_15410);
or U19004 (N_19004,N_15219,N_15173);
nor U19005 (N_19005,N_15546,N_15855);
or U19006 (N_19006,N_15195,N_17390);
nand U19007 (N_19007,N_17202,N_16319);
or U19008 (N_19008,N_16119,N_17321);
nand U19009 (N_19009,N_15169,N_16744);
and U19010 (N_19010,N_16899,N_16394);
nor U19011 (N_19011,N_16558,N_15708);
nand U19012 (N_19012,N_15976,N_16593);
or U19013 (N_19013,N_16391,N_15090);
nor U19014 (N_19014,N_16300,N_15588);
and U19015 (N_19015,N_17080,N_15423);
or U19016 (N_19016,N_17127,N_15131);
and U19017 (N_19017,N_17107,N_16868);
and U19018 (N_19018,N_16121,N_17244);
and U19019 (N_19019,N_17041,N_16352);
and U19020 (N_19020,N_16126,N_15752);
nand U19021 (N_19021,N_17353,N_16314);
nand U19022 (N_19022,N_16879,N_15293);
or U19023 (N_19023,N_16838,N_15307);
and U19024 (N_19024,N_16765,N_15479);
nand U19025 (N_19025,N_15185,N_15498);
or U19026 (N_19026,N_15457,N_17022);
nand U19027 (N_19027,N_17019,N_16700);
nand U19028 (N_19028,N_15728,N_16977);
or U19029 (N_19029,N_17454,N_17424);
nand U19030 (N_19030,N_15079,N_15742);
or U19031 (N_19031,N_16082,N_15756);
nor U19032 (N_19032,N_16845,N_15996);
nand U19033 (N_19033,N_16872,N_16508);
and U19034 (N_19034,N_16152,N_16681);
or U19035 (N_19035,N_16426,N_16840);
and U19036 (N_19036,N_17421,N_15364);
nor U19037 (N_19037,N_15427,N_15547);
nand U19038 (N_19038,N_16530,N_16759);
nor U19039 (N_19039,N_15734,N_16825);
nor U19040 (N_19040,N_16792,N_15157);
nand U19041 (N_19041,N_15084,N_16389);
nor U19042 (N_19042,N_16147,N_15469);
nand U19043 (N_19043,N_15817,N_15024);
nor U19044 (N_19044,N_16631,N_15700);
nor U19045 (N_19045,N_15375,N_16359);
or U19046 (N_19046,N_15290,N_16026);
nand U19047 (N_19047,N_16515,N_16370);
nand U19048 (N_19048,N_15763,N_16030);
nor U19049 (N_19049,N_17109,N_17372);
nand U19050 (N_19050,N_16103,N_15506);
nand U19051 (N_19051,N_16248,N_15780);
nand U19052 (N_19052,N_16405,N_17343);
nor U19053 (N_19053,N_16255,N_17076);
and U19054 (N_19054,N_15789,N_15840);
or U19055 (N_19055,N_15192,N_16284);
and U19056 (N_19056,N_15132,N_16034);
nand U19057 (N_19057,N_15283,N_15478);
xnor U19058 (N_19058,N_16944,N_16375);
nand U19059 (N_19059,N_17472,N_15797);
or U19060 (N_19060,N_16248,N_16102);
or U19061 (N_19061,N_17233,N_15348);
nand U19062 (N_19062,N_17164,N_17401);
nor U19063 (N_19063,N_15067,N_15870);
nor U19064 (N_19064,N_15792,N_15853);
nand U19065 (N_19065,N_17288,N_16864);
nand U19066 (N_19066,N_16474,N_16611);
nand U19067 (N_19067,N_16225,N_17305);
nor U19068 (N_19068,N_15115,N_15306);
nand U19069 (N_19069,N_17010,N_17481);
or U19070 (N_19070,N_16909,N_15725);
or U19071 (N_19071,N_16437,N_17306);
nor U19072 (N_19072,N_15784,N_16130);
and U19073 (N_19073,N_17063,N_15489);
and U19074 (N_19074,N_16664,N_16548);
nand U19075 (N_19075,N_15965,N_17154);
or U19076 (N_19076,N_17148,N_16627);
or U19077 (N_19077,N_16274,N_16625);
nand U19078 (N_19078,N_15234,N_15572);
nor U19079 (N_19079,N_15692,N_16390);
nand U19080 (N_19080,N_16534,N_16676);
or U19081 (N_19081,N_17204,N_17233);
nor U19082 (N_19082,N_15219,N_16123);
and U19083 (N_19083,N_15104,N_15912);
or U19084 (N_19084,N_17066,N_15041);
and U19085 (N_19085,N_16364,N_16098);
nor U19086 (N_19086,N_15285,N_16825);
or U19087 (N_19087,N_16449,N_15357);
or U19088 (N_19088,N_15310,N_16123);
nand U19089 (N_19089,N_16866,N_16783);
or U19090 (N_19090,N_15422,N_15713);
and U19091 (N_19091,N_17318,N_15705);
or U19092 (N_19092,N_15229,N_15755);
or U19093 (N_19093,N_17453,N_15560);
and U19094 (N_19094,N_16587,N_16867);
nand U19095 (N_19095,N_17029,N_15935);
or U19096 (N_19096,N_15137,N_17357);
nor U19097 (N_19097,N_17195,N_15556);
or U19098 (N_19098,N_16456,N_15981);
and U19099 (N_19099,N_17242,N_15628);
and U19100 (N_19100,N_17071,N_16301);
or U19101 (N_19101,N_15996,N_15035);
nand U19102 (N_19102,N_16767,N_16283);
or U19103 (N_19103,N_15818,N_16784);
nor U19104 (N_19104,N_16409,N_17415);
or U19105 (N_19105,N_15314,N_17092);
or U19106 (N_19106,N_15904,N_16927);
or U19107 (N_19107,N_16623,N_16807);
nand U19108 (N_19108,N_15047,N_16608);
and U19109 (N_19109,N_16536,N_15249);
nand U19110 (N_19110,N_15206,N_15690);
nand U19111 (N_19111,N_15472,N_16338);
nor U19112 (N_19112,N_16232,N_15733);
nand U19113 (N_19113,N_16854,N_17168);
or U19114 (N_19114,N_15733,N_16626);
and U19115 (N_19115,N_16004,N_16162);
nand U19116 (N_19116,N_16870,N_16149);
nand U19117 (N_19117,N_15458,N_16919);
and U19118 (N_19118,N_15327,N_16999);
nand U19119 (N_19119,N_16251,N_15604);
and U19120 (N_19120,N_16481,N_15360);
and U19121 (N_19121,N_16959,N_16739);
nor U19122 (N_19122,N_15723,N_15061);
and U19123 (N_19123,N_15816,N_16557);
and U19124 (N_19124,N_16119,N_16654);
nor U19125 (N_19125,N_17220,N_16681);
nand U19126 (N_19126,N_16674,N_15211);
and U19127 (N_19127,N_15396,N_16592);
and U19128 (N_19128,N_17100,N_15300);
or U19129 (N_19129,N_15506,N_15560);
nor U19130 (N_19130,N_15188,N_15184);
xnor U19131 (N_19131,N_16083,N_15701);
nand U19132 (N_19132,N_16225,N_16635);
nand U19133 (N_19133,N_15838,N_17280);
or U19134 (N_19134,N_16021,N_16813);
and U19135 (N_19135,N_17159,N_15501);
nand U19136 (N_19136,N_15058,N_15980);
nand U19137 (N_19137,N_17405,N_17129);
nand U19138 (N_19138,N_17488,N_17164);
nand U19139 (N_19139,N_17021,N_15169);
or U19140 (N_19140,N_16945,N_15849);
nand U19141 (N_19141,N_15890,N_16260);
and U19142 (N_19142,N_16890,N_15459);
and U19143 (N_19143,N_16318,N_15765);
or U19144 (N_19144,N_17199,N_16021);
nand U19145 (N_19145,N_17087,N_17125);
or U19146 (N_19146,N_16148,N_15737);
and U19147 (N_19147,N_16116,N_16164);
and U19148 (N_19148,N_17045,N_15896);
or U19149 (N_19149,N_17382,N_15483);
and U19150 (N_19150,N_16888,N_15639);
and U19151 (N_19151,N_16834,N_15763);
nor U19152 (N_19152,N_17188,N_17009);
nand U19153 (N_19153,N_17350,N_15529);
or U19154 (N_19154,N_16569,N_17141);
or U19155 (N_19155,N_16146,N_16130);
nor U19156 (N_19156,N_15498,N_17289);
nor U19157 (N_19157,N_15334,N_16515);
and U19158 (N_19158,N_17138,N_17331);
or U19159 (N_19159,N_16621,N_15143);
and U19160 (N_19160,N_16492,N_17125);
nand U19161 (N_19161,N_15019,N_17188);
nor U19162 (N_19162,N_15274,N_16097);
or U19163 (N_19163,N_16840,N_17020);
nor U19164 (N_19164,N_17387,N_15744);
or U19165 (N_19165,N_15537,N_16902);
and U19166 (N_19166,N_17003,N_16142);
nor U19167 (N_19167,N_15236,N_15021);
or U19168 (N_19168,N_15839,N_15461);
nand U19169 (N_19169,N_15618,N_16531);
and U19170 (N_19170,N_17071,N_15747);
or U19171 (N_19171,N_16257,N_17472);
nor U19172 (N_19172,N_17499,N_17299);
or U19173 (N_19173,N_15999,N_15602);
nor U19174 (N_19174,N_16363,N_16343);
nand U19175 (N_19175,N_17442,N_16104);
nor U19176 (N_19176,N_15790,N_17235);
or U19177 (N_19177,N_16737,N_17002);
nand U19178 (N_19178,N_17449,N_15111);
or U19179 (N_19179,N_15344,N_15026);
nor U19180 (N_19180,N_16819,N_16948);
or U19181 (N_19181,N_15259,N_15783);
and U19182 (N_19182,N_16591,N_16692);
nand U19183 (N_19183,N_16893,N_16217);
or U19184 (N_19184,N_17424,N_16432);
or U19185 (N_19185,N_15238,N_17324);
and U19186 (N_19186,N_16896,N_16200);
or U19187 (N_19187,N_15863,N_15294);
nand U19188 (N_19188,N_17439,N_15605);
nor U19189 (N_19189,N_15942,N_15537);
nand U19190 (N_19190,N_16239,N_16722);
nand U19191 (N_19191,N_15245,N_16812);
or U19192 (N_19192,N_15007,N_16124);
or U19193 (N_19193,N_15789,N_16613);
nor U19194 (N_19194,N_15232,N_15520);
xor U19195 (N_19195,N_17119,N_15315);
nand U19196 (N_19196,N_15625,N_16928);
nor U19197 (N_19197,N_15410,N_16311);
nor U19198 (N_19198,N_17092,N_16496);
and U19199 (N_19199,N_17016,N_15586);
and U19200 (N_19200,N_17302,N_17054);
nor U19201 (N_19201,N_17034,N_15379);
and U19202 (N_19202,N_17363,N_17244);
nand U19203 (N_19203,N_15498,N_16533);
nor U19204 (N_19204,N_15904,N_15048);
and U19205 (N_19205,N_16223,N_16001);
and U19206 (N_19206,N_15942,N_16053);
and U19207 (N_19207,N_17053,N_17215);
or U19208 (N_19208,N_16198,N_15134);
nor U19209 (N_19209,N_17138,N_15442);
and U19210 (N_19210,N_15129,N_15198);
or U19211 (N_19211,N_15160,N_16109);
and U19212 (N_19212,N_15581,N_17063);
nand U19213 (N_19213,N_17461,N_16603);
nor U19214 (N_19214,N_15422,N_15825);
nor U19215 (N_19215,N_16978,N_15506);
nor U19216 (N_19216,N_16385,N_17146);
nor U19217 (N_19217,N_16858,N_17082);
nor U19218 (N_19218,N_15026,N_16975);
or U19219 (N_19219,N_17383,N_15288);
and U19220 (N_19220,N_16851,N_16946);
or U19221 (N_19221,N_16274,N_16642);
nand U19222 (N_19222,N_17158,N_16624);
or U19223 (N_19223,N_16096,N_17212);
nand U19224 (N_19224,N_17145,N_16155);
or U19225 (N_19225,N_16218,N_17042);
and U19226 (N_19226,N_15600,N_17470);
nand U19227 (N_19227,N_17483,N_16000);
nor U19228 (N_19228,N_16142,N_16996);
or U19229 (N_19229,N_15402,N_16596);
nor U19230 (N_19230,N_15225,N_15724);
xor U19231 (N_19231,N_16726,N_15223);
nor U19232 (N_19232,N_16105,N_17007);
nand U19233 (N_19233,N_15520,N_17071);
nor U19234 (N_19234,N_16817,N_17379);
nand U19235 (N_19235,N_16865,N_15504);
nand U19236 (N_19236,N_17427,N_16149);
nor U19237 (N_19237,N_15179,N_15944);
or U19238 (N_19238,N_15434,N_15974);
and U19239 (N_19239,N_16400,N_15977);
or U19240 (N_19240,N_17038,N_16387);
and U19241 (N_19241,N_17007,N_15631);
nand U19242 (N_19242,N_15581,N_16380);
and U19243 (N_19243,N_16728,N_15116);
nand U19244 (N_19244,N_17039,N_17084);
nor U19245 (N_19245,N_15434,N_15061);
and U19246 (N_19246,N_16360,N_16473);
or U19247 (N_19247,N_16157,N_16294);
or U19248 (N_19248,N_15629,N_16648);
or U19249 (N_19249,N_15036,N_17093);
nor U19250 (N_19250,N_15330,N_16612);
nor U19251 (N_19251,N_17395,N_16176);
or U19252 (N_19252,N_16001,N_15064);
nor U19253 (N_19253,N_15340,N_16864);
and U19254 (N_19254,N_15620,N_16125);
and U19255 (N_19255,N_16531,N_15380);
nor U19256 (N_19256,N_16704,N_16311);
nor U19257 (N_19257,N_17360,N_16760);
xor U19258 (N_19258,N_17046,N_16313);
or U19259 (N_19259,N_15949,N_17033);
and U19260 (N_19260,N_15423,N_16903);
and U19261 (N_19261,N_15995,N_15623);
nor U19262 (N_19262,N_15667,N_17376);
nor U19263 (N_19263,N_17480,N_16230);
and U19264 (N_19264,N_16807,N_16913);
or U19265 (N_19265,N_15847,N_17199);
or U19266 (N_19266,N_16060,N_15570);
and U19267 (N_19267,N_15701,N_15172);
or U19268 (N_19268,N_16347,N_15266);
nand U19269 (N_19269,N_15793,N_16296);
xor U19270 (N_19270,N_16291,N_17363);
and U19271 (N_19271,N_15824,N_15539);
and U19272 (N_19272,N_15959,N_16830);
and U19273 (N_19273,N_15580,N_15415);
nand U19274 (N_19274,N_16507,N_16470);
or U19275 (N_19275,N_15390,N_17466);
nor U19276 (N_19276,N_15061,N_16127);
or U19277 (N_19277,N_17381,N_16579);
and U19278 (N_19278,N_17334,N_16263);
and U19279 (N_19279,N_17435,N_16160);
nand U19280 (N_19280,N_16643,N_15651);
and U19281 (N_19281,N_16936,N_15893);
nor U19282 (N_19282,N_16516,N_15308);
and U19283 (N_19283,N_15825,N_15681);
or U19284 (N_19284,N_16257,N_17113);
or U19285 (N_19285,N_17109,N_17156);
nor U19286 (N_19286,N_15406,N_15217);
nand U19287 (N_19287,N_16503,N_17283);
or U19288 (N_19288,N_15359,N_17219);
or U19289 (N_19289,N_16608,N_16765);
and U19290 (N_19290,N_16147,N_15708);
nand U19291 (N_19291,N_16600,N_16650);
nand U19292 (N_19292,N_15780,N_17228);
nand U19293 (N_19293,N_16930,N_15553);
nand U19294 (N_19294,N_16484,N_15775);
nor U19295 (N_19295,N_17153,N_15318);
or U19296 (N_19296,N_16757,N_16533);
and U19297 (N_19297,N_16767,N_16048);
or U19298 (N_19298,N_15134,N_16678);
or U19299 (N_19299,N_15522,N_15437);
nor U19300 (N_19300,N_16622,N_16983);
nor U19301 (N_19301,N_15949,N_15705);
or U19302 (N_19302,N_15980,N_16035);
nand U19303 (N_19303,N_15866,N_15164);
and U19304 (N_19304,N_15729,N_15401);
or U19305 (N_19305,N_17323,N_15470);
and U19306 (N_19306,N_17307,N_16558);
nand U19307 (N_19307,N_16088,N_17437);
nor U19308 (N_19308,N_17419,N_15993);
nand U19309 (N_19309,N_17257,N_17106);
or U19310 (N_19310,N_16249,N_15186);
and U19311 (N_19311,N_15560,N_15809);
nand U19312 (N_19312,N_17226,N_15198);
xnor U19313 (N_19313,N_16140,N_15034);
nand U19314 (N_19314,N_15103,N_15390);
and U19315 (N_19315,N_15850,N_15669);
or U19316 (N_19316,N_15405,N_16473);
nand U19317 (N_19317,N_16971,N_16805);
nor U19318 (N_19318,N_17410,N_17402);
nor U19319 (N_19319,N_15487,N_17048);
and U19320 (N_19320,N_15668,N_15014);
or U19321 (N_19321,N_15039,N_16402);
or U19322 (N_19322,N_17361,N_15948);
nand U19323 (N_19323,N_16892,N_17479);
nand U19324 (N_19324,N_17312,N_16728);
nand U19325 (N_19325,N_15580,N_15197);
nor U19326 (N_19326,N_15569,N_15748);
or U19327 (N_19327,N_17313,N_17184);
nand U19328 (N_19328,N_15408,N_15246);
nor U19329 (N_19329,N_16854,N_16584);
nor U19330 (N_19330,N_15791,N_17253);
nor U19331 (N_19331,N_16239,N_16281);
nor U19332 (N_19332,N_17479,N_15140);
nor U19333 (N_19333,N_15989,N_16342);
and U19334 (N_19334,N_15431,N_15508);
and U19335 (N_19335,N_17208,N_15323);
and U19336 (N_19336,N_17345,N_17459);
and U19337 (N_19337,N_15481,N_16598);
and U19338 (N_19338,N_16207,N_16874);
nor U19339 (N_19339,N_17298,N_15601);
nor U19340 (N_19340,N_16131,N_15884);
or U19341 (N_19341,N_15128,N_16586);
nor U19342 (N_19342,N_17381,N_17337);
nand U19343 (N_19343,N_15637,N_17080);
nor U19344 (N_19344,N_15786,N_17369);
nor U19345 (N_19345,N_16719,N_16502);
nand U19346 (N_19346,N_16162,N_15871);
or U19347 (N_19347,N_15543,N_16855);
and U19348 (N_19348,N_16955,N_16975);
nand U19349 (N_19349,N_16003,N_15224);
nor U19350 (N_19350,N_15243,N_17493);
nor U19351 (N_19351,N_15415,N_15499);
nor U19352 (N_19352,N_16154,N_15219);
and U19353 (N_19353,N_15376,N_17181);
or U19354 (N_19354,N_16012,N_16432);
or U19355 (N_19355,N_15012,N_15518);
nor U19356 (N_19356,N_15498,N_15543);
and U19357 (N_19357,N_15664,N_15963);
or U19358 (N_19358,N_15244,N_15906);
or U19359 (N_19359,N_16278,N_15645);
nor U19360 (N_19360,N_15719,N_16019);
nand U19361 (N_19361,N_17054,N_16752);
or U19362 (N_19362,N_15840,N_16960);
and U19363 (N_19363,N_15112,N_15730);
and U19364 (N_19364,N_17492,N_15739);
and U19365 (N_19365,N_16385,N_15931);
nand U19366 (N_19366,N_15390,N_17384);
nand U19367 (N_19367,N_17043,N_15291);
or U19368 (N_19368,N_16695,N_16107);
or U19369 (N_19369,N_16405,N_16380);
nand U19370 (N_19370,N_15831,N_17084);
and U19371 (N_19371,N_17085,N_15697);
nand U19372 (N_19372,N_17369,N_16957);
nand U19373 (N_19373,N_15342,N_17289);
nor U19374 (N_19374,N_16541,N_17381);
and U19375 (N_19375,N_16722,N_16931);
nand U19376 (N_19376,N_15811,N_15175);
nand U19377 (N_19377,N_17313,N_17281);
nand U19378 (N_19378,N_15025,N_15651);
and U19379 (N_19379,N_15060,N_16609);
or U19380 (N_19380,N_17451,N_17383);
or U19381 (N_19381,N_17204,N_16595);
nor U19382 (N_19382,N_15341,N_16798);
nand U19383 (N_19383,N_16325,N_16356);
or U19384 (N_19384,N_17004,N_17414);
nand U19385 (N_19385,N_16941,N_16295);
nor U19386 (N_19386,N_17073,N_16887);
or U19387 (N_19387,N_16121,N_15746);
or U19388 (N_19388,N_17297,N_16081);
and U19389 (N_19389,N_15149,N_15522);
nor U19390 (N_19390,N_15528,N_17095);
and U19391 (N_19391,N_15144,N_16512);
nand U19392 (N_19392,N_15423,N_16038);
and U19393 (N_19393,N_16282,N_17226);
nor U19394 (N_19394,N_16437,N_16320);
or U19395 (N_19395,N_17405,N_15953);
or U19396 (N_19396,N_15707,N_15278);
nand U19397 (N_19397,N_17186,N_15061);
nor U19398 (N_19398,N_15107,N_15608);
and U19399 (N_19399,N_16144,N_15117);
nor U19400 (N_19400,N_15944,N_16657);
or U19401 (N_19401,N_15558,N_15087);
or U19402 (N_19402,N_15908,N_17044);
and U19403 (N_19403,N_15341,N_16070);
xnor U19404 (N_19404,N_17486,N_15869);
nor U19405 (N_19405,N_16540,N_15126);
or U19406 (N_19406,N_16206,N_15335);
and U19407 (N_19407,N_16325,N_17072);
nand U19408 (N_19408,N_16026,N_15586);
and U19409 (N_19409,N_15985,N_17481);
or U19410 (N_19410,N_15578,N_16001);
and U19411 (N_19411,N_17428,N_16484);
nor U19412 (N_19412,N_15090,N_15290);
or U19413 (N_19413,N_16180,N_17179);
nor U19414 (N_19414,N_16299,N_16349);
nand U19415 (N_19415,N_15363,N_17403);
nor U19416 (N_19416,N_16071,N_16896);
nor U19417 (N_19417,N_15903,N_15895);
nor U19418 (N_19418,N_15300,N_17299);
nand U19419 (N_19419,N_15613,N_16703);
and U19420 (N_19420,N_16684,N_16744);
and U19421 (N_19421,N_15281,N_15186);
nor U19422 (N_19422,N_16105,N_16760);
or U19423 (N_19423,N_15401,N_16077);
nand U19424 (N_19424,N_15450,N_15090);
or U19425 (N_19425,N_15243,N_15917);
nor U19426 (N_19426,N_16042,N_15234);
nand U19427 (N_19427,N_16332,N_17375);
nor U19428 (N_19428,N_17436,N_16218);
nand U19429 (N_19429,N_15069,N_16750);
nand U19430 (N_19430,N_15717,N_17495);
and U19431 (N_19431,N_15792,N_15580);
nor U19432 (N_19432,N_15607,N_17058);
xor U19433 (N_19433,N_17359,N_16470);
nand U19434 (N_19434,N_16506,N_16127);
and U19435 (N_19435,N_15795,N_15539);
or U19436 (N_19436,N_17220,N_16494);
and U19437 (N_19437,N_15650,N_17051);
or U19438 (N_19438,N_15262,N_15166);
xnor U19439 (N_19439,N_15229,N_16320);
nand U19440 (N_19440,N_16294,N_15480);
nor U19441 (N_19441,N_15192,N_15945);
nor U19442 (N_19442,N_16256,N_16206);
nand U19443 (N_19443,N_17274,N_16169);
and U19444 (N_19444,N_15339,N_16425);
nor U19445 (N_19445,N_16762,N_15171);
nand U19446 (N_19446,N_15691,N_17130);
nor U19447 (N_19447,N_16679,N_17305);
and U19448 (N_19448,N_16039,N_17369);
nor U19449 (N_19449,N_16165,N_15112);
nand U19450 (N_19450,N_16942,N_17351);
nand U19451 (N_19451,N_15557,N_15562);
and U19452 (N_19452,N_17030,N_15809);
nand U19453 (N_19453,N_16598,N_16127);
nor U19454 (N_19454,N_17239,N_15139);
and U19455 (N_19455,N_16656,N_16786);
or U19456 (N_19456,N_17416,N_15781);
and U19457 (N_19457,N_16475,N_15275);
nor U19458 (N_19458,N_16775,N_17035);
nand U19459 (N_19459,N_15207,N_17119);
and U19460 (N_19460,N_15243,N_16096);
or U19461 (N_19461,N_16853,N_17251);
or U19462 (N_19462,N_15207,N_16338);
or U19463 (N_19463,N_15752,N_17425);
and U19464 (N_19464,N_17331,N_16482);
nor U19465 (N_19465,N_17289,N_17422);
and U19466 (N_19466,N_16899,N_15321);
and U19467 (N_19467,N_15584,N_16733);
nor U19468 (N_19468,N_16355,N_17056);
or U19469 (N_19469,N_15274,N_17191);
and U19470 (N_19470,N_17189,N_16118);
and U19471 (N_19471,N_17123,N_15603);
nor U19472 (N_19472,N_15165,N_15683);
nand U19473 (N_19473,N_16939,N_15150);
nor U19474 (N_19474,N_17416,N_16754);
and U19475 (N_19475,N_16314,N_15104);
nor U19476 (N_19476,N_16869,N_15847);
nand U19477 (N_19477,N_16264,N_16088);
and U19478 (N_19478,N_16898,N_15413);
or U19479 (N_19479,N_17323,N_15676);
or U19480 (N_19480,N_15597,N_17050);
xor U19481 (N_19481,N_16820,N_15515);
nand U19482 (N_19482,N_15200,N_16993);
or U19483 (N_19483,N_15498,N_16827);
and U19484 (N_19484,N_15699,N_16802);
nor U19485 (N_19485,N_16545,N_16600);
nor U19486 (N_19486,N_15906,N_16084);
or U19487 (N_19487,N_17283,N_17109);
or U19488 (N_19488,N_16432,N_16100);
or U19489 (N_19489,N_15625,N_15488);
nor U19490 (N_19490,N_17499,N_16665);
and U19491 (N_19491,N_15344,N_17229);
nand U19492 (N_19492,N_16245,N_16801);
and U19493 (N_19493,N_16709,N_16963);
and U19494 (N_19494,N_15381,N_15371);
and U19495 (N_19495,N_15229,N_16075);
nor U19496 (N_19496,N_16531,N_15838);
nand U19497 (N_19497,N_15744,N_16664);
nand U19498 (N_19498,N_15895,N_17140);
and U19499 (N_19499,N_17437,N_15509);
xor U19500 (N_19500,N_16623,N_15332);
and U19501 (N_19501,N_15531,N_15005);
and U19502 (N_19502,N_16792,N_16081);
and U19503 (N_19503,N_16222,N_17170);
nor U19504 (N_19504,N_15543,N_16334);
or U19505 (N_19505,N_16071,N_17319);
xor U19506 (N_19506,N_17142,N_16285);
or U19507 (N_19507,N_17411,N_16329);
or U19508 (N_19508,N_16401,N_16169);
xnor U19509 (N_19509,N_16896,N_15936);
nor U19510 (N_19510,N_16013,N_15528);
and U19511 (N_19511,N_15377,N_16601);
or U19512 (N_19512,N_16584,N_16236);
or U19513 (N_19513,N_17360,N_16538);
nor U19514 (N_19514,N_15133,N_15502);
nor U19515 (N_19515,N_17055,N_16999);
or U19516 (N_19516,N_16543,N_17265);
nor U19517 (N_19517,N_15700,N_17245);
or U19518 (N_19518,N_16330,N_16185);
or U19519 (N_19519,N_15370,N_15896);
and U19520 (N_19520,N_15098,N_16290);
or U19521 (N_19521,N_16775,N_15061);
and U19522 (N_19522,N_17272,N_15277);
nor U19523 (N_19523,N_16892,N_15131);
nand U19524 (N_19524,N_15779,N_16195);
and U19525 (N_19525,N_16303,N_16664);
or U19526 (N_19526,N_16208,N_16945);
and U19527 (N_19527,N_17346,N_16571);
nor U19528 (N_19528,N_16085,N_16580);
nor U19529 (N_19529,N_15035,N_17373);
nand U19530 (N_19530,N_16759,N_15224);
and U19531 (N_19531,N_16535,N_16819);
and U19532 (N_19532,N_15642,N_16060);
and U19533 (N_19533,N_17472,N_15095);
nand U19534 (N_19534,N_17073,N_16920);
nor U19535 (N_19535,N_16468,N_16908);
nor U19536 (N_19536,N_15302,N_15412);
and U19537 (N_19537,N_16893,N_16632);
or U19538 (N_19538,N_15501,N_15190);
or U19539 (N_19539,N_16074,N_17149);
or U19540 (N_19540,N_16076,N_16799);
or U19541 (N_19541,N_15656,N_16675);
or U19542 (N_19542,N_16555,N_15665);
nor U19543 (N_19543,N_16376,N_16965);
or U19544 (N_19544,N_16334,N_15772);
and U19545 (N_19545,N_15688,N_17306);
nand U19546 (N_19546,N_17343,N_15327);
and U19547 (N_19547,N_15948,N_17484);
or U19548 (N_19548,N_17131,N_15775);
and U19549 (N_19549,N_15790,N_15785);
or U19550 (N_19550,N_15496,N_16802);
or U19551 (N_19551,N_15176,N_16809);
or U19552 (N_19552,N_15794,N_15821);
and U19553 (N_19553,N_16427,N_17246);
and U19554 (N_19554,N_16595,N_15271);
nor U19555 (N_19555,N_15816,N_15513);
or U19556 (N_19556,N_15706,N_15465);
nor U19557 (N_19557,N_15110,N_15926);
nor U19558 (N_19558,N_16049,N_17282);
nand U19559 (N_19559,N_15302,N_15031);
nand U19560 (N_19560,N_15416,N_16646);
and U19561 (N_19561,N_16894,N_16343);
or U19562 (N_19562,N_15702,N_17158);
or U19563 (N_19563,N_17167,N_16319);
or U19564 (N_19564,N_16801,N_17420);
and U19565 (N_19565,N_15103,N_15408);
or U19566 (N_19566,N_15996,N_15870);
nand U19567 (N_19567,N_16394,N_16203);
and U19568 (N_19568,N_16905,N_16350);
nand U19569 (N_19569,N_17069,N_17084);
or U19570 (N_19570,N_15682,N_15035);
or U19571 (N_19571,N_15368,N_17388);
and U19572 (N_19572,N_16225,N_16411);
nor U19573 (N_19573,N_16024,N_16759);
nor U19574 (N_19574,N_17093,N_16195);
or U19575 (N_19575,N_16269,N_16210);
nand U19576 (N_19576,N_16724,N_17461);
or U19577 (N_19577,N_15678,N_16369);
and U19578 (N_19578,N_16350,N_17052);
nor U19579 (N_19579,N_15662,N_15562);
nor U19580 (N_19580,N_16387,N_16029);
nand U19581 (N_19581,N_16106,N_15219);
and U19582 (N_19582,N_17433,N_17046);
nor U19583 (N_19583,N_17387,N_15911);
nand U19584 (N_19584,N_17348,N_15591);
and U19585 (N_19585,N_17115,N_15465);
or U19586 (N_19586,N_17128,N_16765);
nor U19587 (N_19587,N_16005,N_16976);
nand U19588 (N_19588,N_15181,N_16438);
or U19589 (N_19589,N_15358,N_16509);
or U19590 (N_19590,N_16631,N_15720);
nor U19591 (N_19591,N_16389,N_17369);
and U19592 (N_19592,N_15586,N_17134);
xnor U19593 (N_19593,N_15061,N_15937);
nand U19594 (N_19594,N_15932,N_16427);
nand U19595 (N_19595,N_17322,N_15389);
nor U19596 (N_19596,N_15270,N_15552);
nand U19597 (N_19597,N_17106,N_15068);
and U19598 (N_19598,N_17230,N_16927);
or U19599 (N_19599,N_17198,N_17358);
or U19600 (N_19600,N_15745,N_15548);
nor U19601 (N_19601,N_16936,N_15202);
or U19602 (N_19602,N_15871,N_15793);
nand U19603 (N_19603,N_15021,N_16794);
nor U19604 (N_19604,N_15192,N_16159);
or U19605 (N_19605,N_16567,N_16330);
nand U19606 (N_19606,N_15780,N_15172);
nand U19607 (N_19607,N_16620,N_17214);
or U19608 (N_19608,N_16736,N_15407);
nand U19609 (N_19609,N_15058,N_15700);
nor U19610 (N_19610,N_15631,N_15959);
nand U19611 (N_19611,N_15879,N_17299);
nand U19612 (N_19612,N_15165,N_16138);
nor U19613 (N_19613,N_16990,N_17199);
nand U19614 (N_19614,N_17334,N_16065);
and U19615 (N_19615,N_15002,N_15776);
and U19616 (N_19616,N_17089,N_15145);
and U19617 (N_19617,N_15323,N_15355);
nor U19618 (N_19618,N_15785,N_16014);
xor U19619 (N_19619,N_16960,N_16118);
or U19620 (N_19620,N_17226,N_16001);
or U19621 (N_19621,N_16744,N_16171);
and U19622 (N_19622,N_15564,N_17358);
or U19623 (N_19623,N_16384,N_16918);
and U19624 (N_19624,N_15321,N_15560);
and U19625 (N_19625,N_15131,N_15648);
and U19626 (N_19626,N_17348,N_17130);
nand U19627 (N_19627,N_15162,N_16942);
nand U19628 (N_19628,N_17259,N_17479);
nor U19629 (N_19629,N_15611,N_16545);
and U19630 (N_19630,N_15778,N_15136);
nand U19631 (N_19631,N_15613,N_15935);
and U19632 (N_19632,N_16330,N_15085);
nand U19633 (N_19633,N_16187,N_15412);
nor U19634 (N_19634,N_16013,N_15147);
nand U19635 (N_19635,N_15640,N_16333);
nor U19636 (N_19636,N_16518,N_15277);
nand U19637 (N_19637,N_15026,N_16492);
nor U19638 (N_19638,N_15961,N_16061);
nand U19639 (N_19639,N_17347,N_17031);
and U19640 (N_19640,N_16933,N_15213);
or U19641 (N_19641,N_15272,N_16969);
nand U19642 (N_19642,N_15504,N_15694);
nor U19643 (N_19643,N_15155,N_16836);
or U19644 (N_19644,N_15434,N_16335);
or U19645 (N_19645,N_15961,N_16518);
nor U19646 (N_19646,N_16905,N_15830);
nor U19647 (N_19647,N_16629,N_16546);
and U19648 (N_19648,N_17226,N_15238);
nand U19649 (N_19649,N_15466,N_16798);
nor U19650 (N_19650,N_15187,N_17217);
nor U19651 (N_19651,N_16310,N_15648);
xor U19652 (N_19652,N_16451,N_17255);
nand U19653 (N_19653,N_16696,N_16200);
and U19654 (N_19654,N_15880,N_16188);
nand U19655 (N_19655,N_16231,N_16725);
xnor U19656 (N_19656,N_15779,N_15603);
or U19657 (N_19657,N_16842,N_15196);
or U19658 (N_19658,N_16424,N_15954);
and U19659 (N_19659,N_16655,N_17459);
nand U19660 (N_19660,N_17250,N_15417);
nand U19661 (N_19661,N_17095,N_15930);
and U19662 (N_19662,N_16756,N_15312);
nand U19663 (N_19663,N_17188,N_15281);
or U19664 (N_19664,N_15898,N_16687);
or U19665 (N_19665,N_15054,N_16565);
nor U19666 (N_19666,N_17197,N_17435);
and U19667 (N_19667,N_17186,N_16000);
nor U19668 (N_19668,N_16853,N_17129);
nand U19669 (N_19669,N_15159,N_16633);
nand U19670 (N_19670,N_16747,N_15098);
nand U19671 (N_19671,N_15742,N_15635);
nor U19672 (N_19672,N_16181,N_15499);
nand U19673 (N_19673,N_17219,N_15762);
nor U19674 (N_19674,N_15368,N_16197);
and U19675 (N_19675,N_16799,N_15348);
nor U19676 (N_19676,N_15705,N_16777);
and U19677 (N_19677,N_17268,N_15945);
and U19678 (N_19678,N_15503,N_15371);
nor U19679 (N_19679,N_16918,N_15992);
and U19680 (N_19680,N_17103,N_15087);
or U19681 (N_19681,N_15000,N_16499);
nand U19682 (N_19682,N_15696,N_16980);
nand U19683 (N_19683,N_15769,N_17234);
and U19684 (N_19684,N_15155,N_16921);
or U19685 (N_19685,N_15136,N_17052);
nand U19686 (N_19686,N_16571,N_16264);
nand U19687 (N_19687,N_16902,N_16748);
nand U19688 (N_19688,N_15468,N_17333);
or U19689 (N_19689,N_15060,N_15684);
nor U19690 (N_19690,N_16843,N_15607);
nor U19691 (N_19691,N_17016,N_17214);
and U19692 (N_19692,N_17438,N_15782);
nand U19693 (N_19693,N_17058,N_17431);
nand U19694 (N_19694,N_15450,N_17396);
and U19695 (N_19695,N_17251,N_15653);
nand U19696 (N_19696,N_16390,N_15504);
and U19697 (N_19697,N_15071,N_15180);
nor U19698 (N_19698,N_17409,N_16382);
and U19699 (N_19699,N_16669,N_17057);
and U19700 (N_19700,N_16979,N_15235);
nand U19701 (N_19701,N_15173,N_15096);
nand U19702 (N_19702,N_16881,N_17008);
nor U19703 (N_19703,N_17049,N_15943);
nor U19704 (N_19704,N_16487,N_16643);
nor U19705 (N_19705,N_16724,N_17332);
nor U19706 (N_19706,N_15955,N_15764);
nor U19707 (N_19707,N_16373,N_15879);
nand U19708 (N_19708,N_16430,N_15474);
and U19709 (N_19709,N_16520,N_17379);
or U19710 (N_19710,N_16370,N_16977);
and U19711 (N_19711,N_15022,N_17398);
nand U19712 (N_19712,N_16415,N_17151);
nor U19713 (N_19713,N_16884,N_15215);
nor U19714 (N_19714,N_17162,N_17038);
nor U19715 (N_19715,N_16406,N_16793);
or U19716 (N_19716,N_16732,N_17332);
or U19717 (N_19717,N_17165,N_15141);
nor U19718 (N_19718,N_16237,N_16057);
or U19719 (N_19719,N_17400,N_16850);
or U19720 (N_19720,N_16891,N_16907);
nand U19721 (N_19721,N_15074,N_16669);
and U19722 (N_19722,N_17287,N_15403);
or U19723 (N_19723,N_17271,N_17147);
nor U19724 (N_19724,N_16713,N_15053);
and U19725 (N_19725,N_16353,N_15084);
xor U19726 (N_19726,N_16881,N_15960);
nand U19727 (N_19727,N_17208,N_15292);
or U19728 (N_19728,N_15981,N_16415);
nand U19729 (N_19729,N_17087,N_16108);
or U19730 (N_19730,N_16710,N_15798);
nor U19731 (N_19731,N_15440,N_15728);
xnor U19732 (N_19732,N_15624,N_15455);
nor U19733 (N_19733,N_16949,N_15061);
or U19734 (N_19734,N_17302,N_15648);
nor U19735 (N_19735,N_15885,N_17248);
nor U19736 (N_19736,N_16971,N_15938);
or U19737 (N_19737,N_16660,N_17333);
and U19738 (N_19738,N_15824,N_16735);
or U19739 (N_19739,N_15279,N_16103);
nand U19740 (N_19740,N_16607,N_16971);
or U19741 (N_19741,N_16083,N_16108);
nor U19742 (N_19742,N_16994,N_17311);
and U19743 (N_19743,N_17174,N_15783);
nor U19744 (N_19744,N_15660,N_16439);
and U19745 (N_19745,N_16692,N_17366);
or U19746 (N_19746,N_16341,N_16578);
nand U19747 (N_19747,N_15935,N_15375);
or U19748 (N_19748,N_16510,N_16666);
nor U19749 (N_19749,N_15092,N_16282);
xor U19750 (N_19750,N_15131,N_16823);
nand U19751 (N_19751,N_16098,N_15907);
xnor U19752 (N_19752,N_15557,N_15086);
nand U19753 (N_19753,N_15937,N_15458);
nand U19754 (N_19754,N_15888,N_16998);
and U19755 (N_19755,N_15213,N_16432);
or U19756 (N_19756,N_16944,N_16038);
and U19757 (N_19757,N_16164,N_17450);
nand U19758 (N_19758,N_16152,N_17218);
and U19759 (N_19759,N_15438,N_15015);
xnor U19760 (N_19760,N_15249,N_16021);
nand U19761 (N_19761,N_15719,N_16138);
and U19762 (N_19762,N_16146,N_16404);
and U19763 (N_19763,N_15198,N_16658);
or U19764 (N_19764,N_15126,N_15937);
and U19765 (N_19765,N_15159,N_15833);
nand U19766 (N_19766,N_16367,N_16272);
and U19767 (N_19767,N_17351,N_16432);
nand U19768 (N_19768,N_15789,N_17159);
xnor U19769 (N_19769,N_15067,N_17223);
nand U19770 (N_19770,N_16853,N_15278);
nand U19771 (N_19771,N_15561,N_16386);
nand U19772 (N_19772,N_15129,N_15420);
nand U19773 (N_19773,N_17300,N_17253);
nand U19774 (N_19774,N_16551,N_16359);
or U19775 (N_19775,N_16786,N_17439);
nor U19776 (N_19776,N_16812,N_15407);
and U19777 (N_19777,N_16082,N_17377);
and U19778 (N_19778,N_17450,N_16903);
or U19779 (N_19779,N_16533,N_15553);
or U19780 (N_19780,N_16430,N_15023);
nor U19781 (N_19781,N_16179,N_15543);
or U19782 (N_19782,N_17159,N_16399);
and U19783 (N_19783,N_16508,N_16197);
nor U19784 (N_19784,N_16546,N_15030);
xnor U19785 (N_19785,N_15967,N_16396);
and U19786 (N_19786,N_16701,N_16168);
nor U19787 (N_19787,N_16404,N_16333);
or U19788 (N_19788,N_15982,N_16332);
nor U19789 (N_19789,N_16314,N_16289);
nor U19790 (N_19790,N_16895,N_17368);
nand U19791 (N_19791,N_15807,N_15878);
nand U19792 (N_19792,N_15809,N_15980);
or U19793 (N_19793,N_17125,N_16163);
or U19794 (N_19794,N_15039,N_16512);
nand U19795 (N_19795,N_15668,N_15008);
nand U19796 (N_19796,N_15564,N_16634);
and U19797 (N_19797,N_16473,N_16406);
nor U19798 (N_19798,N_16961,N_16953);
nor U19799 (N_19799,N_15125,N_15390);
nand U19800 (N_19800,N_15920,N_15010);
or U19801 (N_19801,N_17346,N_15379);
or U19802 (N_19802,N_15248,N_15060);
and U19803 (N_19803,N_15017,N_15299);
nand U19804 (N_19804,N_15625,N_17274);
nand U19805 (N_19805,N_17145,N_15450);
and U19806 (N_19806,N_15396,N_16721);
nand U19807 (N_19807,N_16541,N_16549);
and U19808 (N_19808,N_17203,N_17252);
nand U19809 (N_19809,N_16564,N_15883);
or U19810 (N_19810,N_17034,N_15819);
nor U19811 (N_19811,N_15237,N_15136);
or U19812 (N_19812,N_17446,N_16407);
nor U19813 (N_19813,N_15048,N_15026);
or U19814 (N_19814,N_15986,N_15082);
nor U19815 (N_19815,N_16338,N_16138);
nor U19816 (N_19816,N_15706,N_16444);
or U19817 (N_19817,N_15993,N_17377);
nor U19818 (N_19818,N_15147,N_16485);
nand U19819 (N_19819,N_17219,N_15164);
nand U19820 (N_19820,N_17042,N_16131);
nand U19821 (N_19821,N_16783,N_15442);
nor U19822 (N_19822,N_16882,N_15350);
or U19823 (N_19823,N_16332,N_15909);
and U19824 (N_19824,N_17415,N_16407);
or U19825 (N_19825,N_16661,N_15532);
nor U19826 (N_19826,N_17339,N_15075);
nor U19827 (N_19827,N_15329,N_15033);
nand U19828 (N_19828,N_16582,N_15776);
nor U19829 (N_19829,N_17388,N_16219);
nand U19830 (N_19830,N_17208,N_16798);
nor U19831 (N_19831,N_16375,N_17182);
nor U19832 (N_19832,N_16690,N_15451);
xnor U19833 (N_19833,N_17054,N_16188);
or U19834 (N_19834,N_16032,N_17011);
and U19835 (N_19835,N_15750,N_16339);
or U19836 (N_19836,N_16386,N_15900);
nor U19837 (N_19837,N_15726,N_15419);
and U19838 (N_19838,N_15573,N_17364);
or U19839 (N_19839,N_15073,N_16110);
or U19840 (N_19840,N_15526,N_15055);
nor U19841 (N_19841,N_15159,N_16786);
nor U19842 (N_19842,N_15155,N_15509);
nand U19843 (N_19843,N_16901,N_16617);
and U19844 (N_19844,N_16022,N_16530);
nand U19845 (N_19845,N_15251,N_15921);
or U19846 (N_19846,N_16091,N_17236);
and U19847 (N_19847,N_17088,N_15928);
nor U19848 (N_19848,N_16630,N_16704);
or U19849 (N_19849,N_15740,N_16247);
nand U19850 (N_19850,N_16825,N_16434);
nor U19851 (N_19851,N_16942,N_15497);
or U19852 (N_19852,N_17334,N_16397);
or U19853 (N_19853,N_16193,N_17358);
or U19854 (N_19854,N_17047,N_17347);
or U19855 (N_19855,N_16664,N_17193);
and U19856 (N_19856,N_16749,N_15369);
nand U19857 (N_19857,N_16819,N_17110);
and U19858 (N_19858,N_17203,N_16409);
and U19859 (N_19859,N_16931,N_15164);
or U19860 (N_19860,N_16275,N_17479);
or U19861 (N_19861,N_16563,N_15049);
and U19862 (N_19862,N_17291,N_15233);
or U19863 (N_19863,N_15493,N_16383);
nand U19864 (N_19864,N_15907,N_15369);
nand U19865 (N_19865,N_17370,N_17153);
and U19866 (N_19866,N_17389,N_15848);
or U19867 (N_19867,N_16693,N_16927);
or U19868 (N_19868,N_16964,N_15167);
xor U19869 (N_19869,N_15810,N_17351);
and U19870 (N_19870,N_17335,N_16863);
nand U19871 (N_19871,N_15992,N_16105);
nand U19872 (N_19872,N_16907,N_15560);
nor U19873 (N_19873,N_17487,N_15879);
and U19874 (N_19874,N_16594,N_17351);
nand U19875 (N_19875,N_15606,N_16589);
nand U19876 (N_19876,N_15500,N_16267);
nor U19877 (N_19877,N_16942,N_15709);
nor U19878 (N_19878,N_17411,N_15353);
nand U19879 (N_19879,N_15174,N_16857);
and U19880 (N_19880,N_16167,N_15007);
or U19881 (N_19881,N_16944,N_15237);
nor U19882 (N_19882,N_17402,N_15638);
and U19883 (N_19883,N_17212,N_15587);
and U19884 (N_19884,N_17493,N_15786);
nand U19885 (N_19885,N_16516,N_16813);
nand U19886 (N_19886,N_15857,N_16915);
xnor U19887 (N_19887,N_17080,N_17020);
nor U19888 (N_19888,N_16958,N_15017);
nand U19889 (N_19889,N_17492,N_15713);
nand U19890 (N_19890,N_16438,N_15930);
or U19891 (N_19891,N_15221,N_15618);
nand U19892 (N_19892,N_15539,N_15826);
nand U19893 (N_19893,N_15952,N_15379);
or U19894 (N_19894,N_16591,N_17318);
or U19895 (N_19895,N_15786,N_16375);
or U19896 (N_19896,N_15183,N_17045);
or U19897 (N_19897,N_15082,N_15896);
nor U19898 (N_19898,N_15590,N_17248);
and U19899 (N_19899,N_16246,N_15263);
nand U19900 (N_19900,N_16693,N_15169);
nor U19901 (N_19901,N_16532,N_16742);
nand U19902 (N_19902,N_15834,N_15657);
nor U19903 (N_19903,N_17117,N_16908);
and U19904 (N_19904,N_16427,N_15880);
and U19905 (N_19905,N_16325,N_16823);
or U19906 (N_19906,N_16180,N_15774);
nor U19907 (N_19907,N_17052,N_15918);
and U19908 (N_19908,N_15777,N_15470);
and U19909 (N_19909,N_17115,N_15839);
nand U19910 (N_19910,N_17472,N_17404);
nand U19911 (N_19911,N_15545,N_15492);
nor U19912 (N_19912,N_15974,N_15086);
nand U19913 (N_19913,N_15804,N_15082);
and U19914 (N_19914,N_15261,N_17415);
and U19915 (N_19915,N_15251,N_16763);
nand U19916 (N_19916,N_16758,N_16785);
nor U19917 (N_19917,N_17185,N_15430);
or U19918 (N_19918,N_15789,N_16365);
or U19919 (N_19919,N_15033,N_17438);
or U19920 (N_19920,N_15930,N_16280);
nand U19921 (N_19921,N_16989,N_16299);
nor U19922 (N_19922,N_17002,N_17327);
nand U19923 (N_19923,N_17410,N_15976);
nor U19924 (N_19924,N_15034,N_15978);
nor U19925 (N_19925,N_17162,N_16870);
nand U19926 (N_19926,N_17069,N_16590);
and U19927 (N_19927,N_17247,N_15362);
and U19928 (N_19928,N_16577,N_15939);
nor U19929 (N_19929,N_17095,N_15588);
and U19930 (N_19930,N_17111,N_16979);
nor U19931 (N_19931,N_15350,N_15623);
nand U19932 (N_19932,N_16395,N_15043);
nand U19933 (N_19933,N_16726,N_15401);
nand U19934 (N_19934,N_17387,N_16910);
nand U19935 (N_19935,N_17086,N_17099);
nor U19936 (N_19936,N_16818,N_16121);
nor U19937 (N_19937,N_16982,N_15515);
and U19938 (N_19938,N_15379,N_16939);
nand U19939 (N_19939,N_16341,N_16021);
and U19940 (N_19940,N_15067,N_17428);
and U19941 (N_19941,N_16319,N_16287);
and U19942 (N_19942,N_16879,N_17078);
and U19943 (N_19943,N_17398,N_15794);
nor U19944 (N_19944,N_15343,N_16496);
and U19945 (N_19945,N_17393,N_16065);
nand U19946 (N_19946,N_15096,N_15814);
and U19947 (N_19947,N_16402,N_17165);
and U19948 (N_19948,N_16809,N_16955);
or U19949 (N_19949,N_15409,N_15173);
nor U19950 (N_19950,N_16509,N_16094);
nor U19951 (N_19951,N_16399,N_15509);
nand U19952 (N_19952,N_15192,N_15670);
and U19953 (N_19953,N_16485,N_15164);
and U19954 (N_19954,N_16485,N_16669);
nor U19955 (N_19955,N_16898,N_15598);
or U19956 (N_19956,N_17280,N_17298);
xnor U19957 (N_19957,N_15686,N_15649);
nand U19958 (N_19958,N_15652,N_17244);
and U19959 (N_19959,N_15800,N_15911);
or U19960 (N_19960,N_15646,N_16903);
nor U19961 (N_19961,N_16492,N_16004);
nand U19962 (N_19962,N_17221,N_17354);
nor U19963 (N_19963,N_16604,N_15390);
or U19964 (N_19964,N_15724,N_16606);
nand U19965 (N_19965,N_16241,N_16140);
nand U19966 (N_19966,N_15908,N_17144);
and U19967 (N_19967,N_15741,N_15951);
or U19968 (N_19968,N_15732,N_17084);
nand U19969 (N_19969,N_16846,N_16612);
and U19970 (N_19970,N_15054,N_17223);
or U19971 (N_19971,N_15229,N_15496);
nand U19972 (N_19972,N_16801,N_16248);
nand U19973 (N_19973,N_15068,N_15298);
and U19974 (N_19974,N_17247,N_15508);
nand U19975 (N_19975,N_15846,N_16503);
and U19976 (N_19976,N_16769,N_16765);
and U19977 (N_19977,N_17389,N_15009);
nor U19978 (N_19978,N_15611,N_16678);
nand U19979 (N_19979,N_16672,N_16481);
nor U19980 (N_19980,N_15384,N_16377);
nor U19981 (N_19981,N_16759,N_16540);
nor U19982 (N_19982,N_15280,N_15590);
nand U19983 (N_19983,N_15954,N_17227);
nor U19984 (N_19984,N_17122,N_17430);
nor U19985 (N_19985,N_16626,N_15983);
or U19986 (N_19986,N_15062,N_16064);
xnor U19987 (N_19987,N_15868,N_15831);
and U19988 (N_19988,N_16672,N_17056);
nand U19989 (N_19989,N_15853,N_15632);
and U19990 (N_19990,N_16421,N_16745);
nor U19991 (N_19991,N_16506,N_16515);
and U19992 (N_19992,N_16127,N_17144);
or U19993 (N_19993,N_17390,N_16877);
and U19994 (N_19994,N_16450,N_17489);
and U19995 (N_19995,N_17071,N_16104);
nor U19996 (N_19996,N_16086,N_15750);
nand U19997 (N_19997,N_16566,N_15781);
nor U19998 (N_19998,N_17401,N_16876);
nor U19999 (N_19999,N_16394,N_15306);
nor U20000 (N_20000,N_17920,N_17971);
or U20001 (N_20001,N_19567,N_18622);
nor U20002 (N_20002,N_19236,N_19182);
nor U20003 (N_20003,N_19310,N_17879);
or U20004 (N_20004,N_18572,N_17760);
or U20005 (N_20005,N_19848,N_18555);
or U20006 (N_20006,N_18278,N_19270);
nor U20007 (N_20007,N_18995,N_17703);
and U20008 (N_20008,N_17610,N_19880);
nand U20009 (N_20009,N_18432,N_19554);
nand U20010 (N_20010,N_18292,N_19139);
or U20011 (N_20011,N_17738,N_18894);
nor U20012 (N_20012,N_19418,N_18792);
and U20013 (N_20013,N_18635,N_17652);
or U20014 (N_20014,N_18575,N_18545);
nor U20015 (N_20015,N_17687,N_18322);
or U20016 (N_20016,N_18263,N_18990);
or U20017 (N_20017,N_19950,N_18946);
nand U20018 (N_20018,N_19608,N_18939);
nor U20019 (N_20019,N_17656,N_19108);
or U20020 (N_20020,N_17836,N_18380);
or U20021 (N_20021,N_18436,N_18455);
nand U20022 (N_20022,N_19187,N_18236);
or U20023 (N_20023,N_18513,N_18906);
nand U20024 (N_20024,N_18174,N_19477);
nand U20025 (N_20025,N_17605,N_17705);
nand U20026 (N_20026,N_19250,N_17748);
or U20027 (N_20027,N_19279,N_18066);
nor U20028 (N_20028,N_18962,N_18546);
nand U20029 (N_20029,N_17981,N_18918);
xor U20030 (N_20030,N_18431,N_19438);
or U20031 (N_20031,N_17990,N_19348);
or U20032 (N_20032,N_18003,N_19873);
or U20033 (N_20033,N_18532,N_18331);
nor U20034 (N_20034,N_19160,N_18435);
nand U20035 (N_20035,N_19206,N_17997);
nand U20036 (N_20036,N_18045,N_19266);
nor U20037 (N_20037,N_18330,N_19845);
and U20038 (N_20038,N_18352,N_18379);
nand U20039 (N_20039,N_19213,N_19053);
or U20040 (N_20040,N_17778,N_19753);
or U20041 (N_20041,N_19945,N_19927);
nand U20042 (N_20042,N_17823,N_18320);
and U20043 (N_20043,N_18130,N_17860);
or U20044 (N_20044,N_19530,N_18626);
nand U20045 (N_20045,N_19051,N_19374);
and U20046 (N_20046,N_18531,N_19469);
or U20047 (N_20047,N_18613,N_17507);
nor U20048 (N_20048,N_19178,N_18447);
and U20049 (N_20049,N_19722,N_18863);
nand U20050 (N_20050,N_19289,N_18468);
nor U20051 (N_20051,N_19100,N_18762);
nor U20052 (N_20052,N_17890,N_18599);
nor U20053 (N_20053,N_19508,N_18262);
or U20054 (N_20054,N_19898,N_18820);
nor U20055 (N_20055,N_18516,N_18275);
nor U20056 (N_20056,N_18473,N_17794);
nand U20057 (N_20057,N_19842,N_18344);
and U20058 (N_20058,N_19410,N_18543);
or U20059 (N_20059,N_18267,N_18534);
and U20060 (N_20060,N_18580,N_18654);
and U20061 (N_20061,N_18084,N_18961);
nand U20062 (N_20062,N_19587,N_19037);
or U20063 (N_20063,N_18803,N_19023);
or U20064 (N_20064,N_19937,N_19624);
and U20065 (N_20065,N_17555,N_18073);
or U20066 (N_20066,N_19303,N_19204);
and U20067 (N_20067,N_18249,N_18835);
nand U20068 (N_20068,N_18878,N_19293);
nand U20069 (N_20069,N_17742,N_18289);
nor U20070 (N_20070,N_19866,N_18999);
nand U20071 (N_20071,N_19308,N_19776);
nor U20072 (N_20072,N_17668,N_18602);
nor U20073 (N_20073,N_19474,N_19288);
nand U20074 (N_20074,N_18731,N_18479);
nor U20075 (N_20075,N_17943,N_18807);
and U20076 (N_20076,N_19851,N_18250);
nor U20077 (N_20077,N_18783,N_17887);
and U20078 (N_20078,N_17780,N_19603);
nand U20079 (N_20079,N_18065,N_17775);
nor U20080 (N_20080,N_17945,N_19249);
and U20081 (N_20081,N_19847,N_18884);
nor U20082 (N_20082,N_18472,N_19328);
or U20083 (N_20083,N_17609,N_19292);
nand U20084 (N_20084,N_18858,N_17913);
nand U20085 (N_20085,N_19782,N_18154);
nand U20086 (N_20086,N_17632,N_19315);
nand U20087 (N_20087,N_18893,N_18719);
nor U20088 (N_20088,N_18649,N_19616);
nor U20089 (N_20089,N_17786,N_18035);
nor U20090 (N_20090,N_18897,N_19370);
and U20091 (N_20091,N_19853,N_19179);
nor U20092 (N_20092,N_19617,N_19432);
or U20093 (N_20093,N_19783,N_18218);
and U20094 (N_20094,N_18451,N_19714);
and U20095 (N_20095,N_19985,N_19505);
and U20096 (N_20096,N_18286,N_18606);
or U20097 (N_20097,N_17895,N_18007);
nand U20098 (N_20098,N_19277,N_19844);
nor U20099 (N_20099,N_19883,N_19174);
and U20100 (N_20100,N_17772,N_17639);
or U20101 (N_20101,N_19925,N_19181);
nor U20102 (N_20102,N_18378,N_18509);
or U20103 (N_20103,N_19107,N_18681);
nand U20104 (N_20104,N_19611,N_18216);
and U20105 (N_20105,N_19345,N_19635);
and U20106 (N_20106,N_19124,N_18389);
nand U20107 (N_20107,N_19291,N_18070);
nand U20108 (N_20108,N_19788,N_19045);
or U20109 (N_20109,N_19922,N_18665);
and U20110 (N_20110,N_17935,N_18430);
and U20111 (N_20111,N_18462,N_18709);
or U20112 (N_20112,N_17532,N_19800);
or U20113 (N_20113,N_17807,N_18584);
nor U20114 (N_20114,N_19907,N_18326);
nor U20115 (N_20115,N_19369,N_19614);
nor U20116 (N_20116,N_19669,N_19579);
and U20117 (N_20117,N_18197,N_19425);
or U20118 (N_20118,N_18177,N_19490);
or U20119 (N_20119,N_19994,N_18147);
nor U20120 (N_20120,N_18253,N_18679);
or U20121 (N_20121,N_18283,N_17922);
nor U20122 (N_20122,N_19149,N_19175);
or U20123 (N_20123,N_17741,N_18198);
or U20124 (N_20124,N_19378,N_17592);
and U20125 (N_20125,N_19830,N_19817);
nand U20126 (N_20126,N_17688,N_19522);
nand U20127 (N_20127,N_19426,N_19073);
and U20128 (N_20128,N_19860,N_19736);
nand U20129 (N_20129,N_19028,N_18865);
nand U20130 (N_20130,N_17842,N_18195);
nand U20131 (N_20131,N_19928,N_18520);
nand U20132 (N_20132,N_18176,N_18241);
nor U20133 (N_20133,N_18500,N_18089);
or U20134 (N_20134,N_19271,N_18772);
nor U20135 (N_20135,N_19706,N_18421);
or U20136 (N_20136,N_19365,N_17675);
and U20137 (N_20137,N_18975,N_18202);
nor U20138 (N_20138,N_18490,N_18661);
nor U20139 (N_20139,N_19713,N_19742);
nor U20140 (N_20140,N_18412,N_19029);
or U20141 (N_20141,N_18456,N_18629);
or U20142 (N_20142,N_19155,N_19584);
nor U20143 (N_20143,N_18190,N_18055);
nor U20144 (N_20144,N_19738,N_17865);
or U20145 (N_20145,N_17541,N_17928);
and U20146 (N_20146,N_18640,N_19779);
and U20147 (N_20147,N_18603,N_18439);
or U20148 (N_20148,N_19440,N_19524);
and U20149 (N_20149,N_19699,N_17726);
nor U20150 (N_20150,N_18789,N_17502);
or U20151 (N_20151,N_19083,N_19523);
and U20152 (N_20152,N_18794,N_17663);
and U20153 (N_20153,N_17607,N_18028);
and U20154 (N_20154,N_19599,N_19209);
nor U20155 (N_20155,N_17916,N_18862);
or U20156 (N_20156,N_18644,N_17638);
or U20157 (N_20157,N_19252,N_19919);
or U20158 (N_20158,N_17902,N_18598);
and U20159 (N_20159,N_18301,N_18127);
and U20160 (N_20160,N_17646,N_18419);
nor U20161 (N_20161,N_18461,N_17699);
or U20162 (N_20162,N_18597,N_17702);
or U20163 (N_20163,N_19461,N_17722);
and U20164 (N_20164,N_19493,N_18978);
xnor U20165 (N_20165,N_18014,N_17771);
and U20166 (N_20166,N_19480,N_17736);
nor U20167 (N_20167,N_18312,N_18240);
and U20168 (N_20168,N_19034,N_19887);
nand U20169 (N_20169,N_18033,N_17826);
and U20170 (N_20170,N_19897,N_19006);
nand U20171 (N_20171,N_19752,N_17729);
nand U20172 (N_20172,N_18328,N_19420);
nand U20173 (N_20173,N_17783,N_18778);
or U20174 (N_20174,N_18566,N_17521);
nor U20175 (N_20175,N_18082,N_18837);
and U20176 (N_20176,N_17657,N_18132);
or U20177 (N_20177,N_19543,N_18025);
and U20178 (N_20178,N_18417,N_17658);
nor U20179 (N_20179,N_18487,N_18986);
or U20180 (N_20180,N_18282,N_17882);
or U20181 (N_20181,N_17923,N_19711);
nand U20182 (N_20182,N_18032,N_18185);
and U20183 (N_20183,N_19970,N_18738);
nor U20184 (N_20184,N_18929,N_19122);
and U20185 (N_20185,N_18227,N_18041);
nor U20186 (N_20186,N_19437,N_19721);
nor U20187 (N_20187,N_19105,N_19473);
nor U20188 (N_20188,N_19785,N_19416);
and U20189 (N_20189,N_18392,N_18610);
nand U20190 (N_20190,N_19342,N_19615);
nand U20191 (N_20191,N_19824,N_18518);
nand U20192 (N_20192,N_18735,N_17701);
and U20193 (N_20193,N_19453,N_18887);
nand U20194 (N_20194,N_19217,N_19839);
nor U20195 (N_20195,N_18471,N_19757);
nor U20196 (N_20196,N_19843,N_17975);
nor U20197 (N_20197,N_17861,N_18446);
nor U20198 (N_20198,N_18406,N_18400);
nand U20199 (N_20199,N_18120,N_18433);
nand U20200 (N_20200,N_18579,N_18495);
and U20201 (N_20201,N_19835,N_19192);
nand U20202 (N_20202,N_19668,N_18600);
or U20203 (N_20203,N_17665,N_18036);
and U20204 (N_20204,N_19056,N_18104);
nor U20205 (N_20205,N_17549,N_18601);
nand U20206 (N_20206,N_19991,N_19933);
and U20207 (N_20207,N_19406,N_18424);
nand U20208 (N_20208,N_18034,N_18558);
nor U20209 (N_20209,N_18335,N_18274);
and U20210 (N_20210,N_18113,N_18444);
nor U20211 (N_20211,N_19322,N_19232);
nor U20212 (N_20212,N_18496,N_19156);
or U20213 (N_20213,N_19872,N_17603);
and U20214 (N_20214,N_17968,N_19557);
nand U20215 (N_20215,N_18364,N_18768);
or U20216 (N_20216,N_17613,N_18616);
nand U20217 (N_20217,N_19952,N_18111);
nand U20218 (N_20218,N_18739,N_17561);
nor U20219 (N_20219,N_19899,N_19085);
or U20220 (N_20220,N_19273,N_19309);
nand U20221 (N_20221,N_19349,N_19526);
nor U20222 (N_20222,N_17501,N_17846);
nand U20223 (N_20223,N_19311,N_18022);
or U20224 (N_20224,N_18145,N_18757);
nand U20225 (N_20225,N_18503,N_18058);
and U20226 (N_20226,N_19988,N_17661);
or U20227 (N_20227,N_19906,N_19534);
nand U20228 (N_20228,N_19749,N_18481);
or U20229 (N_20229,N_17801,N_18742);
or U20230 (N_20230,N_17996,N_19093);
and U20231 (N_20231,N_18376,N_19226);
nor U20232 (N_20232,N_17941,N_19072);
or U20233 (N_20233,N_19591,N_17966);
nand U20234 (N_20234,N_18146,N_19704);
nor U20235 (N_20235,N_17531,N_19948);
and U20236 (N_20236,N_18996,N_19185);
nand U20237 (N_20237,N_19459,N_18830);
or U20238 (N_20238,N_18220,N_18829);
and U20239 (N_20239,N_18221,N_19119);
or U20240 (N_20240,N_18623,N_18970);
and U20241 (N_20241,N_19069,N_18729);
nor U20242 (N_20242,N_17550,N_18839);
and U20243 (N_20243,N_19304,N_19816);
or U20244 (N_20244,N_19087,N_19402);
nor U20245 (N_20245,N_18510,N_19917);
nand U20246 (N_20246,N_18779,N_19316);
nand U20247 (N_20247,N_18404,N_17522);
or U20248 (N_20248,N_18697,N_18454);
nor U20249 (N_20249,N_18165,N_17799);
nor U20250 (N_20250,N_19641,N_18402);
or U20251 (N_20251,N_18126,N_19542);
nor U20252 (N_20252,N_19986,N_18491);
and U20253 (N_20253,N_19705,N_18234);
nand U20254 (N_20254,N_17875,N_19483);
or U20255 (N_20255,N_19904,N_19680);
nand U20256 (N_20256,N_17811,N_18838);
nand U20257 (N_20257,N_18269,N_17958);
or U20258 (N_20258,N_19622,N_17690);
nor U20259 (N_20259,N_18016,N_19665);
nand U20260 (N_20260,N_17510,N_18641);
nand U20261 (N_20261,N_19381,N_18337);
nor U20262 (N_20262,N_19797,N_17595);
nor U20263 (N_20263,N_18748,N_18690);
nand U20264 (N_20264,N_17654,N_19081);
nand U20265 (N_20265,N_18909,N_18116);
nand U20266 (N_20266,N_19750,N_18314);
or U20267 (N_20267,N_18067,N_18692);
or U20268 (N_20268,N_18932,N_17999);
or U20269 (N_20269,N_17960,N_18916);
nor U20270 (N_20270,N_17969,N_19772);
or U20271 (N_20271,N_18694,N_18179);
or U20272 (N_20272,N_18426,N_19013);
nand U20273 (N_20273,N_19257,N_19141);
nor U20274 (N_20274,N_17924,N_17641);
nand U20275 (N_20275,N_18215,N_17871);
or U20276 (N_20276,N_19261,N_19215);
and U20277 (N_20277,N_19565,N_18342);
nor U20278 (N_20278,N_19214,N_18828);
nor U20279 (N_20279,N_17535,N_17863);
xor U20280 (N_20280,N_17925,N_18756);
nand U20281 (N_20281,N_17979,N_19334);
or U20282 (N_20282,N_17853,N_18467);
nand U20283 (N_20283,N_17538,N_19900);
nor U20284 (N_20284,N_18955,N_18105);
or U20285 (N_20285,N_17504,N_19339);
nor U20286 (N_20286,N_18798,N_17758);
nand U20287 (N_20287,N_18360,N_18740);
and U20288 (N_20288,N_17708,N_19965);
nor U20289 (N_20289,N_17795,N_18877);
nor U20290 (N_20290,N_17998,N_19696);
nor U20291 (N_20291,N_19022,N_18581);
nand U20292 (N_20292,N_18637,N_17956);
nor U20293 (N_20293,N_18098,N_18853);
or U20294 (N_20294,N_17570,N_18153);
and U20295 (N_20295,N_18158,N_18031);
nor U20296 (N_20296,N_18879,N_18128);
nand U20297 (N_20297,N_18081,N_17844);
and U20298 (N_20298,N_18663,N_19300);
nand U20299 (N_20299,N_19167,N_18268);
or U20300 (N_20300,N_18407,N_19693);
and U20301 (N_20301,N_18137,N_19643);
nor U20302 (N_20302,N_17988,N_19688);
nand U20303 (N_20303,N_18965,N_18046);
and U20304 (N_20304,N_18605,N_19133);
or U20305 (N_20305,N_18166,N_19077);
nand U20306 (N_20306,N_18323,N_19039);
nor U20307 (N_20307,N_18056,N_19092);
and U20308 (N_20308,N_18614,N_17877);
nand U20309 (N_20309,N_18291,N_17528);
nor U20310 (N_20310,N_19755,N_19640);
and U20311 (N_20311,N_18273,N_18733);
nand U20312 (N_20312,N_18437,N_19594);
nand U20313 (N_20313,N_18121,N_19687);
or U20314 (N_20314,N_17757,N_19347);
nor U20315 (N_20315,N_18907,N_19434);
xor U20316 (N_20316,N_17662,N_19208);
or U20317 (N_20317,N_18876,N_19690);
or U20318 (N_20318,N_19126,N_19732);
or U20319 (N_20319,N_19756,N_17822);
or U20320 (N_20320,N_19198,N_19949);
or U20321 (N_20321,N_19487,N_19613);
xor U20322 (N_20322,N_19150,N_17731);
or U20323 (N_20323,N_18673,N_19358);
nand U20324 (N_20324,N_17961,N_18397);
nand U20325 (N_20325,N_18355,N_19313);
and U20326 (N_20326,N_19511,N_17608);
or U20327 (N_20327,N_17914,N_18949);
or U20328 (N_20328,N_19592,N_18152);
nand U20329 (N_20329,N_18134,N_19963);
nand U20330 (N_20330,N_17749,N_18148);
or U20331 (N_20331,N_18464,N_18813);
nor U20332 (N_20332,N_19514,N_17596);
or U20333 (N_20333,N_18560,N_18396);
and U20334 (N_20334,N_19244,N_18325);
nand U20335 (N_20335,N_18948,N_17855);
and U20336 (N_20336,N_18873,N_18085);
or U20337 (N_20337,N_17568,N_18173);
nand U20338 (N_20338,N_19955,N_18911);
and U20339 (N_20339,N_19443,N_18901);
nor U20340 (N_20340,N_18125,N_18213);
nor U20341 (N_20341,N_18724,N_19819);
nor U20342 (N_20342,N_19326,N_18765);
and U20343 (N_20343,N_19216,N_19612);
or U20344 (N_20344,N_18769,N_17536);
or U20345 (N_20345,N_18094,N_18786);
nor U20346 (N_20346,N_19417,N_18280);
or U20347 (N_20347,N_18875,N_18676);
and U20348 (N_20348,N_17830,N_19509);
or U20349 (N_20349,N_19912,N_19810);
or U20350 (N_20350,N_19660,N_18574);
xor U20351 (N_20351,N_19503,N_17972);
or U20352 (N_20352,N_18315,N_19803);
nand U20353 (N_20353,N_17857,N_18339);
or U20354 (N_20354,N_17874,N_19507);
nor U20355 (N_20355,N_18140,N_19692);
xnor U20356 (N_20356,N_19131,N_19791);
or U20357 (N_20357,N_18974,N_19938);
nand U20358 (N_20358,N_17982,N_19058);
nand U20359 (N_20359,N_19106,N_17557);
nor U20360 (N_20360,N_18882,N_19063);
and U20361 (N_20361,N_19829,N_19833);
or U20362 (N_20362,N_19243,N_18488);
nand U20363 (N_20363,N_18504,N_18744);
and U20364 (N_20364,N_18931,N_19778);
and U20365 (N_20365,N_18867,N_19003);
nand U20366 (N_20366,N_18009,N_18167);
or U20367 (N_20367,N_19506,N_17859);
nand U20368 (N_20368,N_18633,N_18141);
and U20369 (N_20369,N_19537,N_17746);
nand U20370 (N_20370,N_18149,N_18874);
or U20371 (N_20371,N_19158,N_18217);
nor U20372 (N_20372,N_19301,N_19993);
and U20373 (N_20373,N_17851,N_19205);
nor U20374 (N_20374,N_19005,N_19637);
and U20375 (N_20375,N_19307,N_17560);
nor U20376 (N_20376,N_19852,N_18420);
and U20377 (N_20377,N_17985,N_19578);
nand U20378 (N_20378,N_19202,N_19893);
or U20379 (N_20379,N_19685,N_17910);
or U20380 (N_20380,N_18170,N_19921);
and U20381 (N_20381,N_17674,N_18136);
nor U20382 (N_20382,N_19413,N_18366);
nand U20383 (N_20383,N_18764,N_19343);
nand U20384 (N_20384,N_18992,N_18701);
nor U20385 (N_20385,N_18880,N_19553);
nand U20386 (N_20386,N_18747,N_18212);
nor U20387 (N_20387,N_19821,N_18394);
or U20388 (N_20388,N_17798,N_19923);
nor U20389 (N_20389,N_18211,N_17569);
nand U20390 (N_20390,N_19762,N_18319);
nand U20391 (N_20391,N_19414,N_19324);
nand U20392 (N_20392,N_19362,N_17947);
xnor U20393 (N_20393,N_17710,N_19541);
nand U20394 (N_20394,N_18452,N_17745);
and U20395 (N_20395,N_19212,N_19954);
or U20396 (N_20396,N_19449,N_17542);
or U20397 (N_20397,N_19391,N_19951);
xor U20398 (N_20398,N_19740,N_19653);
nand U20399 (N_20399,N_19916,N_18725);
nand U20400 (N_20400,N_18252,N_19428);
xor U20401 (N_20401,N_18703,N_18717);
and U20402 (N_20402,N_17625,N_18316);
nor U20403 (N_20403,N_18691,N_17606);
nor U20404 (N_20404,N_19700,N_17586);
and U20405 (N_20405,N_19930,N_18434);
and U20406 (N_20406,N_19684,N_18311);
nor U20407 (N_20407,N_17559,N_19364);
or U20408 (N_20408,N_19451,N_19059);
or U20409 (N_20409,N_19744,N_19229);
or U20410 (N_20410,N_17964,N_18832);
nand U20411 (N_20411,N_18287,N_18243);
and U20412 (N_20412,N_17653,N_17724);
or U20413 (N_20413,N_17636,N_17571);
nand U20414 (N_20414,N_18357,N_19177);
nand U20415 (N_20415,N_19666,N_19082);
nor U20416 (N_20416,N_19476,N_19529);
and U20417 (N_20417,N_18458,N_17770);
nor U20418 (N_20418,N_19392,N_19395);
nor U20419 (N_20419,N_19642,N_18642);
or U20420 (N_20420,N_19136,N_19040);
nor U20421 (N_20421,N_19114,N_18037);
and U20422 (N_20422,N_19784,N_18760);
or U20423 (N_20423,N_18296,N_19892);
and U20424 (N_20424,N_19444,N_18675);
nor U20425 (N_20425,N_19164,N_19387);
xor U20426 (N_20426,N_18964,N_19290);
nor U20427 (N_20427,N_18460,N_19066);
and U20428 (N_20428,N_17752,N_17949);
or U20429 (N_20429,N_18505,N_18550);
and U20430 (N_20430,N_18827,N_18030);
or U20431 (N_20431,N_18059,N_19036);
nand U20432 (N_20432,N_18963,N_19423);
or U20433 (N_20433,N_18369,N_19330);
nand U20434 (N_20434,N_17683,N_19630);
or U20435 (N_20435,N_17616,N_18811);
and U20436 (N_20436,N_19457,N_18684);
nor U20437 (N_20437,N_17644,N_19074);
nand U20438 (N_20438,N_18398,N_19329);
nor U20439 (N_20439,N_18973,N_19065);
or U20440 (N_20440,N_18423,N_18161);
nor U20441 (N_20441,N_19075,N_18743);
nand U20442 (N_20442,N_18934,N_17919);
or U20443 (N_20443,N_18205,N_19723);
and U20444 (N_20444,N_19947,N_17589);
nor U20445 (N_20445,N_19761,N_18303);
nand U20446 (N_20446,N_18203,N_18809);
nor U20447 (N_20447,N_17552,N_17951);
and U20448 (N_20448,N_19148,N_19739);
and U20449 (N_20449,N_17691,N_17727);
nand U20450 (N_20450,N_18567,N_18308);
nor U20451 (N_20451,N_18449,N_18448);
and U20452 (N_20452,N_19559,N_18947);
nor U20453 (N_20453,N_17516,N_17647);
nand U20454 (N_20454,N_19814,N_19184);
nor U20455 (N_20455,N_19794,N_18441);
nand U20456 (N_20456,N_18770,N_18371);
and U20457 (N_20457,N_18191,N_19445);
nor U20458 (N_20458,N_19815,N_19836);
nand U20459 (N_20459,N_19720,N_19936);
or U20460 (N_20460,N_18621,N_19707);
and U20461 (N_20461,N_17679,N_18808);
or U20462 (N_20462,N_17720,N_18395);
nor U20463 (N_20463,N_18727,N_18206);
nand U20464 (N_20464,N_18453,N_19881);
nand U20465 (N_20465,N_18549,N_19863);
or U20466 (N_20466,N_18662,N_18494);
nand U20467 (N_20467,N_19263,N_19850);
nor U20468 (N_20468,N_19396,N_18069);
nand U20469 (N_20469,N_17634,N_19468);
nor U20470 (N_20470,N_19754,N_19060);
xor U20471 (N_20471,N_19371,N_18834);
and U20472 (N_20472,N_19317,N_17723);
and U20473 (N_20473,N_17962,N_17527);
or U20474 (N_20474,N_17917,N_19403);
nand U20475 (N_20475,N_19546,N_17824);
and U20476 (N_20476,N_18515,N_19191);
or U20477 (N_20477,N_19671,N_18324);
nand U20478 (N_20478,N_18302,N_19419);
nor U20479 (N_20479,N_19446,N_17987);
nor U20480 (N_20480,N_19780,N_19605);
or U20481 (N_20481,N_19787,N_18902);
nand U20482 (N_20482,N_19268,N_19078);
and U20483 (N_20483,N_18024,N_18840);
nor U20484 (N_20484,N_18960,N_19424);
nor U20485 (N_20485,N_18443,N_19398);
xnor U20486 (N_20486,N_19549,N_18848);
and U20487 (N_20487,N_18864,N_17944);
or U20488 (N_20488,N_18338,N_19356);
nand U20489 (N_20489,N_18557,N_19016);
nor U20490 (N_20490,N_19966,N_17953);
and U20491 (N_20491,N_17832,N_19352);
or U20492 (N_20492,N_18264,N_18358);
nor U20493 (N_20493,N_19799,N_18092);
or U20494 (N_20494,N_19677,N_17614);
and U20495 (N_20495,N_17548,N_19463);
or U20496 (N_20496,N_17933,N_19781);
nor U20497 (N_20497,N_19974,N_18784);
and U20498 (N_20498,N_19128,N_17707);
or U20499 (N_20499,N_17854,N_18068);
and U20500 (N_20500,N_17900,N_17566);
and U20501 (N_20501,N_18224,N_17986);
and U20502 (N_20502,N_17983,N_19832);
nand U20503 (N_20503,N_18971,N_18083);
or U20504 (N_20504,N_18896,N_18817);
nor U20505 (N_20505,N_18966,N_19068);
nand U20506 (N_20506,N_18010,N_19021);
and U20507 (N_20507,N_19441,N_18791);
or U20508 (N_20508,N_19589,N_18917);
nor U20509 (N_20509,N_18925,N_18524);
and U20510 (N_20510,N_19411,N_19193);
or U20511 (N_20511,N_18271,N_17974);
or U20512 (N_20512,N_19110,N_19602);
nor U20513 (N_20513,N_17980,N_17565);
nor U20514 (N_20514,N_19601,N_19935);
or U20515 (N_20515,N_18983,N_19547);
and U20516 (N_20516,N_18255,N_18321);
or U20517 (N_20517,N_18984,N_19001);
or U20518 (N_20518,N_19327,N_18410);
or U20519 (N_20519,N_18053,N_19975);
or U20520 (N_20520,N_17624,N_18670);
and U20521 (N_20521,N_18525,N_18793);
nand U20522 (N_20522,N_17893,N_17930);
nor U20523 (N_20523,N_17828,N_19535);
nor U20524 (N_20524,N_17831,N_18306);
nand U20525 (N_20525,N_19450,N_18680);
nor U20526 (N_20526,N_17623,N_18645);
nand U20527 (N_20527,N_19929,N_19626);
and U20528 (N_20528,N_18821,N_17880);
or U20529 (N_20529,N_19295,N_19636);
and U20530 (N_20530,N_19885,N_17734);
nand U20531 (N_20531,N_19196,N_18698);
nand U20532 (N_20532,N_17777,N_19401);
nand U20533 (N_20533,N_18699,N_19980);
nand U20534 (N_20534,N_18365,N_19240);
nand U20535 (N_20535,N_18776,N_17881);
or U20536 (N_20536,N_17627,N_19294);
or U20537 (N_20537,N_19404,N_17897);
and U20538 (N_20538,N_18209,N_18559);
nand U20539 (N_20539,N_19305,N_17789);
or U20540 (N_20540,N_18142,N_18841);
nand U20541 (N_20541,N_17575,N_17792);
or U20542 (N_20542,N_19276,N_18079);
nand U20543 (N_20543,N_18736,N_18329);
nand U20544 (N_20544,N_18785,N_17588);
nand U20545 (N_20545,N_17782,N_18425);
nor U20546 (N_20546,N_19090,N_19763);
and U20547 (N_20547,N_17906,N_18801);
nor U20548 (N_20548,N_18539,N_19109);
and U20549 (N_20549,N_19248,N_19030);
and U20550 (N_20550,N_19698,N_17747);
nand U20551 (N_20551,N_19009,N_19415);
nand U20552 (N_20552,N_19153,N_18115);
and U20553 (N_20553,N_19353,N_19499);
or U20554 (N_20554,N_17954,N_18753);
and U20555 (N_20555,N_19484,N_18954);
or U20556 (N_20556,N_18989,N_17655);
and U20557 (N_20557,N_18478,N_18427);
nand U20558 (N_20558,N_18886,N_19801);
and U20559 (N_20559,N_17939,N_17915);
and U20560 (N_20560,N_19517,N_17977);
or U20561 (N_20561,N_18233,N_18232);
or U20562 (N_20562,N_18415,N_19373);
or U20563 (N_20563,N_19321,N_17615);
nor U20564 (N_20564,N_18002,N_18889);
and U20565 (N_20565,N_17909,N_17709);
nand U20566 (N_20566,N_17808,N_17730);
nand U20567 (N_20567,N_19768,N_18568);
and U20568 (N_20568,N_18668,N_19050);
nor U20569 (N_20569,N_19338,N_19501);
and U20570 (N_20570,N_19017,N_19627);
or U20571 (N_20571,N_18728,N_19681);
or U20572 (N_20572,N_18799,N_17682);
nand U20573 (N_20573,N_19325,N_19176);
or U20574 (N_20574,N_17685,N_19355);
or U20575 (N_20575,N_19368,N_18502);
nor U20576 (N_20576,N_19746,N_18522);
or U20577 (N_20577,N_17650,N_19572);
nand U20578 (N_20578,N_17684,N_19489);
or U20579 (N_20579,N_17837,N_17768);
nand U20580 (N_20580,N_18006,N_19224);
or U20581 (N_20581,N_19598,N_18377);
or U20582 (N_20582,N_17574,N_19606);
nand U20583 (N_20583,N_18225,N_19725);
or U20584 (N_20584,N_18595,N_18475);
and U20585 (N_20585,N_18956,N_19151);
or U20586 (N_20586,N_19910,N_18871);
or U20587 (N_20587,N_19046,N_19442);
nor U20588 (N_20588,N_19905,N_18573);
nand U20589 (N_20589,N_19767,N_17660);
and U20590 (N_20590,N_18470,N_18285);
or U20591 (N_20591,N_17719,N_19867);
nor U20592 (N_20592,N_18570,N_18386);
and U20593 (N_20593,N_18771,N_19569);
nor U20594 (N_20594,N_18553,N_18348);
nor U20595 (N_20595,N_19032,N_18001);
and U20596 (N_20596,N_19375,N_19247);
nand U20597 (N_20597,N_18766,N_19597);
or U20598 (N_20598,N_17843,N_18571);
nand U20599 (N_20599,N_18288,N_19094);
or U20600 (N_20600,N_19519,N_19532);
nand U20601 (N_20601,N_19841,N_19510);
or U20602 (N_20602,N_18354,N_19858);
and U20603 (N_20603,N_18457,N_19741);
or U20604 (N_20604,N_19895,N_18235);
nor U20605 (N_20605,N_17523,N_19550);
or U20606 (N_20606,N_18938,N_18124);
and U20607 (N_20607,N_18293,N_18755);
nand U20608 (N_20608,N_18936,N_19154);
nor U20609 (N_20609,N_19113,N_18178);
or U20610 (N_20610,N_18155,N_17677);
nor U20611 (N_20611,N_19724,N_17689);
nand U20612 (N_20612,N_18843,N_18825);
or U20613 (N_20613,N_19429,N_19272);
or U20614 (N_20614,N_19943,N_19967);
nor U20615 (N_20615,N_18281,N_19171);
or U20616 (N_20616,N_19939,N_17567);
or U20617 (N_20617,N_18474,N_19566);
or U20618 (N_20618,N_18492,N_17847);
nand U20619 (N_20619,N_19982,N_17812);
or U20620 (N_20620,N_19871,N_17927);
or U20621 (N_20621,N_18972,N_18556);
or U20622 (N_20622,N_17602,N_18831);
nor U20623 (N_20623,N_18101,N_19431);
nor U20624 (N_20624,N_18688,N_18815);
xor U20625 (N_20625,N_17587,N_18796);
nand U20626 (N_20626,N_19971,N_18594);
or U20627 (N_20627,N_18721,N_19104);
nor U20628 (N_20628,N_18563,N_19765);
and U20629 (N_20629,N_18223,N_19393);
nor U20630 (N_20630,N_19173,N_17676);
nor U20631 (N_20631,N_19708,N_17553);
nor U20632 (N_20632,N_19211,N_19663);
xnor U20633 (N_20633,N_19709,N_19436);
nor U20634 (N_20634,N_19513,N_18781);
or U20635 (N_20635,N_19129,N_19710);
nor U20636 (N_20636,N_19486,N_18135);
or U20637 (N_20637,N_18707,N_19235);
and U20638 (N_20638,N_17876,N_19258);
nor U20639 (N_20639,N_19528,N_18849);
or U20640 (N_20640,N_17643,N_18257);
nor U20641 (N_20641,N_18928,N_19593);
nand U20642 (N_20642,N_18591,N_17993);
nor U20643 (N_20643,N_18270,N_19227);
nor U20644 (N_20644,N_18533,N_18585);
nor U20645 (N_20645,N_18200,N_18657);
or U20646 (N_20646,N_19043,N_17884);
or U20647 (N_20647,N_19674,N_17989);
and U20648 (N_20648,N_19525,N_18912);
or U20649 (N_20649,N_19332,N_19727);
and U20650 (N_20650,N_18171,N_19464);
or U20651 (N_20651,N_17649,N_19882);
nor U20652 (N_20652,N_17803,N_18469);
and U20653 (N_20653,N_18265,N_18933);
nor U20654 (N_20654,N_17963,N_17862);
nor U20655 (N_20655,N_19498,N_17728);
nor U20656 (N_20656,N_17576,N_17821);
nor U20657 (N_20657,N_19804,N_18163);
and U20658 (N_20658,N_18899,N_18501);
and U20659 (N_20659,N_18790,N_19269);
or U20660 (N_20660,N_18484,N_19639);
nand U20661 (N_20661,N_18669,N_19977);
xor U20662 (N_20662,N_18100,N_19618);
and U20663 (N_20663,N_18123,N_18833);
nor U20664 (N_20664,N_18418,N_19968);
nor U20665 (N_20665,N_17835,N_17878);
or U20666 (N_20666,N_19102,N_19112);
nor U20667 (N_20667,N_19408,N_17942);
and U20668 (N_20668,N_18112,N_18183);
nand U20669 (N_20669,N_17889,N_18761);
nor U20670 (N_20670,N_19973,N_17590);
nand U20671 (N_20671,N_17713,N_17716);
and U20672 (N_20672,N_18162,N_19664);
and U20673 (N_20673,N_17692,N_17815);
or U20674 (N_20674,N_17904,N_17899);
and U20675 (N_20675,N_17766,N_18888);
nor U20676 (N_20676,N_17503,N_19629);
nor U20677 (N_20677,N_19076,N_19878);
nor U20678 (N_20678,N_18967,N_19035);
nand U20679 (N_20679,N_17744,N_17908);
nor U20680 (N_20680,N_19691,N_18847);
nand U20681 (N_20681,N_18299,N_19253);
nor U20682 (N_20682,N_18959,N_19287);
nor U20683 (N_20683,N_19806,N_18023);
nor U20684 (N_20684,N_19452,N_17666);
nor U20685 (N_20685,N_17537,N_19336);
and U20686 (N_20686,N_18438,N_19152);
nand U20687 (N_20687,N_19701,N_18199);
nor U20688 (N_20688,N_17721,N_17845);
and U20689 (N_20689,N_18246,N_18682);
nand U20690 (N_20690,N_19827,N_19071);
and U20691 (N_20691,N_19978,N_19735);
and U20692 (N_20692,N_19831,N_19989);
nor U20693 (N_20693,N_18751,N_19686);
and U20694 (N_20694,N_19564,N_19990);
nor U20695 (N_20695,N_17711,N_18695);
and U20696 (N_20696,N_19837,N_17793);
and U20697 (N_20697,N_19716,N_18686);
and U20698 (N_20698,N_18088,N_18548);
or U20699 (N_20699,N_17604,N_17905);
and U20700 (N_20700,N_18741,N_19284);
nand U20701 (N_20701,N_18231,N_17848);
nor U20702 (N_20702,N_17769,N_19957);
nand U20703 (N_20703,N_17978,N_18908);
or U20704 (N_20704,N_19222,N_18393);
nand U20705 (N_20705,N_18655,N_19054);
nor U20706 (N_20706,N_19251,N_19798);
nand U20707 (N_20707,N_17543,N_19625);
nand U20708 (N_20708,N_18618,N_17820);
nor U20709 (N_20709,N_19760,N_18589);
nor U20710 (N_20710,N_19683,N_18011);
or U20711 (N_20711,N_18957,N_19274);
and U20712 (N_20712,N_17519,N_19747);
nor U20713 (N_20713,N_17888,N_19582);
and U20714 (N_20714,N_19813,N_19091);
or U20715 (N_20715,N_18512,N_19047);
nor U20716 (N_20716,N_18054,N_19748);
or U20717 (N_20717,N_18683,N_18745);
or U20718 (N_20718,N_17539,N_17695);
nand U20719 (N_20719,N_17864,N_18582);
nor U20720 (N_20720,N_18208,N_17858);
or U20721 (N_20721,N_18726,N_19361);
nor U20722 (N_20722,N_19228,N_19552);
and U20723 (N_20723,N_17582,N_18856);
and U20724 (N_20724,N_18511,N_19770);
and U20725 (N_20725,N_19659,N_17694);
nor U20726 (N_20726,N_17669,N_18489);
nand U20727 (N_20727,N_19588,N_18071);
nor U20728 (N_20728,N_19166,N_18653);
nor U20729 (N_20729,N_18646,N_19654);
nor U20730 (N_20730,N_17957,N_19633);
nor U20731 (N_20731,N_19427,N_18541);
nor U20732 (N_20732,N_19766,N_19676);
nor U20733 (N_20733,N_18696,N_19646);
and U20734 (N_20734,N_17513,N_18005);
nand U20735 (N_20735,N_19143,N_19998);
nand U20736 (N_20736,N_18295,N_18632);
nor U20737 (N_20737,N_19734,N_18845);
nand U20738 (N_20738,N_19577,N_19793);
nor U20739 (N_20739,N_18693,N_18102);
nand U20740 (N_20740,N_19479,N_18968);
or U20741 (N_20741,N_17506,N_19096);
and U20742 (N_20742,N_19834,N_19254);
nand U20743 (N_20743,N_19127,N_19354);
nand U20744 (N_20744,N_17819,N_18251);
and U20745 (N_20745,N_18440,N_18040);
nor U20746 (N_20746,N_17809,N_19041);
and U20747 (N_20747,N_19377,N_19231);
nand U20748 (N_20748,N_18349,N_17733);
and U20749 (N_20749,N_19052,N_18861);
nand U20750 (N_20750,N_18343,N_17551);
nand U20751 (N_20751,N_19718,N_18866);
or U20752 (N_20752,N_17667,N_18577);
nor U20753 (N_20753,N_18483,N_18008);
and U20754 (N_20754,N_19619,N_18506);
nand U20755 (N_20755,N_18099,N_19849);
nor U20756 (N_20756,N_19840,N_17585);
and U20757 (N_20757,N_17563,N_17976);
nand U20758 (N_20758,N_19568,N_19379);
nor U20759 (N_20759,N_17991,N_19826);
nand U20760 (N_20760,N_19080,N_18997);
nor U20761 (N_20761,N_17754,N_19482);
or U20762 (N_20762,N_19264,N_19786);
and U20763 (N_20763,N_19574,N_19575);
or U20764 (N_20764,N_17594,N_18576);
or U20765 (N_20765,N_18844,N_18802);
and U20766 (N_20766,N_17620,N_17773);
nor U20767 (N_20767,N_18730,N_19521);
or U20768 (N_20768,N_18363,N_19372);
nand U20769 (N_20769,N_19246,N_17883);
and U20770 (N_20770,N_18648,N_18131);
or U20771 (N_20771,N_19366,N_18952);
nand U20772 (N_20772,N_19048,N_19632);
nor U20773 (N_20773,N_17950,N_19015);
nor U20774 (N_20774,N_17918,N_19456);
nor U20775 (N_20775,N_18043,N_18258);
nor U20776 (N_20776,N_18651,N_17583);
nand U20777 (N_20777,N_19194,N_18588);
nor U20778 (N_20778,N_18327,N_19344);
nand U20779 (N_20779,N_18565,N_18836);
or U20780 (N_20780,N_19667,N_18259);
nand U20781 (N_20781,N_17671,N_17621);
nand U20782 (N_20782,N_18596,N_18222);
nand U20783 (N_20783,N_19245,N_18800);
or U20784 (N_20784,N_17802,N_18854);
and U20785 (N_20785,N_19011,N_19055);
nand U20786 (N_20786,N_19859,N_18535);
nand U20787 (N_20787,N_17712,N_18180);
and U20788 (N_20788,N_17931,N_17852);
nand U20789 (N_20789,N_17929,N_18075);
and U20790 (N_20790,N_17952,N_18226);
and U20791 (N_20791,N_18150,N_19884);
nand U20792 (N_20792,N_19759,N_18544);
or U20793 (N_20793,N_19694,N_19702);
nand U20794 (N_20794,N_17737,N_17630);
or U20795 (N_20795,N_19189,N_18117);
and U20796 (N_20796,N_19485,N_17540);
and U20797 (N_20797,N_18168,N_19610);
nor U20798 (N_20798,N_19675,N_19407);
nor U20799 (N_20799,N_17645,N_19942);
nor U20800 (N_20800,N_18850,N_19186);
or U20801 (N_20801,N_19491,N_18237);
nor U20802 (N_20802,N_18156,N_18752);
nor U20803 (N_20803,N_19679,N_18528);
or U20804 (N_20804,N_17508,N_17697);
nor U20805 (N_20805,N_18787,N_18746);
nand U20806 (N_20806,N_17816,N_18373);
nor U20807 (N_20807,N_18562,N_18611);
and U20808 (N_20808,N_18712,N_18076);
nand U20809 (N_20809,N_17759,N_17651);
or U20810 (N_20810,N_18405,N_19019);
nor U20811 (N_20811,N_18976,N_18388);
nor U20812 (N_20812,N_18587,N_19961);
or U20813 (N_20813,N_17781,N_18937);
nor U20814 (N_20814,N_19538,N_18172);
nor U20815 (N_20815,N_18248,N_19044);
and U20816 (N_20816,N_18788,N_19823);
nor U20817 (N_20817,N_19281,N_19771);
xor U20818 (N_20818,N_17868,N_18777);
nand U20819 (N_20819,N_19421,N_18521);
nand U20820 (N_20820,N_19137,N_19996);
nand U20821 (N_20821,N_19282,N_18750);
nand U20822 (N_20822,N_19825,N_17946);
or U20823 (N_20823,N_18718,N_17896);
nor U20824 (N_20824,N_19465,N_17764);
or U20825 (N_20825,N_19380,N_17619);
or U20826 (N_20826,N_19296,N_19855);
and U20827 (N_20827,N_19869,N_18298);
nor U20828 (N_20828,N_19623,N_17948);
and U20829 (N_20829,N_19773,N_18164);
and U20830 (N_20830,N_18716,N_19726);
and U20831 (N_20831,N_19376,N_17765);
or U20832 (N_20832,N_18151,N_18507);
nand U20833 (N_20833,N_18710,N_18977);
nor U20834 (N_20834,N_18926,N_19544);
nand U20835 (N_20835,N_18993,N_17529);
nand U20836 (N_20836,N_17813,N_17995);
and U20837 (N_20837,N_18175,N_18869);
nand U20838 (N_20838,N_18353,N_17732);
or U20839 (N_20839,N_19638,N_19225);
nor U20840 (N_20840,N_17901,N_18051);
or U20841 (N_20841,N_19312,N_18536);
or U20842 (N_20842,N_18026,N_19042);
nor U20843 (N_20843,N_19820,N_19239);
or U20844 (N_20844,N_17776,N_18368);
nor U20845 (N_20845,N_17869,N_17584);
or U20846 (N_20846,N_19631,N_19168);
or U20847 (N_20847,N_17579,N_17788);
and U20848 (N_20848,N_17870,N_18390);
nand U20849 (N_20849,N_19828,N_17779);
or U20850 (N_20850,N_19323,N_19969);
or U20851 (N_20851,N_18660,N_18279);
or U20852 (N_20852,N_19242,N_19777);
nand U20853 (N_20853,N_19908,N_17753);
nand U20854 (N_20854,N_19033,N_19031);
nor U20855 (N_20855,N_19648,N_18892);
nand U20856 (N_20856,N_19117,N_17829);
and U20857 (N_20857,N_18643,N_18921);
nor U20858 (N_20858,N_19703,N_18333);
nor U20859 (N_20859,N_19218,N_18229);
nor U20860 (N_20860,N_18486,N_18647);
nand U20861 (N_20861,N_18704,N_17664);
nand U20862 (N_20862,N_19838,N_17743);
nand U20863 (N_20863,N_19914,N_18945);
or U20864 (N_20864,N_19651,N_19596);
and U20865 (N_20865,N_18340,N_17670);
and U20866 (N_20866,N_17696,N_19874);
or U20867 (N_20867,N_18941,N_17500);
nor U20868 (N_20868,N_19237,N_19576);
or U20869 (N_20869,N_19586,N_19430);
nor U20870 (N_20870,N_17926,N_18919);
or U20871 (N_20871,N_17706,N_18119);
nor U20872 (N_20872,N_19570,N_18318);
or U20873 (N_20873,N_18855,N_18107);
or U20874 (N_20874,N_18261,N_19733);
and U20875 (N_20875,N_18715,N_19846);
nand U20876 (N_20876,N_19868,N_18980);
nand U20877 (N_20877,N_19560,N_18019);
nand U20878 (N_20878,N_17693,N_17700);
or U20879 (N_20879,N_17635,N_18628);
or U20880 (N_20880,N_19628,N_19103);
nand U20881 (N_20881,N_17546,N_19983);
and U20882 (N_20882,N_19944,N_18722);
or U20883 (N_20883,N_17938,N_18759);
or U20884 (N_20884,N_19337,N_17762);
and U20885 (N_20885,N_17903,N_18810);
nand U20886 (N_20886,N_18450,N_19650);
or U20887 (N_20887,N_19875,N_17959);
and U20888 (N_20888,N_19573,N_19609);
and U20889 (N_20889,N_19495,N_18276);
or U20890 (N_20890,N_18561,N_17714);
and U20891 (N_20891,N_19647,N_17784);
or U20892 (N_20892,N_19255,N_17856);
nor U20893 (N_20893,N_18416,N_17867);
or U20894 (N_20894,N_17626,N_18950);
nor U20895 (N_20895,N_19161,N_19590);
and U20896 (N_20896,N_17518,N_17628);
or U20897 (N_20897,N_19233,N_18630);
nand U20898 (N_20898,N_18685,N_19147);
nor U20899 (N_20899,N_18403,N_18093);
nand U20900 (N_20900,N_19162,N_19333);
nor U20901 (N_20901,N_17573,N_17787);
and U20902 (N_20902,N_19891,N_19556);
nor U20903 (N_20903,N_17600,N_17810);
or U20904 (N_20904,N_17681,N_17740);
nand U20905 (N_20905,N_18658,N_19913);
nand U20906 (N_20906,N_17827,N_19120);
xnor U20907 (N_20907,N_19811,N_19689);
or U20908 (N_20908,N_17517,N_18814);
or U20909 (N_20909,N_18823,N_18375);
and U20910 (N_20910,N_18004,N_19712);
or U20911 (N_20911,N_19447,N_17839);
nand U20912 (N_20912,N_19774,N_17886);
nor U20913 (N_20913,N_18077,N_17800);
and U20914 (N_20914,N_19607,N_17642);
nand U20915 (N_20915,N_18370,N_19796);
nand U20916 (N_20916,N_19494,N_17672);
and U20917 (N_20917,N_18617,N_19210);
nand U20918 (N_20918,N_19644,N_17814);
or U20919 (N_20919,N_17841,N_18074);
and U20920 (N_20920,N_18372,N_18188);
nor U20921 (N_20921,N_19673,N_19879);
nand U20922 (N_20922,N_18114,N_19862);
and U20923 (N_20923,N_18080,N_19458);
nor U20924 (N_20924,N_19024,N_19512);
or U20925 (N_20925,N_18898,N_17755);
or U20926 (N_20926,N_18204,N_19382);
or U20927 (N_20927,N_19331,N_18219);
nor U20928 (N_20928,N_18000,N_18636);
nor U20929 (N_20929,N_18890,N_17761);
nand U20930 (N_20930,N_19918,N_19864);
nor U20931 (N_20931,N_17698,N_19920);
and U20932 (N_20932,N_17562,N_19719);
and U20933 (N_20933,N_18341,N_19956);
nor U20934 (N_20934,N_18795,N_18018);
and U20935 (N_20935,N_18775,N_17631);
or U20936 (N_20936,N_18891,N_17525);
and U20937 (N_20937,N_18214,N_19062);
nand U20938 (N_20938,N_19002,N_19995);
xnor U20939 (N_20939,N_17850,N_19769);
nand U20940 (N_20940,N_18819,N_19561);
nor U20941 (N_20941,N_19518,N_19902);
nor U20942 (N_20942,N_18860,N_18294);
nor U20943 (N_20943,N_17796,N_19238);
or U20944 (N_20944,N_19367,N_17750);
nand U20945 (N_20945,N_17756,N_19488);
or U20946 (N_20946,N_17790,N_17785);
nand U20947 (N_20947,N_19115,N_19079);
nor U20948 (N_20948,N_19388,N_18072);
nand U20949 (N_20949,N_19497,N_19394);
nor U20950 (N_20950,N_19941,N_19581);
and U20951 (N_20951,N_19405,N_18408);
nor U20952 (N_20952,N_17598,N_18608);
or U20953 (N_20953,N_18091,N_18210);
nor U20954 (N_20954,N_18384,N_18578);
nor U20955 (N_20955,N_19987,N_19014);
xor U20956 (N_20956,N_19010,N_18552);
nand U20957 (N_20957,N_18181,N_18466);
nor U20958 (N_20958,N_19737,N_18242);
nor U20959 (N_20959,N_18064,N_19932);
nor U20960 (N_20960,N_18797,N_18953);
or U20961 (N_20961,N_19234,N_19386);
and U20962 (N_20962,N_18422,N_18737);
nand U20963 (N_20963,N_18913,N_18714);
or U20964 (N_20964,N_19125,N_17817);
and U20965 (N_20965,N_19889,N_19924);
or U20966 (N_20966,N_18583,N_18998);
and U20967 (N_20967,N_18309,N_18182);
nand U20968 (N_20968,N_19717,N_17572);
or U20969 (N_20969,N_18090,N_18895);
or U20970 (N_20970,N_18391,N_19390);
nor U20971 (N_20971,N_17805,N_19715);
or U20972 (N_20972,N_19805,N_19265);
or U20973 (N_20973,N_18846,N_19682);
or U20974 (N_20974,N_17648,N_17520);
or U20975 (N_20975,N_17833,N_18592);
nor U20976 (N_20976,N_19462,N_18050);
and U20977 (N_20977,N_19397,N_18186);
nand U20978 (N_20978,N_18332,N_17545);
nand U20979 (N_20979,N_19502,N_18915);
nor U20980 (N_20980,N_18244,N_19992);
and U20981 (N_20981,N_17637,N_18157);
nand U20982 (N_20982,N_19634,N_19241);
or U20983 (N_20983,N_18910,N_18767);
or U20984 (N_20984,N_18414,N_18129);
nand U20985 (N_20985,N_18256,N_18052);
and U20986 (N_20986,N_18564,N_18805);
and U20987 (N_20987,N_19539,N_17524);
and U20988 (N_20988,N_19548,N_18480);
nor U20989 (N_20989,N_19795,N_18409);
nand U20990 (N_20990,N_18144,N_17597);
nor U20991 (N_20991,N_18678,N_18445);
or U20992 (N_20992,N_18228,N_19306);
or U20993 (N_20993,N_19200,N_17804);
nand U20994 (N_20994,N_18870,N_18277);
and U20995 (N_20995,N_18029,N_18590);
or U20996 (N_20996,N_19822,N_17791);
nor U20997 (N_20997,N_18593,N_18526);
or U20998 (N_20998,N_19555,N_17885);
nor U20999 (N_20999,N_19435,N_19400);
or U21000 (N_21000,N_19964,N_18192);
xor U21001 (N_21001,N_18904,N_17955);
nor U21002 (N_21002,N_17678,N_19645);
and U21003 (N_21003,N_18477,N_18359);
nand U21004 (N_21004,N_18297,N_18554);
and U21005 (N_21005,N_19500,N_18763);
nor U21006 (N_21006,N_19571,N_18720);
and U21007 (N_21007,N_18300,N_17715);
or U21008 (N_21008,N_18061,N_19562);
or U21009 (N_21009,N_19384,N_19142);
and U21010 (N_21010,N_19360,N_18988);
nand U21011 (N_21011,N_17725,N_17511);
or U21012 (N_21012,N_19460,N_18201);
nand U21013 (N_21013,N_17515,N_19807);
nor U21014 (N_21014,N_19764,N_18304);
and U21015 (N_21015,N_17840,N_19000);
nand U21016 (N_21016,N_17825,N_18885);
or U21017 (N_21017,N_19448,N_19730);
and U21018 (N_21018,N_17892,N_18013);
and U21019 (N_21019,N_19672,N_18060);
or U21020 (N_21020,N_19621,N_18881);
nor U21021 (N_21021,N_18207,N_18924);
xor U21022 (N_21022,N_19319,N_18702);
nand U21023 (N_21023,N_18674,N_19865);
nor U21024 (N_21024,N_19857,N_18758);
or U21025 (N_21025,N_18816,N_17973);
or U21026 (N_21026,N_19466,N_19220);
or U21027 (N_21027,N_18664,N_18542);
nand U21028 (N_21028,N_17509,N_19516);
nor U21029 (N_21029,N_19934,N_18097);
nor U21030 (N_21030,N_17717,N_19604);
nor U21031 (N_21031,N_18350,N_19409);
or U21032 (N_21032,N_19808,N_18987);
nor U21033 (N_21033,N_19472,N_17965);
and U21034 (N_21034,N_19278,N_18822);
or U21035 (N_21035,N_18883,N_17891);
or U21036 (N_21036,N_19064,N_18284);
or U21037 (N_21037,N_19067,N_19188);
and U21038 (N_21038,N_18260,N_19454);
nor U21039 (N_21039,N_19433,N_17577);
or U21040 (N_21040,N_18868,N_19318);
or U21041 (N_21041,N_18982,N_18994);
nand U21042 (N_21042,N_17866,N_19979);
or U21043 (N_21043,N_18160,N_19856);
nor U21044 (N_21044,N_19915,N_18804);
nand U21045 (N_21045,N_19195,N_19169);
and U21046 (N_21046,N_19123,N_17818);
nor U21047 (N_21047,N_19157,N_18604);
nand U21048 (N_21048,N_19199,N_19728);
or U21049 (N_21049,N_17530,N_18346);
nor U21050 (N_21050,N_18429,N_19144);
nor U21051 (N_21051,N_17580,N_18824);
nand U21052 (N_21052,N_17512,N_18413);
and U21053 (N_21053,N_19302,N_19130);
nor U21054 (N_21054,N_18754,N_18842);
or U21055 (N_21055,N_18514,N_18547);
nand U21056 (N_21056,N_17633,N_19809);
xor U21057 (N_21057,N_19854,N_19940);
or U21058 (N_21058,N_17618,N_18620);
or U21059 (N_21059,N_19098,N_19389);
and U21060 (N_21060,N_18711,N_18463);
and U21061 (N_21061,N_19340,N_18872);
nand U21062 (N_21062,N_17967,N_18103);
nor U21063 (N_21063,N_19097,N_18826);
and U21064 (N_21064,N_18499,N_18317);
nor U21065 (N_21065,N_18607,N_18109);
or U21066 (N_21066,N_19049,N_19652);
or U21067 (N_21067,N_18017,N_19999);
or U21068 (N_21068,N_17544,N_19662);
and U21069 (N_21069,N_19190,N_19467);
nor U21070 (N_21070,N_17718,N_18656);
and U21071 (N_21071,N_17735,N_18677);
and U21072 (N_21072,N_19159,N_19267);
nand U21073 (N_21073,N_18619,N_19061);
nand U21074 (N_21074,N_17992,N_17872);
nor U21075 (N_21075,N_18108,N_17554);
nor U21076 (N_21076,N_18272,N_18519);
or U21077 (N_21077,N_18042,N_19399);
nand U21078 (N_21078,N_18266,N_18569);
nand U21079 (N_21079,N_18708,N_18138);
nor U21080 (N_21080,N_19976,N_18852);
nor U21081 (N_21081,N_19901,N_17994);
nand U21082 (N_21082,N_17934,N_18652);
or U21083 (N_21083,N_19583,N_18631);
and U21084 (N_21084,N_19121,N_19089);
nor U21085 (N_21085,N_18383,N_18442);
or U21086 (N_21086,N_19745,N_17578);
nor U21087 (N_21087,N_18290,N_19481);
or U21088 (N_21088,N_18667,N_18122);
and U21089 (N_21089,N_19812,N_18638);
or U21090 (N_21090,N_19086,N_19057);
nor U21091 (N_21091,N_19960,N_19146);
and U21092 (N_21092,N_18687,N_19751);
nand U21093 (N_21093,N_18057,N_19283);
nand U21094 (N_21094,N_18935,N_19743);
nand U21095 (N_21095,N_18922,N_19383);
or U21096 (N_21096,N_19084,N_18465);
nor U21097 (N_21097,N_19135,N_18347);
nor U21098 (N_21098,N_19697,N_18780);
and U21099 (N_21099,N_18900,N_19088);
and U21100 (N_21100,N_17838,N_19478);
nand U21101 (N_21101,N_19953,N_19007);
nand U21102 (N_21102,N_17739,N_19818);
or U21103 (N_21103,N_17581,N_19223);
and U21104 (N_21104,N_19412,N_19180);
nor U21105 (N_21105,N_18254,N_18942);
nand U21106 (N_21106,N_19861,N_18387);
or U21107 (N_21107,N_19649,N_19695);
and U21108 (N_21108,N_19275,N_18095);
nor U21109 (N_21109,N_19661,N_19012);
or U21110 (N_21110,N_19981,N_19870);
nor U21111 (N_21111,N_18639,N_17751);
and U21112 (N_21112,N_18627,N_18194);
nor U21113 (N_21113,N_19280,N_19471);
nand U21114 (N_21114,N_18859,N_17834);
nor U21115 (N_21115,N_17921,N_19203);
and U21116 (N_21116,N_18624,N_18356);
nor U21117 (N_21117,N_18981,N_17984);
and U21118 (N_21118,N_18857,N_17659);
nor U21119 (N_21119,N_17617,N_17970);
nand U21120 (N_21120,N_18774,N_19132);
or U21121 (N_21121,N_18305,N_18723);
nor U21122 (N_21122,N_19256,N_19350);
and U21123 (N_21123,N_18508,N_19335);
or U21124 (N_21124,N_17898,N_19134);
and U21125 (N_21125,N_18374,N_18615);
or U21126 (N_21126,N_17704,N_19931);
and U21127 (N_21127,N_18979,N_19197);
nand U21128 (N_21128,N_17612,N_19789);
nand U21129 (N_21129,N_17601,N_19299);
nand U21130 (N_21130,N_19357,N_18517);
and U21131 (N_21131,N_18943,N_18672);
and U21132 (N_21132,N_17534,N_17558);
and U21133 (N_21133,N_19595,N_19027);
nor U21134 (N_21134,N_18634,N_18143);
nor U21135 (N_21135,N_18012,N_17673);
or U21136 (N_21136,N_19926,N_19116);
and U21137 (N_21137,N_19262,N_17797);
nand U21138 (N_21138,N_18044,N_19138);
or U21139 (N_21139,N_19221,N_19790);
or U21140 (N_21140,N_19958,N_19520);
and U21141 (N_21141,N_19903,N_18914);
nor U21142 (N_21142,N_18086,N_18096);
nand U21143 (N_21143,N_18732,N_18529);
xor U21144 (N_21144,N_18700,N_18193);
nand U21145 (N_21145,N_18351,N_18411);
nor U21146 (N_21146,N_18230,N_18187);
and U21147 (N_21147,N_19670,N_19140);
and U21148 (N_21148,N_19341,N_18485);
nor U21149 (N_21149,N_19515,N_18038);
or U21150 (N_21150,N_17774,N_18021);
nor U21151 (N_21151,N_18903,N_19297);
xor U21152 (N_21152,N_17932,N_17533);
and U21153 (N_21153,N_18940,N_19118);
and U21154 (N_21154,N_18706,N_19385);
and U21155 (N_21155,N_19099,N_19038);
nor U21156 (N_21156,N_18705,N_19531);
nor U21157 (N_21157,N_18020,N_18713);
or U21158 (N_21158,N_17640,N_19580);
nand U21159 (N_21159,N_19020,N_19298);
nand U21160 (N_21160,N_19758,N_19455);
and U21161 (N_21161,N_18540,N_19230);
nand U21162 (N_21162,N_18459,N_18399);
nand U21163 (N_21163,N_19170,N_18015);
nand U21164 (N_21164,N_19496,N_19540);
or U21165 (N_21165,N_18537,N_18345);
and U21166 (N_21166,N_18307,N_18659);
or U21167 (N_21167,N_19492,N_19504);
nand U21168 (N_21168,N_18245,N_19585);
or U21169 (N_21169,N_18336,N_18930);
nor U21170 (N_21170,N_18247,N_19533);
or U21171 (N_21171,N_19876,N_17680);
nand U21172 (N_21172,N_18159,N_18551);
nand U21173 (N_21173,N_18689,N_19775);
or U21174 (N_21174,N_18047,N_17686);
nand U21175 (N_21175,N_19536,N_18782);
or U21176 (N_21176,N_19359,N_17911);
or U21177 (N_21177,N_17526,N_17622);
or U21178 (N_21178,N_18969,N_19792);
or U21179 (N_21179,N_18334,N_18401);
nor U21180 (N_21180,N_18991,N_19025);
or U21181 (N_21181,N_17873,N_17591);
or U21182 (N_21182,N_19984,N_19877);
nand U21183 (N_21183,N_19004,N_19962);
nand U21184 (N_21184,N_17629,N_17767);
xnor U21185 (N_21185,N_18586,N_18773);
xnor U21186 (N_21186,N_17556,N_19890);
nor U21187 (N_21187,N_18428,N_19183);
nand U21188 (N_21188,N_18920,N_17806);
or U21189 (N_21189,N_18476,N_17849);
and U21190 (N_21190,N_19909,N_17564);
and U21191 (N_21191,N_17599,N_19026);
and U21192 (N_21192,N_18062,N_19731);
or U21193 (N_21193,N_19551,N_19545);
nand U21194 (N_21194,N_19656,N_19620);
and U21195 (N_21195,N_18609,N_18650);
and U21196 (N_21196,N_19558,N_19959);
or U21197 (N_21197,N_19363,N_17894);
nand U21198 (N_21198,N_19439,N_18812);
nand U21199 (N_21199,N_19163,N_19314);
nand U21200 (N_21200,N_17547,N_18493);
nor U21201 (N_21201,N_19018,N_18671);
nand U21202 (N_21202,N_18749,N_18313);
or U21203 (N_21203,N_18806,N_18078);
nand U21204 (N_21204,N_18049,N_18985);
and U21205 (N_21205,N_19070,N_19475);
or U21206 (N_21206,N_18196,N_19008);
nand U21207 (N_21207,N_18538,N_18310);
nand U21208 (N_21208,N_19802,N_18498);
nor U21209 (N_21209,N_19172,N_19320);
nand U21210 (N_21210,N_18189,N_18666);
and U21211 (N_21211,N_17937,N_18063);
nand U21212 (N_21212,N_19657,N_18927);
nor U21213 (N_21213,N_19527,N_18362);
nand U21214 (N_21214,N_18958,N_19285);
nand U21215 (N_21215,N_17593,N_19095);
nor U21216 (N_21216,N_17611,N_18048);
or U21217 (N_21217,N_19658,N_19946);
or U21218 (N_21218,N_19470,N_19286);
or U21219 (N_21219,N_18951,N_18497);
nand U21220 (N_21220,N_19422,N_18482);
or U21221 (N_21221,N_19600,N_19563);
nor U21222 (N_21222,N_18184,N_18169);
or U21223 (N_21223,N_18734,N_19888);
and U21224 (N_21224,N_19896,N_18625);
nand U21225 (N_21225,N_18361,N_18133);
or U21226 (N_21226,N_19894,N_18087);
or U21227 (N_21227,N_18239,N_19997);
or U21228 (N_21228,N_19678,N_17763);
nor U21229 (N_21229,N_19886,N_19165);
and U21230 (N_21230,N_18818,N_19972);
nor U21231 (N_21231,N_19219,N_18039);
or U21232 (N_21232,N_18139,N_18118);
and U21233 (N_21233,N_19260,N_19201);
and U21234 (N_21234,N_17514,N_18110);
nand U21235 (N_21235,N_19729,N_18385);
or U21236 (N_21236,N_19145,N_18905);
and U21237 (N_21237,N_18851,N_17936);
and U21238 (N_21238,N_18382,N_19207);
nand U21239 (N_21239,N_19111,N_19259);
nand U21240 (N_21240,N_19911,N_17940);
nand U21241 (N_21241,N_18944,N_18106);
nand U21242 (N_21242,N_19351,N_18367);
nor U21243 (N_21243,N_17912,N_18523);
and U21244 (N_21244,N_18027,N_18238);
and U21245 (N_21245,N_18530,N_19346);
or U21246 (N_21246,N_18612,N_17907);
or U21247 (N_21247,N_18381,N_19655);
and U21248 (N_21248,N_18923,N_17505);
or U21249 (N_21249,N_18527,N_19101);
nor U21250 (N_21250,N_19503,N_18032);
or U21251 (N_21251,N_19435,N_18496);
nor U21252 (N_21252,N_18505,N_18546);
nand U21253 (N_21253,N_18453,N_19519);
nor U21254 (N_21254,N_19342,N_18833);
and U21255 (N_21255,N_18064,N_18061);
nand U21256 (N_21256,N_18405,N_18562);
nand U21257 (N_21257,N_18167,N_18557);
nand U21258 (N_21258,N_18597,N_18120);
nor U21259 (N_21259,N_19402,N_18695);
nor U21260 (N_21260,N_17747,N_19388);
and U21261 (N_21261,N_17923,N_18855);
and U21262 (N_21262,N_17569,N_18070);
and U21263 (N_21263,N_19372,N_17810);
nand U21264 (N_21264,N_17701,N_17909);
and U21265 (N_21265,N_19392,N_19743);
nor U21266 (N_21266,N_19510,N_18313);
and U21267 (N_21267,N_19668,N_19884);
nor U21268 (N_21268,N_19959,N_19908);
nor U21269 (N_21269,N_18766,N_17574);
and U21270 (N_21270,N_18570,N_17964);
nor U21271 (N_21271,N_18808,N_17774);
nor U21272 (N_21272,N_18903,N_18047);
and U21273 (N_21273,N_17991,N_18479);
nand U21274 (N_21274,N_19082,N_18637);
xor U21275 (N_21275,N_19524,N_18471);
nand U21276 (N_21276,N_17702,N_18659);
nand U21277 (N_21277,N_19367,N_19157);
nand U21278 (N_21278,N_19140,N_18371);
or U21279 (N_21279,N_19023,N_19118);
nand U21280 (N_21280,N_18496,N_19995);
or U21281 (N_21281,N_19773,N_19329);
nor U21282 (N_21282,N_19868,N_17664);
or U21283 (N_21283,N_18472,N_18870);
nor U21284 (N_21284,N_19384,N_18998);
and U21285 (N_21285,N_17790,N_18760);
nor U21286 (N_21286,N_19433,N_18569);
nor U21287 (N_21287,N_19380,N_18741);
nor U21288 (N_21288,N_18773,N_18087);
and U21289 (N_21289,N_19604,N_18022);
nand U21290 (N_21290,N_18337,N_19002);
nand U21291 (N_21291,N_19617,N_18309);
or U21292 (N_21292,N_17968,N_18146);
nor U21293 (N_21293,N_19682,N_19170);
nand U21294 (N_21294,N_19223,N_18784);
and U21295 (N_21295,N_18016,N_18138);
or U21296 (N_21296,N_19323,N_19957);
nor U21297 (N_21297,N_18771,N_18908);
nor U21298 (N_21298,N_19656,N_18840);
nand U21299 (N_21299,N_19309,N_19634);
nand U21300 (N_21300,N_19912,N_18691);
and U21301 (N_21301,N_18895,N_19098);
nand U21302 (N_21302,N_18964,N_18736);
nor U21303 (N_21303,N_19041,N_18510);
nor U21304 (N_21304,N_19572,N_18476);
nor U21305 (N_21305,N_19399,N_18836);
or U21306 (N_21306,N_18318,N_19031);
or U21307 (N_21307,N_19215,N_18710);
or U21308 (N_21308,N_19037,N_18090);
nor U21309 (N_21309,N_19023,N_17752);
nand U21310 (N_21310,N_18551,N_19736);
nand U21311 (N_21311,N_18149,N_19193);
or U21312 (N_21312,N_18180,N_17969);
nor U21313 (N_21313,N_18408,N_18675);
nor U21314 (N_21314,N_18042,N_19864);
or U21315 (N_21315,N_17685,N_19338);
nor U21316 (N_21316,N_19656,N_19682);
or U21317 (N_21317,N_19643,N_17585);
or U21318 (N_21318,N_19346,N_19000);
nand U21319 (N_21319,N_17939,N_18829);
nor U21320 (N_21320,N_18440,N_19756);
nor U21321 (N_21321,N_18390,N_19331);
and U21322 (N_21322,N_18249,N_19866);
and U21323 (N_21323,N_17789,N_18431);
nor U21324 (N_21324,N_18865,N_18419);
nand U21325 (N_21325,N_19325,N_19839);
and U21326 (N_21326,N_18185,N_17914);
or U21327 (N_21327,N_18325,N_18407);
and U21328 (N_21328,N_19118,N_17658);
nand U21329 (N_21329,N_19545,N_18723);
nand U21330 (N_21330,N_19461,N_19138);
and U21331 (N_21331,N_19166,N_19291);
nor U21332 (N_21332,N_18320,N_19156);
and U21333 (N_21333,N_19156,N_18049);
and U21334 (N_21334,N_18137,N_17761);
or U21335 (N_21335,N_17645,N_17716);
nor U21336 (N_21336,N_19312,N_18112);
or U21337 (N_21337,N_19020,N_17726);
and U21338 (N_21338,N_18407,N_18759);
and U21339 (N_21339,N_19326,N_17532);
or U21340 (N_21340,N_18227,N_19623);
or U21341 (N_21341,N_18198,N_18686);
nor U21342 (N_21342,N_17751,N_19054);
or U21343 (N_21343,N_19133,N_19549);
and U21344 (N_21344,N_18648,N_18426);
and U21345 (N_21345,N_19864,N_18307);
and U21346 (N_21346,N_19615,N_17989);
or U21347 (N_21347,N_19485,N_19147);
or U21348 (N_21348,N_19222,N_18339);
or U21349 (N_21349,N_18868,N_19254);
nor U21350 (N_21350,N_17681,N_19265);
and U21351 (N_21351,N_17719,N_18841);
and U21352 (N_21352,N_18186,N_19752);
and U21353 (N_21353,N_18775,N_18591);
nand U21354 (N_21354,N_17883,N_19371);
nand U21355 (N_21355,N_19256,N_19405);
or U21356 (N_21356,N_18607,N_19508);
and U21357 (N_21357,N_18683,N_19722);
nand U21358 (N_21358,N_19051,N_17749);
or U21359 (N_21359,N_18594,N_19913);
or U21360 (N_21360,N_18885,N_18947);
nor U21361 (N_21361,N_18378,N_19768);
nand U21362 (N_21362,N_19749,N_19918);
or U21363 (N_21363,N_18953,N_18349);
and U21364 (N_21364,N_19668,N_19425);
nand U21365 (N_21365,N_19545,N_19541);
and U21366 (N_21366,N_18367,N_19992);
nand U21367 (N_21367,N_19602,N_18985);
nand U21368 (N_21368,N_18949,N_19816);
nor U21369 (N_21369,N_19144,N_17646);
and U21370 (N_21370,N_18542,N_17616);
nor U21371 (N_21371,N_17819,N_17988);
nor U21372 (N_21372,N_19739,N_18062);
or U21373 (N_21373,N_17793,N_17844);
and U21374 (N_21374,N_18509,N_18562);
and U21375 (N_21375,N_17502,N_19085);
nand U21376 (N_21376,N_18225,N_17944);
or U21377 (N_21377,N_19519,N_19881);
or U21378 (N_21378,N_19204,N_19325);
nand U21379 (N_21379,N_17896,N_17729);
nand U21380 (N_21380,N_17880,N_18658);
nand U21381 (N_21381,N_18066,N_19024);
or U21382 (N_21382,N_18088,N_19543);
nor U21383 (N_21383,N_19207,N_17579);
nand U21384 (N_21384,N_19554,N_18451);
nand U21385 (N_21385,N_18344,N_19178);
nand U21386 (N_21386,N_19389,N_18123);
nor U21387 (N_21387,N_19189,N_18488);
and U21388 (N_21388,N_17659,N_17819);
or U21389 (N_21389,N_18116,N_18338);
nand U21390 (N_21390,N_18030,N_18246);
and U21391 (N_21391,N_17855,N_18931);
nor U21392 (N_21392,N_19701,N_18532);
or U21393 (N_21393,N_18201,N_17745);
nor U21394 (N_21394,N_17780,N_18020);
and U21395 (N_21395,N_19916,N_19069);
nand U21396 (N_21396,N_18119,N_19117);
nand U21397 (N_21397,N_19807,N_18941);
nand U21398 (N_21398,N_19409,N_19313);
or U21399 (N_21399,N_19325,N_18563);
or U21400 (N_21400,N_18506,N_18103);
and U21401 (N_21401,N_18510,N_19642);
and U21402 (N_21402,N_18011,N_18730);
nor U21403 (N_21403,N_18462,N_18409);
and U21404 (N_21404,N_19580,N_19905);
and U21405 (N_21405,N_17798,N_18627);
nor U21406 (N_21406,N_18803,N_19993);
and U21407 (N_21407,N_19858,N_18061);
and U21408 (N_21408,N_19021,N_18884);
nand U21409 (N_21409,N_17543,N_17905);
nor U21410 (N_21410,N_19386,N_19544);
nor U21411 (N_21411,N_17909,N_18857);
nand U21412 (N_21412,N_18939,N_19279);
nand U21413 (N_21413,N_19100,N_19617);
and U21414 (N_21414,N_17621,N_19573);
or U21415 (N_21415,N_18452,N_19609);
and U21416 (N_21416,N_17863,N_17580);
and U21417 (N_21417,N_19022,N_19331);
nor U21418 (N_21418,N_19297,N_19121);
nand U21419 (N_21419,N_17890,N_18567);
and U21420 (N_21420,N_19438,N_18826);
nor U21421 (N_21421,N_19335,N_18875);
and U21422 (N_21422,N_19679,N_18234);
nand U21423 (N_21423,N_18791,N_19182);
or U21424 (N_21424,N_18689,N_18117);
or U21425 (N_21425,N_17694,N_19457);
nor U21426 (N_21426,N_17848,N_19022);
nand U21427 (N_21427,N_18494,N_17639);
nor U21428 (N_21428,N_19295,N_18460);
or U21429 (N_21429,N_18056,N_19194);
nand U21430 (N_21430,N_17938,N_17592);
nor U21431 (N_21431,N_17599,N_19515);
or U21432 (N_21432,N_19164,N_19747);
nor U21433 (N_21433,N_18958,N_17642);
nand U21434 (N_21434,N_18613,N_17512);
nand U21435 (N_21435,N_19583,N_18571);
and U21436 (N_21436,N_17874,N_18070);
nor U21437 (N_21437,N_19869,N_19919);
and U21438 (N_21438,N_18300,N_17881);
nor U21439 (N_21439,N_18217,N_18637);
nor U21440 (N_21440,N_19655,N_18014);
nand U21441 (N_21441,N_18833,N_18522);
nor U21442 (N_21442,N_19722,N_17722);
nand U21443 (N_21443,N_19379,N_18415);
nor U21444 (N_21444,N_18204,N_18291);
nor U21445 (N_21445,N_18141,N_18567);
nand U21446 (N_21446,N_18466,N_18222);
and U21447 (N_21447,N_18748,N_17771);
and U21448 (N_21448,N_18624,N_17762);
and U21449 (N_21449,N_19532,N_17914);
nor U21450 (N_21450,N_19179,N_17849);
nand U21451 (N_21451,N_18621,N_17502);
nor U21452 (N_21452,N_18846,N_19273);
and U21453 (N_21453,N_18057,N_18859);
or U21454 (N_21454,N_19490,N_19261);
or U21455 (N_21455,N_19302,N_18971);
or U21456 (N_21456,N_18639,N_19143);
and U21457 (N_21457,N_19847,N_18782);
and U21458 (N_21458,N_17878,N_19880);
nand U21459 (N_21459,N_19011,N_19844);
or U21460 (N_21460,N_18265,N_19760);
and U21461 (N_21461,N_18448,N_17757);
nand U21462 (N_21462,N_18490,N_17805);
or U21463 (N_21463,N_17740,N_17932);
or U21464 (N_21464,N_18361,N_18427);
nor U21465 (N_21465,N_18022,N_18386);
or U21466 (N_21466,N_18321,N_18650);
and U21467 (N_21467,N_17680,N_19391);
or U21468 (N_21468,N_17903,N_18441);
or U21469 (N_21469,N_19441,N_18507);
nor U21470 (N_21470,N_18901,N_18667);
nand U21471 (N_21471,N_18981,N_19171);
and U21472 (N_21472,N_19840,N_18627);
nand U21473 (N_21473,N_17859,N_18948);
nor U21474 (N_21474,N_19214,N_19503);
nand U21475 (N_21475,N_19487,N_17598);
nand U21476 (N_21476,N_18177,N_18633);
and U21477 (N_21477,N_17757,N_18071);
nor U21478 (N_21478,N_18511,N_19062);
nand U21479 (N_21479,N_19447,N_18653);
or U21480 (N_21480,N_19920,N_18472);
nand U21481 (N_21481,N_18589,N_18099);
or U21482 (N_21482,N_18164,N_19893);
or U21483 (N_21483,N_18958,N_19655);
or U21484 (N_21484,N_19202,N_19140);
and U21485 (N_21485,N_17991,N_18456);
nand U21486 (N_21486,N_19764,N_19505);
nor U21487 (N_21487,N_17999,N_17837);
xnor U21488 (N_21488,N_17949,N_18716);
nand U21489 (N_21489,N_17806,N_18099);
and U21490 (N_21490,N_18968,N_19776);
nand U21491 (N_21491,N_18062,N_19572);
and U21492 (N_21492,N_18775,N_18585);
nand U21493 (N_21493,N_18286,N_19151);
and U21494 (N_21494,N_17937,N_18458);
nand U21495 (N_21495,N_18511,N_18425);
and U21496 (N_21496,N_17631,N_18132);
and U21497 (N_21497,N_17956,N_19301);
or U21498 (N_21498,N_18438,N_19395);
or U21499 (N_21499,N_18764,N_19871);
and U21500 (N_21500,N_18829,N_19161);
or U21501 (N_21501,N_17769,N_18782);
and U21502 (N_21502,N_19954,N_19120);
nand U21503 (N_21503,N_18302,N_17931);
nand U21504 (N_21504,N_18792,N_17849);
or U21505 (N_21505,N_17745,N_18799);
and U21506 (N_21506,N_18984,N_19983);
nand U21507 (N_21507,N_17690,N_19952);
nor U21508 (N_21508,N_18354,N_18521);
nor U21509 (N_21509,N_17880,N_18133);
or U21510 (N_21510,N_18398,N_18889);
nand U21511 (N_21511,N_19908,N_18855);
xor U21512 (N_21512,N_19661,N_19929);
nand U21513 (N_21513,N_18702,N_19735);
nor U21514 (N_21514,N_18923,N_18913);
nand U21515 (N_21515,N_18701,N_17686);
nor U21516 (N_21516,N_19208,N_19908);
nor U21517 (N_21517,N_18098,N_19116);
nor U21518 (N_21518,N_18757,N_19377);
nor U21519 (N_21519,N_18026,N_19674);
nor U21520 (N_21520,N_19842,N_18893);
or U21521 (N_21521,N_18512,N_19508);
nor U21522 (N_21522,N_19753,N_19789);
and U21523 (N_21523,N_19395,N_19087);
nand U21524 (N_21524,N_19390,N_18688);
nor U21525 (N_21525,N_19204,N_18754);
nand U21526 (N_21526,N_17925,N_19618);
nand U21527 (N_21527,N_19683,N_19526);
nand U21528 (N_21528,N_17626,N_19332);
nand U21529 (N_21529,N_18029,N_19795);
nand U21530 (N_21530,N_18961,N_19255);
and U21531 (N_21531,N_18891,N_18830);
or U21532 (N_21532,N_19686,N_18305);
or U21533 (N_21533,N_17747,N_18419);
nor U21534 (N_21534,N_19853,N_19967);
and U21535 (N_21535,N_18294,N_19372);
nand U21536 (N_21536,N_17677,N_18441);
nor U21537 (N_21537,N_19933,N_18170);
nor U21538 (N_21538,N_17841,N_18112);
nand U21539 (N_21539,N_19154,N_19152);
or U21540 (N_21540,N_19379,N_19611);
and U21541 (N_21541,N_18585,N_19097);
nor U21542 (N_21542,N_19228,N_18214);
or U21543 (N_21543,N_18208,N_18105);
or U21544 (N_21544,N_18636,N_19397);
or U21545 (N_21545,N_18963,N_19447);
nand U21546 (N_21546,N_19326,N_17508);
and U21547 (N_21547,N_18891,N_18495);
and U21548 (N_21548,N_19703,N_19860);
nand U21549 (N_21549,N_18255,N_18626);
nor U21550 (N_21550,N_19909,N_17868);
and U21551 (N_21551,N_18459,N_18187);
or U21552 (N_21552,N_17623,N_19771);
nand U21553 (N_21553,N_19894,N_19612);
and U21554 (N_21554,N_19459,N_19102);
and U21555 (N_21555,N_19078,N_17728);
nor U21556 (N_21556,N_18874,N_19911);
nand U21557 (N_21557,N_18700,N_18655);
nor U21558 (N_21558,N_19917,N_18900);
nand U21559 (N_21559,N_18287,N_19697);
or U21560 (N_21560,N_18025,N_18943);
and U21561 (N_21561,N_18011,N_18441);
and U21562 (N_21562,N_18679,N_18827);
and U21563 (N_21563,N_18759,N_17945);
nand U21564 (N_21564,N_19918,N_18873);
nor U21565 (N_21565,N_18398,N_17661);
and U21566 (N_21566,N_17530,N_18798);
or U21567 (N_21567,N_17660,N_18799);
or U21568 (N_21568,N_19880,N_17997);
nor U21569 (N_21569,N_18809,N_18279);
nand U21570 (N_21570,N_19092,N_18247);
or U21571 (N_21571,N_18216,N_18387);
nor U21572 (N_21572,N_17892,N_19049);
and U21573 (N_21573,N_17964,N_18793);
nand U21574 (N_21574,N_17563,N_18438);
and U21575 (N_21575,N_18753,N_18841);
nor U21576 (N_21576,N_19145,N_18405);
nand U21577 (N_21577,N_19255,N_17610);
and U21578 (N_21578,N_17811,N_18218);
nand U21579 (N_21579,N_19297,N_17964);
nor U21580 (N_21580,N_19701,N_19620);
and U21581 (N_21581,N_18059,N_17788);
nand U21582 (N_21582,N_18715,N_18415);
nor U21583 (N_21583,N_19119,N_19295);
and U21584 (N_21584,N_18326,N_19397);
and U21585 (N_21585,N_18483,N_17946);
nand U21586 (N_21586,N_19224,N_18825);
nor U21587 (N_21587,N_18941,N_17808);
and U21588 (N_21588,N_19413,N_18101);
nand U21589 (N_21589,N_18973,N_17599);
or U21590 (N_21590,N_18104,N_18583);
nand U21591 (N_21591,N_17629,N_17736);
and U21592 (N_21592,N_19209,N_18557);
or U21593 (N_21593,N_19998,N_17860);
or U21594 (N_21594,N_19455,N_18759);
and U21595 (N_21595,N_19602,N_18761);
nand U21596 (N_21596,N_18094,N_18561);
and U21597 (N_21597,N_18293,N_19667);
nor U21598 (N_21598,N_17747,N_19107);
and U21599 (N_21599,N_18118,N_18381);
nor U21600 (N_21600,N_19858,N_18539);
nand U21601 (N_21601,N_18562,N_18421);
or U21602 (N_21602,N_18462,N_17911);
nand U21603 (N_21603,N_19965,N_19490);
nor U21604 (N_21604,N_19975,N_19404);
nor U21605 (N_21605,N_19919,N_18511);
and U21606 (N_21606,N_18050,N_18417);
nand U21607 (N_21607,N_18706,N_18744);
and U21608 (N_21608,N_19182,N_19156);
nor U21609 (N_21609,N_18167,N_19601);
and U21610 (N_21610,N_19900,N_18031);
nor U21611 (N_21611,N_18405,N_17614);
and U21612 (N_21612,N_18091,N_18333);
nand U21613 (N_21613,N_18873,N_17698);
and U21614 (N_21614,N_17819,N_18517);
nand U21615 (N_21615,N_18331,N_17733);
or U21616 (N_21616,N_19249,N_18463);
and U21617 (N_21617,N_19906,N_19568);
nor U21618 (N_21618,N_17777,N_19405);
nor U21619 (N_21619,N_18266,N_19154);
nand U21620 (N_21620,N_19642,N_18318);
and U21621 (N_21621,N_19499,N_18621);
nand U21622 (N_21622,N_18031,N_18673);
or U21623 (N_21623,N_18285,N_17801);
nor U21624 (N_21624,N_17805,N_19611);
and U21625 (N_21625,N_18429,N_19206);
or U21626 (N_21626,N_19866,N_17910);
nor U21627 (N_21627,N_19378,N_17534);
nor U21628 (N_21628,N_18190,N_18322);
nor U21629 (N_21629,N_18213,N_19038);
nand U21630 (N_21630,N_18136,N_19644);
nor U21631 (N_21631,N_17531,N_18704);
and U21632 (N_21632,N_17607,N_19053);
and U21633 (N_21633,N_19485,N_19259);
nor U21634 (N_21634,N_18602,N_18612);
and U21635 (N_21635,N_19192,N_17627);
or U21636 (N_21636,N_19268,N_17761);
nand U21637 (N_21637,N_17898,N_19091);
or U21638 (N_21638,N_18477,N_19645);
nand U21639 (N_21639,N_18381,N_18087);
or U21640 (N_21640,N_19895,N_18353);
and U21641 (N_21641,N_18737,N_18561);
nor U21642 (N_21642,N_18886,N_17596);
nor U21643 (N_21643,N_19864,N_18630);
nand U21644 (N_21644,N_19467,N_18688);
nand U21645 (N_21645,N_19797,N_18075);
or U21646 (N_21646,N_18893,N_19358);
and U21647 (N_21647,N_18233,N_19975);
or U21648 (N_21648,N_17918,N_19740);
nand U21649 (N_21649,N_18052,N_18906);
nor U21650 (N_21650,N_18835,N_18617);
nand U21651 (N_21651,N_19135,N_18834);
or U21652 (N_21652,N_18144,N_17815);
nor U21653 (N_21653,N_19420,N_19121);
or U21654 (N_21654,N_19622,N_19617);
and U21655 (N_21655,N_18154,N_17849);
and U21656 (N_21656,N_18776,N_19852);
nor U21657 (N_21657,N_19112,N_17812);
nand U21658 (N_21658,N_18160,N_19000);
or U21659 (N_21659,N_18767,N_19832);
nand U21660 (N_21660,N_19640,N_19370);
or U21661 (N_21661,N_18744,N_18530);
and U21662 (N_21662,N_17647,N_18431);
nand U21663 (N_21663,N_17589,N_18652);
or U21664 (N_21664,N_19062,N_17895);
nor U21665 (N_21665,N_18462,N_19118);
and U21666 (N_21666,N_19401,N_18730);
nand U21667 (N_21667,N_19040,N_17610);
or U21668 (N_21668,N_18495,N_19407);
and U21669 (N_21669,N_18613,N_18348);
and U21670 (N_21670,N_18357,N_18450);
nand U21671 (N_21671,N_18294,N_19025);
or U21672 (N_21672,N_19411,N_18730);
or U21673 (N_21673,N_17552,N_19968);
or U21674 (N_21674,N_18475,N_17647);
or U21675 (N_21675,N_19084,N_18475);
or U21676 (N_21676,N_18399,N_17555);
and U21677 (N_21677,N_18607,N_19260);
or U21678 (N_21678,N_19370,N_17927);
nand U21679 (N_21679,N_19006,N_17533);
or U21680 (N_21680,N_18837,N_18126);
nand U21681 (N_21681,N_18371,N_19746);
nand U21682 (N_21682,N_18534,N_17918);
and U21683 (N_21683,N_18103,N_18650);
and U21684 (N_21684,N_18079,N_18475);
nand U21685 (N_21685,N_18202,N_19736);
nand U21686 (N_21686,N_19791,N_17531);
nand U21687 (N_21687,N_18853,N_18927);
or U21688 (N_21688,N_17908,N_19112);
nor U21689 (N_21689,N_18733,N_18508);
nand U21690 (N_21690,N_18823,N_17518);
nand U21691 (N_21691,N_17951,N_18037);
nor U21692 (N_21692,N_19385,N_18379);
and U21693 (N_21693,N_17920,N_17717);
and U21694 (N_21694,N_18420,N_19652);
or U21695 (N_21695,N_19049,N_18106);
or U21696 (N_21696,N_19438,N_19448);
or U21697 (N_21697,N_17562,N_19225);
nor U21698 (N_21698,N_19676,N_19204);
or U21699 (N_21699,N_19696,N_19750);
or U21700 (N_21700,N_18717,N_17550);
or U21701 (N_21701,N_19155,N_17820);
or U21702 (N_21702,N_18319,N_19137);
nand U21703 (N_21703,N_19370,N_18383);
nor U21704 (N_21704,N_18015,N_19388);
nand U21705 (N_21705,N_18911,N_18644);
and U21706 (N_21706,N_18131,N_18702);
or U21707 (N_21707,N_18693,N_18623);
or U21708 (N_21708,N_19896,N_18083);
nand U21709 (N_21709,N_19538,N_18146);
or U21710 (N_21710,N_19157,N_19852);
or U21711 (N_21711,N_19554,N_18329);
nand U21712 (N_21712,N_17746,N_17895);
and U21713 (N_21713,N_19366,N_18142);
nor U21714 (N_21714,N_17987,N_19079);
nor U21715 (N_21715,N_18329,N_18709);
or U21716 (N_21716,N_18363,N_19014);
nand U21717 (N_21717,N_18564,N_19155);
and U21718 (N_21718,N_19150,N_17896);
nor U21719 (N_21719,N_19553,N_17953);
or U21720 (N_21720,N_18722,N_18046);
or U21721 (N_21721,N_17676,N_18753);
nor U21722 (N_21722,N_19762,N_18081);
nor U21723 (N_21723,N_17776,N_17654);
or U21724 (N_21724,N_19621,N_19885);
nor U21725 (N_21725,N_18989,N_17661);
nor U21726 (N_21726,N_18970,N_19375);
and U21727 (N_21727,N_19039,N_19006);
and U21728 (N_21728,N_18433,N_18223);
nand U21729 (N_21729,N_17872,N_18406);
and U21730 (N_21730,N_19303,N_19011);
nand U21731 (N_21731,N_19491,N_18034);
nand U21732 (N_21732,N_19888,N_19770);
nor U21733 (N_21733,N_19197,N_19356);
nand U21734 (N_21734,N_18719,N_19934);
nand U21735 (N_21735,N_19639,N_18672);
nor U21736 (N_21736,N_18674,N_18544);
or U21737 (N_21737,N_18734,N_19642);
nor U21738 (N_21738,N_17589,N_19538);
nor U21739 (N_21739,N_17575,N_19915);
or U21740 (N_21740,N_18844,N_18962);
and U21741 (N_21741,N_18863,N_17554);
or U21742 (N_21742,N_18144,N_18589);
and U21743 (N_21743,N_19699,N_19572);
or U21744 (N_21744,N_18132,N_18933);
nor U21745 (N_21745,N_18326,N_18789);
nand U21746 (N_21746,N_19550,N_19601);
or U21747 (N_21747,N_18322,N_18961);
nor U21748 (N_21748,N_17629,N_19667);
nor U21749 (N_21749,N_18885,N_19938);
or U21750 (N_21750,N_18149,N_18691);
or U21751 (N_21751,N_18020,N_17561);
nor U21752 (N_21752,N_19539,N_19654);
or U21753 (N_21753,N_18658,N_19387);
nor U21754 (N_21754,N_19315,N_19714);
or U21755 (N_21755,N_19801,N_19049);
or U21756 (N_21756,N_18703,N_19474);
xnor U21757 (N_21757,N_19430,N_18448);
or U21758 (N_21758,N_19900,N_18181);
and U21759 (N_21759,N_17860,N_19293);
nand U21760 (N_21760,N_18909,N_19713);
or U21761 (N_21761,N_17543,N_19675);
nand U21762 (N_21762,N_18219,N_19865);
or U21763 (N_21763,N_18885,N_18045);
and U21764 (N_21764,N_18338,N_18276);
nor U21765 (N_21765,N_18910,N_19441);
or U21766 (N_21766,N_19112,N_19441);
or U21767 (N_21767,N_18234,N_19894);
nor U21768 (N_21768,N_19040,N_17641);
and U21769 (N_21769,N_19491,N_18495);
nand U21770 (N_21770,N_19668,N_19779);
nand U21771 (N_21771,N_17642,N_19180);
nor U21772 (N_21772,N_18553,N_19755);
and U21773 (N_21773,N_18352,N_19157);
or U21774 (N_21774,N_19084,N_17690);
and U21775 (N_21775,N_17746,N_19592);
nor U21776 (N_21776,N_17963,N_19094);
nand U21777 (N_21777,N_17696,N_17839);
nor U21778 (N_21778,N_19422,N_18466);
nor U21779 (N_21779,N_17529,N_19521);
and U21780 (N_21780,N_18149,N_18075);
or U21781 (N_21781,N_18525,N_17811);
and U21782 (N_21782,N_19936,N_17773);
nand U21783 (N_21783,N_19805,N_18841);
nor U21784 (N_21784,N_18156,N_18487);
nand U21785 (N_21785,N_19961,N_19713);
and U21786 (N_21786,N_18036,N_18884);
and U21787 (N_21787,N_19298,N_17682);
nor U21788 (N_21788,N_17692,N_19573);
and U21789 (N_21789,N_17868,N_19039);
or U21790 (N_21790,N_17957,N_19226);
nand U21791 (N_21791,N_19644,N_18554);
or U21792 (N_21792,N_19258,N_19216);
nor U21793 (N_21793,N_18283,N_19360);
or U21794 (N_21794,N_18518,N_19280);
and U21795 (N_21795,N_19080,N_18964);
and U21796 (N_21796,N_19381,N_18652);
or U21797 (N_21797,N_19806,N_18854);
xnor U21798 (N_21798,N_18487,N_19070);
or U21799 (N_21799,N_17684,N_18519);
or U21800 (N_21800,N_17518,N_18074);
nand U21801 (N_21801,N_17606,N_19778);
nand U21802 (N_21802,N_19769,N_19125);
nor U21803 (N_21803,N_18786,N_17541);
nand U21804 (N_21804,N_18476,N_18762);
and U21805 (N_21805,N_19745,N_18698);
nor U21806 (N_21806,N_18781,N_17932);
nor U21807 (N_21807,N_19578,N_17884);
and U21808 (N_21808,N_18583,N_17821);
and U21809 (N_21809,N_19523,N_17844);
nor U21810 (N_21810,N_18030,N_18707);
nor U21811 (N_21811,N_18344,N_19932);
or U21812 (N_21812,N_18608,N_18633);
nor U21813 (N_21813,N_19526,N_19493);
xor U21814 (N_21814,N_17970,N_17837);
nand U21815 (N_21815,N_18724,N_18684);
or U21816 (N_21816,N_19560,N_18901);
nor U21817 (N_21817,N_19650,N_17789);
nor U21818 (N_21818,N_18655,N_18239);
nor U21819 (N_21819,N_17854,N_19990);
or U21820 (N_21820,N_18627,N_18892);
nor U21821 (N_21821,N_19511,N_19725);
and U21822 (N_21822,N_18157,N_18468);
nand U21823 (N_21823,N_19911,N_17566);
or U21824 (N_21824,N_18141,N_19102);
and U21825 (N_21825,N_18199,N_17566);
nand U21826 (N_21826,N_19459,N_18735);
and U21827 (N_21827,N_17875,N_19289);
and U21828 (N_21828,N_18631,N_19757);
nand U21829 (N_21829,N_18469,N_19630);
nand U21830 (N_21830,N_19721,N_18872);
and U21831 (N_21831,N_18432,N_18888);
and U21832 (N_21832,N_19671,N_17976);
or U21833 (N_21833,N_18500,N_17961);
or U21834 (N_21834,N_17547,N_19331);
nor U21835 (N_21835,N_19088,N_19511);
nor U21836 (N_21836,N_18995,N_17606);
nor U21837 (N_21837,N_17885,N_19727);
nand U21838 (N_21838,N_18973,N_19996);
or U21839 (N_21839,N_19236,N_18892);
nor U21840 (N_21840,N_17696,N_19479);
nand U21841 (N_21841,N_19272,N_18034);
and U21842 (N_21842,N_18534,N_19352);
or U21843 (N_21843,N_18320,N_18048);
nor U21844 (N_21844,N_17897,N_19569);
or U21845 (N_21845,N_18415,N_19309);
nor U21846 (N_21846,N_19703,N_19162);
nand U21847 (N_21847,N_18291,N_18912);
or U21848 (N_21848,N_19178,N_18861);
and U21849 (N_21849,N_18183,N_17874);
or U21850 (N_21850,N_19639,N_19447);
nor U21851 (N_21851,N_19598,N_19642);
or U21852 (N_21852,N_19604,N_18109);
nor U21853 (N_21853,N_19296,N_18196);
or U21854 (N_21854,N_18492,N_19265);
and U21855 (N_21855,N_18796,N_19435);
nor U21856 (N_21856,N_18587,N_17693);
nand U21857 (N_21857,N_19768,N_18718);
nor U21858 (N_21858,N_18544,N_18762);
or U21859 (N_21859,N_19253,N_19957);
nor U21860 (N_21860,N_17691,N_19698);
and U21861 (N_21861,N_18987,N_17759);
xnor U21862 (N_21862,N_17838,N_19999);
and U21863 (N_21863,N_19694,N_19950);
nand U21864 (N_21864,N_18664,N_17924);
or U21865 (N_21865,N_18359,N_17905);
and U21866 (N_21866,N_17840,N_18438);
nand U21867 (N_21867,N_18704,N_17717);
and U21868 (N_21868,N_19270,N_18373);
and U21869 (N_21869,N_18004,N_17921);
nand U21870 (N_21870,N_18993,N_18710);
or U21871 (N_21871,N_18941,N_18631);
nand U21872 (N_21872,N_18607,N_17662);
nand U21873 (N_21873,N_19964,N_18967);
nor U21874 (N_21874,N_19065,N_19840);
nor U21875 (N_21875,N_19450,N_19849);
nand U21876 (N_21876,N_18700,N_19111);
or U21877 (N_21877,N_18401,N_18950);
or U21878 (N_21878,N_18350,N_18217);
nand U21879 (N_21879,N_19366,N_19701);
nor U21880 (N_21880,N_18374,N_18816);
or U21881 (N_21881,N_19048,N_19776);
and U21882 (N_21882,N_18191,N_18720);
nand U21883 (N_21883,N_19961,N_18513);
and U21884 (N_21884,N_17963,N_18178);
and U21885 (N_21885,N_19907,N_19828);
nor U21886 (N_21886,N_18503,N_19636);
nand U21887 (N_21887,N_19757,N_19337);
or U21888 (N_21888,N_19625,N_18923);
or U21889 (N_21889,N_18074,N_18511);
nand U21890 (N_21890,N_19412,N_18827);
nor U21891 (N_21891,N_19903,N_18677);
and U21892 (N_21892,N_18416,N_17624);
nor U21893 (N_21893,N_18243,N_18576);
or U21894 (N_21894,N_19041,N_17827);
or U21895 (N_21895,N_18083,N_17866);
nor U21896 (N_21896,N_18720,N_19590);
nor U21897 (N_21897,N_19278,N_18995);
or U21898 (N_21898,N_19628,N_19152);
and U21899 (N_21899,N_19790,N_17641);
nand U21900 (N_21900,N_19825,N_19541);
or U21901 (N_21901,N_19357,N_18334);
nand U21902 (N_21902,N_17813,N_19550);
nor U21903 (N_21903,N_18886,N_18685);
nor U21904 (N_21904,N_19679,N_18673);
and U21905 (N_21905,N_18291,N_19361);
nor U21906 (N_21906,N_18563,N_18362);
and U21907 (N_21907,N_19166,N_19479);
nand U21908 (N_21908,N_18975,N_17869);
nor U21909 (N_21909,N_18830,N_19907);
or U21910 (N_21910,N_19866,N_19841);
or U21911 (N_21911,N_18137,N_18899);
and U21912 (N_21912,N_19111,N_19982);
nor U21913 (N_21913,N_17850,N_19778);
and U21914 (N_21914,N_18075,N_19814);
or U21915 (N_21915,N_18103,N_19557);
or U21916 (N_21916,N_18340,N_18557);
and U21917 (N_21917,N_19594,N_19694);
and U21918 (N_21918,N_19536,N_19701);
nor U21919 (N_21919,N_19908,N_19993);
nand U21920 (N_21920,N_19949,N_19055);
xor U21921 (N_21921,N_17562,N_18757);
nand U21922 (N_21922,N_19234,N_18215);
and U21923 (N_21923,N_19019,N_18937);
and U21924 (N_21924,N_19535,N_18436);
or U21925 (N_21925,N_19361,N_19612);
and U21926 (N_21926,N_19901,N_18363);
nor U21927 (N_21927,N_18038,N_19640);
or U21928 (N_21928,N_19044,N_19258);
nand U21929 (N_21929,N_18696,N_18700);
nand U21930 (N_21930,N_18324,N_19846);
or U21931 (N_21931,N_18230,N_19684);
or U21932 (N_21932,N_19087,N_19231);
or U21933 (N_21933,N_18498,N_18877);
or U21934 (N_21934,N_17788,N_18354);
nor U21935 (N_21935,N_18610,N_17547);
nand U21936 (N_21936,N_19221,N_18533);
nand U21937 (N_21937,N_17733,N_19539);
nor U21938 (N_21938,N_18570,N_19556);
nand U21939 (N_21939,N_19558,N_19166);
or U21940 (N_21940,N_19581,N_18693);
nand U21941 (N_21941,N_18753,N_18674);
and U21942 (N_21942,N_18826,N_19141);
nor U21943 (N_21943,N_18535,N_18221);
or U21944 (N_21944,N_17773,N_17850);
and U21945 (N_21945,N_18227,N_18918);
nor U21946 (N_21946,N_19855,N_17810);
or U21947 (N_21947,N_18770,N_19247);
nand U21948 (N_21948,N_19154,N_18287);
nand U21949 (N_21949,N_19103,N_18055);
and U21950 (N_21950,N_19167,N_17685);
or U21951 (N_21951,N_19855,N_18026);
nor U21952 (N_21952,N_18026,N_18858);
nor U21953 (N_21953,N_18183,N_18074);
nor U21954 (N_21954,N_19966,N_19036);
xor U21955 (N_21955,N_19710,N_18339);
or U21956 (N_21956,N_18116,N_17529);
or U21957 (N_21957,N_19735,N_17957);
or U21958 (N_21958,N_19455,N_18787);
or U21959 (N_21959,N_18147,N_19054);
nand U21960 (N_21960,N_19170,N_19136);
or U21961 (N_21961,N_17875,N_19060);
nand U21962 (N_21962,N_19431,N_19723);
and U21963 (N_21963,N_19219,N_17717);
and U21964 (N_21964,N_19198,N_18816);
and U21965 (N_21965,N_18559,N_19724);
nor U21966 (N_21966,N_19910,N_17908);
and U21967 (N_21967,N_19405,N_17877);
and U21968 (N_21968,N_18306,N_17667);
nand U21969 (N_21969,N_18430,N_17930);
or U21970 (N_21970,N_18932,N_18448);
nand U21971 (N_21971,N_19857,N_17588);
or U21972 (N_21972,N_18914,N_17665);
or U21973 (N_21973,N_18310,N_18430);
nor U21974 (N_21974,N_19833,N_19933);
nor U21975 (N_21975,N_19571,N_17707);
or U21976 (N_21976,N_18374,N_19373);
nand U21977 (N_21977,N_19140,N_17873);
nand U21978 (N_21978,N_19157,N_18065);
nand U21979 (N_21979,N_19345,N_19652);
nor U21980 (N_21980,N_18274,N_19610);
or U21981 (N_21981,N_19780,N_19385);
or U21982 (N_21982,N_17971,N_18922);
nand U21983 (N_21983,N_19592,N_19127);
or U21984 (N_21984,N_18660,N_18552);
and U21985 (N_21985,N_19718,N_19513);
or U21986 (N_21986,N_19187,N_19593);
nor U21987 (N_21987,N_19286,N_18058);
and U21988 (N_21988,N_19719,N_19621);
and U21989 (N_21989,N_18720,N_19599);
or U21990 (N_21990,N_19157,N_19139);
nor U21991 (N_21991,N_18712,N_19466);
nor U21992 (N_21992,N_19240,N_19615);
and U21993 (N_21993,N_18252,N_19975);
or U21994 (N_21994,N_18427,N_18315);
xor U21995 (N_21995,N_17519,N_17850);
and U21996 (N_21996,N_17702,N_17964);
and U21997 (N_21997,N_18547,N_18759);
or U21998 (N_21998,N_18330,N_19998);
nor U21999 (N_21999,N_18309,N_19584);
nor U22000 (N_22000,N_19308,N_18998);
and U22001 (N_22001,N_18171,N_19451);
and U22002 (N_22002,N_17888,N_18678);
or U22003 (N_22003,N_19563,N_17981);
nor U22004 (N_22004,N_19988,N_19265);
or U22005 (N_22005,N_18282,N_19498);
nor U22006 (N_22006,N_17962,N_17875);
and U22007 (N_22007,N_18083,N_18260);
nor U22008 (N_22008,N_19338,N_19069);
nand U22009 (N_22009,N_19696,N_18950);
and U22010 (N_22010,N_17920,N_18273);
and U22011 (N_22011,N_17687,N_17556);
and U22012 (N_22012,N_17968,N_18892);
nor U22013 (N_22013,N_18161,N_19424);
or U22014 (N_22014,N_19135,N_19803);
or U22015 (N_22015,N_19122,N_18676);
nor U22016 (N_22016,N_19023,N_18862);
nor U22017 (N_22017,N_19906,N_17549);
nor U22018 (N_22018,N_18390,N_17670);
and U22019 (N_22019,N_18296,N_18142);
nand U22020 (N_22020,N_18810,N_19184);
and U22021 (N_22021,N_17820,N_19134);
or U22022 (N_22022,N_18749,N_18931);
or U22023 (N_22023,N_19126,N_18203);
and U22024 (N_22024,N_19869,N_18762);
nor U22025 (N_22025,N_18209,N_19095);
nand U22026 (N_22026,N_19472,N_18586);
or U22027 (N_22027,N_19707,N_19466);
and U22028 (N_22028,N_18184,N_18733);
nand U22029 (N_22029,N_18559,N_19169);
nor U22030 (N_22030,N_19220,N_18434);
or U22031 (N_22031,N_18560,N_17608);
nor U22032 (N_22032,N_18648,N_18901);
or U22033 (N_22033,N_19055,N_18167);
nand U22034 (N_22034,N_18982,N_19597);
nand U22035 (N_22035,N_19429,N_18072);
and U22036 (N_22036,N_19616,N_19008);
or U22037 (N_22037,N_18202,N_18044);
nor U22038 (N_22038,N_17577,N_17540);
and U22039 (N_22039,N_18475,N_18100);
nor U22040 (N_22040,N_19342,N_18427);
nor U22041 (N_22041,N_18245,N_18322);
nand U22042 (N_22042,N_18068,N_17535);
or U22043 (N_22043,N_19967,N_19601);
or U22044 (N_22044,N_19034,N_19608);
nor U22045 (N_22045,N_17919,N_18908);
and U22046 (N_22046,N_18084,N_19510);
or U22047 (N_22047,N_19585,N_18285);
nand U22048 (N_22048,N_17783,N_19707);
nor U22049 (N_22049,N_18221,N_19127);
or U22050 (N_22050,N_18077,N_19152);
nand U22051 (N_22051,N_19656,N_18017);
or U22052 (N_22052,N_19047,N_19038);
nand U22053 (N_22053,N_19735,N_18051);
and U22054 (N_22054,N_18032,N_17517);
or U22055 (N_22055,N_19246,N_19822);
nor U22056 (N_22056,N_17526,N_18538);
nand U22057 (N_22057,N_19549,N_18161);
and U22058 (N_22058,N_18360,N_19554);
and U22059 (N_22059,N_18567,N_19517);
nand U22060 (N_22060,N_18299,N_18718);
and U22061 (N_22061,N_18153,N_19384);
nand U22062 (N_22062,N_19159,N_18071);
and U22063 (N_22063,N_19048,N_19251);
and U22064 (N_22064,N_19935,N_17998);
nand U22065 (N_22065,N_19066,N_18952);
nor U22066 (N_22066,N_19536,N_17748);
nand U22067 (N_22067,N_18055,N_18592);
nand U22068 (N_22068,N_17850,N_18185);
nor U22069 (N_22069,N_19545,N_18188);
nand U22070 (N_22070,N_19896,N_18363);
nand U22071 (N_22071,N_18088,N_19457);
or U22072 (N_22072,N_19150,N_18937);
nor U22073 (N_22073,N_18307,N_19479);
nor U22074 (N_22074,N_18111,N_19795);
nor U22075 (N_22075,N_19172,N_17892);
and U22076 (N_22076,N_19191,N_19898);
nand U22077 (N_22077,N_18769,N_18659);
nand U22078 (N_22078,N_18679,N_17585);
nand U22079 (N_22079,N_19076,N_18341);
nor U22080 (N_22080,N_18117,N_19577);
or U22081 (N_22081,N_18425,N_19824);
and U22082 (N_22082,N_19035,N_19834);
and U22083 (N_22083,N_19658,N_18311);
or U22084 (N_22084,N_17557,N_17767);
and U22085 (N_22085,N_18758,N_18429);
and U22086 (N_22086,N_19004,N_17626);
nand U22087 (N_22087,N_17683,N_17866);
nand U22088 (N_22088,N_19509,N_19244);
and U22089 (N_22089,N_17856,N_19844);
and U22090 (N_22090,N_17928,N_18150);
and U22091 (N_22091,N_17936,N_17661);
nor U22092 (N_22092,N_19486,N_18779);
and U22093 (N_22093,N_18175,N_19544);
nor U22094 (N_22094,N_18117,N_19415);
nand U22095 (N_22095,N_19498,N_17544);
nand U22096 (N_22096,N_17691,N_17896);
or U22097 (N_22097,N_17752,N_17660);
and U22098 (N_22098,N_19024,N_17824);
and U22099 (N_22099,N_18335,N_18571);
nand U22100 (N_22100,N_17877,N_19759);
nand U22101 (N_22101,N_18124,N_18948);
nand U22102 (N_22102,N_19828,N_19199);
nand U22103 (N_22103,N_17503,N_17950);
nor U22104 (N_22104,N_18963,N_18667);
or U22105 (N_22105,N_17859,N_18384);
and U22106 (N_22106,N_18895,N_19480);
nand U22107 (N_22107,N_17626,N_19320);
and U22108 (N_22108,N_19670,N_19292);
or U22109 (N_22109,N_17500,N_19403);
and U22110 (N_22110,N_17789,N_19810);
nand U22111 (N_22111,N_19587,N_17934);
or U22112 (N_22112,N_17965,N_18312);
nor U22113 (N_22113,N_19636,N_18704);
or U22114 (N_22114,N_19144,N_19895);
nor U22115 (N_22115,N_17926,N_18355);
nor U22116 (N_22116,N_18310,N_18236);
and U22117 (N_22117,N_19960,N_18882);
or U22118 (N_22118,N_19170,N_18079);
or U22119 (N_22119,N_19848,N_17520);
or U22120 (N_22120,N_19680,N_17605);
nor U22121 (N_22121,N_19463,N_18586);
nor U22122 (N_22122,N_17996,N_18664);
or U22123 (N_22123,N_19494,N_17956);
nor U22124 (N_22124,N_19248,N_17583);
nand U22125 (N_22125,N_17897,N_17835);
or U22126 (N_22126,N_17987,N_18062);
nor U22127 (N_22127,N_18897,N_19932);
or U22128 (N_22128,N_18781,N_19472);
and U22129 (N_22129,N_18827,N_19897);
nor U22130 (N_22130,N_18958,N_19600);
or U22131 (N_22131,N_18773,N_18589);
nand U22132 (N_22132,N_18092,N_19356);
nand U22133 (N_22133,N_19258,N_19761);
and U22134 (N_22134,N_19739,N_18999);
and U22135 (N_22135,N_19439,N_18123);
nand U22136 (N_22136,N_19553,N_18028);
and U22137 (N_22137,N_18192,N_18891);
and U22138 (N_22138,N_17870,N_18286);
nor U22139 (N_22139,N_18873,N_19457);
nand U22140 (N_22140,N_18271,N_19331);
or U22141 (N_22141,N_19094,N_19444);
or U22142 (N_22142,N_19700,N_18496);
nand U22143 (N_22143,N_19031,N_19142);
nand U22144 (N_22144,N_19833,N_19715);
nor U22145 (N_22145,N_19261,N_18694);
or U22146 (N_22146,N_17594,N_19947);
nand U22147 (N_22147,N_18258,N_17739);
nand U22148 (N_22148,N_18042,N_19795);
or U22149 (N_22149,N_17839,N_19113);
and U22150 (N_22150,N_17587,N_18531);
nand U22151 (N_22151,N_19072,N_18558);
and U22152 (N_22152,N_18182,N_19111);
nand U22153 (N_22153,N_19390,N_18681);
nor U22154 (N_22154,N_19452,N_19428);
and U22155 (N_22155,N_19262,N_18373);
and U22156 (N_22156,N_18553,N_18681);
nand U22157 (N_22157,N_18681,N_19375);
or U22158 (N_22158,N_17808,N_18159);
nand U22159 (N_22159,N_18756,N_18332);
nor U22160 (N_22160,N_18669,N_17573);
nand U22161 (N_22161,N_19285,N_19421);
or U22162 (N_22162,N_19334,N_19189);
or U22163 (N_22163,N_18478,N_18707);
nand U22164 (N_22164,N_19649,N_19516);
and U22165 (N_22165,N_18156,N_19331);
and U22166 (N_22166,N_17817,N_17625);
or U22167 (N_22167,N_18650,N_17706);
and U22168 (N_22168,N_17657,N_18479);
or U22169 (N_22169,N_19623,N_18351);
and U22170 (N_22170,N_18735,N_17838);
nand U22171 (N_22171,N_19267,N_19379);
nand U22172 (N_22172,N_18861,N_19642);
and U22173 (N_22173,N_19882,N_19626);
nor U22174 (N_22174,N_19602,N_19912);
nor U22175 (N_22175,N_19138,N_17533);
or U22176 (N_22176,N_19688,N_17753);
nor U22177 (N_22177,N_19042,N_19542);
or U22178 (N_22178,N_18439,N_17761);
or U22179 (N_22179,N_19304,N_18763);
or U22180 (N_22180,N_19659,N_18918);
or U22181 (N_22181,N_19901,N_19708);
nand U22182 (N_22182,N_19123,N_17598);
and U22183 (N_22183,N_19269,N_19810);
and U22184 (N_22184,N_17870,N_18535);
nand U22185 (N_22185,N_19072,N_17644);
nor U22186 (N_22186,N_18342,N_18593);
or U22187 (N_22187,N_18121,N_18985);
or U22188 (N_22188,N_19571,N_19185);
or U22189 (N_22189,N_17676,N_19839);
nor U22190 (N_22190,N_18264,N_17518);
nor U22191 (N_22191,N_18834,N_18647);
or U22192 (N_22192,N_18137,N_17722);
and U22193 (N_22193,N_18474,N_18292);
nand U22194 (N_22194,N_19848,N_19602);
nand U22195 (N_22195,N_19107,N_18209);
nand U22196 (N_22196,N_19023,N_17669);
and U22197 (N_22197,N_19304,N_19546);
and U22198 (N_22198,N_18109,N_18968);
nand U22199 (N_22199,N_19007,N_17953);
nor U22200 (N_22200,N_17788,N_18130);
nand U22201 (N_22201,N_19874,N_18265);
and U22202 (N_22202,N_19869,N_19473);
or U22203 (N_22203,N_19278,N_19115);
nor U22204 (N_22204,N_18824,N_17829);
nand U22205 (N_22205,N_19600,N_17548);
nand U22206 (N_22206,N_18858,N_19978);
and U22207 (N_22207,N_19753,N_19602);
or U22208 (N_22208,N_18937,N_18135);
or U22209 (N_22209,N_17881,N_18114);
or U22210 (N_22210,N_19402,N_18178);
nand U22211 (N_22211,N_19269,N_19308);
and U22212 (N_22212,N_17503,N_19294);
nor U22213 (N_22213,N_17538,N_18838);
and U22214 (N_22214,N_18832,N_19161);
nor U22215 (N_22215,N_19225,N_18088);
nand U22216 (N_22216,N_18704,N_18726);
nor U22217 (N_22217,N_18800,N_17941);
nor U22218 (N_22218,N_19280,N_18937);
nor U22219 (N_22219,N_17977,N_18309);
xor U22220 (N_22220,N_17685,N_19433);
and U22221 (N_22221,N_18611,N_19629);
or U22222 (N_22222,N_19994,N_18307);
and U22223 (N_22223,N_19075,N_19993);
nand U22224 (N_22224,N_18183,N_18325);
nand U22225 (N_22225,N_19654,N_19582);
nand U22226 (N_22226,N_19122,N_18427);
nor U22227 (N_22227,N_19708,N_18451);
and U22228 (N_22228,N_19441,N_18038);
or U22229 (N_22229,N_18774,N_18347);
nand U22230 (N_22230,N_17508,N_18907);
and U22231 (N_22231,N_17720,N_18207);
and U22232 (N_22232,N_17782,N_19798);
nor U22233 (N_22233,N_17807,N_19779);
or U22234 (N_22234,N_19162,N_17598);
or U22235 (N_22235,N_19102,N_18207);
nor U22236 (N_22236,N_19480,N_17778);
nor U22237 (N_22237,N_17989,N_19764);
xnor U22238 (N_22238,N_19013,N_19285);
and U22239 (N_22239,N_18143,N_18038);
and U22240 (N_22240,N_18344,N_18263);
nor U22241 (N_22241,N_17926,N_19600);
or U22242 (N_22242,N_19796,N_18229);
nor U22243 (N_22243,N_18349,N_19706);
nor U22244 (N_22244,N_19896,N_17786);
nand U22245 (N_22245,N_19550,N_17989);
or U22246 (N_22246,N_17806,N_18812);
and U22247 (N_22247,N_17752,N_18578);
and U22248 (N_22248,N_18567,N_18264);
or U22249 (N_22249,N_18950,N_18632);
nand U22250 (N_22250,N_19630,N_19200);
and U22251 (N_22251,N_19292,N_18233);
nor U22252 (N_22252,N_19725,N_18205);
nand U22253 (N_22253,N_18217,N_17660);
nor U22254 (N_22254,N_18213,N_19722);
nand U22255 (N_22255,N_17778,N_19272);
or U22256 (N_22256,N_19627,N_18435);
nor U22257 (N_22257,N_18874,N_19289);
and U22258 (N_22258,N_19027,N_17769);
nand U22259 (N_22259,N_18693,N_19779);
and U22260 (N_22260,N_19655,N_19053);
and U22261 (N_22261,N_17616,N_19035);
nand U22262 (N_22262,N_18175,N_18121);
nor U22263 (N_22263,N_18823,N_19244);
and U22264 (N_22264,N_17832,N_18078);
and U22265 (N_22265,N_19802,N_18872);
and U22266 (N_22266,N_19460,N_19320);
nor U22267 (N_22267,N_17551,N_18165);
nor U22268 (N_22268,N_19211,N_18149);
or U22269 (N_22269,N_18195,N_18885);
nand U22270 (N_22270,N_18221,N_19471);
and U22271 (N_22271,N_19151,N_18050);
or U22272 (N_22272,N_17572,N_17918);
nand U22273 (N_22273,N_18537,N_19072);
nor U22274 (N_22274,N_17649,N_18527);
nand U22275 (N_22275,N_19254,N_19341);
and U22276 (N_22276,N_17558,N_17855);
and U22277 (N_22277,N_19051,N_19794);
nand U22278 (N_22278,N_19849,N_17855);
or U22279 (N_22279,N_17543,N_17903);
nand U22280 (N_22280,N_18954,N_17821);
nand U22281 (N_22281,N_19084,N_19010);
or U22282 (N_22282,N_18665,N_19908);
nor U22283 (N_22283,N_18929,N_19269);
nor U22284 (N_22284,N_17512,N_18013);
and U22285 (N_22285,N_17979,N_19562);
nor U22286 (N_22286,N_18606,N_18633);
or U22287 (N_22287,N_17660,N_18524);
or U22288 (N_22288,N_18633,N_19986);
or U22289 (N_22289,N_19297,N_18705);
nor U22290 (N_22290,N_19592,N_17580);
and U22291 (N_22291,N_18923,N_19934);
nand U22292 (N_22292,N_17820,N_18530);
and U22293 (N_22293,N_18040,N_18148);
nor U22294 (N_22294,N_19147,N_19064);
nor U22295 (N_22295,N_19978,N_18153);
nand U22296 (N_22296,N_18043,N_19619);
and U22297 (N_22297,N_18374,N_18906);
nand U22298 (N_22298,N_19911,N_17768);
and U22299 (N_22299,N_17947,N_19926);
nand U22300 (N_22300,N_17862,N_19058);
and U22301 (N_22301,N_18768,N_18191);
nor U22302 (N_22302,N_18956,N_17563);
or U22303 (N_22303,N_18954,N_17907);
nor U22304 (N_22304,N_19881,N_17998);
and U22305 (N_22305,N_18227,N_18542);
or U22306 (N_22306,N_19602,N_18279);
nor U22307 (N_22307,N_18903,N_17805);
nand U22308 (N_22308,N_18594,N_18079);
and U22309 (N_22309,N_18264,N_19026);
nand U22310 (N_22310,N_19029,N_19114);
or U22311 (N_22311,N_18553,N_17512);
nand U22312 (N_22312,N_18708,N_19443);
nand U22313 (N_22313,N_19322,N_19437);
nand U22314 (N_22314,N_18575,N_18003);
or U22315 (N_22315,N_19223,N_19366);
or U22316 (N_22316,N_19511,N_19203);
and U22317 (N_22317,N_19485,N_19555);
or U22318 (N_22318,N_17756,N_19593);
nor U22319 (N_22319,N_19171,N_18463);
nand U22320 (N_22320,N_19900,N_19475);
nor U22321 (N_22321,N_18981,N_18872);
nand U22322 (N_22322,N_19640,N_17908);
or U22323 (N_22323,N_18498,N_19108);
nor U22324 (N_22324,N_18008,N_19368);
nand U22325 (N_22325,N_18614,N_19938);
or U22326 (N_22326,N_18330,N_18981);
nor U22327 (N_22327,N_18773,N_18161);
and U22328 (N_22328,N_19976,N_18176);
or U22329 (N_22329,N_18036,N_17847);
nand U22330 (N_22330,N_19832,N_17916);
nor U22331 (N_22331,N_19084,N_19658);
and U22332 (N_22332,N_18031,N_19288);
or U22333 (N_22333,N_18003,N_18890);
nor U22334 (N_22334,N_17903,N_19214);
nand U22335 (N_22335,N_18111,N_19183);
and U22336 (N_22336,N_17788,N_19526);
and U22337 (N_22337,N_18063,N_19538);
and U22338 (N_22338,N_18591,N_18415);
nor U22339 (N_22339,N_19381,N_17776);
xnor U22340 (N_22340,N_17591,N_18088);
nand U22341 (N_22341,N_17960,N_18778);
nor U22342 (N_22342,N_18926,N_18919);
and U22343 (N_22343,N_17966,N_17776);
nand U22344 (N_22344,N_18345,N_19594);
nor U22345 (N_22345,N_17603,N_19792);
or U22346 (N_22346,N_18242,N_18993);
nand U22347 (N_22347,N_19976,N_17557);
and U22348 (N_22348,N_18078,N_19925);
or U22349 (N_22349,N_19984,N_19979);
xor U22350 (N_22350,N_18464,N_18403);
nor U22351 (N_22351,N_17603,N_19422);
nand U22352 (N_22352,N_19832,N_18894);
nor U22353 (N_22353,N_18136,N_19901);
nand U22354 (N_22354,N_17513,N_17903);
nor U22355 (N_22355,N_19937,N_19800);
or U22356 (N_22356,N_17576,N_19268);
nor U22357 (N_22357,N_18893,N_18681);
nor U22358 (N_22358,N_18611,N_17949);
nand U22359 (N_22359,N_18940,N_19125);
and U22360 (N_22360,N_19517,N_19070);
or U22361 (N_22361,N_19107,N_17965);
or U22362 (N_22362,N_18822,N_19844);
and U22363 (N_22363,N_18930,N_18500);
nor U22364 (N_22364,N_18391,N_19557);
nand U22365 (N_22365,N_19619,N_19682);
and U22366 (N_22366,N_18052,N_17953);
or U22367 (N_22367,N_19010,N_18484);
and U22368 (N_22368,N_17766,N_19677);
nand U22369 (N_22369,N_18729,N_18155);
nand U22370 (N_22370,N_17642,N_18521);
xnor U22371 (N_22371,N_18573,N_19707);
nor U22372 (N_22372,N_18774,N_19108);
nor U22373 (N_22373,N_17972,N_19902);
nand U22374 (N_22374,N_18961,N_19909);
and U22375 (N_22375,N_19721,N_19784);
and U22376 (N_22376,N_19330,N_18421);
nor U22377 (N_22377,N_17646,N_19003);
nor U22378 (N_22378,N_18407,N_17736);
and U22379 (N_22379,N_18031,N_19392);
nor U22380 (N_22380,N_18749,N_19717);
and U22381 (N_22381,N_18030,N_19591);
nand U22382 (N_22382,N_19420,N_19606);
or U22383 (N_22383,N_18606,N_18261);
xor U22384 (N_22384,N_19112,N_19483);
nand U22385 (N_22385,N_19252,N_17950);
and U22386 (N_22386,N_17567,N_18692);
or U22387 (N_22387,N_18413,N_19256);
nand U22388 (N_22388,N_17831,N_19734);
nand U22389 (N_22389,N_17851,N_19101);
or U22390 (N_22390,N_18617,N_17860);
and U22391 (N_22391,N_18709,N_17602);
nand U22392 (N_22392,N_19685,N_19789);
nand U22393 (N_22393,N_19708,N_17578);
or U22394 (N_22394,N_19010,N_18997);
or U22395 (N_22395,N_19681,N_18133);
nand U22396 (N_22396,N_17915,N_17598);
nand U22397 (N_22397,N_19136,N_19376);
or U22398 (N_22398,N_19390,N_18168);
or U22399 (N_22399,N_17539,N_18791);
nand U22400 (N_22400,N_18642,N_18525);
nand U22401 (N_22401,N_18798,N_19267);
nor U22402 (N_22402,N_18815,N_17615);
nand U22403 (N_22403,N_19979,N_19841);
nand U22404 (N_22404,N_19576,N_19027);
nand U22405 (N_22405,N_18179,N_19179);
and U22406 (N_22406,N_18125,N_18540);
nor U22407 (N_22407,N_19069,N_18647);
nor U22408 (N_22408,N_18631,N_19519);
nor U22409 (N_22409,N_18557,N_17831);
nand U22410 (N_22410,N_18656,N_18729);
nor U22411 (N_22411,N_19176,N_18476);
nor U22412 (N_22412,N_18430,N_19639);
nor U22413 (N_22413,N_18161,N_19573);
or U22414 (N_22414,N_18213,N_18648);
and U22415 (N_22415,N_18544,N_19128);
or U22416 (N_22416,N_19226,N_19207);
nand U22417 (N_22417,N_17546,N_18769);
or U22418 (N_22418,N_18200,N_19899);
nor U22419 (N_22419,N_19088,N_19376);
nor U22420 (N_22420,N_18977,N_18877);
and U22421 (N_22421,N_17737,N_19609);
nor U22422 (N_22422,N_17884,N_18515);
or U22423 (N_22423,N_17525,N_19430);
nand U22424 (N_22424,N_17976,N_18347);
or U22425 (N_22425,N_18849,N_17620);
nor U22426 (N_22426,N_18920,N_18649);
nand U22427 (N_22427,N_19234,N_19890);
and U22428 (N_22428,N_19970,N_17638);
and U22429 (N_22429,N_17824,N_18911);
nor U22430 (N_22430,N_18209,N_19754);
nand U22431 (N_22431,N_17799,N_19055);
and U22432 (N_22432,N_19914,N_17897);
and U22433 (N_22433,N_19923,N_17837);
or U22434 (N_22434,N_19302,N_17929);
or U22435 (N_22435,N_19054,N_19385);
nand U22436 (N_22436,N_17603,N_18223);
nand U22437 (N_22437,N_17820,N_19505);
or U22438 (N_22438,N_17544,N_18228);
nand U22439 (N_22439,N_19028,N_17617);
nor U22440 (N_22440,N_17638,N_19615);
or U22441 (N_22441,N_19886,N_19240);
nor U22442 (N_22442,N_18819,N_18852);
or U22443 (N_22443,N_19596,N_18913);
nand U22444 (N_22444,N_18906,N_18754);
nor U22445 (N_22445,N_19946,N_17716);
and U22446 (N_22446,N_18897,N_18902);
nor U22447 (N_22447,N_19671,N_18315);
nand U22448 (N_22448,N_19142,N_17627);
or U22449 (N_22449,N_18668,N_17896);
nor U22450 (N_22450,N_18256,N_18696);
or U22451 (N_22451,N_19926,N_19623);
or U22452 (N_22452,N_18262,N_18086);
nor U22453 (N_22453,N_18029,N_18342);
or U22454 (N_22454,N_17565,N_17776);
xor U22455 (N_22455,N_19893,N_19359);
nand U22456 (N_22456,N_19085,N_17817);
nor U22457 (N_22457,N_18695,N_18455);
nand U22458 (N_22458,N_17681,N_18089);
nor U22459 (N_22459,N_18767,N_18060);
or U22460 (N_22460,N_19815,N_19958);
nand U22461 (N_22461,N_19972,N_18571);
or U22462 (N_22462,N_18260,N_17966);
or U22463 (N_22463,N_19778,N_17747);
nor U22464 (N_22464,N_19035,N_18315);
or U22465 (N_22465,N_18862,N_18700);
nand U22466 (N_22466,N_18420,N_19025);
and U22467 (N_22467,N_18797,N_17683);
or U22468 (N_22468,N_19926,N_18201);
and U22469 (N_22469,N_18103,N_18309);
nand U22470 (N_22470,N_17798,N_18653);
nand U22471 (N_22471,N_17822,N_17689);
and U22472 (N_22472,N_18958,N_18716);
and U22473 (N_22473,N_17843,N_19970);
nand U22474 (N_22474,N_19788,N_19520);
nor U22475 (N_22475,N_18915,N_19657);
or U22476 (N_22476,N_19756,N_17887);
or U22477 (N_22477,N_19099,N_19226);
nand U22478 (N_22478,N_19176,N_18189);
or U22479 (N_22479,N_18411,N_17883);
nor U22480 (N_22480,N_19903,N_19475);
nor U22481 (N_22481,N_17507,N_19260);
and U22482 (N_22482,N_19157,N_19245);
or U22483 (N_22483,N_19053,N_18112);
nor U22484 (N_22484,N_19364,N_17755);
nand U22485 (N_22485,N_19787,N_19140);
nand U22486 (N_22486,N_17943,N_18197);
nor U22487 (N_22487,N_19470,N_18813);
nand U22488 (N_22488,N_18928,N_18193);
nor U22489 (N_22489,N_19933,N_18673);
nand U22490 (N_22490,N_18787,N_18901);
or U22491 (N_22491,N_19745,N_17918);
or U22492 (N_22492,N_17759,N_18918);
nand U22493 (N_22493,N_19747,N_17760);
or U22494 (N_22494,N_19766,N_17992);
nand U22495 (N_22495,N_18554,N_19633);
and U22496 (N_22496,N_19313,N_18002);
and U22497 (N_22497,N_19160,N_18975);
and U22498 (N_22498,N_17890,N_18040);
or U22499 (N_22499,N_18814,N_18765);
and U22500 (N_22500,N_22263,N_22226);
and U22501 (N_22501,N_21311,N_21159);
nand U22502 (N_22502,N_22425,N_22008);
or U22503 (N_22503,N_21546,N_20449);
and U22504 (N_22504,N_21548,N_21732);
nor U22505 (N_22505,N_20756,N_21240);
nor U22506 (N_22506,N_20819,N_21230);
nand U22507 (N_22507,N_22113,N_21082);
and U22508 (N_22508,N_20336,N_21619);
nor U22509 (N_22509,N_22371,N_21487);
nor U22510 (N_22510,N_21584,N_21410);
or U22511 (N_22511,N_21865,N_20679);
nor U22512 (N_22512,N_20689,N_21258);
and U22513 (N_22513,N_21696,N_20417);
and U22514 (N_22514,N_21947,N_22122);
and U22515 (N_22515,N_22393,N_22396);
or U22516 (N_22516,N_22229,N_20140);
or U22517 (N_22517,N_21892,N_21228);
nor U22518 (N_22518,N_22088,N_21201);
or U22519 (N_22519,N_20943,N_22168);
and U22520 (N_22520,N_21436,N_21925);
nand U22521 (N_22521,N_20793,N_22043);
nand U22522 (N_22522,N_21362,N_20419);
and U22523 (N_22523,N_20164,N_21848);
nand U22524 (N_22524,N_21090,N_21132);
nor U22525 (N_22525,N_22038,N_22417);
nor U22526 (N_22526,N_22323,N_20452);
nand U22527 (N_22527,N_21708,N_20080);
and U22528 (N_22528,N_22055,N_21611);
nor U22529 (N_22529,N_20945,N_21941);
nand U22530 (N_22530,N_20811,N_21239);
and U22531 (N_22531,N_22162,N_20127);
xnor U22532 (N_22532,N_20940,N_20575);
or U22533 (N_22533,N_20663,N_21167);
or U22534 (N_22534,N_20493,N_21828);
and U22535 (N_22535,N_22490,N_21023);
nand U22536 (N_22536,N_20055,N_20720);
nand U22537 (N_22537,N_20172,N_21782);
or U22538 (N_22538,N_20455,N_22000);
nand U22539 (N_22539,N_21525,N_20406);
and U22540 (N_22540,N_21147,N_20602);
or U22541 (N_22541,N_20077,N_20938);
nand U22542 (N_22542,N_21886,N_20827);
and U22543 (N_22543,N_20657,N_20246);
and U22544 (N_22544,N_21571,N_21531);
and U22545 (N_22545,N_21823,N_20537);
nand U22546 (N_22546,N_21615,N_20622);
xor U22547 (N_22547,N_21261,N_21797);
and U22548 (N_22548,N_20761,N_22197);
or U22549 (N_22549,N_20754,N_21118);
or U22550 (N_22550,N_21687,N_21538);
or U22551 (N_22551,N_20571,N_20021);
and U22552 (N_22552,N_20705,N_21363);
and U22553 (N_22553,N_21209,N_21432);
or U22554 (N_22554,N_20374,N_20932);
nand U22555 (N_22555,N_20195,N_21857);
nand U22556 (N_22556,N_21924,N_20381);
and U22557 (N_22557,N_22296,N_20005);
and U22558 (N_22558,N_21214,N_20597);
nand U22559 (N_22559,N_22165,N_21177);
and U22560 (N_22560,N_22073,N_20105);
and U22561 (N_22561,N_22030,N_20652);
nor U22562 (N_22562,N_22255,N_22437);
nor U22563 (N_22563,N_22138,N_20111);
nand U22564 (N_22564,N_20759,N_21497);
and U22565 (N_22565,N_20796,N_20368);
or U22566 (N_22566,N_20716,N_20881);
and U22567 (N_22567,N_21370,N_21256);
or U22568 (N_22568,N_20250,N_21157);
or U22569 (N_22569,N_22488,N_20068);
nand U22570 (N_22570,N_20821,N_21065);
nor U22571 (N_22571,N_21578,N_22314);
nor U22572 (N_22572,N_22014,N_20697);
nand U22573 (N_22573,N_21437,N_21547);
and U22574 (N_22574,N_20243,N_22140);
and U22575 (N_22575,N_21260,N_21472);
nor U22576 (N_22576,N_22430,N_20865);
nand U22577 (N_22577,N_20890,N_21383);
or U22578 (N_22578,N_21073,N_22114);
and U22579 (N_22579,N_21496,N_21698);
nand U22580 (N_22580,N_20109,N_22006);
nand U22581 (N_22581,N_21489,N_21255);
and U22582 (N_22582,N_20792,N_20364);
nand U22583 (N_22583,N_21229,N_21701);
or U22584 (N_22584,N_22119,N_21544);
nand U22585 (N_22585,N_22147,N_21286);
xnor U22586 (N_22586,N_20560,N_20453);
nor U22587 (N_22587,N_20191,N_20846);
and U22588 (N_22588,N_21169,N_21498);
and U22589 (N_22589,N_20825,N_20334);
nand U22590 (N_22590,N_21481,N_21406);
nand U22591 (N_22591,N_21816,N_20545);
xor U22592 (N_22592,N_20682,N_21199);
or U22593 (N_22593,N_20201,N_21354);
and U22594 (N_22594,N_20040,N_22280);
and U22595 (N_22595,N_20313,N_21815);
nor U22596 (N_22596,N_21694,N_21749);
nand U22597 (N_22597,N_21098,N_20123);
nor U22598 (N_22598,N_21898,N_21558);
nor U22599 (N_22599,N_22325,N_20902);
or U22600 (N_22600,N_21478,N_20516);
and U22601 (N_22601,N_21306,N_21699);
nor U22602 (N_22602,N_20808,N_20726);
nor U22603 (N_22603,N_21665,N_21689);
or U22604 (N_22604,N_21096,N_22341);
nand U22605 (N_22605,N_21483,N_21474);
nand U22606 (N_22606,N_22268,N_21996);
or U22607 (N_22607,N_20521,N_21453);
or U22608 (N_22608,N_20408,N_21355);
or U22609 (N_22609,N_20850,N_21331);
or U22610 (N_22610,N_21566,N_21770);
or U22611 (N_22611,N_21289,N_22290);
and U22612 (N_22612,N_21500,N_20060);
nor U22613 (N_22613,N_22368,N_21248);
nand U22614 (N_22614,N_22466,N_21019);
or U22615 (N_22615,N_20971,N_22433);
nor U22616 (N_22616,N_21275,N_20215);
and U22617 (N_22617,N_22460,N_22481);
and U22618 (N_22618,N_20658,N_20848);
or U22619 (N_22619,N_21024,N_21549);
and U22620 (N_22620,N_20703,N_22413);
xnor U22621 (N_22621,N_20376,N_20511);
or U22622 (N_22622,N_22126,N_20740);
and U22623 (N_22623,N_21902,N_20183);
nand U22624 (N_22624,N_22192,N_21590);
and U22625 (N_22625,N_21008,N_20310);
nand U22626 (N_22626,N_21322,N_20042);
nand U22627 (N_22627,N_20024,N_21787);
nand U22628 (N_22628,N_20931,N_21655);
or U22629 (N_22629,N_21780,N_20712);
or U22630 (N_22630,N_20169,N_21644);
and U22631 (N_22631,N_20507,N_22007);
and U22632 (N_22632,N_20648,N_21343);
or U22633 (N_22633,N_20803,N_21979);
nand U22634 (N_22634,N_20830,N_21802);
and U22635 (N_22635,N_20016,N_20446);
or U22636 (N_22636,N_22467,N_21287);
nand U22637 (N_22637,N_21541,N_20157);
nand U22638 (N_22638,N_20676,N_22064);
nand U22639 (N_22639,N_20952,N_20563);
nand U22640 (N_22640,N_21397,N_20221);
nor U22641 (N_22641,N_22306,N_20096);
or U22642 (N_22642,N_20866,N_21367);
or U22643 (N_22643,N_20829,N_20568);
or U22644 (N_22644,N_22106,N_20581);
nand U22645 (N_22645,N_21299,N_21969);
or U22646 (N_22646,N_20908,N_20847);
or U22647 (N_22647,N_21338,N_20822);
or U22648 (N_22648,N_21326,N_20473);
or U22649 (N_22649,N_20779,N_21845);
or U22650 (N_22650,N_21217,N_21552);
and U22651 (N_22651,N_21904,N_21409);
or U22652 (N_22652,N_21658,N_21743);
nor U22653 (N_22653,N_20503,N_22358);
and U22654 (N_22654,N_21234,N_21637);
and U22655 (N_22655,N_21262,N_21804);
and U22656 (N_22656,N_21746,N_22435);
nand U22657 (N_22657,N_22065,N_21106);
and U22658 (N_22658,N_21404,N_22241);
nor U22659 (N_22659,N_20724,N_21358);
or U22660 (N_22660,N_21585,N_22427);
nand U22661 (N_22661,N_20423,N_22407);
and U22662 (N_22662,N_20693,N_21029);
nor U22663 (N_22663,N_21610,N_22134);
nor U22664 (N_22664,N_21955,N_21891);
nand U22665 (N_22665,N_20818,N_21994);
nand U22666 (N_22666,N_20506,N_22482);
nand U22667 (N_22667,N_21309,N_21622);
nor U22668 (N_22668,N_21020,N_21282);
and U22669 (N_22669,N_22209,N_20284);
and U22670 (N_22670,N_20546,N_20889);
nor U22671 (N_22671,N_21545,N_21194);
and U22672 (N_22672,N_22201,N_20566);
or U22673 (N_22673,N_21009,N_20324);
nor U22674 (N_22674,N_20441,N_20135);
xor U22675 (N_22675,N_20508,N_21308);
and U22676 (N_22676,N_20861,N_21168);
nor U22677 (N_22677,N_20162,N_21401);
nor U22678 (N_22678,N_21920,N_20177);
or U22679 (N_22679,N_22117,N_21012);
and U22680 (N_22680,N_20986,N_20667);
and U22681 (N_22681,N_21219,N_20458);
or U22682 (N_22682,N_21965,N_20262);
nand U22683 (N_22683,N_21120,N_21321);
nor U22684 (N_22684,N_21928,N_20628);
nand U22685 (N_22685,N_21606,N_20029);
and U22686 (N_22686,N_22356,N_20443);
nor U22687 (N_22687,N_22269,N_21860);
or U22688 (N_22688,N_20450,N_20460);
nand U22689 (N_22689,N_21609,N_21036);
and U22690 (N_22690,N_21963,N_22077);
nor U22691 (N_22691,N_21115,N_20263);
nor U22692 (N_22692,N_21893,N_21442);
or U22693 (N_22693,N_21257,N_20231);
nor U22694 (N_22694,N_20949,N_20348);
nand U22695 (N_22695,N_21390,N_21136);
nand U22696 (N_22696,N_21433,N_22003);
nor U22697 (N_22697,N_20681,N_22054);
nand U22698 (N_22698,N_22202,N_20817);
nor U22699 (N_22699,N_20744,N_20130);
nor U22700 (N_22700,N_20100,N_20468);
nand U22701 (N_22701,N_21706,N_20565);
xor U22702 (N_22702,N_21456,N_20015);
nand U22703 (N_22703,N_20656,N_20690);
and U22704 (N_22704,N_22087,N_21420);
nor U22705 (N_22705,N_21464,N_21573);
nor U22706 (N_22706,N_20337,N_21365);
or U22707 (N_22707,N_20812,N_21883);
or U22708 (N_22708,N_20256,N_21919);
and U22709 (N_22709,N_22431,N_20207);
or U22710 (N_22710,N_20107,N_20877);
nand U22711 (N_22711,N_20240,N_22342);
and U22712 (N_22712,N_20139,N_21600);
or U22713 (N_22713,N_22136,N_21441);
nand U22714 (N_22714,N_22385,N_21164);
nand U22715 (N_22715,N_21897,N_20067);
nor U22716 (N_22716,N_22154,N_20646);
and U22717 (N_22717,N_22419,N_21274);
or U22718 (N_22718,N_21810,N_20594);
nand U22719 (N_22719,N_20849,N_21128);
or U22720 (N_22720,N_22259,N_20126);
nor U22721 (N_22721,N_22072,N_20141);
or U22722 (N_22722,N_22124,N_20110);
nor U22723 (N_22723,N_21907,N_21182);
xor U22724 (N_22724,N_21844,N_20739);
or U22725 (N_22725,N_22182,N_22352);
nand U22726 (N_22726,N_21447,N_22232);
nand U22727 (N_22727,N_20244,N_21055);
or U22728 (N_22728,N_20317,N_21723);
or U22729 (N_22729,N_22053,N_22378);
nand U22730 (N_22730,N_22292,N_22452);
and U22731 (N_22731,N_21779,N_20813);
nor U22732 (N_22732,N_21466,N_20721);
or U22733 (N_22733,N_20996,N_20403);
or U22734 (N_22734,N_20731,N_20969);
or U22735 (N_22735,N_20483,N_20580);
and U22736 (N_22736,N_21396,N_20416);
or U22737 (N_22737,N_20979,N_20843);
and U22738 (N_22738,N_22468,N_20367);
or U22739 (N_22739,N_20853,N_20878);
nand U22740 (N_22740,N_22019,N_21042);
nand U22741 (N_22741,N_21330,N_22079);
nor U22742 (N_22742,N_22102,N_21625);
nand U22743 (N_22743,N_22455,N_22370);
and U22744 (N_22744,N_20644,N_22061);
or U22745 (N_22745,N_22223,N_21051);
or U22746 (N_22746,N_22098,N_21097);
nor U22747 (N_22747,N_21430,N_21601);
nand U22748 (N_22748,N_22066,N_20194);
nor U22749 (N_22749,N_20289,N_22476);
or U22750 (N_22750,N_20586,N_20701);
nand U22751 (N_22751,N_21943,N_22274);
or U22752 (N_22752,N_21266,N_22365);
or U22753 (N_22753,N_21825,N_21849);
nand U22754 (N_22754,N_20467,N_20729);
or U22755 (N_22755,N_22367,N_20610);
nand U22756 (N_22756,N_22277,N_21236);
or U22757 (N_22757,N_21554,N_22236);
and U22758 (N_22758,N_21081,N_21197);
nand U22759 (N_22759,N_22028,N_21369);
or U22760 (N_22760,N_20944,N_20227);
nor U22761 (N_22761,N_22057,N_21010);
nor U22762 (N_22762,N_21163,N_20746);
nand U22763 (N_22763,N_22491,N_22278);
nand U22764 (N_22764,N_20218,N_21711);
nand U22765 (N_22765,N_20688,N_21649);
nand U22766 (N_22766,N_21948,N_21681);
or U22767 (N_22767,N_20420,N_21087);
or U22768 (N_22768,N_20014,N_21707);
or U22769 (N_22769,N_20909,N_21833);
or U22770 (N_22770,N_21412,N_20981);
nor U22771 (N_22771,N_21271,N_22382);
nand U22772 (N_22772,N_21543,N_21461);
and U22773 (N_22773,N_20736,N_20444);
nand U22774 (N_22774,N_21469,N_21284);
xor U22775 (N_22775,N_21068,N_21334);
or U22776 (N_22776,N_21937,N_21421);
and U22777 (N_22777,N_21517,N_21524);
nor U22778 (N_22778,N_21374,N_21423);
and U22779 (N_22779,N_21613,N_21105);
or U22780 (N_22780,N_20540,N_20894);
or U22781 (N_22781,N_22373,N_21521);
nor U22782 (N_22782,N_21672,N_20457);
nor U22783 (N_22783,N_21803,N_20327);
nor U22784 (N_22784,N_21853,N_21734);
or U22785 (N_22785,N_20903,N_21705);
nand U22786 (N_22786,N_22027,N_22004);
nor U22787 (N_22787,N_21726,N_21424);
nand U22788 (N_22788,N_20750,N_20200);
nand U22789 (N_22789,N_20926,N_20351);
and U22790 (N_22790,N_20344,N_20907);
nor U22791 (N_22791,N_20155,N_20053);
and U22792 (N_22792,N_20501,N_20412);
nor U22793 (N_22793,N_21301,N_22118);
or U22794 (N_22794,N_22123,N_21627);
nor U22795 (N_22795,N_20091,N_22010);
or U22796 (N_22796,N_20020,N_20895);
nor U22797 (N_22797,N_20333,N_22400);
nor U22798 (N_22798,N_20097,N_22001);
and U22799 (N_22799,N_20770,N_22258);
and U22800 (N_22800,N_20871,N_20249);
nand U22801 (N_22801,N_21434,N_22275);
and U22802 (N_22802,N_20185,N_20884);
or U22803 (N_22803,N_20113,N_20066);
or U22804 (N_22804,N_20561,N_21473);
and U22805 (N_22805,N_20255,N_21567);
nand U22806 (N_22806,N_20839,N_20767);
xnor U22807 (N_22807,N_20478,N_20046);
nand U22808 (N_22808,N_21686,N_20976);
or U22809 (N_22809,N_20003,N_21360);
nor U22810 (N_22810,N_22357,N_20612);
nor U22811 (N_22811,N_20842,N_20598);
and U22812 (N_22812,N_21504,N_20181);
nand U22813 (N_22813,N_20384,N_21302);
nor U22814 (N_22814,N_20790,N_20522);
and U22815 (N_22815,N_21104,N_21288);
or U22816 (N_22816,N_20558,N_22234);
nor U22817 (N_22817,N_21313,N_20763);
nor U22818 (N_22818,N_21427,N_22015);
or U22819 (N_22819,N_20677,N_20136);
nor U22820 (N_22820,N_21646,N_21133);
or U22821 (N_22821,N_21942,N_20772);
nand U22822 (N_22822,N_21206,N_22059);
or U22823 (N_22823,N_21911,N_20858);
or U22824 (N_22824,N_20248,N_20947);
and U22825 (N_22825,N_20574,N_22409);
and U22826 (N_22826,N_22011,N_20121);
and U22827 (N_22827,N_21344,N_20474);
or U22828 (N_22828,N_20094,N_22181);
nand U22829 (N_22829,N_20271,N_22206);
and U22830 (N_22830,N_21908,N_22375);
nand U22831 (N_22831,N_22330,N_22288);
or U22832 (N_22832,N_20439,N_21636);
and U22833 (N_22833,N_21179,N_21704);
or U22834 (N_22834,N_20623,N_20189);
and U22835 (N_22835,N_21916,N_22249);
nand U22836 (N_22836,N_20259,N_20809);
nand U22837 (N_22837,N_20859,N_22170);
or U22838 (N_22838,N_20707,N_21186);
or U22839 (N_22839,N_20421,N_20799);
nand U22840 (N_22840,N_20708,N_21913);
and U22841 (N_22841,N_20319,N_22498);
nand U22842 (N_22842,N_20553,N_21414);
or U22843 (N_22843,N_20620,N_20922);
and U22844 (N_22844,N_20448,N_20335);
and U22845 (N_22845,N_21112,N_22097);
nand U22846 (N_22846,N_20711,N_22369);
nand U22847 (N_22847,N_20192,N_22312);
nand U22848 (N_22848,N_22089,N_20974);
or U22849 (N_22849,N_21131,N_22013);
nor U22850 (N_22850,N_20175,N_20517);
nand U22851 (N_22851,N_20424,N_20983);
or U22852 (N_22852,N_21737,N_21822);
or U22853 (N_22853,N_21176,N_21030);
nand U22854 (N_22854,N_20409,N_21086);
or U22855 (N_22855,N_21091,N_21751);
or U22856 (N_22856,N_21006,N_20395);
nor U22857 (N_22857,N_20436,N_22096);
and U22858 (N_22858,N_20524,N_21259);
nand U22859 (N_22859,N_21623,N_20340);
nand U22860 (N_22860,N_20965,N_20230);
or U22861 (N_22861,N_20329,N_20975);
or U22862 (N_22862,N_22132,N_21858);
and U22863 (N_22863,N_20788,N_20445);
or U22864 (N_22864,N_21820,N_22456);
or U22865 (N_22865,N_20959,N_21912);
nor U22866 (N_22866,N_20869,N_22142);
nand U22867 (N_22867,N_22276,N_20299);
nand U22868 (N_22868,N_22345,N_20685);
nand U22869 (N_22869,N_22063,N_21038);
nand U22870 (N_22870,N_21842,N_21034);
nor U22871 (N_22871,N_21189,N_22465);
and U22872 (N_22872,N_22026,N_21570);
or U22873 (N_22873,N_21568,N_21027);
and U22874 (N_22874,N_20190,N_20519);
nor U22875 (N_22875,N_20341,N_22475);
and U22876 (N_22876,N_21675,N_20011);
and U22877 (N_22877,N_22387,N_21639);
or U22878 (N_22878,N_21642,N_20209);
nor U22879 (N_22879,N_20151,N_22494);
nor U22880 (N_22880,N_22046,N_21993);
or U22881 (N_22881,N_21516,N_22443);
nor U22882 (N_22882,N_20125,N_22076);
nand U22883 (N_22883,N_21298,N_20213);
nand U22884 (N_22884,N_21628,N_20397);
nand U22885 (N_22885,N_21475,N_22025);
nor U22886 (N_22886,N_20228,N_21031);
nand U22887 (N_22887,N_20533,N_20738);
nand U22888 (N_22888,N_22024,N_20485);
and U22889 (N_22889,N_21740,N_21754);
and U22890 (N_22890,N_20592,N_21018);
nor U22891 (N_22891,N_21867,N_20806);
or U22892 (N_22892,N_21975,N_22362);
or U22893 (N_22893,N_20325,N_20480);
nand U22894 (N_22894,N_21514,N_21297);
nor U22895 (N_22895,N_21022,N_21764);
or U22896 (N_22896,N_20290,N_21633);
or U22897 (N_22897,N_22203,N_20165);
or U22898 (N_22898,N_20856,N_22211);
and U22899 (N_22899,N_20010,N_21371);
and U22900 (N_22900,N_20518,N_20318);
nor U22901 (N_22901,N_20783,N_21184);
nand U22902 (N_22902,N_20840,N_21494);
and U22903 (N_22903,N_20224,N_20834);
nand U22904 (N_22904,N_22354,N_21515);
nor U22905 (N_22905,N_21263,N_20713);
and U22906 (N_22906,N_21805,N_20961);
nor U22907 (N_22907,N_22484,N_20810);
nor U22908 (N_22908,N_21528,N_21641);
nand U22909 (N_22909,N_22085,N_20893);
xor U22910 (N_22910,N_21922,N_21890);
nor U22911 (N_22911,N_22225,N_20860);
or U22912 (N_22912,N_20124,N_21812);
and U22913 (N_22913,N_22086,N_20321);
or U22914 (N_22914,N_20929,N_21089);
or U22915 (N_22915,N_22462,N_21368);
and U22916 (N_22916,N_20208,N_22381);
nand U22917 (N_22917,N_21763,N_20528);
and U22918 (N_22918,N_21772,N_20063);
nand U22919 (N_22919,N_20393,N_21232);
or U22920 (N_22920,N_21443,N_21620);
or U22921 (N_22921,N_20304,N_20339);
and U22922 (N_22922,N_20857,N_22439);
nand U22923 (N_22923,N_21793,N_21391);
or U22924 (N_22924,N_22398,N_20596);
nor U22925 (N_22925,N_21002,N_22247);
nand U22926 (N_22926,N_20252,N_22084);
or U22927 (N_22927,N_21603,N_20167);
and U22928 (N_22928,N_20923,N_21878);
nand U22929 (N_22929,N_20733,N_22374);
or U22930 (N_22930,N_21663,N_21088);
nor U22931 (N_22931,N_20674,N_20489);
nand U22932 (N_22932,N_21250,N_20999);
nor U22933 (N_22933,N_22295,N_20615);
nand U22934 (N_22934,N_20088,N_20780);
nor U22935 (N_22935,N_21114,N_20650);
nor U22936 (N_22936,N_20116,N_20178);
nand U22937 (N_22937,N_22451,N_22218);
or U22938 (N_22938,N_21332,N_20163);
and U22939 (N_22939,N_20129,N_22036);
or U22940 (N_22940,N_21831,N_20358);
nor U22941 (N_22941,N_21945,N_22472);
and U22942 (N_22942,N_20548,N_21551);
xor U22943 (N_22943,N_22188,N_21231);
and U22944 (N_22944,N_22399,N_22405);
and U22945 (N_22945,N_20216,N_20146);
and U22946 (N_22946,N_20757,N_22320);
nor U22947 (N_22947,N_20862,N_21621);
nand U22948 (N_22948,N_22442,N_20948);
nand U22949 (N_22949,N_21691,N_21914);
nand U22950 (N_22950,N_21951,N_21617);
nand U22951 (N_22951,N_20970,N_20653);
and U22952 (N_22952,N_20312,N_22331);
and U22953 (N_22953,N_20437,N_21565);
nor U22954 (N_22954,N_20741,N_22139);
nor U22955 (N_22955,N_20914,N_21773);
and U22956 (N_22956,N_22023,N_22155);
and U22957 (N_22957,N_21191,N_21821);
nand U22958 (N_22958,N_21973,N_21265);
or U22959 (N_22959,N_21645,N_20702);
and U22960 (N_22960,N_22291,N_20265);
nor U22961 (N_22961,N_20211,N_20638);
nand U22962 (N_22962,N_21840,N_21539);
nand U22963 (N_22963,N_21003,N_21300);
nand U22964 (N_22964,N_21653,N_20845);
nor U22965 (N_22965,N_21974,N_22128);
and U22966 (N_22966,N_20589,N_20203);
nand U22967 (N_22967,N_20085,N_21340);
nor U22968 (N_22968,N_20936,N_22366);
nand U22969 (N_22969,N_20634,N_22480);
and U22970 (N_22970,N_22394,N_21053);
or U22971 (N_22971,N_20535,N_20432);
and U22972 (N_22972,N_21195,N_21079);
nor U22973 (N_22973,N_20306,N_21569);
nor U22974 (N_22974,N_21372,N_20018);
and U22975 (N_22975,N_21353,N_20924);
and U22976 (N_22976,N_21192,N_22340);
and U22977 (N_22977,N_21956,N_21083);
or U22978 (N_22978,N_20798,N_21151);
and U22979 (N_22979,N_20916,N_22304);
nor U22980 (N_22980,N_20766,N_21015);
nor U22981 (N_22981,N_20104,N_22108);
or U22982 (N_22982,N_22099,N_20009);
xnor U22983 (N_22983,N_21373,N_20267);
or U22984 (N_22984,N_20198,N_22347);
or U22985 (N_22985,N_22219,N_21238);
nor U22986 (N_22986,N_20082,N_20268);
nand U22987 (N_22987,N_21638,N_20315);
nor U22988 (N_22988,N_20987,N_20785);
nor U22989 (N_22989,N_20876,N_20314);
nand U22990 (N_22990,N_21839,N_21760);
and U22991 (N_22991,N_22095,N_20283);
or U22992 (N_22992,N_22074,N_20300);
or U22993 (N_22993,N_21519,N_21064);
and U22994 (N_22994,N_20606,N_21455);
nor U22995 (N_22995,N_21341,N_20138);
and U22996 (N_22996,N_21060,N_20214);
and U22997 (N_22997,N_20673,N_20044);
nand U22998 (N_22998,N_20173,N_20301);
nor U22999 (N_22999,N_22176,N_21605);
nor U23000 (N_23000,N_21594,N_21431);
nand U23001 (N_23001,N_22260,N_20980);
nand U23002 (N_23002,N_21440,N_20715);
or U23003 (N_23003,N_20826,N_21438);
nor U23004 (N_23004,N_20150,N_20614);
or U23005 (N_23005,N_21210,N_20831);
nand U23006 (N_23006,N_22309,N_22440);
and U23007 (N_23007,N_20514,N_20680);
nor U23008 (N_23008,N_21887,N_20035);
nand U23009 (N_23009,N_20418,N_20002);
or U23010 (N_23010,N_21972,N_22174);
and U23011 (N_23011,N_20611,N_22233);
or U23012 (N_23012,N_21101,N_20982);
nor U23013 (N_23013,N_20649,N_20805);
and U23014 (N_23014,N_21612,N_20801);
or U23015 (N_23015,N_21715,N_21318);
or U23016 (N_23016,N_22078,N_21211);
or U23017 (N_23017,N_20699,N_22208);
or U23018 (N_23018,N_21856,N_20905);
nand U23019 (N_23019,N_20539,N_20920);
nor U23020 (N_23020,N_20631,N_21185);
nor U23021 (N_23021,N_20219,N_22293);
nor U23022 (N_23022,N_21884,N_21540);
or U23023 (N_23023,N_20128,N_22080);
or U23024 (N_23024,N_21561,N_21119);
or U23025 (N_23025,N_22322,N_20472);
nand U23026 (N_23026,N_21767,N_22056);
nand U23027 (N_23027,N_21335,N_20059);
nand U23028 (N_23028,N_21005,N_20991);
nor U23029 (N_23029,N_21664,N_21792);
xnor U23030 (N_23030,N_20311,N_20710);
and U23031 (N_23031,N_21870,N_21624);
or U23032 (N_23032,N_20081,N_21327);
nand U23033 (N_23033,N_21033,N_21063);
nand U23034 (N_23034,N_21011,N_21968);
nand U23035 (N_23035,N_21953,N_22346);
nor U23036 (N_23036,N_20242,N_21523);
nand U23037 (N_23037,N_21932,N_21819);
and U23038 (N_23038,N_21534,N_21673);
and U23039 (N_23039,N_20771,N_22163);
nor U23040 (N_23040,N_21074,N_20885);
nand U23041 (N_23041,N_20547,N_21137);
or U23042 (N_23042,N_22483,N_20717);
nor U23043 (N_23043,N_21467,N_20919);
or U23044 (N_23044,N_21807,N_21276);
nor U23045 (N_23045,N_21451,N_22067);
nor U23046 (N_23046,N_21439,N_22121);
or U23047 (N_23047,N_21058,N_21149);
nand U23048 (N_23048,N_21283,N_20755);
or U23049 (N_23049,N_20600,N_21786);
nor U23050 (N_23050,N_21801,N_20669);
or U23051 (N_23051,N_20355,N_20133);
nand U23052 (N_23052,N_22224,N_21241);
xnor U23053 (N_23053,N_21589,N_20692);
or U23054 (N_23054,N_22446,N_21224);
or U23055 (N_23055,N_21529,N_21315);
or U23056 (N_23056,N_21762,N_21385);
and U23057 (N_23057,N_20237,N_22071);
nor U23058 (N_23058,N_22069,N_21852);
or U23059 (N_23059,N_21889,N_21425);
nand U23060 (N_23060,N_21962,N_21480);
nor U23061 (N_23061,N_21400,N_20202);
nand U23062 (N_23062,N_21868,N_21741);
or U23063 (N_23063,N_22459,N_20451);
nand U23064 (N_23064,N_20502,N_20171);
or U23065 (N_23065,N_20095,N_22495);
or U23066 (N_23066,N_21560,N_21952);
nand U23067 (N_23067,N_21290,N_22110);
nor U23068 (N_23068,N_20698,N_21862);
and U23069 (N_23069,N_21143,N_20621);
or U23070 (N_23070,N_21277,N_21346);
and U23071 (N_23071,N_22423,N_21895);
or U23072 (N_23072,N_20027,N_20512);
nand U23073 (N_23073,N_22469,N_22227);
or U23074 (N_23074,N_22426,N_20595);
and U23075 (N_23075,N_21099,N_21505);
nand U23076 (N_23076,N_20398,N_21316);
nand U23077 (N_23077,N_21971,N_22130);
nand U23078 (N_23078,N_21142,N_21317);
and U23079 (N_23079,N_20030,N_21435);
xnor U23080 (N_23080,N_20782,N_22415);
or U23081 (N_23081,N_20937,N_20353);
nand U23082 (N_23082,N_21382,N_20049);
nor U23083 (N_23083,N_22017,N_20001);
or U23084 (N_23084,N_22081,N_20365);
and U23085 (N_23085,N_22364,N_20573);
nand U23086 (N_23086,N_20307,N_21499);
nor U23087 (N_23087,N_21304,N_20605);
and U23088 (N_23088,N_20401,N_22305);
or U23089 (N_23089,N_20769,N_21669);
nor U23090 (N_23090,N_21426,N_21196);
and U23091 (N_23091,N_20544,N_20977);
or U23092 (N_23092,N_20686,N_22094);
nand U23093 (N_23093,N_21678,N_21513);
nor U23094 (N_23094,N_21864,N_20781);
nand U23095 (N_23095,N_21449,N_20402);
and U23096 (N_23096,N_21748,N_20072);
and U23097 (N_23097,N_21724,N_22169);
nand U23098 (N_23098,N_21285,N_22457);
and U23099 (N_23099,N_20156,N_20273);
nand U23100 (N_23100,N_20559,N_20051);
nand U23101 (N_23101,N_20748,N_20582);
nand U23102 (N_23102,N_22416,N_22020);
nand U23103 (N_23103,N_21900,N_21959);
and U23104 (N_23104,N_21312,N_21781);
or U23105 (N_23105,N_20466,N_20554);
and U23106 (N_23106,N_22334,N_20394);
nand U23107 (N_23107,N_20238,N_21488);
and U23108 (N_23108,N_22104,N_21491);
nor U23109 (N_23109,N_20700,N_21398);
and U23110 (N_23110,N_20170,N_20400);
nand U23111 (N_23111,N_22436,N_20260);
or U23112 (N_23112,N_21542,N_20967);
nor U23113 (N_23113,N_20297,N_20978);
nand U23114 (N_23114,N_21808,N_20050);
nand U23115 (N_23115,N_22270,N_22049);
and U23116 (N_23116,N_20490,N_21931);
or U23117 (N_23117,N_22153,N_20593);
nor U23118 (N_23118,N_21486,N_20637);
nor U23119 (N_23119,N_20430,N_20671);
nand U23120 (N_23120,N_21084,N_21124);
or U23121 (N_23121,N_21061,N_20863);
nor U23122 (N_23122,N_20281,N_22105);
or U23123 (N_23123,N_21991,N_21918);
or U23124 (N_23124,N_21555,N_21927);
or U23125 (N_23125,N_20617,N_22199);
or U23126 (N_23126,N_21180,N_21154);
nor U23127 (N_23127,N_21938,N_20052);
nand U23128 (N_23128,N_21934,N_20504);
and U23129 (N_23129,N_21223,N_21685);
nand U23130 (N_23130,N_20662,N_20530);
or U23131 (N_23131,N_22207,N_20873);
and U23132 (N_23132,N_22316,N_22383);
or U23133 (N_23133,N_22133,N_21450);
or U23134 (N_23134,N_20407,N_21272);
nand U23135 (N_23135,N_22044,N_21183);
and U23136 (N_23136,N_22404,N_21647);
and U23137 (N_23137,N_21880,N_21843);
nand U23138 (N_23138,N_22496,N_21243);
or U23139 (N_23139,N_20386,N_22177);
and U23140 (N_23140,N_20017,N_21752);
or U23141 (N_23141,N_21307,N_22264);
nand U23142 (N_23142,N_20352,N_20405);
nand U23143 (N_23143,N_21817,N_20426);
nand U23144 (N_23144,N_22411,N_21377);
or U23145 (N_23145,N_22324,N_21745);
nor U23146 (N_23146,N_21403,N_20206);
and U23147 (N_23147,N_21459,N_22235);
or U23148 (N_23148,N_21855,N_22350);
xnor U23149 (N_23149,N_20795,N_22244);
nand U23150 (N_23150,N_20226,N_21946);
or U23151 (N_23151,N_21085,N_20901);
nor U23152 (N_23152,N_20882,N_21755);
or U23153 (N_23153,N_22172,N_21987);
and U23154 (N_23154,N_21056,N_22256);
or U23155 (N_23155,N_20481,N_20168);
nor U23156 (N_23156,N_22447,N_21742);
and U23157 (N_23157,N_21107,N_20435);
nor U23158 (N_23158,N_22198,N_21399);
or U23159 (N_23159,N_21983,N_22402);
nand U23160 (N_23160,N_21050,N_21683);
or U23161 (N_23161,N_22307,N_20347);
nand U23162 (N_23162,N_21203,N_20342);
or U23163 (N_23163,N_20910,N_20515);
or U23164 (N_23164,N_20973,N_22180);
nor U23165 (N_23165,N_20666,N_20851);
nand U23166 (N_23166,N_21725,N_20935);
nand U23167 (N_23167,N_21458,N_20531);
nor U23168 (N_23168,N_20934,N_22361);
and U23169 (N_23169,N_21493,N_21417);
nor U23170 (N_23170,N_20643,N_21126);
and U23171 (N_23171,N_21198,N_21632);
and U23172 (N_23172,N_20989,N_21445);
nand U23173 (N_23173,N_21837,N_20143);
nand U23174 (N_23174,N_22157,N_21503);
nor U23175 (N_23175,N_20205,N_21452);
and U23176 (N_23176,N_20784,N_21387);
or U23177 (N_23177,N_20388,N_21325);
nor U23178 (N_23178,N_20278,N_21045);
or U23179 (N_23179,N_22392,N_20193);
nor U23180 (N_23180,N_22294,N_20664);
or U23181 (N_23181,N_22377,N_20529);
or U23182 (N_23182,N_20870,N_22444);
or U23183 (N_23183,N_20180,N_20261);
nand U23184 (N_23184,N_22418,N_22388);
nor U23185 (N_23185,N_21882,N_22461);
and U23186 (N_23186,N_20253,N_21511);
and U23187 (N_23187,N_21593,N_20122);
or U23188 (N_23188,N_21794,N_21273);
and U23189 (N_23189,N_21877,N_21854);
or U23190 (N_23190,N_21502,N_20036);
and U23191 (N_23191,N_22485,N_20727);
nor U23192 (N_23192,N_20963,N_20641);
or U23193 (N_23193,N_22441,N_20494);
nor U23194 (N_23194,N_21170,N_20098);
and U23195 (N_23195,N_20147,N_21608);
or U23196 (N_23196,N_20158,N_20349);
nor U23197 (N_23197,N_22487,N_22363);
and U23198 (N_23198,N_20118,N_21830);
nand U23199 (N_23199,N_21001,N_21293);
or U23200 (N_23200,N_21885,N_21092);
xor U23201 (N_23201,N_21879,N_22301);
or U23202 (N_23202,N_20232,N_21140);
or U23203 (N_23203,N_20429,N_21465);
or U23204 (N_23204,N_21032,N_20387);
or U23205 (N_23205,N_20469,N_22336);
nor U23206 (N_23206,N_21654,N_21630);
nor U23207 (N_23207,N_22252,N_20745);
or U23208 (N_23208,N_21981,N_20904);
and U23209 (N_23209,N_21957,N_21629);
nor U23210 (N_23210,N_21379,N_21933);
and U23211 (N_23211,N_20758,N_21233);
or U23212 (N_23212,N_21139,N_20824);
and U23213 (N_23213,N_21949,N_20816);
nand U23214 (N_23214,N_20921,N_20026);
nor U23215 (N_23215,N_20655,N_22047);
nor U23216 (N_23216,N_20275,N_22230);
nor U23217 (N_23217,N_22389,N_21251);
and U23218 (N_23218,N_21881,N_20951);
and U23219 (N_23219,N_20350,N_20411);
nor U23220 (N_23220,N_22279,N_20102);
and U23221 (N_23221,N_21249,N_20953);
nand U23222 (N_23222,N_20968,N_20955);
nand U23223 (N_23223,N_22329,N_21408);
nor U23224 (N_23224,N_22231,N_20765);
or U23225 (N_23225,N_20120,N_20835);
or U23226 (N_23226,N_22445,N_21471);
nand U23227 (N_23227,N_21025,N_20837);
or U23228 (N_23228,N_20526,N_20078);
nor U23229 (N_23229,N_20629,N_20234);
and U23230 (N_23230,N_20061,N_20694);
nor U23231 (N_23231,N_20995,N_20000);
nand U23232 (N_23232,N_20119,N_22317);
nand U23233 (N_23233,N_21342,N_21574);
nor U23234 (N_23234,N_22173,N_21359);
nand U23235 (N_23235,N_21215,N_21677);
nand U23236 (N_23236,N_20564,N_22204);
nand U23237 (N_23237,N_20089,N_20872);
nor U23238 (N_23238,N_22332,N_21294);
nor U23239 (N_23239,N_20804,N_20532);
nand U23240 (N_23240,N_21530,N_20266);
and U23241 (N_23241,N_20294,N_20279);
and U23242 (N_23242,N_20245,N_20964);
or U23243 (N_23243,N_20499,N_21418);
and U23244 (N_23244,N_20584,N_20775);
nor U23245 (N_23245,N_20990,N_21989);
or U23246 (N_23246,N_21429,N_22300);
nor U23247 (N_23247,N_20090,N_21366);
and U23248 (N_23248,N_20389,N_21872);
xnor U23249 (N_23249,N_20251,N_21731);
nor U23250 (N_23250,N_22262,N_21832);
and U23251 (N_23251,N_20187,N_20607);
or U23252 (N_23252,N_20379,N_21329);
and U23253 (N_23253,N_20092,N_21044);
or U23254 (N_23254,N_22189,N_22179);
nor U23255 (N_23255,N_20370,N_21572);
nor U23256 (N_23256,N_22131,N_21407);
nand U23257 (N_23257,N_21468,N_21970);
or U23258 (N_23258,N_20022,N_22283);
and U23259 (N_23259,N_20627,N_22448);
nand U23260 (N_23260,N_22303,N_21495);
nor U23261 (N_23261,N_21361,N_22239);
or U23262 (N_23262,N_22009,N_20956);
and U23263 (N_23263,N_20008,N_22380);
nand U23264 (N_23264,N_20199,N_20323);
and U23265 (N_23265,N_20391,N_22171);
or U23266 (N_23266,N_22438,N_22052);
nor U23267 (N_23267,N_21591,N_20186);
and U23268 (N_23268,N_22434,N_22037);
xnor U23269 (N_23269,N_21671,N_22159);
and U23270 (N_23270,N_20985,N_20390);
nor U23271 (N_23271,N_21247,N_21905);
nand U23272 (N_23272,N_20288,N_21462);
nand U23273 (N_23273,N_20070,N_22251);
nor U23274 (N_23274,N_22175,N_21692);
or U23275 (N_23275,N_20286,N_22339);
nand U23276 (N_23276,N_21988,N_21982);
nand U23277 (N_23277,N_20383,N_21730);
or U23278 (N_23278,N_20047,N_21328);
nand U23279 (N_23279,N_21700,N_22166);
nand U23280 (N_23280,N_20645,N_20569);
nor U23281 (N_23281,N_20496,N_20960);
and U23282 (N_23282,N_21166,N_20241);
or U23283 (N_23283,N_22343,N_21292);
or U23284 (N_23284,N_20484,N_20380);
or U23285 (N_23285,N_22187,N_21047);
nand U23286 (N_23286,N_20883,N_21657);
and U23287 (N_23287,N_20425,N_21007);
nand U23288 (N_23288,N_21109,N_21990);
nor U23289 (N_23289,N_21966,N_21227);
and U23290 (N_23290,N_20159,N_21016);
nand U23291 (N_23291,N_20728,N_20075);
or U23292 (N_23292,N_20625,N_20332);
or U23293 (N_23293,N_22183,N_22298);
nand U23294 (N_23294,N_21759,N_20678);
nand U23295 (N_23295,N_21216,N_21835);
nand U23296 (N_23296,N_20103,N_20897);
nor U23297 (N_23297,N_20371,N_21077);
nor U23298 (N_23298,N_20852,N_21237);
nor U23299 (N_23299,N_20357,N_21204);
nor U23300 (N_23300,N_21798,N_20354);
nand U23301 (N_23301,N_22284,N_21757);
or U23302 (N_23302,N_21130,N_21536);
and U23303 (N_23303,N_21846,N_21618);
nand U23304 (N_23304,N_22246,N_22478);
nand U23305 (N_23305,N_22261,N_22101);
nor U23306 (N_23306,N_22286,N_22315);
or U23307 (N_23307,N_21080,N_21446);
nor U23308 (N_23308,N_22149,N_22449);
nand U23309 (N_23309,N_20776,N_21225);
or U23310 (N_23310,N_20233,N_22031);
and U23311 (N_23311,N_20101,N_20025);
or U23312 (N_23312,N_22144,N_20298);
and U23313 (N_23313,N_21037,N_20773);
nand U23314 (N_23314,N_21896,N_20555);
nor U23315 (N_23315,N_21716,N_20972);
nand U23316 (N_23316,N_20112,N_22308);
and U23317 (N_23317,N_21576,N_21894);
nor U23318 (N_23318,N_20800,N_21588);
nand U23319 (N_23319,N_20235,N_20399);
or U23320 (N_23320,N_22410,N_20557);
or U23321 (N_23321,N_21871,N_21869);
or U23322 (N_23322,N_21771,N_21604);
and U23323 (N_23323,N_20456,N_21679);
nor U23324 (N_23324,N_21796,N_21181);
nand U23325 (N_23325,N_22191,N_21643);
or U23326 (N_23326,N_20048,N_20854);
nor U23327 (N_23327,N_20647,N_20917);
nand U23328 (N_23328,N_21220,N_20326);
or U23329 (N_23329,N_20043,N_22160);
nand U23330 (N_23330,N_20742,N_21861);
nand U23331 (N_23331,N_20293,N_21656);
or U23332 (N_23332,N_20875,N_22158);
and U23333 (N_23333,N_21859,N_21936);
nand U23334 (N_23334,N_21799,N_20012);
nor U23335 (N_23335,N_21111,N_21134);
nand U23336 (N_23336,N_20217,N_21875);
nor U23337 (N_23337,N_21146,N_20604);
nand U23338 (N_23338,N_20032,N_20309);
or U23339 (N_23339,N_22091,N_20672);
or U23340 (N_23340,N_21717,N_22116);
and U23341 (N_23341,N_21939,N_20749);
or U23342 (N_23342,N_21785,N_21205);
or U23343 (N_23343,N_20148,N_20718);
or U23344 (N_23344,N_20887,N_20879);
nor U23345 (N_23345,N_20642,N_22248);
or U23346 (N_23346,N_20958,N_21776);
and U23347 (N_23347,N_21910,N_20491);
nand U23348 (N_23348,N_20372,N_21626);
nand U23349 (N_23349,N_21135,N_20639);
nand U23350 (N_23350,N_21125,N_22302);
nand U23351 (N_23351,N_22464,N_21153);
or U23352 (N_23352,N_22486,N_20520);
and U23353 (N_23353,N_21836,N_22111);
nand U23354 (N_23354,N_22338,N_20486);
nor U23355 (N_23355,N_20659,N_21270);
nor U23356 (N_23356,N_20320,N_20925);
nor U23357 (N_23357,N_21944,N_20410);
or U23358 (N_23358,N_21721,N_21336);
nand U23359 (N_23359,N_21512,N_21392);
nor U23360 (N_23360,N_20154,N_21017);
nand U23361 (N_23361,N_21769,N_21155);
and U23362 (N_23362,N_21697,N_22178);
nand U23363 (N_23363,N_20303,N_21428);
and U23364 (N_23364,N_20464,N_20099);
or U23365 (N_23365,N_21508,N_20867);
and U23366 (N_23366,N_22386,N_20844);
and U23367 (N_23367,N_22390,N_21758);
and U23368 (N_23368,N_20404,N_20142);
and U23369 (N_23369,N_20131,N_21026);
nor U23370 (N_23370,N_22022,N_20019);
nor U23371 (N_23371,N_21718,N_21661);
and U23372 (N_23372,N_22271,N_21659);
or U23373 (N_23373,N_20950,N_22406);
or U23374 (N_23374,N_21254,N_22002);
nand U23375 (N_23375,N_21533,N_20590);
and U23376 (N_23376,N_21651,N_21635);
and U23377 (N_23377,N_20006,N_20220);
nor U23378 (N_23378,N_20360,N_21800);
and U23379 (N_23379,N_21774,N_20762);
nor U23380 (N_23380,N_20461,N_22479);
or U23381 (N_23381,N_21863,N_21667);
and U23382 (N_23382,N_22215,N_21784);
and U23383 (N_23383,N_22299,N_22474);
nor U23384 (N_23384,N_21123,N_20687);
nor U23385 (N_23385,N_21094,N_22125);
xnor U23386 (N_23386,N_21122,N_22429);
nand U23387 (N_23387,N_21129,N_20463);
nand U23388 (N_23388,N_21834,N_20704);
nor U23389 (N_23389,N_21527,N_20363);
nor U23390 (N_23390,N_22266,N_20556);
nand U23391 (N_23391,N_22035,N_20459);
nor U23392 (N_23392,N_22051,N_22217);
nor U23393 (N_23393,N_20322,N_22222);
nor U23394 (N_23394,N_20369,N_21349);
nand U23395 (N_23395,N_21788,N_20087);
nand U23396 (N_23396,N_21350,N_21980);
or U23397 (N_23397,N_21103,N_21553);
nand U23398 (N_23398,N_20176,N_20064);
and U23399 (N_23399,N_20828,N_20037);
nand U23400 (N_23400,N_21506,N_20802);
or U23401 (N_23401,N_21356,N_20079);
and U23402 (N_23402,N_21518,N_22384);
or U23403 (N_23403,N_21419,N_20855);
or U23404 (N_23404,N_21648,N_21484);
nor U23405 (N_23405,N_21559,N_22422);
and U23406 (N_23406,N_22214,N_22297);
nand U23407 (N_23407,N_21100,N_20734);
nand U23408 (N_23408,N_21490,N_20747);
nand U23409 (N_23409,N_22428,N_22040);
and U23410 (N_23410,N_21977,N_21909);
nor U23411 (N_23411,N_20338,N_20254);
nor U23412 (N_23412,N_22355,N_20719);
and U23413 (N_23413,N_21244,N_22412);
or U23414 (N_23414,N_21324,N_22210);
nor U23415 (N_23415,N_21014,N_20285);
nor U23416 (N_23416,N_22470,N_20635);
nand U23417 (N_23417,N_20495,N_20505);
nor U23418 (N_23418,N_22042,N_21413);
or U23419 (N_23419,N_20295,N_22333);
or U23420 (N_23420,N_20276,N_21305);
nand U23421 (N_23421,N_21507,N_20696);
nand U23422 (N_23422,N_20777,N_20477);
nor U23423 (N_23423,N_21479,N_20892);
or U23424 (N_23424,N_20609,N_21278);
or U23425 (N_23425,N_20114,N_21454);
nor U23426 (N_23426,N_22190,N_22327);
and U23427 (N_23427,N_20542,N_20149);
or U23428 (N_23428,N_20482,N_21761);
nand U23429 (N_23429,N_20913,N_21556);
or U23430 (N_23430,N_20045,N_21950);
nor U23431 (N_23431,N_20906,N_20392);
or U23432 (N_23432,N_20161,N_21127);
nand U23433 (N_23433,N_21826,N_21386);
or U23434 (N_23434,N_22041,N_21470);
nand U23435 (N_23435,N_22242,N_20918);
nor U23436 (N_23436,N_21463,N_21818);
nor U23437 (N_23437,N_21448,N_21158);
and U23438 (N_23438,N_21888,N_21940);
and U23439 (N_23439,N_20117,N_21253);
nand U23440 (N_23440,N_21720,N_20382);
nor U23441 (N_23441,N_20270,N_22103);
and U23442 (N_23442,N_20134,N_22265);
or U23443 (N_23443,N_20626,N_20069);
and U23444 (N_23444,N_20891,N_20927);
nand U23445 (N_23445,N_20137,N_21162);
xor U23446 (N_23446,N_20838,N_22250);
nor U23447 (N_23447,N_20651,N_21174);
nor U23448 (N_23448,N_21598,N_21827);
nand U23449 (N_23449,N_21668,N_21674);
and U23450 (N_23450,N_21066,N_21188);
and U23451 (N_23451,N_21457,N_20223);
or U23452 (N_23452,N_21562,N_21915);
and U23453 (N_23453,N_22045,N_20552);
or U23454 (N_23454,N_21710,N_20670);
nand U23455 (N_23455,N_20534,N_20868);
and U23456 (N_23456,N_22070,N_22090);
or U23457 (N_23457,N_21145,N_20427);
and U23458 (N_23458,N_20613,N_21175);
nand U23459 (N_23459,N_22107,N_21733);
or U23460 (N_23460,N_20660,N_20106);
or U23461 (N_23461,N_21337,N_20510);
and U23462 (N_23462,N_22152,N_22205);
nand U23463 (N_23463,N_21476,N_22414);
or U23464 (N_23464,N_21921,N_20841);
or U23465 (N_23465,N_21713,N_20730);
nand U23466 (N_23466,N_22313,N_22360);
nor U23467 (N_23467,N_21580,N_20272);
nor U23468 (N_23468,N_22167,N_21492);
nand U23469 (N_23469,N_20084,N_20823);
nor U23470 (N_23470,N_21739,N_22353);
or U23471 (N_23471,N_20257,N_22319);
and U23472 (N_23472,N_22141,N_21116);
nor U23473 (N_23473,N_20076,N_22238);
nand U23474 (N_23474,N_21348,N_21319);
nor U23475 (N_23475,N_21670,N_20433);
nor U23476 (N_23476,N_20440,N_22237);
or U23477 (N_23477,N_21690,N_20930);
nor U23478 (N_23478,N_21178,N_21958);
or U23479 (N_23479,N_21597,N_21688);
and U23480 (N_23480,N_20362,N_21778);
nor U23481 (N_23481,N_22492,N_21703);
nand U23482 (N_23482,N_21000,N_20056);
and U23483 (N_23483,N_21395,N_21043);
and U23484 (N_23484,N_20152,N_21999);
nor U23485 (N_23485,N_20587,N_20536);
or U23486 (N_23486,N_21520,N_22109);
nand U23487 (N_23487,N_22115,N_21035);
and U23488 (N_23488,N_22083,N_22403);
or U23489 (N_23489,N_21917,N_21333);
nand U23490 (N_23490,N_21550,N_20998);
nor U23491 (N_23491,N_21695,N_21873);
or U23492 (N_23492,N_20328,N_20465);
and U23493 (N_23493,N_21193,N_20874);
or U23494 (N_23494,N_20994,N_21200);
nor U23495 (N_23495,N_21650,N_22075);
nor U23496 (N_23496,N_20471,N_20188);
nor U23497 (N_23497,N_20588,N_20331);
and U23498 (N_23498,N_20709,N_22289);
or U23499 (N_23499,N_20683,N_21213);
nor U23500 (N_23500,N_21595,N_21156);
and U23501 (N_23501,N_21121,N_21202);
nor U23502 (N_23502,N_21744,N_20007);
nand U23503 (N_23503,N_22245,N_20661);
or U23504 (N_23504,N_20305,N_21041);
and U23505 (N_23505,N_20396,N_21535);
nand U23506 (N_23506,N_20632,N_22082);
nor U23507 (N_23507,N_21736,N_20880);
nand U23508 (N_23508,N_22143,N_22408);
nand U23509 (N_23509,N_21264,N_22454);
nand U23510 (N_23510,N_22151,N_21095);
nor U23511 (N_23511,N_20296,N_21824);
or U23512 (N_23512,N_21165,N_22146);
and U23513 (N_23513,N_21575,N_20033);
nand U23514 (N_23514,N_20737,N_20576);
and U23515 (N_23515,N_21930,N_20023);
nand U23516 (N_23516,N_22050,N_21728);
or U23517 (N_23517,N_21537,N_20359);
or U23518 (N_23518,N_20236,N_20601);
nand U23519 (N_23519,N_20108,N_21783);
nor U23520 (N_23520,N_20166,N_22432);
or U23521 (N_23521,N_20414,N_20229);
and U23522 (N_23522,N_20836,N_20422);
nor U23523 (N_23523,N_20413,N_22471);
xor U23524 (N_23524,N_21389,N_20280);
nor U23525 (N_23525,N_20442,N_21906);
and U23526 (N_23526,N_22489,N_21960);
nand U23527 (N_23527,N_21738,N_21067);
nand U23528 (N_23528,N_22493,N_20665);
nand U23529 (N_23529,N_22473,N_21352);
nor U23530 (N_23530,N_22112,N_20791);
nand U23531 (N_23531,N_20086,N_20434);
nor U23532 (N_23532,N_22257,N_21161);
nor U23533 (N_23533,N_20570,N_22391);
or U23534 (N_23534,N_21268,N_22193);
nor U23535 (N_23535,N_20939,N_22137);
nor U23536 (N_23536,N_20196,N_21222);
or U23537 (N_23537,N_22326,N_20210);
and U23538 (N_23538,N_21485,N_22379);
and U23539 (N_23539,N_21314,N_20222);
or U23540 (N_23540,N_20668,N_21666);
nor U23541 (N_23541,N_21719,N_20274);
nor U23542 (N_23542,N_20438,N_21693);
nor U23543 (N_23543,N_22243,N_21347);
nor U23544 (N_23544,N_20492,N_21790);
nor U23545 (N_23545,N_21660,N_22135);
nand U23546 (N_23546,N_21985,N_22216);
nor U23547 (N_23547,N_20291,N_21267);
nand U23548 (N_23548,N_21351,N_22150);
or U23549 (N_23549,N_21381,N_20366);
and U23550 (N_23550,N_21777,N_22318);
nor U23551 (N_23551,N_22029,N_20247);
or U23552 (N_23552,N_21422,N_22282);
and U23553 (N_23553,N_20864,N_21766);
nor U23554 (N_23554,N_21411,N_20345);
nand U23555 (N_23555,N_21582,N_20551);
or U23556 (N_23556,N_20083,N_20786);
and U23557 (N_23557,N_21303,N_21416);
and U23558 (N_23558,N_21393,N_20488);
nor U23559 (N_23559,N_20578,N_20572);
and U23560 (N_23560,N_22328,N_22058);
or U23561 (N_23561,N_21402,N_20753);
nor U23562 (N_23562,N_21935,N_20225);
and U23563 (N_23563,N_20900,N_22337);
nor U23564 (N_23564,N_20993,N_21923);
nand U23565 (N_23565,N_22344,N_20912);
and U23566 (N_23566,N_20764,N_20454);
or U23567 (N_23567,N_21676,N_20509);
nand U23568 (N_23568,N_20039,N_21477);
and U23569 (N_23569,N_21150,N_21460);
nand U23570 (N_23570,N_20527,N_20538);
or U23571 (N_23571,N_21187,N_21841);
and U23572 (N_23572,N_20330,N_20984);
or U23573 (N_23573,N_20498,N_21702);
nand U23574 (N_23574,N_21607,N_21364);
and U23575 (N_23575,N_22376,N_20093);
nor U23576 (N_23576,N_20957,N_21501);
nor U23577 (N_23577,N_20691,N_20292);
and U23578 (N_23578,N_22184,N_20479);
or U23579 (N_23579,N_22185,N_21997);
nor U23580 (N_23580,N_20277,N_20184);
and U23581 (N_23581,N_20487,N_20212);
or U23582 (N_23582,N_20896,N_21526);
nor U23583 (N_23583,N_21069,N_21978);
nand U23584 (N_23584,N_21281,N_21052);
and U23585 (N_23585,N_21652,N_21814);
nor U23586 (N_23586,N_20239,N_20316);
or U23587 (N_23587,N_20041,N_21093);
nor U23588 (N_23588,N_20778,N_20378);
nand U23589 (N_23589,N_20144,N_20583);
or U23590 (N_23590,N_20525,N_21075);
nor U23591 (N_23591,N_22092,N_20911);
nor U23592 (N_23592,N_22401,N_22359);
or U23593 (N_23593,N_20549,N_20058);
nand U23594 (N_23594,N_20567,N_20732);
nor U23595 (N_23595,N_21405,N_20385);
xor U23596 (N_23596,N_21899,N_21684);
or U23597 (N_23597,N_21384,N_20898);
or U23598 (N_23598,N_22424,N_20065);
or U23599 (N_23599,N_21599,N_21040);
nand U23600 (N_23600,N_20807,N_22253);
nand U23601 (N_23601,N_21110,N_20722);
nor U23602 (N_23602,N_20475,N_21727);
nand U23603 (N_23603,N_21850,N_21735);
or U23604 (N_23604,N_20640,N_20591);
and U23605 (N_23605,N_21986,N_22349);
nor U23606 (N_23606,N_20282,N_21838);
or U23607 (N_23607,N_20373,N_20820);
nor U23608 (N_23608,N_21753,N_20579);
xor U23609 (N_23609,N_21813,N_21280);
nor U23610 (N_23610,N_20073,N_21070);
and U23611 (N_23611,N_20675,N_22016);
nand U23612 (N_23612,N_20004,N_20462);
nand U23613 (N_23613,N_20428,N_22497);
nor U23614 (N_23614,N_20608,N_20714);
nand U23615 (N_23615,N_22220,N_20375);
and U23616 (N_23616,N_21596,N_21173);
nor U23617 (N_23617,N_20343,N_20057);
and U23618 (N_23618,N_20774,N_21226);
nand U23619 (N_23619,N_20179,N_20361);
nand U23620 (N_23620,N_20954,N_20616);
and U23621 (N_23621,N_20550,N_21102);
and U23622 (N_23622,N_21614,N_21984);
and U23623 (N_23623,N_22195,N_21059);
nand U23624 (N_23624,N_21964,N_21722);
or U23625 (N_23625,N_22093,N_21252);
and U23626 (N_23626,N_21172,N_20497);
nor U23627 (N_23627,N_20346,N_20752);
nor U23628 (N_23628,N_20899,N_21510);
and U23629 (N_23629,N_22200,N_21357);
nor U23630 (N_23630,N_22453,N_21108);
nor U23631 (N_23631,N_21747,N_22156);
or U23632 (N_23632,N_21054,N_20760);
nor U23633 (N_23633,N_22039,N_20966);
or U23634 (N_23634,N_22310,N_21138);
nor U23635 (N_23635,N_21750,N_22228);
nand U23636 (N_23636,N_21113,N_22005);
nand U23637 (N_23637,N_21581,N_20062);
and U23638 (N_23638,N_20541,N_20992);
nor U23639 (N_23639,N_22060,N_22372);
and U23640 (N_23640,N_20132,N_22335);
nand U23641 (N_23641,N_21078,N_22463);
or U23642 (N_23642,N_22062,N_20287);
or U23643 (N_23643,N_22194,N_21929);
and U23644 (N_23644,N_21926,N_21152);
and U23645 (N_23645,N_20470,N_21415);
and U23646 (N_23646,N_21212,N_21557);
nand U23647 (N_23647,N_21587,N_20182);
and U23648 (N_23648,N_20269,N_20725);
and U23649 (N_23649,N_21235,N_21004);
nand U23650 (N_23650,N_21388,N_21046);
or U23651 (N_23651,N_20145,N_22351);
and U23652 (N_23652,N_21532,N_20946);
nand U23653 (N_23653,N_21394,N_21954);
or U23654 (N_23654,N_20160,N_21320);
nor U23655 (N_23655,N_20204,N_22145);
nor U23656 (N_23656,N_20447,N_22254);
and U23657 (N_23657,N_20476,N_22272);
or U23658 (N_23658,N_20603,N_20997);
and U23659 (N_23659,N_22127,N_21028);
nor U23660 (N_23660,N_21829,N_20833);
and U23661 (N_23661,N_22021,N_22450);
nor U23662 (N_23662,N_21295,N_20513);
nand U23663 (N_23663,N_20933,N_20886);
nor U23664 (N_23664,N_21345,N_21339);
nand U23665 (N_23665,N_21117,N_21039);
and U23666 (N_23666,N_21072,N_21901);
or U23667 (N_23667,N_22213,N_21874);
nor U23668 (N_23668,N_20258,N_22267);
or U23669 (N_23669,N_21768,N_22068);
or U23670 (N_23670,N_21775,N_20074);
nand U23671 (N_23671,N_21579,N_21634);
and U23672 (N_23672,N_22397,N_20034);
or U23673 (N_23673,N_21071,N_21586);
and U23674 (N_23674,N_22395,N_21714);
nand U23675 (N_23675,N_22321,N_21992);
and U23676 (N_23676,N_21013,N_20815);
nor U23677 (N_23677,N_21809,N_20706);
and U23678 (N_23678,N_22421,N_20038);
and U23679 (N_23679,N_20942,N_21310);
and U23680 (N_23680,N_21246,N_21242);
nand U23681 (N_23681,N_22034,N_21144);
nand U23682 (N_23682,N_20523,N_21791);
or U23683 (N_23683,N_20789,N_20624);
nor U23684 (N_23684,N_21729,N_21998);
nand U23685 (N_23685,N_20431,N_21221);
or U23686 (N_23686,N_21380,N_21851);
or U23687 (N_23687,N_22018,N_21049);
or U23688 (N_23688,N_22161,N_22032);
nor U23689 (N_23689,N_20028,N_21509);
and U23690 (N_23690,N_20988,N_22240);
or U23691 (N_23691,N_20814,N_21712);
nand U23692 (N_23692,N_20356,N_20633);
nand U23693 (N_23693,N_22273,N_21564);
nand U23694 (N_23694,N_21378,N_22221);
nand U23695 (N_23695,N_21961,N_21207);
and U23696 (N_23696,N_21208,N_20619);
and U23697 (N_23697,N_21806,N_21682);
or U23698 (N_23698,N_20174,N_21141);
or U23699 (N_23699,N_22012,N_21148);
nor U23700 (N_23700,N_21245,N_20797);
and U23701 (N_23701,N_21765,N_21876);
and U23702 (N_23702,N_20654,N_22281);
and U23703 (N_23703,N_22196,N_22148);
or U23704 (N_23704,N_22285,N_21976);
or U23705 (N_23705,N_21444,N_22348);
and U23706 (N_23706,N_20768,N_20787);
nand U23707 (N_23707,N_20751,N_20794);
nand U23708 (N_23708,N_20618,N_21218);
nand U23709 (N_23709,N_20888,N_20500);
or U23710 (N_23710,N_20308,N_22287);
nor U23711 (N_23711,N_21375,N_21811);
or U23712 (N_23712,N_20684,N_22477);
nor U23713 (N_23713,N_21995,N_22212);
and U23714 (N_23714,N_20377,N_20543);
or U23715 (N_23715,N_21866,N_21376);
xnor U23716 (N_23716,N_20013,N_22186);
nor U23717 (N_23717,N_20962,N_21057);
nand U23718 (N_23718,N_21680,N_21076);
or U23719 (N_23719,N_21789,N_20941);
nand U23720 (N_23720,N_21592,N_20115);
nand U23721 (N_23721,N_22048,N_21160);
nor U23722 (N_23722,N_22129,N_20054);
or U23723 (N_23723,N_20723,N_20743);
or U23724 (N_23724,N_20585,N_20630);
or U23725 (N_23725,N_22100,N_21482);
and U23726 (N_23726,N_21847,N_21903);
and U23727 (N_23727,N_21279,N_21602);
and U23728 (N_23728,N_22033,N_20153);
nor U23729 (N_23729,N_20832,N_21709);
nor U23730 (N_23730,N_21171,N_20031);
nor U23731 (N_23731,N_20071,N_21662);
or U23732 (N_23732,N_20415,N_21062);
nor U23733 (N_23733,N_22120,N_21631);
nor U23734 (N_23734,N_21323,N_21967);
nand U23735 (N_23735,N_20928,N_21296);
or U23736 (N_23736,N_21577,N_21522);
nand U23737 (N_23737,N_20599,N_20264);
or U23738 (N_23738,N_22458,N_21795);
nor U23739 (N_23739,N_21048,N_20915);
xor U23740 (N_23740,N_21583,N_21563);
nand U23741 (N_23741,N_22420,N_20577);
nor U23742 (N_23742,N_22499,N_22311);
nand U23743 (N_23743,N_21190,N_21640);
and U23744 (N_23744,N_20197,N_21756);
xor U23745 (N_23745,N_22164,N_20636);
and U23746 (N_23746,N_20302,N_20695);
and U23747 (N_23747,N_21616,N_21021);
nand U23748 (N_23748,N_21269,N_20735);
or U23749 (N_23749,N_21291,N_20562);
nor U23750 (N_23750,N_20548,N_21011);
and U23751 (N_23751,N_21508,N_21779);
or U23752 (N_23752,N_22343,N_20962);
nand U23753 (N_23753,N_22096,N_20366);
and U23754 (N_23754,N_20627,N_21243);
or U23755 (N_23755,N_21405,N_22069);
nor U23756 (N_23756,N_20114,N_21837);
and U23757 (N_23757,N_21501,N_22375);
or U23758 (N_23758,N_21357,N_22263);
nand U23759 (N_23759,N_20412,N_21711);
and U23760 (N_23760,N_20277,N_20667);
nand U23761 (N_23761,N_21108,N_21449);
or U23762 (N_23762,N_20005,N_20875);
nor U23763 (N_23763,N_21402,N_21301);
and U23764 (N_23764,N_20755,N_22381);
nand U23765 (N_23765,N_20690,N_20701);
or U23766 (N_23766,N_21113,N_21143);
or U23767 (N_23767,N_20307,N_20936);
nand U23768 (N_23768,N_20106,N_22475);
nand U23769 (N_23769,N_20573,N_20784);
nand U23770 (N_23770,N_20449,N_21345);
nand U23771 (N_23771,N_21856,N_21455);
and U23772 (N_23772,N_21636,N_20830);
or U23773 (N_23773,N_20892,N_21094);
or U23774 (N_23774,N_20490,N_20173);
or U23775 (N_23775,N_20548,N_22261);
nor U23776 (N_23776,N_22108,N_22364);
and U23777 (N_23777,N_21807,N_20221);
nand U23778 (N_23778,N_20679,N_20497);
nor U23779 (N_23779,N_22043,N_22410);
and U23780 (N_23780,N_22368,N_21699);
or U23781 (N_23781,N_22452,N_20129);
xor U23782 (N_23782,N_21212,N_20246);
or U23783 (N_23783,N_22032,N_21188);
and U23784 (N_23784,N_21544,N_22165);
or U23785 (N_23785,N_20164,N_20568);
nand U23786 (N_23786,N_21769,N_22278);
or U23787 (N_23787,N_21221,N_21676);
nand U23788 (N_23788,N_20418,N_22346);
or U23789 (N_23789,N_20464,N_21981);
and U23790 (N_23790,N_21295,N_21822);
nor U23791 (N_23791,N_21686,N_22470);
xnor U23792 (N_23792,N_20808,N_21578);
and U23793 (N_23793,N_20630,N_21239);
and U23794 (N_23794,N_20497,N_20343);
and U23795 (N_23795,N_20608,N_21218);
xnor U23796 (N_23796,N_20014,N_20218);
and U23797 (N_23797,N_22452,N_22161);
nand U23798 (N_23798,N_22028,N_21105);
nor U23799 (N_23799,N_21228,N_21604);
and U23800 (N_23800,N_20655,N_20053);
nor U23801 (N_23801,N_20874,N_21507);
nor U23802 (N_23802,N_21299,N_20824);
nand U23803 (N_23803,N_20710,N_20978);
and U23804 (N_23804,N_21575,N_20435);
nor U23805 (N_23805,N_20813,N_20257);
nand U23806 (N_23806,N_20681,N_21434);
nand U23807 (N_23807,N_21081,N_20206);
nand U23808 (N_23808,N_20141,N_22078);
nor U23809 (N_23809,N_21672,N_21433);
nor U23810 (N_23810,N_20625,N_21174);
or U23811 (N_23811,N_22137,N_21778);
or U23812 (N_23812,N_21216,N_20266);
nand U23813 (N_23813,N_21483,N_22195);
or U23814 (N_23814,N_21663,N_20030);
nor U23815 (N_23815,N_21624,N_20731);
nand U23816 (N_23816,N_20470,N_21187);
nor U23817 (N_23817,N_22166,N_20519);
or U23818 (N_23818,N_20461,N_21614);
or U23819 (N_23819,N_21518,N_21529);
nand U23820 (N_23820,N_21744,N_21763);
and U23821 (N_23821,N_21873,N_22346);
and U23822 (N_23822,N_20330,N_21375);
and U23823 (N_23823,N_21243,N_22004);
nand U23824 (N_23824,N_20969,N_20436);
or U23825 (N_23825,N_22270,N_20605);
and U23826 (N_23826,N_22215,N_21227);
or U23827 (N_23827,N_22027,N_22166);
nor U23828 (N_23828,N_22260,N_21050);
nor U23829 (N_23829,N_20369,N_22289);
nand U23830 (N_23830,N_20688,N_21375);
nor U23831 (N_23831,N_22362,N_21840);
nor U23832 (N_23832,N_20135,N_20584);
nor U23833 (N_23833,N_22409,N_20714);
nor U23834 (N_23834,N_20513,N_21438);
nor U23835 (N_23835,N_21368,N_20555);
nand U23836 (N_23836,N_22303,N_20935);
or U23837 (N_23837,N_21305,N_20934);
nor U23838 (N_23838,N_20004,N_21002);
xor U23839 (N_23839,N_20143,N_22249);
nand U23840 (N_23840,N_21081,N_21468);
or U23841 (N_23841,N_21539,N_20202);
and U23842 (N_23842,N_20749,N_21108);
nor U23843 (N_23843,N_20357,N_20818);
and U23844 (N_23844,N_21747,N_21286);
or U23845 (N_23845,N_21021,N_22357);
and U23846 (N_23846,N_21590,N_20650);
xnor U23847 (N_23847,N_20169,N_20286);
and U23848 (N_23848,N_22245,N_22049);
nor U23849 (N_23849,N_20512,N_22211);
nand U23850 (N_23850,N_22070,N_21743);
nor U23851 (N_23851,N_22337,N_22061);
and U23852 (N_23852,N_21610,N_20623);
or U23853 (N_23853,N_20190,N_21643);
or U23854 (N_23854,N_22245,N_21533);
or U23855 (N_23855,N_20289,N_21078);
nand U23856 (N_23856,N_22119,N_21038);
or U23857 (N_23857,N_21515,N_22023);
nand U23858 (N_23858,N_21444,N_20856);
or U23859 (N_23859,N_20403,N_21616);
nand U23860 (N_23860,N_20102,N_22087);
and U23861 (N_23861,N_21548,N_20930);
nand U23862 (N_23862,N_21660,N_20794);
nand U23863 (N_23863,N_20743,N_22041);
nand U23864 (N_23864,N_20862,N_20152);
and U23865 (N_23865,N_21581,N_20633);
and U23866 (N_23866,N_20176,N_21042);
nor U23867 (N_23867,N_20532,N_21807);
nor U23868 (N_23868,N_22031,N_21995);
and U23869 (N_23869,N_20464,N_21385);
nor U23870 (N_23870,N_20134,N_21844);
nand U23871 (N_23871,N_21853,N_22252);
nand U23872 (N_23872,N_20532,N_21165);
or U23873 (N_23873,N_21257,N_21932);
nor U23874 (N_23874,N_20720,N_20253);
or U23875 (N_23875,N_20208,N_20402);
nor U23876 (N_23876,N_22166,N_20239);
nor U23877 (N_23877,N_21997,N_20224);
nand U23878 (N_23878,N_20598,N_20306);
nor U23879 (N_23879,N_20615,N_20513);
nor U23880 (N_23880,N_20839,N_20882);
nand U23881 (N_23881,N_22395,N_20295);
or U23882 (N_23882,N_21203,N_20872);
and U23883 (N_23883,N_20961,N_20468);
nor U23884 (N_23884,N_20431,N_21499);
nand U23885 (N_23885,N_20530,N_20902);
or U23886 (N_23886,N_20636,N_21880);
or U23887 (N_23887,N_21092,N_20092);
nor U23888 (N_23888,N_20602,N_21777);
or U23889 (N_23889,N_21648,N_20331);
or U23890 (N_23890,N_22196,N_20179);
or U23891 (N_23891,N_20916,N_21250);
nor U23892 (N_23892,N_22067,N_21574);
and U23893 (N_23893,N_20045,N_20637);
nand U23894 (N_23894,N_21178,N_21931);
nor U23895 (N_23895,N_20113,N_21144);
or U23896 (N_23896,N_21984,N_20266);
nand U23897 (N_23897,N_20400,N_20399);
nor U23898 (N_23898,N_21432,N_22377);
nand U23899 (N_23899,N_20417,N_22028);
nor U23900 (N_23900,N_21221,N_21893);
or U23901 (N_23901,N_21508,N_21211);
and U23902 (N_23902,N_21744,N_20449);
nand U23903 (N_23903,N_20089,N_21645);
nor U23904 (N_23904,N_21691,N_22406);
or U23905 (N_23905,N_20719,N_20627);
and U23906 (N_23906,N_20732,N_22053);
nand U23907 (N_23907,N_21785,N_21033);
or U23908 (N_23908,N_20894,N_21656);
nor U23909 (N_23909,N_21839,N_20595);
nor U23910 (N_23910,N_20667,N_20742);
nand U23911 (N_23911,N_21044,N_21357);
nand U23912 (N_23912,N_21527,N_20156);
and U23913 (N_23913,N_20323,N_21695);
or U23914 (N_23914,N_20580,N_20167);
nor U23915 (N_23915,N_20882,N_21752);
nand U23916 (N_23916,N_20596,N_22366);
and U23917 (N_23917,N_20346,N_21470);
or U23918 (N_23918,N_21737,N_20818);
nand U23919 (N_23919,N_21648,N_22405);
and U23920 (N_23920,N_20984,N_22294);
nor U23921 (N_23921,N_20592,N_20231);
nor U23922 (N_23922,N_21276,N_21811);
or U23923 (N_23923,N_20884,N_22136);
nor U23924 (N_23924,N_21329,N_20035);
nand U23925 (N_23925,N_21086,N_21672);
or U23926 (N_23926,N_20141,N_20026);
nor U23927 (N_23927,N_21590,N_21391);
and U23928 (N_23928,N_22078,N_20638);
and U23929 (N_23929,N_21844,N_21495);
nor U23930 (N_23930,N_20100,N_21363);
nand U23931 (N_23931,N_21181,N_20426);
nor U23932 (N_23932,N_21209,N_20932);
nand U23933 (N_23933,N_20909,N_22053);
or U23934 (N_23934,N_21656,N_22084);
nand U23935 (N_23935,N_21800,N_20158);
nor U23936 (N_23936,N_22395,N_22495);
and U23937 (N_23937,N_22372,N_21794);
and U23938 (N_23938,N_20248,N_21361);
nor U23939 (N_23939,N_22299,N_21568);
nor U23940 (N_23940,N_20829,N_21436);
or U23941 (N_23941,N_20662,N_20590);
nor U23942 (N_23942,N_21377,N_20389);
nor U23943 (N_23943,N_20184,N_20097);
nand U23944 (N_23944,N_20043,N_21929);
or U23945 (N_23945,N_22326,N_20230);
nand U23946 (N_23946,N_20981,N_21032);
and U23947 (N_23947,N_21978,N_21776);
nand U23948 (N_23948,N_20868,N_21294);
nand U23949 (N_23949,N_20019,N_20579);
or U23950 (N_23950,N_20667,N_22111);
xnor U23951 (N_23951,N_21209,N_20790);
and U23952 (N_23952,N_22077,N_21692);
and U23953 (N_23953,N_20507,N_20564);
and U23954 (N_23954,N_21740,N_21915);
nand U23955 (N_23955,N_20410,N_21745);
nor U23956 (N_23956,N_21857,N_22347);
nand U23957 (N_23957,N_20968,N_21161);
or U23958 (N_23958,N_22488,N_21676);
nor U23959 (N_23959,N_21783,N_21469);
nor U23960 (N_23960,N_20726,N_22120);
and U23961 (N_23961,N_20706,N_20525);
nand U23962 (N_23962,N_21982,N_22208);
nor U23963 (N_23963,N_22166,N_21752);
and U23964 (N_23964,N_20050,N_20448);
or U23965 (N_23965,N_21875,N_20633);
and U23966 (N_23966,N_22419,N_20855);
or U23967 (N_23967,N_20985,N_22209);
and U23968 (N_23968,N_22318,N_20019);
nand U23969 (N_23969,N_20462,N_20985);
or U23970 (N_23970,N_21649,N_20527);
and U23971 (N_23971,N_20663,N_21269);
nor U23972 (N_23972,N_20598,N_22421);
and U23973 (N_23973,N_20329,N_20839);
nand U23974 (N_23974,N_20075,N_21691);
or U23975 (N_23975,N_21286,N_20776);
or U23976 (N_23976,N_22359,N_20841);
nor U23977 (N_23977,N_21553,N_21252);
or U23978 (N_23978,N_20994,N_20485);
and U23979 (N_23979,N_20102,N_21540);
or U23980 (N_23980,N_22180,N_22256);
and U23981 (N_23981,N_21856,N_20620);
and U23982 (N_23982,N_21781,N_20495);
nor U23983 (N_23983,N_21312,N_21165);
nor U23984 (N_23984,N_20487,N_22429);
nor U23985 (N_23985,N_20211,N_22468);
nand U23986 (N_23986,N_21586,N_20827);
nand U23987 (N_23987,N_21746,N_20278);
nor U23988 (N_23988,N_21015,N_21585);
nor U23989 (N_23989,N_21855,N_20970);
nor U23990 (N_23990,N_20886,N_20031);
and U23991 (N_23991,N_21631,N_21079);
nor U23992 (N_23992,N_21951,N_20856);
nand U23993 (N_23993,N_20396,N_21918);
xnor U23994 (N_23994,N_21753,N_21122);
and U23995 (N_23995,N_22410,N_21411);
or U23996 (N_23996,N_20493,N_20969);
and U23997 (N_23997,N_20318,N_20771);
nor U23998 (N_23998,N_21102,N_21830);
nor U23999 (N_23999,N_21782,N_22450);
nand U24000 (N_24000,N_22167,N_21056);
nand U24001 (N_24001,N_21746,N_21536);
nand U24002 (N_24002,N_20791,N_21506);
nor U24003 (N_24003,N_21684,N_21670);
nand U24004 (N_24004,N_21097,N_22326);
nand U24005 (N_24005,N_21874,N_21819);
nor U24006 (N_24006,N_20273,N_21652);
or U24007 (N_24007,N_20299,N_20612);
or U24008 (N_24008,N_20945,N_21162);
nor U24009 (N_24009,N_22443,N_21715);
or U24010 (N_24010,N_21991,N_20619);
nand U24011 (N_24011,N_21404,N_21494);
nand U24012 (N_24012,N_20841,N_20313);
or U24013 (N_24013,N_20216,N_20263);
nand U24014 (N_24014,N_20259,N_20077);
nor U24015 (N_24015,N_21148,N_22456);
nor U24016 (N_24016,N_21677,N_22107);
and U24017 (N_24017,N_22020,N_20443);
nand U24018 (N_24018,N_20493,N_20083);
or U24019 (N_24019,N_20103,N_21609);
nand U24020 (N_24020,N_22297,N_20023);
nand U24021 (N_24021,N_21236,N_20362);
and U24022 (N_24022,N_22340,N_20052);
nor U24023 (N_24023,N_21682,N_20575);
nor U24024 (N_24024,N_22156,N_20491);
nand U24025 (N_24025,N_22153,N_21014);
nand U24026 (N_24026,N_21851,N_20133);
nand U24027 (N_24027,N_20851,N_20869);
or U24028 (N_24028,N_21135,N_21149);
nor U24029 (N_24029,N_20396,N_20931);
and U24030 (N_24030,N_20328,N_20100);
or U24031 (N_24031,N_21767,N_20931);
nand U24032 (N_24032,N_20893,N_21416);
or U24033 (N_24033,N_20483,N_21622);
xor U24034 (N_24034,N_20654,N_20975);
nand U24035 (N_24035,N_22159,N_20580);
nor U24036 (N_24036,N_21429,N_20256);
nor U24037 (N_24037,N_22301,N_22071);
or U24038 (N_24038,N_20171,N_20248);
or U24039 (N_24039,N_22391,N_20556);
nand U24040 (N_24040,N_22299,N_21073);
nor U24041 (N_24041,N_22399,N_20062);
nand U24042 (N_24042,N_21374,N_20124);
nor U24043 (N_24043,N_20025,N_20650);
and U24044 (N_24044,N_22143,N_20640);
or U24045 (N_24045,N_20913,N_20191);
and U24046 (N_24046,N_21346,N_22112);
and U24047 (N_24047,N_22084,N_20644);
or U24048 (N_24048,N_20122,N_20909);
or U24049 (N_24049,N_21977,N_20981);
nand U24050 (N_24050,N_20515,N_22393);
or U24051 (N_24051,N_21262,N_21787);
or U24052 (N_24052,N_22193,N_21165);
or U24053 (N_24053,N_20687,N_22173);
nor U24054 (N_24054,N_22191,N_21226);
and U24055 (N_24055,N_21424,N_21101);
nor U24056 (N_24056,N_21706,N_21572);
and U24057 (N_24057,N_20731,N_21364);
or U24058 (N_24058,N_20153,N_22404);
or U24059 (N_24059,N_22074,N_20472);
and U24060 (N_24060,N_22275,N_21394);
nor U24061 (N_24061,N_21566,N_21781);
nand U24062 (N_24062,N_20654,N_21353);
nor U24063 (N_24063,N_20498,N_21183);
or U24064 (N_24064,N_21934,N_20381);
nor U24065 (N_24065,N_20522,N_20728);
and U24066 (N_24066,N_22100,N_21304);
nor U24067 (N_24067,N_21799,N_22156);
nor U24068 (N_24068,N_22181,N_21779);
and U24069 (N_24069,N_21913,N_22423);
nand U24070 (N_24070,N_21026,N_21687);
and U24071 (N_24071,N_21502,N_20552);
nand U24072 (N_24072,N_21472,N_22480);
nand U24073 (N_24073,N_21197,N_21736);
and U24074 (N_24074,N_21304,N_21749);
or U24075 (N_24075,N_21533,N_21946);
and U24076 (N_24076,N_20166,N_20510);
nand U24077 (N_24077,N_21682,N_21671);
nand U24078 (N_24078,N_21315,N_21187);
or U24079 (N_24079,N_20621,N_20929);
nand U24080 (N_24080,N_20207,N_20907);
nand U24081 (N_24081,N_20954,N_22090);
nor U24082 (N_24082,N_21911,N_22268);
or U24083 (N_24083,N_21888,N_20297);
or U24084 (N_24084,N_22199,N_20375);
and U24085 (N_24085,N_22006,N_20823);
nand U24086 (N_24086,N_22194,N_21478);
and U24087 (N_24087,N_21294,N_21732);
and U24088 (N_24088,N_22269,N_21124);
nand U24089 (N_24089,N_20379,N_22222);
nand U24090 (N_24090,N_20997,N_20017);
nand U24091 (N_24091,N_21620,N_21736);
and U24092 (N_24092,N_22456,N_21872);
and U24093 (N_24093,N_21102,N_21608);
xor U24094 (N_24094,N_21743,N_21332);
and U24095 (N_24095,N_21811,N_21907);
nor U24096 (N_24096,N_21925,N_22087);
or U24097 (N_24097,N_21934,N_20246);
nand U24098 (N_24098,N_20611,N_21270);
nor U24099 (N_24099,N_20340,N_20585);
nor U24100 (N_24100,N_21410,N_21079);
xor U24101 (N_24101,N_21890,N_20129);
nand U24102 (N_24102,N_20052,N_21418);
nand U24103 (N_24103,N_20274,N_21848);
and U24104 (N_24104,N_22372,N_21042);
nand U24105 (N_24105,N_22391,N_21319);
nor U24106 (N_24106,N_21762,N_20513);
nor U24107 (N_24107,N_20125,N_21017);
or U24108 (N_24108,N_21714,N_20049);
nor U24109 (N_24109,N_22453,N_22243);
nand U24110 (N_24110,N_22427,N_21769);
nor U24111 (N_24111,N_20807,N_21562);
nor U24112 (N_24112,N_21826,N_20130);
nand U24113 (N_24113,N_22315,N_21207);
nor U24114 (N_24114,N_20312,N_22230);
or U24115 (N_24115,N_21633,N_20633);
xnor U24116 (N_24116,N_22201,N_20585);
or U24117 (N_24117,N_20965,N_20633);
nor U24118 (N_24118,N_20221,N_21558);
or U24119 (N_24119,N_20204,N_21965);
nor U24120 (N_24120,N_21482,N_21552);
or U24121 (N_24121,N_22222,N_21233);
nand U24122 (N_24122,N_20724,N_21037);
or U24123 (N_24123,N_20822,N_20552);
nand U24124 (N_24124,N_20737,N_21061);
and U24125 (N_24125,N_20048,N_20615);
and U24126 (N_24126,N_20757,N_22313);
nor U24127 (N_24127,N_22473,N_20200);
and U24128 (N_24128,N_20138,N_21831);
nand U24129 (N_24129,N_20151,N_20657);
and U24130 (N_24130,N_21279,N_22144);
nand U24131 (N_24131,N_22387,N_21723);
xor U24132 (N_24132,N_21082,N_21857);
or U24133 (N_24133,N_22111,N_21591);
or U24134 (N_24134,N_20433,N_21687);
nor U24135 (N_24135,N_21713,N_20049);
or U24136 (N_24136,N_20636,N_21272);
nor U24137 (N_24137,N_20872,N_20969);
or U24138 (N_24138,N_20753,N_22210);
nand U24139 (N_24139,N_20503,N_20642);
nand U24140 (N_24140,N_20351,N_22327);
and U24141 (N_24141,N_21967,N_21633);
nor U24142 (N_24142,N_21040,N_20046);
or U24143 (N_24143,N_20136,N_21454);
or U24144 (N_24144,N_22050,N_20567);
nand U24145 (N_24145,N_21629,N_20638);
xor U24146 (N_24146,N_20719,N_21175);
and U24147 (N_24147,N_22214,N_20528);
nor U24148 (N_24148,N_20961,N_20851);
nand U24149 (N_24149,N_20349,N_21545);
or U24150 (N_24150,N_22024,N_21734);
and U24151 (N_24151,N_21885,N_21481);
nor U24152 (N_24152,N_20419,N_21556);
nor U24153 (N_24153,N_20624,N_21897);
and U24154 (N_24154,N_20806,N_20756);
nand U24155 (N_24155,N_20762,N_21474);
nor U24156 (N_24156,N_22291,N_20234);
nand U24157 (N_24157,N_20460,N_21703);
and U24158 (N_24158,N_22204,N_20573);
or U24159 (N_24159,N_22126,N_21753);
and U24160 (N_24160,N_21381,N_22430);
and U24161 (N_24161,N_21581,N_21279);
nor U24162 (N_24162,N_20400,N_21828);
or U24163 (N_24163,N_20671,N_22422);
nor U24164 (N_24164,N_21318,N_22063);
nand U24165 (N_24165,N_21316,N_21905);
nor U24166 (N_24166,N_20768,N_20479);
xnor U24167 (N_24167,N_20431,N_20433);
or U24168 (N_24168,N_20855,N_21330);
nor U24169 (N_24169,N_21062,N_21203);
nor U24170 (N_24170,N_21380,N_20683);
nor U24171 (N_24171,N_20087,N_20699);
nor U24172 (N_24172,N_21366,N_20473);
nor U24173 (N_24173,N_21141,N_21183);
nor U24174 (N_24174,N_21244,N_22252);
nor U24175 (N_24175,N_20111,N_20541);
nor U24176 (N_24176,N_20160,N_20691);
and U24177 (N_24177,N_20227,N_20641);
and U24178 (N_24178,N_22219,N_21461);
and U24179 (N_24179,N_21087,N_22331);
nand U24180 (N_24180,N_20614,N_22191);
nor U24181 (N_24181,N_22241,N_22122);
nor U24182 (N_24182,N_22419,N_21863);
nor U24183 (N_24183,N_21812,N_20354);
nand U24184 (N_24184,N_21336,N_21654);
or U24185 (N_24185,N_21738,N_21837);
or U24186 (N_24186,N_20599,N_20953);
nor U24187 (N_24187,N_21106,N_20448);
nor U24188 (N_24188,N_20038,N_21771);
or U24189 (N_24189,N_20387,N_22235);
and U24190 (N_24190,N_21823,N_22020);
and U24191 (N_24191,N_22273,N_21594);
and U24192 (N_24192,N_20314,N_21545);
and U24193 (N_24193,N_21027,N_20432);
or U24194 (N_24194,N_20832,N_20058);
or U24195 (N_24195,N_20483,N_20511);
or U24196 (N_24196,N_20431,N_20161);
or U24197 (N_24197,N_21280,N_20409);
and U24198 (N_24198,N_21556,N_20021);
and U24199 (N_24199,N_20711,N_20782);
nand U24200 (N_24200,N_20769,N_22329);
and U24201 (N_24201,N_20213,N_20031);
and U24202 (N_24202,N_21346,N_22272);
or U24203 (N_24203,N_22325,N_20531);
nand U24204 (N_24204,N_22233,N_20117);
or U24205 (N_24205,N_21868,N_20684);
and U24206 (N_24206,N_20162,N_22318);
and U24207 (N_24207,N_21707,N_20060);
nor U24208 (N_24208,N_20638,N_21664);
or U24209 (N_24209,N_22394,N_22418);
nand U24210 (N_24210,N_21792,N_22171);
or U24211 (N_24211,N_20450,N_21154);
nor U24212 (N_24212,N_22415,N_21642);
nor U24213 (N_24213,N_21241,N_21135);
and U24214 (N_24214,N_21562,N_21718);
nor U24215 (N_24215,N_21965,N_20099);
or U24216 (N_24216,N_20349,N_22303);
and U24217 (N_24217,N_21653,N_20191);
nor U24218 (N_24218,N_20355,N_21539);
nor U24219 (N_24219,N_22236,N_20258);
nor U24220 (N_24220,N_22039,N_21354);
and U24221 (N_24221,N_22364,N_20611);
nor U24222 (N_24222,N_21708,N_22491);
or U24223 (N_24223,N_20704,N_21270);
nand U24224 (N_24224,N_20027,N_21506);
nor U24225 (N_24225,N_21232,N_20955);
or U24226 (N_24226,N_22270,N_20265);
nand U24227 (N_24227,N_22329,N_21584);
nand U24228 (N_24228,N_21869,N_20943);
or U24229 (N_24229,N_20428,N_21829);
nor U24230 (N_24230,N_22199,N_20185);
nor U24231 (N_24231,N_22445,N_21808);
or U24232 (N_24232,N_22125,N_20063);
nor U24233 (N_24233,N_20134,N_20609);
or U24234 (N_24234,N_21342,N_21683);
nor U24235 (N_24235,N_21007,N_21041);
nand U24236 (N_24236,N_22367,N_20298);
nand U24237 (N_24237,N_21779,N_20577);
xor U24238 (N_24238,N_20642,N_20456);
nand U24239 (N_24239,N_21468,N_21463);
nand U24240 (N_24240,N_22332,N_21994);
or U24241 (N_24241,N_21981,N_21561);
nor U24242 (N_24242,N_20777,N_21019);
nand U24243 (N_24243,N_22276,N_20841);
and U24244 (N_24244,N_21060,N_20297);
or U24245 (N_24245,N_20868,N_21095);
nor U24246 (N_24246,N_21799,N_20351);
and U24247 (N_24247,N_20631,N_21818);
nor U24248 (N_24248,N_21276,N_20808);
or U24249 (N_24249,N_21848,N_20163);
nor U24250 (N_24250,N_21965,N_22111);
or U24251 (N_24251,N_22080,N_21873);
nor U24252 (N_24252,N_22434,N_20234);
nor U24253 (N_24253,N_21303,N_21099);
xnor U24254 (N_24254,N_22088,N_22142);
nand U24255 (N_24255,N_21884,N_22063);
nand U24256 (N_24256,N_21744,N_20208);
xnor U24257 (N_24257,N_20443,N_20132);
or U24258 (N_24258,N_21027,N_21010);
nor U24259 (N_24259,N_21462,N_21550);
or U24260 (N_24260,N_21453,N_21218);
nor U24261 (N_24261,N_20220,N_22374);
nand U24262 (N_24262,N_20203,N_22039);
nor U24263 (N_24263,N_21372,N_21409);
or U24264 (N_24264,N_21546,N_20207);
nand U24265 (N_24265,N_20068,N_22168);
nand U24266 (N_24266,N_20322,N_21302);
or U24267 (N_24267,N_20498,N_21048);
nand U24268 (N_24268,N_20867,N_22044);
and U24269 (N_24269,N_20527,N_20260);
nand U24270 (N_24270,N_21304,N_20360);
nand U24271 (N_24271,N_20411,N_20808);
nor U24272 (N_24272,N_21341,N_21304);
nor U24273 (N_24273,N_22206,N_22007);
nor U24274 (N_24274,N_20225,N_22197);
or U24275 (N_24275,N_21020,N_20912);
and U24276 (N_24276,N_21824,N_20825);
or U24277 (N_24277,N_20430,N_20491);
nor U24278 (N_24278,N_22266,N_21582);
and U24279 (N_24279,N_20963,N_21720);
or U24280 (N_24280,N_22174,N_22020);
or U24281 (N_24281,N_20167,N_20985);
nand U24282 (N_24282,N_20642,N_22332);
nor U24283 (N_24283,N_20845,N_21858);
nand U24284 (N_24284,N_21521,N_21538);
or U24285 (N_24285,N_20733,N_20111);
nand U24286 (N_24286,N_20980,N_21932);
or U24287 (N_24287,N_20281,N_22140);
nand U24288 (N_24288,N_20558,N_21121);
nor U24289 (N_24289,N_21996,N_21112);
nor U24290 (N_24290,N_22025,N_21507);
and U24291 (N_24291,N_21945,N_22079);
or U24292 (N_24292,N_21268,N_21843);
nor U24293 (N_24293,N_22097,N_20938);
nor U24294 (N_24294,N_20332,N_22269);
nor U24295 (N_24295,N_20780,N_21598);
and U24296 (N_24296,N_21349,N_21803);
nand U24297 (N_24297,N_21211,N_20040);
nand U24298 (N_24298,N_22293,N_21122);
or U24299 (N_24299,N_22000,N_22182);
nor U24300 (N_24300,N_22040,N_20823);
and U24301 (N_24301,N_22238,N_22036);
nor U24302 (N_24302,N_21778,N_21524);
or U24303 (N_24303,N_21528,N_20570);
nand U24304 (N_24304,N_20823,N_22498);
and U24305 (N_24305,N_20244,N_20975);
xnor U24306 (N_24306,N_20927,N_20951);
and U24307 (N_24307,N_20502,N_20096);
nor U24308 (N_24308,N_21206,N_20783);
and U24309 (N_24309,N_21805,N_22369);
nand U24310 (N_24310,N_20624,N_21279);
nor U24311 (N_24311,N_21762,N_20136);
nor U24312 (N_24312,N_20160,N_21532);
nor U24313 (N_24313,N_21956,N_21766);
nand U24314 (N_24314,N_22361,N_22384);
xnor U24315 (N_24315,N_21079,N_21547);
nor U24316 (N_24316,N_21775,N_21330);
nor U24317 (N_24317,N_20433,N_21938);
or U24318 (N_24318,N_21452,N_20822);
nor U24319 (N_24319,N_20431,N_21130);
nand U24320 (N_24320,N_21839,N_20196);
nor U24321 (N_24321,N_20294,N_22050);
or U24322 (N_24322,N_22225,N_21836);
nor U24323 (N_24323,N_21769,N_21994);
nor U24324 (N_24324,N_22385,N_21262);
nand U24325 (N_24325,N_21081,N_20916);
and U24326 (N_24326,N_20030,N_22084);
nand U24327 (N_24327,N_21753,N_20704);
nand U24328 (N_24328,N_20460,N_20170);
nand U24329 (N_24329,N_20701,N_21747);
nor U24330 (N_24330,N_21197,N_20670);
and U24331 (N_24331,N_20483,N_21945);
and U24332 (N_24332,N_21476,N_22011);
nor U24333 (N_24333,N_22440,N_21566);
or U24334 (N_24334,N_20257,N_21754);
and U24335 (N_24335,N_20277,N_22383);
nand U24336 (N_24336,N_22426,N_21285);
and U24337 (N_24337,N_20031,N_22325);
and U24338 (N_24338,N_20522,N_20634);
and U24339 (N_24339,N_20711,N_22472);
nor U24340 (N_24340,N_22048,N_21078);
nor U24341 (N_24341,N_22132,N_22091);
or U24342 (N_24342,N_20812,N_22420);
nand U24343 (N_24343,N_21660,N_22082);
or U24344 (N_24344,N_21300,N_22189);
and U24345 (N_24345,N_22372,N_20712);
or U24346 (N_24346,N_20234,N_21096);
nor U24347 (N_24347,N_20919,N_21457);
and U24348 (N_24348,N_20282,N_20391);
nor U24349 (N_24349,N_20202,N_20801);
and U24350 (N_24350,N_20348,N_20554);
nand U24351 (N_24351,N_20166,N_22374);
or U24352 (N_24352,N_21988,N_21620);
nand U24353 (N_24353,N_21643,N_20462);
nor U24354 (N_24354,N_21828,N_21128);
nand U24355 (N_24355,N_22282,N_22286);
nor U24356 (N_24356,N_21855,N_22204);
nand U24357 (N_24357,N_22423,N_20510);
or U24358 (N_24358,N_20252,N_21895);
and U24359 (N_24359,N_21185,N_22313);
nand U24360 (N_24360,N_21670,N_21812);
nand U24361 (N_24361,N_22153,N_22365);
and U24362 (N_24362,N_21833,N_21451);
nand U24363 (N_24363,N_21235,N_22239);
nor U24364 (N_24364,N_21476,N_21923);
nand U24365 (N_24365,N_22401,N_20294);
and U24366 (N_24366,N_21312,N_20663);
or U24367 (N_24367,N_21269,N_20463);
or U24368 (N_24368,N_21968,N_20560);
and U24369 (N_24369,N_21141,N_21439);
and U24370 (N_24370,N_21353,N_20424);
or U24371 (N_24371,N_22288,N_21882);
nor U24372 (N_24372,N_22331,N_20789);
nor U24373 (N_24373,N_20643,N_21593);
nand U24374 (N_24374,N_20973,N_20779);
nor U24375 (N_24375,N_21131,N_21151);
nor U24376 (N_24376,N_21055,N_20413);
nand U24377 (N_24377,N_21762,N_20515);
nand U24378 (N_24378,N_21600,N_20673);
nor U24379 (N_24379,N_20162,N_20306);
nand U24380 (N_24380,N_21382,N_20917);
or U24381 (N_24381,N_20707,N_21713);
nand U24382 (N_24382,N_22121,N_20815);
nand U24383 (N_24383,N_21508,N_21637);
nand U24384 (N_24384,N_20434,N_20762);
or U24385 (N_24385,N_20031,N_21565);
nand U24386 (N_24386,N_21293,N_22133);
or U24387 (N_24387,N_20698,N_21049);
nand U24388 (N_24388,N_20620,N_20168);
nor U24389 (N_24389,N_21458,N_21488);
nor U24390 (N_24390,N_20893,N_21780);
nor U24391 (N_24391,N_20112,N_21769);
and U24392 (N_24392,N_20607,N_21093);
xnor U24393 (N_24393,N_22317,N_21786);
or U24394 (N_24394,N_22242,N_20367);
nor U24395 (N_24395,N_21018,N_21423);
nand U24396 (N_24396,N_21510,N_20663);
or U24397 (N_24397,N_22091,N_21008);
nand U24398 (N_24398,N_20099,N_22171);
nand U24399 (N_24399,N_22345,N_22355);
and U24400 (N_24400,N_21996,N_21255);
or U24401 (N_24401,N_20960,N_20337);
nor U24402 (N_24402,N_21888,N_21884);
nand U24403 (N_24403,N_20799,N_20882);
and U24404 (N_24404,N_22003,N_20149);
or U24405 (N_24405,N_21523,N_20045);
or U24406 (N_24406,N_21537,N_21695);
nand U24407 (N_24407,N_21387,N_20184);
or U24408 (N_24408,N_20292,N_20328);
nand U24409 (N_24409,N_21803,N_20331);
nor U24410 (N_24410,N_21127,N_22203);
nor U24411 (N_24411,N_20798,N_21144);
or U24412 (N_24412,N_20919,N_21655);
and U24413 (N_24413,N_21475,N_21332);
or U24414 (N_24414,N_21386,N_20716);
nor U24415 (N_24415,N_20025,N_20759);
and U24416 (N_24416,N_22406,N_20323);
or U24417 (N_24417,N_20582,N_20051);
nor U24418 (N_24418,N_20222,N_20632);
nor U24419 (N_24419,N_21759,N_20198);
nor U24420 (N_24420,N_21699,N_20850);
nand U24421 (N_24421,N_21015,N_22400);
nor U24422 (N_24422,N_22134,N_22290);
and U24423 (N_24423,N_21741,N_22038);
and U24424 (N_24424,N_22202,N_20133);
or U24425 (N_24425,N_21580,N_20417);
nor U24426 (N_24426,N_22185,N_20653);
or U24427 (N_24427,N_22075,N_20357);
or U24428 (N_24428,N_20528,N_21191);
nor U24429 (N_24429,N_20098,N_22305);
nor U24430 (N_24430,N_20699,N_21081);
nor U24431 (N_24431,N_20008,N_21151);
and U24432 (N_24432,N_20380,N_21207);
and U24433 (N_24433,N_21975,N_21137);
or U24434 (N_24434,N_21807,N_20127);
nand U24435 (N_24435,N_21293,N_20195);
nand U24436 (N_24436,N_21153,N_21347);
nor U24437 (N_24437,N_21338,N_22096);
nand U24438 (N_24438,N_22393,N_21405);
and U24439 (N_24439,N_21410,N_22129);
nand U24440 (N_24440,N_22072,N_20874);
and U24441 (N_24441,N_21564,N_21335);
and U24442 (N_24442,N_20631,N_22099);
or U24443 (N_24443,N_20569,N_22258);
and U24444 (N_24444,N_20704,N_20517);
nand U24445 (N_24445,N_20862,N_22279);
or U24446 (N_24446,N_22168,N_22205);
nand U24447 (N_24447,N_21998,N_21810);
or U24448 (N_24448,N_21569,N_22329);
nor U24449 (N_24449,N_20829,N_20280);
nand U24450 (N_24450,N_22435,N_20499);
and U24451 (N_24451,N_21981,N_20093);
and U24452 (N_24452,N_22139,N_20233);
nand U24453 (N_24453,N_21604,N_20177);
nand U24454 (N_24454,N_21714,N_20646);
or U24455 (N_24455,N_21680,N_22137);
nor U24456 (N_24456,N_21084,N_20911);
nand U24457 (N_24457,N_22253,N_21515);
and U24458 (N_24458,N_20416,N_20131);
nand U24459 (N_24459,N_21486,N_22483);
nor U24460 (N_24460,N_20935,N_22371);
and U24461 (N_24461,N_21889,N_21166);
nor U24462 (N_24462,N_21131,N_21160);
nor U24463 (N_24463,N_20903,N_20041);
nor U24464 (N_24464,N_21241,N_21532);
and U24465 (N_24465,N_20201,N_20271);
or U24466 (N_24466,N_20286,N_22163);
and U24467 (N_24467,N_21236,N_20834);
nand U24468 (N_24468,N_20505,N_22300);
or U24469 (N_24469,N_21816,N_21251);
nand U24470 (N_24470,N_21350,N_21241);
nor U24471 (N_24471,N_21730,N_20664);
xor U24472 (N_24472,N_21437,N_20815);
and U24473 (N_24473,N_21077,N_21129);
or U24474 (N_24474,N_21553,N_20776);
nand U24475 (N_24475,N_22485,N_22280);
nor U24476 (N_24476,N_20226,N_21982);
or U24477 (N_24477,N_21446,N_21876);
or U24478 (N_24478,N_20099,N_20226);
or U24479 (N_24479,N_20854,N_21971);
or U24480 (N_24480,N_20624,N_21036);
nor U24481 (N_24481,N_22308,N_21526);
nor U24482 (N_24482,N_20743,N_21216);
and U24483 (N_24483,N_20285,N_21826);
and U24484 (N_24484,N_20934,N_22437);
nor U24485 (N_24485,N_20219,N_21445);
nand U24486 (N_24486,N_20463,N_20073);
and U24487 (N_24487,N_21395,N_21377);
nand U24488 (N_24488,N_22085,N_20599);
nor U24489 (N_24489,N_20162,N_21701);
nand U24490 (N_24490,N_22453,N_22160);
and U24491 (N_24491,N_20598,N_22129);
nand U24492 (N_24492,N_21531,N_21618);
nor U24493 (N_24493,N_20154,N_21924);
nor U24494 (N_24494,N_21716,N_20552);
nand U24495 (N_24495,N_21207,N_20523);
and U24496 (N_24496,N_21092,N_20167);
nand U24497 (N_24497,N_20628,N_20673);
and U24498 (N_24498,N_21904,N_22444);
or U24499 (N_24499,N_21787,N_20072);
or U24500 (N_24500,N_20224,N_20043);
nand U24501 (N_24501,N_21925,N_22421);
nand U24502 (N_24502,N_21426,N_21772);
or U24503 (N_24503,N_20755,N_22491);
nor U24504 (N_24504,N_21313,N_20416);
or U24505 (N_24505,N_20894,N_20154);
or U24506 (N_24506,N_20407,N_20247);
and U24507 (N_24507,N_21720,N_20128);
nor U24508 (N_24508,N_21602,N_20036);
nand U24509 (N_24509,N_20616,N_22090);
nand U24510 (N_24510,N_22090,N_20403);
and U24511 (N_24511,N_21365,N_20846);
nor U24512 (N_24512,N_22218,N_20923);
nand U24513 (N_24513,N_21495,N_22435);
nand U24514 (N_24514,N_21339,N_22041);
nand U24515 (N_24515,N_22432,N_21752);
nand U24516 (N_24516,N_20563,N_22068);
nand U24517 (N_24517,N_20252,N_20403);
nand U24518 (N_24518,N_21608,N_21085);
nor U24519 (N_24519,N_22193,N_20245);
and U24520 (N_24520,N_20297,N_21401);
and U24521 (N_24521,N_20082,N_21614);
nor U24522 (N_24522,N_22496,N_20326);
and U24523 (N_24523,N_22181,N_20576);
and U24524 (N_24524,N_20901,N_22009);
or U24525 (N_24525,N_20054,N_20087);
nand U24526 (N_24526,N_20626,N_21811);
nand U24527 (N_24527,N_21950,N_22275);
and U24528 (N_24528,N_21114,N_22390);
nor U24529 (N_24529,N_21481,N_22104);
or U24530 (N_24530,N_20616,N_20190);
and U24531 (N_24531,N_22248,N_20654);
or U24532 (N_24532,N_20693,N_20508);
or U24533 (N_24533,N_22342,N_21981);
or U24534 (N_24534,N_20048,N_22360);
nand U24535 (N_24535,N_20951,N_21264);
and U24536 (N_24536,N_22400,N_22054);
nor U24537 (N_24537,N_21719,N_21744);
and U24538 (N_24538,N_21673,N_20085);
or U24539 (N_24539,N_22081,N_21022);
nor U24540 (N_24540,N_20658,N_21680);
nand U24541 (N_24541,N_22329,N_22459);
nand U24542 (N_24542,N_21229,N_22083);
nand U24543 (N_24543,N_21563,N_21355);
or U24544 (N_24544,N_22187,N_21925);
nand U24545 (N_24545,N_21349,N_20779);
and U24546 (N_24546,N_20330,N_20744);
or U24547 (N_24547,N_21772,N_21976);
or U24548 (N_24548,N_20499,N_22056);
nor U24549 (N_24549,N_22484,N_21094);
or U24550 (N_24550,N_20545,N_20763);
nor U24551 (N_24551,N_20131,N_21062);
and U24552 (N_24552,N_22415,N_20836);
or U24553 (N_24553,N_20348,N_21134);
nor U24554 (N_24554,N_21455,N_20494);
or U24555 (N_24555,N_22095,N_21659);
nor U24556 (N_24556,N_22365,N_21385);
nor U24557 (N_24557,N_22288,N_20379);
and U24558 (N_24558,N_20813,N_22065);
xor U24559 (N_24559,N_22274,N_21497);
or U24560 (N_24560,N_21931,N_20686);
nand U24561 (N_24561,N_20474,N_20540);
and U24562 (N_24562,N_21581,N_20281);
nand U24563 (N_24563,N_21345,N_21923);
and U24564 (N_24564,N_20354,N_21520);
and U24565 (N_24565,N_22473,N_21615);
nand U24566 (N_24566,N_21693,N_22314);
and U24567 (N_24567,N_20589,N_22141);
nor U24568 (N_24568,N_21883,N_20730);
or U24569 (N_24569,N_21077,N_21220);
or U24570 (N_24570,N_20981,N_20371);
or U24571 (N_24571,N_21845,N_21917);
nor U24572 (N_24572,N_21916,N_21009);
nor U24573 (N_24573,N_21973,N_20254);
or U24574 (N_24574,N_21053,N_20805);
or U24575 (N_24575,N_22248,N_21940);
or U24576 (N_24576,N_20609,N_22266);
or U24577 (N_24577,N_21093,N_20054);
or U24578 (N_24578,N_22359,N_21516);
nor U24579 (N_24579,N_20071,N_21742);
nor U24580 (N_24580,N_20495,N_22183);
nor U24581 (N_24581,N_22341,N_21244);
and U24582 (N_24582,N_22134,N_21499);
nand U24583 (N_24583,N_20870,N_22336);
and U24584 (N_24584,N_20204,N_20389);
nor U24585 (N_24585,N_20823,N_22332);
nor U24586 (N_24586,N_20658,N_21681);
xnor U24587 (N_24587,N_22488,N_20570);
and U24588 (N_24588,N_20546,N_22253);
or U24589 (N_24589,N_21232,N_20221);
and U24590 (N_24590,N_20256,N_20093);
and U24591 (N_24591,N_21173,N_21395);
or U24592 (N_24592,N_20954,N_20339);
nand U24593 (N_24593,N_22038,N_20401);
nand U24594 (N_24594,N_21956,N_22215);
or U24595 (N_24595,N_21535,N_20869);
or U24596 (N_24596,N_20305,N_21296);
nand U24597 (N_24597,N_20750,N_20029);
and U24598 (N_24598,N_21195,N_20064);
nor U24599 (N_24599,N_20241,N_20579);
and U24600 (N_24600,N_22078,N_21210);
nor U24601 (N_24601,N_20911,N_21843);
nand U24602 (N_24602,N_21962,N_21254);
nor U24603 (N_24603,N_21646,N_20694);
nor U24604 (N_24604,N_21772,N_22160);
nand U24605 (N_24605,N_21576,N_22220);
nand U24606 (N_24606,N_21903,N_22437);
nand U24607 (N_24607,N_21833,N_20836);
and U24608 (N_24608,N_21733,N_21665);
nor U24609 (N_24609,N_21845,N_21937);
and U24610 (N_24610,N_20120,N_21757);
or U24611 (N_24611,N_21051,N_21442);
or U24612 (N_24612,N_21706,N_22048);
and U24613 (N_24613,N_22288,N_22153);
and U24614 (N_24614,N_22128,N_20169);
and U24615 (N_24615,N_22235,N_20119);
and U24616 (N_24616,N_20842,N_20530);
and U24617 (N_24617,N_20806,N_20989);
or U24618 (N_24618,N_21883,N_20169);
or U24619 (N_24619,N_21978,N_21007);
nand U24620 (N_24620,N_22190,N_21878);
or U24621 (N_24621,N_20591,N_20426);
nor U24622 (N_24622,N_21340,N_22025);
and U24623 (N_24623,N_21818,N_20024);
or U24624 (N_24624,N_20614,N_21575);
and U24625 (N_24625,N_20872,N_22315);
and U24626 (N_24626,N_22176,N_20153);
nor U24627 (N_24627,N_21142,N_22031);
nor U24628 (N_24628,N_21260,N_20593);
nand U24629 (N_24629,N_21246,N_20735);
and U24630 (N_24630,N_21939,N_20409);
nand U24631 (N_24631,N_22139,N_20768);
and U24632 (N_24632,N_20846,N_22467);
nor U24633 (N_24633,N_22037,N_21096);
and U24634 (N_24634,N_21232,N_20761);
nand U24635 (N_24635,N_20098,N_22166);
and U24636 (N_24636,N_20036,N_20713);
nand U24637 (N_24637,N_20497,N_21875);
or U24638 (N_24638,N_21481,N_20655);
nor U24639 (N_24639,N_20552,N_20482);
nor U24640 (N_24640,N_21886,N_20125);
and U24641 (N_24641,N_21595,N_20779);
nand U24642 (N_24642,N_21450,N_20098);
and U24643 (N_24643,N_20778,N_21465);
and U24644 (N_24644,N_21245,N_22319);
nor U24645 (N_24645,N_21197,N_20583);
or U24646 (N_24646,N_21518,N_21564);
nand U24647 (N_24647,N_20401,N_20894);
or U24648 (N_24648,N_20426,N_20744);
or U24649 (N_24649,N_20575,N_20866);
nand U24650 (N_24650,N_22260,N_20819);
or U24651 (N_24651,N_21842,N_21928);
nor U24652 (N_24652,N_22487,N_20287);
and U24653 (N_24653,N_21410,N_21200);
nor U24654 (N_24654,N_20662,N_20548);
or U24655 (N_24655,N_22276,N_20365);
or U24656 (N_24656,N_20744,N_20627);
xor U24657 (N_24657,N_20762,N_20055);
or U24658 (N_24658,N_21283,N_20547);
and U24659 (N_24659,N_22039,N_20240);
nand U24660 (N_24660,N_22076,N_21971);
or U24661 (N_24661,N_20145,N_20611);
nand U24662 (N_24662,N_22136,N_20318);
or U24663 (N_24663,N_21462,N_21657);
or U24664 (N_24664,N_22331,N_22114);
nand U24665 (N_24665,N_21542,N_20419);
nand U24666 (N_24666,N_21263,N_21959);
nor U24667 (N_24667,N_20185,N_22142);
or U24668 (N_24668,N_22047,N_20236);
or U24669 (N_24669,N_20322,N_20412);
nor U24670 (N_24670,N_20476,N_22400);
and U24671 (N_24671,N_21494,N_20204);
or U24672 (N_24672,N_21662,N_22195);
nand U24673 (N_24673,N_21782,N_21415);
and U24674 (N_24674,N_21625,N_21951);
nand U24675 (N_24675,N_22287,N_21805);
nor U24676 (N_24676,N_21094,N_21826);
nor U24677 (N_24677,N_20295,N_20140);
nor U24678 (N_24678,N_22241,N_22036);
or U24679 (N_24679,N_21374,N_21412);
and U24680 (N_24680,N_20391,N_20069);
and U24681 (N_24681,N_21377,N_20114);
nand U24682 (N_24682,N_22492,N_22212);
nand U24683 (N_24683,N_20167,N_21532);
and U24684 (N_24684,N_20566,N_22404);
or U24685 (N_24685,N_21250,N_20325);
nand U24686 (N_24686,N_21618,N_21352);
and U24687 (N_24687,N_22374,N_21843);
or U24688 (N_24688,N_21953,N_22312);
nand U24689 (N_24689,N_20309,N_21593);
nand U24690 (N_24690,N_20511,N_21097);
or U24691 (N_24691,N_21320,N_20362);
nand U24692 (N_24692,N_22104,N_22065);
or U24693 (N_24693,N_21763,N_21032);
nand U24694 (N_24694,N_21415,N_21984);
and U24695 (N_24695,N_20710,N_21921);
or U24696 (N_24696,N_21940,N_20118);
nor U24697 (N_24697,N_21920,N_22465);
nor U24698 (N_24698,N_20033,N_21167);
nor U24699 (N_24699,N_21660,N_20331);
nand U24700 (N_24700,N_21185,N_20695);
and U24701 (N_24701,N_21408,N_22437);
nand U24702 (N_24702,N_20151,N_22016);
nand U24703 (N_24703,N_20574,N_20572);
and U24704 (N_24704,N_20079,N_21624);
and U24705 (N_24705,N_21485,N_21269);
nand U24706 (N_24706,N_21964,N_20357);
nor U24707 (N_24707,N_21684,N_22136);
nor U24708 (N_24708,N_22039,N_22274);
nor U24709 (N_24709,N_22413,N_22150);
and U24710 (N_24710,N_22448,N_21813);
nor U24711 (N_24711,N_20192,N_22247);
and U24712 (N_24712,N_20619,N_20804);
and U24713 (N_24713,N_22229,N_20361);
or U24714 (N_24714,N_20522,N_20051);
and U24715 (N_24715,N_21415,N_20352);
and U24716 (N_24716,N_22202,N_20235);
or U24717 (N_24717,N_20041,N_22262);
or U24718 (N_24718,N_21009,N_22342);
and U24719 (N_24719,N_21030,N_22499);
nor U24720 (N_24720,N_22421,N_21515);
or U24721 (N_24721,N_20757,N_21780);
nor U24722 (N_24722,N_20506,N_20629);
nand U24723 (N_24723,N_21065,N_20104);
nor U24724 (N_24724,N_20832,N_20261);
and U24725 (N_24725,N_21316,N_20373);
or U24726 (N_24726,N_20032,N_22249);
and U24727 (N_24727,N_21961,N_20579);
nor U24728 (N_24728,N_22334,N_21482);
and U24729 (N_24729,N_21229,N_20584);
or U24730 (N_24730,N_21320,N_21269);
nor U24731 (N_24731,N_20722,N_20007);
or U24732 (N_24732,N_20124,N_20768);
nor U24733 (N_24733,N_21893,N_21467);
nor U24734 (N_24734,N_21660,N_20100);
nand U24735 (N_24735,N_22061,N_20829);
nand U24736 (N_24736,N_21851,N_21345);
or U24737 (N_24737,N_20794,N_21458);
nor U24738 (N_24738,N_20756,N_20372);
and U24739 (N_24739,N_21804,N_20623);
and U24740 (N_24740,N_21067,N_22117);
nor U24741 (N_24741,N_20202,N_21411);
or U24742 (N_24742,N_20609,N_20058);
nand U24743 (N_24743,N_21263,N_22107);
nand U24744 (N_24744,N_22472,N_20872);
and U24745 (N_24745,N_22308,N_21475);
nand U24746 (N_24746,N_22010,N_22475);
and U24747 (N_24747,N_20180,N_20074);
and U24748 (N_24748,N_22282,N_22062);
nand U24749 (N_24749,N_21325,N_21926);
and U24750 (N_24750,N_20460,N_20999);
nor U24751 (N_24751,N_20698,N_21948);
nand U24752 (N_24752,N_20734,N_22410);
nand U24753 (N_24753,N_21117,N_21460);
nor U24754 (N_24754,N_20762,N_21338);
nand U24755 (N_24755,N_21500,N_21587);
or U24756 (N_24756,N_20059,N_20792);
nand U24757 (N_24757,N_22393,N_21731);
nand U24758 (N_24758,N_20057,N_22485);
or U24759 (N_24759,N_22023,N_20535);
xnor U24760 (N_24760,N_21079,N_21493);
nor U24761 (N_24761,N_20137,N_20917);
or U24762 (N_24762,N_20727,N_20522);
or U24763 (N_24763,N_20574,N_20293);
or U24764 (N_24764,N_21850,N_22495);
nand U24765 (N_24765,N_21735,N_20724);
nor U24766 (N_24766,N_20341,N_20700);
and U24767 (N_24767,N_20241,N_22335);
nand U24768 (N_24768,N_22037,N_20380);
and U24769 (N_24769,N_20949,N_20646);
or U24770 (N_24770,N_21120,N_22387);
nor U24771 (N_24771,N_20311,N_20698);
nand U24772 (N_24772,N_21583,N_22451);
nor U24773 (N_24773,N_21435,N_20193);
nand U24774 (N_24774,N_22224,N_22326);
and U24775 (N_24775,N_20963,N_20509);
nand U24776 (N_24776,N_21302,N_22192);
and U24777 (N_24777,N_20136,N_22261);
nor U24778 (N_24778,N_21020,N_22265);
and U24779 (N_24779,N_22196,N_21497);
and U24780 (N_24780,N_20760,N_21237);
and U24781 (N_24781,N_20963,N_20159);
or U24782 (N_24782,N_20431,N_20420);
nor U24783 (N_24783,N_21594,N_21691);
nand U24784 (N_24784,N_21298,N_20839);
or U24785 (N_24785,N_21890,N_22417);
or U24786 (N_24786,N_20137,N_21219);
nor U24787 (N_24787,N_20642,N_20094);
and U24788 (N_24788,N_21660,N_21332);
and U24789 (N_24789,N_21454,N_21533);
and U24790 (N_24790,N_20183,N_22238);
and U24791 (N_24791,N_22327,N_20185);
or U24792 (N_24792,N_20533,N_20555);
nand U24793 (N_24793,N_21035,N_22422);
and U24794 (N_24794,N_20420,N_21481);
nor U24795 (N_24795,N_20119,N_22380);
nand U24796 (N_24796,N_22309,N_21769);
or U24797 (N_24797,N_21695,N_21896);
and U24798 (N_24798,N_21065,N_22235);
or U24799 (N_24799,N_21273,N_21286);
nand U24800 (N_24800,N_22300,N_21431);
nor U24801 (N_24801,N_20645,N_22272);
and U24802 (N_24802,N_22320,N_20940);
and U24803 (N_24803,N_22388,N_20018);
nand U24804 (N_24804,N_21874,N_22480);
xor U24805 (N_24805,N_21737,N_22332);
or U24806 (N_24806,N_21632,N_20388);
and U24807 (N_24807,N_20558,N_22340);
and U24808 (N_24808,N_21205,N_21362);
or U24809 (N_24809,N_20558,N_22226);
and U24810 (N_24810,N_21600,N_22168);
nand U24811 (N_24811,N_21475,N_20215);
or U24812 (N_24812,N_21893,N_21059);
and U24813 (N_24813,N_20997,N_20473);
or U24814 (N_24814,N_22128,N_21371);
and U24815 (N_24815,N_21061,N_21410);
and U24816 (N_24816,N_20363,N_21786);
and U24817 (N_24817,N_20451,N_21841);
and U24818 (N_24818,N_22016,N_22362);
nand U24819 (N_24819,N_22022,N_20812);
and U24820 (N_24820,N_21397,N_20430);
nor U24821 (N_24821,N_20510,N_20868);
or U24822 (N_24822,N_21178,N_21504);
and U24823 (N_24823,N_20079,N_21622);
or U24824 (N_24824,N_21295,N_22107);
or U24825 (N_24825,N_20527,N_21419);
nor U24826 (N_24826,N_20785,N_22314);
and U24827 (N_24827,N_20288,N_20457);
or U24828 (N_24828,N_21792,N_21544);
and U24829 (N_24829,N_21767,N_20719);
xnor U24830 (N_24830,N_20905,N_21494);
nand U24831 (N_24831,N_22381,N_20963);
nand U24832 (N_24832,N_20853,N_22158);
or U24833 (N_24833,N_20121,N_21166);
nand U24834 (N_24834,N_21751,N_20066);
or U24835 (N_24835,N_21177,N_21049);
and U24836 (N_24836,N_20109,N_21726);
and U24837 (N_24837,N_21126,N_21080);
nand U24838 (N_24838,N_22345,N_21751);
nand U24839 (N_24839,N_21248,N_21199);
and U24840 (N_24840,N_20121,N_20884);
or U24841 (N_24841,N_20005,N_20632);
nor U24842 (N_24842,N_22282,N_21248);
nor U24843 (N_24843,N_21163,N_21135);
or U24844 (N_24844,N_21744,N_20232);
or U24845 (N_24845,N_21630,N_20714);
nor U24846 (N_24846,N_20789,N_20725);
nor U24847 (N_24847,N_21349,N_20108);
nand U24848 (N_24848,N_22481,N_20530);
and U24849 (N_24849,N_20179,N_21904);
and U24850 (N_24850,N_22455,N_20447);
nor U24851 (N_24851,N_20136,N_22035);
nand U24852 (N_24852,N_21361,N_21938);
and U24853 (N_24853,N_21989,N_22328);
nand U24854 (N_24854,N_22008,N_21777);
or U24855 (N_24855,N_20852,N_21960);
and U24856 (N_24856,N_21621,N_21587);
and U24857 (N_24857,N_22110,N_21367);
or U24858 (N_24858,N_20511,N_21627);
nor U24859 (N_24859,N_20157,N_20531);
nor U24860 (N_24860,N_21108,N_22392);
and U24861 (N_24861,N_22090,N_21488);
and U24862 (N_24862,N_22204,N_22303);
nor U24863 (N_24863,N_20224,N_22471);
nor U24864 (N_24864,N_21688,N_20551);
or U24865 (N_24865,N_20213,N_20351);
and U24866 (N_24866,N_21422,N_20851);
and U24867 (N_24867,N_20918,N_21627);
and U24868 (N_24868,N_20005,N_21384);
nand U24869 (N_24869,N_22377,N_20256);
nand U24870 (N_24870,N_20085,N_22281);
and U24871 (N_24871,N_21942,N_22460);
nand U24872 (N_24872,N_20945,N_21215);
nor U24873 (N_24873,N_20951,N_20921);
nor U24874 (N_24874,N_22018,N_21689);
and U24875 (N_24875,N_21898,N_22137);
xor U24876 (N_24876,N_21267,N_22093);
nand U24877 (N_24877,N_21394,N_22099);
or U24878 (N_24878,N_20947,N_20702);
or U24879 (N_24879,N_20071,N_22354);
nor U24880 (N_24880,N_21547,N_20729);
and U24881 (N_24881,N_20705,N_20257);
or U24882 (N_24882,N_20038,N_20141);
nor U24883 (N_24883,N_22206,N_20961);
or U24884 (N_24884,N_21240,N_21120);
and U24885 (N_24885,N_20731,N_22295);
or U24886 (N_24886,N_21660,N_22133);
nand U24887 (N_24887,N_21976,N_20014);
or U24888 (N_24888,N_20720,N_21100);
and U24889 (N_24889,N_20438,N_22483);
nand U24890 (N_24890,N_22436,N_20630);
and U24891 (N_24891,N_21003,N_22250);
and U24892 (N_24892,N_20890,N_21736);
and U24893 (N_24893,N_21117,N_20753);
and U24894 (N_24894,N_21490,N_20918);
nor U24895 (N_24895,N_20284,N_21693);
nor U24896 (N_24896,N_21815,N_22244);
and U24897 (N_24897,N_21813,N_22354);
nand U24898 (N_24898,N_22221,N_20641);
nor U24899 (N_24899,N_20902,N_22341);
nor U24900 (N_24900,N_21805,N_20614);
nand U24901 (N_24901,N_22091,N_21052);
or U24902 (N_24902,N_20694,N_20570);
nand U24903 (N_24903,N_20522,N_20684);
and U24904 (N_24904,N_20058,N_22481);
or U24905 (N_24905,N_21845,N_22333);
nor U24906 (N_24906,N_22170,N_21332);
and U24907 (N_24907,N_22251,N_21238);
nor U24908 (N_24908,N_21650,N_20773);
or U24909 (N_24909,N_20471,N_21259);
nand U24910 (N_24910,N_20047,N_20433);
and U24911 (N_24911,N_20007,N_21902);
nor U24912 (N_24912,N_20179,N_20403);
and U24913 (N_24913,N_21280,N_20999);
nor U24914 (N_24914,N_22233,N_21580);
or U24915 (N_24915,N_20222,N_20928);
or U24916 (N_24916,N_21030,N_22239);
and U24917 (N_24917,N_20046,N_20901);
nand U24918 (N_24918,N_20389,N_20494);
nor U24919 (N_24919,N_22164,N_20789);
nand U24920 (N_24920,N_20337,N_20284);
or U24921 (N_24921,N_22373,N_20279);
and U24922 (N_24922,N_22481,N_21150);
or U24923 (N_24923,N_20448,N_22473);
nand U24924 (N_24924,N_22296,N_22114);
nor U24925 (N_24925,N_21058,N_21840);
and U24926 (N_24926,N_21236,N_22213);
or U24927 (N_24927,N_21917,N_22030);
or U24928 (N_24928,N_22452,N_20669);
nand U24929 (N_24929,N_21368,N_21413);
nand U24930 (N_24930,N_20749,N_22468);
and U24931 (N_24931,N_21309,N_21407);
nand U24932 (N_24932,N_20786,N_21666);
nand U24933 (N_24933,N_21510,N_21599);
nand U24934 (N_24934,N_20955,N_21049);
nor U24935 (N_24935,N_22176,N_20838);
nand U24936 (N_24936,N_22280,N_22430);
nor U24937 (N_24937,N_22292,N_20756);
nor U24938 (N_24938,N_20635,N_20417);
or U24939 (N_24939,N_21316,N_20949);
nand U24940 (N_24940,N_22051,N_22035);
or U24941 (N_24941,N_22134,N_20627);
nor U24942 (N_24942,N_22088,N_21801);
or U24943 (N_24943,N_20053,N_21996);
or U24944 (N_24944,N_20485,N_20010);
and U24945 (N_24945,N_20600,N_21904);
nor U24946 (N_24946,N_21813,N_21543);
and U24947 (N_24947,N_20341,N_20396);
or U24948 (N_24948,N_20076,N_21277);
nor U24949 (N_24949,N_20378,N_20545);
nor U24950 (N_24950,N_21177,N_21446);
nand U24951 (N_24951,N_21532,N_20944);
and U24952 (N_24952,N_20118,N_20109);
or U24953 (N_24953,N_21496,N_21940);
or U24954 (N_24954,N_21482,N_20612);
and U24955 (N_24955,N_21244,N_22062);
or U24956 (N_24956,N_22307,N_21200);
and U24957 (N_24957,N_21684,N_21937);
or U24958 (N_24958,N_21823,N_20318);
nor U24959 (N_24959,N_20926,N_20965);
nand U24960 (N_24960,N_20369,N_21223);
nand U24961 (N_24961,N_20451,N_22048);
nand U24962 (N_24962,N_20412,N_20240);
xnor U24963 (N_24963,N_20373,N_21954);
nand U24964 (N_24964,N_21804,N_20870);
nor U24965 (N_24965,N_20780,N_20064);
and U24966 (N_24966,N_22360,N_21872);
or U24967 (N_24967,N_21602,N_20783);
or U24968 (N_24968,N_20728,N_21172);
or U24969 (N_24969,N_20922,N_20481);
and U24970 (N_24970,N_20552,N_22298);
and U24971 (N_24971,N_21528,N_20895);
or U24972 (N_24972,N_20179,N_20902);
nor U24973 (N_24973,N_21104,N_20781);
or U24974 (N_24974,N_22210,N_21993);
nand U24975 (N_24975,N_20167,N_22207);
or U24976 (N_24976,N_21855,N_20290);
or U24977 (N_24977,N_21270,N_20993);
and U24978 (N_24978,N_21413,N_20800);
or U24979 (N_24979,N_20906,N_22492);
nand U24980 (N_24980,N_21462,N_20802);
nand U24981 (N_24981,N_21909,N_20672);
nor U24982 (N_24982,N_21976,N_21993);
and U24983 (N_24983,N_21597,N_21179);
nor U24984 (N_24984,N_22361,N_21416);
nand U24985 (N_24985,N_20292,N_20327);
nor U24986 (N_24986,N_21880,N_20661);
nor U24987 (N_24987,N_21510,N_21894);
nor U24988 (N_24988,N_21073,N_22251);
nor U24989 (N_24989,N_21946,N_20872);
nand U24990 (N_24990,N_20352,N_22025);
and U24991 (N_24991,N_22441,N_21213);
and U24992 (N_24992,N_22052,N_20907);
or U24993 (N_24993,N_22467,N_21338);
nor U24994 (N_24994,N_21079,N_21625);
nor U24995 (N_24995,N_20333,N_20956);
or U24996 (N_24996,N_21724,N_22413);
and U24997 (N_24997,N_22228,N_20317);
nand U24998 (N_24998,N_20829,N_20222);
nor U24999 (N_24999,N_21127,N_20742);
nand UO_0 (O_0,N_22839,N_23442);
and UO_1 (O_1,N_23460,N_23778);
or UO_2 (O_2,N_24015,N_24115);
or UO_3 (O_3,N_22502,N_24507);
nand UO_4 (O_4,N_23530,N_23286);
and UO_5 (O_5,N_23779,N_24354);
nand UO_6 (O_6,N_24261,N_23647);
nor UO_7 (O_7,N_23316,N_24135);
nor UO_8 (O_8,N_24552,N_23449);
nand UO_9 (O_9,N_24240,N_24383);
or UO_10 (O_10,N_23043,N_22773);
nor UO_11 (O_11,N_23477,N_22876);
nand UO_12 (O_12,N_23904,N_22826);
and UO_13 (O_13,N_22781,N_24230);
and UO_14 (O_14,N_24620,N_24708);
or UO_15 (O_15,N_24503,N_24168);
or UO_16 (O_16,N_23083,N_23329);
or UO_17 (O_17,N_23894,N_24066);
or UO_18 (O_18,N_22527,N_24361);
or UO_19 (O_19,N_22565,N_23932);
and UO_20 (O_20,N_24975,N_23057);
and UO_21 (O_21,N_23523,N_24526);
or UO_22 (O_22,N_24497,N_24282);
and UO_23 (O_23,N_24810,N_23721);
and UO_24 (O_24,N_24114,N_24273);
nand UO_25 (O_25,N_24349,N_23342);
nor UO_26 (O_26,N_24903,N_24221);
nand UO_27 (O_27,N_22886,N_24757);
nor UO_28 (O_28,N_24428,N_24622);
or UO_29 (O_29,N_23405,N_24625);
nor UO_30 (O_30,N_24921,N_23123);
nand UO_31 (O_31,N_22637,N_23787);
and UO_32 (O_32,N_24938,N_23609);
and UO_33 (O_33,N_22896,N_22512);
nand UO_34 (O_34,N_22589,N_24063);
nor UO_35 (O_35,N_24642,N_24953);
nor UO_36 (O_36,N_23989,N_24351);
xor UO_37 (O_37,N_23847,N_22847);
or UO_38 (O_38,N_22689,N_23125);
nand UO_39 (O_39,N_23545,N_24774);
nand UO_40 (O_40,N_23351,N_24889);
nand UO_41 (O_41,N_23438,N_24659);
nor UO_42 (O_42,N_24617,N_23914);
and UO_43 (O_43,N_23614,N_24485);
nand UO_44 (O_44,N_22966,N_23980);
nor UO_45 (O_45,N_22842,N_23168);
and UO_46 (O_46,N_23106,N_22569);
or UO_47 (O_47,N_24258,N_22771);
and UO_48 (O_48,N_24731,N_24974);
or UO_49 (O_49,N_24170,N_23754);
nand UO_50 (O_50,N_23866,N_22718);
nand UO_51 (O_51,N_22632,N_23166);
nand UO_52 (O_52,N_23469,N_24207);
or UO_53 (O_53,N_23134,N_22756);
nor UO_54 (O_54,N_24246,N_23941);
xnor UO_55 (O_55,N_24250,N_24236);
and UO_56 (O_56,N_23666,N_24465);
and UO_57 (O_57,N_24105,N_24064);
nor UO_58 (O_58,N_23875,N_24884);
nand UO_59 (O_59,N_24068,N_23433);
nor UO_60 (O_60,N_24329,N_22529);
or UO_61 (O_61,N_23455,N_24511);
and UO_62 (O_62,N_23317,N_24430);
nand UO_63 (O_63,N_23985,N_24618);
or UO_64 (O_64,N_23293,N_23148);
nor UO_65 (O_65,N_22892,N_22963);
or UO_66 (O_66,N_23312,N_24054);
nand UO_67 (O_67,N_24188,N_23174);
nor UO_68 (O_68,N_24784,N_24123);
and UO_69 (O_69,N_22938,N_24101);
nand UO_70 (O_70,N_24277,N_23809);
and UO_71 (O_71,N_23885,N_23256);
or UO_72 (O_72,N_24893,N_23745);
and UO_73 (O_73,N_22902,N_23384);
and UO_74 (O_74,N_22812,N_22526);
or UO_75 (O_75,N_24519,N_24256);
nor UO_76 (O_76,N_24720,N_24461);
nor UO_77 (O_77,N_24022,N_23109);
nor UO_78 (O_78,N_24514,N_23473);
nor UO_79 (O_79,N_24513,N_24588);
nor UO_80 (O_80,N_24728,N_23390);
or UO_81 (O_81,N_23430,N_22647);
and UO_82 (O_82,N_24646,N_24786);
nand UO_83 (O_83,N_24152,N_22720);
or UO_84 (O_84,N_24594,N_23295);
and UO_85 (O_85,N_24881,N_24819);
nor UO_86 (O_86,N_23300,N_24451);
and UO_87 (O_87,N_23600,N_24761);
nor UO_88 (O_88,N_22764,N_23482);
nor UO_89 (O_89,N_24539,N_22926);
and UO_90 (O_90,N_24968,N_24342);
nand UO_91 (O_91,N_23297,N_24362);
nor UO_92 (O_92,N_22624,N_24704);
or UO_93 (O_93,N_23187,N_23006);
and UO_94 (O_94,N_24477,N_22581);
nor UO_95 (O_95,N_24981,N_23465);
or UO_96 (O_96,N_24025,N_22711);
or UO_97 (O_97,N_24865,N_23518);
nand UO_98 (O_98,N_24072,N_23574);
or UO_99 (O_99,N_24885,N_23815);
and UO_100 (O_100,N_23713,N_24689);
and UO_101 (O_101,N_23697,N_24749);
and UO_102 (O_102,N_23284,N_23749);
nor UO_103 (O_103,N_22804,N_22783);
nand UO_104 (O_104,N_22823,N_22753);
nand UO_105 (O_105,N_24472,N_23146);
nor UO_106 (O_106,N_24125,N_22957);
nand UO_107 (O_107,N_22913,N_22878);
or UO_108 (O_108,N_22874,N_22664);
and UO_109 (O_109,N_23507,N_24009);
nand UO_110 (O_110,N_23045,N_22734);
and UO_111 (O_111,N_23004,N_22777);
nor UO_112 (O_112,N_23956,N_24032);
nor UO_113 (O_113,N_23694,N_22815);
or UO_114 (O_114,N_22920,N_24755);
and UO_115 (O_115,N_23436,N_24779);
nor UO_116 (O_116,N_23247,N_24409);
or UO_117 (O_117,N_23893,N_23868);
nor UO_118 (O_118,N_23009,N_24076);
nor UO_119 (O_119,N_22633,N_23192);
and UO_120 (O_120,N_24290,N_24667);
and UO_121 (O_121,N_23539,N_24458);
nor UO_122 (O_122,N_24845,N_24260);
nor UO_123 (O_123,N_23205,N_22542);
nand UO_124 (O_124,N_24883,N_23526);
and UO_125 (O_125,N_23343,N_24565);
nand UO_126 (O_126,N_24281,N_24356);
and UO_127 (O_127,N_23199,N_24510);
or UO_128 (O_128,N_24661,N_24346);
or UO_129 (O_129,N_23828,N_23688);
and UO_130 (O_130,N_22736,N_24985);
nand UO_131 (O_131,N_24946,N_23546);
or UO_132 (O_132,N_23226,N_23493);
nand UO_133 (O_133,N_24426,N_24532);
and UO_134 (O_134,N_22727,N_22610);
and UO_135 (O_135,N_23578,N_24542);
nor UO_136 (O_136,N_23413,N_24644);
or UO_137 (O_137,N_22662,N_23221);
or UO_138 (O_138,N_24099,N_24536);
nand UO_139 (O_139,N_23764,N_24355);
or UO_140 (O_140,N_23997,N_24449);
nor UO_141 (O_141,N_23494,N_23562);
nand UO_142 (O_142,N_24219,N_22821);
or UO_143 (O_143,N_22970,N_24039);
nand UO_144 (O_144,N_24504,N_24665);
nor UO_145 (O_145,N_22803,N_22560);
nand UO_146 (O_146,N_22616,N_24705);
or UO_147 (O_147,N_23726,N_22747);
or UO_148 (O_148,N_23063,N_24190);
or UO_149 (O_149,N_24943,N_22940);
or UO_150 (O_150,N_23008,N_22788);
nor UO_151 (O_151,N_22950,N_24977);
nor UO_152 (O_152,N_24210,N_24994);
nor UO_153 (O_153,N_24827,N_24085);
and UO_154 (O_154,N_22939,N_22574);
and UO_155 (O_155,N_22546,N_23890);
nor UO_156 (O_156,N_23440,N_23037);
nand UO_157 (O_157,N_23087,N_22779);
or UO_158 (O_158,N_22690,N_23102);
and UO_159 (O_159,N_23658,N_22922);
nand UO_160 (O_160,N_22754,N_23708);
and UO_161 (O_161,N_22930,N_24494);
or UO_162 (O_162,N_23266,N_22854);
and UO_163 (O_163,N_24577,N_23039);
nor UO_164 (O_164,N_23097,N_23733);
and UO_165 (O_165,N_24136,N_24529);
or UO_166 (O_166,N_22895,N_24636);
or UO_167 (O_167,N_23085,N_24442);
or UO_168 (O_168,N_24008,N_24991);
nand UO_169 (O_169,N_23068,N_24331);
and UO_170 (O_170,N_24959,N_24386);
nor UO_171 (O_171,N_23821,N_23158);
or UO_172 (O_172,N_24655,N_23521);
and UO_173 (O_173,N_23371,N_24359);
nor UO_174 (O_174,N_23982,N_22983);
and UO_175 (O_175,N_22794,N_22699);
nor UO_176 (O_176,N_24028,N_23589);
or UO_177 (O_177,N_23816,N_23432);
and UO_178 (O_178,N_23865,N_23591);
nand UO_179 (O_179,N_23330,N_24538);
or UO_180 (O_180,N_22873,N_23054);
nand UO_181 (O_181,N_23717,N_23527);
and UO_182 (O_182,N_24487,N_24293);
and UO_183 (O_183,N_22732,N_24723);
or UO_184 (O_184,N_24399,N_22654);
and UO_185 (O_185,N_22918,N_23543);
or UO_186 (O_186,N_23977,N_22620);
nand UO_187 (O_187,N_23558,N_23129);
nor UO_188 (O_188,N_24753,N_24450);
nand UO_189 (O_189,N_23459,N_23281);
nand UO_190 (O_190,N_23595,N_23116);
nand UO_191 (O_191,N_24590,N_24247);
and UO_192 (O_192,N_23217,N_24204);
nand UO_193 (O_193,N_23958,N_22658);
nand UO_194 (O_194,N_23888,N_24264);
xor UO_195 (O_195,N_23800,N_22679);
nor UO_196 (O_196,N_23921,N_24972);
or UO_197 (O_197,N_23775,N_24104);
and UO_198 (O_198,N_23251,N_23711);
nor UO_199 (O_199,N_23328,N_22894);
and UO_200 (O_200,N_24730,N_24651);
nor UO_201 (O_201,N_23567,N_24906);
nor UO_202 (O_202,N_24948,N_22543);
nand UO_203 (O_203,N_24817,N_23499);
nor UO_204 (O_204,N_24295,N_24671);
nor UO_205 (O_205,N_22887,N_23786);
nand UO_206 (O_206,N_22669,N_23916);
nand UO_207 (O_207,N_23246,N_24433);
or UO_208 (O_208,N_24463,N_22937);
or UO_209 (O_209,N_22760,N_23321);
and UO_210 (O_210,N_24806,N_22719);
nor UO_211 (O_211,N_23627,N_24026);
and UO_212 (O_212,N_24815,N_23423);
and UO_213 (O_213,N_24719,N_24111);
or UO_214 (O_214,N_24982,N_24678);
nand UO_215 (O_215,N_23279,N_23783);
nor UO_216 (O_216,N_23684,N_23025);
and UO_217 (O_217,N_24822,N_23065);
nand UO_218 (O_218,N_24910,N_24852);
and UO_219 (O_219,N_24986,N_22622);
nor UO_220 (O_220,N_24058,N_22525);
and UO_221 (O_221,N_23468,N_22671);
and UO_222 (O_222,N_24096,N_24267);
nand UO_223 (O_223,N_23495,N_24838);
and UO_224 (O_224,N_23963,N_22538);
or UO_225 (O_225,N_22712,N_23356);
or UO_226 (O_226,N_24425,N_23796);
or UO_227 (O_227,N_23644,N_23632);
and UO_228 (O_228,N_24711,N_23705);
nor UO_229 (O_229,N_23415,N_24467);
and UO_230 (O_230,N_22717,N_24133);
and UO_231 (O_231,N_23970,N_23502);
or UO_232 (O_232,N_24656,N_22865);
nor UO_233 (O_233,N_24447,N_22776);
nand UO_234 (O_234,N_23616,N_24887);
nand UO_235 (O_235,N_22630,N_22591);
or UO_236 (O_236,N_24189,N_23292);
nor UO_237 (O_237,N_23124,N_23912);
or UO_238 (O_238,N_23793,N_22891);
nand UO_239 (O_239,N_23555,N_23906);
nor UO_240 (O_240,N_23731,N_24375);
nor UO_241 (O_241,N_23664,N_24621);
and UO_242 (O_242,N_24302,N_23603);
nor UO_243 (O_243,N_23770,N_24602);
or UO_244 (O_244,N_22688,N_22784);
and UO_245 (O_245,N_22915,N_24927);
and UO_246 (O_246,N_24162,N_24106);
or UO_247 (O_247,N_23145,N_23996);
or UO_248 (O_248,N_24769,N_23748);
nor UO_249 (O_249,N_23104,N_24307);
or UO_250 (O_250,N_23092,N_23190);
or UO_251 (O_251,N_23178,N_22566);
and UO_252 (O_252,N_23425,N_22659);
nand UO_253 (O_253,N_22617,N_22841);
nor UO_254 (O_254,N_23824,N_23451);
and UO_255 (O_255,N_23325,N_24309);
or UO_256 (O_256,N_23951,N_23795);
nand UO_257 (O_257,N_24951,N_22822);
nor UO_258 (O_258,N_22604,N_24081);
or UO_259 (O_259,N_24225,N_23736);
nand UO_260 (O_260,N_24854,N_23061);
and UO_261 (O_261,N_24398,N_23575);
nand UO_262 (O_262,N_24183,N_24431);
or UO_263 (O_263,N_24117,N_23806);
or UO_264 (O_264,N_24151,N_23386);
nor UO_265 (O_265,N_23271,N_24462);
nor UO_266 (O_266,N_23219,N_24460);
and UO_267 (O_267,N_23805,N_23245);
and UO_268 (O_268,N_23995,N_24148);
and UO_269 (O_269,N_23298,N_23119);
and UO_270 (O_270,N_24814,N_24306);
nor UO_271 (O_271,N_24147,N_24229);
nand UO_272 (O_272,N_24448,N_22917);
or UO_273 (O_273,N_24262,N_23262);
nor UO_274 (O_274,N_23464,N_24645);
or UO_275 (O_275,N_24562,N_24792);
and UO_276 (O_276,N_23275,N_24097);
nand UO_277 (O_277,N_24721,N_23725);
or UO_278 (O_278,N_23872,N_24495);
nor UO_279 (O_279,N_22818,N_24088);
nor UO_280 (O_280,N_22737,N_24227);
or UO_281 (O_281,N_24443,N_24003);
nor UO_282 (O_282,N_22971,N_23566);
nor UO_283 (O_283,N_23743,N_22640);
nand UO_284 (O_284,N_23602,N_23968);
nand UO_285 (O_285,N_22710,N_24777);
or UO_286 (O_286,N_23703,N_23659);
nand UO_287 (O_287,N_23819,N_22641);
and UO_288 (O_288,N_23269,N_24706);
or UO_289 (O_289,N_23784,N_23619);
nand UO_290 (O_290,N_23024,N_24019);
nand UO_291 (O_291,N_23311,N_22868);
or UO_292 (O_292,N_23570,N_22549);
and UO_293 (O_293,N_23623,N_22676);
nor UO_294 (O_294,N_24836,N_23841);
nor UO_295 (O_295,N_23204,N_22749);
and UO_296 (O_296,N_22986,N_22834);
nand UO_297 (O_297,N_23840,N_22909);
xnor UO_298 (O_298,N_24652,N_23042);
nor UO_299 (O_299,N_24904,N_24967);
nor UO_300 (O_300,N_22927,N_24298);
nor UO_301 (O_301,N_23224,N_22999);
nand UO_302 (O_302,N_22994,N_22511);
nor UO_303 (O_303,N_23058,N_24175);
or UO_304 (O_304,N_24549,N_24805);
nor UO_305 (O_305,N_23206,N_23887);
nor UO_306 (O_306,N_22725,N_23755);
nand UO_307 (O_307,N_23699,N_23301);
nand UO_308 (O_308,N_22800,N_24924);
nand UO_309 (O_309,N_23794,N_23480);
or UO_310 (O_310,N_24427,N_23362);
or UO_311 (O_311,N_23277,N_24186);
or UO_312 (O_312,N_22523,N_24547);
or UO_313 (O_313,N_22739,N_24080);
nand UO_314 (O_314,N_24216,N_23698);
and UO_315 (O_315,N_24898,N_23072);
nand UO_316 (O_316,N_24205,N_23565);
and UO_317 (O_317,N_22849,N_22837);
nor UO_318 (O_318,N_23674,N_24568);
and UO_319 (O_319,N_24128,N_22573);
nand UO_320 (O_320,N_23047,N_24929);
or UO_321 (O_321,N_24046,N_23454);
nand UO_322 (O_322,N_23090,N_22905);
or UO_323 (O_323,N_23142,N_24479);
and UO_324 (O_324,N_22979,N_22504);
nor UO_325 (O_325,N_23988,N_24034);
or UO_326 (O_326,N_22792,N_24209);
nor UO_327 (O_327,N_24336,N_23797);
nor UO_328 (O_328,N_23303,N_24103);
nand UO_329 (O_329,N_22738,N_24597);
and UO_330 (O_330,N_24319,N_23859);
and UO_331 (O_331,N_23533,N_22976);
nor UO_332 (O_332,N_23457,N_24082);
or UO_333 (O_333,N_23948,N_23990);
nor UO_334 (O_334,N_24434,N_24373);
nand UO_335 (O_335,N_23727,N_23690);
nor UO_336 (O_336,N_22869,N_23155);
nor UO_337 (O_337,N_22608,N_23926);
and UO_338 (O_338,N_22974,N_22772);
nand UO_339 (O_339,N_24158,N_23902);
nand UO_340 (O_340,N_24680,N_24275);
nor UO_341 (O_341,N_23599,N_22934);
nor UO_342 (O_342,N_22809,N_24376);
nand UO_343 (O_343,N_23769,N_23126);
and UO_344 (O_344,N_22584,N_23829);
and UO_345 (O_345,N_24614,N_23248);
nor UO_346 (O_346,N_24478,N_22893);
nand UO_347 (O_347,N_24998,N_24217);
nand UO_348 (O_348,N_23392,N_24238);
or UO_349 (O_349,N_24452,N_23525);
nor UO_350 (O_350,N_23896,N_22515);
nand UO_351 (O_351,N_23572,N_23992);
and UO_352 (O_352,N_24759,N_23244);
and UO_353 (O_353,N_22899,N_24722);
nand UO_354 (O_354,N_22724,N_22948);
nand UO_355 (O_355,N_24741,N_23804);
and UO_356 (O_356,N_22645,N_23376);
and UO_357 (O_357,N_23663,N_23642);
nand UO_358 (O_358,N_24368,N_23290);
and UO_359 (O_359,N_22706,N_22572);
nand UO_360 (O_360,N_24473,N_24969);
nor UO_361 (O_361,N_23895,N_23400);
and UO_362 (O_362,N_23772,N_23452);
or UO_363 (O_363,N_23856,N_23541);
and UO_364 (O_364,N_22838,N_23188);
nand UO_365 (O_365,N_23515,N_24658);
or UO_366 (O_366,N_24412,N_23511);
nand UO_367 (O_367,N_23274,N_22859);
and UO_368 (O_368,N_22588,N_24595);
or UO_369 (O_369,N_22721,N_23216);
nand UO_370 (O_370,N_22817,N_24846);
and UO_371 (O_371,N_23193,N_24591);
nor UO_372 (O_372,N_24695,N_22852);
and UO_373 (O_373,N_23514,N_24876);
and UO_374 (O_374,N_24573,N_22656);
and UO_375 (O_375,N_23782,N_22614);
and UO_376 (O_376,N_23680,N_22889);
or UO_377 (O_377,N_22746,N_23503);
nor UO_378 (O_378,N_22594,N_23822);
or UO_379 (O_379,N_22672,N_22975);
or UO_380 (O_380,N_24897,N_22703);
nor UO_381 (O_381,N_23422,N_23978);
and UO_382 (O_382,N_24469,N_23931);
nand UO_383 (O_383,N_23594,N_23167);
nand UO_384 (O_384,N_23471,N_24740);
or UO_385 (O_385,N_24592,N_23969);
nor UO_386 (O_386,N_23634,N_23676);
nand UO_387 (O_387,N_24253,N_23681);
and UO_388 (O_388,N_24560,N_24920);
and UO_389 (O_389,N_23751,N_22908);
or UO_390 (O_390,N_24407,N_24043);
nor UO_391 (O_391,N_23682,N_23673);
nor UO_392 (O_392,N_24699,N_22516);
nand UO_393 (O_393,N_23689,N_24065);
nand UO_394 (O_394,N_22980,N_22661);
nor UO_395 (O_395,N_23542,N_23304);
or UO_396 (O_396,N_23767,N_22805);
and UO_397 (O_397,N_23774,N_23552);
nor UO_398 (O_398,N_23173,N_24006);
nand UO_399 (O_399,N_23287,N_23496);
nand UO_400 (O_400,N_24013,N_23508);
nand UO_401 (O_401,N_24036,N_22879);
nand UO_402 (O_402,N_23876,N_23839);
or UO_403 (O_403,N_24608,N_22613);
nand UO_404 (O_404,N_22530,N_23428);
nor UO_405 (O_405,N_23818,N_22621);
nor UO_406 (O_406,N_23777,N_24596);
and UO_407 (O_407,N_23345,N_24167);
or UO_408 (O_408,N_22555,N_23406);
or UO_409 (O_409,N_23848,N_23021);
or UO_410 (O_410,N_24773,N_23463);
nor UO_411 (O_411,N_23122,N_24341);
nor UO_412 (O_412,N_23537,N_24856);
or UO_413 (O_413,N_23625,N_23346);
nor UO_414 (O_414,N_22600,N_23975);
or UO_415 (O_415,N_23007,N_24795);
or UO_416 (O_416,N_22864,N_24131);
nand UO_417 (O_417,N_23149,N_23947);
and UO_418 (O_418,N_22607,N_24489);
and UO_419 (O_419,N_23320,N_23746);
or UO_420 (O_420,N_24796,N_23110);
or UO_421 (O_421,N_24453,N_24886);
nor UO_422 (O_422,N_23453,N_24482);
nand UO_423 (O_423,N_24138,N_24401);
nand UO_424 (O_424,N_23823,N_22929);
nand UO_425 (O_425,N_24014,N_23660);
nor UO_426 (O_426,N_23240,N_24875);
or UO_427 (O_427,N_23112,N_24687);
nor UO_428 (O_428,N_23089,N_24987);
nand UO_429 (O_429,N_23111,N_23984);
nor UO_430 (O_430,N_24701,N_24669);
nand UO_431 (O_431,N_24793,N_23863);
and UO_432 (O_432,N_24402,N_24191);
or UO_433 (O_433,N_24824,N_24696);
or UO_434 (O_434,N_22977,N_23280);
or UO_435 (O_435,N_23225,N_22820);
or UO_436 (O_436,N_23040,N_23027);
and UO_437 (O_437,N_23466,N_22844);
and UO_438 (O_438,N_23079,N_23185);
and UO_439 (O_439,N_23762,N_22666);
or UO_440 (O_440,N_22537,N_23137);
or UO_441 (O_441,N_24691,N_22623);
nand UO_442 (O_442,N_23165,N_24871);
nor UO_443 (O_443,N_24768,N_24571);
nor UO_444 (O_444,N_23852,N_22593);
and UO_445 (O_445,N_23186,N_24564);
and UO_446 (O_446,N_23074,N_24055);
nor UO_447 (O_447,N_23568,N_23812);
and UO_448 (O_448,N_24629,N_23944);
and UO_449 (O_449,N_22642,N_24844);
nor UO_450 (O_450,N_23522,N_23189);
nor UO_451 (O_451,N_23488,N_24962);
nor UO_452 (O_452,N_23234,N_23909);
or UO_453 (O_453,N_23366,N_23624);
and UO_454 (O_454,N_23484,N_24024);
or UO_455 (O_455,N_24772,N_24382);
and UO_456 (O_456,N_22914,N_24095);
or UO_457 (O_457,N_22846,N_24446);
nand UO_458 (O_458,N_24187,N_22660);
nand UO_459 (O_459,N_22557,N_24094);
nor UO_460 (O_460,N_23882,N_24421);
or UO_461 (O_461,N_23781,N_24098);
or UO_462 (O_462,N_23309,N_24734);
nand UO_463 (O_463,N_23322,N_22603);
nor UO_464 (O_464,N_22707,N_22545);
and UO_465 (O_465,N_22997,N_24270);
nand UO_466 (O_466,N_24234,N_24289);
nor UO_467 (O_467,N_24387,N_24454);
or UO_468 (O_468,N_23100,N_22968);
nand UO_469 (O_469,N_23691,N_24177);
and UO_470 (O_470,N_24956,N_24949);
nor UO_471 (O_471,N_22933,N_23214);
nor UO_472 (O_472,N_23831,N_23949);
or UO_473 (O_473,N_23613,N_24126);
nand UO_474 (O_474,N_24931,N_23593);
and UO_475 (O_475,N_23842,N_24141);
or UO_476 (O_476,N_23263,N_22995);
or UO_477 (O_477,N_23272,N_24850);
or UO_478 (O_478,N_22984,N_24603);
or UO_479 (O_479,N_22579,N_23587);
nor UO_480 (O_480,N_24196,N_22518);
and UO_481 (O_481,N_24650,N_24320);
nand UO_482 (O_482,N_22925,N_23826);
and UO_483 (O_483,N_22759,N_24628);
nor UO_484 (O_484,N_24563,N_22575);
nor UO_485 (O_485,N_24727,N_24067);
and UO_486 (O_486,N_22670,N_23737);
and UO_487 (O_487,N_24278,N_22558);
nor UO_488 (O_488,N_24251,N_24149);
or UO_489 (O_489,N_24914,N_23446);
and UO_490 (O_490,N_24411,N_23845);
or UO_491 (O_491,N_24647,N_23260);
xnor UO_492 (O_492,N_24010,N_23242);
nor UO_493 (O_493,N_23472,N_24345);
or UO_494 (O_494,N_22881,N_23348);
nor UO_495 (O_495,N_24798,N_24000);
or UO_496 (O_496,N_22836,N_24089);
nor UO_497 (O_497,N_24505,N_24410);
nor UO_498 (O_498,N_22851,N_24056);
nand UO_499 (O_499,N_24107,N_24957);
and UO_500 (O_500,N_24702,N_23837);
and UO_501 (O_501,N_24352,N_23924);
nand UO_502 (O_502,N_23981,N_23210);
nor UO_503 (O_503,N_24609,N_24829);
nor UO_504 (O_504,N_24780,N_24809);
and UO_505 (O_505,N_24124,N_23971);
and UO_506 (O_506,N_24760,N_22714);
or UO_507 (O_507,N_24002,N_24093);
and UO_508 (O_508,N_22816,N_23067);
nand UO_509 (O_509,N_24005,N_23195);
nor UO_510 (O_510,N_24794,N_24173);
or UO_511 (O_511,N_24422,N_22978);
nand UO_512 (O_512,N_23763,N_23475);
nor UO_513 (O_513,N_24276,N_23732);
nor UO_514 (O_514,N_24900,N_24820);
or UO_515 (O_515,N_23291,N_23055);
nor UO_516 (O_516,N_23907,N_23018);
and UO_517 (O_517,N_23285,N_24976);
nand UO_518 (O_518,N_23633,N_23441);
and UO_519 (O_519,N_23490,N_24709);
nand UO_520 (O_520,N_23636,N_23002);
nand UO_521 (O_521,N_23138,N_23177);
or UO_522 (O_522,N_24841,N_23709);
nor UO_523 (O_523,N_24041,N_24634);
nand UO_524 (O_524,N_23060,N_23294);
nand UO_525 (O_525,N_22677,N_24470);
and UO_526 (O_526,N_23255,N_23005);
and UO_527 (O_527,N_23540,N_24747);
xor UO_528 (O_528,N_24733,N_24330);
or UO_529 (O_529,N_23030,N_24633);
and UO_530 (O_530,N_24861,N_22735);
and UO_531 (O_531,N_23077,N_24828);
nand UO_532 (O_532,N_24582,N_23991);
nor UO_533 (O_533,N_23427,N_24990);
nor UO_534 (O_534,N_23654,N_24812);
nand UO_535 (O_535,N_23563,N_24537);
and UO_536 (O_536,N_23117,N_24979);
nor UO_537 (O_537,N_23296,N_24218);
nand UO_538 (O_538,N_23231,N_22882);
or UO_539 (O_539,N_24159,N_24688);
and UO_540 (O_540,N_22629,N_22653);
nor UO_541 (O_541,N_23960,N_22903);
and UO_542 (O_542,N_22901,N_23897);
nand UO_543 (O_543,N_24388,N_22769);
or UO_544 (O_544,N_23966,N_22990);
or UO_545 (O_545,N_24243,N_23922);
nand UO_546 (O_546,N_24580,N_24530);
or UO_547 (O_547,N_22907,N_24715);
nor UO_548 (O_548,N_24807,N_24630);
or UO_549 (O_549,N_23015,N_23326);
and UO_550 (O_550,N_24857,N_23757);
nor UO_551 (O_551,N_23605,N_22952);
nand UO_552 (O_552,N_24649,N_23598);
nor UO_553 (O_553,N_24804,N_24996);
nor UO_554 (O_554,N_22988,N_23344);
or UO_555 (O_555,N_22953,N_23588);
nand UO_556 (O_556,N_22626,N_23157);
or UO_557 (O_557,N_24508,N_24619);
or UO_558 (O_558,N_22531,N_23535);
nand UO_559 (O_559,N_23373,N_22643);
nand UO_560 (O_560,N_24344,N_24703);
nand UO_561 (O_561,N_22682,N_24848);
or UO_562 (O_562,N_23808,N_24791);
nor UO_563 (O_563,N_24120,N_23728);
and UO_564 (O_564,N_23378,N_22789);
or UO_565 (O_565,N_22540,N_24843);
or UO_566 (O_566,N_24864,N_24308);
and UO_567 (O_567,N_23282,N_24129);
nor UO_568 (O_568,N_24265,N_23678);
nand UO_569 (O_569,N_23722,N_24783);
or UO_570 (O_570,N_22539,N_24380);
or UO_571 (O_571,N_22942,N_23959);
and UO_572 (O_572,N_24683,N_22742);
and UO_573 (O_573,N_23456,N_23032);
nand UO_574 (O_574,N_23053,N_23807);
nor UO_575 (O_575,N_22931,N_22571);
nand UO_576 (O_576,N_24555,N_23756);
and UO_577 (O_577,N_23132,N_24941);
or UO_578 (O_578,N_24860,N_24203);
or UO_579 (O_579,N_24685,N_24377);
nor UO_580 (O_580,N_23445,N_23233);
and UO_581 (O_581,N_24821,N_23569);
and UO_582 (O_582,N_22861,N_24310);
nor UO_583 (O_583,N_22715,N_22528);
nor UO_584 (O_584,N_23892,N_22701);
and UO_585 (O_585,N_22618,N_24285);
or UO_586 (O_586,N_23986,N_23374);
or UO_587 (O_587,N_24775,N_24598);
or UO_588 (O_588,N_23412,N_24586);
nand UO_589 (O_589,N_24954,N_24403);
nand UO_590 (O_590,N_24574,N_24788);
nand UO_591 (O_591,N_23520,N_24559);
and UO_592 (O_592,N_23476,N_22947);
and UO_593 (O_593,N_24880,N_23814);
and UO_594 (O_594,N_24764,N_22919);
and UO_595 (O_595,N_24263,N_24512);
nor UO_596 (O_596,N_24926,N_23820);
nor UO_597 (O_597,N_23967,N_23093);
nor UO_598 (O_598,N_24936,N_24280);
or UO_599 (O_599,N_22833,N_23340);
nor UO_600 (O_600,N_23900,N_24578);
or UO_601 (O_601,N_24961,N_24789);
and UO_602 (O_602,N_23364,N_23798);
nand UO_603 (O_603,N_23611,N_23631);
and UO_604 (O_604,N_24390,N_24488);
or UO_605 (O_605,N_24474,N_22687);
nand UO_606 (O_606,N_22787,N_24127);
or UO_607 (O_607,N_22883,N_23404);
nor UO_608 (O_608,N_24363,N_24315);
nor UO_609 (O_609,N_24917,N_23113);
nand UO_610 (O_610,N_23147,N_24992);
nor UO_611 (O_611,N_24500,N_22855);
and UO_612 (O_612,N_24413,N_23538);
and UO_613 (O_613,N_22795,N_24327);
or UO_614 (O_614,N_23127,N_23864);
or UO_615 (O_615,N_23942,N_23648);
nand UO_616 (O_616,N_24616,N_22774);
and UO_617 (O_617,N_22704,N_23857);
or UO_618 (O_618,N_23750,N_24269);
nor UO_619 (O_619,N_23369,N_23038);
or UO_620 (O_620,N_24561,N_23861);
nor UO_621 (O_621,N_24660,N_24553);
nand UO_622 (O_622,N_24831,N_23954);
or UO_623 (O_623,N_24575,N_23898);
nor UO_624 (O_624,N_22763,N_22806);
nor UO_625 (O_625,N_24397,N_24928);
nand UO_626 (O_626,N_24012,N_24185);
nand UO_627 (O_627,N_22989,N_24208);
nor UO_628 (O_628,N_23141,N_24323);
nand UO_629 (O_629,N_23687,N_24932);
or UO_630 (O_630,N_24862,N_23091);
nor UO_631 (O_631,N_24299,N_23385);
nand UO_632 (O_632,N_22683,N_24045);
or UO_633 (O_633,N_23355,N_24551);
nor UO_634 (O_634,N_24973,N_23154);
nor UO_635 (O_635,N_24358,N_23319);
and UO_636 (O_636,N_23099,N_22951);
or UO_637 (O_637,N_24483,N_24697);
and UO_638 (O_638,N_22972,N_24778);
and UO_639 (O_639,N_22595,N_22731);
nand UO_640 (O_640,N_23076,N_23801);
or UO_641 (O_641,N_22508,N_24692);
nand UO_642 (O_642,N_23923,N_24057);
or UO_643 (O_643,N_24134,N_23318);
nand UO_644 (O_644,N_23817,N_24161);
and UO_645 (O_645,N_23640,N_24601);
or UO_646 (O_646,N_24899,N_23012);
nand UO_647 (O_647,N_24326,N_23509);
nand UO_648 (O_648,N_24109,N_22567);
or UO_649 (O_649,N_24021,N_22541);
and UO_650 (O_650,N_24414,N_24077);
nand UO_651 (O_651,N_23544,N_22559);
or UO_652 (O_652,N_23270,N_24653);
or UO_653 (O_653,N_24916,N_23891);
nor UO_654 (O_654,N_22906,N_23785);
or UO_655 (O_655,N_23347,N_24882);
and UO_656 (O_656,N_24690,N_24370);
nor UO_657 (O_657,N_24184,N_23396);
nand UO_658 (O_658,N_24391,N_23419);
and UO_659 (O_659,N_24237,N_23046);
nor UO_660 (O_660,N_24673,N_22944);
or UO_661 (O_661,N_24394,N_24666);
or UO_662 (O_662,N_24714,N_22709);
and UO_663 (O_663,N_23610,N_23229);
nand UO_664 (O_664,N_22563,N_23435);
nand UO_665 (O_665,N_23649,N_24766);
and UO_666 (O_666,N_24737,N_22685);
and UO_667 (O_667,N_23353,N_23843);
and UO_668 (O_668,N_23661,N_22561);
or UO_669 (O_669,N_24018,N_24360);
and UO_670 (O_670,N_24762,N_23656);
or UO_671 (O_671,N_24392,N_24842);
nand UO_672 (O_672,N_22730,N_22577);
nand UO_673 (O_673,N_24940,N_23026);
nand UO_674 (O_674,N_24569,N_23213);
nor UO_675 (O_675,N_22862,N_24318);
nand UO_676 (O_676,N_23331,N_23761);
nor UO_677 (O_677,N_24501,N_24070);
or UO_678 (O_678,N_23360,N_23780);
and UO_679 (O_679,N_23034,N_23152);
or UO_680 (O_680,N_24746,N_24677);
or UO_681 (O_681,N_23792,N_24863);
nor UO_682 (O_682,N_24266,N_24220);
nor UO_683 (O_683,N_24545,N_22912);
and UO_684 (O_684,N_24739,N_23972);
and UO_685 (O_685,N_23813,N_24132);
or UO_686 (O_686,N_22649,N_24027);
nor UO_687 (O_687,N_22520,N_22568);
or UO_688 (O_688,N_24423,N_23879);
and UO_689 (O_689,N_24249,N_23000);
or UO_690 (O_690,N_24053,N_22954);
and UO_691 (O_691,N_24178,N_24393);
nor UO_692 (O_692,N_23510,N_22619);
nor UO_693 (O_693,N_24767,N_23497);
or UO_694 (O_694,N_23044,N_22580);
and UO_695 (O_695,N_23439,N_24211);
or UO_696 (O_696,N_23197,N_23918);
nor UO_697 (O_697,N_23409,N_23159);
nand UO_698 (O_698,N_23228,N_23715);
or UO_699 (O_699,N_24901,N_22723);
nor UO_700 (O_700,N_24137,N_24605);
nor UO_701 (O_701,N_23930,N_24441);
nand UO_702 (O_702,N_24455,N_23953);
or UO_703 (O_703,N_23833,N_24415);
nor UO_704 (O_704,N_23937,N_23665);
and UO_705 (O_705,N_23939,N_24700);
or UO_706 (O_706,N_22797,N_24771);
or UO_707 (O_707,N_22596,N_23434);
and UO_708 (O_708,N_22863,N_24781);
or UO_709 (O_709,N_22770,N_23714);
and UO_710 (O_710,N_23903,N_23095);
or UO_711 (O_711,N_23337,N_22923);
or UO_712 (O_712,N_23066,N_22716);
and UO_713 (O_713,N_23685,N_23003);
and UO_714 (O_714,N_24016,N_24406);
nand UO_715 (O_715,N_23500,N_23171);
nand UO_716 (O_716,N_24051,N_24222);
and UO_717 (O_717,N_23580,N_22503);
nand UO_718 (O_718,N_24044,N_22981);
nor UO_719 (O_719,N_24166,N_22514);
nand UO_720 (O_720,N_24419,N_24520);
or UO_721 (O_721,N_23420,N_24623);
nand UO_722 (O_722,N_23230,N_22991);
nor UO_723 (O_723,N_23788,N_24763);
and UO_724 (O_724,N_23050,N_23928);
nor UO_725 (O_725,N_23470,N_22536);
and UO_726 (O_726,N_23261,N_24548);
nand UO_727 (O_727,N_23252,N_23744);
nand UO_728 (O_728,N_23880,N_23606);
nor UO_729 (O_729,N_22967,N_23001);
and UO_730 (O_730,N_23128,N_24934);
or UO_731 (O_731,N_23408,N_24142);
nor UO_732 (O_732,N_24833,N_23519);
or UO_733 (O_733,N_24984,N_23388);
nor UO_734 (O_734,N_23107,N_22585);
or UO_735 (O_735,N_23164,N_23629);
nor UO_736 (O_736,N_22612,N_24400);
or UO_737 (O_737,N_24632,N_22830);
and UO_738 (O_738,N_23448,N_24579);
and UO_739 (O_739,N_23144,N_24585);
nor UO_740 (O_740,N_22631,N_22713);
nand UO_741 (O_741,N_23267,N_23354);
and UO_742 (O_742,N_23652,N_24213);
nor UO_743 (O_743,N_23410,N_23051);
nand UO_744 (O_744,N_24365,N_23375);
nor UO_745 (O_745,N_24287,N_22884);
and UO_746 (O_746,N_24242,N_23431);
and UO_747 (O_747,N_23965,N_24896);
or UO_748 (O_748,N_22521,N_23908);
or UO_749 (O_749,N_24086,N_23747);
nor UO_750 (O_750,N_22576,N_23115);
and UO_751 (O_751,N_22761,N_24670);
or UO_752 (O_752,N_23802,N_23056);
or UO_753 (O_753,N_22693,N_24826);
and UO_754 (O_754,N_23583,N_22888);
and UO_755 (O_755,N_24525,N_23925);
nand UO_756 (O_756,N_24797,N_23220);
nor UO_757 (O_757,N_22740,N_23334);
nor UO_758 (O_758,N_23249,N_24599);
and UO_759 (O_759,N_24654,N_23597);
and UO_760 (O_760,N_23169,N_24785);
nand UO_761 (O_761,N_23049,N_24790);
and UO_762 (O_762,N_23288,N_23421);
nand UO_763 (O_763,N_24366,N_23974);
nor UO_764 (O_764,N_24292,N_23998);
and UO_765 (O_765,N_23424,N_23667);
nor UO_766 (O_766,N_24338,N_23462);
nand UO_767 (O_767,N_23310,N_24084);
or UO_768 (O_768,N_24745,N_23194);
nor UO_769 (O_769,N_23564,N_24515);
nand UO_770 (O_770,N_23628,N_23639);
and UO_771 (O_771,N_24075,N_23671);
and UO_772 (O_772,N_24684,N_22959);
and UO_773 (O_773,N_23911,N_22814);
or UO_774 (O_774,N_23283,N_24321);
nor UO_775 (O_775,N_23517,N_22733);
nand UO_776 (O_776,N_24541,N_23478);
or UO_777 (O_777,N_24395,N_23993);
or UO_778 (O_778,N_24439,N_22767);
nor UO_779 (O_779,N_22729,N_23414);
or UO_780 (O_780,N_24118,N_23098);
or UO_781 (O_781,N_24257,N_24374);
nand UO_782 (O_782,N_23243,N_22924);
nor UO_783 (O_783,N_22945,N_24923);
or UO_784 (O_784,N_24248,N_23940);
and UO_785 (O_785,N_23361,N_22665);
and UO_786 (O_786,N_23612,N_24892);
nor UO_787 (O_787,N_24228,N_22802);
nor UO_788 (O_788,N_24966,N_23182);
and UO_789 (O_789,N_22877,N_23114);
or UO_790 (O_790,N_22694,N_23871);
or UO_791 (O_791,N_23417,N_23550);
nand UO_792 (O_792,N_23913,N_24197);
nor UO_793 (O_793,N_23172,N_24496);
or UO_794 (O_794,N_24176,N_23150);
nand UO_795 (O_795,N_23437,N_24935);
nor UO_796 (O_796,N_23212,N_24194);
and UO_797 (O_797,N_24182,N_23683);
nor UO_798 (O_798,N_23069,N_24584);
and UO_799 (O_799,N_22611,N_22965);
nand UO_800 (O_800,N_24847,N_22973);
nand UO_801 (O_801,N_23604,N_23759);
or UO_802 (O_802,N_24459,N_24637);
nand UO_803 (O_803,N_23306,N_23945);
and UO_804 (O_804,N_24988,N_23582);
or UO_805 (O_805,N_24372,N_24333);
nand UO_806 (O_806,N_24353,N_23869);
nor UO_807 (O_807,N_22866,N_23179);
nor UO_808 (O_808,N_23429,N_24878);
nand UO_809 (O_809,N_22936,N_24890);
or UO_810 (O_810,N_24201,N_22548);
nand UO_811 (O_811,N_24100,N_23622);
and UO_812 (O_812,N_24384,N_23516);
or UO_813 (O_813,N_24802,N_22609);
nand UO_814 (O_814,N_24030,N_22858);
nand UO_815 (O_815,N_24980,N_23983);
or UO_816 (O_816,N_22582,N_24726);
and UO_817 (O_817,N_22639,N_23483);
or UO_818 (O_818,N_24866,N_22638);
nand UO_819 (O_819,N_23140,N_23101);
nor UO_820 (O_820,N_23467,N_22790);
xor UO_821 (O_821,N_23036,N_24799);
and UO_822 (O_822,N_24533,N_23211);
nor UO_823 (O_823,N_23258,N_23191);
nand UO_824 (O_824,N_23586,N_24233);
or UO_825 (O_825,N_24212,N_22897);
and UO_826 (O_826,N_23153,N_24676);
nor UO_827 (O_827,N_23335,N_23062);
and UO_828 (O_828,N_23810,N_24963);
and UO_829 (O_829,N_24324,N_22708);
nand UO_830 (O_830,N_22819,N_23834);
nor UO_831 (O_831,N_24832,N_23359);
or UO_832 (O_832,N_23692,N_23706);
and UO_833 (O_833,N_23679,N_23492);
and UO_834 (O_834,N_23601,N_23118);
or UO_835 (O_835,N_23838,N_22780);
nor UO_836 (O_836,N_24523,N_24235);
nand UO_837 (O_837,N_24823,N_24522);
nand UO_838 (O_838,N_24995,N_24499);
nor UO_839 (O_839,N_24516,N_24589);
or UO_840 (O_840,N_23741,N_24787);
nor UO_841 (O_841,N_24540,N_24983);
nor UO_842 (O_842,N_23608,N_24020);
nand UO_843 (O_843,N_23082,N_22599);
or UO_844 (O_844,N_24435,N_24083);
nor UO_845 (O_845,N_23052,N_22684);
nand UO_846 (O_846,N_24710,N_23175);
nor UO_847 (O_847,N_22627,N_24156);
or UO_848 (O_848,N_23668,N_23554);
and UO_849 (O_849,N_24071,N_24417);
or UO_850 (O_850,N_23657,N_24146);
nor UO_851 (O_851,N_24029,N_24751);
nor UO_852 (O_852,N_24813,N_24416);
or UO_853 (O_853,N_24364,N_24017);
nor UO_854 (O_854,N_23324,N_24905);
nor UO_855 (O_855,N_23200,N_24808);
or UO_856 (O_856,N_24301,N_23235);
nor UO_857 (O_857,N_24909,N_22885);
nor UO_858 (O_858,N_23776,N_23208);
nand UO_859 (O_859,N_24074,N_24748);
and UO_860 (O_860,N_24060,N_23830);
nand UO_861 (O_861,N_22636,N_23299);
or UO_862 (O_862,N_23307,N_23278);
nor UO_863 (O_863,N_23162,N_22831);
nor UO_864 (O_864,N_23135,N_24648);
and UO_865 (O_865,N_24337,N_24919);
nand UO_866 (O_866,N_24311,N_23402);
or UO_867 (O_867,N_24180,N_24830);
nand UO_868 (O_868,N_23081,N_24576);
or UO_869 (O_869,N_24873,N_24252);
nand UO_870 (O_870,N_24037,N_23506);
and UO_871 (O_871,N_24059,N_24312);
and UO_872 (O_872,N_24404,N_24554);
and UO_873 (O_873,N_23273,N_23854);
or UO_874 (O_874,N_22726,N_23073);
or UO_875 (O_875,N_23367,N_24042);
nor UO_876 (O_876,N_23017,N_23742);
nor UO_877 (O_877,N_23712,N_22534);
nor UO_878 (O_878,N_24078,N_22875);
or UO_879 (O_879,N_24879,N_24305);
or UO_880 (O_880,N_23827,N_24268);
nor UO_881 (O_881,N_22996,N_24707);
nand UO_882 (O_882,N_23529,N_23915);
or UO_883 (O_883,N_23693,N_23444);
and UO_884 (O_884,N_22801,N_23336);
xnor UO_885 (O_885,N_23227,N_23920);
nand UO_886 (O_886,N_23710,N_23237);
nand UO_887 (O_887,N_23389,N_22547);
or UO_888 (O_888,N_23096,N_22513);
xnor UO_889 (O_889,N_23846,N_23724);
or UO_890 (O_890,N_23350,N_24999);
nand UO_891 (O_891,N_22741,N_24432);
and UO_892 (O_892,N_23677,N_23976);
and UO_893 (O_893,N_23702,N_23655);
nor UO_894 (O_894,N_24486,N_22668);
nor UO_895 (O_895,N_24544,N_24466);
and UO_896 (O_896,N_24145,N_24534);
nand UO_897 (O_897,N_24557,N_24288);
and UO_898 (O_898,N_23013,N_24456);
or UO_899 (O_899,N_24206,N_24693);
and UO_900 (O_900,N_23927,N_24997);
or UO_901 (O_901,N_23254,N_24004);
nor UO_902 (O_902,N_22755,N_22583);
nor UO_903 (O_903,N_24121,N_23315);
nand UO_904 (O_904,N_23377,N_22757);
and UO_905 (O_905,N_23513,N_23753);
or UO_906 (O_906,N_22964,N_23729);
nor UO_907 (O_907,N_22813,N_23370);
nand UO_908 (O_908,N_24918,N_23016);
xnor UO_909 (O_909,N_23305,N_23080);
or UO_910 (O_910,N_23870,N_24912);
and UO_911 (O_911,N_24335,N_23474);
or UO_912 (O_912,N_22867,N_24468);
nand UO_913 (O_913,N_24853,N_24993);
nor UO_914 (O_914,N_23238,N_23084);
nor UO_915 (O_915,N_23064,N_23962);
or UO_916 (O_916,N_22598,N_22681);
nor UO_917 (O_917,N_23874,N_24718);
and UO_918 (O_918,N_24837,N_24294);
nor UO_919 (O_919,N_23094,N_24079);
nor UO_920 (O_920,N_24930,N_24140);
and UO_921 (O_921,N_23549,N_23391);
or UO_922 (O_922,N_22969,N_24765);
and UO_923 (O_923,N_22606,N_23120);
and UO_924 (O_924,N_24743,N_22646);
nand UO_925 (O_925,N_22910,N_24955);
nor UO_926 (O_926,N_23707,N_22848);
or UO_927 (O_927,N_23403,N_23257);
and UO_928 (O_928,N_24471,N_23265);
nor UO_929 (O_929,N_22562,N_24214);
nor UO_930 (O_930,N_24153,N_24895);
and UO_931 (O_931,N_22960,N_24389);
and UO_932 (O_932,N_24570,N_23368);
nand UO_933 (O_933,N_23791,N_24581);
and UO_934 (O_934,N_23180,N_23617);
nand UO_935 (O_935,N_23130,N_24475);
nor UO_936 (O_936,N_24224,N_23607);
and UO_937 (O_937,N_24322,N_23579);
nor UO_938 (O_938,N_23393,N_24908);
nor UO_939 (O_939,N_23498,N_23646);
and UO_940 (O_940,N_23524,N_23917);
nor UO_941 (O_941,N_23592,N_23136);
nor UO_942 (O_942,N_23853,N_23650);
or UO_943 (O_943,N_24521,N_24937);
nor UO_944 (O_944,N_23950,N_24834);
and UO_945 (O_945,N_22799,N_23620);
and UO_946 (O_946,N_22890,N_22958);
or UO_947 (O_947,N_24849,N_23103);
nor UO_948 (O_948,N_23638,N_22552);
and UO_949 (O_949,N_24202,N_22840);
nor UO_950 (O_950,N_23489,N_24102);
nor UO_951 (O_951,N_23020,N_24877);
nand UO_952 (O_952,N_23730,N_22916);
nand UO_953 (O_953,N_23719,N_23860);
or UO_954 (O_954,N_24241,N_22722);
and UO_955 (O_955,N_22832,N_22752);
nand UO_956 (O_956,N_22615,N_24160);
and UO_957 (O_957,N_23618,N_24090);
nand UO_958 (O_958,N_23910,N_23536);
nor UO_959 (O_959,N_23486,N_23250);
nand UO_960 (O_960,N_23070,N_23669);
nor UO_961 (O_961,N_24942,N_23383);
nand UO_962 (O_962,N_24284,N_24035);
nand UO_963 (O_963,N_23653,N_24113);
nand UO_964 (O_964,N_24332,N_24524);
or UO_965 (O_965,N_22768,N_23443);
nor UO_966 (O_966,N_24112,N_22828);
or UO_967 (O_967,N_24215,N_24314);
nor UO_968 (O_968,N_22824,N_24662);
nand UO_969 (O_969,N_23339,N_24150);
or UO_970 (O_970,N_22962,N_24199);
or UO_971 (O_971,N_24933,N_23028);
nor UO_972 (O_972,N_24583,N_22961);
and UO_973 (O_973,N_23528,N_24907);
nor UO_974 (O_974,N_24756,N_22766);
nor UO_975 (O_975,N_23718,N_23556);
nor UO_976 (O_976,N_24668,N_24776);
nor UO_977 (O_977,N_24436,N_24283);
or UO_978 (O_978,N_24169,N_23143);
and UO_979 (O_979,N_24543,N_22856);
nor UO_980 (O_980,N_22554,N_22696);
nand UO_981 (O_981,N_23695,N_23553);
and UO_982 (O_982,N_23979,N_24750);
nand UO_983 (O_983,N_23630,N_22551);
nand UO_984 (O_984,N_22998,N_24255);
or UO_985 (O_985,N_23716,N_24157);
and UO_986 (O_986,N_23557,N_22850);
or UO_987 (O_987,N_23071,N_23615);
nand UO_988 (O_988,N_24960,N_23789);
and UO_989 (O_989,N_22762,N_24816);
and UO_990 (O_990,N_23901,N_23771);
or UO_991 (O_991,N_22845,N_23201);
nand UO_992 (O_992,N_24627,N_23873);
or UO_993 (O_993,N_24558,N_22651);
or UO_994 (O_994,N_24556,N_22904);
and UO_995 (O_995,N_23259,N_24334);
nor UO_996 (O_996,N_23176,N_23399);
or UO_997 (O_997,N_24742,N_24424);
nand UO_998 (O_998,N_22871,N_23851);
nand UO_999 (O_999,N_23987,N_24339);
or UO_1000 (O_1000,N_22692,N_24163);
nor UO_1001 (O_1001,N_24550,N_22946);
or UO_1002 (O_1002,N_22829,N_22592);
or UO_1003 (O_1003,N_23323,N_23670);
and UO_1004 (O_1004,N_22705,N_23957);
nor UO_1005 (O_1005,N_22853,N_22745);
nor UO_1006 (O_1006,N_24947,N_22602);
or UO_1007 (O_1007,N_23332,N_24989);
or UO_1008 (O_1008,N_24172,N_23662);
nand UO_1009 (O_1009,N_22898,N_24193);
and UO_1010 (O_1010,N_24945,N_22807);
or UO_1011 (O_1011,N_24818,N_23407);
nand UO_1012 (O_1012,N_22993,N_24092);
nor UO_1013 (O_1013,N_23723,N_22956);
and UO_1014 (O_1014,N_24343,N_24481);
or UO_1015 (O_1015,N_24567,N_22785);
nor UO_1016 (O_1016,N_24007,N_22544);
and UO_1017 (O_1017,N_23551,N_23264);
and UO_1018 (O_1018,N_22810,N_23672);
nor UO_1019 (O_1019,N_23041,N_22680);
nand UO_1020 (O_1020,N_23836,N_23884);
or UO_1021 (O_1021,N_24445,N_23382);
and UO_1022 (O_1022,N_24572,N_24405);
or UO_1023 (O_1023,N_22793,N_24378);
and UO_1024 (O_1024,N_23867,N_22786);
or UO_1025 (O_1025,N_24958,N_23581);
and UO_1026 (O_1026,N_24232,N_24350);
nand UO_1027 (O_1027,N_23704,N_24640);
nand UO_1028 (O_1028,N_22928,N_22870);
nand UO_1029 (O_1029,N_23014,N_23577);
or UO_1030 (O_1030,N_24610,N_24717);
nor UO_1031 (O_1031,N_23160,N_22825);
nand UO_1032 (O_1032,N_23720,N_23547);
nand UO_1033 (O_1033,N_23163,N_23207);
or UO_1034 (O_1034,N_24870,N_22533);
or UO_1035 (O_1035,N_24638,N_22675);
nor UO_1036 (O_1036,N_24888,N_22985);
nand UO_1037 (O_1037,N_23576,N_24171);
or UO_1038 (O_1038,N_24724,N_23881);
or UO_1039 (O_1039,N_24357,N_24752);
or UO_1040 (O_1040,N_24297,N_23078);
nand UO_1041 (O_1041,N_23203,N_24840);
or UO_1042 (O_1042,N_22955,N_23905);
nor UO_1043 (O_1043,N_22791,N_23973);
and UO_1044 (O_1044,N_24174,N_24231);
nand UO_1045 (O_1045,N_23202,N_24744);
nor UO_1046 (O_1046,N_24379,N_22506);
nor UO_1047 (O_1047,N_23858,N_24438);
nand UO_1048 (O_1048,N_23450,N_24296);
and UO_1049 (O_1049,N_24429,N_24155);
nor UO_1050 (O_1050,N_24518,N_23961);
or UO_1051 (O_1051,N_24492,N_23491);
nor UO_1052 (O_1052,N_24328,N_22691);
nand UO_1053 (O_1053,N_23561,N_22798);
nand UO_1054 (O_1054,N_24851,N_23946);
and UO_1055 (O_1055,N_24011,N_24444);
nand UO_1056 (O_1056,N_24922,N_24279);
and UO_1057 (O_1057,N_22605,N_23534);
nand UO_1058 (O_1058,N_24566,N_24872);
nand UO_1059 (O_1059,N_22587,N_23411);
or UO_1060 (O_1060,N_24663,N_24825);
nor UO_1061 (O_1061,N_22921,N_22827);
nand UO_1062 (O_1062,N_22748,N_24272);
nand UO_1063 (O_1063,N_24672,N_23701);
and UO_1064 (O_1064,N_24970,N_23398);
and UO_1065 (O_1065,N_23560,N_24073);
nand UO_1066 (O_1066,N_23241,N_22758);
nand UO_1067 (O_1067,N_22992,N_22652);
and UO_1068 (O_1068,N_23481,N_23327);
and UO_1069 (O_1069,N_22648,N_24643);
nor UO_1070 (O_1070,N_24062,N_23268);
and UO_1071 (O_1071,N_23358,N_24770);
or UO_1072 (O_1072,N_23849,N_24729);
or UO_1073 (O_1073,N_23308,N_23585);
xnor UO_1074 (O_1074,N_23811,N_24535);
nor UO_1075 (O_1075,N_24498,N_24165);
and UO_1076 (O_1076,N_24340,N_24048);
nor UO_1077 (O_1077,N_24313,N_24517);
and UO_1078 (O_1078,N_23531,N_22564);
and UO_1079 (O_1079,N_23752,N_22522);
nand UO_1080 (O_1080,N_24835,N_23395);
and UO_1081 (O_1081,N_22634,N_23416);
nand UO_1082 (O_1082,N_22550,N_24600);
or UO_1083 (O_1083,N_23302,N_22808);
nand UO_1084 (O_1084,N_22625,N_23532);
nand UO_1085 (O_1085,N_24604,N_23033);
nand UO_1086 (O_1086,N_24682,N_22586);
nand UO_1087 (O_1087,N_23253,N_23236);
or UO_1088 (O_1088,N_23825,N_22860);
nand UO_1089 (O_1089,N_23029,N_24894);
nor UO_1090 (O_1090,N_24801,N_24593);
or UO_1091 (O_1091,N_24952,N_23151);
nor UO_1092 (O_1092,N_24052,N_23121);
nand UO_1093 (O_1093,N_23548,N_24891);
nor UO_1094 (O_1094,N_23994,N_23832);
or UO_1095 (O_1095,N_23105,N_22695);
or UO_1096 (O_1096,N_23333,N_22932);
nor UO_1097 (O_1097,N_24925,N_24300);
nor UO_1098 (O_1098,N_22674,N_23883);
or UO_1099 (O_1099,N_24713,N_22880);
nand UO_1100 (O_1100,N_24348,N_23365);
and UO_1101 (O_1101,N_22597,N_24939);
and UO_1102 (O_1102,N_24527,N_23855);
and UO_1103 (O_1103,N_22811,N_24758);
and UO_1104 (O_1104,N_24502,N_24800);
nand UO_1105 (O_1105,N_24867,N_23485);
or UO_1106 (O_1106,N_23479,N_24040);
and UO_1107 (O_1107,N_24239,N_23696);
or UO_1108 (O_1108,N_23381,N_24490);
nand UO_1109 (O_1109,N_24631,N_24782);
nor UO_1110 (O_1110,N_23170,N_23862);
nand UO_1111 (O_1111,N_22751,N_24108);
nand UO_1112 (O_1112,N_24738,N_23289);
or UO_1113 (O_1113,N_24480,N_24144);
and UO_1114 (O_1114,N_24245,N_23760);
nor UO_1115 (O_1115,N_22744,N_24303);
and UO_1116 (O_1116,N_24087,N_22535);
or UO_1117 (O_1117,N_23765,N_22655);
and UO_1118 (O_1118,N_22678,N_22601);
nand UO_1119 (O_1119,N_22775,N_24271);
nor UO_1120 (O_1120,N_22507,N_24418);
or UO_1121 (O_1121,N_24244,N_23426);
nand UO_1122 (O_1122,N_22700,N_24033);
and UO_1123 (O_1123,N_23936,N_23232);
and UO_1124 (O_1124,N_22500,N_23276);
nor UO_1125 (O_1125,N_23766,N_24913);
nor UO_1126 (O_1126,N_23086,N_24050);
or UO_1127 (O_1127,N_24179,N_23735);
and UO_1128 (O_1128,N_24681,N_23758);
or UO_1129 (O_1129,N_24674,N_24259);
nand UO_1130 (O_1130,N_24735,N_24286);
or UO_1131 (O_1131,N_23571,N_23139);
and UO_1132 (O_1132,N_24061,N_22900);
nor UO_1133 (O_1133,N_23803,N_24615);
or UO_1134 (O_1134,N_24440,N_22663);
nor UO_1135 (O_1135,N_24859,N_24130);
nor UO_1136 (O_1136,N_23621,N_24420);
or UO_1137 (O_1137,N_23239,N_23338);
and UO_1138 (O_1138,N_24304,N_24611);
or UO_1139 (O_1139,N_23938,N_24484);
and UO_1140 (O_1140,N_22796,N_23019);
and UO_1141 (O_1141,N_23401,N_24347);
nor UO_1142 (O_1142,N_22556,N_23379);
nor UO_1143 (O_1143,N_23773,N_24119);
and UO_1144 (O_1144,N_23352,N_24316);
and UO_1145 (O_1145,N_24736,N_23686);
nor UO_1146 (O_1146,N_24437,N_24110);
or UO_1147 (O_1147,N_24198,N_24811);
and UO_1148 (O_1148,N_23738,N_23573);
and UO_1149 (O_1149,N_22843,N_23501);
nor UO_1150 (O_1150,N_24716,N_23596);
and UO_1151 (O_1151,N_23461,N_24978);
or UO_1152 (O_1152,N_22673,N_23850);
and UO_1153 (O_1153,N_22943,N_23929);
nor UO_1154 (O_1154,N_24291,N_23889);
nand UO_1155 (O_1155,N_23899,N_24915);
nand UO_1156 (O_1156,N_24408,N_23878);
and UO_1157 (O_1157,N_22509,N_22644);
and UO_1158 (O_1158,N_23133,N_22941);
and UO_1159 (O_1159,N_23131,N_24223);
and UO_1160 (O_1160,N_23357,N_23011);
or UO_1161 (O_1161,N_24457,N_22553);
and UO_1162 (O_1162,N_24274,N_23218);
nand UO_1163 (O_1163,N_23512,N_23313);
nand UO_1164 (O_1164,N_23048,N_22570);
and UO_1165 (O_1165,N_24143,N_24396);
and UO_1166 (O_1166,N_23739,N_24911);
and UO_1167 (O_1167,N_23626,N_22628);
or UO_1168 (O_1168,N_24635,N_23675);
nor UO_1169 (O_1169,N_23209,N_23504);
nand UO_1170 (O_1170,N_24694,N_24116);
nor UO_1171 (O_1171,N_24122,N_24686);
nor UO_1172 (O_1172,N_22949,N_23635);
nor UO_1173 (O_1173,N_23964,N_22782);
and UO_1174 (O_1174,N_22650,N_23088);
or UO_1175 (O_1175,N_22510,N_23181);
or UO_1176 (O_1176,N_24254,N_22728);
nand UO_1177 (O_1177,N_24531,N_23387);
or UO_1178 (O_1178,N_22743,N_23886);
nor UO_1179 (O_1179,N_24200,N_23031);
and UO_1180 (O_1180,N_24506,N_22667);
or UO_1181 (O_1181,N_23418,N_23799);
and UO_1182 (O_1182,N_24712,N_24971);
or UO_1183 (O_1183,N_24839,N_23108);
nand UO_1184 (O_1184,N_24858,N_24732);
nor UO_1185 (O_1185,N_24675,N_24031);
or UO_1186 (O_1186,N_23934,N_22982);
nor UO_1187 (O_1187,N_22501,N_22532);
nand UO_1188 (O_1188,N_24491,N_23183);
and UO_1189 (O_1189,N_23156,N_24868);
and UO_1190 (O_1190,N_22778,N_23458);
and UO_1191 (O_1191,N_24038,N_24612);
or UO_1192 (O_1192,N_23877,N_24869);
or UO_1193 (O_1193,N_24001,N_24139);
or UO_1194 (O_1194,N_24964,N_24855);
nor UO_1195 (O_1195,N_23651,N_23999);
and UO_1196 (O_1196,N_22872,N_24528);
and UO_1197 (O_1197,N_22697,N_24679);
or UO_1198 (O_1198,N_23394,N_24069);
or UO_1199 (O_1199,N_24657,N_24950);
and UO_1200 (O_1200,N_23935,N_23955);
and UO_1201 (O_1201,N_22519,N_22765);
nor UO_1202 (O_1202,N_23184,N_23559);
nor UO_1203 (O_1203,N_23790,N_22578);
nor UO_1204 (O_1204,N_24195,N_24226);
nor UO_1205 (O_1205,N_24047,N_24371);
nand UO_1206 (O_1206,N_24626,N_24546);
nor UO_1207 (O_1207,N_24944,N_24587);
and UO_1208 (O_1208,N_24965,N_23643);
or UO_1209 (O_1209,N_24664,N_22517);
nand UO_1210 (O_1210,N_23314,N_23075);
or UO_1211 (O_1211,N_24624,N_23952);
or UO_1212 (O_1212,N_23341,N_24641);
and UO_1213 (O_1213,N_22698,N_24464);
nand UO_1214 (O_1214,N_24091,N_24192);
nor UO_1215 (O_1215,N_23222,N_22857);
and UO_1216 (O_1216,N_23023,N_23505);
nor UO_1217 (O_1217,N_23645,N_23215);
nor UO_1218 (O_1218,N_23349,N_23919);
and UO_1219 (O_1219,N_24607,N_23590);
and UO_1220 (O_1220,N_23487,N_24509);
nand UO_1221 (O_1221,N_23223,N_23768);
or UO_1222 (O_1222,N_23740,N_24874);
nor UO_1223 (O_1223,N_24325,N_23943);
nand UO_1224 (O_1224,N_23196,N_22686);
and UO_1225 (O_1225,N_23035,N_24023);
or UO_1226 (O_1226,N_24476,N_23022);
and UO_1227 (O_1227,N_24367,N_22935);
nand UO_1228 (O_1228,N_23844,N_23584);
or UO_1229 (O_1229,N_23198,N_23637);
or UO_1230 (O_1230,N_23010,N_24381);
nand UO_1231 (O_1231,N_24154,N_24369);
nand UO_1232 (O_1232,N_24698,N_23059);
or UO_1233 (O_1233,N_22505,N_22750);
or UO_1234 (O_1234,N_24049,N_24317);
nor UO_1235 (O_1235,N_23835,N_22590);
nor UO_1236 (O_1236,N_24639,N_24754);
nand UO_1237 (O_1237,N_22987,N_22835);
nand UO_1238 (O_1238,N_24606,N_22657);
nor UO_1239 (O_1239,N_22911,N_23447);
and UO_1240 (O_1240,N_23161,N_24164);
or UO_1241 (O_1241,N_23734,N_22702);
and UO_1242 (O_1242,N_24385,N_23363);
or UO_1243 (O_1243,N_23380,N_22524);
nand UO_1244 (O_1244,N_23397,N_22635);
nor UO_1245 (O_1245,N_24902,N_23933);
and UO_1246 (O_1246,N_24493,N_24613);
xor UO_1247 (O_1247,N_24181,N_23700);
nand UO_1248 (O_1248,N_24725,N_24803);
nor UO_1249 (O_1249,N_23641,N_23372);
or UO_1250 (O_1250,N_23641,N_22542);
nor UO_1251 (O_1251,N_24959,N_24745);
nor UO_1252 (O_1252,N_23839,N_22725);
nand UO_1253 (O_1253,N_22503,N_23080);
xor UO_1254 (O_1254,N_23399,N_24071);
and UO_1255 (O_1255,N_23973,N_23432);
and UO_1256 (O_1256,N_24814,N_24703);
nor UO_1257 (O_1257,N_22745,N_24180);
and UO_1258 (O_1258,N_24595,N_24112);
nand UO_1259 (O_1259,N_22963,N_24024);
or UO_1260 (O_1260,N_24547,N_23175);
and UO_1261 (O_1261,N_23638,N_23252);
nand UO_1262 (O_1262,N_23440,N_24858);
or UO_1263 (O_1263,N_22650,N_24689);
nor UO_1264 (O_1264,N_23800,N_24515);
nand UO_1265 (O_1265,N_24291,N_24122);
or UO_1266 (O_1266,N_22932,N_24133);
xor UO_1267 (O_1267,N_23118,N_24858);
nand UO_1268 (O_1268,N_22847,N_23399);
or UO_1269 (O_1269,N_22704,N_24482);
nor UO_1270 (O_1270,N_24304,N_22619);
xnor UO_1271 (O_1271,N_24016,N_23961);
or UO_1272 (O_1272,N_23523,N_23734);
or UO_1273 (O_1273,N_24853,N_23947);
or UO_1274 (O_1274,N_23015,N_23871);
nor UO_1275 (O_1275,N_22888,N_24540);
and UO_1276 (O_1276,N_22624,N_22919);
or UO_1277 (O_1277,N_24370,N_24015);
nor UO_1278 (O_1278,N_22921,N_24932);
nand UO_1279 (O_1279,N_22554,N_22620);
nor UO_1280 (O_1280,N_23935,N_23756);
nor UO_1281 (O_1281,N_23330,N_23348);
and UO_1282 (O_1282,N_23299,N_22532);
nand UO_1283 (O_1283,N_24976,N_22826);
and UO_1284 (O_1284,N_23244,N_24299);
nand UO_1285 (O_1285,N_22629,N_24279);
or UO_1286 (O_1286,N_24474,N_23869);
nand UO_1287 (O_1287,N_22690,N_23616);
and UO_1288 (O_1288,N_24679,N_22768);
and UO_1289 (O_1289,N_22972,N_22585);
or UO_1290 (O_1290,N_24318,N_23082);
nand UO_1291 (O_1291,N_24668,N_22677);
nand UO_1292 (O_1292,N_24731,N_24721);
nand UO_1293 (O_1293,N_24002,N_23504);
nor UO_1294 (O_1294,N_24247,N_23030);
nand UO_1295 (O_1295,N_22740,N_23716);
nor UO_1296 (O_1296,N_24921,N_24616);
and UO_1297 (O_1297,N_22971,N_24957);
or UO_1298 (O_1298,N_24084,N_22613);
nor UO_1299 (O_1299,N_24739,N_23075);
and UO_1300 (O_1300,N_23691,N_24981);
or UO_1301 (O_1301,N_24040,N_24888);
or UO_1302 (O_1302,N_22847,N_22616);
and UO_1303 (O_1303,N_22728,N_24794);
or UO_1304 (O_1304,N_23821,N_23733);
and UO_1305 (O_1305,N_22863,N_23955);
or UO_1306 (O_1306,N_23959,N_22966);
and UO_1307 (O_1307,N_23387,N_24984);
or UO_1308 (O_1308,N_23320,N_22894);
nand UO_1309 (O_1309,N_23293,N_24821);
and UO_1310 (O_1310,N_24996,N_24662);
or UO_1311 (O_1311,N_24139,N_24217);
nand UO_1312 (O_1312,N_24064,N_22636);
nand UO_1313 (O_1313,N_24629,N_24864);
and UO_1314 (O_1314,N_22762,N_24461);
and UO_1315 (O_1315,N_24425,N_24686);
nor UO_1316 (O_1316,N_23565,N_23803);
nor UO_1317 (O_1317,N_23719,N_23196);
and UO_1318 (O_1318,N_24020,N_22689);
nand UO_1319 (O_1319,N_23970,N_22779);
and UO_1320 (O_1320,N_23288,N_24659);
nor UO_1321 (O_1321,N_24748,N_24949);
and UO_1322 (O_1322,N_23624,N_24565);
nor UO_1323 (O_1323,N_24004,N_23543);
and UO_1324 (O_1324,N_23385,N_24298);
or UO_1325 (O_1325,N_24723,N_24831);
and UO_1326 (O_1326,N_23717,N_24709);
nand UO_1327 (O_1327,N_22675,N_24734);
and UO_1328 (O_1328,N_23438,N_24727);
or UO_1329 (O_1329,N_23612,N_22765);
or UO_1330 (O_1330,N_24801,N_24726);
xnor UO_1331 (O_1331,N_22820,N_23569);
nor UO_1332 (O_1332,N_22536,N_24041);
nand UO_1333 (O_1333,N_23048,N_24454);
or UO_1334 (O_1334,N_23783,N_24789);
nor UO_1335 (O_1335,N_24073,N_23372);
and UO_1336 (O_1336,N_23719,N_23825);
or UO_1337 (O_1337,N_23089,N_24136);
or UO_1338 (O_1338,N_23985,N_24403);
nor UO_1339 (O_1339,N_22669,N_22661);
or UO_1340 (O_1340,N_22840,N_24919);
nor UO_1341 (O_1341,N_23169,N_23894);
nand UO_1342 (O_1342,N_23468,N_22665);
nor UO_1343 (O_1343,N_22509,N_24732);
and UO_1344 (O_1344,N_24245,N_24137);
nor UO_1345 (O_1345,N_24572,N_24802);
nand UO_1346 (O_1346,N_23038,N_24157);
xor UO_1347 (O_1347,N_22864,N_24885);
nand UO_1348 (O_1348,N_22716,N_23539);
nor UO_1349 (O_1349,N_23505,N_23633);
and UO_1350 (O_1350,N_23540,N_24136);
or UO_1351 (O_1351,N_23328,N_22838);
or UO_1352 (O_1352,N_23232,N_24122);
nor UO_1353 (O_1353,N_24134,N_22597);
or UO_1354 (O_1354,N_24937,N_24929);
nand UO_1355 (O_1355,N_23949,N_22548);
and UO_1356 (O_1356,N_23104,N_23265);
or UO_1357 (O_1357,N_24360,N_24226);
nand UO_1358 (O_1358,N_23910,N_24743);
nand UO_1359 (O_1359,N_24831,N_23816);
nand UO_1360 (O_1360,N_24990,N_24321);
or UO_1361 (O_1361,N_22691,N_23878);
and UO_1362 (O_1362,N_23773,N_22952);
and UO_1363 (O_1363,N_23344,N_23900);
nand UO_1364 (O_1364,N_24328,N_24550);
or UO_1365 (O_1365,N_22696,N_23756);
or UO_1366 (O_1366,N_23055,N_24029);
nand UO_1367 (O_1367,N_22656,N_24678);
nand UO_1368 (O_1368,N_24524,N_22552);
or UO_1369 (O_1369,N_22747,N_24461);
nor UO_1370 (O_1370,N_24945,N_23397);
and UO_1371 (O_1371,N_22896,N_24248);
and UO_1372 (O_1372,N_24280,N_22976);
or UO_1373 (O_1373,N_23843,N_22992);
and UO_1374 (O_1374,N_23991,N_24060);
nor UO_1375 (O_1375,N_23401,N_23970);
nand UO_1376 (O_1376,N_23109,N_23469);
or UO_1377 (O_1377,N_23202,N_22737);
and UO_1378 (O_1378,N_22582,N_23291);
or UO_1379 (O_1379,N_24199,N_24055);
nor UO_1380 (O_1380,N_24803,N_23523);
nor UO_1381 (O_1381,N_22537,N_23501);
nand UO_1382 (O_1382,N_23654,N_23157);
nand UO_1383 (O_1383,N_24303,N_23620);
or UO_1384 (O_1384,N_24399,N_24739);
and UO_1385 (O_1385,N_24020,N_22644);
nand UO_1386 (O_1386,N_24866,N_23613);
or UO_1387 (O_1387,N_24387,N_24976);
nor UO_1388 (O_1388,N_24473,N_24387);
or UO_1389 (O_1389,N_24873,N_22784);
or UO_1390 (O_1390,N_24804,N_23662);
nand UO_1391 (O_1391,N_23211,N_23581);
or UO_1392 (O_1392,N_24536,N_22628);
nor UO_1393 (O_1393,N_24793,N_23428);
nand UO_1394 (O_1394,N_24733,N_24908);
and UO_1395 (O_1395,N_22521,N_24906);
nor UO_1396 (O_1396,N_23418,N_24430);
nor UO_1397 (O_1397,N_22875,N_23483);
nor UO_1398 (O_1398,N_22730,N_23849);
nor UO_1399 (O_1399,N_22926,N_24984);
or UO_1400 (O_1400,N_23272,N_24579);
nor UO_1401 (O_1401,N_24674,N_23373);
or UO_1402 (O_1402,N_24459,N_24806);
nand UO_1403 (O_1403,N_23219,N_24278);
or UO_1404 (O_1404,N_23487,N_23229);
and UO_1405 (O_1405,N_22922,N_23359);
and UO_1406 (O_1406,N_23394,N_22921);
xor UO_1407 (O_1407,N_24827,N_23452);
and UO_1408 (O_1408,N_24968,N_24115);
or UO_1409 (O_1409,N_24491,N_22743);
and UO_1410 (O_1410,N_24795,N_24199);
and UO_1411 (O_1411,N_24382,N_24857);
and UO_1412 (O_1412,N_23719,N_22549);
or UO_1413 (O_1413,N_23153,N_23322);
and UO_1414 (O_1414,N_23398,N_23041);
nor UO_1415 (O_1415,N_24987,N_23734);
and UO_1416 (O_1416,N_24175,N_22872);
or UO_1417 (O_1417,N_24879,N_23133);
nand UO_1418 (O_1418,N_23143,N_23569);
and UO_1419 (O_1419,N_24622,N_24633);
nor UO_1420 (O_1420,N_23604,N_24467);
nand UO_1421 (O_1421,N_24219,N_23510);
and UO_1422 (O_1422,N_22630,N_23978);
and UO_1423 (O_1423,N_23659,N_24597);
or UO_1424 (O_1424,N_23227,N_24085);
and UO_1425 (O_1425,N_24238,N_24526);
and UO_1426 (O_1426,N_22716,N_22561);
nor UO_1427 (O_1427,N_22887,N_24668);
nand UO_1428 (O_1428,N_23319,N_22837);
nor UO_1429 (O_1429,N_23479,N_23483);
and UO_1430 (O_1430,N_24363,N_24164);
and UO_1431 (O_1431,N_24043,N_22597);
or UO_1432 (O_1432,N_23877,N_23555);
and UO_1433 (O_1433,N_22781,N_22767);
or UO_1434 (O_1434,N_23279,N_23089);
and UO_1435 (O_1435,N_23696,N_24760);
nand UO_1436 (O_1436,N_23022,N_24856);
or UO_1437 (O_1437,N_23116,N_23793);
nor UO_1438 (O_1438,N_24485,N_22742);
nand UO_1439 (O_1439,N_23508,N_24656);
or UO_1440 (O_1440,N_24455,N_22795);
or UO_1441 (O_1441,N_24698,N_24097);
nand UO_1442 (O_1442,N_24297,N_24269);
nor UO_1443 (O_1443,N_23108,N_23312);
and UO_1444 (O_1444,N_22740,N_23140);
and UO_1445 (O_1445,N_24975,N_24218);
nand UO_1446 (O_1446,N_24474,N_24463);
nand UO_1447 (O_1447,N_24257,N_24035);
nor UO_1448 (O_1448,N_24847,N_23690);
nor UO_1449 (O_1449,N_24609,N_23984);
nand UO_1450 (O_1450,N_23344,N_22716);
nand UO_1451 (O_1451,N_22563,N_24867);
or UO_1452 (O_1452,N_24825,N_24180);
nor UO_1453 (O_1453,N_24976,N_24448);
nor UO_1454 (O_1454,N_23245,N_23638);
or UO_1455 (O_1455,N_23391,N_22865);
nor UO_1456 (O_1456,N_24599,N_23199);
or UO_1457 (O_1457,N_23381,N_24525);
nor UO_1458 (O_1458,N_22606,N_23970);
and UO_1459 (O_1459,N_23848,N_23114);
and UO_1460 (O_1460,N_23664,N_22862);
or UO_1461 (O_1461,N_24110,N_23173);
nor UO_1462 (O_1462,N_23902,N_24304);
or UO_1463 (O_1463,N_24112,N_23308);
or UO_1464 (O_1464,N_23514,N_24366);
and UO_1465 (O_1465,N_24703,N_24294);
nand UO_1466 (O_1466,N_23604,N_23155);
nor UO_1467 (O_1467,N_24635,N_22642);
nor UO_1468 (O_1468,N_23085,N_24491);
nand UO_1469 (O_1469,N_24216,N_23216);
and UO_1470 (O_1470,N_24495,N_23943);
and UO_1471 (O_1471,N_23181,N_24848);
and UO_1472 (O_1472,N_24433,N_23671);
and UO_1473 (O_1473,N_24989,N_24272);
nand UO_1474 (O_1474,N_24193,N_22526);
nor UO_1475 (O_1475,N_24733,N_24393);
and UO_1476 (O_1476,N_23350,N_24746);
nor UO_1477 (O_1477,N_24469,N_23932);
and UO_1478 (O_1478,N_22761,N_22939);
and UO_1479 (O_1479,N_23284,N_24115);
nor UO_1480 (O_1480,N_22629,N_24723);
nor UO_1481 (O_1481,N_24646,N_23577);
or UO_1482 (O_1482,N_24447,N_24298);
nand UO_1483 (O_1483,N_24841,N_23510);
nor UO_1484 (O_1484,N_24024,N_24362);
nor UO_1485 (O_1485,N_23339,N_23548);
or UO_1486 (O_1486,N_23585,N_24830);
nand UO_1487 (O_1487,N_24413,N_24266);
and UO_1488 (O_1488,N_22729,N_24050);
nand UO_1489 (O_1489,N_24809,N_23422);
nand UO_1490 (O_1490,N_23194,N_23322);
nand UO_1491 (O_1491,N_23947,N_24440);
nor UO_1492 (O_1492,N_23157,N_23877);
and UO_1493 (O_1493,N_23652,N_22748);
or UO_1494 (O_1494,N_24102,N_23507);
and UO_1495 (O_1495,N_22796,N_24933);
nor UO_1496 (O_1496,N_24393,N_24932);
nor UO_1497 (O_1497,N_24590,N_23962);
and UO_1498 (O_1498,N_24522,N_24593);
nor UO_1499 (O_1499,N_23123,N_24634);
nor UO_1500 (O_1500,N_22991,N_23133);
or UO_1501 (O_1501,N_22526,N_24641);
nand UO_1502 (O_1502,N_23367,N_22943);
and UO_1503 (O_1503,N_23336,N_24785);
nand UO_1504 (O_1504,N_24600,N_24210);
nand UO_1505 (O_1505,N_24015,N_24781);
and UO_1506 (O_1506,N_22948,N_22659);
nor UO_1507 (O_1507,N_23061,N_23398);
nor UO_1508 (O_1508,N_22834,N_22639);
or UO_1509 (O_1509,N_23684,N_24085);
nor UO_1510 (O_1510,N_22798,N_22521);
or UO_1511 (O_1511,N_23620,N_24096);
nor UO_1512 (O_1512,N_23618,N_23322);
nor UO_1513 (O_1513,N_23594,N_23201);
nor UO_1514 (O_1514,N_23105,N_24992);
or UO_1515 (O_1515,N_23642,N_23726);
or UO_1516 (O_1516,N_23245,N_24078);
nand UO_1517 (O_1517,N_22750,N_23134);
nand UO_1518 (O_1518,N_24659,N_24588);
and UO_1519 (O_1519,N_22961,N_24111);
and UO_1520 (O_1520,N_23346,N_24513);
and UO_1521 (O_1521,N_23594,N_24403);
or UO_1522 (O_1522,N_24994,N_24286);
and UO_1523 (O_1523,N_23185,N_23107);
nor UO_1524 (O_1524,N_23713,N_23552);
nand UO_1525 (O_1525,N_23277,N_23882);
nand UO_1526 (O_1526,N_22556,N_24348);
nand UO_1527 (O_1527,N_22673,N_23329);
nor UO_1528 (O_1528,N_22871,N_23904);
or UO_1529 (O_1529,N_22540,N_22938);
and UO_1530 (O_1530,N_23472,N_24645);
nand UO_1531 (O_1531,N_22946,N_23383);
nor UO_1532 (O_1532,N_24614,N_23327);
and UO_1533 (O_1533,N_22574,N_22663);
xnor UO_1534 (O_1534,N_23381,N_23823);
and UO_1535 (O_1535,N_24994,N_24805);
nor UO_1536 (O_1536,N_22766,N_24178);
and UO_1537 (O_1537,N_23177,N_22728);
or UO_1538 (O_1538,N_22896,N_22703);
nand UO_1539 (O_1539,N_23042,N_24809);
nand UO_1540 (O_1540,N_24483,N_23822);
nor UO_1541 (O_1541,N_24643,N_24855);
nor UO_1542 (O_1542,N_24997,N_23080);
and UO_1543 (O_1543,N_23660,N_24380);
and UO_1544 (O_1544,N_24740,N_24987);
or UO_1545 (O_1545,N_24102,N_22578);
nor UO_1546 (O_1546,N_23043,N_23192);
and UO_1547 (O_1547,N_22722,N_24140);
nand UO_1548 (O_1548,N_24245,N_24323);
nor UO_1549 (O_1549,N_23761,N_22660);
xor UO_1550 (O_1550,N_22874,N_23049);
or UO_1551 (O_1551,N_23659,N_24696);
nor UO_1552 (O_1552,N_24946,N_24926);
nor UO_1553 (O_1553,N_22952,N_24770);
and UO_1554 (O_1554,N_23216,N_23990);
nand UO_1555 (O_1555,N_23775,N_22950);
and UO_1556 (O_1556,N_23553,N_23476);
nor UO_1557 (O_1557,N_23270,N_23324);
and UO_1558 (O_1558,N_23225,N_22770);
nand UO_1559 (O_1559,N_23412,N_23787);
or UO_1560 (O_1560,N_23900,N_24442);
or UO_1561 (O_1561,N_24390,N_23082);
nand UO_1562 (O_1562,N_23088,N_23982);
nand UO_1563 (O_1563,N_22749,N_22654);
nor UO_1564 (O_1564,N_24424,N_24966);
or UO_1565 (O_1565,N_23331,N_24648);
and UO_1566 (O_1566,N_23929,N_23434);
nand UO_1567 (O_1567,N_23690,N_22521);
nor UO_1568 (O_1568,N_23381,N_24761);
and UO_1569 (O_1569,N_23945,N_22740);
and UO_1570 (O_1570,N_24758,N_23264);
and UO_1571 (O_1571,N_24888,N_24096);
nor UO_1572 (O_1572,N_23031,N_22649);
nand UO_1573 (O_1573,N_23629,N_24160);
nand UO_1574 (O_1574,N_22838,N_23012);
or UO_1575 (O_1575,N_24095,N_23613);
or UO_1576 (O_1576,N_24979,N_23542);
nor UO_1577 (O_1577,N_24392,N_23811);
nor UO_1578 (O_1578,N_22660,N_24398);
or UO_1579 (O_1579,N_22931,N_24598);
and UO_1580 (O_1580,N_23401,N_24657);
or UO_1581 (O_1581,N_24726,N_23549);
and UO_1582 (O_1582,N_24673,N_24679);
nand UO_1583 (O_1583,N_22534,N_24091);
nor UO_1584 (O_1584,N_24533,N_23029);
nor UO_1585 (O_1585,N_22836,N_24037);
or UO_1586 (O_1586,N_22515,N_23719);
nand UO_1587 (O_1587,N_22667,N_23210);
nand UO_1588 (O_1588,N_23149,N_23518);
or UO_1589 (O_1589,N_24005,N_24800);
nand UO_1590 (O_1590,N_23512,N_23090);
nor UO_1591 (O_1591,N_23853,N_22636);
nor UO_1592 (O_1592,N_24957,N_23674);
nand UO_1593 (O_1593,N_24156,N_22932);
nand UO_1594 (O_1594,N_22705,N_24884);
nor UO_1595 (O_1595,N_23431,N_24497);
and UO_1596 (O_1596,N_23460,N_24056);
or UO_1597 (O_1597,N_23640,N_23220);
nor UO_1598 (O_1598,N_23580,N_23482);
nand UO_1599 (O_1599,N_22882,N_24425);
and UO_1600 (O_1600,N_23798,N_22505);
nand UO_1601 (O_1601,N_24613,N_23580);
nor UO_1602 (O_1602,N_22979,N_23336);
or UO_1603 (O_1603,N_24614,N_24247);
or UO_1604 (O_1604,N_24307,N_23241);
nor UO_1605 (O_1605,N_24121,N_23240);
nor UO_1606 (O_1606,N_22604,N_22641);
nor UO_1607 (O_1607,N_23392,N_24727);
nand UO_1608 (O_1608,N_23203,N_23909);
nor UO_1609 (O_1609,N_23758,N_22753);
or UO_1610 (O_1610,N_22746,N_24951);
nand UO_1611 (O_1611,N_24721,N_23089);
or UO_1612 (O_1612,N_24453,N_23528);
nand UO_1613 (O_1613,N_24882,N_23986);
or UO_1614 (O_1614,N_23793,N_24674);
or UO_1615 (O_1615,N_23298,N_24996);
and UO_1616 (O_1616,N_22877,N_22707);
and UO_1617 (O_1617,N_23119,N_24439);
or UO_1618 (O_1618,N_22572,N_24917);
nand UO_1619 (O_1619,N_23256,N_22849);
or UO_1620 (O_1620,N_24992,N_24366);
nor UO_1621 (O_1621,N_23388,N_24180);
or UO_1622 (O_1622,N_24934,N_23452);
or UO_1623 (O_1623,N_24123,N_24730);
nor UO_1624 (O_1624,N_22993,N_24077);
nand UO_1625 (O_1625,N_22798,N_23139);
nor UO_1626 (O_1626,N_24485,N_24499);
and UO_1627 (O_1627,N_24375,N_23838);
or UO_1628 (O_1628,N_23051,N_23144);
nand UO_1629 (O_1629,N_23971,N_22833);
and UO_1630 (O_1630,N_23354,N_23548);
or UO_1631 (O_1631,N_23071,N_22561);
and UO_1632 (O_1632,N_22737,N_22558);
or UO_1633 (O_1633,N_24469,N_23435);
nor UO_1634 (O_1634,N_24055,N_24645);
nor UO_1635 (O_1635,N_23137,N_23897);
xnor UO_1636 (O_1636,N_23426,N_23497);
or UO_1637 (O_1637,N_22953,N_24061);
nor UO_1638 (O_1638,N_23222,N_23955);
nand UO_1639 (O_1639,N_24275,N_23526);
nand UO_1640 (O_1640,N_23675,N_24486);
nand UO_1641 (O_1641,N_24228,N_22988);
nand UO_1642 (O_1642,N_22520,N_22722);
nor UO_1643 (O_1643,N_24244,N_24278);
nor UO_1644 (O_1644,N_24486,N_24409);
nand UO_1645 (O_1645,N_23584,N_23441);
or UO_1646 (O_1646,N_22799,N_24257);
and UO_1647 (O_1647,N_22930,N_24917);
nand UO_1648 (O_1648,N_23951,N_22606);
nor UO_1649 (O_1649,N_23442,N_23903);
nand UO_1650 (O_1650,N_24903,N_24917);
and UO_1651 (O_1651,N_22610,N_24293);
nor UO_1652 (O_1652,N_23087,N_22794);
or UO_1653 (O_1653,N_24308,N_23243);
nand UO_1654 (O_1654,N_22943,N_23535);
and UO_1655 (O_1655,N_23360,N_23343);
or UO_1656 (O_1656,N_22744,N_24481);
nand UO_1657 (O_1657,N_24186,N_24273);
nand UO_1658 (O_1658,N_22558,N_22705);
and UO_1659 (O_1659,N_22673,N_23652);
nand UO_1660 (O_1660,N_22615,N_24049);
nor UO_1661 (O_1661,N_24500,N_22976);
and UO_1662 (O_1662,N_23131,N_22800);
xnor UO_1663 (O_1663,N_24519,N_22931);
and UO_1664 (O_1664,N_22503,N_24944);
nor UO_1665 (O_1665,N_23312,N_24834);
or UO_1666 (O_1666,N_22712,N_23361);
or UO_1667 (O_1667,N_22789,N_23768);
nor UO_1668 (O_1668,N_22527,N_22992);
and UO_1669 (O_1669,N_22661,N_24528);
or UO_1670 (O_1670,N_24354,N_23478);
or UO_1671 (O_1671,N_23119,N_24096);
or UO_1672 (O_1672,N_24507,N_24590);
nor UO_1673 (O_1673,N_24721,N_24107);
nand UO_1674 (O_1674,N_23185,N_23031);
nand UO_1675 (O_1675,N_24747,N_23121);
or UO_1676 (O_1676,N_23442,N_24231);
or UO_1677 (O_1677,N_22742,N_23674);
or UO_1678 (O_1678,N_24044,N_24302);
nand UO_1679 (O_1679,N_24903,N_23357);
nand UO_1680 (O_1680,N_24851,N_24582);
nor UO_1681 (O_1681,N_24240,N_23777);
xor UO_1682 (O_1682,N_23434,N_23254);
or UO_1683 (O_1683,N_22646,N_24782);
nand UO_1684 (O_1684,N_24339,N_23908);
nand UO_1685 (O_1685,N_22523,N_23129);
nand UO_1686 (O_1686,N_23240,N_22913);
nand UO_1687 (O_1687,N_23868,N_22523);
and UO_1688 (O_1688,N_24375,N_22874);
or UO_1689 (O_1689,N_24834,N_23247);
nor UO_1690 (O_1690,N_24201,N_24168);
nor UO_1691 (O_1691,N_24737,N_23043);
and UO_1692 (O_1692,N_23281,N_24526);
nand UO_1693 (O_1693,N_22599,N_23807);
and UO_1694 (O_1694,N_24333,N_23761);
or UO_1695 (O_1695,N_23838,N_22723);
nand UO_1696 (O_1696,N_23753,N_23373);
nand UO_1697 (O_1697,N_22876,N_23869);
or UO_1698 (O_1698,N_24809,N_24386);
or UO_1699 (O_1699,N_23316,N_24177);
nor UO_1700 (O_1700,N_24526,N_23370);
nor UO_1701 (O_1701,N_23324,N_22612);
or UO_1702 (O_1702,N_23869,N_24057);
and UO_1703 (O_1703,N_23656,N_23437);
and UO_1704 (O_1704,N_22521,N_23946);
nor UO_1705 (O_1705,N_24059,N_23718);
nand UO_1706 (O_1706,N_23035,N_24312);
nor UO_1707 (O_1707,N_23166,N_23007);
nor UO_1708 (O_1708,N_22566,N_23070);
or UO_1709 (O_1709,N_23185,N_23791);
and UO_1710 (O_1710,N_23516,N_24945);
nor UO_1711 (O_1711,N_24074,N_24388);
or UO_1712 (O_1712,N_23518,N_23876);
or UO_1713 (O_1713,N_23667,N_23288);
and UO_1714 (O_1714,N_22520,N_24223);
nand UO_1715 (O_1715,N_24795,N_24912);
and UO_1716 (O_1716,N_22660,N_23263);
nand UO_1717 (O_1717,N_22656,N_23627);
nand UO_1718 (O_1718,N_23184,N_22912);
nor UO_1719 (O_1719,N_23311,N_23310);
nor UO_1720 (O_1720,N_22697,N_24810);
nand UO_1721 (O_1721,N_22752,N_24492);
or UO_1722 (O_1722,N_24905,N_23402);
nand UO_1723 (O_1723,N_23402,N_22942);
and UO_1724 (O_1724,N_22925,N_22761);
and UO_1725 (O_1725,N_23499,N_23756);
nand UO_1726 (O_1726,N_24007,N_24523);
nor UO_1727 (O_1727,N_24509,N_23155);
and UO_1728 (O_1728,N_22821,N_23066);
nor UO_1729 (O_1729,N_23379,N_22958);
or UO_1730 (O_1730,N_23632,N_24688);
nand UO_1731 (O_1731,N_23494,N_23305);
nor UO_1732 (O_1732,N_24687,N_22512);
and UO_1733 (O_1733,N_23165,N_24575);
nand UO_1734 (O_1734,N_22724,N_22944);
nor UO_1735 (O_1735,N_23011,N_24542);
nand UO_1736 (O_1736,N_23782,N_23613);
and UO_1737 (O_1737,N_23758,N_24783);
nand UO_1738 (O_1738,N_22712,N_24052);
nand UO_1739 (O_1739,N_24828,N_23245);
nor UO_1740 (O_1740,N_24242,N_23449);
nand UO_1741 (O_1741,N_22739,N_22607);
or UO_1742 (O_1742,N_24931,N_23344);
nand UO_1743 (O_1743,N_24084,N_23158);
nand UO_1744 (O_1744,N_22594,N_23558);
or UO_1745 (O_1745,N_24968,N_24609);
xor UO_1746 (O_1746,N_24070,N_24329);
nor UO_1747 (O_1747,N_24842,N_24154);
nand UO_1748 (O_1748,N_23725,N_23019);
nand UO_1749 (O_1749,N_23800,N_23544);
and UO_1750 (O_1750,N_22607,N_23167);
nand UO_1751 (O_1751,N_24595,N_24784);
nor UO_1752 (O_1752,N_23164,N_24702);
nand UO_1753 (O_1753,N_22679,N_23749);
or UO_1754 (O_1754,N_24756,N_23134);
and UO_1755 (O_1755,N_24760,N_23433);
and UO_1756 (O_1756,N_24005,N_24127);
or UO_1757 (O_1757,N_24596,N_23443);
nand UO_1758 (O_1758,N_23755,N_24451);
and UO_1759 (O_1759,N_22909,N_23905);
xnor UO_1760 (O_1760,N_22597,N_24787);
nand UO_1761 (O_1761,N_24246,N_24435);
or UO_1762 (O_1762,N_24964,N_23834);
or UO_1763 (O_1763,N_24636,N_22679);
nand UO_1764 (O_1764,N_22824,N_22561);
and UO_1765 (O_1765,N_22530,N_23913);
nor UO_1766 (O_1766,N_24037,N_24978);
or UO_1767 (O_1767,N_24904,N_22999);
nand UO_1768 (O_1768,N_23772,N_23606);
nand UO_1769 (O_1769,N_22600,N_24392);
or UO_1770 (O_1770,N_22631,N_22604);
nor UO_1771 (O_1771,N_22912,N_24563);
nand UO_1772 (O_1772,N_23537,N_24455);
nor UO_1773 (O_1773,N_23411,N_23143);
or UO_1774 (O_1774,N_23203,N_23663);
nor UO_1775 (O_1775,N_24781,N_24582);
nand UO_1776 (O_1776,N_22500,N_23809);
nand UO_1777 (O_1777,N_22565,N_23316);
or UO_1778 (O_1778,N_24632,N_23085);
nor UO_1779 (O_1779,N_23452,N_22930);
and UO_1780 (O_1780,N_24466,N_23445);
nor UO_1781 (O_1781,N_23540,N_24345);
nor UO_1782 (O_1782,N_22709,N_23928);
or UO_1783 (O_1783,N_24589,N_22947);
and UO_1784 (O_1784,N_23388,N_24632);
nand UO_1785 (O_1785,N_22524,N_23418);
or UO_1786 (O_1786,N_24693,N_24632);
nand UO_1787 (O_1787,N_22583,N_23630);
nor UO_1788 (O_1788,N_24665,N_24174);
nor UO_1789 (O_1789,N_22583,N_24344);
and UO_1790 (O_1790,N_22869,N_23119);
nor UO_1791 (O_1791,N_24298,N_24564);
nor UO_1792 (O_1792,N_23572,N_22539);
nor UO_1793 (O_1793,N_22573,N_24622);
and UO_1794 (O_1794,N_24168,N_24361);
or UO_1795 (O_1795,N_24474,N_23945);
or UO_1796 (O_1796,N_23005,N_23990);
and UO_1797 (O_1797,N_22926,N_24602);
nor UO_1798 (O_1798,N_23441,N_24049);
or UO_1799 (O_1799,N_22707,N_23387);
nor UO_1800 (O_1800,N_22676,N_22667);
or UO_1801 (O_1801,N_23899,N_24196);
and UO_1802 (O_1802,N_24894,N_24513);
or UO_1803 (O_1803,N_23721,N_23539);
nand UO_1804 (O_1804,N_23873,N_24238);
nor UO_1805 (O_1805,N_24848,N_23423);
and UO_1806 (O_1806,N_23611,N_22905);
nor UO_1807 (O_1807,N_24269,N_23734);
nand UO_1808 (O_1808,N_24840,N_24151);
nand UO_1809 (O_1809,N_24271,N_24296);
and UO_1810 (O_1810,N_22902,N_24352);
and UO_1811 (O_1811,N_24930,N_24286);
nand UO_1812 (O_1812,N_23050,N_24696);
and UO_1813 (O_1813,N_23164,N_23979);
nor UO_1814 (O_1814,N_22888,N_24784);
nor UO_1815 (O_1815,N_24260,N_24292);
or UO_1816 (O_1816,N_22815,N_23201);
and UO_1817 (O_1817,N_23632,N_23131);
nor UO_1818 (O_1818,N_23350,N_24120);
and UO_1819 (O_1819,N_24427,N_23238);
nor UO_1820 (O_1820,N_23808,N_22734);
nor UO_1821 (O_1821,N_23259,N_24057);
nor UO_1822 (O_1822,N_23815,N_22695);
or UO_1823 (O_1823,N_22740,N_22543);
or UO_1824 (O_1824,N_24614,N_23083);
nand UO_1825 (O_1825,N_23370,N_23604);
nand UO_1826 (O_1826,N_24578,N_23948);
and UO_1827 (O_1827,N_23272,N_24344);
and UO_1828 (O_1828,N_24704,N_22727);
nand UO_1829 (O_1829,N_24703,N_23600);
nand UO_1830 (O_1830,N_24834,N_24341);
nor UO_1831 (O_1831,N_23915,N_24917);
nor UO_1832 (O_1832,N_22657,N_23172);
and UO_1833 (O_1833,N_24556,N_24719);
nor UO_1834 (O_1834,N_23999,N_23731);
nor UO_1835 (O_1835,N_22603,N_24533);
nand UO_1836 (O_1836,N_22845,N_24699);
nand UO_1837 (O_1837,N_23619,N_23188);
and UO_1838 (O_1838,N_24206,N_22545);
and UO_1839 (O_1839,N_24517,N_23662);
nor UO_1840 (O_1840,N_24389,N_22622);
and UO_1841 (O_1841,N_24121,N_24316);
nor UO_1842 (O_1842,N_23996,N_24959);
nand UO_1843 (O_1843,N_22528,N_24290);
or UO_1844 (O_1844,N_24796,N_24825);
and UO_1845 (O_1845,N_24157,N_23773);
nor UO_1846 (O_1846,N_23677,N_22512);
nand UO_1847 (O_1847,N_23986,N_23513);
nor UO_1848 (O_1848,N_22565,N_24273);
or UO_1849 (O_1849,N_24793,N_22926);
nand UO_1850 (O_1850,N_23839,N_24473);
nor UO_1851 (O_1851,N_22537,N_24559);
or UO_1852 (O_1852,N_23363,N_22962);
nor UO_1853 (O_1853,N_24168,N_22574);
nand UO_1854 (O_1854,N_23154,N_23518);
nand UO_1855 (O_1855,N_23153,N_23784);
nand UO_1856 (O_1856,N_24220,N_23551);
and UO_1857 (O_1857,N_24888,N_23853);
nand UO_1858 (O_1858,N_24511,N_23190);
nand UO_1859 (O_1859,N_24666,N_22505);
nand UO_1860 (O_1860,N_23710,N_22697);
or UO_1861 (O_1861,N_24377,N_23381);
or UO_1862 (O_1862,N_22652,N_23486);
nor UO_1863 (O_1863,N_24729,N_23117);
nor UO_1864 (O_1864,N_24398,N_23199);
or UO_1865 (O_1865,N_23010,N_24528);
or UO_1866 (O_1866,N_24845,N_24267);
or UO_1867 (O_1867,N_24359,N_22573);
nor UO_1868 (O_1868,N_24723,N_22722);
nand UO_1869 (O_1869,N_23150,N_23197);
nand UO_1870 (O_1870,N_23714,N_24076);
nand UO_1871 (O_1871,N_23787,N_22818);
nand UO_1872 (O_1872,N_22793,N_23241);
nand UO_1873 (O_1873,N_22706,N_24952);
nor UO_1874 (O_1874,N_23200,N_22976);
nor UO_1875 (O_1875,N_24757,N_23137);
nor UO_1876 (O_1876,N_24570,N_23688);
nand UO_1877 (O_1877,N_24077,N_24695);
and UO_1878 (O_1878,N_24041,N_24412);
and UO_1879 (O_1879,N_22719,N_23253);
or UO_1880 (O_1880,N_23055,N_23371);
or UO_1881 (O_1881,N_23052,N_23641);
nor UO_1882 (O_1882,N_24170,N_23601);
nor UO_1883 (O_1883,N_23087,N_24414);
or UO_1884 (O_1884,N_22998,N_24437);
nand UO_1885 (O_1885,N_22632,N_23637);
nand UO_1886 (O_1886,N_22889,N_24156);
and UO_1887 (O_1887,N_23890,N_23012);
nand UO_1888 (O_1888,N_24025,N_22733);
nor UO_1889 (O_1889,N_24462,N_24502);
nand UO_1890 (O_1890,N_22873,N_24363);
nand UO_1891 (O_1891,N_23360,N_23593);
nor UO_1892 (O_1892,N_23688,N_24619);
or UO_1893 (O_1893,N_22723,N_24097);
nand UO_1894 (O_1894,N_24384,N_23463);
and UO_1895 (O_1895,N_23492,N_23402);
and UO_1896 (O_1896,N_24309,N_23360);
and UO_1897 (O_1897,N_24533,N_24101);
and UO_1898 (O_1898,N_24570,N_23832);
or UO_1899 (O_1899,N_22939,N_23617);
or UO_1900 (O_1900,N_23975,N_24141);
or UO_1901 (O_1901,N_23186,N_24374);
or UO_1902 (O_1902,N_24644,N_23613);
nor UO_1903 (O_1903,N_24627,N_23544);
nand UO_1904 (O_1904,N_22875,N_22999);
and UO_1905 (O_1905,N_24528,N_23404);
or UO_1906 (O_1906,N_24549,N_24950);
nand UO_1907 (O_1907,N_24470,N_24655);
or UO_1908 (O_1908,N_24123,N_22729);
or UO_1909 (O_1909,N_22992,N_24686);
nand UO_1910 (O_1910,N_23193,N_22985);
nand UO_1911 (O_1911,N_23337,N_23291);
or UO_1912 (O_1912,N_24402,N_24161);
nor UO_1913 (O_1913,N_24574,N_24210);
and UO_1914 (O_1914,N_24798,N_23980);
and UO_1915 (O_1915,N_22642,N_23060);
nand UO_1916 (O_1916,N_23484,N_23745);
nand UO_1917 (O_1917,N_22959,N_23557);
nor UO_1918 (O_1918,N_22616,N_24033);
and UO_1919 (O_1919,N_22516,N_22812);
nor UO_1920 (O_1920,N_23745,N_24601);
and UO_1921 (O_1921,N_23419,N_24643);
and UO_1922 (O_1922,N_24901,N_23807);
or UO_1923 (O_1923,N_24571,N_24240);
or UO_1924 (O_1924,N_23517,N_24537);
nand UO_1925 (O_1925,N_23783,N_24312);
nor UO_1926 (O_1926,N_24103,N_23214);
nor UO_1927 (O_1927,N_23960,N_24787);
and UO_1928 (O_1928,N_23471,N_23410);
nor UO_1929 (O_1929,N_24872,N_23402);
nor UO_1930 (O_1930,N_24103,N_23088);
and UO_1931 (O_1931,N_23657,N_23844);
or UO_1932 (O_1932,N_23195,N_24829);
and UO_1933 (O_1933,N_24050,N_24434);
nor UO_1934 (O_1934,N_24994,N_24360);
nand UO_1935 (O_1935,N_24191,N_23074);
nor UO_1936 (O_1936,N_24346,N_22654);
nand UO_1937 (O_1937,N_23155,N_24596);
nor UO_1938 (O_1938,N_24312,N_22510);
nand UO_1939 (O_1939,N_23973,N_24339);
and UO_1940 (O_1940,N_24852,N_24380);
and UO_1941 (O_1941,N_22774,N_24325);
nand UO_1942 (O_1942,N_24453,N_24049);
and UO_1943 (O_1943,N_24817,N_23397);
nand UO_1944 (O_1944,N_23424,N_23095);
or UO_1945 (O_1945,N_24259,N_24308);
or UO_1946 (O_1946,N_24307,N_24962);
or UO_1947 (O_1947,N_24291,N_24532);
and UO_1948 (O_1948,N_24797,N_24715);
nor UO_1949 (O_1949,N_23953,N_23036);
nor UO_1950 (O_1950,N_22854,N_23777);
or UO_1951 (O_1951,N_22918,N_23453);
nand UO_1952 (O_1952,N_23582,N_23474);
nor UO_1953 (O_1953,N_22814,N_24288);
nand UO_1954 (O_1954,N_24854,N_22788);
or UO_1955 (O_1955,N_22631,N_23919);
nand UO_1956 (O_1956,N_23370,N_24084);
nor UO_1957 (O_1957,N_24738,N_22772);
nor UO_1958 (O_1958,N_23612,N_23054);
and UO_1959 (O_1959,N_24176,N_22715);
and UO_1960 (O_1960,N_24010,N_22595);
or UO_1961 (O_1961,N_23248,N_23061);
and UO_1962 (O_1962,N_22879,N_24137);
nand UO_1963 (O_1963,N_22634,N_24410);
and UO_1964 (O_1964,N_24034,N_24824);
and UO_1965 (O_1965,N_24893,N_23358);
nand UO_1966 (O_1966,N_23139,N_23273);
or UO_1967 (O_1967,N_22691,N_23817);
nor UO_1968 (O_1968,N_24954,N_22995);
nand UO_1969 (O_1969,N_23247,N_22515);
nor UO_1970 (O_1970,N_24106,N_23577);
nor UO_1971 (O_1971,N_24920,N_22634);
nor UO_1972 (O_1972,N_23789,N_22897);
and UO_1973 (O_1973,N_24344,N_23812);
and UO_1974 (O_1974,N_23434,N_23021);
nor UO_1975 (O_1975,N_24824,N_24755);
nand UO_1976 (O_1976,N_24595,N_22598);
and UO_1977 (O_1977,N_24995,N_24238);
nor UO_1978 (O_1978,N_24684,N_24968);
nand UO_1979 (O_1979,N_24766,N_22995);
nand UO_1980 (O_1980,N_24625,N_23675);
or UO_1981 (O_1981,N_24803,N_22756);
or UO_1982 (O_1982,N_24136,N_24744);
and UO_1983 (O_1983,N_23821,N_23969);
and UO_1984 (O_1984,N_23315,N_23258);
or UO_1985 (O_1985,N_23217,N_22538);
nand UO_1986 (O_1986,N_23331,N_23099);
nor UO_1987 (O_1987,N_23511,N_24178);
nor UO_1988 (O_1988,N_22965,N_23745);
nor UO_1989 (O_1989,N_24049,N_23213);
or UO_1990 (O_1990,N_24143,N_22623);
nor UO_1991 (O_1991,N_24713,N_24595);
and UO_1992 (O_1992,N_23024,N_22862);
nor UO_1993 (O_1993,N_23808,N_23034);
nand UO_1994 (O_1994,N_24217,N_23457);
and UO_1995 (O_1995,N_24621,N_23986);
nor UO_1996 (O_1996,N_24703,N_23485);
nor UO_1997 (O_1997,N_22573,N_22560);
and UO_1998 (O_1998,N_24254,N_24836);
and UO_1999 (O_1999,N_23248,N_23281);
and UO_2000 (O_2000,N_23433,N_24003);
or UO_2001 (O_2001,N_24697,N_23738);
nand UO_2002 (O_2002,N_24478,N_24949);
nand UO_2003 (O_2003,N_23175,N_23967);
or UO_2004 (O_2004,N_23228,N_22809);
nand UO_2005 (O_2005,N_24922,N_24953);
or UO_2006 (O_2006,N_23612,N_23445);
and UO_2007 (O_2007,N_23714,N_22794);
nor UO_2008 (O_2008,N_24627,N_24576);
nor UO_2009 (O_2009,N_24815,N_22625);
or UO_2010 (O_2010,N_23961,N_24488);
or UO_2011 (O_2011,N_23600,N_23078);
nand UO_2012 (O_2012,N_23245,N_23617);
nand UO_2013 (O_2013,N_23539,N_24241);
or UO_2014 (O_2014,N_23366,N_23984);
nand UO_2015 (O_2015,N_22754,N_24897);
or UO_2016 (O_2016,N_24061,N_23187);
nand UO_2017 (O_2017,N_24669,N_24129);
or UO_2018 (O_2018,N_24943,N_23549);
or UO_2019 (O_2019,N_22554,N_22798);
nand UO_2020 (O_2020,N_24201,N_24413);
and UO_2021 (O_2021,N_24262,N_23515);
nor UO_2022 (O_2022,N_24164,N_23555);
or UO_2023 (O_2023,N_24283,N_23010);
nor UO_2024 (O_2024,N_24859,N_23600);
nor UO_2025 (O_2025,N_22683,N_22977);
nand UO_2026 (O_2026,N_23234,N_24491);
nor UO_2027 (O_2027,N_24088,N_23823);
and UO_2028 (O_2028,N_22956,N_23035);
nor UO_2029 (O_2029,N_24101,N_23672);
nand UO_2030 (O_2030,N_22971,N_22605);
nor UO_2031 (O_2031,N_23037,N_23965);
or UO_2032 (O_2032,N_23770,N_24708);
nand UO_2033 (O_2033,N_24667,N_24880);
or UO_2034 (O_2034,N_22550,N_23471);
or UO_2035 (O_2035,N_23892,N_23731);
nand UO_2036 (O_2036,N_24915,N_24453);
and UO_2037 (O_2037,N_24663,N_23018);
or UO_2038 (O_2038,N_22641,N_24698);
and UO_2039 (O_2039,N_23825,N_22668);
or UO_2040 (O_2040,N_23837,N_23004);
nand UO_2041 (O_2041,N_23810,N_23477);
and UO_2042 (O_2042,N_23391,N_24199);
or UO_2043 (O_2043,N_23065,N_24526);
or UO_2044 (O_2044,N_24869,N_23119);
xnor UO_2045 (O_2045,N_23996,N_22532);
or UO_2046 (O_2046,N_23797,N_24402);
or UO_2047 (O_2047,N_23863,N_23796);
nand UO_2048 (O_2048,N_24787,N_24008);
and UO_2049 (O_2049,N_24334,N_24544);
or UO_2050 (O_2050,N_24834,N_24871);
and UO_2051 (O_2051,N_23327,N_24250);
and UO_2052 (O_2052,N_24123,N_22982);
and UO_2053 (O_2053,N_22560,N_24144);
and UO_2054 (O_2054,N_23540,N_23936);
or UO_2055 (O_2055,N_23707,N_24395);
or UO_2056 (O_2056,N_23569,N_23596);
nand UO_2057 (O_2057,N_23352,N_24133);
and UO_2058 (O_2058,N_23703,N_23658);
nand UO_2059 (O_2059,N_22939,N_24358);
or UO_2060 (O_2060,N_23696,N_23381);
and UO_2061 (O_2061,N_24058,N_22739);
nor UO_2062 (O_2062,N_24430,N_23810);
and UO_2063 (O_2063,N_23605,N_24248);
or UO_2064 (O_2064,N_24208,N_23101);
or UO_2065 (O_2065,N_24655,N_23556);
nand UO_2066 (O_2066,N_22599,N_22965);
nor UO_2067 (O_2067,N_24281,N_23406);
and UO_2068 (O_2068,N_24380,N_24808);
nor UO_2069 (O_2069,N_22526,N_24452);
and UO_2070 (O_2070,N_23118,N_22651);
or UO_2071 (O_2071,N_24962,N_23672);
nor UO_2072 (O_2072,N_23867,N_22550);
or UO_2073 (O_2073,N_23074,N_23979);
and UO_2074 (O_2074,N_24700,N_24681);
or UO_2075 (O_2075,N_24981,N_24944);
and UO_2076 (O_2076,N_22587,N_22719);
nor UO_2077 (O_2077,N_23481,N_22555);
nand UO_2078 (O_2078,N_23237,N_22592);
and UO_2079 (O_2079,N_23813,N_24890);
or UO_2080 (O_2080,N_22805,N_23363);
or UO_2081 (O_2081,N_24719,N_24864);
and UO_2082 (O_2082,N_22776,N_23176);
nor UO_2083 (O_2083,N_23650,N_24570);
nor UO_2084 (O_2084,N_22924,N_23830);
or UO_2085 (O_2085,N_24593,N_24741);
or UO_2086 (O_2086,N_23684,N_22905);
nand UO_2087 (O_2087,N_23477,N_23069);
and UO_2088 (O_2088,N_23244,N_23883);
and UO_2089 (O_2089,N_24382,N_24397);
and UO_2090 (O_2090,N_23711,N_24592);
or UO_2091 (O_2091,N_23005,N_23903);
nand UO_2092 (O_2092,N_22582,N_22737);
or UO_2093 (O_2093,N_22729,N_24575);
or UO_2094 (O_2094,N_23622,N_24978);
nor UO_2095 (O_2095,N_22905,N_24645);
or UO_2096 (O_2096,N_24687,N_23630);
or UO_2097 (O_2097,N_22522,N_23889);
or UO_2098 (O_2098,N_23829,N_24625);
nor UO_2099 (O_2099,N_24987,N_23789);
and UO_2100 (O_2100,N_24289,N_24498);
nor UO_2101 (O_2101,N_23763,N_23911);
and UO_2102 (O_2102,N_24070,N_24736);
nand UO_2103 (O_2103,N_23534,N_24571);
and UO_2104 (O_2104,N_24422,N_24608);
nor UO_2105 (O_2105,N_24871,N_23253);
nand UO_2106 (O_2106,N_22996,N_23877);
nand UO_2107 (O_2107,N_23179,N_24898);
and UO_2108 (O_2108,N_24861,N_24015);
or UO_2109 (O_2109,N_22563,N_23369);
or UO_2110 (O_2110,N_23566,N_23769);
and UO_2111 (O_2111,N_23111,N_24763);
nand UO_2112 (O_2112,N_23304,N_23273);
nand UO_2113 (O_2113,N_23523,N_23055);
nand UO_2114 (O_2114,N_24195,N_23622);
nand UO_2115 (O_2115,N_23795,N_22566);
nand UO_2116 (O_2116,N_23213,N_23024);
and UO_2117 (O_2117,N_23055,N_22655);
nor UO_2118 (O_2118,N_23220,N_23690);
and UO_2119 (O_2119,N_23105,N_22638);
and UO_2120 (O_2120,N_24554,N_22581);
nor UO_2121 (O_2121,N_23669,N_24397);
and UO_2122 (O_2122,N_23784,N_23466);
nor UO_2123 (O_2123,N_24636,N_24256);
nand UO_2124 (O_2124,N_23398,N_23970);
or UO_2125 (O_2125,N_24577,N_24735);
nand UO_2126 (O_2126,N_23623,N_23317);
nand UO_2127 (O_2127,N_23976,N_23230);
and UO_2128 (O_2128,N_23321,N_24801);
nor UO_2129 (O_2129,N_23615,N_23321);
nor UO_2130 (O_2130,N_24757,N_22629);
and UO_2131 (O_2131,N_24049,N_23710);
nor UO_2132 (O_2132,N_24040,N_22689);
nor UO_2133 (O_2133,N_24128,N_23427);
nor UO_2134 (O_2134,N_22646,N_24843);
and UO_2135 (O_2135,N_23246,N_23067);
xor UO_2136 (O_2136,N_23687,N_24731);
or UO_2137 (O_2137,N_23980,N_22608);
or UO_2138 (O_2138,N_24369,N_22668);
and UO_2139 (O_2139,N_23872,N_24337);
and UO_2140 (O_2140,N_24233,N_22946);
nor UO_2141 (O_2141,N_23189,N_23804);
nor UO_2142 (O_2142,N_24757,N_22795);
nor UO_2143 (O_2143,N_22676,N_24129);
and UO_2144 (O_2144,N_22551,N_24962);
and UO_2145 (O_2145,N_22857,N_23777);
nand UO_2146 (O_2146,N_24028,N_24625);
nand UO_2147 (O_2147,N_24938,N_23230);
and UO_2148 (O_2148,N_24266,N_24976);
or UO_2149 (O_2149,N_24053,N_23597);
nand UO_2150 (O_2150,N_24257,N_22816);
nand UO_2151 (O_2151,N_23368,N_24681);
and UO_2152 (O_2152,N_23836,N_24988);
and UO_2153 (O_2153,N_24680,N_23428);
or UO_2154 (O_2154,N_23799,N_23348);
nor UO_2155 (O_2155,N_23127,N_22995);
nor UO_2156 (O_2156,N_23609,N_24983);
or UO_2157 (O_2157,N_24917,N_23344);
and UO_2158 (O_2158,N_22884,N_23871);
nand UO_2159 (O_2159,N_24135,N_24065);
and UO_2160 (O_2160,N_22623,N_23307);
and UO_2161 (O_2161,N_24432,N_23322);
and UO_2162 (O_2162,N_22807,N_22669);
nand UO_2163 (O_2163,N_23953,N_24807);
nor UO_2164 (O_2164,N_23556,N_23979);
nand UO_2165 (O_2165,N_23719,N_24146);
nor UO_2166 (O_2166,N_22574,N_23806);
and UO_2167 (O_2167,N_23044,N_23334);
nor UO_2168 (O_2168,N_24898,N_23437);
or UO_2169 (O_2169,N_24930,N_23967);
nor UO_2170 (O_2170,N_23928,N_24206);
nand UO_2171 (O_2171,N_23827,N_24700);
or UO_2172 (O_2172,N_24593,N_22843);
or UO_2173 (O_2173,N_23204,N_22989);
and UO_2174 (O_2174,N_24027,N_24717);
and UO_2175 (O_2175,N_23980,N_22784);
nor UO_2176 (O_2176,N_24261,N_24465);
and UO_2177 (O_2177,N_22633,N_23650);
and UO_2178 (O_2178,N_24535,N_23613);
nand UO_2179 (O_2179,N_23258,N_22615);
and UO_2180 (O_2180,N_24353,N_22537);
nor UO_2181 (O_2181,N_24406,N_22857);
and UO_2182 (O_2182,N_23217,N_23657);
or UO_2183 (O_2183,N_23652,N_24003);
or UO_2184 (O_2184,N_23642,N_24478);
nand UO_2185 (O_2185,N_24977,N_23785);
nand UO_2186 (O_2186,N_24660,N_23334);
and UO_2187 (O_2187,N_24415,N_23920);
or UO_2188 (O_2188,N_24417,N_23984);
and UO_2189 (O_2189,N_23349,N_22729);
xnor UO_2190 (O_2190,N_24431,N_23501);
nor UO_2191 (O_2191,N_24667,N_24994);
and UO_2192 (O_2192,N_23098,N_24308);
or UO_2193 (O_2193,N_23033,N_24922);
or UO_2194 (O_2194,N_24900,N_22638);
or UO_2195 (O_2195,N_22789,N_23772);
and UO_2196 (O_2196,N_24020,N_23164);
nor UO_2197 (O_2197,N_24624,N_23677);
or UO_2198 (O_2198,N_22677,N_24813);
nor UO_2199 (O_2199,N_23230,N_24770);
or UO_2200 (O_2200,N_24832,N_23186);
and UO_2201 (O_2201,N_24314,N_23787);
xnor UO_2202 (O_2202,N_23565,N_22512);
nor UO_2203 (O_2203,N_24746,N_22599);
nor UO_2204 (O_2204,N_23850,N_22555);
and UO_2205 (O_2205,N_23961,N_23074);
nand UO_2206 (O_2206,N_24255,N_23655);
or UO_2207 (O_2207,N_23375,N_22663);
or UO_2208 (O_2208,N_22830,N_24199);
nor UO_2209 (O_2209,N_22745,N_24805);
nand UO_2210 (O_2210,N_24044,N_23997);
nand UO_2211 (O_2211,N_24339,N_23522);
or UO_2212 (O_2212,N_24366,N_24071);
or UO_2213 (O_2213,N_24809,N_24461);
nor UO_2214 (O_2214,N_22925,N_22737);
or UO_2215 (O_2215,N_24667,N_24731);
or UO_2216 (O_2216,N_24596,N_23999);
nand UO_2217 (O_2217,N_23284,N_23990);
nor UO_2218 (O_2218,N_22970,N_24107);
or UO_2219 (O_2219,N_23539,N_22763);
nor UO_2220 (O_2220,N_24584,N_22968);
or UO_2221 (O_2221,N_23533,N_24669);
and UO_2222 (O_2222,N_24910,N_23006);
nor UO_2223 (O_2223,N_22530,N_24466);
nor UO_2224 (O_2224,N_22964,N_23018);
and UO_2225 (O_2225,N_22902,N_22523);
nor UO_2226 (O_2226,N_23652,N_23524);
nor UO_2227 (O_2227,N_23320,N_24160);
and UO_2228 (O_2228,N_22702,N_23583);
and UO_2229 (O_2229,N_23249,N_23919);
nor UO_2230 (O_2230,N_22812,N_23653);
nor UO_2231 (O_2231,N_23444,N_23061);
nor UO_2232 (O_2232,N_24676,N_23469);
nand UO_2233 (O_2233,N_22564,N_23596);
or UO_2234 (O_2234,N_23121,N_24618);
nand UO_2235 (O_2235,N_23194,N_23850);
or UO_2236 (O_2236,N_23749,N_23560);
nand UO_2237 (O_2237,N_22583,N_22516);
nor UO_2238 (O_2238,N_24216,N_24475);
and UO_2239 (O_2239,N_24870,N_22955);
and UO_2240 (O_2240,N_23756,N_24978);
nand UO_2241 (O_2241,N_24279,N_22671);
nor UO_2242 (O_2242,N_23626,N_22636);
and UO_2243 (O_2243,N_23584,N_23706);
and UO_2244 (O_2244,N_24452,N_23819);
nand UO_2245 (O_2245,N_24631,N_24718);
or UO_2246 (O_2246,N_22531,N_24208);
nand UO_2247 (O_2247,N_23485,N_22843);
nand UO_2248 (O_2248,N_22741,N_23645);
nand UO_2249 (O_2249,N_22881,N_24182);
nand UO_2250 (O_2250,N_24906,N_24515);
or UO_2251 (O_2251,N_23600,N_23513);
or UO_2252 (O_2252,N_23677,N_24615);
and UO_2253 (O_2253,N_23737,N_23649);
and UO_2254 (O_2254,N_23671,N_23350);
nor UO_2255 (O_2255,N_23023,N_22876);
nand UO_2256 (O_2256,N_24498,N_23569);
or UO_2257 (O_2257,N_22642,N_22673);
or UO_2258 (O_2258,N_23182,N_23144);
and UO_2259 (O_2259,N_23340,N_22574);
or UO_2260 (O_2260,N_23041,N_23264);
nand UO_2261 (O_2261,N_23645,N_23012);
and UO_2262 (O_2262,N_24627,N_23189);
nor UO_2263 (O_2263,N_23494,N_23399);
nand UO_2264 (O_2264,N_24478,N_22783);
nor UO_2265 (O_2265,N_24975,N_24461);
or UO_2266 (O_2266,N_23677,N_24208);
and UO_2267 (O_2267,N_24085,N_23364);
nand UO_2268 (O_2268,N_22543,N_24907);
or UO_2269 (O_2269,N_24501,N_24504);
nor UO_2270 (O_2270,N_23820,N_23938);
xor UO_2271 (O_2271,N_24547,N_24514);
and UO_2272 (O_2272,N_24942,N_23832);
or UO_2273 (O_2273,N_23700,N_23883);
and UO_2274 (O_2274,N_24873,N_22734);
and UO_2275 (O_2275,N_23146,N_22818);
or UO_2276 (O_2276,N_22986,N_22665);
nor UO_2277 (O_2277,N_23083,N_24685);
nand UO_2278 (O_2278,N_23869,N_24383);
nor UO_2279 (O_2279,N_23098,N_22813);
nand UO_2280 (O_2280,N_24898,N_24470);
or UO_2281 (O_2281,N_23598,N_22840);
nor UO_2282 (O_2282,N_24020,N_23514);
or UO_2283 (O_2283,N_23659,N_23430);
and UO_2284 (O_2284,N_22576,N_23356);
or UO_2285 (O_2285,N_23071,N_23425);
nor UO_2286 (O_2286,N_23240,N_23122);
and UO_2287 (O_2287,N_24177,N_24434);
nand UO_2288 (O_2288,N_23205,N_22798);
or UO_2289 (O_2289,N_24529,N_24914);
nand UO_2290 (O_2290,N_23208,N_22770);
nor UO_2291 (O_2291,N_22779,N_23251);
or UO_2292 (O_2292,N_22925,N_22538);
xnor UO_2293 (O_2293,N_23938,N_24458);
and UO_2294 (O_2294,N_24487,N_24593);
and UO_2295 (O_2295,N_23057,N_24007);
and UO_2296 (O_2296,N_23512,N_22857);
nand UO_2297 (O_2297,N_22661,N_23859);
or UO_2298 (O_2298,N_24145,N_23479);
or UO_2299 (O_2299,N_24324,N_22855);
nor UO_2300 (O_2300,N_23337,N_24025);
nor UO_2301 (O_2301,N_22660,N_24712);
or UO_2302 (O_2302,N_22916,N_23359);
nand UO_2303 (O_2303,N_24583,N_22989);
nor UO_2304 (O_2304,N_24402,N_24762);
nand UO_2305 (O_2305,N_24579,N_23146);
or UO_2306 (O_2306,N_22624,N_22752);
nor UO_2307 (O_2307,N_23589,N_23894);
or UO_2308 (O_2308,N_24908,N_24328);
nor UO_2309 (O_2309,N_23912,N_23518);
nor UO_2310 (O_2310,N_23916,N_23960);
nor UO_2311 (O_2311,N_22954,N_24362);
nor UO_2312 (O_2312,N_22989,N_24577);
or UO_2313 (O_2313,N_23526,N_23122);
or UO_2314 (O_2314,N_24247,N_22949);
or UO_2315 (O_2315,N_24152,N_23422);
or UO_2316 (O_2316,N_23553,N_24837);
or UO_2317 (O_2317,N_24883,N_23465);
and UO_2318 (O_2318,N_24142,N_22502);
or UO_2319 (O_2319,N_22531,N_24301);
nor UO_2320 (O_2320,N_23743,N_24882);
nor UO_2321 (O_2321,N_23798,N_24831);
nor UO_2322 (O_2322,N_22609,N_24908);
or UO_2323 (O_2323,N_24127,N_24212);
and UO_2324 (O_2324,N_24103,N_23199);
or UO_2325 (O_2325,N_22809,N_22702);
and UO_2326 (O_2326,N_24367,N_23284);
and UO_2327 (O_2327,N_23898,N_23287);
or UO_2328 (O_2328,N_24551,N_22869);
and UO_2329 (O_2329,N_23853,N_24685);
xor UO_2330 (O_2330,N_22876,N_22827);
and UO_2331 (O_2331,N_23918,N_22522);
and UO_2332 (O_2332,N_24262,N_23183);
nor UO_2333 (O_2333,N_22801,N_23801);
nand UO_2334 (O_2334,N_24777,N_24615);
nand UO_2335 (O_2335,N_23194,N_23131);
or UO_2336 (O_2336,N_22667,N_24579);
or UO_2337 (O_2337,N_24904,N_23029);
or UO_2338 (O_2338,N_23309,N_24815);
nand UO_2339 (O_2339,N_24188,N_24134);
nor UO_2340 (O_2340,N_24351,N_22996);
nand UO_2341 (O_2341,N_24488,N_24920);
and UO_2342 (O_2342,N_24838,N_24005);
nor UO_2343 (O_2343,N_22959,N_23352);
nand UO_2344 (O_2344,N_23293,N_23279);
nor UO_2345 (O_2345,N_24090,N_24006);
nand UO_2346 (O_2346,N_23707,N_22699);
nor UO_2347 (O_2347,N_23833,N_22659);
nand UO_2348 (O_2348,N_23986,N_23713);
nand UO_2349 (O_2349,N_23682,N_24666);
or UO_2350 (O_2350,N_24778,N_24497);
nand UO_2351 (O_2351,N_24543,N_23486);
and UO_2352 (O_2352,N_23407,N_22890);
and UO_2353 (O_2353,N_24332,N_23607);
nor UO_2354 (O_2354,N_24532,N_23193);
and UO_2355 (O_2355,N_23707,N_23856);
nand UO_2356 (O_2356,N_23224,N_23186);
and UO_2357 (O_2357,N_23545,N_22946);
nor UO_2358 (O_2358,N_22885,N_22755);
nand UO_2359 (O_2359,N_23893,N_22658);
nand UO_2360 (O_2360,N_22777,N_23180);
or UO_2361 (O_2361,N_23971,N_22977);
nand UO_2362 (O_2362,N_22836,N_23356);
nand UO_2363 (O_2363,N_23376,N_24341);
or UO_2364 (O_2364,N_24988,N_24759);
nor UO_2365 (O_2365,N_24627,N_23661);
and UO_2366 (O_2366,N_23921,N_24243);
nor UO_2367 (O_2367,N_23229,N_22745);
nor UO_2368 (O_2368,N_24739,N_23953);
and UO_2369 (O_2369,N_24247,N_23240);
or UO_2370 (O_2370,N_23456,N_24463);
nand UO_2371 (O_2371,N_22807,N_23061);
nand UO_2372 (O_2372,N_23565,N_22905);
or UO_2373 (O_2373,N_22695,N_24988);
and UO_2374 (O_2374,N_23169,N_22524);
or UO_2375 (O_2375,N_24205,N_24043);
and UO_2376 (O_2376,N_24278,N_22673);
nor UO_2377 (O_2377,N_23828,N_24550);
or UO_2378 (O_2378,N_24470,N_24322);
or UO_2379 (O_2379,N_23076,N_24264);
or UO_2380 (O_2380,N_23581,N_24965);
nand UO_2381 (O_2381,N_23212,N_22592);
nor UO_2382 (O_2382,N_23929,N_24660);
and UO_2383 (O_2383,N_22500,N_23427);
nor UO_2384 (O_2384,N_24218,N_24772);
nand UO_2385 (O_2385,N_24501,N_24481);
and UO_2386 (O_2386,N_24982,N_24092);
nor UO_2387 (O_2387,N_23550,N_22721);
and UO_2388 (O_2388,N_22652,N_22993);
nand UO_2389 (O_2389,N_22688,N_24236);
nand UO_2390 (O_2390,N_22584,N_23384);
nand UO_2391 (O_2391,N_24095,N_22672);
nand UO_2392 (O_2392,N_23204,N_23902);
or UO_2393 (O_2393,N_24754,N_22988);
nand UO_2394 (O_2394,N_22922,N_23720);
nor UO_2395 (O_2395,N_24433,N_24089);
nor UO_2396 (O_2396,N_23619,N_23256);
or UO_2397 (O_2397,N_23652,N_23106);
or UO_2398 (O_2398,N_23011,N_22825);
and UO_2399 (O_2399,N_22643,N_23313);
xor UO_2400 (O_2400,N_24534,N_23336);
nand UO_2401 (O_2401,N_23759,N_23513);
or UO_2402 (O_2402,N_24230,N_23918);
nor UO_2403 (O_2403,N_24676,N_24668);
nand UO_2404 (O_2404,N_22994,N_24257);
or UO_2405 (O_2405,N_23917,N_22632);
and UO_2406 (O_2406,N_23837,N_22786);
nor UO_2407 (O_2407,N_24953,N_22860);
or UO_2408 (O_2408,N_23395,N_22656);
or UO_2409 (O_2409,N_23743,N_23505);
nand UO_2410 (O_2410,N_22792,N_23906);
nand UO_2411 (O_2411,N_23312,N_24087);
nand UO_2412 (O_2412,N_23201,N_23865);
and UO_2413 (O_2413,N_24992,N_23470);
or UO_2414 (O_2414,N_23943,N_24619);
nand UO_2415 (O_2415,N_24882,N_23394);
or UO_2416 (O_2416,N_24332,N_24950);
or UO_2417 (O_2417,N_24231,N_24004);
nor UO_2418 (O_2418,N_22929,N_24285);
nand UO_2419 (O_2419,N_22771,N_24531);
nor UO_2420 (O_2420,N_22537,N_24974);
or UO_2421 (O_2421,N_23077,N_23274);
and UO_2422 (O_2422,N_23209,N_22803);
nand UO_2423 (O_2423,N_24319,N_23123);
or UO_2424 (O_2424,N_24046,N_23847);
or UO_2425 (O_2425,N_23961,N_23982);
and UO_2426 (O_2426,N_24112,N_22769);
nor UO_2427 (O_2427,N_24149,N_23229);
or UO_2428 (O_2428,N_23984,N_24271);
nor UO_2429 (O_2429,N_23714,N_24247);
nand UO_2430 (O_2430,N_23339,N_23378);
nor UO_2431 (O_2431,N_23786,N_23153);
or UO_2432 (O_2432,N_22869,N_22980);
and UO_2433 (O_2433,N_23507,N_24640);
nor UO_2434 (O_2434,N_24349,N_23528);
nor UO_2435 (O_2435,N_23009,N_24397);
nor UO_2436 (O_2436,N_24388,N_22543);
or UO_2437 (O_2437,N_24982,N_23212);
or UO_2438 (O_2438,N_24295,N_24191);
or UO_2439 (O_2439,N_24409,N_22511);
and UO_2440 (O_2440,N_24790,N_23790);
and UO_2441 (O_2441,N_23866,N_23617);
nor UO_2442 (O_2442,N_24050,N_22894);
nand UO_2443 (O_2443,N_23726,N_24910);
nand UO_2444 (O_2444,N_23465,N_24462);
nand UO_2445 (O_2445,N_24090,N_23834);
or UO_2446 (O_2446,N_24993,N_23849);
and UO_2447 (O_2447,N_24050,N_24960);
or UO_2448 (O_2448,N_23075,N_23336);
nand UO_2449 (O_2449,N_23839,N_22587);
nor UO_2450 (O_2450,N_24054,N_23367);
nand UO_2451 (O_2451,N_23661,N_22643);
and UO_2452 (O_2452,N_24871,N_24860);
or UO_2453 (O_2453,N_23687,N_23854);
nor UO_2454 (O_2454,N_24673,N_24565);
and UO_2455 (O_2455,N_23165,N_23155);
nand UO_2456 (O_2456,N_23107,N_23337);
and UO_2457 (O_2457,N_24338,N_22742);
and UO_2458 (O_2458,N_24697,N_23513);
or UO_2459 (O_2459,N_22751,N_23862);
nand UO_2460 (O_2460,N_24351,N_24916);
nand UO_2461 (O_2461,N_24134,N_23481);
nand UO_2462 (O_2462,N_23345,N_23010);
nor UO_2463 (O_2463,N_22862,N_23612);
and UO_2464 (O_2464,N_24635,N_24172);
nor UO_2465 (O_2465,N_23341,N_24083);
nand UO_2466 (O_2466,N_23515,N_24701);
and UO_2467 (O_2467,N_22521,N_22620);
and UO_2468 (O_2468,N_23656,N_24648);
and UO_2469 (O_2469,N_24973,N_24584);
and UO_2470 (O_2470,N_24162,N_23537);
or UO_2471 (O_2471,N_23380,N_22992);
or UO_2472 (O_2472,N_24108,N_23046);
or UO_2473 (O_2473,N_24167,N_23142);
nor UO_2474 (O_2474,N_23041,N_22513);
nand UO_2475 (O_2475,N_24247,N_22682);
nor UO_2476 (O_2476,N_23594,N_24836);
and UO_2477 (O_2477,N_23085,N_22618);
nor UO_2478 (O_2478,N_24139,N_23240);
nor UO_2479 (O_2479,N_23730,N_23223);
and UO_2480 (O_2480,N_24915,N_23604);
and UO_2481 (O_2481,N_22525,N_23225);
or UO_2482 (O_2482,N_23852,N_23890);
xor UO_2483 (O_2483,N_24494,N_24809);
nand UO_2484 (O_2484,N_24207,N_22931);
or UO_2485 (O_2485,N_23033,N_24914);
and UO_2486 (O_2486,N_24228,N_23373);
nand UO_2487 (O_2487,N_24485,N_23246);
nand UO_2488 (O_2488,N_24352,N_24107);
nand UO_2489 (O_2489,N_24956,N_23004);
nand UO_2490 (O_2490,N_24126,N_23836);
nor UO_2491 (O_2491,N_24882,N_22763);
or UO_2492 (O_2492,N_23972,N_23392);
and UO_2493 (O_2493,N_24043,N_24237);
nor UO_2494 (O_2494,N_24504,N_22548);
and UO_2495 (O_2495,N_23288,N_22527);
or UO_2496 (O_2496,N_23284,N_24374);
and UO_2497 (O_2497,N_23793,N_23983);
and UO_2498 (O_2498,N_24888,N_23169);
nor UO_2499 (O_2499,N_24828,N_23879);
or UO_2500 (O_2500,N_23892,N_24980);
nand UO_2501 (O_2501,N_23652,N_23374);
or UO_2502 (O_2502,N_23087,N_24618);
nor UO_2503 (O_2503,N_23299,N_24806);
or UO_2504 (O_2504,N_24768,N_22808);
and UO_2505 (O_2505,N_23537,N_24398);
and UO_2506 (O_2506,N_23506,N_23562);
nand UO_2507 (O_2507,N_24369,N_23082);
or UO_2508 (O_2508,N_23477,N_22951);
or UO_2509 (O_2509,N_23155,N_24065);
and UO_2510 (O_2510,N_24905,N_23732);
or UO_2511 (O_2511,N_22541,N_24001);
nor UO_2512 (O_2512,N_23782,N_24219);
or UO_2513 (O_2513,N_24674,N_23965);
and UO_2514 (O_2514,N_23733,N_23678);
nand UO_2515 (O_2515,N_24869,N_22882);
and UO_2516 (O_2516,N_23746,N_22971);
or UO_2517 (O_2517,N_24426,N_23900);
and UO_2518 (O_2518,N_24542,N_23416);
nor UO_2519 (O_2519,N_24053,N_24388);
or UO_2520 (O_2520,N_23538,N_23342);
nor UO_2521 (O_2521,N_23295,N_23823);
nand UO_2522 (O_2522,N_24470,N_22549);
and UO_2523 (O_2523,N_24981,N_24200);
nor UO_2524 (O_2524,N_24288,N_24294);
nand UO_2525 (O_2525,N_24630,N_23352);
or UO_2526 (O_2526,N_23270,N_23291);
or UO_2527 (O_2527,N_23692,N_24911);
or UO_2528 (O_2528,N_23892,N_24609);
nand UO_2529 (O_2529,N_24486,N_24007);
nor UO_2530 (O_2530,N_23893,N_23408);
or UO_2531 (O_2531,N_23263,N_23349);
nand UO_2532 (O_2532,N_23395,N_23496);
nor UO_2533 (O_2533,N_24353,N_22667);
nor UO_2534 (O_2534,N_23179,N_24868);
or UO_2535 (O_2535,N_23582,N_22870);
nand UO_2536 (O_2536,N_22811,N_24679);
nand UO_2537 (O_2537,N_24685,N_24695);
nand UO_2538 (O_2538,N_23780,N_24639);
and UO_2539 (O_2539,N_23417,N_23178);
xor UO_2540 (O_2540,N_23105,N_22848);
nand UO_2541 (O_2541,N_24262,N_23219);
and UO_2542 (O_2542,N_24631,N_23454);
nor UO_2543 (O_2543,N_22541,N_22858);
nand UO_2544 (O_2544,N_23981,N_23926);
nor UO_2545 (O_2545,N_24552,N_24121);
and UO_2546 (O_2546,N_22626,N_23375);
nand UO_2547 (O_2547,N_24203,N_24555);
nor UO_2548 (O_2548,N_23431,N_23898);
or UO_2549 (O_2549,N_23641,N_24024);
or UO_2550 (O_2550,N_24181,N_22819);
or UO_2551 (O_2551,N_22673,N_24415);
or UO_2552 (O_2552,N_22851,N_24614);
and UO_2553 (O_2553,N_23888,N_23734);
or UO_2554 (O_2554,N_22531,N_22673);
or UO_2555 (O_2555,N_22846,N_24097);
nor UO_2556 (O_2556,N_23037,N_23260);
nand UO_2557 (O_2557,N_24099,N_24648);
and UO_2558 (O_2558,N_24177,N_24697);
nor UO_2559 (O_2559,N_22863,N_24254);
nand UO_2560 (O_2560,N_23733,N_24278);
nor UO_2561 (O_2561,N_23587,N_24841);
nor UO_2562 (O_2562,N_23518,N_24423);
nor UO_2563 (O_2563,N_24586,N_24930);
or UO_2564 (O_2564,N_22569,N_24319);
nand UO_2565 (O_2565,N_24045,N_22611);
nor UO_2566 (O_2566,N_24181,N_23295);
or UO_2567 (O_2567,N_24066,N_22676);
nor UO_2568 (O_2568,N_22592,N_24875);
and UO_2569 (O_2569,N_23932,N_23426);
or UO_2570 (O_2570,N_23856,N_23738);
nand UO_2571 (O_2571,N_22698,N_24771);
and UO_2572 (O_2572,N_23520,N_22604);
or UO_2573 (O_2573,N_24492,N_24991);
nand UO_2574 (O_2574,N_23087,N_24823);
xnor UO_2575 (O_2575,N_24553,N_22759);
or UO_2576 (O_2576,N_22863,N_24816);
or UO_2577 (O_2577,N_23815,N_24424);
or UO_2578 (O_2578,N_23615,N_24374);
nor UO_2579 (O_2579,N_23951,N_23636);
and UO_2580 (O_2580,N_22640,N_24669);
and UO_2581 (O_2581,N_24204,N_23029);
or UO_2582 (O_2582,N_22721,N_22852);
nor UO_2583 (O_2583,N_22542,N_23513);
and UO_2584 (O_2584,N_24903,N_22650);
or UO_2585 (O_2585,N_23388,N_23747);
nor UO_2586 (O_2586,N_22568,N_22654);
or UO_2587 (O_2587,N_24235,N_22657);
and UO_2588 (O_2588,N_22573,N_22887);
or UO_2589 (O_2589,N_24181,N_23058);
nand UO_2590 (O_2590,N_22554,N_22527);
nand UO_2591 (O_2591,N_22982,N_22508);
nand UO_2592 (O_2592,N_23569,N_24479);
nand UO_2593 (O_2593,N_23514,N_23948);
nand UO_2594 (O_2594,N_23236,N_23148);
and UO_2595 (O_2595,N_23908,N_24906);
or UO_2596 (O_2596,N_23710,N_24053);
nor UO_2597 (O_2597,N_24878,N_24582);
nand UO_2598 (O_2598,N_23089,N_24067);
or UO_2599 (O_2599,N_23989,N_24178);
nor UO_2600 (O_2600,N_24184,N_23111);
or UO_2601 (O_2601,N_23856,N_24899);
nor UO_2602 (O_2602,N_24079,N_24863);
nor UO_2603 (O_2603,N_23438,N_22965);
nand UO_2604 (O_2604,N_23155,N_22688);
nand UO_2605 (O_2605,N_24675,N_23528);
or UO_2606 (O_2606,N_22713,N_23455);
and UO_2607 (O_2607,N_23981,N_23769);
or UO_2608 (O_2608,N_24736,N_24063);
nand UO_2609 (O_2609,N_24801,N_24048);
nor UO_2610 (O_2610,N_24544,N_24818);
nor UO_2611 (O_2611,N_23832,N_23522);
nor UO_2612 (O_2612,N_22971,N_23556);
or UO_2613 (O_2613,N_23487,N_24931);
or UO_2614 (O_2614,N_24584,N_23337);
or UO_2615 (O_2615,N_23649,N_24798);
nor UO_2616 (O_2616,N_24199,N_24234);
xor UO_2617 (O_2617,N_23077,N_24728);
and UO_2618 (O_2618,N_24158,N_24842);
nor UO_2619 (O_2619,N_24694,N_24713);
nor UO_2620 (O_2620,N_24572,N_23327);
nand UO_2621 (O_2621,N_23054,N_23977);
and UO_2622 (O_2622,N_23912,N_24243);
nand UO_2623 (O_2623,N_22816,N_23195);
nand UO_2624 (O_2624,N_23472,N_23677);
nor UO_2625 (O_2625,N_23678,N_23955);
nand UO_2626 (O_2626,N_24827,N_23483);
or UO_2627 (O_2627,N_24895,N_24702);
nor UO_2628 (O_2628,N_23604,N_23822);
nand UO_2629 (O_2629,N_23767,N_22804);
and UO_2630 (O_2630,N_22589,N_23879);
nor UO_2631 (O_2631,N_24443,N_23833);
xor UO_2632 (O_2632,N_23542,N_23684);
nor UO_2633 (O_2633,N_24980,N_24154);
or UO_2634 (O_2634,N_22698,N_22990);
nor UO_2635 (O_2635,N_24002,N_22986);
and UO_2636 (O_2636,N_23433,N_23477);
and UO_2637 (O_2637,N_23518,N_24920);
xnor UO_2638 (O_2638,N_22994,N_22781);
nand UO_2639 (O_2639,N_24332,N_22612);
or UO_2640 (O_2640,N_24595,N_23741);
nand UO_2641 (O_2641,N_23680,N_22805);
xor UO_2642 (O_2642,N_24572,N_24290);
nand UO_2643 (O_2643,N_22999,N_23391);
nand UO_2644 (O_2644,N_23787,N_22949);
and UO_2645 (O_2645,N_23011,N_22953);
nor UO_2646 (O_2646,N_23510,N_24258);
xnor UO_2647 (O_2647,N_24294,N_23902);
or UO_2648 (O_2648,N_23423,N_22727);
or UO_2649 (O_2649,N_24577,N_23011);
nor UO_2650 (O_2650,N_24561,N_23198);
nand UO_2651 (O_2651,N_23611,N_24522);
nor UO_2652 (O_2652,N_23849,N_23060);
nand UO_2653 (O_2653,N_24613,N_24546);
or UO_2654 (O_2654,N_24772,N_23250);
and UO_2655 (O_2655,N_24484,N_24283);
and UO_2656 (O_2656,N_23297,N_23317);
or UO_2657 (O_2657,N_23563,N_23342);
nand UO_2658 (O_2658,N_23682,N_23193);
or UO_2659 (O_2659,N_23326,N_23854);
nand UO_2660 (O_2660,N_23171,N_24920);
or UO_2661 (O_2661,N_22511,N_24560);
nor UO_2662 (O_2662,N_24373,N_24959);
and UO_2663 (O_2663,N_24154,N_23948);
nor UO_2664 (O_2664,N_24855,N_23919);
nor UO_2665 (O_2665,N_24234,N_23012);
nor UO_2666 (O_2666,N_23277,N_24763);
or UO_2667 (O_2667,N_24412,N_24078);
nor UO_2668 (O_2668,N_23682,N_24839);
or UO_2669 (O_2669,N_23000,N_23960);
nor UO_2670 (O_2670,N_24213,N_23061);
nand UO_2671 (O_2671,N_23490,N_24739);
xnor UO_2672 (O_2672,N_24785,N_23145);
or UO_2673 (O_2673,N_23129,N_24191);
nor UO_2674 (O_2674,N_22823,N_24526);
and UO_2675 (O_2675,N_24681,N_24383);
or UO_2676 (O_2676,N_24570,N_22717);
nand UO_2677 (O_2677,N_23167,N_23538);
or UO_2678 (O_2678,N_24980,N_22956);
nor UO_2679 (O_2679,N_22616,N_23001);
or UO_2680 (O_2680,N_24803,N_23047);
nor UO_2681 (O_2681,N_24616,N_23338);
or UO_2682 (O_2682,N_23966,N_24401);
nand UO_2683 (O_2683,N_23712,N_24648);
nor UO_2684 (O_2684,N_24093,N_24920);
or UO_2685 (O_2685,N_22741,N_23814);
nand UO_2686 (O_2686,N_23072,N_24042);
and UO_2687 (O_2687,N_23342,N_23046);
nor UO_2688 (O_2688,N_24108,N_24550);
nor UO_2689 (O_2689,N_22548,N_22689);
or UO_2690 (O_2690,N_24866,N_22934);
and UO_2691 (O_2691,N_23685,N_24279);
and UO_2692 (O_2692,N_24132,N_24385);
nand UO_2693 (O_2693,N_23564,N_24103);
and UO_2694 (O_2694,N_23801,N_23029);
nand UO_2695 (O_2695,N_24655,N_24838);
nor UO_2696 (O_2696,N_23717,N_24028);
or UO_2697 (O_2697,N_24225,N_24118);
nand UO_2698 (O_2698,N_24806,N_24138);
nand UO_2699 (O_2699,N_22680,N_24369);
nand UO_2700 (O_2700,N_24275,N_23469);
nand UO_2701 (O_2701,N_22876,N_22602);
nor UO_2702 (O_2702,N_23125,N_24497);
or UO_2703 (O_2703,N_24108,N_23357);
or UO_2704 (O_2704,N_23398,N_24534);
and UO_2705 (O_2705,N_22561,N_24805);
nor UO_2706 (O_2706,N_24553,N_24009);
nor UO_2707 (O_2707,N_24153,N_23272);
nor UO_2708 (O_2708,N_23275,N_23007);
and UO_2709 (O_2709,N_23485,N_24476);
nor UO_2710 (O_2710,N_23420,N_22549);
nor UO_2711 (O_2711,N_23024,N_24027);
nor UO_2712 (O_2712,N_24315,N_24524);
or UO_2713 (O_2713,N_22547,N_24159);
nand UO_2714 (O_2714,N_24357,N_23675);
or UO_2715 (O_2715,N_22886,N_22808);
nand UO_2716 (O_2716,N_22995,N_24470);
or UO_2717 (O_2717,N_23598,N_23645);
nor UO_2718 (O_2718,N_23650,N_24915);
nand UO_2719 (O_2719,N_24652,N_24310);
xor UO_2720 (O_2720,N_23801,N_23769);
nand UO_2721 (O_2721,N_22562,N_23310);
or UO_2722 (O_2722,N_22655,N_23780);
nor UO_2723 (O_2723,N_24056,N_22717);
nor UO_2724 (O_2724,N_24454,N_24066);
or UO_2725 (O_2725,N_23956,N_24682);
and UO_2726 (O_2726,N_22558,N_24609);
or UO_2727 (O_2727,N_24911,N_22907);
nand UO_2728 (O_2728,N_24573,N_24620);
nand UO_2729 (O_2729,N_22699,N_24482);
nor UO_2730 (O_2730,N_22612,N_22825);
and UO_2731 (O_2731,N_22796,N_23898);
nand UO_2732 (O_2732,N_23902,N_22717);
or UO_2733 (O_2733,N_22942,N_22756);
nor UO_2734 (O_2734,N_24439,N_24437);
or UO_2735 (O_2735,N_24893,N_24298);
nand UO_2736 (O_2736,N_24222,N_23998);
nor UO_2737 (O_2737,N_23637,N_22578);
nor UO_2738 (O_2738,N_23610,N_24649);
nor UO_2739 (O_2739,N_24389,N_22707);
and UO_2740 (O_2740,N_23543,N_23530);
or UO_2741 (O_2741,N_24377,N_23755);
or UO_2742 (O_2742,N_23865,N_24426);
and UO_2743 (O_2743,N_23683,N_24188);
nand UO_2744 (O_2744,N_24858,N_22563);
or UO_2745 (O_2745,N_22665,N_24347);
nand UO_2746 (O_2746,N_24477,N_24676);
nand UO_2747 (O_2747,N_23579,N_23982);
nand UO_2748 (O_2748,N_24438,N_24085);
and UO_2749 (O_2749,N_23949,N_23939);
or UO_2750 (O_2750,N_22980,N_24690);
and UO_2751 (O_2751,N_23220,N_23825);
and UO_2752 (O_2752,N_23079,N_24942);
or UO_2753 (O_2753,N_23060,N_24486);
nor UO_2754 (O_2754,N_24163,N_24042);
and UO_2755 (O_2755,N_24429,N_22796);
nor UO_2756 (O_2756,N_24994,N_24931);
nand UO_2757 (O_2757,N_22829,N_24022);
or UO_2758 (O_2758,N_23182,N_23595);
nand UO_2759 (O_2759,N_24696,N_23349);
nand UO_2760 (O_2760,N_24935,N_23514);
nand UO_2761 (O_2761,N_24991,N_24668);
nor UO_2762 (O_2762,N_23903,N_22505);
or UO_2763 (O_2763,N_23387,N_22523);
nor UO_2764 (O_2764,N_23186,N_23778);
nor UO_2765 (O_2765,N_23186,N_23574);
and UO_2766 (O_2766,N_24965,N_22550);
or UO_2767 (O_2767,N_23797,N_23151);
nand UO_2768 (O_2768,N_23953,N_23433);
nand UO_2769 (O_2769,N_24687,N_23784);
nor UO_2770 (O_2770,N_24432,N_22889);
or UO_2771 (O_2771,N_24960,N_23627);
nor UO_2772 (O_2772,N_23703,N_23146);
or UO_2773 (O_2773,N_23705,N_23410);
nor UO_2774 (O_2774,N_23466,N_23116);
and UO_2775 (O_2775,N_23038,N_23903);
or UO_2776 (O_2776,N_24613,N_24399);
or UO_2777 (O_2777,N_24411,N_24297);
nand UO_2778 (O_2778,N_22883,N_23793);
or UO_2779 (O_2779,N_23329,N_23145);
nor UO_2780 (O_2780,N_24021,N_24324);
nand UO_2781 (O_2781,N_23188,N_22577);
or UO_2782 (O_2782,N_22815,N_23499);
nor UO_2783 (O_2783,N_22804,N_24645);
and UO_2784 (O_2784,N_24921,N_23246);
nand UO_2785 (O_2785,N_22965,N_23659);
and UO_2786 (O_2786,N_24102,N_22631);
nor UO_2787 (O_2787,N_23485,N_23994);
nand UO_2788 (O_2788,N_23422,N_24554);
or UO_2789 (O_2789,N_23553,N_24453);
nor UO_2790 (O_2790,N_24630,N_23494);
and UO_2791 (O_2791,N_24233,N_23095);
and UO_2792 (O_2792,N_24310,N_24657);
and UO_2793 (O_2793,N_22596,N_22995);
nor UO_2794 (O_2794,N_23423,N_24132);
and UO_2795 (O_2795,N_22593,N_23790);
nor UO_2796 (O_2796,N_23862,N_22531);
nor UO_2797 (O_2797,N_22804,N_24185);
or UO_2798 (O_2798,N_23140,N_22614);
or UO_2799 (O_2799,N_24177,N_23195);
or UO_2800 (O_2800,N_22704,N_24397);
nand UO_2801 (O_2801,N_23521,N_23380);
or UO_2802 (O_2802,N_22639,N_22768);
and UO_2803 (O_2803,N_23329,N_23542);
and UO_2804 (O_2804,N_22630,N_24363);
nor UO_2805 (O_2805,N_24911,N_23249);
nand UO_2806 (O_2806,N_23153,N_22522);
nor UO_2807 (O_2807,N_24724,N_22956);
nand UO_2808 (O_2808,N_22860,N_23563);
and UO_2809 (O_2809,N_23271,N_24902);
and UO_2810 (O_2810,N_23401,N_24489);
or UO_2811 (O_2811,N_23359,N_24243);
and UO_2812 (O_2812,N_22625,N_22977);
nand UO_2813 (O_2813,N_24164,N_23801);
or UO_2814 (O_2814,N_24480,N_24006);
nor UO_2815 (O_2815,N_24580,N_22734);
or UO_2816 (O_2816,N_22890,N_24023);
and UO_2817 (O_2817,N_22649,N_24731);
and UO_2818 (O_2818,N_23164,N_23690);
and UO_2819 (O_2819,N_23303,N_22660);
or UO_2820 (O_2820,N_24924,N_22837);
nor UO_2821 (O_2821,N_24727,N_22920);
nand UO_2822 (O_2822,N_23776,N_23934);
or UO_2823 (O_2823,N_24498,N_24748);
nor UO_2824 (O_2824,N_24111,N_24965);
nor UO_2825 (O_2825,N_23476,N_23912);
and UO_2826 (O_2826,N_24668,N_24634);
and UO_2827 (O_2827,N_24741,N_22547);
and UO_2828 (O_2828,N_22660,N_23426);
nand UO_2829 (O_2829,N_23381,N_23533);
and UO_2830 (O_2830,N_24229,N_24990);
or UO_2831 (O_2831,N_23925,N_23968);
nor UO_2832 (O_2832,N_24531,N_24247);
nor UO_2833 (O_2833,N_22927,N_24110);
and UO_2834 (O_2834,N_22694,N_23180);
nor UO_2835 (O_2835,N_24212,N_23182);
and UO_2836 (O_2836,N_24504,N_22948);
nand UO_2837 (O_2837,N_23882,N_24856);
nor UO_2838 (O_2838,N_22820,N_23454);
nand UO_2839 (O_2839,N_23602,N_23572);
or UO_2840 (O_2840,N_22540,N_23514);
and UO_2841 (O_2841,N_23200,N_23671);
and UO_2842 (O_2842,N_24370,N_23338);
nand UO_2843 (O_2843,N_23194,N_24386);
nand UO_2844 (O_2844,N_23379,N_24788);
or UO_2845 (O_2845,N_24950,N_22907);
or UO_2846 (O_2846,N_22948,N_24930);
and UO_2847 (O_2847,N_23831,N_23662);
nand UO_2848 (O_2848,N_22912,N_23036);
or UO_2849 (O_2849,N_24811,N_24621);
nand UO_2850 (O_2850,N_23402,N_23491);
and UO_2851 (O_2851,N_23069,N_24557);
nor UO_2852 (O_2852,N_23825,N_24622);
nand UO_2853 (O_2853,N_24719,N_23327);
nor UO_2854 (O_2854,N_22634,N_23923);
or UO_2855 (O_2855,N_24887,N_24617);
nor UO_2856 (O_2856,N_24651,N_24273);
and UO_2857 (O_2857,N_24557,N_24676);
nor UO_2858 (O_2858,N_22560,N_24956);
nor UO_2859 (O_2859,N_24832,N_24247);
nand UO_2860 (O_2860,N_24259,N_23242);
nor UO_2861 (O_2861,N_24382,N_22539);
and UO_2862 (O_2862,N_24657,N_22949);
and UO_2863 (O_2863,N_22927,N_22711);
nor UO_2864 (O_2864,N_23914,N_24762);
or UO_2865 (O_2865,N_23957,N_23415);
nand UO_2866 (O_2866,N_23403,N_24281);
nand UO_2867 (O_2867,N_22835,N_23515);
nor UO_2868 (O_2868,N_23578,N_24536);
nor UO_2869 (O_2869,N_22846,N_22682);
nor UO_2870 (O_2870,N_22683,N_23441);
or UO_2871 (O_2871,N_22922,N_24555);
or UO_2872 (O_2872,N_23464,N_22937);
and UO_2873 (O_2873,N_24651,N_22907);
or UO_2874 (O_2874,N_23747,N_23999);
nand UO_2875 (O_2875,N_24092,N_23066);
nor UO_2876 (O_2876,N_22933,N_23894);
nor UO_2877 (O_2877,N_22608,N_22846);
nand UO_2878 (O_2878,N_24497,N_22960);
or UO_2879 (O_2879,N_23610,N_23435);
nand UO_2880 (O_2880,N_23670,N_23618);
nand UO_2881 (O_2881,N_22848,N_24058);
nor UO_2882 (O_2882,N_23346,N_24216);
xor UO_2883 (O_2883,N_24473,N_24564);
and UO_2884 (O_2884,N_24419,N_24463);
and UO_2885 (O_2885,N_22764,N_22966);
or UO_2886 (O_2886,N_22811,N_24964);
or UO_2887 (O_2887,N_22966,N_23745);
and UO_2888 (O_2888,N_22713,N_23459);
nand UO_2889 (O_2889,N_23050,N_23333);
or UO_2890 (O_2890,N_24594,N_23165);
nand UO_2891 (O_2891,N_23299,N_23208);
and UO_2892 (O_2892,N_23746,N_24331);
nand UO_2893 (O_2893,N_22848,N_24569);
or UO_2894 (O_2894,N_22953,N_23730);
and UO_2895 (O_2895,N_24604,N_24631);
and UO_2896 (O_2896,N_24505,N_22722);
or UO_2897 (O_2897,N_24993,N_24166);
or UO_2898 (O_2898,N_24960,N_23817);
and UO_2899 (O_2899,N_24100,N_22835);
or UO_2900 (O_2900,N_23406,N_23187);
and UO_2901 (O_2901,N_23682,N_24337);
nand UO_2902 (O_2902,N_23287,N_24232);
or UO_2903 (O_2903,N_23234,N_23210);
or UO_2904 (O_2904,N_24056,N_24364);
nor UO_2905 (O_2905,N_24550,N_23967);
nand UO_2906 (O_2906,N_23793,N_23925);
nand UO_2907 (O_2907,N_24959,N_23536);
nand UO_2908 (O_2908,N_22904,N_22525);
or UO_2909 (O_2909,N_24600,N_24336);
and UO_2910 (O_2910,N_23838,N_24858);
nor UO_2911 (O_2911,N_24927,N_24866);
and UO_2912 (O_2912,N_22567,N_23234);
nand UO_2913 (O_2913,N_22534,N_23946);
nand UO_2914 (O_2914,N_23130,N_22601);
or UO_2915 (O_2915,N_22734,N_23358);
or UO_2916 (O_2916,N_24963,N_22775);
nand UO_2917 (O_2917,N_23004,N_23243);
nand UO_2918 (O_2918,N_24997,N_23383);
nand UO_2919 (O_2919,N_24834,N_23358);
and UO_2920 (O_2920,N_22738,N_23243);
nor UO_2921 (O_2921,N_22826,N_22781);
nand UO_2922 (O_2922,N_23361,N_23913);
nor UO_2923 (O_2923,N_23701,N_24704);
or UO_2924 (O_2924,N_23637,N_24042);
nor UO_2925 (O_2925,N_24664,N_23722);
nand UO_2926 (O_2926,N_23553,N_23868);
or UO_2927 (O_2927,N_23765,N_24374);
nor UO_2928 (O_2928,N_24746,N_24138);
nor UO_2929 (O_2929,N_23719,N_24290);
or UO_2930 (O_2930,N_23024,N_22953);
and UO_2931 (O_2931,N_24424,N_23261);
and UO_2932 (O_2932,N_23040,N_24029);
nor UO_2933 (O_2933,N_23109,N_24173);
nand UO_2934 (O_2934,N_24472,N_23681);
nor UO_2935 (O_2935,N_23605,N_24784);
or UO_2936 (O_2936,N_23609,N_24508);
nand UO_2937 (O_2937,N_22519,N_24337);
nand UO_2938 (O_2938,N_24215,N_24476);
and UO_2939 (O_2939,N_23726,N_22923);
nand UO_2940 (O_2940,N_24193,N_24130);
nor UO_2941 (O_2941,N_23287,N_24272);
nand UO_2942 (O_2942,N_23080,N_24645);
or UO_2943 (O_2943,N_24874,N_24099);
or UO_2944 (O_2944,N_23739,N_22684);
nand UO_2945 (O_2945,N_24047,N_23425);
and UO_2946 (O_2946,N_22957,N_23814);
or UO_2947 (O_2947,N_23808,N_24679);
nand UO_2948 (O_2948,N_24346,N_23121);
nand UO_2949 (O_2949,N_24367,N_24639);
or UO_2950 (O_2950,N_23976,N_23939);
nand UO_2951 (O_2951,N_24929,N_23761);
and UO_2952 (O_2952,N_24295,N_23709);
or UO_2953 (O_2953,N_23879,N_24968);
nand UO_2954 (O_2954,N_22612,N_23364);
and UO_2955 (O_2955,N_22515,N_24192);
or UO_2956 (O_2956,N_23016,N_24170);
nor UO_2957 (O_2957,N_24135,N_23696);
nand UO_2958 (O_2958,N_24574,N_24958);
and UO_2959 (O_2959,N_23832,N_24651);
nor UO_2960 (O_2960,N_23538,N_24214);
or UO_2961 (O_2961,N_23303,N_23359);
nand UO_2962 (O_2962,N_23736,N_23446);
or UO_2963 (O_2963,N_22743,N_23427);
and UO_2964 (O_2964,N_22618,N_24052);
or UO_2965 (O_2965,N_23168,N_23569);
nor UO_2966 (O_2966,N_23597,N_24103);
nor UO_2967 (O_2967,N_24909,N_23608);
or UO_2968 (O_2968,N_22687,N_22981);
nor UO_2969 (O_2969,N_22981,N_24181);
or UO_2970 (O_2970,N_22871,N_23935);
and UO_2971 (O_2971,N_24874,N_24879);
and UO_2972 (O_2972,N_24498,N_23792);
and UO_2973 (O_2973,N_23078,N_22516);
nor UO_2974 (O_2974,N_24202,N_22990);
and UO_2975 (O_2975,N_24805,N_23353);
nor UO_2976 (O_2976,N_22972,N_22642);
nor UO_2977 (O_2977,N_24657,N_23666);
or UO_2978 (O_2978,N_23010,N_24989);
and UO_2979 (O_2979,N_23911,N_24618);
nand UO_2980 (O_2980,N_24401,N_23805);
and UO_2981 (O_2981,N_23434,N_22720);
or UO_2982 (O_2982,N_23483,N_22846);
and UO_2983 (O_2983,N_24538,N_23369);
nand UO_2984 (O_2984,N_23437,N_23053);
or UO_2985 (O_2985,N_22747,N_23581);
nand UO_2986 (O_2986,N_23073,N_23548);
xor UO_2987 (O_2987,N_24664,N_24198);
nand UO_2988 (O_2988,N_23433,N_23640);
nor UO_2989 (O_2989,N_23791,N_23537);
or UO_2990 (O_2990,N_23682,N_23659);
and UO_2991 (O_2991,N_23989,N_23532);
nand UO_2992 (O_2992,N_24084,N_23337);
and UO_2993 (O_2993,N_22575,N_24080);
or UO_2994 (O_2994,N_24055,N_22558);
or UO_2995 (O_2995,N_23041,N_24595);
and UO_2996 (O_2996,N_23386,N_23263);
and UO_2997 (O_2997,N_22524,N_24488);
and UO_2998 (O_2998,N_22839,N_24396);
and UO_2999 (O_2999,N_23000,N_23012);
endmodule