module basic_1000_10000_1500_4_levels_2xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
nand U0 (N_0,In_629,In_893);
nor U1 (N_1,In_744,In_392);
or U2 (N_2,In_244,In_367);
nor U3 (N_3,In_647,In_427);
or U4 (N_4,In_37,In_612);
nor U5 (N_5,In_884,In_762);
nand U6 (N_6,In_257,In_987);
and U7 (N_7,In_325,In_695);
nand U8 (N_8,In_761,In_313);
or U9 (N_9,In_352,In_596);
and U10 (N_10,In_890,In_779);
and U11 (N_11,In_384,In_318);
or U12 (N_12,In_930,In_804);
nor U13 (N_13,In_64,In_30);
or U14 (N_14,In_599,In_56);
nor U15 (N_15,In_93,In_946);
nor U16 (N_16,In_232,In_404);
nor U17 (N_17,In_171,In_640);
and U18 (N_18,In_721,In_788);
or U19 (N_19,In_792,In_44);
and U20 (N_20,In_403,In_219);
and U21 (N_21,In_678,In_197);
and U22 (N_22,In_148,In_113);
or U23 (N_23,In_110,In_593);
nor U24 (N_24,In_9,In_388);
nor U25 (N_25,In_862,In_674);
nand U26 (N_26,In_787,In_574);
and U27 (N_27,In_423,In_133);
nand U28 (N_28,In_181,In_769);
or U29 (N_29,In_322,In_875);
or U30 (N_30,In_157,In_940);
or U31 (N_31,In_797,In_477);
nor U32 (N_32,In_342,In_880);
or U33 (N_33,In_752,In_253);
and U34 (N_34,In_434,In_357);
nor U35 (N_35,In_786,In_141);
nor U36 (N_36,In_425,In_421);
and U37 (N_37,In_311,In_484);
nand U38 (N_38,In_962,In_20);
nand U39 (N_39,In_233,In_487);
nand U40 (N_40,In_859,In_591);
nor U41 (N_41,In_334,In_570);
and U42 (N_42,In_132,In_210);
xor U43 (N_43,In_472,In_346);
or U44 (N_44,In_745,In_530);
and U45 (N_45,In_691,In_700);
nand U46 (N_46,In_422,In_290);
nand U47 (N_47,In_375,In_843);
and U48 (N_48,In_662,In_348);
nand U49 (N_49,In_77,In_5);
xor U50 (N_50,In_426,In_920);
nand U51 (N_51,In_852,In_383);
nand U52 (N_52,In_672,In_904);
nor U53 (N_53,In_925,In_807);
nand U54 (N_54,In_551,In_619);
nand U55 (N_55,In_517,In_473);
or U56 (N_56,In_305,In_448);
xnor U57 (N_57,In_659,In_889);
and U58 (N_58,In_588,In_833);
xnor U59 (N_59,In_496,In_12);
nor U60 (N_60,In_306,In_255);
and U61 (N_61,In_708,In_319);
xor U62 (N_62,In_623,In_967);
and U63 (N_63,In_160,In_541);
nor U64 (N_64,In_656,In_768);
nand U65 (N_65,In_784,In_193);
xor U66 (N_66,In_853,In_929);
nor U67 (N_67,In_846,In_83);
nor U68 (N_68,In_989,In_568);
or U69 (N_69,In_870,In_598);
nor U70 (N_70,In_349,In_312);
and U71 (N_71,In_912,In_43);
or U72 (N_72,In_972,In_370);
and U73 (N_73,In_54,In_380);
or U74 (N_74,In_543,In_876);
nor U75 (N_75,In_918,In_275);
nand U76 (N_76,In_184,In_478);
nor U77 (N_77,In_634,In_394);
nor U78 (N_78,In_10,In_158);
nor U79 (N_79,In_699,In_41);
nand U80 (N_80,In_605,In_172);
nor U81 (N_81,In_379,In_645);
and U82 (N_82,In_594,In_213);
nand U83 (N_83,In_439,In_958);
nand U84 (N_84,In_316,In_980);
nand U85 (N_85,In_838,In_268);
xor U86 (N_86,In_636,In_653);
nor U87 (N_87,In_2,In_65);
and U88 (N_88,In_327,In_463);
nor U89 (N_89,In_207,In_152);
nor U90 (N_90,In_242,In_888);
nor U91 (N_91,In_39,In_821);
and U92 (N_92,In_75,In_916);
or U93 (N_93,In_240,In_173);
or U94 (N_94,In_990,In_664);
nand U95 (N_95,In_883,In_225);
or U96 (N_96,In_715,In_983);
nand U97 (N_97,In_975,In_446);
nand U98 (N_98,In_732,In_302);
or U99 (N_99,In_187,In_33);
nand U100 (N_100,In_999,In_689);
nor U101 (N_101,In_597,In_581);
and U102 (N_102,In_651,In_707);
nor U103 (N_103,In_694,In_80);
nor U104 (N_104,In_239,In_615);
nand U105 (N_105,In_696,In_856);
and U106 (N_106,In_750,In_292);
and U107 (N_107,In_776,In_974);
and U108 (N_108,In_410,In_996);
xor U109 (N_109,In_397,In_498);
and U110 (N_110,In_964,In_151);
or U111 (N_111,In_419,In_176);
nor U112 (N_112,In_330,In_886);
or U113 (N_113,In_993,In_355);
or U114 (N_114,In_481,In_587);
nand U115 (N_115,In_770,In_16);
and U116 (N_116,In_931,In_328);
and U117 (N_117,In_222,In_680);
and U118 (N_118,In_248,In_402);
nor U119 (N_119,In_21,In_516);
nor U120 (N_120,In_848,In_278);
nand U121 (N_121,In_50,In_351);
nor U122 (N_122,In_710,In_178);
nor U123 (N_123,In_923,In_329);
nand U124 (N_124,In_280,In_238);
nor U125 (N_125,In_430,In_542);
and U126 (N_126,In_153,In_466);
or U127 (N_127,In_345,In_72);
nand U128 (N_128,In_569,In_897);
nand U129 (N_129,In_970,In_869);
nor U130 (N_130,In_87,In_376);
and U131 (N_131,In_725,In_910);
nand U132 (N_132,In_857,In_147);
or U133 (N_133,In_17,In_631);
nor U134 (N_134,In_953,In_417);
nor U135 (N_135,In_648,In_438);
or U136 (N_136,In_604,In_489);
or U137 (N_137,In_566,In_561);
nor U138 (N_138,In_727,In_298);
or U139 (N_139,In_456,In_667);
nor U140 (N_140,In_200,In_584);
nor U141 (N_141,In_373,In_411);
and U142 (N_142,In_490,In_296);
nand U143 (N_143,In_76,In_390);
and U144 (N_144,In_690,In_511);
or U145 (N_145,In_978,In_994);
or U146 (N_146,In_703,In_709);
nand U147 (N_147,In_803,In_23);
nand U148 (N_148,In_465,In_524);
xor U149 (N_149,In_191,In_682);
or U150 (N_150,In_767,In_273);
and U151 (N_151,In_717,In_464);
nor U152 (N_152,In_102,In_673);
nor U153 (N_153,In_670,In_863);
nor U154 (N_154,In_722,In_865);
xnor U155 (N_155,In_266,In_36);
nor U156 (N_156,In_704,In_63);
nand U157 (N_157,In_228,In_968);
nand U158 (N_158,In_576,In_751);
or U159 (N_159,In_476,In_227);
and U160 (N_160,In_378,In_74);
nand U161 (N_161,In_186,In_557);
and U162 (N_162,In_168,In_189);
nand U163 (N_163,In_250,In_830);
or U164 (N_164,In_733,In_909);
nor U165 (N_165,In_795,In_208);
nand U166 (N_166,In_161,In_97);
nor U167 (N_167,In_766,In_494);
nor U168 (N_168,In_461,In_272);
nor U169 (N_169,In_179,In_201);
nor U170 (N_170,In_510,In_553);
and U171 (N_171,In_354,In_501);
nor U172 (N_172,In_130,In_933);
and U173 (N_173,In_560,In_523);
and U174 (N_174,In_460,In_3);
or U175 (N_175,In_131,In_22);
or U176 (N_176,In_149,In_229);
nand U177 (N_177,In_984,In_7);
nor U178 (N_178,In_366,In_395);
and U179 (N_179,In_337,In_190);
nor U180 (N_180,In_760,In_246);
nand U181 (N_181,In_895,In_881);
and U182 (N_182,In_300,In_961);
nor U183 (N_183,In_457,In_572);
or U184 (N_184,In_121,In_163);
xnor U185 (N_185,In_669,In_42);
nor U186 (N_186,In_365,In_264);
and U187 (N_187,In_758,In_861);
nor U188 (N_188,In_416,In_998);
nand U189 (N_189,In_782,In_374);
nand U190 (N_190,In_981,In_759);
and U191 (N_191,In_467,In_332);
and U192 (N_192,In_155,In_814);
nor U193 (N_193,In_84,In_8);
nor U194 (N_194,In_538,In_661);
and U195 (N_195,In_211,In_741);
nand U196 (N_196,In_536,In_199);
and U197 (N_197,In_724,In_844);
or U198 (N_198,In_169,In_713);
nor U199 (N_199,In_559,In_632);
nor U200 (N_200,In_735,In_217);
or U201 (N_201,In_982,In_934);
and U202 (N_202,In_548,In_164);
or U203 (N_203,In_486,In_19);
and U204 (N_204,In_205,In_748);
and U205 (N_205,In_714,In_407);
and U206 (N_206,In_79,In_364);
and U207 (N_207,In_522,In_252);
nor U208 (N_208,In_877,In_847);
or U209 (N_209,In_595,In_618);
nand U210 (N_210,In_668,In_116);
and U211 (N_211,In_837,In_726);
or U212 (N_212,In_474,In_124);
or U213 (N_213,In_902,In_635);
nor U214 (N_214,In_317,In_13);
or U215 (N_215,In_91,In_399);
nor U216 (N_216,In_798,In_59);
or U217 (N_217,In_96,In_879);
and U218 (N_218,In_765,In_772);
nor U219 (N_219,In_192,In_85);
or U220 (N_220,In_749,In_582);
or U221 (N_221,In_125,In_256);
nor U222 (N_222,In_675,In_224);
or U223 (N_223,In_254,In_815);
nor U224 (N_224,In_137,In_127);
and U225 (N_225,In_260,In_420);
or U226 (N_226,In_545,In_734);
and U227 (N_227,In_401,In_949);
and U228 (N_228,In_90,In_347);
or U229 (N_229,In_601,In_550);
or U230 (N_230,In_747,In_284);
and U231 (N_231,In_488,In_663);
nor U232 (N_232,In_534,In_61);
or U233 (N_233,In_445,In_796);
and U234 (N_234,In_14,In_406);
nand U235 (N_235,In_180,In_681);
or U236 (N_236,In_204,In_114);
xnor U237 (N_237,In_485,In_607);
nor U238 (N_238,In_819,In_447);
nor U239 (N_239,In_68,In_899);
or U240 (N_240,In_976,In_0);
nor U241 (N_241,In_515,In_697);
nand U242 (N_242,In_908,In_692);
nor U243 (N_243,In_756,In_941);
or U244 (N_244,In_808,In_389);
and U245 (N_245,In_927,In_780);
and U246 (N_246,In_73,In_633);
or U247 (N_247,In_391,In_297);
nor U248 (N_248,In_509,In_138);
nand U249 (N_249,In_109,In_602);
nand U250 (N_250,In_665,In_649);
xor U251 (N_251,In_156,In_939);
or U252 (N_252,In_269,In_450);
nand U253 (N_253,In_911,In_47);
nor U254 (N_254,In_282,In_757);
or U255 (N_255,In_362,In_935);
or U256 (N_256,In_644,In_236);
nor U257 (N_257,In_52,In_818);
or U258 (N_258,In_276,In_554);
or U259 (N_259,In_105,In_740);
nand U260 (N_260,In_202,In_432);
nand U261 (N_261,In_616,In_608);
nand U262 (N_262,In_754,In_951);
nand U263 (N_263,In_177,In_531);
nor U264 (N_264,In_431,In_965);
or U265 (N_265,In_475,In_556);
and U266 (N_266,In_359,In_95);
nor U267 (N_267,In_834,In_907);
or U268 (N_268,In_307,In_314);
nand U269 (N_269,In_851,In_283);
nand U270 (N_270,In_539,In_995);
nand U271 (N_271,In_251,In_88);
nor U272 (N_272,In_781,In_519);
nor U273 (N_273,In_145,In_791);
nor U274 (N_274,In_643,In_94);
nand U275 (N_275,In_209,In_288);
or U276 (N_276,In_57,In_973);
and U277 (N_277,In_705,In_492);
nor U278 (N_278,In_241,In_583);
nand U279 (N_279,In_112,In_957);
nand U280 (N_280,In_926,In_600);
nand U281 (N_281,In_919,In_26);
nor U282 (N_282,In_728,In_777);
nor U283 (N_283,In_353,In_736);
and U284 (N_284,In_514,In_885);
nor U285 (N_285,In_706,In_529);
nor U286 (N_286,In_55,In_943);
or U287 (N_287,In_111,In_398);
and U288 (N_288,In_455,In_773);
or U289 (N_289,In_842,In_100);
or U290 (N_290,In_140,In_563);
nand U291 (N_291,In_482,In_413);
nor U292 (N_292,In_986,In_646);
and U293 (N_293,In_118,In_535);
and U294 (N_294,In_45,In_136);
and U295 (N_295,In_997,In_294);
and U296 (N_296,In_945,In_469);
and U297 (N_297,In_866,In_611);
and U298 (N_298,In_871,In_533);
or U299 (N_299,In_462,In_28);
nand U300 (N_300,In_743,In_609);
nor U301 (N_301,In_360,In_99);
nand U302 (N_302,In_580,In_960);
or U303 (N_303,In_753,In_723);
and U304 (N_304,In_279,In_579);
nand U305 (N_305,In_237,In_82);
or U306 (N_306,In_428,In_142);
nand U307 (N_307,In_258,In_154);
and U308 (N_308,In_104,In_340);
and U309 (N_309,In_32,In_120);
or U310 (N_310,In_840,In_805);
or U311 (N_311,In_738,In_433);
nor U312 (N_312,In_825,In_820);
and U313 (N_313,In_11,In_67);
or U314 (N_314,In_234,In_70);
and U315 (N_315,In_684,In_301);
nor U316 (N_316,In_249,In_746);
and U317 (N_317,In_513,In_954);
and U318 (N_318,In_671,In_122);
nand U319 (N_319,In_15,In_339);
nand U320 (N_320,In_443,In_129);
or U321 (N_321,In_764,In_547);
nor U322 (N_322,In_48,In_686);
nor U323 (N_323,In_285,In_414);
nand U324 (N_324,In_552,In_144);
nor U325 (N_325,In_265,In_737);
nor U326 (N_326,In_409,In_827);
and U327 (N_327,In_385,In_799);
nor U328 (N_328,In_702,In_29);
nor U329 (N_329,In_679,In_898);
and U330 (N_330,In_849,In_206);
nor U331 (N_331,In_626,In_326);
or U332 (N_332,In_274,In_40);
nand U333 (N_333,In_216,In_991);
and U334 (N_334,In_261,In_742);
or U335 (N_335,In_162,In_66);
and U336 (N_336,In_310,In_377);
and U337 (N_337,In_625,In_549);
nand U338 (N_338,In_226,In_315);
or U339 (N_339,In_677,In_698);
or U340 (N_340,In_812,In_590);
nand U341 (N_341,In_182,In_174);
nor U342 (N_342,In_215,In_525);
and U343 (N_343,In_247,In_537);
nand U344 (N_344,In_882,In_555);
nand U345 (N_345,In_540,In_719);
or U346 (N_346,In_658,In_18);
nand U347 (N_347,In_586,In_324);
nor U348 (N_348,In_175,In_829);
nor U349 (N_349,In_165,In_836);
nand U350 (N_350,In_654,In_720);
nor U351 (N_351,In_143,In_763);
or U352 (N_352,In_624,In_495);
or U353 (N_353,In_676,In_135);
or U354 (N_354,In_578,In_277);
and U355 (N_355,In_458,In_195);
or U356 (N_356,In_518,In_436);
nor U357 (N_357,In_491,In_824);
nand U358 (N_358,In_955,In_479);
and U359 (N_359,In_243,In_900);
and U360 (N_360,In_128,In_739);
or U361 (N_361,In_166,In_860);
and U362 (N_362,In_71,In_103);
and U363 (N_363,In_755,In_874);
and U364 (N_364,In_299,In_89);
nand U365 (N_365,In_571,In_235);
nand U366 (N_366,In_901,In_544);
nor U367 (N_367,In_321,In_230);
or U368 (N_368,In_429,In_785);
and U369 (N_369,In_817,In_31);
nand U370 (N_370,In_139,In_577);
nand U371 (N_371,In_183,In_630);
nor U372 (N_372,In_850,In_873);
nor U373 (N_373,In_521,In_731);
nor U374 (N_374,In_221,In_650);
nor U375 (N_375,In_712,In_813);
nand U376 (N_376,In_453,In_564);
xor U377 (N_377,In_49,In_614);
nor U378 (N_378,In_903,In_454);
nand U379 (N_379,In_638,In_620);
and U380 (N_380,In_198,In_948);
or U381 (N_381,In_203,In_683);
or U382 (N_382,In_642,In_592);
or U383 (N_383,In_444,In_471);
and U384 (N_384,In_778,In_959);
nor U385 (N_385,In_977,In_368);
nor U386 (N_386,In_69,In_641);
nand U387 (N_387,In_497,In_358);
nand U388 (N_388,In_98,In_854);
nor U389 (N_389,In_335,In_214);
or U390 (N_390,In_988,In_942);
nor U391 (N_391,In_480,In_46);
or U392 (N_392,In_452,In_532);
and U393 (N_393,In_24,In_966);
nand U394 (N_394,In_503,In_361);
nor U395 (N_395,In_412,In_979);
or U396 (N_396,In_822,In_839);
and U397 (N_397,In_101,In_891);
and U398 (N_398,In_371,In_286);
or U399 (N_399,In_526,In_639);
nand U400 (N_400,In_470,In_304);
or U401 (N_401,In_387,In_505);
nor U402 (N_402,In_499,In_864);
and U403 (N_403,In_915,In_652);
or U404 (N_404,In_701,In_573);
or U405 (N_405,In_4,In_126);
nand U406 (N_406,In_685,In_231);
nor U407 (N_407,In_621,In_35);
nand U408 (N_408,In_336,In_905);
or U409 (N_409,In_78,In_372);
and U410 (N_410,In_159,In_655);
or U411 (N_411,In_194,In_937);
or U412 (N_412,In_341,In_562);
and U413 (N_413,In_938,In_528);
and U414 (N_414,In_1,In_693);
or U415 (N_415,In_393,In_289);
nand U416 (N_416,In_123,In_944);
nand U417 (N_417,In_867,In_802);
and U418 (N_418,In_892,In_567);
nand U419 (N_419,In_134,In_512);
and U420 (N_420,In_783,In_263);
or U421 (N_421,In_811,In_823);
nor U422 (N_422,In_558,In_350);
and U423 (N_423,In_502,In_504);
or U424 (N_424,In_841,In_382);
nor U425 (N_425,In_493,In_921);
nor U426 (N_426,In_343,In_107);
or U427 (N_427,In_603,In_459);
nand U428 (N_428,In_575,In_223);
or U429 (N_429,In_483,In_320);
nand U430 (N_430,In_947,In_500);
nor U431 (N_431,In_188,In_212);
nand U432 (N_432,In_245,In_323);
nor U433 (N_433,In_51,In_441);
and U434 (N_434,In_952,In_657);
or U435 (N_435,In_449,In_170);
nor U436 (N_436,In_333,In_809);
nor U437 (N_437,In_917,In_816);
or U438 (N_438,In_622,In_25);
and U439 (N_439,In_950,In_344);
and U440 (N_440,In_932,In_381);
or U441 (N_441,In_58,In_878);
and U442 (N_442,In_868,In_295);
nand U443 (N_443,In_936,In_971);
nand U444 (N_444,In_828,In_835);
nor U445 (N_445,In_303,In_271);
or U446 (N_446,In_309,In_218);
nand U447 (N_447,In_716,In_627);
nor U448 (N_448,In_424,In_331);
nand U449 (N_449,In_565,In_196);
nand U450 (N_450,In_363,In_806);
nor U451 (N_451,In_281,In_356);
nand U452 (N_452,In_106,In_775);
nand U453 (N_453,In_771,In_270);
and U454 (N_454,In_914,In_53);
or U455 (N_455,In_985,In_27);
nand U456 (N_456,In_418,In_287);
nand U457 (N_457,In_913,In_831);
xor U458 (N_458,In_220,In_963);
or U459 (N_459,In_338,In_34);
and U460 (N_460,In_117,In_589);
xor U461 (N_461,In_86,In_400);
and U462 (N_462,In_832,In_520);
nor U463 (N_463,In_546,In_660);
or U464 (N_464,In_845,In_527);
and U465 (N_465,In_794,In_992);
nand U466 (N_466,In_408,In_506);
and U467 (N_467,In_451,In_711);
and U468 (N_468,In_606,In_826);
nand U469 (N_469,In_508,In_872);
nor U470 (N_470,In_617,In_60);
or U471 (N_471,In_688,In_896);
and U472 (N_472,In_293,In_810);
and U473 (N_473,In_259,In_793);
nand U474 (N_474,In_415,In_774);
nand U475 (N_475,In_610,In_790);
nor U476 (N_476,In_146,In_718);
or U477 (N_477,In_800,In_887);
or U478 (N_478,In_92,In_115);
nand U479 (N_479,In_185,In_396);
and U480 (N_480,In_405,In_730);
and U481 (N_481,In_922,In_167);
and U482 (N_482,In_291,In_894);
nand U483 (N_483,In_442,In_150);
and U484 (N_484,In_858,In_855);
nor U485 (N_485,In_308,In_507);
or U486 (N_486,In_613,In_628);
nand U487 (N_487,In_369,In_440);
and U488 (N_488,In_687,In_38);
nor U489 (N_489,In_6,In_267);
and U490 (N_490,In_801,In_435);
or U491 (N_491,In_956,In_62);
nand U492 (N_492,In_437,In_262);
nor U493 (N_493,In_906,In_969);
nand U494 (N_494,In_468,In_119);
nand U495 (N_495,In_928,In_637);
and U496 (N_496,In_924,In_81);
nand U497 (N_497,In_585,In_729);
nand U498 (N_498,In_108,In_666);
and U499 (N_499,In_789,In_386);
or U500 (N_500,In_914,In_782);
and U501 (N_501,In_431,In_368);
or U502 (N_502,In_944,In_827);
or U503 (N_503,In_312,In_100);
nand U504 (N_504,In_559,In_482);
nand U505 (N_505,In_836,In_865);
and U506 (N_506,In_332,In_347);
nor U507 (N_507,In_210,In_138);
or U508 (N_508,In_365,In_880);
nand U509 (N_509,In_421,In_643);
or U510 (N_510,In_967,In_872);
xor U511 (N_511,In_99,In_899);
nand U512 (N_512,In_70,In_940);
and U513 (N_513,In_935,In_483);
or U514 (N_514,In_271,In_4);
nand U515 (N_515,In_27,In_541);
and U516 (N_516,In_206,In_82);
or U517 (N_517,In_652,In_55);
and U518 (N_518,In_894,In_820);
nand U519 (N_519,In_216,In_556);
and U520 (N_520,In_438,In_552);
and U521 (N_521,In_474,In_352);
and U522 (N_522,In_867,In_902);
and U523 (N_523,In_414,In_175);
nor U524 (N_524,In_783,In_796);
nor U525 (N_525,In_246,In_891);
nand U526 (N_526,In_515,In_430);
nor U527 (N_527,In_224,In_535);
nand U528 (N_528,In_94,In_759);
nand U529 (N_529,In_53,In_465);
xor U530 (N_530,In_563,In_268);
or U531 (N_531,In_143,In_294);
and U532 (N_532,In_119,In_314);
nor U533 (N_533,In_199,In_30);
nor U534 (N_534,In_91,In_422);
nor U535 (N_535,In_925,In_604);
nand U536 (N_536,In_64,In_79);
or U537 (N_537,In_605,In_242);
or U538 (N_538,In_17,In_694);
or U539 (N_539,In_638,In_347);
nor U540 (N_540,In_364,In_474);
and U541 (N_541,In_960,In_407);
nand U542 (N_542,In_791,In_555);
nor U543 (N_543,In_796,In_669);
and U544 (N_544,In_151,In_708);
nand U545 (N_545,In_858,In_358);
and U546 (N_546,In_925,In_945);
or U547 (N_547,In_900,In_892);
nor U548 (N_548,In_226,In_959);
xor U549 (N_549,In_393,In_59);
nand U550 (N_550,In_114,In_34);
nand U551 (N_551,In_245,In_89);
or U552 (N_552,In_546,In_932);
nor U553 (N_553,In_847,In_660);
nor U554 (N_554,In_485,In_887);
and U555 (N_555,In_788,In_929);
nand U556 (N_556,In_207,In_421);
nor U557 (N_557,In_265,In_499);
and U558 (N_558,In_166,In_319);
xor U559 (N_559,In_952,In_32);
nor U560 (N_560,In_981,In_494);
nand U561 (N_561,In_942,In_25);
or U562 (N_562,In_612,In_742);
nor U563 (N_563,In_435,In_455);
nor U564 (N_564,In_155,In_25);
or U565 (N_565,In_14,In_716);
or U566 (N_566,In_185,In_61);
nor U567 (N_567,In_149,In_807);
nor U568 (N_568,In_848,In_781);
nor U569 (N_569,In_809,In_172);
and U570 (N_570,In_318,In_708);
nor U571 (N_571,In_272,In_267);
or U572 (N_572,In_493,In_49);
nand U573 (N_573,In_756,In_657);
nor U574 (N_574,In_974,In_468);
nor U575 (N_575,In_78,In_338);
nor U576 (N_576,In_247,In_182);
nand U577 (N_577,In_213,In_154);
nand U578 (N_578,In_515,In_959);
nand U579 (N_579,In_673,In_450);
and U580 (N_580,In_918,In_803);
nand U581 (N_581,In_256,In_337);
and U582 (N_582,In_563,In_865);
nand U583 (N_583,In_544,In_226);
and U584 (N_584,In_143,In_997);
nand U585 (N_585,In_216,In_590);
nand U586 (N_586,In_373,In_700);
nand U587 (N_587,In_874,In_746);
or U588 (N_588,In_153,In_234);
or U589 (N_589,In_53,In_961);
and U590 (N_590,In_454,In_89);
nand U591 (N_591,In_391,In_269);
nor U592 (N_592,In_98,In_111);
and U593 (N_593,In_120,In_772);
and U594 (N_594,In_1,In_201);
or U595 (N_595,In_397,In_905);
or U596 (N_596,In_573,In_13);
nor U597 (N_597,In_432,In_983);
nand U598 (N_598,In_614,In_442);
and U599 (N_599,In_274,In_479);
nor U600 (N_600,In_543,In_462);
or U601 (N_601,In_976,In_647);
nor U602 (N_602,In_969,In_635);
nor U603 (N_603,In_588,In_505);
nand U604 (N_604,In_334,In_976);
and U605 (N_605,In_790,In_655);
nand U606 (N_606,In_369,In_975);
or U607 (N_607,In_905,In_55);
nand U608 (N_608,In_863,In_616);
nor U609 (N_609,In_873,In_99);
nand U610 (N_610,In_740,In_232);
nand U611 (N_611,In_668,In_266);
and U612 (N_612,In_706,In_13);
nand U613 (N_613,In_525,In_407);
nor U614 (N_614,In_111,In_920);
and U615 (N_615,In_631,In_106);
and U616 (N_616,In_300,In_105);
nor U617 (N_617,In_634,In_969);
and U618 (N_618,In_354,In_246);
or U619 (N_619,In_123,In_117);
nand U620 (N_620,In_819,In_480);
and U621 (N_621,In_476,In_449);
and U622 (N_622,In_882,In_173);
and U623 (N_623,In_879,In_861);
nand U624 (N_624,In_194,In_140);
nor U625 (N_625,In_523,In_550);
and U626 (N_626,In_594,In_575);
nor U627 (N_627,In_137,In_854);
and U628 (N_628,In_893,In_86);
nor U629 (N_629,In_23,In_505);
nor U630 (N_630,In_997,In_176);
or U631 (N_631,In_100,In_606);
nand U632 (N_632,In_129,In_574);
and U633 (N_633,In_639,In_984);
or U634 (N_634,In_961,In_104);
nand U635 (N_635,In_444,In_658);
or U636 (N_636,In_322,In_331);
and U637 (N_637,In_874,In_414);
nand U638 (N_638,In_575,In_828);
nand U639 (N_639,In_482,In_3);
nor U640 (N_640,In_771,In_992);
nand U641 (N_641,In_353,In_442);
or U642 (N_642,In_255,In_405);
nand U643 (N_643,In_507,In_975);
nand U644 (N_644,In_449,In_118);
or U645 (N_645,In_859,In_282);
nand U646 (N_646,In_738,In_36);
or U647 (N_647,In_929,In_516);
nor U648 (N_648,In_438,In_615);
nor U649 (N_649,In_182,In_705);
and U650 (N_650,In_410,In_495);
nand U651 (N_651,In_615,In_780);
nand U652 (N_652,In_264,In_940);
xnor U653 (N_653,In_730,In_670);
nor U654 (N_654,In_364,In_336);
nor U655 (N_655,In_978,In_597);
nor U656 (N_656,In_958,In_851);
nor U657 (N_657,In_956,In_514);
nand U658 (N_658,In_220,In_438);
nand U659 (N_659,In_216,In_827);
nor U660 (N_660,In_353,In_947);
nand U661 (N_661,In_618,In_50);
nand U662 (N_662,In_489,In_704);
or U663 (N_663,In_748,In_536);
nor U664 (N_664,In_765,In_815);
and U665 (N_665,In_14,In_593);
nand U666 (N_666,In_476,In_434);
or U667 (N_667,In_367,In_164);
or U668 (N_668,In_38,In_724);
nand U669 (N_669,In_709,In_754);
or U670 (N_670,In_778,In_979);
nor U671 (N_671,In_281,In_985);
and U672 (N_672,In_646,In_688);
xor U673 (N_673,In_677,In_135);
or U674 (N_674,In_32,In_168);
nand U675 (N_675,In_436,In_510);
and U676 (N_676,In_44,In_695);
or U677 (N_677,In_345,In_270);
and U678 (N_678,In_211,In_563);
nand U679 (N_679,In_739,In_920);
nor U680 (N_680,In_791,In_114);
nor U681 (N_681,In_861,In_505);
nand U682 (N_682,In_428,In_953);
or U683 (N_683,In_325,In_229);
nor U684 (N_684,In_968,In_294);
nor U685 (N_685,In_784,In_356);
nand U686 (N_686,In_366,In_168);
nand U687 (N_687,In_353,In_914);
nand U688 (N_688,In_600,In_51);
and U689 (N_689,In_629,In_687);
and U690 (N_690,In_256,In_910);
nor U691 (N_691,In_29,In_710);
nand U692 (N_692,In_345,In_529);
nand U693 (N_693,In_332,In_15);
and U694 (N_694,In_509,In_528);
or U695 (N_695,In_447,In_403);
nand U696 (N_696,In_996,In_127);
or U697 (N_697,In_391,In_34);
nand U698 (N_698,In_565,In_979);
and U699 (N_699,In_493,In_38);
and U700 (N_700,In_177,In_637);
nor U701 (N_701,In_525,In_827);
nand U702 (N_702,In_948,In_801);
and U703 (N_703,In_707,In_987);
and U704 (N_704,In_758,In_245);
xor U705 (N_705,In_880,In_251);
nor U706 (N_706,In_17,In_876);
or U707 (N_707,In_596,In_715);
nor U708 (N_708,In_218,In_365);
nor U709 (N_709,In_204,In_499);
or U710 (N_710,In_293,In_823);
nand U711 (N_711,In_586,In_724);
nor U712 (N_712,In_939,In_344);
and U713 (N_713,In_991,In_116);
or U714 (N_714,In_525,In_797);
or U715 (N_715,In_866,In_209);
and U716 (N_716,In_534,In_441);
and U717 (N_717,In_336,In_638);
nor U718 (N_718,In_310,In_705);
nand U719 (N_719,In_211,In_788);
nor U720 (N_720,In_831,In_949);
nand U721 (N_721,In_883,In_597);
nand U722 (N_722,In_668,In_849);
nor U723 (N_723,In_39,In_256);
or U724 (N_724,In_43,In_941);
and U725 (N_725,In_868,In_856);
and U726 (N_726,In_426,In_629);
or U727 (N_727,In_715,In_973);
nand U728 (N_728,In_154,In_631);
nand U729 (N_729,In_886,In_504);
and U730 (N_730,In_593,In_645);
or U731 (N_731,In_483,In_979);
and U732 (N_732,In_624,In_730);
or U733 (N_733,In_8,In_347);
and U734 (N_734,In_377,In_809);
xnor U735 (N_735,In_145,In_506);
or U736 (N_736,In_818,In_579);
and U737 (N_737,In_725,In_719);
nand U738 (N_738,In_889,In_777);
and U739 (N_739,In_967,In_535);
or U740 (N_740,In_680,In_975);
nor U741 (N_741,In_193,In_600);
nor U742 (N_742,In_781,In_856);
and U743 (N_743,In_681,In_879);
nand U744 (N_744,In_500,In_74);
or U745 (N_745,In_627,In_844);
nand U746 (N_746,In_247,In_291);
xnor U747 (N_747,In_333,In_233);
nand U748 (N_748,In_276,In_363);
and U749 (N_749,In_464,In_791);
and U750 (N_750,In_711,In_981);
nor U751 (N_751,In_903,In_848);
or U752 (N_752,In_992,In_301);
nor U753 (N_753,In_614,In_725);
or U754 (N_754,In_795,In_181);
nor U755 (N_755,In_533,In_170);
nand U756 (N_756,In_512,In_89);
nand U757 (N_757,In_93,In_901);
and U758 (N_758,In_223,In_64);
or U759 (N_759,In_687,In_279);
nor U760 (N_760,In_325,In_261);
nor U761 (N_761,In_304,In_119);
nor U762 (N_762,In_567,In_234);
nor U763 (N_763,In_661,In_182);
nand U764 (N_764,In_771,In_416);
or U765 (N_765,In_714,In_735);
nand U766 (N_766,In_525,In_983);
or U767 (N_767,In_503,In_989);
and U768 (N_768,In_650,In_848);
or U769 (N_769,In_906,In_654);
nor U770 (N_770,In_982,In_154);
nand U771 (N_771,In_690,In_698);
or U772 (N_772,In_938,In_232);
or U773 (N_773,In_282,In_964);
and U774 (N_774,In_468,In_304);
or U775 (N_775,In_866,In_751);
and U776 (N_776,In_117,In_349);
nand U777 (N_777,In_142,In_538);
nor U778 (N_778,In_848,In_289);
xnor U779 (N_779,In_784,In_86);
nand U780 (N_780,In_985,In_635);
nand U781 (N_781,In_938,In_350);
and U782 (N_782,In_368,In_243);
and U783 (N_783,In_909,In_3);
nor U784 (N_784,In_762,In_616);
nor U785 (N_785,In_499,In_563);
nand U786 (N_786,In_794,In_79);
and U787 (N_787,In_929,In_767);
or U788 (N_788,In_121,In_136);
or U789 (N_789,In_359,In_55);
nand U790 (N_790,In_935,In_415);
nor U791 (N_791,In_538,In_245);
or U792 (N_792,In_824,In_643);
or U793 (N_793,In_752,In_180);
nor U794 (N_794,In_268,In_252);
or U795 (N_795,In_710,In_187);
nor U796 (N_796,In_967,In_414);
and U797 (N_797,In_221,In_191);
nand U798 (N_798,In_233,In_175);
nand U799 (N_799,In_248,In_909);
or U800 (N_800,In_808,In_382);
nand U801 (N_801,In_844,In_924);
and U802 (N_802,In_798,In_60);
nor U803 (N_803,In_651,In_32);
and U804 (N_804,In_104,In_805);
or U805 (N_805,In_399,In_29);
nand U806 (N_806,In_140,In_794);
nor U807 (N_807,In_151,In_309);
nor U808 (N_808,In_451,In_313);
and U809 (N_809,In_39,In_810);
and U810 (N_810,In_926,In_314);
nand U811 (N_811,In_892,In_100);
nand U812 (N_812,In_623,In_364);
nand U813 (N_813,In_421,In_43);
or U814 (N_814,In_354,In_227);
or U815 (N_815,In_411,In_612);
nand U816 (N_816,In_508,In_958);
nor U817 (N_817,In_722,In_890);
or U818 (N_818,In_389,In_593);
nand U819 (N_819,In_103,In_483);
and U820 (N_820,In_839,In_52);
nor U821 (N_821,In_774,In_52);
nand U822 (N_822,In_19,In_899);
and U823 (N_823,In_701,In_5);
or U824 (N_824,In_778,In_539);
nand U825 (N_825,In_991,In_922);
or U826 (N_826,In_13,In_561);
or U827 (N_827,In_317,In_645);
and U828 (N_828,In_125,In_908);
nor U829 (N_829,In_125,In_494);
and U830 (N_830,In_881,In_173);
nor U831 (N_831,In_298,In_293);
or U832 (N_832,In_990,In_821);
and U833 (N_833,In_890,In_767);
nand U834 (N_834,In_496,In_261);
and U835 (N_835,In_119,In_626);
nand U836 (N_836,In_113,In_691);
nor U837 (N_837,In_571,In_63);
and U838 (N_838,In_883,In_688);
nand U839 (N_839,In_633,In_202);
and U840 (N_840,In_714,In_890);
nor U841 (N_841,In_226,In_880);
or U842 (N_842,In_476,In_636);
nor U843 (N_843,In_480,In_330);
nor U844 (N_844,In_127,In_228);
nand U845 (N_845,In_834,In_491);
and U846 (N_846,In_974,In_546);
and U847 (N_847,In_179,In_998);
nor U848 (N_848,In_646,In_289);
or U849 (N_849,In_597,In_744);
xor U850 (N_850,In_26,In_781);
nand U851 (N_851,In_222,In_947);
or U852 (N_852,In_207,In_751);
or U853 (N_853,In_809,In_810);
or U854 (N_854,In_514,In_805);
nand U855 (N_855,In_232,In_22);
and U856 (N_856,In_327,In_186);
nor U857 (N_857,In_151,In_22);
and U858 (N_858,In_587,In_589);
or U859 (N_859,In_946,In_282);
nand U860 (N_860,In_345,In_646);
nor U861 (N_861,In_690,In_387);
or U862 (N_862,In_904,In_620);
or U863 (N_863,In_986,In_294);
nor U864 (N_864,In_959,In_39);
or U865 (N_865,In_969,In_513);
nand U866 (N_866,In_251,In_323);
and U867 (N_867,In_736,In_52);
nand U868 (N_868,In_371,In_711);
xnor U869 (N_869,In_257,In_583);
xnor U870 (N_870,In_840,In_969);
and U871 (N_871,In_372,In_853);
nor U872 (N_872,In_187,In_0);
nand U873 (N_873,In_341,In_287);
nor U874 (N_874,In_225,In_695);
or U875 (N_875,In_17,In_911);
and U876 (N_876,In_214,In_76);
or U877 (N_877,In_827,In_142);
nand U878 (N_878,In_513,In_510);
nand U879 (N_879,In_38,In_206);
nand U880 (N_880,In_705,In_984);
or U881 (N_881,In_226,In_345);
or U882 (N_882,In_734,In_646);
nand U883 (N_883,In_371,In_227);
nand U884 (N_884,In_777,In_865);
or U885 (N_885,In_725,In_608);
nand U886 (N_886,In_345,In_428);
nor U887 (N_887,In_371,In_530);
nand U888 (N_888,In_352,In_22);
or U889 (N_889,In_524,In_600);
and U890 (N_890,In_740,In_97);
and U891 (N_891,In_823,In_940);
nand U892 (N_892,In_559,In_479);
nor U893 (N_893,In_775,In_412);
or U894 (N_894,In_310,In_511);
or U895 (N_895,In_290,In_204);
and U896 (N_896,In_457,In_657);
nor U897 (N_897,In_994,In_93);
and U898 (N_898,In_395,In_838);
xnor U899 (N_899,In_938,In_217);
and U900 (N_900,In_419,In_557);
and U901 (N_901,In_59,In_610);
or U902 (N_902,In_328,In_629);
and U903 (N_903,In_258,In_935);
and U904 (N_904,In_929,In_990);
and U905 (N_905,In_352,In_39);
nand U906 (N_906,In_910,In_469);
nand U907 (N_907,In_729,In_776);
or U908 (N_908,In_220,In_79);
and U909 (N_909,In_250,In_908);
nor U910 (N_910,In_250,In_364);
nor U911 (N_911,In_558,In_801);
and U912 (N_912,In_984,In_870);
and U913 (N_913,In_463,In_462);
and U914 (N_914,In_987,In_762);
and U915 (N_915,In_332,In_541);
nor U916 (N_916,In_212,In_516);
and U917 (N_917,In_246,In_232);
or U918 (N_918,In_342,In_923);
and U919 (N_919,In_194,In_740);
or U920 (N_920,In_252,In_181);
or U921 (N_921,In_492,In_389);
or U922 (N_922,In_184,In_536);
or U923 (N_923,In_486,In_762);
nand U924 (N_924,In_399,In_902);
or U925 (N_925,In_417,In_994);
nor U926 (N_926,In_514,In_502);
or U927 (N_927,In_196,In_524);
and U928 (N_928,In_820,In_12);
and U929 (N_929,In_37,In_323);
nand U930 (N_930,In_9,In_978);
nor U931 (N_931,In_543,In_869);
and U932 (N_932,In_622,In_733);
nand U933 (N_933,In_829,In_432);
and U934 (N_934,In_819,In_163);
nor U935 (N_935,In_450,In_918);
or U936 (N_936,In_319,In_958);
nor U937 (N_937,In_657,In_827);
nor U938 (N_938,In_750,In_179);
or U939 (N_939,In_743,In_754);
and U940 (N_940,In_566,In_716);
xor U941 (N_941,In_897,In_644);
nor U942 (N_942,In_22,In_892);
or U943 (N_943,In_565,In_428);
or U944 (N_944,In_546,In_422);
nand U945 (N_945,In_402,In_739);
and U946 (N_946,In_492,In_196);
nand U947 (N_947,In_690,In_746);
and U948 (N_948,In_737,In_425);
nand U949 (N_949,In_662,In_280);
nor U950 (N_950,In_745,In_923);
or U951 (N_951,In_936,In_899);
nor U952 (N_952,In_257,In_866);
and U953 (N_953,In_764,In_456);
or U954 (N_954,In_232,In_935);
and U955 (N_955,In_320,In_561);
or U956 (N_956,In_455,In_482);
or U957 (N_957,In_295,In_238);
or U958 (N_958,In_787,In_157);
nor U959 (N_959,In_892,In_881);
and U960 (N_960,In_739,In_745);
or U961 (N_961,In_364,In_232);
nor U962 (N_962,In_877,In_670);
or U963 (N_963,In_96,In_455);
nor U964 (N_964,In_239,In_685);
nor U965 (N_965,In_902,In_136);
and U966 (N_966,In_461,In_235);
or U967 (N_967,In_306,In_471);
or U968 (N_968,In_146,In_990);
and U969 (N_969,In_500,In_667);
or U970 (N_970,In_323,In_69);
and U971 (N_971,In_788,In_235);
nor U972 (N_972,In_25,In_952);
nor U973 (N_973,In_925,In_85);
or U974 (N_974,In_50,In_486);
xor U975 (N_975,In_867,In_976);
and U976 (N_976,In_793,In_105);
nand U977 (N_977,In_44,In_963);
or U978 (N_978,In_510,In_431);
and U979 (N_979,In_231,In_464);
nand U980 (N_980,In_711,In_934);
nor U981 (N_981,In_161,In_972);
or U982 (N_982,In_88,In_45);
and U983 (N_983,In_418,In_647);
and U984 (N_984,In_274,In_622);
or U985 (N_985,In_44,In_148);
and U986 (N_986,In_694,In_742);
or U987 (N_987,In_959,In_584);
nand U988 (N_988,In_662,In_94);
nor U989 (N_989,In_124,In_55);
or U990 (N_990,In_263,In_130);
nor U991 (N_991,In_679,In_809);
xnor U992 (N_992,In_25,In_639);
nand U993 (N_993,In_397,In_644);
or U994 (N_994,In_246,In_383);
nand U995 (N_995,In_271,In_415);
nor U996 (N_996,In_409,In_925);
nor U997 (N_997,In_612,In_970);
nand U998 (N_998,In_474,In_858);
or U999 (N_999,In_392,In_741);
nor U1000 (N_1000,In_831,In_943);
nand U1001 (N_1001,In_512,In_772);
or U1002 (N_1002,In_2,In_83);
or U1003 (N_1003,In_470,In_790);
or U1004 (N_1004,In_474,In_47);
xor U1005 (N_1005,In_109,In_865);
and U1006 (N_1006,In_648,In_690);
and U1007 (N_1007,In_996,In_341);
nand U1008 (N_1008,In_135,In_652);
and U1009 (N_1009,In_107,In_694);
or U1010 (N_1010,In_807,In_196);
xor U1011 (N_1011,In_481,In_26);
nand U1012 (N_1012,In_753,In_424);
nor U1013 (N_1013,In_843,In_25);
nand U1014 (N_1014,In_440,In_243);
nor U1015 (N_1015,In_495,In_521);
nor U1016 (N_1016,In_413,In_785);
or U1017 (N_1017,In_19,In_742);
xnor U1018 (N_1018,In_757,In_254);
or U1019 (N_1019,In_833,In_573);
nand U1020 (N_1020,In_328,In_151);
nand U1021 (N_1021,In_711,In_429);
nand U1022 (N_1022,In_362,In_109);
or U1023 (N_1023,In_917,In_592);
nand U1024 (N_1024,In_397,In_505);
or U1025 (N_1025,In_650,In_59);
nor U1026 (N_1026,In_402,In_109);
or U1027 (N_1027,In_572,In_200);
nor U1028 (N_1028,In_129,In_545);
or U1029 (N_1029,In_370,In_117);
or U1030 (N_1030,In_460,In_548);
and U1031 (N_1031,In_638,In_943);
or U1032 (N_1032,In_439,In_275);
and U1033 (N_1033,In_838,In_719);
nor U1034 (N_1034,In_213,In_598);
nand U1035 (N_1035,In_529,In_988);
nor U1036 (N_1036,In_220,In_216);
nor U1037 (N_1037,In_688,In_3);
nor U1038 (N_1038,In_754,In_106);
and U1039 (N_1039,In_6,In_614);
nand U1040 (N_1040,In_510,In_212);
nand U1041 (N_1041,In_263,In_937);
nor U1042 (N_1042,In_259,In_757);
nand U1043 (N_1043,In_734,In_48);
nand U1044 (N_1044,In_472,In_439);
or U1045 (N_1045,In_164,In_700);
nand U1046 (N_1046,In_873,In_722);
nor U1047 (N_1047,In_236,In_256);
nor U1048 (N_1048,In_891,In_619);
or U1049 (N_1049,In_971,In_336);
nor U1050 (N_1050,In_27,In_922);
nand U1051 (N_1051,In_415,In_529);
nand U1052 (N_1052,In_393,In_595);
and U1053 (N_1053,In_206,In_647);
and U1054 (N_1054,In_851,In_240);
nand U1055 (N_1055,In_202,In_382);
or U1056 (N_1056,In_764,In_280);
and U1057 (N_1057,In_25,In_995);
nand U1058 (N_1058,In_522,In_674);
and U1059 (N_1059,In_795,In_599);
xor U1060 (N_1060,In_902,In_647);
and U1061 (N_1061,In_454,In_315);
nand U1062 (N_1062,In_863,In_884);
and U1063 (N_1063,In_18,In_118);
nor U1064 (N_1064,In_955,In_786);
nand U1065 (N_1065,In_560,In_803);
and U1066 (N_1066,In_78,In_834);
nor U1067 (N_1067,In_93,In_789);
nor U1068 (N_1068,In_540,In_504);
or U1069 (N_1069,In_361,In_350);
nor U1070 (N_1070,In_830,In_49);
and U1071 (N_1071,In_702,In_599);
or U1072 (N_1072,In_194,In_989);
nand U1073 (N_1073,In_300,In_307);
nand U1074 (N_1074,In_165,In_22);
nor U1075 (N_1075,In_177,In_856);
and U1076 (N_1076,In_250,In_196);
nor U1077 (N_1077,In_703,In_571);
nand U1078 (N_1078,In_461,In_367);
nand U1079 (N_1079,In_323,In_382);
or U1080 (N_1080,In_365,In_593);
nand U1081 (N_1081,In_24,In_40);
and U1082 (N_1082,In_18,In_556);
nor U1083 (N_1083,In_368,In_657);
nand U1084 (N_1084,In_239,In_302);
and U1085 (N_1085,In_888,In_618);
and U1086 (N_1086,In_213,In_303);
or U1087 (N_1087,In_873,In_225);
nand U1088 (N_1088,In_994,In_684);
and U1089 (N_1089,In_202,In_297);
nand U1090 (N_1090,In_537,In_532);
or U1091 (N_1091,In_794,In_626);
nand U1092 (N_1092,In_895,In_855);
and U1093 (N_1093,In_957,In_718);
xor U1094 (N_1094,In_9,In_860);
nand U1095 (N_1095,In_72,In_358);
nor U1096 (N_1096,In_702,In_175);
nand U1097 (N_1097,In_237,In_930);
or U1098 (N_1098,In_783,In_850);
nand U1099 (N_1099,In_317,In_24);
or U1100 (N_1100,In_228,In_171);
and U1101 (N_1101,In_895,In_702);
nand U1102 (N_1102,In_876,In_854);
nor U1103 (N_1103,In_442,In_78);
or U1104 (N_1104,In_310,In_468);
and U1105 (N_1105,In_891,In_562);
nor U1106 (N_1106,In_246,In_982);
nor U1107 (N_1107,In_851,In_393);
nor U1108 (N_1108,In_703,In_501);
nand U1109 (N_1109,In_765,In_826);
nor U1110 (N_1110,In_699,In_489);
nor U1111 (N_1111,In_346,In_542);
and U1112 (N_1112,In_185,In_354);
nand U1113 (N_1113,In_909,In_975);
or U1114 (N_1114,In_618,In_763);
or U1115 (N_1115,In_562,In_914);
nor U1116 (N_1116,In_268,In_233);
nand U1117 (N_1117,In_654,In_705);
nand U1118 (N_1118,In_495,In_800);
nor U1119 (N_1119,In_19,In_285);
nand U1120 (N_1120,In_238,In_294);
and U1121 (N_1121,In_250,In_228);
xor U1122 (N_1122,In_436,In_326);
and U1123 (N_1123,In_312,In_542);
or U1124 (N_1124,In_311,In_867);
nor U1125 (N_1125,In_718,In_412);
nand U1126 (N_1126,In_529,In_427);
nand U1127 (N_1127,In_928,In_731);
and U1128 (N_1128,In_504,In_471);
or U1129 (N_1129,In_147,In_760);
nor U1130 (N_1130,In_449,In_414);
and U1131 (N_1131,In_592,In_978);
nand U1132 (N_1132,In_152,In_106);
and U1133 (N_1133,In_621,In_842);
or U1134 (N_1134,In_365,In_845);
nor U1135 (N_1135,In_53,In_433);
and U1136 (N_1136,In_686,In_130);
xor U1137 (N_1137,In_99,In_34);
nand U1138 (N_1138,In_344,In_79);
and U1139 (N_1139,In_852,In_782);
nor U1140 (N_1140,In_182,In_126);
nor U1141 (N_1141,In_837,In_638);
nand U1142 (N_1142,In_502,In_880);
nor U1143 (N_1143,In_700,In_814);
and U1144 (N_1144,In_228,In_522);
and U1145 (N_1145,In_307,In_580);
nand U1146 (N_1146,In_25,In_679);
nand U1147 (N_1147,In_100,In_298);
and U1148 (N_1148,In_139,In_674);
or U1149 (N_1149,In_174,In_507);
or U1150 (N_1150,In_388,In_428);
or U1151 (N_1151,In_830,In_328);
nor U1152 (N_1152,In_811,In_780);
and U1153 (N_1153,In_843,In_620);
and U1154 (N_1154,In_746,In_862);
or U1155 (N_1155,In_327,In_301);
and U1156 (N_1156,In_414,In_795);
and U1157 (N_1157,In_388,In_872);
or U1158 (N_1158,In_100,In_74);
nand U1159 (N_1159,In_293,In_496);
xnor U1160 (N_1160,In_51,In_230);
or U1161 (N_1161,In_403,In_731);
nor U1162 (N_1162,In_310,In_669);
or U1163 (N_1163,In_236,In_698);
or U1164 (N_1164,In_871,In_472);
or U1165 (N_1165,In_826,In_687);
or U1166 (N_1166,In_593,In_374);
nand U1167 (N_1167,In_722,In_831);
nor U1168 (N_1168,In_417,In_501);
and U1169 (N_1169,In_266,In_183);
or U1170 (N_1170,In_494,In_999);
nand U1171 (N_1171,In_928,In_940);
nand U1172 (N_1172,In_620,In_517);
nand U1173 (N_1173,In_669,In_634);
and U1174 (N_1174,In_733,In_771);
and U1175 (N_1175,In_980,In_468);
nand U1176 (N_1176,In_412,In_282);
or U1177 (N_1177,In_353,In_280);
nor U1178 (N_1178,In_965,In_780);
nor U1179 (N_1179,In_934,In_116);
nand U1180 (N_1180,In_317,In_629);
nor U1181 (N_1181,In_462,In_52);
or U1182 (N_1182,In_311,In_403);
and U1183 (N_1183,In_38,In_988);
or U1184 (N_1184,In_809,In_608);
nor U1185 (N_1185,In_6,In_952);
and U1186 (N_1186,In_429,In_778);
nor U1187 (N_1187,In_906,In_162);
and U1188 (N_1188,In_996,In_958);
nand U1189 (N_1189,In_248,In_978);
nor U1190 (N_1190,In_620,In_636);
and U1191 (N_1191,In_266,In_862);
or U1192 (N_1192,In_375,In_466);
nand U1193 (N_1193,In_107,In_545);
or U1194 (N_1194,In_433,In_811);
and U1195 (N_1195,In_63,In_628);
nor U1196 (N_1196,In_92,In_789);
and U1197 (N_1197,In_290,In_604);
nand U1198 (N_1198,In_10,In_301);
nor U1199 (N_1199,In_218,In_198);
nand U1200 (N_1200,In_721,In_35);
nand U1201 (N_1201,In_305,In_903);
nand U1202 (N_1202,In_979,In_282);
xnor U1203 (N_1203,In_429,In_57);
and U1204 (N_1204,In_667,In_711);
or U1205 (N_1205,In_857,In_841);
xor U1206 (N_1206,In_103,In_31);
nand U1207 (N_1207,In_41,In_170);
and U1208 (N_1208,In_571,In_393);
or U1209 (N_1209,In_161,In_734);
or U1210 (N_1210,In_786,In_529);
xor U1211 (N_1211,In_689,In_802);
and U1212 (N_1212,In_483,In_631);
and U1213 (N_1213,In_965,In_637);
nand U1214 (N_1214,In_92,In_108);
nor U1215 (N_1215,In_319,In_47);
and U1216 (N_1216,In_80,In_432);
or U1217 (N_1217,In_385,In_579);
or U1218 (N_1218,In_525,In_478);
nor U1219 (N_1219,In_747,In_162);
nand U1220 (N_1220,In_233,In_770);
nor U1221 (N_1221,In_957,In_970);
xor U1222 (N_1222,In_109,In_278);
and U1223 (N_1223,In_978,In_608);
and U1224 (N_1224,In_335,In_537);
nor U1225 (N_1225,In_945,In_345);
xor U1226 (N_1226,In_770,In_329);
or U1227 (N_1227,In_172,In_501);
nand U1228 (N_1228,In_956,In_625);
nor U1229 (N_1229,In_260,In_133);
nand U1230 (N_1230,In_421,In_626);
and U1231 (N_1231,In_481,In_564);
nand U1232 (N_1232,In_653,In_721);
nor U1233 (N_1233,In_432,In_783);
nor U1234 (N_1234,In_863,In_48);
nand U1235 (N_1235,In_517,In_2);
nor U1236 (N_1236,In_924,In_499);
or U1237 (N_1237,In_144,In_965);
or U1238 (N_1238,In_542,In_263);
nor U1239 (N_1239,In_871,In_123);
nor U1240 (N_1240,In_195,In_65);
nand U1241 (N_1241,In_673,In_778);
nand U1242 (N_1242,In_336,In_347);
nor U1243 (N_1243,In_733,In_331);
or U1244 (N_1244,In_712,In_360);
or U1245 (N_1245,In_501,In_240);
nor U1246 (N_1246,In_75,In_199);
and U1247 (N_1247,In_250,In_419);
or U1248 (N_1248,In_716,In_782);
or U1249 (N_1249,In_503,In_485);
nor U1250 (N_1250,In_825,In_409);
and U1251 (N_1251,In_418,In_79);
and U1252 (N_1252,In_813,In_45);
and U1253 (N_1253,In_154,In_103);
nand U1254 (N_1254,In_237,In_831);
and U1255 (N_1255,In_989,In_632);
or U1256 (N_1256,In_441,In_862);
or U1257 (N_1257,In_152,In_94);
nand U1258 (N_1258,In_653,In_368);
nand U1259 (N_1259,In_992,In_756);
nor U1260 (N_1260,In_107,In_46);
nor U1261 (N_1261,In_401,In_319);
nand U1262 (N_1262,In_182,In_684);
nand U1263 (N_1263,In_729,In_815);
nand U1264 (N_1264,In_467,In_572);
or U1265 (N_1265,In_221,In_12);
and U1266 (N_1266,In_279,In_774);
nand U1267 (N_1267,In_731,In_832);
nor U1268 (N_1268,In_179,In_969);
nor U1269 (N_1269,In_728,In_472);
nand U1270 (N_1270,In_620,In_696);
and U1271 (N_1271,In_535,In_116);
nand U1272 (N_1272,In_796,In_594);
and U1273 (N_1273,In_672,In_860);
or U1274 (N_1274,In_114,In_667);
or U1275 (N_1275,In_482,In_401);
or U1276 (N_1276,In_847,In_986);
nor U1277 (N_1277,In_552,In_160);
or U1278 (N_1278,In_772,In_733);
and U1279 (N_1279,In_788,In_297);
nand U1280 (N_1280,In_545,In_412);
nand U1281 (N_1281,In_352,In_497);
nand U1282 (N_1282,In_63,In_821);
nand U1283 (N_1283,In_240,In_352);
nand U1284 (N_1284,In_716,In_290);
nor U1285 (N_1285,In_931,In_341);
nand U1286 (N_1286,In_566,In_940);
or U1287 (N_1287,In_718,In_660);
nand U1288 (N_1288,In_348,In_629);
or U1289 (N_1289,In_464,In_855);
nor U1290 (N_1290,In_240,In_536);
nor U1291 (N_1291,In_982,In_255);
and U1292 (N_1292,In_174,In_512);
and U1293 (N_1293,In_557,In_599);
xnor U1294 (N_1294,In_745,In_197);
nand U1295 (N_1295,In_858,In_749);
and U1296 (N_1296,In_67,In_383);
nand U1297 (N_1297,In_650,In_872);
or U1298 (N_1298,In_245,In_179);
or U1299 (N_1299,In_793,In_230);
nand U1300 (N_1300,In_460,In_758);
or U1301 (N_1301,In_13,In_491);
or U1302 (N_1302,In_81,In_713);
nor U1303 (N_1303,In_128,In_922);
and U1304 (N_1304,In_383,In_430);
nor U1305 (N_1305,In_505,In_307);
nor U1306 (N_1306,In_204,In_294);
nor U1307 (N_1307,In_955,In_122);
or U1308 (N_1308,In_1,In_158);
nor U1309 (N_1309,In_811,In_898);
nand U1310 (N_1310,In_556,In_85);
xor U1311 (N_1311,In_526,In_12);
nand U1312 (N_1312,In_105,In_413);
nand U1313 (N_1313,In_239,In_348);
nand U1314 (N_1314,In_26,In_928);
nor U1315 (N_1315,In_497,In_303);
nand U1316 (N_1316,In_465,In_882);
nand U1317 (N_1317,In_608,In_643);
nor U1318 (N_1318,In_963,In_947);
nand U1319 (N_1319,In_838,In_403);
nor U1320 (N_1320,In_971,In_20);
nor U1321 (N_1321,In_92,In_812);
nor U1322 (N_1322,In_722,In_788);
xor U1323 (N_1323,In_914,In_328);
nand U1324 (N_1324,In_683,In_296);
nor U1325 (N_1325,In_484,In_385);
or U1326 (N_1326,In_666,In_869);
nand U1327 (N_1327,In_660,In_192);
or U1328 (N_1328,In_31,In_303);
nor U1329 (N_1329,In_218,In_843);
nor U1330 (N_1330,In_304,In_513);
or U1331 (N_1331,In_173,In_63);
or U1332 (N_1332,In_881,In_811);
nand U1333 (N_1333,In_488,In_143);
nand U1334 (N_1334,In_611,In_255);
nor U1335 (N_1335,In_973,In_98);
and U1336 (N_1336,In_735,In_515);
nor U1337 (N_1337,In_637,In_805);
nor U1338 (N_1338,In_101,In_329);
nor U1339 (N_1339,In_780,In_3);
nand U1340 (N_1340,In_210,In_672);
or U1341 (N_1341,In_197,In_171);
and U1342 (N_1342,In_254,In_46);
or U1343 (N_1343,In_963,In_365);
nor U1344 (N_1344,In_656,In_16);
nor U1345 (N_1345,In_984,In_652);
and U1346 (N_1346,In_908,In_678);
and U1347 (N_1347,In_184,In_992);
and U1348 (N_1348,In_349,In_414);
xnor U1349 (N_1349,In_32,In_163);
nand U1350 (N_1350,In_295,In_925);
nand U1351 (N_1351,In_527,In_774);
or U1352 (N_1352,In_791,In_206);
or U1353 (N_1353,In_623,In_27);
or U1354 (N_1354,In_128,In_360);
or U1355 (N_1355,In_288,In_369);
or U1356 (N_1356,In_600,In_672);
nand U1357 (N_1357,In_566,In_443);
or U1358 (N_1358,In_614,In_768);
and U1359 (N_1359,In_144,In_924);
or U1360 (N_1360,In_951,In_274);
or U1361 (N_1361,In_646,In_476);
nor U1362 (N_1362,In_17,In_77);
nor U1363 (N_1363,In_339,In_750);
nand U1364 (N_1364,In_326,In_248);
and U1365 (N_1365,In_659,In_226);
nor U1366 (N_1366,In_368,In_626);
and U1367 (N_1367,In_875,In_331);
and U1368 (N_1368,In_342,In_670);
nand U1369 (N_1369,In_617,In_805);
nor U1370 (N_1370,In_320,In_97);
and U1371 (N_1371,In_185,In_109);
and U1372 (N_1372,In_261,In_616);
xnor U1373 (N_1373,In_600,In_282);
or U1374 (N_1374,In_100,In_431);
and U1375 (N_1375,In_138,In_923);
nor U1376 (N_1376,In_991,In_834);
nand U1377 (N_1377,In_144,In_816);
nand U1378 (N_1378,In_352,In_650);
nand U1379 (N_1379,In_590,In_908);
or U1380 (N_1380,In_850,In_223);
and U1381 (N_1381,In_725,In_283);
or U1382 (N_1382,In_303,In_460);
nand U1383 (N_1383,In_314,In_722);
nand U1384 (N_1384,In_747,In_198);
and U1385 (N_1385,In_458,In_209);
and U1386 (N_1386,In_4,In_330);
or U1387 (N_1387,In_42,In_943);
or U1388 (N_1388,In_299,In_607);
nor U1389 (N_1389,In_839,In_921);
xnor U1390 (N_1390,In_804,In_726);
or U1391 (N_1391,In_864,In_2);
and U1392 (N_1392,In_840,In_980);
or U1393 (N_1393,In_114,In_678);
nor U1394 (N_1394,In_412,In_698);
xnor U1395 (N_1395,In_532,In_80);
or U1396 (N_1396,In_684,In_191);
nor U1397 (N_1397,In_819,In_48);
nand U1398 (N_1398,In_122,In_564);
nor U1399 (N_1399,In_67,In_574);
nand U1400 (N_1400,In_675,In_543);
and U1401 (N_1401,In_12,In_798);
nor U1402 (N_1402,In_395,In_942);
nand U1403 (N_1403,In_724,In_279);
nor U1404 (N_1404,In_227,In_483);
and U1405 (N_1405,In_375,In_103);
and U1406 (N_1406,In_329,In_599);
and U1407 (N_1407,In_196,In_661);
or U1408 (N_1408,In_544,In_484);
xnor U1409 (N_1409,In_766,In_88);
and U1410 (N_1410,In_490,In_354);
or U1411 (N_1411,In_195,In_45);
nand U1412 (N_1412,In_93,In_434);
and U1413 (N_1413,In_634,In_800);
or U1414 (N_1414,In_90,In_113);
or U1415 (N_1415,In_818,In_266);
or U1416 (N_1416,In_540,In_588);
or U1417 (N_1417,In_41,In_807);
nor U1418 (N_1418,In_459,In_72);
nand U1419 (N_1419,In_318,In_495);
and U1420 (N_1420,In_832,In_759);
nor U1421 (N_1421,In_342,In_114);
or U1422 (N_1422,In_850,In_784);
nand U1423 (N_1423,In_715,In_292);
nor U1424 (N_1424,In_248,In_132);
nand U1425 (N_1425,In_402,In_431);
or U1426 (N_1426,In_79,In_560);
and U1427 (N_1427,In_984,In_401);
or U1428 (N_1428,In_24,In_874);
or U1429 (N_1429,In_569,In_797);
nor U1430 (N_1430,In_852,In_349);
nor U1431 (N_1431,In_437,In_616);
and U1432 (N_1432,In_200,In_353);
nand U1433 (N_1433,In_487,In_720);
or U1434 (N_1434,In_271,In_790);
nor U1435 (N_1435,In_668,In_60);
nor U1436 (N_1436,In_200,In_611);
nand U1437 (N_1437,In_899,In_967);
or U1438 (N_1438,In_730,In_656);
nand U1439 (N_1439,In_810,In_769);
nand U1440 (N_1440,In_465,In_996);
or U1441 (N_1441,In_964,In_541);
nor U1442 (N_1442,In_139,In_786);
nand U1443 (N_1443,In_634,In_351);
nor U1444 (N_1444,In_630,In_701);
nor U1445 (N_1445,In_301,In_828);
or U1446 (N_1446,In_368,In_231);
and U1447 (N_1447,In_470,In_172);
nand U1448 (N_1448,In_17,In_457);
and U1449 (N_1449,In_515,In_580);
or U1450 (N_1450,In_264,In_425);
and U1451 (N_1451,In_5,In_861);
nand U1452 (N_1452,In_992,In_692);
and U1453 (N_1453,In_655,In_708);
nor U1454 (N_1454,In_796,In_214);
and U1455 (N_1455,In_629,In_283);
nand U1456 (N_1456,In_84,In_121);
or U1457 (N_1457,In_369,In_723);
or U1458 (N_1458,In_447,In_928);
nand U1459 (N_1459,In_825,In_389);
nor U1460 (N_1460,In_207,In_49);
nor U1461 (N_1461,In_230,In_49);
nor U1462 (N_1462,In_913,In_345);
nand U1463 (N_1463,In_321,In_981);
or U1464 (N_1464,In_675,In_890);
and U1465 (N_1465,In_379,In_964);
or U1466 (N_1466,In_930,In_999);
nor U1467 (N_1467,In_671,In_113);
nand U1468 (N_1468,In_975,In_427);
nand U1469 (N_1469,In_12,In_351);
nor U1470 (N_1470,In_686,In_858);
nor U1471 (N_1471,In_977,In_449);
or U1472 (N_1472,In_295,In_119);
nor U1473 (N_1473,In_973,In_655);
or U1474 (N_1474,In_420,In_139);
nand U1475 (N_1475,In_797,In_481);
nor U1476 (N_1476,In_635,In_720);
xor U1477 (N_1477,In_849,In_294);
or U1478 (N_1478,In_551,In_833);
and U1479 (N_1479,In_654,In_237);
and U1480 (N_1480,In_818,In_151);
xnor U1481 (N_1481,In_63,In_512);
or U1482 (N_1482,In_56,In_828);
and U1483 (N_1483,In_790,In_223);
nand U1484 (N_1484,In_712,In_262);
or U1485 (N_1485,In_945,In_417);
or U1486 (N_1486,In_921,In_741);
or U1487 (N_1487,In_711,In_491);
nand U1488 (N_1488,In_42,In_306);
nor U1489 (N_1489,In_35,In_768);
and U1490 (N_1490,In_992,In_354);
nand U1491 (N_1491,In_782,In_762);
or U1492 (N_1492,In_910,In_173);
or U1493 (N_1493,In_671,In_546);
or U1494 (N_1494,In_33,In_804);
or U1495 (N_1495,In_858,In_783);
nor U1496 (N_1496,In_334,In_233);
or U1497 (N_1497,In_380,In_197);
nand U1498 (N_1498,In_524,In_695);
nor U1499 (N_1499,In_857,In_287);
nor U1500 (N_1500,In_217,In_845);
or U1501 (N_1501,In_681,In_654);
or U1502 (N_1502,In_148,In_0);
nor U1503 (N_1503,In_362,In_466);
nor U1504 (N_1504,In_911,In_546);
nand U1505 (N_1505,In_484,In_90);
and U1506 (N_1506,In_447,In_142);
nand U1507 (N_1507,In_435,In_149);
nand U1508 (N_1508,In_324,In_42);
and U1509 (N_1509,In_825,In_340);
and U1510 (N_1510,In_811,In_817);
xnor U1511 (N_1511,In_412,In_571);
nand U1512 (N_1512,In_306,In_624);
nand U1513 (N_1513,In_828,In_186);
or U1514 (N_1514,In_931,In_467);
or U1515 (N_1515,In_365,In_210);
or U1516 (N_1516,In_739,In_618);
and U1517 (N_1517,In_314,In_374);
or U1518 (N_1518,In_273,In_47);
or U1519 (N_1519,In_598,In_107);
or U1520 (N_1520,In_521,In_334);
and U1521 (N_1521,In_762,In_58);
and U1522 (N_1522,In_567,In_671);
nand U1523 (N_1523,In_651,In_269);
nand U1524 (N_1524,In_615,In_1);
nor U1525 (N_1525,In_264,In_506);
nand U1526 (N_1526,In_878,In_110);
nor U1527 (N_1527,In_634,In_54);
and U1528 (N_1528,In_20,In_19);
or U1529 (N_1529,In_343,In_349);
or U1530 (N_1530,In_241,In_688);
or U1531 (N_1531,In_123,In_463);
nor U1532 (N_1532,In_884,In_390);
xor U1533 (N_1533,In_311,In_124);
xnor U1534 (N_1534,In_933,In_577);
nor U1535 (N_1535,In_941,In_928);
or U1536 (N_1536,In_768,In_548);
or U1537 (N_1537,In_33,In_42);
and U1538 (N_1538,In_30,In_567);
or U1539 (N_1539,In_798,In_832);
nand U1540 (N_1540,In_109,In_172);
nand U1541 (N_1541,In_147,In_15);
and U1542 (N_1542,In_35,In_50);
nor U1543 (N_1543,In_940,In_777);
nor U1544 (N_1544,In_410,In_313);
or U1545 (N_1545,In_142,In_287);
nor U1546 (N_1546,In_447,In_110);
nor U1547 (N_1547,In_358,In_975);
or U1548 (N_1548,In_697,In_583);
nor U1549 (N_1549,In_35,In_739);
nor U1550 (N_1550,In_144,In_360);
and U1551 (N_1551,In_970,In_291);
nand U1552 (N_1552,In_266,In_460);
or U1553 (N_1553,In_241,In_163);
nor U1554 (N_1554,In_234,In_969);
or U1555 (N_1555,In_537,In_677);
nand U1556 (N_1556,In_344,In_608);
nor U1557 (N_1557,In_531,In_995);
nor U1558 (N_1558,In_986,In_934);
or U1559 (N_1559,In_406,In_678);
or U1560 (N_1560,In_132,In_876);
or U1561 (N_1561,In_47,In_836);
nand U1562 (N_1562,In_195,In_742);
or U1563 (N_1563,In_794,In_715);
or U1564 (N_1564,In_476,In_508);
and U1565 (N_1565,In_460,In_490);
nand U1566 (N_1566,In_883,In_114);
nand U1567 (N_1567,In_724,In_866);
nand U1568 (N_1568,In_203,In_316);
and U1569 (N_1569,In_975,In_828);
and U1570 (N_1570,In_681,In_678);
nand U1571 (N_1571,In_519,In_10);
nor U1572 (N_1572,In_605,In_603);
nor U1573 (N_1573,In_643,In_522);
xnor U1574 (N_1574,In_825,In_600);
nand U1575 (N_1575,In_133,In_880);
or U1576 (N_1576,In_696,In_469);
nor U1577 (N_1577,In_316,In_423);
nand U1578 (N_1578,In_377,In_721);
nor U1579 (N_1579,In_133,In_578);
xnor U1580 (N_1580,In_875,In_967);
xor U1581 (N_1581,In_242,In_532);
nor U1582 (N_1582,In_434,In_147);
or U1583 (N_1583,In_774,In_716);
nand U1584 (N_1584,In_169,In_350);
and U1585 (N_1585,In_388,In_517);
or U1586 (N_1586,In_384,In_10);
or U1587 (N_1587,In_828,In_240);
nand U1588 (N_1588,In_216,In_59);
and U1589 (N_1589,In_429,In_436);
or U1590 (N_1590,In_203,In_813);
or U1591 (N_1591,In_471,In_968);
nand U1592 (N_1592,In_762,In_667);
nor U1593 (N_1593,In_61,In_784);
or U1594 (N_1594,In_844,In_778);
and U1595 (N_1595,In_346,In_170);
or U1596 (N_1596,In_339,In_826);
nor U1597 (N_1597,In_160,In_322);
nand U1598 (N_1598,In_29,In_706);
nand U1599 (N_1599,In_169,In_75);
and U1600 (N_1600,In_652,In_902);
nor U1601 (N_1601,In_505,In_96);
nand U1602 (N_1602,In_879,In_956);
or U1603 (N_1603,In_319,In_356);
and U1604 (N_1604,In_631,In_107);
nor U1605 (N_1605,In_451,In_453);
nor U1606 (N_1606,In_507,In_751);
and U1607 (N_1607,In_85,In_134);
nor U1608 (N_1608,In_703,In_854);
or U1609 (N_1609,In_570,In_701);
nand U1610 (N_1610,In_563,In_837);
nor U1611 (N_1611,In_371,In_523);
nand U1612 (N_1612,In_936,In_254);
and U1613 (N_1613,In_692,In_385);
or U1614 (N_1614,In_979,In_980);
and U1615 (N_1615,In_615,In_982);
nand U1616 (N_1616,In_267,In_338);
and U1617 (N_1617,In_540,In_799);
and U1618 (N_1618,In_688,In_14);
nand U1619 (N_1619,In_226,In_772);
and U1620 (N_1620,In_847,In_641);
and U1621 (N_1621,In_347,In_504);
or U1622 (N_1622,In_301,In_921);
nor U1623 (N_1623,In_4,In_647);
or U1624 (N_1624,In_50,In_413);
and U1625 (N_1625,In_838,In_509);
nor U1626 (N_1626,In_688,In_102);
or U1627 (N_1627,In_575,In_855);
or U1628 (N_1628,In_80,In_111);
nand U1629 (N_1629,In_970,In_265);
or U1630 (N_1630,In_535,In_757);
nand U1631 (N_1631,In_182,In_375);
nand U1632 (N_1632,In_789,In_47);
or U1633 (N_1633,In_635,In_207);
and U1634 (N_1634,In_10,In_882);
or U1635 (N_1635,In_556,In_31);
nand U1636 (N_1636,In_409,In_986);
nand U1637 (N_1637,In_540,In_35);
or U1638 (N_1638,In_105,In_779);
or U1639 (N_1639,In_986,In_54);
nor U1640 (N_1640,In_127,In_556);
nor U1641 (N_1641,In_857,In_432);
and U1642 (N_1642,In_521,In_369);
nand U1643 (N_1643,In_140,In_67);
and U1644 (N_1644,In_376,In_442);
nor U1645 (N_1645,In_538,In_202);
nor U1646 (N_1646,In_105,In_797);
nor U1647 (N_1647,In_941,In_80);
nand U1648 (N_1648,In_905,In_521);
or U1649 (N_1649,In_567,In_413);
nor U1650 (N_1650,In_176,In_447);
or U1651 (N_1651,In_576,In_286);
and U1652 (N_1652,In_922,In_679);
nor U1653 (N_1653,In_723,In_808);
or U1654 (N_1654,In_259,In_514);
nor U1655 (N_1655,In_378,In_608);
or U1656 (N_1656,In_566,In_247);
nand U1657 (N_1657,In_467,In_914);
nand U1658 (N_1658,In_438,In_576);
nand U1659 (N_1659,In_75,In_884);
and U1660 (N_1660,In_105,In_61);
nand U1661 (N_1661,In_756,In_833);
nand U1662 (N_1662,In_213,In_471);
nand U1663 (N_1663,In_770,In_139);
nand U1664 (N_1664,In_556,In_869);
nand U1665 (N_1665,In_711,In_17);
or U1666 (N_1666,In_960,In_34);
or U1667 (N_1667,In_271,In_37);
nor U1668 (N_1668,In_932,In_564);
nor U1669 (N_1669,In_496,In_694);
xnor U1670 (N_1670,In_506,In_115);
nand U1671 (N_1671,In_974,In_497);
nand U1672 (N_1672,In_564,In_637);
nor U1673 (N_1673,In_567,In_122);
and U1674 (N_1674,In_69,In_263);
nor U1675 (N_1675,In_345,In_213);
or U1676 (N_1676,In_276,In_10);
or U1677 (N_1677,In_681,In_869);
and U1678 (N_1678,In_773,In_227);
or U1679 (N_1679,In_175,In_767);
xor U1680 (N_1680,In_49,In_180);
or U1681 (N_1681,In_986,In_80);
nand U1682 (N_1682,In_192,In_783);
nor U1683 (N_1683,In_219,In_64);
nor U1684 (N_1684,In_957,In_128);
or U1685 (N_1685,In_902,In_373);
nor U1686 (N_1686,In_779,In_480);
or U1687 (N_1687,In_283,In_665);
and U1688 (N_1688,In_63,In_703);
nand U1689 (N_1689,In_835,In_912);
nor U1690 (N_1690,In_977,In_476);
nor U1691 (N_1691,In_150,In_705);
or U1692 (N_1692,In_51,In_367);
or U1693 (N_1693,In_966,In_190);
or U1694 (N_1694,In_226,In_397);
nand U1695 (N_1695,In_33,In_152);
nand U1696 (N_1696,In_257,In_983);
nor U1697 (N_1697,In_728,In_249);
or U1698 (N_1698,In_991,In_855);
or U1699 (N_1699,In_58,In_490);
and U1700 (N_1700,In_903,In_298);
nand U1701 (N_1701,In_226,In_187);
nor U1702 (N_1702,In_762,In_950);
nand U1703 (N_1703,In_939,In_886);
nor U1704 (N_1704,In_720,In_90);
and U1705 (N_1705,In_301,In_575);
nor U1706 (N_1706,In_713,In_307);
nor U1707 (N_1707,In_179,In_996);
and U1708 (N_1708,In_551,In_627);
nand U1709 (N_1709,In_91,In_533);
nand U1710 (N_1710,In_541,In_707);
nor U1711 (N_1711,In_156,In_876);
and U1712 (N_1712,In_263,In_153);
nor U1713 (N_1713,In_223,In_749);
nand U1714 (N_1714,In_302,In_162);
nand U1715 (N_1715,In_768,In_914);
and U1716 (N_1716,In_182,In_518);
nor U1717 (N_1717,In_257,In_168);
nor U1718 (N_1718,In_238,In_248);
nor U1719 (N_1719,In_781,In_229);
nand U1720 (N_1720,In_823,In_62);
or U1721 (N_1721,In_602,In_232);
nand U1722 (N_1722,In_166,In_183);
nand U1723 (N_1723,In_603,In_954);
or U1724 (N_1724,In_576,In_862);
nand U1725 (N_1725,In_327,In_7);
and U1726 (N_1726,In_101,In_112);
and U1727 (N_1727,In_650,In_891);
nand U1728 (N_1728,In_186,In_407);
nand U1729 (N_1729,In_102,In_393);
nand U1730 (N_1730,In_123,In_927);
or U1731 (N_1731,In_840,In_194);
xnor U1732 (N_1732,In_117,In_802);
nand U1733 (N_1733,In_78,In_174);
nor U1734 (N_1734,In_272,In_817);
nand U1735 (N_1735,In_271,In_150);
nand U1736 (N_1736,In_238,In_662);
nand U1737 (N_1737,In_531,In_83);
and U1738 (N_1738,In_723,In_997);
nor U1739 (N_1739,In_317,In_111);
nor U1740 (N_1740,In_391,In_321);
or U1741 (N_1741,In_997,In_413);
and U1742 (N_1742,In_426,In_196);
or U1743 (N_1743,In_498,In_570);
and U1744 (N_1744,In_533,In_241);
or U1745 (N_1745,In_35,In_895);
nor U1746 (N_1746,In_178,In_915);
and U1747 (N_1747,In_665,In_403);
or U1748 (N_1748,In_803,In_593);
or U1749 (N_1749,In_418,In_945);
nand U1750 (N_1750,In_55,In_481);
or U1751 (N_1751,In_496,In_499);
and U1752 (N_1752,In_840,In_395);
nor U1753 (N_1753,In_556,In_644);
nand U1754 (N_1754,In_635,In_95);
and U1755 (N_1755,In_390,In_476);
nand U1756 (N_1756,In_990,In_931);
and U1757 (N_1757,In_726,In_592);
nor U1758 (N_1758,In_689,In_856);
xor U1759 (N_1759,In_365,In_788);
nand U1760 (N_1760,In_544,In_4);
or U1761 (N_1761,In_493,In_719);
and U1762 (N_1762,In_838,In_714);
and U1763 (N_1763,In_807,In_943);
nor U1764 (N_1764,In_378,In_610);
and U1765 (N_1765,In_896,In_20);
nand U1766 (N_1766,In_29,In_640);
and U1767 (N_1767,In_588,In_899);
nand U1768 (N_1768,In_959,In_495);
nor U1769 (N_1769,In_412,In_258);
nand U1770 (N_1770,In_41,In_189);
or U1771 (N_1771,In_979,In_295);
nand U1772 (N_1772,In_171,In_559);
nand U1773 (N_1773,In_864,In_770);
and U1774 (N_1774,In_257,In_212);
and U1775 (N_1775,In_511,In_555);
and U1776 (N_1776,In_241,In_424);
and U1777 (N_1777,In_631,In_92);
or U1778 (N_1778,In_246,In_33);
nor U1779 (N_1779,In_888,In_900);
nor U1780 (N_1780,In_182,In_381);
nand U1781 (N_1781,In_398,In_574);
nor U1782 (N_1782,In_781,In_244);
and U1783 (N_1783,In_131,In_400);
nor U1784 (N_1784,In_670,In_213);
nor U1785 (N_1785,In_535,In_912);
nand U1786 (N_1786,In_498,In_80);
or U1787 (N_1787,In_224,In_0);
or U1788 (N_1788,In_933,In_590);
and U1789 (N_1789,In_815,In_972);
nor U1790 (N_1790,In_453,In_830);
nor U1791 (N_1791,In_846,In_132);
and U1792 (N_1792,In_408,In_660);
nor U1793 (N_1793,In_555,In_664);
or U1794 (N_1794,In_638,In_324);
nor U1795 (N_1795,In_176,In_555);
nor U1796 (N_1796,In_2,In_903);
and U1797 (N_1797,In_708,In_680);
nand U1798 (N_1798,In_211,In_120);
and U1799 (N_1799,In_198,In_898);
and U1800 (N_1800,In_412,In_272);
and U1801 (N_1801,In_593,In_540);
nor U1802 (N_1802,In_137,In_975);
or U1803 (N_1803,In_530,In_257);
nand U1804 (N_1804,In_906,In_144);
nand U1805 (N_1805,In_603,In_115);
nor U1806 (N_1806,In_697,In_896);
or U1807 (N_1807,In_588,In_431);
and U1808 (N_1808,In_400,In_759);
nand U1809 (N_1809,In_756,In_247);
nor U1810 (N_1810,In_186,In_664);
nand U1811 (N_1811,In_549,In_49);
nand U1812 (N_1812,In_276,In_315);
nand U1813 (N_1813,In_534,In_360);
xnor U1814 (N_1814,In_122,In_408);
or U1815 (N_1815,In_350,In_686);
or U1816 (N_1816,In_164,In_939);
and U1817 (N_1817,In_404,In_93);
nand U1818 (N_1818,In_300,In_36);
nor U1819 (N_1819,In_863,In_718);
and U1820 (N_1820,In_378,In_609);
nand U1821 (N_1821,In_869,In_359);
nand U1822 (N_1822,In_200,In_713);
nand U1823 (N_1823,In_755,In_671);
nand U1824 (N_1824,In_168,In_932);
and U1825 (N_1825,In_525,In_996);
nand U1826 (N_1826,In_992,In_590);
nor U1827 (N_1827,In_509,In_444);
nor U1828 (N_1828,In_821,In_205);
nand U1829 (N_1829,In_529,In_587);
and U1830 (N_1830,In_419,In_223);
and U1831 (N_1831,In_154,In_236);
and U1832 (N_1832,In_705,In_185);
nor U1833 (N_1833,In_371,In_239);
and U1834 (N_1834,In_285,In_535);
and U1835 (N_1835,In_147,In_161);
nand U1836 (N_1836,In_626,In_496);
and U1837 (N_1837,In_69,In_89);
xor U1838 (N_1838,In_542,In_808);
nand U1839 (N_1839,In_516,In_280);
and U1840 (N_1840,In_766,In_810);
or U1841 (N_1841,In_6,In_166);
nor U1842 (N_1842,In_233,In_401);
nor U1843 (N_1843,In_279,In_602);
or U1844 (N_1844,In_973,In_111);
nor U1845 (N_1845,In_980,In_419);
and U1846 (N_1846,In_527,In_659);
and U1847 (N_1847,In_669,In_247);
and U1848 (N_1848,In_336,In_527);
xor U1849 (N_1849,In_72,In_670);
xnor U1850 (N_1850,In_418,In_841);
nor U1851 (N_1851,In_720,In_415);
nor U1852 (N_1852,In_439,In_868);
and U1853 (N_1853,In_60,In_56);
nand U1854 (N_1854,In_776,In_349);
or U1855 (N_1855,In_989,In_469);
or U1856 (N_1856,In_872,In_9);
and U1857 (N_1857,In_353,In_21);
nor U1858 (N_1858,In_692,In_518);
nand U1859 (N_1859,In_139,In_390);
nor U1860 (N_1860,In_350,In_489);
nand U1861 (N_1861,In_399,In_281);
or U1862 (N_1862,In_189,In_857);
and U1863 (N_1863,In_889,In_243);
nor U1864 (N_1864,In_17,In_758);
and U1865 (N_1865,In_505,In_682);
nand U1866 (N_1866,In_833,In_562);
or U1867 (N_1867,In_688,In_50);
or U1868 (N_1868,In_143,In_195);
xnor U1869 (N_1869,In_703,In_169);
nor U1870 (N_1870,In_367,In_393);
nand U1871 (N_1871,In_162,In_88);
or U1872 (N_1872,In_136,In_864);
nor U1873 (N_1873,In_957,In_355);
or U1874 (N_1874,In_987,In_709);
or U1875 (N_1875,In_481,In_590);
and U1876 (N_1876,In_908,In_492);
and U1877 (N_1877,In_0,In_100);
or U1878 (N_1878,In_484,In_554);
nor U1879 (N_1879,In_389,In_577);
and U1880 (N_1880,In_369,In_201);
nor U1881 (N_1881,In_321,In_75);
or U1882 (N_1882,In_79,In_189);
or U1883 (N_1883,In_580,In_149);
nor U1884 (N_1884,In_318,In_657);
and U1885 (N_1885,In_734,In_43);
nand U1886 (N_1886,In_801,In_986);
nor U1887 (N_1887,In_821,In_192);
nand U1888 (N_1888,In_929,In_19);
and U1889 (N_1889,In_280,In_315);
nor U1890 (N_1890,In_178,In_196);
and U1891 (N_1891,In_475,In_23);
or U1892 (N_1892,In_668,In_392);
or U1893 (N_1893,In_258,In_430);
nand U1894 (N_1894,In_856,In_365);
nor U1895 (N_1895,In_402,In_383);
or U1896 (N_1896,In_887,In_38);
and U1897 (N_1897,In_324,In_232);
and U1898 (N_1898,In_286,In_738);
nand U1899 (N_1899,In_240,In_91);
nor U1900 (N_1900,In_449,In_323);
or U1901 (N_1901,In_509,In_642);
nor U1902 (N_1902,In_818,In_142);
and U1903 (N_1903,In_500,In_856);
and U1904 (N_1904,In_540,In_70);
xor U1905 (N_1905,In_50,In_91);
and U1906 (N_1906,In_562,In_264);
nand U1907 (N_1907,In_470,In_528);
nor U1908 (N_1908,In_65,In_467);
or U1909 (N_1909,In_659,In_986);
nand U1910 (N_1910,In_973,In_651);
and U1911 (N_1911,In_563,In_374);
nand U1912 (N_1912,In_377,In_320);
xnor U1913 (N_1913,In_697,In_597);
and U1914 (N_1914,In_636,In_600);
nor U1915 (N_1915,In_976,In_231);
nand U1916 (N_1916,In_270,In_90);
nor U1917 (N_1917,In_765,In_5);
or U1918 (N_1918,In_218,In_96);
nand U1919 (N_1919,In_51,In_818);
and U1920 (N_1920,In_136,In_114);
or U1921 (N_1921,In_161,In_263);
nand U1922 (N_1922,In_992,In_31);
or U1923 (N_1923,In_302,In_187);
nand U1924 (N_1924,In_841,In_665);
and U1925 (N_1925,In_51,In_69);
nand U1926 (N_1926,In_726,In_969);
nand U1927 (N_1927,In_329,In_449);
nand U1928 (N_1928,In_358,In_882);
nand U1929 (N_1929,In_453,In_643);
or U1930 (N_1930,In_791,In_938);
and U1931 (N_1931,In_491,In_293);
and U1932 (N_1932,In_384,In_848);
or U1933 (N_1933,In_266,In_857);
or U1934 (N_1934,In_156,In_122);
nand U1935 (N_1935,In_54,In_224);
or U1936 (N_1936,In_649,In_90);
and U1937 (N_1937,In_531,In_372);
nand U1938 (N_1938,In_467,In_543);
and U1939 (N_1939,In_925,In_886);
or U1940 (N_1940,In_107,In_683);
xnor U1941 (N_1941,In_676,In_917);
or U1942 (N_1942,In_694,In_187);
or U1943 (N_1943,In_923,In_997);
nand U1944 (N_1944,In_882,In_402);
nor U1945 (N_1945,In_877,In_454);
or U1946 (N_1946,In_937,In_70);
or U1947 (N_1947,In_217,In_805);
nor U1948 (N_1948,In_688,In_332);
and U1949 (N_1949,In_242,In_380);
and U1950 (N_1950,In_622,In_917);
and U1951 (N_1951,In_889,In_152);
nor U1952 (N_1952,In_987,In_339);
nor U1953 (N_1953,In_448,In_251);
nor U1954 (N_1954,In_4,In_801);
and U1955 (N_1955,In_669,In_864);
or U1956 (N_1956,In_682,In_129);
nor U1957 (N_1957,In_895,In_265);
nand U1958 (N_1958,In_136,In_488);
nor U1959 (N_1959,In_343,In_80);
nor U1960 (N_1960,In_824,In_0);
xor U1961 (N_1961,In_483,In_343);
nand U1962 (N_1962,In_712,In_417);
nor U1963 (N_1963,In_52,In_360);
or U1964 (N_1964,In_468,In_485);
nand U1965 (N_1965,In_542,In_167);
and U1966 (N_1966,In_514,In_865);
and U1967 (N_1967,In_793,In_400);
and U1968 (N_1968,In_826,In_34);
nor U1969 (N_1969,In_789,In_660);
and U1970 (N_1970,In_492,In_565);
or U1971 (N_1971,In_309,In_457);
or U1972 (N_1972,In_492,In_479);
nor U1973 (N_1973,In_750,In_266);
or U1974 (N_1974,In_13,In_372);
nor U1975 (N_1975,In_223,In_500);
xnor U1976 (N_1976,In_495,In_803);
and U1977 (N_1977,In_659,In_128);
or U1978 (N_1978,In_482,In_741);
or U1979 (N_1979,In_650,In_484);
nor U1980 (N_1980,In_876,In_46);
or U1981 (N_1981,In_212,In_514);
or U1982 (N_1982,In_483,In_642);
nand U1983 (N_1983,In_275,In_390);
nand U1984 (N_1984,In_453,In_329);
nor U1985 (N_1985,In_140,In_201);
xnor U1986 (N_1986,In_13,In_79);
xor U1987 (N_1987,In_712,In_576);
and U1988 (N_1988,In_494,In_776);
and U1989 (N_1989,In_336,In_120);
xor U1990 (N_1990,In_482,In_902);
and U1991 (N_1991,In_815,In_311);
and U1992 (N_1992,In_614,In_677);
nand U1993 (N_1993,In_127,In_545);
and U1994 (N_1994,In_451,In_693);
nand U1995 (N_1995,In_840,In_252);
and U1996 (N_1996,In_780,In_98);
and U1997 (N_1997,In_230,In_434);
nand U1998 (N_1998,In_378,In_976);
or U1999 (N_1999,In_223,In_761);
nand U2000 (N_2000,In_928,In_125);
nand U2001 (N_2001,In_120,In_783);
nor U2002 (N_2002,In_451,In_573);
nor U2003 (N_2003,In_664,In_515);
nor U2004 (N_2004,In_657,In_541);
nor U2005 (N_2005,In_882,In_735);
xor U2006 (N_2006,In_297,In_570);
nor U2007 (N_2007,In_250,In_990);
nor U2008 (N_2008,In_793,In_800);
nor U2009 (N_2009,In_13,In_1);
nor U2010 (N_2010,In_707,In_184);
and U2011 (N_2011,In_618,In_312);
nand U2012 (N_2012,In_684,In_565);
or U2013 (N_2013,In_431,In_481);
nor U2014 (N_2014,In_248,In_962);
or U2015 (N_2015,In_757,In_307);
nor U2016 (N_2016,In_65,In_405);
or U2017 (N_2017,In_132,In_110);
nand U2018 (N_2018,In_869,In_549);
and U2019 (N_2019,In_385,In_277);
or U2020 (N_2020,In_91,In_639);
nand U2021 (N_2021,In_590,In_882);
xor U2022 (N_2022,In_581,In_44);
nor U2023 (N_2023,In_700,In_996);
or U2024 (N_2024,In_8,In_398);
nand U2025 (N_2025,In_749,In_851);
nor U2026 (N_2026,In_291,In_343);
or U2027 (N_2027,In_945,In_725);
nor U2028 (N_2028,In_379,In_617);
nand U2029 (N_2029,In_728,In_803);
and U2030 (N_2030,In_656,In_749);
and U2031 (N_2031,In_947,In_32);
nand U2032 (N_2032,In_325,In_454);
or U2033 (N_2033,In_364,In_128);
or U2034 (N_2034,In_558,In_653);
nand U2035 (N_2035,In_512,In_10);
nor U2036 (N_2036,In_944,In_945);
nor U2037 (N_2037,In_659,In_619);
xor U2038 (N_2038,In_443,In_287);
nand U2039 (N_2039,In_383,In_591);
and U2040 (N_2040,In_766,In_197);
nor U2041 (N_2041,In_358,In_269);
and U2042 (N_2042,In_625,In_370);
or U2043 (N_2043,In_153,In_576);
or U2044 (N_2044,In_90,In_861);
nor U2045 (N_2045,In_406,In_998);
xnor U2046 (N_2046,In_642,In_52);
nand U2047 (N_2047,In_235,In_722);
nand U2048 (N_2048,In_213,In_92);
nand U2049 (N_2049,In_102,In_847);
or U2050 (N_2050,In_754,In_261);
and U2051 (N_2051,In_524,In_383);
nand U2052 (N_2052,In_250,In_76);
and U2053 (N_2053,In_665,In_208);
xnor U2054 (N_2054,In_323,In_9);
or U2055 (N_2055,In_636,In_795);
or U2056 (N_2056,In_449,In_557);
xnor U2057 (N_2057,In_326,In_227);
nand U2058 (N_2058,In_305,In_510);
and U2059 (N_2059,In_658,In_301);
nand U2060 (N_2060,In_765,In_683);
nor U2061 (N_2061,In_593,In_684);
nor U2062 (N_2062,In_777,In_522);
or U2063 (N_2063,In_488,In_965);
or U2064 (N_2064,In_17,In_564);
nor U2065 (N_2065,In_711,In_529);
nor U2066 (N_2066,In_392,In_799);
and U2067 (N_2067,In_674,In_328);
nor U2068 (N_2068,In_940,In_86);
nand U2069 (N_2069,In_323,In_578);
nor U2070 (N_2070,In_15,In_839);
nor U2071 (N_2071,In_230,In_614);
nor U2072 (N_2072,In_49,In_31);
nand U2073 (N_2073,In_901,In_921);
nand U2074 (N_2074,In_123,In_866);
nand U2075 (N_2075,In_704,In_124);
nor U2076 (N_2076,In_100,In_324);
or U2077 (N_2077,In_149,In_242);
or U2078 (N_2078,In_66,In_951);
nand U2079 (N_2079,In_439,In_779);
nor U2080 (N_2080,In_745,In_540);
or U2081 (N_2081,In_873,In_141);
nand U2082 (N_2082,In_210,In_59);
or U2083 (N_2083,In_713,In_356);
and U2084 (N_2084,In_909,In_466);
nand U2085 (N_2085,In_465,In_407);
and U2086 (N_2086,In_546,In_412);
nand U2087 (N_2087,In_250,In_813);
and U2088 (N_2088,In_895,In_997);
and U2089 (N_2089,In_769,In_977);
and U2090 (N_2090,In_122,In_819);
or U2091 (N_2091,In_125,In_910);
nor U2092 (N_2092,In_9,In_80);
or U2093 (N_2093,In_804,In_655);
or U2094 (N_2094,In_324,In_652);
and U2095 (N_2095,In_809,In_900);
and U2096 (N_2096,In_878,In_726);
or U2097 (N_2097,In_231,In_781);
and U2098 (N_2098,In_888,In_674);
and U2099 (N_2099,In_459,In_616);
nor U2100 (N_2100,In_790,In_909);
or U2101 (N_2101,In_406,In_969);
nand U2102 (N_2102,In_999,In_52);
and U2103 (N_2103,In_442,In_738);
and U2104 (N_2104,In_807,In_525);
nand U2105 (N_2105,In_159,In_782);
and U2106 (N_2106,In_769,In_512);
and U2107 (N_2107,In_306,In_679);
nand U2108 (N_2108,In_163,In_384);
xor U2109 (N_2109,In_29,In_809);
nand U2110 (N_2110,In_238,In_304);
xor U2111 (N_2111,In_345,In_514);
or U2112 (N_2112,In_66,In_235);
xnor U2113 (N_2113,In_918,In_877);
nand U2114 (N_2114,In_337,In_24);
or U2115 (N_2115,In_19,In_829);
or U2116 (N_2116,In_901,In_242);
nor U2117 (N_2117,In_372,In_236);
or U2118 (N_2118,In_644,In_917);
or U2119 (N_2119,In_821,In_246);
and U2120 (N_2120,In_56,In_206);
nor U2121 (N_2121,In_660,In_816);
nand U2122 (N_2122,In_305,In_983);
or U2123 (N_2123,In_785,In_463);
nand U2124 (N_2124,In_944,In_31);
nor U2125 (N_2125,In_661,In_198);
or U2126 (N_2126,In_205,In_347);
nor U2127 (N_2127,In_163,In_302);
and U2128 (N_2128,In_307,In_65);
nor U2129 (N_2129,In_460,In_739);
nand U2130 (N_2130,In_891,In_913);
nor U2131 (N_2131,In_237,In_551);
nor U2132 (N_2132,In_540,In_908);
and U2133 (N_2133,In_438,In_479);
and U2134 (N_2134,In_496,In_7);
and U2135 (N_2135,In_517,In_189);
or U2136 (N_2136,In_283,In_917);
and U2137 (N_2137,In_375,In_43);
and U2138 (N_2138,In_388,In_27);
or U2139 (N_2139,In_290,In_825);
and U2140 (N_2140,In_502,In_803);
nor U2141 (N_2141,In_859,In_102);
xnor U2142 (N_2142,In_857,In_245);
and U2143 (N_2143,In_303,In_574);
or U2144 (N_2144,In_120,In_43);
and U2145 (N_2145,In_622,In_250);
xnor U2146 (N_2146,In_376,In_216);
nor U2147 (N_2147,In_530,In_981);
nor U2148 (N_2148,In_65,In_339);
or U2149 (N_2149,In_666,In_877);
nor U2150 (N_2150,In_544,In_470);
nor U2151 (N_2151,In_696,In_192);
nor U2152 (N_2152,In_759,In_980);
nor U2153 (N_2153,In_690,In_916);
nor U2154 (N_2154,In_450,In_688);
or U2155 (N_2155,In_854,In_911);
nand U2156 (N_2156,In_171,In_514);
nor U2157 (N_2157,In_419,In_746);
and U2158 (N_2158,In_404,In_880);
nor U2159 (N_2159,In_800,In_985);
and U2160 (N_2160,In_864,In_998);
and U2161 (N_2161,In_533,In_274);
or U2162 (N_2162,In_20,In_156);
or U2163 (N_2163,In_727,In_855);
nor U2164 (N_2164,In_860,In_405);
nor U2165 (N_2165,In_847,In_836);
and U2166 (N_2166,In_620,In_119);
and U2167 (N_2167,In_728,In_843);
nor U2168 (N_2168,In_771,In_657);
nand U2169 (N_2169,In_579,In_386);
nor U2170 (N_2170,In_875,In_897);
nand U2171 (N_2171,In_889,In_694);
nor U2172 (N_2172,In_589,In_516);
and U2173 (N_2173,In_113,In_516);
or U2174 (N_2174,In_698,In_764);
or U2175 (N_2175,In_194,In_738);
nand U2176 (N_2176,In_993,In_436);
or U2177 (N_2177,In_688,In_353);
nor U2178 (N_2178,In_294,In_802);
and U2179 (N_2179,In_652,In_594);
nor U2180 (N_2180,In_400,In_918);
and U2181 (N_2181,In_950,In_413);
and U2182 (N_2182,In_498,In_379);
nor U2183 (N_2183,In_293,In_978);
or U2184 (N_2184,In_92,In_971);
or U2185 (N_2185,In_997,In_510);
nand U2186 (N_2186,In_789,In_27);
and U2187 (N_2187,In_382,In_72);
or U2188 (N_2188,In_517,In_634);
or U2189 (N_2189,In_151,In_944);
nand U2190 (N_2190,In_145,In_309);
nor U2191 (N_2191,In_880,In_410);
or U2192 (N_2192,In_28,In_57);
or U2193 (N_2193,In_184,In_247);
nor U2194 (N_2194,In_694,In_832);
nand U2195 (N_2195,In_15,In_866);
nand U2196 (N_2196,In_838,In_145);
xor U2197 (N_2197,In_723,In_623);
and U2198 (N_2198,In_311,In_15);
nand U2199 (N_2199,In_650,In_263);
nor U2200 (N_2200,In_700,In_378);
nand U2201 (N_2201,In_125,In_390);
xnor U2202 (N_2202,In_985,In_814);
or U2203 (N_2203,In_359,In_993);
nor U2204 (N_2204,In_643,In_970);
xor U2205 (N_2205,In_66,In_260);
and U2206 (N_2206,In_913,In_759);
nand U2207 (N_2207,In_440,In_424);
nand U2208 (N_2208,In_551,In_919);
or U2209 (N_2209,In_39,In_58);
and U2210 (N_2210,In_362,In_241);
or U2211 (N_2211,In_870,In_877);
or U2212 (N_2212,In_337,In_710);
and U2213 (N_2213,In_93,In_795);
nand U2214 (N_2214,In_570,In_55);
or U2215 (N_2215,In_876,In_959);
nor U2216 (N_2216,In_462,In_935);
and U2217 (N_2217,In_677,In_153);
nor U2218 (N_2218,In_531,In_497);
and U2219 (N_2219,In_131,In_662);
nand U2220 (N_2220,In_607,In_554);
nand U2221 (N_2221,In_539,In_867);
nor U2222 (N_2222,In_759,In_819);
and U2223 (N_2223,In_758,In_351);
and U2224 (N_2224,In_581,In_619);
nor U2225 (N_2225,In_727,In_240);
nand U2226 (N_2226,In_785,In_149);
nor U2227 (N_2227,In_596,In_180);
and U2228 (N_2228,In_255,In_595);
or U2229 (N_2229,In_75,In_353);
nor U2230 (N_2230,In_746,In_28);
nor U2231 (N_2231,In_845,In_386);
and U2232 (N_2232,In_451,In_607);
and U2233 (N_2233,In_684,In_595);
and U2234 (N_2234,In_95,In_819);
or U2235 (N_2235,In_101,In_337);
nor U2236 (N_2236,In_630,In_315);
nand U2237 (N_2237,In_265,In_941);
or U2238 (N_2238,In_154,In_458);
or U2239 (N_2239,In_289,In_948);
nor U2240 (N_2240,In_216,In_327);
nor U2241 (N_2241,In_420,In_105);
nand U2242 (N_2242,In_957,In_383);
nor U2243 (N_2243,In_865,In_686);
and U2244 (N_2244,In_105,In_506);
or U2245 (N_2245,In_982,In_81);
and U2246 (N_2246,In_598,In_447);
or U2247 (N_2247,In_841,In_603);
and U2248 (N_2248,In_815,In_492);
nand U2249 (N_2249,In_333,In_262);
nor U2250 (N_2250,In_172,In_735);
or U2251 (N_2251,In_834,In_79);
nor U2252 (N_2252,In_994,In_281);
and U2253 (N_2253,In_521,In_797);
nor U2254 (N_2254,In_791,In_835);
nand U2255 (N_2255,In_402,In_119);
nor U2256 (N_2256,In_389,In_826);
and U2257 (N_2257,In_525,In_221);
nor U2258 (N_2258,In_323,In_559);
nor U2259 (N_2259,In_889,In_980);
xnor U2260 (N_2260,In_382,In_959);
or U2261 (N_2261,In_329,In_298);
nand U2262 (N_2262,In_915,In_722);
nand U2263 (N_2263,In_131,In_690);
and U2264 (N_2264,In_775,In_699);
and U2265 (N_2265,In_363,In_11);
nor U2266 (N_2266,In_796,In_24);
and U2267 (N_2267,In_284,In_343);
or U2268 (N_2268,In_966,In_207);
nor U2269 (N_2269,In_870,In_307);
or U2270 (N_2270,In_122,In_971);
or U2271 (N_2271,In_284,In_514);
or U2272 (N_2272,In_840,In_741);
nor U2273 (N_2273,In_168,In_504);
or U2274 (N_2274,In_250,In_154);
nor U2275 (N_2275,In_562,In_854);
or U2276 (N_2276,In_440,In_307);
nor U2277 (N_2277,In_429,In_330);
or U2278 (N_2278,In_136,In_198);
nor U2279 (N_2279,In_444,In_812);
nor U2280 (N_2280,In_335,In_464);
nor U2281 (N_2281,In_685,In_940);
and U2282 (N_2282,In_219,In_720);
nor U2283 (N_2283,In_487,In_153);
nand U2284 (N_2284,In_727,In_837);
and U2285 (N_2285,In_483,In_176);
nor U2286 (N_2286,In_841,In_201);
or U2287 (N_2287,In_632,In_975);
nand U2288 (N_2288,In_474,In_392);
or U2289 (N_2289,In_601,In_228);
nor U2290 (N_2290,In_695,In_809);
nor U2291 (N_2291,In_159,In_924);
nand U2292 (N_2292,In_952,In_46);
or U2293 (N_2293,In_960,In_810);
nor U2294 (N_2294,In_663,In_62);
and U2295 (N_2295,In_770,In_347);
and U2296 (N_2296,In_672,In_754);
or U2297 (N_2297,In_267,In_543);
and U2298 (N_2298,In_95,In_69);
or U2299 (N_2299,In_517,In_905);
and U2300 (N_2300,In_413,In_386);
nand U2301 (N_2301,In_258,In_474);
nor U2302 (N_2302,In_832,In_841);
nor U2303 (N_2303,In_405,In_723);
or U2304 (N_2304,In_584,In_276);
and U2305 (N_2305,In_404,In_669);
and U2306 (N_2306,In_700,In_537);
or U2307 (N_2307,In_93,In_704);
and U2308 (N_2308,In_980,In_802);
or U2309 (N_2309,In_148,In_325);
nand U2310 (N_2310,In_520,In_91);
nor U2311 (N_2311,In_397,In_823);
and U2312 (N_2312,In_486,In_69);
nor U2313 (N_2313,In_204,In_983);
nand U2314 (N_2314,In_966,In_748);
or U2315 (N_2315,In_407,In_837);
and U2316 (N_2316,In_306,In_569);
nor U2317 (N_2317,In_473,In_783);
and U2318 (N_2318,In_379,In_616);
and U2319 (N_2319,In_721,In_36);
nor U2320 (N_2320,In_391,In_965);
or U2321 (N_2321,In_964,In_367);
nor U2322 (N_2322,In_825,In_78);
xnor U2323 (N_2323,In_399,In_75);
nand U2324 (N_2324,In_713,In_292);
nor U2325 (N_2325,In_280,In_824);
nor U2326 (N_2326,In_621,In_839);
and U2327 (N_2327,In_43,In_554);
nand U2328 (N_2328,In_54,In_994);
nand U2329 (N_2329,In_193,In_212);
and U2330 (N_2330,In_215,In_454);
or U2331 (N_2331,In_885,In_747);
or U2332 (N_2332,In_744,In_514);
nand U2333 (N_2333,In_849,In_900);
and U2334 (N_2334,In_514,In_730);
nor U2335 (N_2335,In_641,In_576);
and U2336 (N_2336,In_805,In_382);
nor U2337 (N_2337,In_447,In_131);
nand U2338 (N_2338,In_541,In_215);
nand U2339 (N_2339,In_730,In_995);
nor U2340 (N_2340,In_902,In_195);
nor U2341 (N_2341,In_518,In_323);
and U2342 (N_2342,In_283,In_869);
and U2343 (N_2343,In_290,In_35);
nand U2344 (N_2344,In_18,In_773);
nor U2345 (N_2345,In_573,In_123);
nand U2346 (N_2346,In_136,In_474);
and U2347 (N_2347,In_731,In_886);
nor U2348 (N_2348,In_980,In_582);
or U2349 (N_2349,In_1,In_663);
nor U2350 (N_2350,In_674,In_440);
nand U2351 (N_2351,In_972,In_448);
and U2352 (N_2352,In_605,In_908);
nor U2353 (N_2353,In_347,In_911);
and U2354 (N_2354,In_216,In_796);
nand U2355 (N_2355,In_865,In_490);
nand U2356 (N_2356,In_385,In_995);
nor U2357 (N_2357,In_282,In_501);
and U2358 (N_2358,In_158,In_996);
nor U2359 (N_2359,In_722,In_166);
or U2360 (N_2360,In_812,In_895);
and U2361 (N_2361,In_484,In_440);
nand U2362 (N_2362,In_872,In_716);
xnor U2363 (N_2363,In_181,In_266);
or U2364 (N_2364,In_703,In_168);
nand U2365 (N_2365,In_496,In_467);
xnor U2366 (N_2366,In_552,In_82);
or U2367 (N_2367,In_803,In_984);
nand U2368 (N_2368,In_986,In_189);
nand U2369 (N_2369,In_888,In_819);
nor U2370 (N_2370,In_900,In_22);
nand U2371 (N_2371,In_930,In_958);
nor U2372 (N_2372,In_13,In_758);
nor U2373 (N_2373,In_684,In_76);
nor U2374 (N_2374,In_571,In_317);
or U2375 (N_2375,In_140,In_28);
nand U2376 (N_2376,In_895,In_0);
or U2377 (N_2377,In_147,In_455);
nand U2378 (N_2378,In_554,In_583);
or U2379 (N_2379,In_552,In_794);
nand U2380 (N_2380,In_450,In_260);
and U2381 (N_2381,In_455,In_5);
xor U2382 (N_2382,In_308,In_17);
and U2383 (N_2383,In_368,In_515);
or U2384 (N_2384,In_31,In_465);
nand U2385 (N_2385,In_142,In_160);
and U2386 (N_2386,In_183,In_943);
or U2387 (N_2387,In_898,In_769);
nor U2388 (N_2388,In_336,In_236);
nand U2389 (N_2389,In_112,In_388);
or U2390 (N_2390,In_346,In_801);
and U2391 (N_2391,In_320,In_546);
and U2392 (N_2392,In_72,In_592);
and U2393 (N_2393,In_308,In_499);
nand U2394 (N_2394,In_97,In_243);
or U2395 (N_2395,In_715,In_395);
and U2396 (N_2396,In_417,In_371);
and U2397 (N_2397,In_696,In_80);
nor U2398 (N_2398,In_326,In_346);
or U2399 (N_2399,In_118,In_511);
nor U2400 (N_2400,In_823,In_296);
nor U2401 (N_2401,In_318,In_878);
and U2402 (N_2402,In_871,In_64);
nand U2403 (N_2403,In_136,In_771);
nor U2404 (N_2404,In_47,In_143);
nor U2405 (N_2405,In_235,In_666);
nand U2406 (N_2406,In_382,In_490);
and U2407 (N_2407,In_408,In_472);
nand U2408 (N_2408,In_528,In_194);
nand U2409 (N_2409,In_81,In_973);
or U2410 (N_2410,In_224,In_14);
nor U2411 (N_2411,In_88,In_290);
or U2412 (N_2412,In_811,In_288);
xnor U2413 (N_2413,In_453,In_242);
and U2414 (N_2414,In_249,In_369);
nor U2415 (N_2415,In_129,In_744);
or U2416 (N_2416,In_929,In_364);
and U2417 (N_2417,In_732,In_141);
or U2418 (N_2418,In_22,In_600);
or U2419 (N_2419,In_759,In_312);
nor U2420 (N_2420,In_711,In_113);
and U2421 (N_2421,In_278,In_573);
xnor U2422 (N_2422,In_258,In_185);
and U2423 (N_2423,In_840,In_545);
or U2424 (N_2424,In_429,In_340);
nand U2425 (N_2425,In_249,In_580);
xnor U2426 (N_2426,In_397,In_593);
nor U2427 (N_2427,In_21,In_767);
nor U2428 (N_2428,In_576,In_804);
or U2429 (N_2429,In_26,In_943);
nand U2430 (N_2430,In_357,In_824);
nand U2431 (N_2431,In_290,In_380);
nand U2432 (N_2432,In_65,In_157);
nand U2433 (N_2433,In_222,In_927);
nand U2434 (N_2434,In_325,In_983);
and U2435 (N_2435,In_256,In_282);
and U2436 (N_2436,In_781,In_517);
nand U2437 (N_2437,In_826,In_90);
or U2438 (N_2438,In_349,In_859);
or U2439 (N_2439,In_684,In_63);
nand U2440 (N_2440,In_798,In_687);
and U2441 (N_2441,In_433,In_490);
and U2442 (N_2442,In_514,In_350);
and U2443 (N_2443,In_77,In_2);
nand U2444 (N_2444,In_142,In_397);
nand U2445 (N_2445,In_47,In_875);
nand U2446 (N_2446,In_515,In_589);
and U2447 (N_2447,In_748,In_192);
xnor U2448 (N_2448,In_851,In_895);
nand U2449 (N_2449,In_398,In_902);
xnor U2450 (N_2450,In_788,In_480);
nor U2451 (N_2451,In_340,In_207);
or U2452 (N_2452,In_429,In_909);
nand U2453 (N_2453,In_843,In_361);
and U2454 (N_2454,In_939,In_931);
nand U2455 (N_2455,In_990,In_270);
nand U2456 (N_2456,In_330,In_168);
and U2457 (N_2457,In_701,In_436);
nor U2458 (N_2458,In_19,In_192);
and U2459 (N_2459,In_598,In_177);
or U2460 (N_2460,In_571,In_457);
nor U2461 (N_2461,In_34,In_5);
nand U2462 (N_2462,In_260,In_836);
or U2463 (N_2463,In_108,In_201);
nor U2464 (N_2464,In_891,In_718);
and U2465 (N_2465,In_134,In_437);
and U2466 (N_2466,In_883,In_324);
nor U2467 (N_2467,In_586,In_320);
or U2468 (N_2468,In_258,In_501);
or U2469 (N_2469,In_920,In_986);
nor U2470 (N_2470,In_214,In_514);
and U2471 (N_2471,In_747,In_256);
or U2472 (N_2472,In_867,In_210);
nand U2473 (N_2473,In_468,In_237);
nor U2474 (N_2474,In_688,In_934);
nor U2475 (N_2475,In_727,In_454);
and U2476 (N_2476,In_966,In_791);
nand U2477 (N_2477,In_209,In_386);
or U2478 (N_2478,In_551,In_865);
nor U2479 (N_2479,In_812,In_28);
nand U2480 (N_2480,In_884,In_1);
nand U2481 (N_2481,In_553,In_597);
nor U2482 (N_2482,In_392,In_777);
nand U2483 (N_2483,In_159,In_906);
nand U2484 (N_2484,In_978,In_387);
or U2485 (N_2485,In_248,In_342);
or U2486 (N_2486,In_861,In_166);
or U2487 (N_2487,In_374,In_292);
and U2488 (N_2488,In_482,In_120);
or U2489 (N_2489,In_141,In_742);
nand U2490 (N_2490,In_25,In_519);
nor U2491 (N_2491,In_628,In_534);
nor U2492 (N_2492,In_152,In_321);
nor U2493 (N_2493,In_201,In_932);
nand U2494 (N_2494,In_73,In_687);
and U2495 (N_2495,In_735,In_871);
and U2496 (N_2496,In_264,In_976);
and U2497 (N_2497,In_720,In_10);
or U2498 (N_2498,In_830,In_813);
nor U2499 (N_2499,In_600,In_758);
or U2500 (N_2500,N_2468,N_134);
nor U2501 (N_2501,N_2258,N_2201);
nor U2502 (N_2502,N_1468,N_2026);
and U2503 (N_2503,N_1327,N_1058);
or U2504 (N_2504,N_469,N_1068);
and U2505 (N_2505,N_428,N_1105);
nor U2506 (N_2506,N_2248,N_2017);
and U2507 (N_2507,N_889,N_636);
xor U2508 (N_2508,N_1528,N_239);
nand U2509 (N_2509,N_1510,N_1989);
or U2510 (N_2510,N_475,N_2305);
nor U2511 (N_2511,N_753,N_1939);
and U2512 (N_2512,N_1849,N_40);
nand U2513 (N_2513,N_850,N_2157);
or U2514 (N_2514,N_1474,N_1863);
nand U2515 (N_2515,N_1493,N_1031);
nand U2516 (N_2516,N_711,N_162);
and U2517 (N_2517,N_1577,N_1896);
and U2518 (N_2518,N_1888,N_839);
or U2519 (N_2519,N_863,N_446);
nor U2520 (N_2520,N_1312,N_2125);
nand U2521 (N_2521,N_315,N_2287);
nand U2522 (N_2522,N_1171,N_525);
nand U2523 (N_2523,N_1672,N_2316);
xnor U2524 (N_2524,N_627,N_1937);
and U2525 (N_2525,N_1842,N_1460);
xnor U2526 (N_2526,N_2373,N_356);
nand U2527 (N_2527,N_188,N_985);
nor U2528 (N_2528,N_30,N_922);
nand U2529 (N_2529,N_1366,N_614);
nand U2530 (N_2530,N_258,N_398);
nand U2531 (N_2531,N_1355,N_1913);
xnor U2532 (N_2532,N_524,N_1673);
nor U2533 (N_2533,N_1783,N_909);
and U2534 (N_2534,N_2033,N_1763);
nand U2535 (N_2535,N_2035,N_1648);
nor U2536 (N_2536,N_1950,N_2318);
and U2537 (N_2537,N_2402,N_1288);
nand U2538 (N_2538,N_399,N_1554);
nand U2539 (N_2539,N_1889,N_759);
nand U2540 (N_2540,N_1419,N_1008);
nand U2541 (N_2541,N_632,N_2296);
nand U2542 (N_2542,N_2431,N_267);
nand U2543 (N_2543,N_2022,N_384);
nand U2544 (N_2544,N_146,N_370);
nand U2545 (N_2545,N_1906,N_1866);
or U2546 (N_2546,N_2218,N_1861);
and U2547 (N_2547,N_2117,N_89);
nand U2548 (N_2548,N_1152,N_198);
nor U2549 (N_2549,N_2036,N_1582);
nor U2550 (N_2550,N_2114,N_1848);
nor U2551 (N_2551,N_1410,N_1765);
and U2552 (N_2552,N_713,N_1162);
nand U2553 (N_2553,N_184,N_447);
nand U2554 (N_2554,N_876,N_715);
nor U2555 (N_2555,N_859,N_2052);
nor U2556 (N_2556,N_2369,N_1604);
nand U2557 (N_2557,N_1575,N_63);
or U2558 (N_2558,N_1340,N_1482);
nand U2559 (N_2559,N_799,N_1702);
nand U2560 (N_2560,N_435,N_246);
or U2561 (N_2561,N_893,N_2070);
nor U2562 (N_2562,N_987,N_1453);
or U2563 (N_2563,N_76,N_301);
and U2564 (N_2564,N_642,N_1051);
nand U2565 (N_2565,N_942,N_2029);
and U2566 (N_2566,N_1285,N_275);
or U2567 (N_2567,N_982,N_1155);
and U2568 (N_2568,N_2471,N_328);
and U2569 (N_2569,N_169,N_1899);
or U2570 (N_2570,N_66,N_1801);
nand U2571 (N_2571,N_2365,N_2105);
nand U2572 (N_2572,N_1643,N_1103);
and U2573 (N_2573,N_2192,N_1235);
nand U2574 (N_2574,N_1274,N_1841);
nor U2575 (N_2575,N_2356,N_1399);
or U2576 (N_2576,N_760,N_490);
nand U2577 (N_2577,N_1484,N_453);
nand U2578 (N_2578,N_718,N_564);
and U2579 (N_2579,N_686,N_758);
or U2580 (N_2580,N_1886,N_459);
and U2581 (N_2581,N_1465,N_1398);
nand U2582 (N_2582,N_928,N_1443);
or U2583 (N_2583,N_2412,N_1876);
or U2584 (N_2584,N_113,N_828);
and U2585 (N_2585,N_923,N_2133);
or U2586 (N_2586,N_941,N_1033);
nand U2587 (N_2587,N_1471,N_1035);
or U2588 (N_2588,N_242,N_1266);
nor U2589 (N_2589,N_2185,N_515);
or U2590 (N_2590,N_41,N_61);
or U2591 (N_2591,N_350,N_1494);
or U2592 (N_2592,N_875,N_1233);
and U2593 (N_2593,N_628,N_1978);
and U2594 (N_2594,N_1588,N_1722);
nand U2595 (N_2595,N_1855,N_694);
or U2596 (N_2596,N_1160,N_1319);
nand U2597 (N_2597,N_1001,N_1979);
and U2598 (N_2598,N_741,N_764);
or U2599 (N_2599,N_1902,N_1810);
or U2600 (N_2600,N_196,N_1418);
or U2601 (N_2601,N_1449,N_96);
nand U2602 (N_2602,N_1167,N_1628);
nand U2603 (N_2603,N_2443,N_1436);
nand U2604 (N_2604,N_2415,N_426);
and U2605 (N_2605,N_2380,N_1789);
and U2606 (N_2606,N_331,N_1372);
nor U2607 (N_2607,N_1074,N_556);
nor U2608 (N_2608,N_818,N_2276);
nand U2609 (N_2609,N_699,N_1712);
or U2610 (N_2610,N_354,N_2233);
and U2611 (N_2611,N_379,N_1873);
or U2612 (N_2612,N_1395,N_1935);
nor U2613 (N_2613,N_28,N_245);
nand U2614 (N_2614,N_1748,N_2224);
or U2615 (N_2615,N_927,N_1469);
nor U2616 (N_2616,N_1335,N_1788);
and U2617 (N_2617,N_2436,N_199);
or U2618 (N_2618,N_974,N_705);
and U2619 (N_2619,N_1703,N_1870);
nand U2620 (N_2620,N_665,N_2271);
and U2621 (N_2621,N_268,N_2165);
or U2622 (N_2622,N_1428,N_794);
and U2623 (N_2623,N_164,N_1557);
xor U2624 (N_2624,N_259,N_2363);
xnor U2625 (N_2625,N_429,N_2025);
or U2626 (N_2626,N_1751,N_93);
or U2627 (N_2627,N_1221,N_58);
or U2628 (N_2628,N_406,N_2068);
and U2629 (N_2629,N_1202,N_809);
nor U2630 (N_2630,N_1097,N_1324);
nand U2631 (N_2631,N_1017,N_1151);
and U2632 (N_2632,N_1323,N_2190);
or U2633 (N_2633,N_948,N_1424);
or U2634 (N_2634,N_1691,N_170);
or U2635 (N_2635,N_717,N_1574);
or U2636 (N_2636,N_731,N_810);
nand U2637 (N_2637,N_1804,N_656);
nand U2638 (N_2638,N_579,N_53);
and U2639 (N_2639,N_119,N_658);
or U2640 (N_2640,N_1214,N_2067);
and U2641 (N_2641,N_1966,N_473);
or U2642 (N_2642,N_86,N_1882);
and U2643 (N_2643,N_885,N_1178);
nand U2644 (N_2644,N_357,N_880);
nor U2645 (N_2645,N_1367,N_1525);
nor U2646 (N_2646,N_1927,N_795);
nand U2647 (N_2647,N_770,N_2394);
nand U2648 (N_2648,N_1715,N_445);
and U2649 (N_2649,N_1364,N_1092);
and U2650 (N_2650,N_1096,N_2166);
xor U2651 (N_2651,N_1857,N_270);
nor U2652 (N_2652,N_2262,N_299);
nor U2653 (N_2653,N_2191,N_1706);
and U2654 (N_2654,N_1153,N_156);
or U2655 (N_2655,N_913,N_1503);
nor U2656 (N_2656,N_844,N_1807);
nor U2657 (N_2657,N_2461,N_1511);
nand U2658 (N_2658,N_2331,N_266);
and U2659 (N_2659,N_787,N_1635);
and U2660 (N_2660,N_819,N_2348);
nor U2661 (N_2661,N_1800,N_2072);
nand U2662 (N_2662,N_1346,N_434);
nand U2663 (N_2663,N_975,N_1980);
nand U2664 (N_2664,N_2354,N_1455);
nor U2665 (N_2665,N_2139,N_1618);
or U2666 (N_2666,N_1417,N_2441);
nand U2667 (N_2667,N_2328,N_1144);
or U2668 (N_2668,N_683,N_1191);
or U2669 (N_2669,N_1249,N_2132);
nand U2670 (N_2670,N_1523,N_1661);
nand U2671 (N_2671,N_1206,N_1885);
or U2672 (N_2672,N_1388,N_444);
nor U2673 (N_2673,N_931,N_2372);
and U2674 (N_2674,N_2249,N_521);
and U2675 (N_2675,N_1678,N_405);
or U2676 (N_2676,N_1595,N_36);
nand U2677 (N_2677,N_4,N_1081);
or U2678 (N_2678,N_827,N_1006);
nor U2679 (N_2679,N_565,N_2102);
and U2680 (N_2680,N_211,N_2491);
or U2681 (N_2681,N_2315,N_1229);
nand U2682 (N_2682,N_771,N_286);
nor U2683 (N_2683,N_1599,N_1542);
and U2684 (N_2684,N_2288,N_281);
or U2685 (N_2685,N_1687,N_2307);
nor U2686 (N_2686,N_19,N_804);
nand U2687 (N_2687,N_1490,N_1454);
or U2688 (N_2688,N_2155,N_1560);
nand U2689 (N_2689,N_2217,N_414);
or U2690 (N_2690,N_2278,N_1875);
nor U2691 (N_2691,N_1723,N_652);
nand U2692 (N_2692,N_2467,N_2416);
xnor U2693 (N_2693,N_1272,N_674);
nor U2694 (N_2694,N_2,N_495);
nand U2695 (N_2695,N_411,N_1117);
or U2696 (N_2696,N_176,N_892);
and U2697 (N_2697,N_905,N_1883);
nand U2698 (N_2698,N_2175,N_2401);
nand U2699 (N_2699,N_1880,N_2024);
or U2700 (N_2700,N_1287,N_1948);
or U2701 (N_2701,N_1034,N_786);
or U2702 (N_2702,N_2069,N_2489);
and U2703 (N_2703,N_99,N_750);
or U2704 (N_2704,N_2213,N_1425);
or U2705 (N_2705,N_1743,N_236);
nor U2706 (N_2706,N_2140,N_1086);
nor U2707 (N_2707,N_333,N_1492);
nand U2708 (N_2708,N_825,N_1241);
and U2709 (N_2709,N_1878,N_2339);
or U2710 (N_2710,N_2151,N_1015);
or U2711 (N_2711,N_820,N_531);
nor U2712 (N_2712,N_1853,N_1548);
or U2713 (N_2713,N_327,N_836);
or U2714 (N_2714,N_2014,N_580);
and U2715 (N_2715,N_1351,N_597);
nand U2716 (N_2716,N_75,N_70);
and U2717 (N_2717,N_1124,N_2089);
nand U2718 (N_2718,N_371,N_882);
nand U2719 (N_2719,N_373,N_18);
and U2720 (N_2720,N_486,N_765);
or U2721 (N_2721,N_2194,N_2368);
nor U2722 (N_2722,N_1243,N_639);
nor U2723 (N_2723,N_2388,N_846);
nand U2724 (N_2724,N_2426,N_2205);
nor U2725 (N_2725,N_952,N_1964);
and U2726 (N_2726,N_1467,N_623);
and U2727 (N_2727,N_1383,N_1688);
xnor U2728 (N_2728,N_2223,N_2381);
or U2729 (N_2729,N_2138,N_142);
or U2730 (N_2730,N_569,N_1255);
and U2731 (N_2731,N_1877,N_132);
nand U2732 (N_2732,N_547,N_1825);
nor U2733 (N_2733,N_2438,N_2281);
or U2734 (N_2734,N_568,N_374);
or U2735 (N_2735,N_1063,N_1440);
and U2736 (N_2736,N_1738,N_1573);
and U2737 (N_2737,N_1282,N_1529);
nor U2738 (N_2738,N_2387,N_1023);
and U2739 (N_2739,N_462,N_265);
and U2740 (N_2740,N_90,N_34);
and U2741 (N_2741,N_1251,N_180);
nand U2742 (N_2742,N_1048,N_210);
or U2743 (N_2743,N_2337,N_2392);
nand U2744 (N_2744,N_944,N_8);
or U2745 (N_2745,N_995,N_141);
nand U2746 (N_2746,N_2285,N_2207);
nor U2747 (N_2747,N_1971,N_1742);
nor U2748 (N_2748,N_1683,N_1594);
nand U2749 (N_2749,N_2150,N_79);
and U2750 (N_2750,N_480,N_1280);
and U2751 (N_2751,N_2179,N_1815);
or U2752 (N_2752,N_601,N_1375);
nand U2753 (N_2753,N_672,N_1495);
or U2754 (N_2754,N_1836,N_872);
and U2755 (N_2755,N_62,N_2290);
nor U2756 (N_2756,N_26,N_467);
nor U2757 (N_2757,N_822,N_1333);
nand U2758 (N_2758,N_575,N_2172);
nor U2759 (N_2759,N_2108,N_2044);
and U2760 (N_2760,N_1159,N_71);
nand U2761 (N_2761,N_2366,N_2259);
or U2762 (N_2762,N_342,N_2228);
nand U2763 (N_2763,N_2286,N_2349);
nand U2764 (N_2764,N_2264,N_2367);
nor U2765 (N_2765,N_1360,N_386);
or U2766 (N_2766,N_1318,N_365);
nand U2767 (N_2767,N_1727,N_1504);
nand U2768 (N_2768,N_2031,N_2137);
and U2769 (N_2769,N_360,N_1201);
and U2770 (N_2770,N_121,N_2235);
nor U2771 (N_2771,N_1596,N_687);
and U2772 (N_2772,N_1128,N_1970);
and U2773 (N_2773,N_2393,N_1309);
nand U2774 (N_2774,N_1275,N_830);
and U2775 (N_2775,N_1865,N_1326);
and U2776 (N_2776,N_2209,N_899);
or U2777 (N_2777,N_51,N_910);
nor U2778 (N_2778,N_1030,N_408);
and U2779 (N_2779,N_324,N_845);
nor U2780 (N_2780,N_2481,N_1717);
and U2781 (N_2781,N_1580,N_1371);
nor U2782 (N_2782,N_2109,N_2230);
and U2783 (N_2783,N_2147,N_1852);
and U2784 (N_2784,N_898,N_1037);
nor U2785 (N_2785,N_2314,N_229);
nor U2786 (N_2786,N_805,N_2016);
or U2787 (N_2787,N_917,N_92);
or U2788 (N_2788,N_938,N_2239);
xnor U2789 (N_2789,N_2263,N_1046);
and U2790 (N_2790,N_341,N_2162);
xnor U2791 (N_2791,N_91,N_1342);
and U2792 (N_2792,N_1354,N_1150);
or U2793 (N_2793,N_904,N_2008);
nor U2794 (N_2794,N_1666,N_1983);
nand U2795 (N_2795,N_1986,N_730);
or U2796 (N_2796,N_529,N_1294);
and U2797 (N_2797,N_1085,N_2126);
nor U2798 (N_2798,N_349,N_282);
nand U2799 (N_2799,N_1846,N_2340);
nor U2800 (N_2800,N_663,N_1115);
nand U2801 (N_2801,N_477,N_271);
nand U2802 (N_2802,N_2289,N_769);
or U2803 (N_2803,N_2304,N_2360);
and U2804 (N_2804,N_1403,N_930);
or U2805 (N_2805,N_1740,N_305);
nand U2806 (N_2806,N_2066,N_2028);
nor U2807 (N_2807,N_1920,N_743);
nor U2808 (N_2808,N_864,N_1479);
nor U2809 (N_2809,N_1791,N_1600);
or U2810 (N_2810,N_1695,N_2232);
and U2811 (N_2811,N_138,N_2435);
nor U2812 (N_2812,N_2269,N_744);
and U2813 (N_2813,N_310,N_1969);
or U2814 (N_2814,N_207,N_1129);
and U2815 (N_2815,N_650,N_693);
or U2816 (N_2816,N_849,N_1427);
and U2817 (N_2817,N_1158,N_46);
or U2818 (N_2818,N_1502,N_1644);
nor U2819 (N_2819,N_1254,N_842);
nor U2820 (N_2820,N_1198,N_961);
or U2821 (N_2821,N_32,N_158);
nor U2822 (N_2822,N_2127,N_500);
and U2823 (N_2823,N_1918,N_1689);
nor U2824 (N_2824,N_1653,N_599);
nor U2825 (N_2825,N_1378,N_1116);
and U2826 (N_2826,N_1382,N_60);
nor U2827 (N_2827,N_127,N_782);
or U2828 (N_2828,N_2374,N_2032);
nor U2829 (N_2829,N_998,N_56);
nor U2830 (N_2830,N_2414,N_1820);
or U2831 (N_2831,N_1140,N_817);
or U2832 (N_2832,N_11,N_746);
or U2833 (N_2833,N_2479,N_2274);
and U2834 (N_2834,N_867,N_122);
nor U2835 (N_2835,N_102,N_1154);
or U2836 (N_2836,N_755,N_1212);
nor U2837 (N_2837,N_83,N_1929);
and U2838 (N_2838,N_1990,N_2131);
or U2839 (N_2839,N_219,N_1619);
nand U2840 (N_2840,N_111,N_1744);
and U2841 (N_2841,N_424,N_1515);
and U2842 (N_2842,N_2265,N_1387);
nor U2843 (N_2843,N_2445,N_2427);
and U2844 (N_2844,N_726,N_1268);
and U2845 (N_2845,N_322,N_307);
or U2846 (N_2846,N_317,N_1615);
or U2847 (N_2847,N_1328,N_692);
or U2848 (N_2848,N_1559,N_2112);
and U2849 (N_2849,N_277,N_958);
or U2850 (N_2850,N_50,N_689);
or U2851 (N_2851,N_1397,N_213);
or U2852 (N_2852,N_1640,N_2247);
nand U2853 (N_2853,N_1322,N_816);
nor U2854 (N_2854,N_2189,N_1071);
and U2855 (N_2855,N_1414,N_1442);
and U2856 (N_2856,N_708,N_1208);
or U2857 (N_2857,N_654,N_668);
xnor U2858 (N_2858,N_410,N_609);
xnor U2859 (N_2859,N_2227,N_478);
nand U2860 (N_2860,N_1112,N_465);
nor U2861 (N_2861,N_2483,N_318);
or U2862 (N_2862,N_2335,N_1977);
xnor U2863 (N_2863,N_1729,N_800);
or U2864 (N_2864,N_971,N_82);
nor U2865 (N_2865,N_588,N_773);
nor U2866 (N_2866,N_1834,N_2183);
nand U2867 (N_2867,N_1924,N_1812);
nand U2868 (N_2868,N_1100,N_2094);
nand U2869 (N_2869,N_811,N_1499);
or U2870 (N_2870,N_77,N_544);
xnor U2871 (N_2871,N_130,N_681);
nor U2872 (N_2872,N_796,N_2152);
and U2873 (N_2873,N_2219,N_1752);
nand U2874 (N_2874,N_2425,N_1148);
and U2875 (N_2875,N_1405,N_1130);
and U2876 (N_2876,N_1769,N_707);
and U2877 (N_2877,N_1172,N_712);
nor U2878 (N_2878,N_2007,N_1125);
nor U2879 (N_2879,N_437,N_1463);
nor U2880 (N_2880,N_664,N_2496);
and U2881 (N_2881,N_2176,N_181);
nor U2882 (N_2882,N_2199,N_352);
and U2883 (N_2883,N_95,N_545);
nand U2884 (N_2884,N_2330,N_631);
and U2885 (N_2885,N_2055,N_857);
nand U2886 (N_2886,N_2297,N_1697);
and U2887 (N_2887,N_1291,N_27);
or U2888 (N_2888,N_1185,N_1018);
and U2889 (N_2889,N_1612,N_1536);
and U2890 (N_2890,N_204,N_438);
or U2891 (N_2891,N_1867,N_1407);
or U2892 (N_2892,N_1753,N_716);
nand U2893 (N_2893,N_367,N_725);
and U2894 (N_2894,N_1331,N_49);
nor U2895 (N_2895,N_1524,N_2364);
xnor U2896 (N_2896,N_2119,N_695);
nor U2897 (N_2897,N_2204,N_1358);
nor U2898 (N_2898,N_749,N_1147);
xnor U2899 (N_2899,N_202,N_418);
nor U2900 (N_2900,N_291,N_596);
or U2901 (N_2901,N_402,N_1664);
nor U2902 (N_2902,N_2423,N_1713);
and U2903 (N_2903,N_485,N_1591);
nor U2904 (N_2904,N_1416,N_1222);
and U2905 (N_2905,N_835,N_2193);
nor U2906 (N_2906,N_284,N_651);
or U2907 (N_2907,N_2039,N_906);
or U2908 (N_2908,N_2107,N_1119);
and U2909 (N_2909,N_1660,N_1728);
or U2910 (N_2910,N_807,N_1634);
nand U2911 (N_2911,N_2391,N_1982);
or U2912 (N_2912,N_1337,N_1109);
and U2913 (N_2913,N_1451,N_432);
and U2914 (N_2914,N_570,N_1802);
or U2915 (N_2915,N_2073,N_574);
and U2916 (N_2916,N_2341,N_1256);
and U2917 (N_2917,N_2148,N_2000);
nor U2918 (N_2918,N_2211,N_598);
nand U2919 (N_2919,N_1607,N_368);
nor U2920 (N_2920,N_1512,N_1163);
nand U2921 (N_2921,N_1146,N_375);
nor U2922 (N_2922,N_673,N_2319);
or U2923 (N_2923,N_1265,N_612);
nor U2924 (N_2924,N_1393,N_611);
nand U2925 (N_2925,N_1078,N_983);
and U2926 (N_2926,N_1283,N_458);
or U2927 (N_2927,N_1408,N_1556);
or U2928 (N_2928,N_513,N_2096);
nor U2929 (N_2929,N_552,N_2455);
or U2930 (N_2930,N_1317,N_1052);
xnor U2931 (N_2931,N_1149,N_1350);
nor U2932 (N_2932,N_748,N_2499);
and U2933 (N_2933,N_516,N_780);
and U2934 (N_2934,N_355,N_1749);
or U2935 (N_2935,N_1731,N_1624);
nand U2936 (N_2936,N_2384,N_2111);
nor U2937 (N_2937,N_1516,N_319);
and U2938 (N_2938,N_1422,N_582);
or U2939 (N_2939,N_2011,N_2283);
nor U2940 (N_2940,N_172,N_263);
or U2941 (N_2941,N_1083,N_1627);
nand U2942 (N_2942,N_2236,N_2180);
or U2943 (N_2943,N_1002,N_562);
nor U2944 (N_2944,N_676,N_511);
nor U2945 (N_2945,N_2267,N_359);
nor U2946 (N_2946,N_2163,N_874);
nand U2947 (N_2947,N_2103,N_1796);
or U2948 (N_2948,N_273,N_1064);
nor U2949 (N_2949,N_363,N_39);
nand U2950 (N_2950,N_2434,N_1025);
or U2951 (N_2951,N_1082,N_2303);
and U2952 (N_2952,N_577,N_926);
or U2953 (N_2953,N_969,N_289);
and U2954 (N_2954,N_1781,N_260);
nand U2955 (N_2955,N_2170,N_2018);
nand U2956 (N_2956,N_2083,N_72);
and U2957 (N_2957,N_2167,N_1385);
or U2958 (N_2958,N_1629,N_996);
and U2959 (N_2959,N_1923,N_1381);
nor U2960 (N_2960,N_2085,N_2306);
nand U2961 (N_2961,N_1677,N_422);
nand U2962 (N_2962,N_540,N_1497);
and U2963 (N_2963,N_100,N_1633);
nor U2964 (N_2964,N_1551,N_616);
and U2965 (N_2965,N_1281,N_152);
and U2966 (N_2966,N_1872,N_756);
and U2967 (N_2967,N_1732,N_933);
nand U2968 (N_2968,N_1412,N_973);
or U2969 (N_2969,N_585,N_1997);
nand U2970 (N_2970,N_1338,N_2023);
or U2971 (N_2971,N_2473,N_2317);
and U2972 (N_2972,N_806,N_157);
nand U2973 (N_2973,N_1278,N_655);
nor U2974 (N_2974,N_228,N_230);
nor U2975 (N_2975,N_205,N_2399);
nand U2976 (N_2976,N_514,N_1754);
nand U2977 (N_2977,N_1180,N_225);
or U2978 (N_2978,N_1795,N_2203);
nor U2979 (N_2979,N_881,N_1726);
nand U2980 (N_2980,N_2336,N_1840);
xnor U2981 (N_2981,N_1332,N_2400);
or U2982 (N_2982,N_1005,N_2327);
nor U2983 (N_2983,N_999,N_2104);
xnor U2984 (N_2984,N_1730,N_54);
or U2985 (N_2985,N_2313,N_1839);
and U2986 (N_2986,N_392,N_1879);
or U2987 (N_2987,N_1404,N_2158);
and U2988 (N_2988,N_2302,N_1797);
or U2989 (N_2989,N_214,N_250);
or U2990 (N_2990,N_1864,N_1194);
or U2991 (N_2991,N_2260,N_518);
or U2992 (N_2992,N_1157,N_1234);
and U2993 (N_2993,N_1674,N_2051);
or U2994 (N_2994,N_1960,N_2418);
nand U2995 (N_2995,N_1306,N_1587);
and U2996 (N_2996,N_1758,N_936);
or U2997 (N_2997,N_1447,N_870);
and U2998 (N_2998,N_419,N_2242);
and U2999 (N_2999,N_1477,N_2338);
and U3000 (N_3000,N_276,N_2160);
and U3001 (N_3001,N_2472,N_182);
and U3002 (N_3002,N_2122,N_1406);
or U3003 (N_3003,N_622,N_2099);
or U3004 (N_3004,N_2145,N_919);
nand U3005 (N_3005,N_866,N_1868);
or U3006 (N_3006,N_2323,N_1696);
or U3007 (N_3007,N_1205,N_2097);
or U3008 (N_3008,N_900,N_1);
nor U3009 (N_3009,N_1122,N_238);
nor U3010 (N_3010,N_1652,N_2293);
and U3011 (N_3011,N_361,N_861);
or U3012 (N_3012,N_1571,N_2053);
nor U3013 (N_3013,N_2298,N_159);
nand U3014 (N_3014,N_1021,N_1799);
xnor U3015 (N_3015,N_733,N_44);
nand U3016 (N_3016,N_346,N_2121);
nor U3017 (N_3017,N_116,N_413);
and U3018 (N_3018,N_1489,N_1223);
or U3019 (N_3019,N_2003,N_1373);
or U3020 (N_3020,N_2240,N_85);
or U3021 (N_3021,N_297,N_1423);
nor U3022 (N_3022,N_1301,N_1993);
nand U3023 (N_3023,N_2272,N_1359);
xnor U3024 (N_3024,N_1597,N_785);
and U3025 (N_3025,N_2474,N_378);
and U3026 (N_3026,N_2347,N_959);
or U3027 (N_3027,N_380,N_1762);
nand U3028 (N_3028,N_2006,N_2406);
nor U3029 (N_3029,N_1922,N_783);
xnor U3030 (N_3030,N_326,N_2291);
nor U3031 (N_3031,N_763,N_624);
nand U3032 (N_3032,N_2020,N_1850);
and U3033 (N_3033,N_1508,N_2322);
nand U3034 (N_3034,N_2404,N_2019);
or U3035 (N_3035,N_979,N_1297);
xor U3036 (N_3036,N_1343,N_620);
or U3037 (N_3037,N_1543,N_2222);
nand U3038 (N_3038,N_912,N_607);
nand U3039 (N_3039,N_934,N_1623);
nor U3040 (N_3040,N_522,N_487);
and U3041 (N_3041,N_548,N_1299);
nor U3042 (N_3042,N_1780,N_1136);
nand U3043 (N_3043,N_339,N_1118);
nand U3044 (N_3044,N_1632,N_1040);
nor U3045 (N_3045,N_1267,N_968);
nor U3046 (N_3046,N_1303,N_1230);
or U3047 (N_3047,N_1057,N_1509);
nor U3048 (N_3048,N_1773,N_212);
and U3049 (N_3049,N_186,N_992);
nand U3050 (N_3050,N_1583,N_421);
nor U3051 (N_3051,N_1290,N_232);
nand U3052 (N_3052,N_1611,N_1028);
xnor U3053 (N_3053,N_1095,N_1253);
and U3054 (N_3054,N_84,N_295);
and U3055 (N_3055,N_1658,N_932);
and U3056 (N_3056,N_1339,N_915);
nand U3057 (N_3057,N_549,N_1625);
nor U3058 (N_3058,N_1061,N_1871);
or U3059 (N_3059,N_550,N_1269);
nor U3060 (N_3060,N_1941,N_1426);
nor U3061 (N_3061,N_221,N_2110);
and U3062 (N_3062,N_1481,N_724);
nor U3063 (N_3063,N_965,N_1998);
and U3064 (N_3064,N_2419,N_394);
or U3065 (N_3065,N_42,N_461);
or U3066 (N_3066,N_136,N_1041);
nand U3067 (N_3067,N_2456,N_166);
nor U3068 (N_3068,N_131,N_1012);
nand U3069 (N_3069,N_1589,N_2346);
and U3070 (N_3070,N_2430,N_1821);
nor U3071 (N_3071,N_1655,N_165);
and U3072 (N_3072,N_1391,N_602);
or U3073 (N_3073,N_1345,N_1485);
or U3074 (N_3074,N_1759,N_1298);
nand U3075 (N_3075,N_2359,N_2250);
and U3076 (N_3076,N_412,N_35);
and U3077 (N_3077,N_645,N_1377);
nand U3078 (N_3078,N_2403,N_593);
nor U3079 (N_3079,N_2476,N_2045);
nor U3080 (N_3080,N_878,N_2396);
nand U3081 (N_3081,N_1507,N_814);
or U3082 (N_3082,N_1321,N_1884);
nor U3083 (N_3083,N_1755,N_2449);
or U3084 (N_3084,N_535,N_2135);
nand U3085 (N_3085,N_2049,N_235);
nor U3086 (N_3086,N_1009,N_2494);
xor U3087 (N_3087,N_1680,N_851);
or U3088 (N_3088,N_1179,N_2161);
nor U3089 (N_3089,N_1362,N_1305);
or U3090 (N_3090,N_248,N_2353);
nor U3091 (N_3091,N_595,N_31);
nor U3092 (N_3092,N_1177,N_2385);
nand U3093 (N_3093,N_1808,N_2141);
nor U3094 (N_3094,N_1374,N_853);
and U3095 (N_3095,N_2464,N_1965);
and U3096 (N_3096,N_252,N_1916);
nor U3097 (N_3097,N_140,N_2310);
nand U3098 (N_3098,N_949,N_55);
and U3099 (N_3099,N_1699,N_902);
nand U3100 (N_3100,N_1325,N_1770);
nor U3101 (N_3101,N_1334,N_2004);
nand U3102 (N_3102,N_454,N_353);
nor U3103 (N_3103,N_358,N_1947);
nand U3104 (N_3104,N_536,N_1681);
nor U3105 (N_3105,N_1522,N_442);
nor U3106 (N_3106,N_2088,N_2226);
or U3107 (N_3107,N_1545,N_1598);
nand U3108 (N_3108,N_1026,N_937);
nand U3109 (N_3109,N_1520,N_951);
nand U3110 (N_3110,N_2320,N_1209);
nor U3111 (N_3111,N_667,N_605);
nor U3112 (N_3112,N_87,N_1707);
and U3113 (N_3113,N_1608,N_2277);
and U3114 (N_3114,N_1761,N_947);
or U3115 (N_3115,N_921,N_2156);
nand U3116 (N_3116,N_1047,N_727);
nor U3117 (N_3117,N_1895,N_2021);
xnor U3118 (N_3118,N_838,N_1537);
and U3119 (N_3119,N_1890,N_1956);
and U3120 (N_3120,N_504,N_1887);
and U3121 (N_3121,N_2345,N_508);
nand U3122 (N_3122,N_366,N_2253);
and U3123 (N_3123,N_1662,N_154);
nand U3124 (N_3124,N_884,N_640);
nor U3125 (N_3125,N_2153,N_1094);
and U3126 (N_3126,N_2100,N_690);
or U3127 (N_3127,N_348,N_1772);
xnor U3128 (N_3128,N_98,N_1131);
and U3129 (N_3129,N_1368,N_1777);
and U3130 (N_3130,N_1838,N_304);
nand U3131 (N_3131,N_431,N_2486);
and U3132 (N_3132,N_2390,N_679);
nand U3133 (N_3133,N_193,N_1356);
nor U3134 (N_3134,N_1475,N_45);
or U3135 (N_3135,N_1996,N_945);
or U3136 (N_3136,N_1987,N_2216);
or U3137 (N_3137,N_869,N_340);
and U3138 (N_3138,N_496,N_555);
nand U3139 (N_3139,N_1832,N_279);
nor U3140 (N_3140,N_124,N_369);
or U3141 (N_3141,N_954,N_1692);
nand U3142 (N_3142,N_244,N_1480);
or U3143 (N_3143,N_1869,N_1891);
xor U3144 (N_3144,N_1682,N_567);
or U3145 (N_3145,N_1219,N_1432);
or U3146 (N_3146,N_2463,N_1705);
nand U3147 (N_3147,N_714,N_2059);
or U3148 (N_3148,N_2352,N_1039);
and U3149 (N_3149,N_1892,N_2241);
or U3150 (N_3150,N_946,N_766);
nor U3151 (N_3151,N_1143,N_1431);
and U3152 (N_3152,N_409,N_2186);
and U3153 (N_3153,N_1073,N_526);
nand U3154 (N_3154,N_1798,N_1530);
nor U3155 (N_3155,N_984,N_37);
or U3156 (N_3156,N_837,N_88);
nor U3157 (N_3157,N_484,N_669);
nor U3158 (N_3158,N_1183,N_854);
or U3159 (N_3159,N_528,N_1390);
nand U3160 (N_3160,N_1976,N_101);
or U3161 (N_3161,N_943,N_2005);
nand U3162 (N_3162,N_865,N_2063);
nor U3163 (N_3163,N_1394,N_190);
or U3164 (N_3164,N_474,N_1854);
and U3165 (N_3165,N_891,N_1365);
and U3166 (N_3166,N_617,N_888);
nand U3167 (N_3167,N_455,N_1273);
or U3168 (N_3168,N_1166,N_1519);
nand U3169 (N_3169,N_2389,N_2038);
nor U3170 (N_3170,N_960,N_1720);
or U3171 (N_3171,N_470,N_704);
nand U3172 (N_3172,N_784,N_2300);
nor U3173 (N_3173,N_1347,N_1622);
and U3174 (N_3174,N_519,N_314);
nand U3175 (N_3175,N_621,N_302);
or U3176 (N_3176,N_290,N_1579);
and U3177 (N_3177,N_1569,N_2065);
and U3178 (N_3178,N_1805,N_613);
or U3179 (N_3179,N_980,N_2355);
or U3180 (N_3180,N_1458,N_29);
or U3181 (N_3181,N_120,N_1540);
xor U3182 (N_3182,N_1909,N_697);
nor U3183 (N_3183,N_1518,N_278);
and U3184 (N_3184,N_231,N_1042);
nor U3185 (N_3185,N_2311,N_2054);
xnor U3186 (N_3186,N_1844,N_739);
or U3187 (N_3187,N_450,N_2212);
nor U3188 (N_3188,N_476,N_194);
or U3189 (N_3189,N_2308,N_2409);
or U3190 (N_3190,N_1544,N_309);
or U3191 (N_3191,N_1491,N_978);
or U3192 (N_3192,N_466,N_1466);
nand U3193 (N_3193,N_1851,N_848);
nand U3194 (N_3194,N_1411,N_343);
nand U3195 (N_3195,N_1803,N_2344);
nand U3196 (N_3196,N_1445,N_2459);
and U3197 (N_3197,N_1488,N_561);
or U3198 (N_3198,N_925,N_2123);
nor U3199 (N_3199,N_1196,N_586);
and U3200 (N_3200,N_2043,N_781);
or U3201 (N_3201,N_1659,N_1113);
nor U3202 (N_3202,N_855,N_761);
nor U3203 (N_3203,N_1231,N_1207);
or U3204 (N_3204,N_1750,N_2234);
and U3205 (N_3205,N_661,N_147);
xor U3206 (N_3206,N_1669,N_790);
nor U3207 (N_3207,N_512,N_815);
and U3208 (N_3208,N_1292,N_407);
and U3209 (N_3209,N_2397,N_2184);
nand U3210 (N_3210,N_1261,N_2309);
or U3211 (N_3211,N_1464,N_557);
or U3212 (N_3212,N_1656,N_2252);
or U3213 (N_3213,N_390,N_554);
nand U3214 (N_3214,N_2256,N_1741);
xnor U3215 (N_3215,N_439,N_584);
nor U3216 (N_3216,N_1736,N_108);
and U3217 (N_3217,N_1771,N_1127);
xor U3218 (N_3218,N_2142,N_1420);
or U3219 (N_3219,N_1814,N_163);
or U3220 (N_3220,N_2268,N_2168);
nor U3221 (N_3221,N_2375,N_1973);
nor U3222 (N_3222,N_115,N_2251);
nand U3223 (N_3223,N_1369,N_1824);
nand U3224 (N_3224,N_2159,N_451);
nand U3225 (N_3225,N_1831,N_1760);
nor U3226 (N_3226,N_887,N_1133);
or U3227 (N_3227,N_1108,N_1019);
nor U3228 (N_3228,N_1262,N_393);
or U3229 (N_3229,N_2057,N_1934);
nor U3230 (N_3230,N_1187,N_993);
nor U3231 (N_3231,N_2453,N_1386);
nor U3232 (N_3232,N_2130,N_1957);
or U3233 (N_3233,N_441,N_1893);
and U3234 (N_3234,N_306,N_737);
and U3235 (N_3235,N_262,N_2002);
and U3236 (N_3236,N_1186,N_1605);
or U3237 (N_3237,N_2221,N_1348);
or U3238 (N_3238,N_1910,N_2086);
nand U3239 (N_3239,N_1470,N_1277);
nor U3240 (N_3240,N_171,N_709);
and U3241 (N_3241,N_576,N_1550);
and U3242 (N_3242,N_1958,N_1329);
or U3243 (N_3243,N_1905,N_2237);
or U3244 (N_3244,N_1258,N_1517);
nand U3245 (N_3245,N_1174,N_387);
nand U3246 (N_3246,N_1237,N_957);
and U3247 (N_3247,N_2299,N_2171);
or U3248 (N_3248,N_862,N_1264);
nor U3249 (N_3249,N_2444,N_1991);
nor U3250 (N_3250,N_1300,N_1921);
nor U3251 (N_3251,N_1224,N_203);
or U3252 (N_3252,N_685,N_777);
nor U3253 (N_3253,N_81,N_729);
nand U3254 (N_3254,N_2273,N_1215);
xor U3255 (N_3255,N_1043,N_1444);
nand U3256 (N_3256,N_1787,N_2332);
nor U3257 (N_3257,N_657,N_2497);
nor U3258 (N_3258,N_956,N_527);
or U3259 (N_3259,N_629,N_1293);
and U3260 (N_3260,N_15,N_372);
xor U3261 (N_3261,N_587,N_2101);
or U3262 (N_3262,N_646,N_2098);
or U3263 (N_3263,N_2116,N_2421);
nand U3264 (N_3264,N_871,N_1062);
nor U3265 (N_3265,N_481,N_560);
nand U3266 (N_3266,N_2410,N_2058);
nor U3267 (N_3267,N_2446,N_499);
or U3268 (N_3268,N_255,N_2238);
or U3269 (N_3269,N_2480,N_149);
xor U3270 (N_3270,N_139,N_220);
or U3271 (N_3271,N_877,N_1252);
or U3272 (N_3272,N_2442,N_991);
nor U3273 (N_3273,N_148,N_660);
nand U3274 (N_3274,N_1483,N_294);
and U3275 (N_3275,N_2246,N_2482);
or U3276 (N_3276,N_966,N_1558);
xor U3277 (N_3277,N_831,N_376);
nor U3278 (N_3278,N_539,N_1188);
or U3279 (N_3279,N_1609,N_312);
or U3280 (N_3280,N_543,N_1059);
nand U3281 (N_3281,N_1932,N_740);
or U3282 (N_3282,N_1693,N_1446);
and U3283 (N_3283,N_1376,N_1650);
and U3284 (N_3284,N_2342,N_2082);
or U3285 (N_3285,N_1942,N_2046);
and U3286 (N_3286,N_59,N_1307);
and U3287 (N_3287,N_1940,N_420);
nor U3288 (N_3288,N_1032,N_1213);
and U3289 (N_3289,N_1793,N_1013);
nand U3290 (N_3290,N_1415,N_313);
or U3291 (N_3291,N_858,N_1190);
nor U3292 (N_3292,N_362,N_1645);
nor U3293 (N_3293,N_907,N_1856);
nand U3294 (N_3294,N_1076,N_1602);
nand U3295 (N_3295,N_1402,N_1606);
nor U3296 (N_3296,N_678,N_103);
and U3297 (N_3297,N_264,N_1944);
or U3298 (N_3298,N_1045,N_216);
and U3299 (N_3299,N_821,N_520);
nand U3300 (N_3300,N_2485,N_509);
and U3301 (N_3301,N_1734,N_1898);
or U3302 (N_3302,N_351,N_791);
and U3303 (N_3303,N_1004,N_2010);
nor U3304 (N_3304,N_1901,N_1690);
nor U3305 (N_3305,N_581,N_114);
or U3306 (N_3306,N_762,N_448);
nand U3307 (N_3307,N_2454,N_2478);
and U3308 (N_3308,N_1457,N_832);
nor U3309 (N_3309,N_2405,N_2093);
or U3310 (N_3310,N_1000,N_2460);
and U3311 (N_3311,N_189,N_940);
nand U3312 (N_3312,N_1829,N_2208);
or U3313 (N_3313,N_1137,N_1984);
nand U3314 (N_3314,N_2437,N_551);
nand U3315 (N_3315,N_2182,N_797);
and U3316 (N_3316,N_734,N_1257);
or U3317 (N_3317,N_1911,N_129);
nand U3318 (N_3318,N_137,N_471);
and U3319 (N_3319,N_1284,N_706);
xor U3320 (N_3320,N_161,N_648);
nand U3321 (N_3321,N_2411,N_338);
nand U3322 (N_3322,N_283,N_977);
or U3323 (N_3323,N_1992,N_1904);
or U3324 (N_3324,N_187,N_1217);
or U3325 (N_3325,N_1240,N_300);
or U3326 (N_3326,N_2181,N_767);
or U3327 (N_3327,N_1572,N_2376);
nand U3328 (N_3328,N_1260,N_1995);
and U3329 (N_3329,N_1708,N_247);
nand U3330 (N_3330,N_2048,N_1534);
nor U3331 (N_3331,N_719,N_2015);
nor U3332 (N_3332,N_1389,N_173);
nor U3333 (N_3333,N_688,N_2477);
nor U3334 (N_3334,N_1698,N_2037);
and U3335 (N_3335,N_1363,N_488);
xnor U3336 (N_3336,N_1933,N_2077);
and U3337 (N_3337,N_1197,N_2370);
or U3338 (N_3338,N_452,N_778);
or U3339 (N_3339,N_1434,N_1259);
and U3340 (N_3340,N_1132,N_227);
nor U3341 (N_3341,N_1271,N_2080);
xnor U3342 (N_3342,N_633,N_1782);
and U3343 (N_3343,N_630,N_1919);
nand U3344 (N_3344,N_2034,N_1286);
and U3345 (N_3345,N_2090,N_153);
or U3346 (N_3346,N_224,N_2056);
nand U3347 (N_3347,N_1450,N_890);
and U3348 (N_3348,N_377,N_873);
nand U3349 (N_3349,N_1289,N_1270);
nor U3350 (N_3350,N_16,N_2062);
or U3351 (N_3351,N_145,N_1437);
or U3352 (N_3352,N_666,N_2371);
nand U3353 (N_3353,N_192,N_856);
and U3354 (N_3354,N_604,N_533);
nand U3355 (N_3355,N_2488,N_69);
and U3356 (N_3356,N_1439,N_1646);
nor U3357 (N_3357,N_578,N_1079);
nand U3358 (N_3358,N_684,N_1737);
or U3359 (N_3359,N_347,N_647);
nor U3360 (N_3360,N_364,N_2198);
and U3361 (N_3361,N_1161,N_2206);
and U3362 (N_3362,N_2136,N_1336);
nand U3363 (N_3363,N_1954,N_1651);
and U3364 (N_3364,N_1352,N_2386);
and U3365 (N_3365,N_1396,N_38);
nor U3366 (N_3366,N_1757,N_2395);
nor U3367 (N_3367,N_506,N_2078);
or U3368 (N_3368,N_1928,N_274);
and U3369 (N_3369,N_1641,N_1401);
or U3370 (N_3370,N_285,N_1370);
xnor U3371 (N_3371,N_1114,N_1601);
and U3372 (N_3372,N_2187,N_1441);
nand U3373 (N_3373,N_970,N_1276);
or U3374 (N_3374,N_234,N_847);
nand U3375 (N_3375,N_1462,N_1620);
and U3376 (N_3376,N_1647,N_1184);
and U3377 (N_3377,N_1003,N_2333);
nor U3378 (N_3378,N_1945,N_1603);
nand U3379 (N_3379,N_68,N_65);
nor U3380 (N_3380,N_1952,N_2270);
and U3381 (N_3381,N_1084,N_48);
or U3382 (N_3382,N_24,N_2429);
nand U3383 (N_3383,N_23,N_1126);
and U3384 (N_3384,N_802,N_2061);
nand U3385 (N_3385,N_415,N_1090);
nand U3386 (N_3386,N_2146,N_3);
or U3387 (N_3387,N_404,N_2027);
nand U3388 (N_3388,N_175,N_2294);
nor U3389 (N_3389,N_1227,N_1218);
and U3390 (N_3390,N_542,N_1704);
and U3391 (N_3391,N_2071,N_497);
or U3392 (N_3392,N_2326,N_840);
and U3393 (N_3393,N_559,N_1675);
nand U3394 (N_3394,N_2301,N_2447);
nand U3395 (N_3395,N_135,N_1776);
xor U3396 (N_3396,N_2173,N_916);
xor U3397 (N_3397,N_257,N_303);
or U3398 (N_3398,N_345,N_1101);
and U3399 (N_3399,N_792,N_1007);
and U3400 (N_3400,N_1341,N_2009);
or U3401 (N_3401,N_1236,N_1181);
or U3402 (N_3402,N_1098,N_2324);
xor U3403 (N_3403,N_774,N_1539);
and U3404 (N_3404,N_1862,N_493);
and U3405 (N_3405,N_583,N_879);
or U3406 (N_3406,N_990,N_710);
or U3407 (N_3407,N_2433,N_736);
and U3408 (N_3408,N_563,N_2106);
and U3409 (N_3409,N_1247,N_0);
nor U3410 (N_3410,N_677,N_517);
and U3411 (N_3411,N_1671,N_638);
and U3412 (N_3412,N_553,N_2282);
nor U3413 (N_3413,N_316,N_150);
xnor U3414 (N_3414,N_33,N_464);
nor U3415 (N_3415,N_494,N_1056);
or U3416 (N_3416,N_1806,N_2493);
and U3417 (N_3417,N_986,N_177);
nor U3418 (N_3418,N_1663,N_1833);
or U3419 (N_3419,N_1204,N_1747);
nor U3420 (N_3420,N_1565,N_2490);
nor U3421 (N_3421,N_237,N_2215);
xor U3422 (N_3422,N_1819,N_1392);
nand U3423 (N_3423,N_2200,N_1139);
or U3424 (N_3424,N_1709,N_2030);
or U3425 (N_3425,N_972,N_671);
and U3426 (N_3426,N_1173,N_1195);
nor U3427 (N_3427,N_1182,N_1562);
nor U3428 (N_3428,N_1087,N_460);
xnor U3429 (N_3429,N_1538,N_843);
nor U3430 (N_3430,N_608,N_1532);
or U3431 (N_3431,N_1448,N_382);
nor U3432 (N_3432,N_1785,N_2129);
nor U3433 (N_3433,N_2245,N_1050);
or U3434 (N_3434,N_2329,N_566);
nor U3435 (N_3435,N_269,N_1828);
nand U3436 (N_3436,N_2280,N_701);
nor U3437 (N_3437,N_292,N_1189);
and U3438 (N_3438,N_682,N_530);
xnor U3439 (N_3439,N_1036,N_1111);
and U3440 (N_3440,N_967,N_963);
and U3441 (N_3441,N_1999,N_2422);
nand U3442 (N_3442,N_1716,N_2383);
nand U3443 (N_3443,N_288,N_2134);
or U3444 (N_3444,N_272,N_144);
nand U3445 (N_3445,N_105,N_125);
or U3446 (N_3446,N_416,N_793);
or U3447 (N_3447,N_502,N_702);
and U3448 (N_3448,N_523,N_1216);
nor U3449 (N_3449,N_1409,N_2432);
nor U3450 (N_3450,N_388,N_1794);
nand U3451 (N_3451,N_1925,N_911);
and U3452 (N_3452,N_2220,N_1764);
and U3453 (N_3453,N_1070,N_1912);
or U3454 (N_3454,N_2149,N_1302);
and U3455 (N_3455,N_1384,N_1353);
nor U3456 (N_3456,N_14,N_1038);
nand U3457 (N_3457,N_788,N_735);
or U3458 (N_3458,N_1121,N_829);
or U3459 (N_3459,N_615,N_179);
or U3460 (N_3460,N_643,N_17);
or U3461 (N_3461,N_1676,N_1584);
nand U3462 (N_3462,N_2177,N_2465);
and U3463 (N_3463,N_573,N_1786);
nand U3464 (N_3464,N_395,N_1859);
nand U3465 (N_3465,N_1244,N_222);
nand U3466 (N_3466,N_720,N_1701);
or U3467 (N_3467,N_2343,N_223);
or U3468 (N_3468,N_696,N_427);
or U3469 (N_3469,N_472,N_254);
and U3470 (N_3470,N_2498,N_1055);
or U3471 (N_3471,N_2458,N_1816);
nand U3472 (N_3472,N_1955,N_1478);
nand U3473 (N_3473,N_1721,N_2284);
or U3474 (N_3474,N_600,N_2041);
or U3475 (N_3475,N_296,N_1308);
nand U3476 (N_3476,N_2484,N_1637);
nor U3477 (N_3477,N_2398,N_308);
and U3478 (N_3478,N_1135,N_1053);
or U3479 (N_3479,N_2254,N_1959);
and U3480 (N_3480,N_1072,N_1200);
nand U3481 (N_3481,N_883,N_64);
nand U3482 (N_3482,N_1226,N_1845);
or U3483 (N_3483,N_1843,N_813);
nor U3484 (N_3484,N_2115,N_2001);
and U3485 (N_3485,N_1361,N_962);
and U3486 (N_3486,N_1900,N_738);
nand U3487 (N_3487,N_1010,N_2074);
nand U3488 (N_3488,N_2120,N_323);
or U3489 (N_3489,N_808,N_2334);
and U3490 (N_3490,N_1822,N_13);
nand U3491 (N_3491,N_2378,N_603);
and U3492 (N_3492,N_1316,N_1250);
nor U3493 (N_3493,N_2079,N_2257);
and U3494 (N_3494,N_2448,N_501);
or U3495 (N_3495,N_1400,N_742);
nor U3496 (N_3496,N_860,N_634);
nor U3497 (N_3497,N_1636,N_2321);
and U3498 (N_3498,N_1089,N_261);
nor U3499 (N_3499,N_178,N_1593);
nor U3500 (N_3500,N_1813,N_21);
or U3501 (N_3501,N_78,N_2361);
nand U3502 (N_3502,N_1080,N_2229);
and U3503 (N_3503,N_920,N_914);
nor U3504 (N_3504,N_381,N_591);
nor U3505 (N_3505,N_757,N_1670);
nand U3506 (N_3506,N_2174,N_498);
nand U3507 (N_3507,N_1176,N_1379);
and U3508 (N_3508,N_155,N_1521);
or U3509 (N_3509,N_2210,N_1165);
nor U3510 (N_3510,N_1547,N_440);
and U3511 (N_3511,N_868,N_1746);
nand U3512 (N_3512,N_479,N_483);
and U3513 (N_3513,N_1242,N_2013);
or U3514 (N_3514,N_482,N_935);
or U3515 (N_3515,N_436,N_2279);
nand U3516 (N_3516,N_1768,N_5);
or U3517 (N_3517,N_1024,N_1473);
nand U3518 (N_3518,N_489,N_1568);
and U3519 (N_3519,N_2407,N_1067);
nand U3520 (N_3520,N_1549,N_2424);
and U3521 (N_3521,N_1429,N_2255);
and U3522 (N_3522,N_1570,N_385);
or U3523 (N_3523,N_1099,N_619);
nor U3524 (N_3524,N_383,N_293);
nor U3525 (N_3525,N_2040,N_1555);
and U3526 (N_3526,N_391,N_1567);
and U3527 (N_3527,N_510,N_1349);
nand U3528 (N_3528,N_929,N_939);
and U3529 (N_3529,N_151,N_1564);
or U3530 (N_3530,N_1320,N_1279);
nor U3531 (N_3531,N_721,N_2012);
or U3532 (N_3532,N_1994,N_1029);
nor U3533 (N_3533,N_1586,N_107);
and U3534 (N_3534,N_834,N_12);
nor U3535 (N_3535,N_1313,N_572);
nor U3536 (N_3536,N_1774,N_776);
nor U3537 (N_3537,N_1874,N_1638);
and U3538 (N_3538,N_964,N_1225);
nor U3539 (N_3539,N_732,N_1566);
and U3540 (N_3540,N_1459,N_330);
and U3541 (N_3541,N_1238,N_1091);
or U3542 (N_3542,N_1894,N_592);
and U3543 (N_3543,N_1535,N_1621);
or U3544 (N_3544,N_1314,N_104);
nor U3545 (N_3545,N_924,N_1718);
nand U3546 (N_3546,N_1413,N_160);
nand U3547 (N_3547,N_2113,N_546);
nor U3548 (N_3548,N_1106,N_1745);
and U3549 (N_3549,N_253,N_779);
or U3550 (N_3550,N_1811,N_1930);
and U3551 (N_3551,N_218,N_1134);
or U3552 (N_3552,N_1430,N_1203);
nand U3553 (N_3553,N_2261,N_803);
or U3554 (N_3554,N_1936,N_1546);
nor U3555 (N_3555,N_52,N_2452);
nor U3556 (N_3556,N_852,N_1296);
nand U3557 (N_3557,N_20,N_2451);
nand U3558 (N_3558,N_80,N_1107);
nor U3559 (N_3559,N_953,N_801);
nand U3560 (N_3560,N_344,N_894);
nand U3561 (N_3561,N_1835,N_1438);
nor U3562 (N_3562,N_1778,N_396);
and U3563 (N_3563,N_594,N_417);
nand U3564 (N_3564,N_2188,N_558);
or U3565 (N_3565,N_1138,N_641);
nand U3566 (N_3566,N_22,N_2428);
and U3567 (N_3567,N_1685,N_1714);
nor U3568 (N_3568,N_1823,N_1654);
nand U3569 (N_3569,N_1093,N_1897);
nor U3570 (N_3570,N_1461,N_2095);
and U3571 (N_3571,N_2042,N_768);
nand U3572 (N_3572,N_1315,N_1248);
nor U3573 (N_3573,N_1561,N_989);
nand U3574 (N_3574,N_745,N_1951);
nor U3575 (N_3575,N_754,N_6);
nor U3576 (N_3576,N_321,N_1792);
and U3577 (N_3577,N_1553,N_9);
or U3578 (N_3578,N_67,N_662);
nor U3579 (N_3579,N_2060,N_1514);
nor U3580 (N_3580,N_1310,N_723);
nand U3581 (N_3581,N_1938,N_886);
nand U3582 (N_3582,N_703,N_507);
nand U3583 (N_3583,N_1860,N_2202);
and U3584 (N_3584,N_1505,N_1102);
nand U3585 (N_3585,N_208,N_2382);
nand U3586 (N_3586,N_2295,N_841);
nor U3587 (N_3587,N_298,N_1907);
nor U3588 (N_3588,N_1830,N_590);
nor U3589 (N_3589,N_1044,N_503);
nor U3590 (N_3590,N_955,N_1120);
nor U3591 (N_3591,N_1421,N_2214);
or U3592 (N_3592,N_981,N_1610);
and U3593 (N_3593,N_1506,N_1330);
nor U3594 (N_3594,N_823,N_538);
or U3595 (N_3595,N_2091,N_226);
nor U3596 (N_3596,N_2169,N_2350);
nand U3597 (N_3597,N_1642,N_1239);
or U3598 (N_3598,N_988,N_468);
nor U3599 (N_3599,N_1541,N_2050);
and U3600 (N_3600,N_1486,N_1668);
and U3601 (N_3601,N_1665,N_2357);
nand U3602 (N_3602,N_618,N_824);
nand U3603 (N_3603,N_329,N_812);
nand U3604 (N_3604,N_789,N_505);
nor U3605 (N_3605,N_209,N_2379);
nor U3606 (N_3606,N_637,N_1263);
or U3607 (N_3607,N_200,N_240);
or U3608 (N_3608,N_571,N_752);
or U3609 (N_3609,N_950,N_1245);
nor U3610 (N_3610,N_1592,N_430);
or U3611 (N_3611,N_1563,N_2154);
or U3612 (N_3612,N_1739,N_1246);
nor U3613 (N_3613,N_903,N_1649);
nor U3614 (N_3614,N_1193,N_1943);
nand U3615 (N_3615,N_1578,N_400);
nand U3616 (N_3616,N_133,N_206);
or U3617 (N_3617,N_1585,N_635);
nand U3618 (N_3618,N_1784,N_2128);
nand U3619 (N_3619,N_1020,N_1501);
nor U3620 (N_3620,N_332,N_233);
nand U3621 (N_3621,N_2244,N_94);
and U3622 (N_3622,N_1630,N_2178);
and U3623 (N_3623,N_1766,N_644);
or U3624 (N_3624,N_1686,N_625);
and U3625 (N_3625,N_2164,N_1049);
or U3626 (N_3626,N_1949,N_1065);
and U3627 (N_3627,N_1531,N_2487);
nand U3628 (N_3628,N_1790,N_1110);
nor U3629 (N_3629,N_1164,N_401);
nor U3630 (N_3630,N_106,N_1613);
nand U3631 (N_3631,N_532,N_1914);
or U3632 (N_3632,N_397,N_492);
and U3633 (N_3633,N_97,N_433);
or U3634 (N_3634,N_1526,N_1903);
and U3635 (N_3635,N_215,N_1066);
and U3636 (N_3636,N_1141,N_700);
and U3637 (N_3637,N_2351,N_117);
or U3638 (N_3638,N_751,N_1527);
or U3639 (N_3639,N_1679,N_1123);
and U3640 (N_3640,N_2457,N_1192);
nand U3641 (N_3641,N_168,N_1775);
nor U3642 (N_3642,N_2417,N_1631);
xor U3643 (N_3643,N_2469,N_143);
nand U3644 (N_3644,N_2075,N_1433);
nor U3645 (N_3645,N_1145,N_1837);
nor U3646 (N_3646,N_1858,N_1500);
or U3647 (N_3647,N_457,N_2144);
and U3648 (N_3648,N_589,N_1220);
xnor U3649 (N_3649,N_1380,N_185);
or U3650 (N_3650,N_1614,N_1170);
and U3651 (N_3651,N_73,N_2225);
nor U3652 (N_3652,N_1552,N_118);
xor U3653 (N_3653,N_997,N_74);
and U3654 (N_3654,N_826,N_1915);
and U3655 (N_3655,N_1169,N_334);
and U3656 (N_3656,N_456,N_1175);
or U3657 (N_3657,N_1199,N_1694);
or U3658 (N_3658,N_775,N_728);
nor U3659 (N_3659,N_1472,N_1156);
nor U3660 (N_3660,N_403,N_320);
or U3661 (N_3661,N_7,N_1168);
or U3662 (N_3662,N_2084,N_2312);
nor U3663 (N_3663,N_1616,N_1626);
and U3664 (N_3664,N_311,N_675);
nand U3665 (N_3665,N_1881,N_1719);
or U3666 (N_3666,N_1826,N_1617);
nor U3667 (N_3667,N_1972,N_691);
nand U3668 (N_3668,N_1953,N_994);
nand U3669 (N_3669,N_653,N_2143);
xnor U3670 (N_3670,N_1908,N_1931);
nand U3671 (N_3671,N_2087,N_1725);
or U3672 (N_3672,N_722,N_1060);
or U3673 (N_3673,N_537,N_425);
or U3674 (N_3674,N_772,N_649);
nor U3675 (N_3675,N_2118,N_606);
xnor U3676 (N_3676,N_57,N_1054);
and U3677 (N_3677,N_389,N_1735);
nor U3678 (N_3678,N_197,N_1232);
or U3679 (N_3679,N_908,N_1963);
or U3680 (N_3680,N_1452,N_1295);
nand U3681 (N_3681,N_610,N_1700);
or U3682 (N_3682,N_1311,N_25);
xor U3683 (N_3683,N_1968,N_423);
and U3684 (N_3684,N_670,N_901);
nor U3685 (N_3685,N_243,N_747);
nor U3686 (N_3686,N_534,N_1435);
and U3687 (N_3687,N_1357,N_2439);
and U3688 (N_3688,N_195,N_2462);
nand U3689 (N_3689,N_918,N_1975);
nor U3690 (N_3690,N_1210,N_2362);
nand U3691 (N_3691,N_1639,N_2440);
nor U3692 (N_3692,N_1756,N_336);
nand U3693 (N_3693,N_1667,N_659);
or U3694 (N_3694,N_698,N_1974);
and U3695 (N_3695,N_126,N_897);
nand U3696 (N_3696,N_1962,N_128);
or U3697 (N_3697,N_2266,N_47);
nor U3698 (N_3698,N_2047,N_2358);
and U3699 (N_3699,N_1581,N_1487);
and U3700 (N_3700,N_2243,N_1657);
and U3701 (N_3701,N_1827,N_895);
nand U3702 (N_3702,N_1088,N_110);
xor U3703 (N_3703,N_2450,N_2081);
or U3704 (N_3704,N_1027,N_1576);
nor U3705 (N_3705,N_217,N_1711);
and U3706 (N_3706,N_1961,N_2275);
and U3707 (N_3707,N_2495,N_1985);
nor U3708 (N_3708,N_2076,N_109);
nor U3709 (N_3709,N_541,N_1847);
nor U3710 (N_3710,N_1069,N_10);
or U3711 (N_3711,N_1724,N_1228);
nand U3712 (N_3712,N_2325,N_256);
nor U3713 (N_3713,N_1476,N_2420);
xnor U3714 (N_3714,N_287,N_43);
and U3715 (N_3715,N_1779,N_2492);
nand U3716 (N_3716,N_167,N_2124);
or U3717 (N_3717,N_2466,N_183);
and U3718 (N_3718,N_1981,N_1022);
or U3719 (N_3719,N_201,N_2195);
or U3720 (N_3720,N_241,N_896);
nor U3721 (N_3721,N_191,N_1498);
and U3722 (N_3722,N_112,N_1926);
nand U3723 (N_3723,N_1211,N_1533);
or U3724 (N_3724,N_174,N_1967);
nand U3725 (N_3725,N_2231,N_2064);
or U3726 (N_3726,N_680,N_1014);
nor U3727 (N_3727,N_2092,N_1988);
nor U3728 (N_3728,N_1946,N_2470);
or U3729 (N_3729,N_1075,N_2292);
nand U3730 (N_3730,N_280,N_1344);
nor U3731 (N_3731,N_976,N_325);
nand U3732 (N_3732,N_1818,N_463);
nor U3733 (N_3733,N_626,N_1104);
nand U3734 (N_3734,N_449,N_1016);
xor U3735 (N_3735,N_443,N_2408);
or U3736 (N_3736,N_1513,N_1710);
nor U3737 (N_3737,N_123,N_251);
nor U3738 (N_3738,N_1733,N_1011);
or U3739 (N_3739,N_337,N_335);
and U3740 (N_3740,N_1456,N_2475);
nor U3741 (N_3741,N_1809,N_2413);
or U3742 (N_3742,N_2377,N_1590);
nor U3743 (N_3743,N_1917,N_2196);
nor U3744 (N_3744,N_1767,N_1304);
or U3745 (N_3745,N_1496,N_249);
or U3746 (N_3746,N_798,N_1142);
and U3747 (N_3747,N_1817,N_1077);
or U3748 (N_3748,N_1684,N_2197);
or U3749 (N_3749,N_491,N_833);
nand U3750 (N_3750,N_1438,N_2360);
nor U3751 (N_3751,N_1446,N_313);
and U3752 (N_3752,N_61,N_2481);
nor U3753 (N_3753,N_132,N_701);
and U3754 (N_3754,N_1146,N_1216);
or U3755 (N_3755,N_2235,N_2454);
nand U3756 (N_3756,N_924,N_308);
nand U3757 (N_3757,N_1779,N_668);
nor U3758 (N_3758,N_341,N_1544);
xnor U3759 (N_3759,N_1944,N_1841);
nor U3760 (N_3760,N_687,N_1912);
nor U3761 (N_3761,N_1713,N_1197);
or U3762 (N_3762,N_2324,N_478);
nand U3763 (N_3763,N_796,N_1055);
nor U3764 (N_3764,N_209,N_1617);
nor U3765 (N_3765,N_2229,N_1547);
and U3766 (N_3766,N_657,N_2019);
and U3767 (N_3767,N_777,N_2119);
or U3768 (N_3768,N_1684,N_491);
nand U3769 (N_3769,N_352,N_462);
and U3770 (N_3770,N_1930,N_2364);
or U3771 (N_3771,N_983,N_602);
xnor U3772 (N_3772,N_996,N_1684);
nand U3773 (N_3773,N_690,N_2353);
nand U3774 (N_3774,N_1457,N_1887);
nor U3775 (N_3775,N_2134,N_1619);
and U3776 (N_3776,N_965,N_1929);
or U3777 (N_3777,N_1776,N_1991);
and U3778 (N_3778,N_785,N_1962);
nor U3779 (N_3779,N_662,N_2411);
nand U3780 (N_3780,N_385,N_674);
nand U3781 (N_3781,N_1252,N_2376);
and U3782 (N_3782,N_1808,N_1579);
and U3783 (N_3783,N_2410,N_2412);
nor U3784 (N_3784,N_2171,N_1382);
nand U3785 (N_3785,N_702,N_2306);
xor U3786 (N_3786,N_831,N_2253);
nor U3787 (N_3787,N_472,N_1718);
and U3788 (N_3788,N_1071,N_1650);
nor U3789 (N_3789,N_1999,N_1330);
nor U3790 (N_3790,N_670,N_2280);
nor U3791 (N_3791,N_1369,N_341);
and U3792 (N_3792,N_1076,N_907);
and U3793 (N_3793,N_635,N_99);
and U3794 (N_3794,N_846,N_1682);
nor U3795 (N_3795,N_1374,N_963);
nor U3796 (N_3796,N_921,N_677);
or U3797 (N_3797,N_1447,N_280);
nand U3798 (N_3798,N_1467,N_1403);
and U3799 (N_3799,N_1705,N_561);
and U3800 (N_3800,N_847,N_1325);
and U3801 (N_3801,N_336,N_283);
nor U3802 (N_3802,N_2102,N_2078);
xor U3803 (N_3803,N_1727,N_2262);
or U3804 (N_3804,N_609,N_2121);
and U3805 (N_3805,N_2001,N_490);
or U3806 (N_3806,N_1842,N_2077);
xor U3807 (N_3807,N_74,N_263);
or U3808 (N_3808,N_1638,N_1335);
or U3809 (N_3809,N_1079,N_2045);
and U3810 (N_3810,N_1413,N_1071);
nor U3811 (N_3811,N_1798,N_169);
and U3812 (N_3812,N_215,N_1450);
nand U3813 (N_3813,N_1035,N_1889);
and U3814 (N_3814,N_1819,N_1239);
and U3815 (N_3815,N_2292,N_2408);
or U3816 (N_3816,N_1673,N_1152);
nand U3817 (N_3817,N_72,N_1745);
nor U3818 (N_3818,N_1090,N_1564);
or U3819 (N_3819,N_249,N_1585);
and U3820 (N_3820,N_273,N_2347);
or U3821 (N_3821,N_2061,N_1230);
or U3822 (N_3822,N_2383,N_451);
or U3823 (N_3823,N_349,N_1341);
nor U3824 (N_3824,N_954,N_1964);
and U3825 (N_3825,N_275,N_1688);
nor U3826 (N_3826,N_1603,N_378);
or U3827 (N_3827,N_2029,N_1511);
nand U3828 (N_3828,N_2423,N_109);
nand U3829 (N_3829,N_1558,N_1722);
nand U3830 (N_3830,N_505,N_301);
or U3831 (N_3831,N_2149,N_37);
or U3832 (N_3832,N_528,N_1374);
and U3833 (N_3833,N_1562,N_1544);
and U3834 (N_3834,N_1436,N_961);
nor U3835 (N_3835,N_418,N_1983);
or U3836 (N_3836,N_1570,N_2016);
and U3837 (N_3837,N_1372,N_751);
nand U3838 (N_3838,N_1404,N_1018);
or U3839 (N_3839,N_2094,N_2044);
nor U3840 (N_3840,N_242,N_1604);
nand U3841 (N_3841,N_1751,N_1219);
nand U3842 (N_3842,N_614,N_2059);
nand U3843 (N_3843,N_397,N_1255);
nand U3844 (N_3844,N_295,N_2005);
and U3845 (N_3845,N_2388,N_951);
xnor U3846 (N_3846,N_76,N_1122);
nand U3847 (N_3847,N_516,N_1810);
and U3848 (N_3848,N_114,N_1595);
and U3849 (N_3849,N_10,N_1241);
xor U3850 (N_3850,N_1994,N_1845);
or U3851 (N_3851,N_1552,N_2001);
or U3852 (N_3852,N_2029,N_968);
nand U3853 (N_3853,N_445,N_1891);
and U3854 (N_3854,N_464,N_276);
or U3855 (N_3855,N_641,N_2062);
nand U3856 (N_3856,N_1709,N_1107);
and U3857 (N_3857,N_965,N_1448);
or U3858 (N_3858,N_931,N_862);
nand U3859 (N_3859,N_2484,N_2171);
or U3860 (N_3860,N_1805,N_1847);
nor U3861 (N_3861,N_629,N_738);
nand U3862 (N_3862,N_961,N_504);
and U3863 (N_3863,N_1727,N_1976);
nand U3864 (N_3864,N_224,N_1946);
nor U3865 (N_3865,N_2090,N_1699);
and U3866 (N_3866,N_128,N_1418);
nor U3867 (N_3867,N_1180,N_666);
nor U3868 (N_3868,N_524,N_745);
and U3869 (N_3869,N_859,N_2320);
nor U3870 (N_3870,N_1995,N_1854);
nand U3871 (N_3871,N_116,N_1452);
nand U3872 (N_3872,N_384,N_338);
nand U3873 (N_3873,N_1984,N_1951);
or U3874 (N_3874,N_735,N_173);
nand U3875 (N_3875,N_744,N_2322);
nor U3876 (N_3876,N_1854,N_845);
nand U3877 (N_3877,N_1062,N_1933);
nor U3878 (N_3878,N_1066,N_1463);
nor U3879 (N_3879,N_2449,N_1641);
xor U3880 (N_3880,N_1278,N_1536);
nand U3881 (N_3881,N_1272,N_857);
or U3882 (N_3882,N_1734,N_228);
or U3883 (N_3883,N_339,N_639);
nand U3884 (N_3884,N_688,N_1029);
nor U3885 (N_3885,N_1425,N_75);
or U3886 (N_3886,N_677,N_1546);
nand U3887 (N_3887,N_2495,N_2135);
and U3888 (N_3888,N_2380,N_1665);
nor U3889 (N_3889,N_211,N_392);
nand U3890 (N_3890,N_1937,N_855);
and U3891 (N_3891,N_1013,N_1755);
or U3892 (N_3892,N_670,N_200);
nand U3893 (N_3893,N_2023,N_1278);
nand U3894 (N_3894,N_1447,N_2141);
nor U3895 (N_3895,N_2018,N_2364);
nand U3896 (N_3896,N_295,N_1628);
nand U3897 (N_3897,N_498,N_2083);
and U3898 (N_3898,N_689,N_1585);
or U3899 (N_3899,N_859,N_1108);
xnor U3900 (N_3900,N_2040,N_969);
nand U3901 (N_3901,N_1170,N_2164);
nor U3902 (N_3902,N_1951,N_1098);
nor U3903 (N_3903,N_2460,N_2255);
or U3904 (N_3904,N_70,N_2158);
and U3905 (N_3905,N_759,N_1513);
nor U3906 (N_3906,N_1166,N_503);
nor U3907 (N_3907,N_867,N_2336);
and U3908 (N_3908,N_804,N_988);
nor U3909 (N_3909,N_1371,N_1832);
nor U3910 (N_3910,N_1301,N_809);
or U3911 (N_3911,N_241,N_1417);
nand U3912 (N_3912,N_1453,N_2496);
and U3913 (N_3913,N_1832,N_2204);
nor U3914 (N_3914,N_695,N_62);
nand U3915 (N_3915,N_1227,N_29);
nor U3916 (N_3916,N_41,N_2353);
or U3917 (N_3917,N_1564,N_1753);
nand U3918 (N_3918,N_7,N_1019);
nor U3919 (N_3919,N_837,N_1362);
and U3920 (N_3920,N_242,N_1378);
or U3921 (N_3921,N_1964,N_881);
nor U3922 (N_3922,N_472,N_2421);
nor U3923 (N_3923,N_1007,N_2308);
or U3924 (N_3924,N_189,N_10);
and U3925 (N_3925,N_1257,N_844);
nand U3926 (N_3926,N_2385,N_1263);
xor U3927 (N_3927,N_1185,N_2168);
nand U3928 (N_3928,N_1380,N_807);
or U3929 (N_3929,N_1723,N_1745);
or U3930 (N_3930,N_2242,N_1530);
nor U3931 (N_3931,N_1657,N_1158);
and U3932 (N_3932,N_179,N_1965);
nand U3933 (N_3933,N_822,N_2488);
and U3934 (N_3934,N_194,N_510);
nand U3935 (N_3935,N_11,N_920);
nand U3936 (N_3936,N_444,N_2483);
and U3937 (N_3937,N_1005,N_272);
nand U3938 (N_3938,N_1911,N_246);
and U3939 (N_3939,N_1186,N_506);
nand U3940 (N_3940,N_742,N_1851);
nor U3941 (N_3941,N_2049,N_1872);
and U3942 (N_3942,N_509,N_393);
or U3943 (N_3943,N_2204,N_826);
or U3944 (N_3944,N_1075,N_1569);
or U3945 (N_3945,N_794,N_1598);
nand U3946 (N_3946,N_1594,N_1128);
nand U3947 (N_3947,N_1402,N_2385);
nor U3948 (N_3948,N_912,N_980);
xnor U3949 (N_3949,N_717,N_2090);
and U3950 (N_3950,N_104,N_517);
and U3951 (N_3951,N_516,N_2335);
or U3952 (N_3952,N_1330,N_88);
or U3953 (N_3953,N_1950,N_875);
nand U3954 (N_3954,N_792,N_972);
nor U3955 (N_3955,N_2149,N_2041);
and U3956 (N_3956,N_348,N_445);
or U3957 (N_3957,N_881,N_346);
or U3958 (N_3958,N_2477,N_915);
nor U3959 (N_3959,N_2075,N_2149);
nand U3960 (N_3960,N_2276,N_1902);
nor U3961 (N_3961,N_1772,N_2146);
nor U3962 (N_3962,N_2238,N_1526);
or U3963 (N_3963,N_1003,N_983);
and U3964 (N_3964,N_406,N_1539);
or U3965 (N_3965,N_1885,N_159);
nor U3966 (N_3966,N_1118,N_1801);
or U3967 (N_3967,N_763,N_2174);
nor U3968 (N_3968,N_2449,N_715);
or U3969 (N_3969,N_882,N_1955);
or U3970 (N_3970,N_82,N_2179);
and U3971 (N_3971,N_2347,N_2282);
or U3972 (N_3972,N_2311,N_1108);
nand U3973 (N_3973,N_2459,N_1312);
and U3974 (N_3974,N_297,N_2471);
or U3975 (N_3975,N_2012,N_242);
nand U3976 (N_3976,N_415,N_888);
nor U3977 (N_3977,N_2162,N_1242);
or U3978 (N_3978,N_2290,N_2181);
nand U3979 (N_3979,N_776,N_2384);
or U3980 (N_3980,N_1075,N_1969);
or U3981 (N_3981,N_2418,N_1249);
nand U3982 (N_3982,N_245,N_351);
nor U3983 (N_3983,N_2191,N_1389);
nand U3984 (N_3984,N_1652,N_690);
xnor U3985 (N_3985,N_469,N_1464);
nand U3986 (N_3986,N_335,N_777);
or U3987 (N_3987,N_1454,N_1163);
nor U3988 (N_3988,N_910,N_911);
and U3989 (N_3989,N_1460,N_2056);
and U3990 (N_3990,N_535,N_1065);
and U3991 (N_3991,N_153,N_1908);
nor U3992 (N_3992,N_987,N_2075);
or U3993 (N_3993,N_1270,N_694);
or U3994 (N_3994,N_831,N_1334);
xnor U3995 (N_3995,N_2108,N_2384);
nor U3996 (N_3996,N_327,N_977);
or U3997 (N_3997,N_1435,N_1775);
nand U3998 (N_3998,N_1877,N_1988);
or U3999 (N_3999,N_754,N_1039);
and U4000 (N_4000,N_763,N_1337);
or U4001 (N_4001,N_111,N_2254);
or U4002 (N_4002,N_876,N_1751);
nand U4003 (N_4003,N_804,N_2022);
and U4004 (N_4004,N_2261,N_586);
nor U4005 (N_4005,N_477,N_1228);
and U4006 (N_4006,N_535,N_2039);
nor U4007 (N_4007,N_1324,N_14);
nand U4008 (N_4008,N_81,N_752);
and U4009 (N_4009,N_49,N_688);
or U4010 (N_4010,N_770,N_1755);
or U4011 (N_4011,N_1605,N_2178);
nand U4012 (N_4012,N_1785,N_1557);
nor U4013 (N_4013,N_26,N_977);
nand U4014 (N_4014,N_229,N_1281);
and U4015 (N_4015,N_565,N_1553);
or U4016 (N_4016,N_548,N_2312);
or U4017 (N_4017,N_991,N_2079);
xnor U4018 (N_4018,N_2352,N_1538);
nand U4019 (N_4019,N_1708,N_997);
or U4020 (N_4020,N_1067,N_486);
and U4021 (N_4021,N_1040,N_2161);
xnor U4022 (N_4022,N_930,N_1734);
and U4023 (N_4023,N_897,N_1112);
and U4024 (N_4024,N_160,N_943);
nor U4025 (N_4025,N_1011,N_2080);
nor U4026 (N_4026,N_1780,N_757);
or U4027 (N_4027,N_899,N_624);
xor U4028 (N_4028,N_684,N_1683);
nand U4029 (N_4029,N_913,N_842);
or U4030 (N_4030,N_244,N_679);
and U4031 (N_4031,N_136,N_1063);
and U4032 (N_4032,N_2282,N_776);
and U4033 (N_4033,N_52,N_1598);
or U4034 (N_4034,N_1344,N_1446);
nor U4035 (N_4035,N_345,N_1461);
nand U4036 (N_4036,N_50,N_1941);
nor U4037 (N_4037,N_1230,N_635);
and U4038 (N_4038,N_327,N_1554);
or U4039 (N_4039,N_1479,N_2335);
nand U4040 (N_4040,N_91,N_1893);
nor U4041 (N_4041,N_2474,N_215);
nand U4042 (N_4042,N_435,N_1379);
and U4043 (N_4043,N_553,N_310);
or U4044 (N_4044,N_46,N_2095);
or U4045 (N_4045,N_808,N_2022);
nor U4046 (N_4046,N_953,N_151);
and U4047 (N_4047,N_1159,N_1221);
nand U4048 (N_4048,N_1356,N_2285);
nand U4049 (N_4049,N_607,N_1635);
and U4050 (N_4050,N_1916,N_406);
nor U4051 (N_4051,N_2037,N_606);
nor U4052 (N_4052,N_704,N_57);
nand U4053 (N_4053,N_1567,N_2112);
nand U4054 (N_4054,N_2208,N_212);
and U4055 (N_4055,N_2356,N_1316);
or U4056 (N_4056,N_2201,N_347);
and U4057 (N_4057,N_967,N_560);
or U4058 (N_4058,N_1434,N_1166);
nor U4059 (N_4059,N_1117,N_93);
and U4060 (N_4060,N_2281,N_2277);
and U4061 (N_4061,N_2398,N_448);
nand U4062 (N_4062,N_2466,N_93);
or U4063 (N_4063,N_2289,N_536);
nor U4064 (N_4064,N_2239,N_1467);
nor U4065 (N_4065,N_2169,N_271);
nor U4066 (N_4066,N_859,N_1736);
nand U4067 (N_4067,N_955,N_1208);
or U4068 (N_4068,N_262,N_614);
or U4069 (N_4069,N_380,N_1275);
nand U4070 (N_4070,N_992,N_962);
xnor U4071 (N_4071,N_2315,N_217);
nor U4072 (N_4072,N_411,N_2374);
and U4073 (N_4073,N_2047,N_424);
or U4074 (N_4074,N_344,N_258);
nand U4075 (N_4075,N_473,N_1465);
and U4076 (N_4076,N_1081,N_1413);
nand U4077 (N_4077,N_1264,N_307);
xnor U4078 (N_4078,N_85,N_2408);
or U4079 (N_4079,N_2035,N_942);
and U4080 (N_4080,N_432,N_1173);
nor U4081 (N_4081,N_450,N_471);
and U4082 (N_4082,N_1194,N_1205);
nand U4083 (N_4083,N_1553,N_989);
or U4084 (N_4084,N_1971,N_2037);
or U4085 (N_4085,N_2411,N_1519);
nand U4086 (N_4086,N_998,N_909);
or U4087 (N_4087,N_136,N_891);
nand U4088 (N_4088,N_1352,N_1021);
and U4089 (N_4089,N_1449,N_710);
nor U4090 (N_4090,N_1962,N_1373);
nand U4091 (N_4091,N_1015,N_108);
or U4092 (N_4092,N_711,N_1656);
and U4093 (N_4093,N_734,N_2142);
nor U4094 (N_4094,N_1982,N_2404);
and U4095 (N_4095,N_350,N_2410);
nor U4096 (N_4096,N_1528,N_1384);
and U4097 (N_4097,N_1509,N_1398);
nand U4098 (N_4098,N_321,N_2352);
nor U4099 (N_4099,N_927,N_1011);
nand U4100 (N_4100,N_2193,N_1029);
nand U4101 (N_4101,N_2105,N_1989);
nand U4102 (N_4102,N_2349,N_1860);
or U4103 (N_4103,N_1425,N_974);
nor U4104 (N_4104,N_1616,N_351);
and U4105 (N_4105,N_432,N_658);
and U4106 (N_4106,N_2462,N_1905);
and U4107 (N_4107,N_1185,N_981);
or U4108 (N_4108,N_2207,N_792);
and U4109 (N_4109,N_2165,N_1403);
or U4110 (N_4110,N_109,N_2111);
and U4111 (N_4111,N_739,N_1281);
nand U4112 (N_4112,N_2430,N_701);
or U4113 (N_4113,N_751,N_2282);
or U4114 (N_4114,N_1894,N_1163);
nand U4115 (N_4115,N_2205,N_1330);
or U4116 (N_4116,N_1102,N_687);
nor U4117 (N_4117,N_1633,N_1257);
and U4118 (N_4118,N_1228,N_612);
nor U4119 (N_4119,N_2154,N_161);
or U4120 (N_4120,N_1212,N_433);
or U4121 (N_4121,N_1552,N_1183);
nor U4122 (N_4122,N_355,N_105);
and U4123 (N_4123,N_699,N_2285);
nand U4124 (N_4124,N_1245,N_114);
nand U4125 (N_4125,N_163,N_2365);
nand U4126 (N_4126,N_1643,N_856);
nand U4127 (N_4127,N_268,N_2223);
nor U4128 (N_4128,N_1623,N_1844);
nor U4129 (N_4129,N_684,N_1758);
or U4130 (N_4130,N_955,N_884);
and U4131 (N_4131,N_247,N_793);
nand U4132 (N_4132,N_2196,N_2374);
or U4133 (N_4133,N_1444,N_2253);
nor U4134 (N_4134,N_1620,N_1943);
or U4135 (N_4135,N_533,N_1575);
nand U4136 (N_4136,N_2227,N_296);
nor U4137 (N_4137,N_2100,N_2259);
or U4138 (N_4138,N_1140,N_1489);
nand U4139 (N_4139,N_1125,N_2174);
nand U4140 (N_4140,N_1568,N_65);
and U4141 (N_4141,N_2272,N_2294);
or U4142 (N_4142,N_512,N_2105);
nand U4143 (N_4143,N_753,N_932);
or U4144 (N_4144,N_1007,N_829);
and U4145 (N_4145,N_1234,N_1241);
or U4146 (N_4146,N_2407,N_399);
nor U4147 (N_4147,N_51,N_2128);
nor U4148 (N_4148,N_2102,N_2260);
nand U4149 (N_4149,N_874,N_2209);
and U4150 (N_4150,N_1198,N_855);
or U4151 (N_4151,N_2237,N_286);
and U4152 (N_4152,N_315,N_2270);
nand U4153 (N_4153,N_137,N_2101);
or U4154 (N_4154,N_380,N_1670);
or U4155 (N_4155,N_878,N_818);
and U4156 (N_4156,N_1816,N_1089);
nor U4157 (N_4157,N_956,N_2270);
and U4158 (N_4158,N_594,N_1199);
nor U4159 (N_4159,N_876,N_946);
and U4160 (N_4160,N_1009,N_1951);
nand U4161 (N_4161,N_986,N_1096);
and U4162 (N_4162,N_2165,N_228);
or U4163 (N_4163,N_2062,N_1962);
or U4164 (N_4164,N_392,N_1385);
or U4165 (N_4165,N_1537,N_248);
nor U4166 (N_4166,N_1788,N_684);
or U4167 (N_4167,N_274,N_579);
and U4168 (N_4168,N_1665,N_340);
and U4169 (N_4169,N_1851,N_2142);
nand U4170 (N_4170,N_2060,N_111);
nor U4171 (N_4171,N_13,N_2074);
and U4172 (N_4172,N_1412,N_521);
and U4173 (N_4173,N_1676,N_1144);
nand U4174 (N_4174,N_414,N_935);
nor U4175 (N_4175,N_1812,N_115);
nor U4176 (N_4176,N_319,N_315);
nand U4177 (N_4177,N_2289,N_132);
and U4178 (N_4178,N_147,N_522);
xor U4179 (N_4179,N_572,N_2346);
or U4180 (N_4180,N_259,N_1621);
nor U4181 (N_4181,N_1979,N_1902);
and U4182 (N_4182,N_1465,N_1602);
and U4183 (N_4183,N_857,N_918);
nor U4184 (N_4184,N_2210,N_1952);
xnor U4185 (N_4185,N_1285,N_1654);
nand U4186 (N_4186,N_2340,N_2135);
nand U4187 (N_4187,N_1395,N_2396);
nor U4188 (N_4188,N_950,N_55);
or U4189 (N_4189,N_0,N_1308);
and U4190 (N_4190,N_2198,N_1096);
or U4191 (N_4191,N_351,N_2393);
nand U4192 (N_4192,N_914,N_2249);
or U4193 (N_4193,N_473,N_1374);
nand U4194 (N_4194,N_1649,N_1381);
nand U4195 (N_4195,N_143,N_1110);
or U4196 (N_4196,N_245,N_684);
or U4197 (N_4197,N_2187,N_1316);
nand U4198 (N_4198,N_2490,N_1995);
and U4199 (N_4199,N_76,N_1748);
or U4200 (N_4200,N_242,N_1436);
nor U4201 (N_4201,N_373,N_674);
and U4202 (N_4202,N_1513,N_211);
and U4203 (N_4203,N_212,N_1182);
nor U4204 (N_4204,N_2223,N_2307);
nand U4205 (N_4205,N_779,N_1969);
and U4206 (N_4206,N_1711,N_2497);
nor U4207 (N_4207,N_1613,N_96);
and U4208 (N_4208,N_108,N_1556);
nor U4209 (N_4209,N_115,N_217);
nor U4210 (N_4210,N_367,N_1036);
nor U4211 (N_4211,N_1242,N_2326);
or U4212 (N_4212,N_791,N_582);
or U4213 (N_4213,N_877,N_1919);
nand U4214 (N_4214,N_1005,N_743);
or U4215 (N_4215,N_889,N_2275);
and U4216 (N_4216,N_855,N_1155);
nor U4217 (N_4217,N_2346,N_698);
or U4218 (N_4218,N_978,N_800);
and U4219 (N_4219,N_756,N_868);
nand U4220 (N_4220,N_1006,N_1121);
xnor U4221 (N_4221,N_1981,N_1473);
or U4222 (N_4222,N_275,N_1407);
and U4223 (N_4223,N_2160,N_299);
and U4224 (N_4224,N_541,N_2352);
and U4225 (N_4225,N_1276,N_101);
and U4226 (N_4226,N_368,N_1096);
and U4227 (N_4227,N_2465,N_206);
nand U4228 (N_4228,N_1542,N_1810);
and U4229 (N_4229,N_1929,N_92);
nor U4230 (N_4230,N_145,N_2317);
nand U4231 (N_4231,N_1212,N_289);
nand U4232 (N_4232,N_454,N_2278);
or U4233 (N_4233,N_802,N_2017);
and U4234 (N_4234,N_1472,N_2095);
and U4235 (N_4235,N_1824,N_1074);
xnor U4236 (N_4236,N_2056,N_650);
nor U4237 (N_4237,N_1624,N_1143);
nor U4238 (N_4238,N_1017,N_2135);
nand U4239 (N_4239,N_2299,N_2261);
and U4240 (N_4240,N_1725,N_1279);
nor U4241 (N_4241,N_1774,N_989);
and U4242 (N_4242,N_1633,N_1203);
and U4243 (N_4243,N_2196,N_8);
and U4244 (N_4244,N_31,N_85);
nand U4245 (N_4245,N_907,N_2422);
xnor U4246 (N_4246,N_1142,N_2011);
or U4247 (N_4247,N_1598,N_2327);
nor U4248 (N_4248,N_389,N_67);
and U4249 (N_4249,N_407,N_836);
and U4250 (N_4250,N_2140,N_84);
nor U4251 (N_4251,N_1894,N_1062);
or U4252 (N_4252,N_2232,N_952);
and U4253 (N_4253,N_2113,N_2401);
nand U4254 (N_4254,N_2032,N_833);
or U4255 (N_4255,N_2107,N_1174);
nand U4256 (N_4256,N_2486,N_2461);
or U4257 (N_4257,N_2048,N_2103);
and U4258 (N_4258,N_752,N_2405);
or U4259 (N_4259,N_2175,N_2367);
and U4260 (N_4260,N_224,N_168);
or U4261 (N_4261,N_1171,N_2137);
nor U4262 (N_4262,N_1099,N_2107);
nand U4263 (N_4263,N_327,N_1072);
and U4264 (N_4264,N_1755,N_103);
nor U4265 (N_4265,N_1285,N_584);
nor U4266 (N_4266,N_2061,N_1580);
nand U4267 (N_4267,N_1692,N_2234);
and U4268 (N_4268,N_1330,N_903);
or U4269 (N_4269,N_265,N_591);
or U4270 (N_4270,N_748,N_2227);
or U4271 (N_4271,N_1985,N_1493);
nor U4272 (N_4272,N_1446,N_1568);
nor U4273 (N_4273,N_1740,N_2164);
and U4274 (N_4274,N_723,N_436);
nor U4275 (N_4275,N_1164,N_1041);
nor U4276 (N_4276,N_1501,N_1552);
or U4277 (N_4277,N_1250,N_652);
and U4278 (N_4278,N_642,N_215);
nand U4279 (N_4279,N_2057,N_2071);
or U4280 (N_4280,N_1461,N_2213);
nand U4281 (N_4281,N_529,N_2265);
and U4282 (N_4282,N_1879,N_418);
nand U4283 (N_4283,N_632,N_1597);
nor U4284 (N_4284,N_1817,N_1547);
nand U4285 (N_4285,N_279,N_166);
and U4286 (N_4286,N_1739,N_1579);
xnor U4287 (N_4287,N_93,N_594);
or U4288 (N_4288,N_291,N_977);
nor U4289 (N_4289,N_510,N_801);
or U4290 (N_4290,N_21,N_1607);
nor U4291 (N_4291,N_111,N_636);
or U4292 (N_4292,N_2066,N_1121);
nand U4293 (N_4293,N_563,N_466);
and U4294 (N_4294,N_2269,N_2388);
nand U4295 (N_4295,N_2348,N_1614);
nor U4296 (N_4296,N_974,N_959);
and U4297 (N_4297,N_1034,N_565);
nand U4298 (N_4298,N_44,N_1943);
and U4299 (N_4299,N_1903,N_1223);
nor U4300 (N_4300,N_1724,N_1903);
or U4301 (N_4301,N_885,N_844);
nor U4302 (N_4302,N_1793,N_812);
nand U4303 (N_4303,N_20,N_2401);
nor U4304 (N_4304,N_452,N_635);
and U4305 (N_4305,N_2328,N_621);
nor U4306 (N_4306,N_2389,N_473);
and U4307 (N_4307,N_2330,N_87);
nand U4308 (N_4308,N_2154,N_745);
or U4309 (N_4309,N_395,N_1586);
xor U4310 (N_4310,N_1621,N_1644);
and U4311 (N_4311,N_1815,N_1589);
or U4312 (N_4312,N_517,N_1819);
or U4313 (N_4313,N_1763,N_2046);
nor U4314 (N_4314,N_1676,N_594);
or U4315 (N_4315,N_175,N_1072);
nor U4316 (N_4316,N_699,N_1871);
or U4317 (N_4317,N_1135,N_1677);
or U4318 (N_4318,N_289,N_1747);
nand U4319 (N_4319,N_605,N_2328);
nor U4320 (N_4320,N_2125,N_2286);
or U4321 (N_4321,N_1753,N_1023);
nand U4322 (N_4322,N_2253,N_2470);
nand U4323 (N_4323,N_2238,N_862);
or U4324 (N_4324,N_214,N_2403);
or U4325 (N_4325,N_69,N_1650);
or U4326 (N_4326,N_1561,N_1810);
nand U4327 (N_4327,N_418,N_1405);
and U4328 (N_4328,N_1330,N_1070);
or U4329 (N_4329,N_580,N_220);
and U4330 (N_4330,N_649,N_1934);
and U4331 (N_4331,N_1754,N_87);
nor U4332 (N_4332,N_1848,N_605);
or U4333 (N_4333,N_2157,N_825);
or U4334 (N_4334,N_2033,N_1561);
nor U4335 (N_4335,N_738,N_1701);
nand U4336 (N_4336,N_694,N_987);
nor U4337 (N_4337,N_1079,N_2333);
nand U4338 (N_4338,N_122,N_1307);
or U4339 (N_4339,N_132,N_35);
nand U4340 (N_4340,N_1158,N_291);
nor U4341 (N_4341,N_2119,N_2495);
nand U4342 (N_4342,N_13,N_1633);
or U4343 (N_4343,N_663,N_1473);
nor U4344 (N_4344,N_1673,N_2492);
nand U4345 (N_4345,N_1857,N_812);
nor U4346 (N_4346,N_282,N_1116);
nand U4347 (N_4347,N_2258,N_634);
nor U4348 (N_4348,N_705,N_123);
or U4349 (N_4349,N_47,N_629);
or U4350 (N_4350,N_587,N_799);
nand U4351 (N_4351,N_855,N_195);
nand U4352 (N_4352,N_756,N_1649);
or U4353 (N_4353,N_861,N_1592);
or U4354 (N_4354,N_2358,N_1953);
nand U4355 (N_4355,N_176,N_1788);
or U4356 (N_4356,N_23,N_56);
nor U4357 (N_4357,N_1907,N_1309);
or U4358 (N_4358,N_498,N_2351);
nand U4359 (N_4359,N_1685,N_552);
or U4360 (N_4360,N_1886,N_1842);
or U4361 (N_4361,N_902,N_1462);
nor U4362 (N_4362,N_615,N_805);
or U4363 (N_4363,N_1784,N_2121);
nand U4364 (N_4364,N_1626,N_1480);
nor U4365 (N_4365,N_741,N_217);
or U4366 (N_4366,N_2216,N_622);
nand U4367 (N_4367,N_1400,N_1443);
and U4368 (N_4368,N_1609,N_1382);
nand U4369 (N_4369,N_1334,N_457);
and U4370 (N_4370,N_1605,N_2472);
or U4371 (N_4371,N_139,N_1634);
or U4372 (N_4372,N_1974,N_1096);
or U4373 (N_4373,N_968,N_1582);
nor U4374 (N_4374,N_2476,N_2344);
and U4375 (N_4375,N_196,N_978);
nor U4376 (N_4376,N_952,N_709);
nor U4377 (N_4377,N_820,N_1251);
nand U4378 (N_4378,N_2493,N_1928);
nand U4379 (N_4379,N_491,N_1451);
nand U4380 (N_4380,N_1615,N_656);
nor U4381 (N_4381,N_859,N_621);
and U4382 (N_4382,N_1172,N_2110);
nor U4383 (N_4383,N_726,N_2446);
or U4384 (N_4384,N_551,N_703);
and U4385 (N_4385,N_1828,N_851);
or U4386 (N_4386,N_923,N_1220);
and U4387 (N_4387,N_260,N_1914);
nor U4388 (N_4388,N_2197,N_1254);
or U4389 (N_4389,N_113,N_701);
or U4390 (N_4390,N_730,N_386);
nand U4391 (N_4391,N_1948,N_919);
and U4392 (N_4392,N_858,N_2242);
nor U4393 (N_4393,N_177,N_1374);
nor U4394 (N_4394,N_1033,N_666);
nor U4395 (N_4395,N_1508,N_2180);
or U4396 (N_4396,N_1665,N_1277);
or U4397 (N_4397,N_1799,N_2464);
or U4398 (N_4398,N_358,N_181);
nor U4399 (N_4399,N_837,N_1736);
nand U4400 (N_4400,N_1734,N_1276);
and U4401 (N_4401,N_397,N_704);
or U4402 (N_4402,N_134,N_766);
nor U4403 (N_4403,N_1108,N_1784);
nand U4404 (N_4404,N_441,N_1733);
nor U4405 (N_4405,N_470,N_318);
nand U4406 (N_4406,N_1915,N_1301);
or U4407 (N_4407,N_1301,N_1888);
nand U4408 (N_4408,N_1895,N_996);
or U4409 (N_4409,N_3,N_178);
nand U4410 (N_4410,N_890,N_2202);
or U4411 (N_4411,N_1712,N_1943);
and U4412 (N_4412,N_2262,N_682);
and U4413 (N_4413,N_1964,N_1024);
nand U4414 (N_4414,N_1013,N_2111);
and U4415 (N_4415,N_2107,N_460);
nand U4416 (N_4416,N_1685,N_542);
nor U4417 (N_4417,N_1509,N_104);
nand U4418 (N_4418,N_476,N_2187);
or U4419 (N_4419,N_2382,N_2087);
and U4420 (N_4420,N_385,N_2313);
and U4421 (N_4421,N_2263,N_1113);
or U4422 (N_4422,N_1669,N_1886);
nand U4423 (N_4423,N_584,N_111);
or U4424 (N_4424,N_806,N_1612);
nor U4425 (N_4425,N_1569,N_2458);
nand U4426 (N_4426,N_286,N_876);
nor U4427 (N_4427,N_195,N_2128);
or U4428 (N_4428,N_1697,N_2057);
or U4429 (N_4429,N_1970,N_1139);
nor U4430 (N_4430,N_908,N_509);
and U4431 (N_4431,N_648,N_414);
or U4432 (N_4432,N_844,N_2445);
nand U4433 (N_4433,N_1324,N_1430);
and U4434 (N_4434,N_129,N_2448);
or U4435 (N_4435,N_1985,N_2465);
nand U4436 (N_4436,N_863,N_437);
or U4437 (N_4437,N_2090,N_224);
and U4438 (N_4438,N_937,N_2239);
nor U4439 (N_4439,N_1227,N_201);
or U4440 (N_4440,N_1477,N_1693);
and U4441 (N_4441,N_1963,N_2074);
or U4442 (N_4442,N_1009,N_2113);
and U4443 (N_4443,N_791,N_2096);
nor U4444 (N_4444,N_1764,N_234);
nor U4445 (N_4445,N_10,N_908);
and U4446 (N_4446,N_2125,N_379);
nor U4447 (N_4447,N_2461,N_935);
nor U4448 (N_4448,N_2029,N_605);
nand U4449 (N_4449,N_2027,N_1812);
or U4450 (N_4450,N_63,N_736);
and U4451 (N_4451,N_2201,N_818);
nand U4452 (N_4452,N_2399,N_931);
nor U4453 (N_4453,N_2230,N_2232);
nand U4454 (N_4454,N_1234,N_1578);
and U4455 (N_4455,N_40,N_709);
or U4456 (N_4456,N_313,N_862);
and U4457 (N_4457,N_855,N_1738);
nor U4458 (N_4458,N_1201,N_1028);
or U4459 (N_4459,N_1309,N_2325);
nand U4460 (N_4460,N_2178,N_1072);
or U4461 (N_4461,N_1315,N_1783);
or U4462 (N_4462,N_932,N_2359);
and U4463 (N_4463,N_139,N_370);
xor U4464 (N_4464,N_292,N_1993);
or U4465 (N_4465,N_635,N_200);
and U4466 (N_4466,N_1947,N_149);
or U4467 (N_4467,N_2324,N_1660);
nand U4468 (N_4468,N_1696,N_1990);
nand U4469 (N_4469,N_2081,N_333);
and U4470 (N_4470,N_734,N_2097);
or U4471 (N_4471,N_413,N_1144);
and U4472 (N_4472,N_2332,N_2329);
or U4473 (N_4473,N_1045,N_93);
nor U4474 (N_4474,N_1071,N_1961);
and U4475 (N_4475,N_1041,N_1792);
and U4476 (N_4476,N_673,N_2456);
nor U4477 (N_4477,N_393,N_1759);
nand U4478 (N_4478,N_1073,N_785);
and U4479 (N_4479,N_317,N_1145);
nand U4480 (N_4480,N_2419,N_1595);
or U4481 (N_4481,N_2214,N_736);
or U4482 (N_4482,N_173,N_2197);
and U4483 (N_4483,N_959,N_570);
or U4484 (N_4484,N_1426,N_1984);
and U4485 (N_4485,N_381,N_700);
nand U4486 (N_4486,N_2420,N_2364);
or U4487 (N_4487,N_386,N_511);
or U4488 (N_4488,N_521,N_2436);
nor U4489 (N_4489,N_1134,N_66);
nand U4490 (N_4490,N_2360,N_2132);
nor U4491 (N_4491,N_1689,N_791);
nand U4492 (N_4492,N_433,N_2164);
and U4493 (N_4493,N_951,N_536);
or U4494 (N_4494,N_809,N_1495);
nand U4495 (N_4495,N_1434,N_725);
nand U4496 (N_4496,N_1211,N_2221);
or U4497 (N_4497,N_584,N_466);
or U4498 (N_4498,N_1882,N_404);
nand U4499 (N_4499,N_1424,N_1769);
and U4500 (N_4500,N_237,N_1639);
or U4501 (N_4501,N_1731,N_2049);
nand U4502 (N_4502,N_1659,N_53);
or U4503 (N_4503,N_1742,N_974);
nor U4504 (N_4504,N_1041,N_50);
and U4505 (N_4505,N_2470,N_55);
or U4506 (N_4506,N_963,N_1933);
and U4507 (N_4507,N_1423,N_961);
or U4508 (N_4508,N_1936,N_1373);
nand U4509 (N_4509,N_1273,N_501);
or U4510 (N_4510,N_799,N_2376);
and U4511 (N_4511,N_512,N_1412);
nand U4512 (N_4512,N_10,N_502);
and U4513 (N_4513,N_98,N_2241);
or U4514 (N_4514,N_1356,N_2035);
nand U4515 (N_4515,N_985,N_582);
or U4516 (N_4516,N_2062,N_1796);
nor U4517 (N_4517,N_719,N_649);
or U4518 (N_4518,N_1684,N_2440);
and U4519 (N_4519,N_529,N_2007);
or U4520 (N_4520,N_2266,N_658);
nand U4521 (N_4521,N_1264,N_1451);
or U4522 (N_4522,N_1639,N_1038);
or U4523 (N_4523,N_475,N_266);
nor U4524 (N_4524,N_1620,N_1331);
or U4525 (N_4525,N_1771,N_33);
or U4526 (N_4526,N_2281,N_2459);
nor U4527 (N_4527,N_1430,N_1678);
nor U4528 (N_4528,N_2236,N_1723);
nand U4529 (N_4529,N_1620,N_1994);
or U4530 (N_4530,N_1025,N_1340);
or U4531 (N_4531,N_150,N_1063);
or U4532 (N_4532,N_1786,N_2256);
or U4533 (N_4533,N_2167,N_1072);
nor U4534 (N_4534,N_2222,N_2009);
and U4535 (N_4535,N_1658,N_1141);
and U4536 (N_4536,N_1316,N_921);
nor U4537 (N_4537,N_512,N_858);
nand U4538 (N_4538,N_17,N_1220);
nand U4539 (N_4539,N_831,N_1612);
and U4540 (N_4540,N_294,N_1596);
nor U4541 (N_4541,N_2059,N_603);
or U4542 (N_4542,N_325,N_533);
and U4543 (N_4543,N_1247,N_1490);
nand U4544 (N_4544,N_1981,N_665);
or U4545 (N_4545,N_1211,N_2280);
or U4546 (N_4546,N_2277,N_1371);
nand U4547 (N_4547,N_1409,N_298);
nand U4548 (N_4548,N_334,N_689);
and U4549 (N_4549,N_845,N_233);
nor U4550 (N_4550,N_191,N_829);
or U4551 (N_4551,N_1642,N_2314);
nor U4552 (N_4552,N_881,N_2029);
or U4553 (N_4553,N_2325,N_1645);
and U4554 (N_4554,N_824,N_1589);
nand U4555 (N_4555,N_1373,N_766);
nor U4556 (N_4556,N_703,N_589);
and U4557 (N_4557,N_1582,N_2365);
nor U4558 (N_4558,N_13,N_502);
or U4559 (N_4559,N_592,N_74);
nand U4560 (N_4560,N_1159,N_2100);
and U4561 (N_4561,N_2392,N_1798);
and U4562 (N_4562,N_1108,N_1478);
xnor U4563 (N_4563,N_405,N_349);
nand U4564 (N_4564,N_134,N_773);
nand U4565 (N_4565,N_1154,N_798);
or U4566 (N_4566,N_223,N_1048);
nand U4567 (N_4567,N_1053,N_1246);
or U4568 (N_4568,N_1029,N_83);
nor U4569 (N_4569,N_2479,N_901);
nor U4570 (N_4570,N_231,N_1515);
or U4571 (N_4571,N_1929,N_2389);
nor U4572 (N_4572,N_988,N_339);
nor U4573 (N_4573,N_1089,N_11);
or U4574 (N_4574,N_1905,N_1241);
and U4575 (N_4575,N_559,N_1987);
and U4576 (N_4576,N_2133,N_2047);
nor U4577 (N_4577,N_1481,N_2166);
xor U4578 (N_4578,N_671,N_791);
or U4579 (N_4579,N_97,N_2290);
or U4580 (N_4580,N_2014,N_531);
nand U4581 (N_4581,N_1242,N_2142);
nor U4582 (N_4582,N_1199,N_188);
nand U4583 (N_4583,N_2164,N_2439);
or U4584 (N_4584,N_1471,N_1103);
nor U4585 (N_4585,N_1204,N_186);
and U4586 (N_4586,N_659,N_261);
or U4587 (N_4587,N_1357,N_1467);
and U4588 (N_4588,N_1915,N_2005);
xnor U4589 (N_4589,N_1192,N_833);
or U4590 (N_4590,N_2354,N_873);
nor U4591 (N_4591,N_134,N_263);
or U4592 (N_4592,N_833,N_1901);
nor U4593 (N_4593,N_236,N_1503);
or U4594 (N_4594,N_1552,N_301);
or U4595 (N_4595,N_573,N_129);
nand U4596 (N_4596,N_1202,N_2271);
and U4597 (N_4597,N_1655,N_103);
nand U4598 (N_4598,N_908,N_1409);
nor U4599 (N_4599,N_130,N_74);
nor U4600 (N_4600,N_1373,N_2189);
or U4601 (N_4601,N_1127,N_173);
nand U4602 (N_4602,N_985,N_505);
and U4603 (N_4603,N_1052,N_2418);
nor U4604 (N_4604,N_1670,N_1623);
nand U4605 (N_4605,N_190,N_1641);
xor U4606 (N_4606,N_85,N_1704);
and U4607 (N_4607,N_1996,N_1311);
nand U4608 (N_4608,N_1879,N_2409);
and U4609 (N_4609,N_196,N_1079);
or U4610 (N_4610,N_388,N_1173);
nor U4611 (N_4611,N_1937,N_2305);
and U4612 (N_4612,N_2147,N_2429);
and U4613 (N_4613,N_2027,N_1386);
or U4614 (N_4614,N_795,N_353);
or U4615 (N_4615,N_62,N_861);
or U4616 (N_4616,N_688,N_528);
or U4617 (N_4617,N_1255,N_2281);
nor U4618 (N_4618,N_1515,N_461);
or U4619 (N_4619,N_131,N_88);
or U4620 (N_4620,N_1924,N_1537);
nor U4621 (N_4621,N_1355,N_1804);
or U4622 (N_4622,N_1096,N_2367);
xor U4623 (N_4623,N_2370,N_1630);
nand U4624 (N_4624,N_1924,N_1428);
and U4625 (N_4625,N_1167,N_1940);
or U4626 (N_4626,N_1571,N_1090);
or U4627 (N_4627,N_778,N_263);
or U4628 (N_4628,N_454,N_1147);
or U4629 (N_4629,N_884,N_343);
and U4630 (N_4630,N_2453,N_1624);
and U4631 (N_4631,N_156,N_1384);
and U4632 (N_4632,N_646,N_1041);
and U4633 (N_4633,N_1795,N_2093);
xnor U4634 (N_4634,N_441,N_660);
nand U4635 (N_4635,N_1020,N_465);
nand U4636 (N_4636,N_618,N_127);
and U4637 (N_4637,N_1282,N_637);
and U4638 (N_4638,N_1267,N_567);
or U4639 (N_4639,N_1673,N_610);
nor U4640 (N_4640,N_615,N_2267);
or U4641 (N_4641,N_50,N_2204);
or U4642 (N_4642,N_1602,N_1281);
or U4643 (N_4643,N_1736,N_930);
nand U4644 (N_4644,N_1899,N_867);
nand U4645 (N_4645,N_1729,N_381);
or U4646 (N_4646,N_1112,N_825);
or U4647 (N_4647,N_1664,N_1062);
nor U4648 (N_4648,N_1432,N_985);
and U4649 (N_4649,N_2165,N_1215);
and U4650 (N_4650,N_2383,N_1430);
nand U4651 (N_4651,N_73,N_643);
xnor U4652 (N_4652,N_450,N_902);
or U4653 (N_4653,N_350,N_2203);
or U4654 (N_4654,N_273,N_551);
xor U4655 (N_4655,N_2383,N_1354);
nand U4656 (N_4656,N_884,N_626);
nor U4657 (N_4657,N_80,N_2210);
and U4658 (N_4658,N_903,N_84);
or U4659 (N_4659,N_535,N_1814);
nor U4660 (N_4660,N_461,N_330);
nor U4661 (N_4661,N_252,N_1630);
and U4662 (N_4662,N_2280,N_536);
nand U4663 (N_4663,N_2347,N_1694);
and U4664 (N_4664,N_1486,N_1406);
and U4665 (N_4665,N_1204,N_117);
or U4666 (N_4666,N_339,N_207);
nor U4667 (N_4667,N_1675,N_2082);
nand U4668 (N_4668,N_1880,N_2243);
nor U4669 (N_4669,N_1439,N_1634);
and U4670 (N_4670,N_1892,N_693);
or U4671 (N_4671,N_691,N_924);
nand U4672 (N_4672,N_1176,N_467);
and U4673 (N_4673,N_2089,N_324);
nor U4674 (N_4674,N_1274,N_1320);
or U4675 (N_4675,N_106,N_381);
nand U4676 (N_4676,N_483,N_2003);
nand U4677 (N_4677,N_24,N_2331);
and U4678 (N_4678,N_1942,N_1296);
nand U4679 (N_4679,N_838,N_2467);
and U4680 (N_4680,N_1433,N_13);
and U4681 (N_4681,N_2176,N_2396);
nand U4682 (N_4682,N_1645,N_1019);
and U4683 (N_4683,N_773,N_839);
nor U4684 (N_4684,N_2014,N_1561);
or U4685 (N_4685,N_1154,N_1484);
or U4686 (N_4686,N_1513,N_1753);
nand U4687 (N_4687,N_1881,N_2035);
or U4688 (N_4688,N_2139,N_643);
and U4689 (N_4689,N_885,N_1626);
nand U4690 (N_4690,N_2250,N_492);
nor U4691 (N_4691,N_569,N_1826);
or U4692 (N_4692,N_1321,N_2118);
xnor U4693 (N_4693,N_352,N_1124);
or U4694 (N_4694,N_2032,N_718);
or U4695 (N_4695,N_385,N_362);
xnor U4696 (N_4696,N_2396,N_1936);
nor U4697 (N_4697,N_652,N_2297);
nand U4698 (N_4698,N_853,N_1533);
nand U4699 (N_4699,N_2443,N_1911);
nand U4700 (N_4700,N_374,N_1143);
or U4701 (N_4701,N_795,N_2288);
or U4702 (N_4702,N_119,N_1542);
or U4703 (N_4703,N_237,N_881);
and U4704 (N_4704,N_1016,N_1546);
nor U4705 (N_4705,N_185,N_1596);
nor U4706 (N_4706,N_1361,N_2318);
and U4707 (N_4707,N_1578,N_1696);
nor U4708 (N_4708,N_2144,N_2105);
and U4709 (N_4709,N_217,N_714);
and U4710 (N_4710,N_2475,N_1135);
nor U4711 (N_4711,N_570,N_2101);
and U4712 (N_4712,N_1307,N_534);
nand U4713 (N_4713,N_2347,N_728);
nor U4714 (N_4714,N_843,N_672);
and U4715 (N_4715,N_1966,N_2074);
xnor U4716 (N_4716,N_1668,N_389);
nand U4717 (N_4717,N_2361,N_1267);
and U4718 (N_4718,N_1501,N_125);
or U4719 (N_4719,N_1320,N_605);
nor U4720 (N_4720,N_54,N_1296);
and U4721 (N_4721,N_159,N_610);
xnor U4722 (N_4722,N_2333,N_1870);
nor U4723 (N_4723,N_970,N_1869);
nor U4724 (N_4724,N_1574,N_1888);
and U4725 (N_4725,N_684,N_584);
or U4726 (N_4726,N_1922,N_2103);
and U4727 (N_4727,N_1309,N_2106);
nand U4728 (N_4728,N_739,N_1638);
nor U4729 (N_4729,N_20,N_1202);
nand U4730 (N_4730,N_991,N_1836);
or U4731 (N_4731,N_271,N_587);
nor U4732 (N_4732,N_1071,N_1032);
or U4733 (N_4733,N_1095,N_1012);
or U4734 (N_4734,N_77,N_2174);
and U4735 (N_4735,N_1729,N_2281);
nor U4736 (N_4736,N_172,N_1852);
or U4737 (N_4737,N_1912,N_2330);
and U4738 (N_4738,N_574,N_738);
nor U4739 (N_4739,N_262,N_21);
nor U4740 (N_4740,N_986,N_564);
nand U4741 (N_4741,N_1523,N_1112);
nor U4742 (N_4742,N_1251,N_691);
nand U4743 (N_4743,N_597,N_556);
nand U4744 (N_4744,N_1884,N_1371);
and U4745 (N_4745,N_449,N_2226);
or U4746 (N_4746,N_983,N_2115);
and U4747 (N_4747,N_1691,N_12);
or U4748 (N_4748,N_2124,N_367);
nand U4749 (N_4749,N_2459,N_1017);
and U4750 (N_4750,N_1022,N_2138);
and U4751 (N_4751,N_2441,N_1796);
nor U4752 (N_4752,N_2160,N_1086);
and U4753 (N_4753,N_2376,N_2107);
and U4754 (N_4754,N_1340,N_2174);
or U4755 (N_4755,N_332,N_944);
nor U4756 (N_4756,N_327,N_1939);
nand U4757 (N_4757,N_1779,N_1982);
and U4758 (N_4758,N_324,N_1614);
nor U4759 (N_4759,N_2010,N_620);
nor U4760 (N_4760,N_2136,N_615);
and U4761 (N_4761,N_1163,N_363);
and U4762 (N_4762,N_604,N_1919);
nor U4763 (N_4763,N_761,N_1279);
nand U4764 (N_4764,N_390,N_1026);
nor U4765 (N_4765,N_129,N_44);
and U4766 (N_4766,N_776,N_64);
nor U4767 (N_4767,N_1621,N_1216);
and U4768 (N_4768,N_989,N_273);
or U4769 (N_4769,N_2389,N_1935);
nor U4770 (N_4770,N_1567,N_2193);
or U4771 (N_4771,N_1719,N_2189);
nor U4772 (N_4772,N_2128,N_1566);
xnor U4773 (N_4773,N_466,N_712);
nand U4774 (N_4774,N_2315,N_134);
nand U4775 (N_4775,N_911,N_970);
or U4776 (N_4776,N_1088,N_886);
and U4777 (N_4777,N_1300,N_1290);
and U4778 (N_4778,N_609,N_1474);
nor U4779 (N_4779,N_677,N_1838);
and U4780 (N_4780,N_2359,N_1357);
xor U4781 (N_4781,N_2108,N_122);
nor U4782 (N_4782,N_1240,N_795);
or U4783 (N_4783,N_607,N_1664);
nor U4784 (N_4784,N_2481,N_609);
xor U4785 (N_4785,N_2380,N_1166);
or U4786 (N_4786,N_349,N_1759);
or U4787 (N_4787,N_1790,N_1698);
nor U4788 (N_4788,N_1937,N_787);
xor U4789 (N_4789,N_2136,N_913);
nand U4790 (N_4790,N_1860,N_1357);
nand U4791 (N_4791,N_344,N_291);
and U4792 (N_4792,N_1424,N_2066);
nor U4793 (N_4793,N_2028,N_363);
and U4794 (N_4794,N_2289,N_600);
or U4795 (N_4795,N_1807,N_2298);
and U4796 (N_4796,N_2435,N_6);
nor U4797 (N_4797,N_1270,N_474);
xnor U4798 (N_4798,N_1229,N_708);
nor U4799 (N_4799,N_2221,N_879);
nor U4800 (N_4800,N_292,N_1238);
xnor U4801 (N_4801,N_920,N_1784);
nand U4802 (N_4802,N_869,N_479);
and U4803 (N_4803,N_57,N_1912);
nor U4804 (N_4804,N_1461,N_2469);
nor U4805 (N_4805,N_1361,N_2185);
nand U4806 (N_4806,N_1609,N_61);
nand U4807 (N_4807,N_966,N_2035);
and U4808 (N_4808,N_2109,N_2204);
and U4809 (N_4809,N_300,N_1411);
nand U4810 (N_4810,N_2073,N_2178);
nand U4811 (N_4811,N_1243,N_1927);
or U4812 (N_4812,N_676,N_2412);
nor U4813 (N_4813,N_2126,N_131);
nand U4814 (N_4814,N_947,N_716);
or U4815 (N_4815,N_1230,N_1899);
or U4816 (N_4816,N_666,N_1603);
nor U4817 (N_4817,N_1,N_1145);
and U4818 (N_4818,N_2068,N_461);
and U4819 (N_4819,N_1171,N_1123);
or U4820 (N_4820,N_2308,N_884);
and U4821 (N_4821,N_1735,N_1102);
nand U4822 (N_4822,N_2466,N_2446);
or U4823 (N_4823,N_1217,N_680);
and U4824 (N_4824,N_1473,N_2268);
nor U4825 (N_4825,N_261,N_1183);
nand U4826 (N_4826,N_99,N_1740);
and U4827 (N_4827,N_667,N_2351);
nand U4828 (N_4828,N_899,N_1675);
and U4829 (N_4829,N_1484,N_357);
nor U4830 (N_4830,N_1956,N_1372);
and U4831 (N_4831,N_2403,N_2351);
nor U4832 (N_4832,N_2085,N_2263);
nand U4833 (N_4833,N_1454,N_126);
or U4834 (N_4834,N_1264,N_551);
nand U4835 (N_4835,N_523,N_2078);
nand U4836 (N_4836,N_1706,N_2139);
or U4837 (N_4837,N_488,N_1087);
nand U4838 (N_4838,N_141,N_1018);
xor U4839 (N_4839,N_2140,N_1479);
nand U4840 (N_4840,N_1363,N_1611);
and U4841 (N_4841,N_1189,N_1126);
and U4842 (N_4842,N_2460,N_2289);
and U4843 (N_4843,N_1746,N_114);
or U4844 (N_4844,N_1750,N_2323);
nand U4845 (N_4845,N_2266,N_1082);
xor U4846 (N_4846,N_1654,N_2390);
nand U4847 (N_4847,N_1601,N_2326);
and U4848 (N_4848,N_2279,N_1141);
or U4849 (N_4849,N_22,N_579);
nor U4850 (N_4850,N_831,N_1096);
nor U4851 (N_4851,N_777,N_1678);
and U4852 (N_4852,N_579,N_163);
or U4853 (N_4853,N_1843,N_1675);
and U4854 (N_4854,N_335,N_1777);
nand U4855 (N_4855,N_1407,N_1418);
and U4856 (N_4856,N_1264,N_845);
or U4857 (N_4857,N_2246,N_2368);
and U4858 (N_4858,N_432,N_938);
nand U4859 (N_4859,N_170,N_1890);
or U4860 (N_4860,N_1670,N_636);
or U4861 (N_4861,N_1466,N_1489);
xnor U4862 (N_4862,N_923,N_2162);
or U4863 (N_4863,N_2491,N_2217);
nand U4864 (N_4864,N_1540,N_178);
nor U4865 (N_4865,N_1915,N_1627);
or U4866 (N_4866,N_1304,N_1376);
and U4867 (N_4867,N_768,N_164);
nand U4868 (N_4868,N_1048,N_1355);
or U4869 (N_4869,N_1602,N_2239);
and U4870 (N_4870,N_1661,N_642);
nand U4871 (N_4871,N_2104,N_1828);
and U4872 (N_4872,N_359,N_1430);
nand U4873 (N_4873,N_2410,N_2371);
nor U4874 (N_4874,N_77,N_523);
nand U4875 (N_4875,N_1667,N_244);
or U4876 (N_4876,N_341,N_1051);
xnor U4877 (N_4877,N_1293,N_1303);
nand U4878 (N_4878,N_2065,N_387);
or U4879 (N_4879,N_1069,N_110);
and U4880 (N_4880,N_311,N_771);
and U4881 (N_4881,N_1690,N_621);
and U4882 (N_4882,N_1625,N_994);
and U4883 (N_4883,N_974,N_1791);
nor U4884 (N_4884,N_485,N_883);
nor U4885 (N_4885,N_627,N_243);
or U4886 (N_4886,N_865,N_2162);
or U4887 (N_4887,N_281,N_2198);
xnor U4888 (N_4888,N_890,N_1646);
or U4889 (N_4889,N_830,N_1700);
nand U4890 (N_4890,N_2468,N_1393);
and U4891 (N_4891,N_1261,N_2172);
nand U4892 (N_4892,N_2011,N_2288);
nand U4893 (N_4893,N_373,N_288);
nor U4894 (N_4894,N_1789,N_1291);
and U4895 (N_4895,N_521,N_571);
or U4896 (N_4896,N_1147,N_2355);
and U4897 (N_4897,N_1560,N_905);
nand U4898 (N_4898,N_818,N_1278);
or U4899 (N_4899,N_2402,N_331);
and U4900 (N_4900,N_1870,N_412);
nor U4901 (N_4901,N_2067,N_1667);
xor U4902 (N_4902,N_1401,N_1222);
nor U4903 (N_4903,N_1246,N_223);
or U4904 (N_4904,N_1686,N_2441);
or U4905 (N_4905,N_100,N_2031);
and U4906 (N_4906,N_670,N_662);
nand U4907 (N_4907,N_64,N_228);
nor U4908 (N_4908,N_2333,N_425);
nor U4909 (N_4909,N_905,N_2287);
and U4910 (N_4910,N_273,N_2478);
nand U4911 (N_4911,N_763,N_2375);
nand U4912 (N_4912,N_2194,N_926);
nand U4913 (N_4913,N_20,N_390);
nor U4914 (N_4914,N_1139,N_2477);
and U4915 (N_4915,N_1045,N_1613);
or U4916 (N_4916,N_183,N_2236);
and U4917 (N_4917,N_1812,N_1361);
nand U4918 (N_4918,N_251,N_894);
nor U4919 (N_4919,N_2039,N_2103);
or U4920 (N_4920,N_2162,N_629);
and U4921 (N_4921,N_1242,N_515);
and U4922 (N_4922,N_373,N_2048);
or U4923 (N_4923,N_342,N_1504);
nand U4924 (N_4924,N_1214,N_153);
nor U4925 (N_4925,N_2027,N_705);
nand U4926 (N_4926,N_1285,N_1866);
nor U4927 (N_4927,N_2202,N_1952);
nand U4928 (N_4928,N_1843,N_401);
nand U4929 (N_4929,N_1641,N_1605);
nand U4930 (N_4930,N_928,N_396);
or U4931 (N_4931,N_982,N_586);
nor U4932 (N_4932,N_121,N_2365);
nand U4933 (N_4933,N_1996,N_802);
and U4934 (N_4934,N_1751,N_2430);
nor U4935 (N_4935,N_2174,N_18);
nand U4936 (N_4936,N_2132,N_566);
or U4937 (N_4937,N_2085,N_1079);
or U4938 (N_4938,N_1748,N_1574);
nand U4939 (N_4939,N_321,N_447);
and U4940 (N_4940,N_485,N_1182);
and U4941 (N_4941,N_2454,N_1931);
xor U4942 (N_4942,N_1105,N_2492);
or U4943 (N_4943,N_850,N_2418);
and U4944 (N_4944,N_1517,N_1295);
nand U4945 (N_4945,N_677,N_1081);
or U4946 (N_4946,N_1661,N_1931);
or U4947 (N_4947,N_2085,N_1136);
nor U4948 (N_4948,N_2212,N_2171);
or U4949 (N_4949,N_2106,N_1893);
nor U4950 (N_4950,N_545,N_1952);
nor U4951 (N_4951,N_868,N_1091);
nor U4952 (N_4952,N_709,N_1589);
nor U4953 (N_4953,N_6,N_2420);
nand U4954 (N_4954,N_139,N_2175);
nor U4955 (N_4955,N_1133,N_2116);
and U4956 (N_4956,N_655,N_2019);
nand U4957 (N_4957,N_787,N_2201);
nand U4958 (N_4958,N_84,N_1847);
nand U4959 (N_4959,N_639,N_2060);
or U4960 (N_4960,N_967,N_1776);
and U4961 (N_4961,N_1619,N_220);
or U4962 (N_4962,N_1620,N_2435);
nand U4963 (N_4963,N_350,N_1279);
or U4964 (N_4964,N_109,N_1562);
or U4965 (N_4965,N_1700,N_1149);
and U4966 (N_4966,N_59,N_167);
or U4967 (N_4967,N_1833,N_781);
and U4968 (N_4968,N_1102,N_1578);
nor U4969 (N_4969,N_158,N_2437);
nand U4970 (N_4970,N_2410,N_123);
nand U4971 (N_4971,N_193,N_397);
and U4972 (N_4972,N_350,N_2371);
nand U4973 (N_4973,N_662,N_1842);
nand U4974 (N_4974,N_1946,N_513);
nand U4975 (N_4975,N_1126,N_2394);
and U4976 (N_4976,N_1781,N_233);
nand U4977 (N_4977,N_1799,N_1249);
nand U4978 (N_4978,N_1542,N_1176);
nor U4979 (N_4979,N_1990,N_501);
and U4980 (N_4980,N_2406,N_858);
nor U4981 (N_4981,N_343,N_1185);
or U4982 (N_4982,N_1242,N_2177);
nor U4983 (N_4983,N_504,N_1743);
and U4984 (N_4984,N_26,N_1826);
nand U4985 (N_4985,N_2311,N_2078);
nand U4986 (N_4986,N_586,N_2420);
nor U4987 (N_4987,N_1788,N_2068);
nor U4988 (N_4988,N_162,N_2361);
nand U4989 (N_4989,N_1455,N_238);
nand U4990 (N_4990,N_323,N_2391);
nand U4991 (N_4991,N_289,N_997);
nand U4992 (N_4992,N_1006,N_30);
and U4993 (N_4993,N_568,N_2427);
nand U4994 (N_4994,N_309,N_2188);
or U4995 (N_4995,N_1083,N_1657);
nand U4996 (N_4996,N_433,N_490);
and U4997 (N_4997,N_1765,N_512);
nand U4998 (N_4998,N_1023,N_1782);
or U4999 (N_4999,N_795,N_2088);
and U5000 (N_5000,N_3692,N_3841);
nor U5001 (N_5001,N_3563,N_3582);
or U5002 (N_5002,N_2541,N_4190);
nand U5003 (N_5003,N_2947,N_4574);
nand U5004 (N_5004,N_4445,N_4439);
or U5005 (N_5005,N_2914,N_4284);
nand U5006 (N_5006,N_2895,N_3088);
or U5007 (N_5007,N_4207,N_3220);
nand U5008 (N_5008,N_2856,N_4116);
or U5009 (N_5009,N_4538,N_3015);
or U5010 (N_5010,N_3074,N_3596);
nor U5011 (N_5011,N_4587,N_3910);
nor U5012 (N_5012,N_4966,N_4949);
xnor U5013 (N_5013,N_4550,N_2571);
nand U5014 (N_5014,N_3265,N_3800);
or U5015 (N_5015,N_4200,N_3001);
or U5016 (N_5016,N_2765,N_4972);
nand U5017 (N_5017,N_4760,N_3566);
and U5018 (N_5018,N_3702,N_3521);
or U5019 (N_5019,N_3039,N_3558);
nand U5020 (N_5020,N_3972,N_4716);
and U5021 (N_5021,N_3327,N_3895);
or U5022 (N_5022,N_3962,N_4344);
or U5023 (N_5023,N_2964,N_2702);
and U5024 (N_5024,N_3365,N_4629);
and U5025 (N_5025,N_3609,N_3701);
or U5026 (N_5026,N_2602,N_3258);
or U5027 (N_5027,N_4916,N_3241);
nand U5028 (N_5028,N_3257,N_4230);
and U5029 (N_5029,N_4301,N_2645);
nand U5030 (N_5030,N_3635,N_3380);
or U5031 (N_5031,N_4479,N_3976);
xnor U5032 (N_5032,N_4177,N_4502);
nor U5033 (N_5033,N_4110,N_3330);
and U5034 (N_5034,N_4299,N_4012);
nand U5035 (N_5035,N_4072,N_3648);
and U5036 (N_5036,N_4215,N_4578);
or U5037 (N_5037,N_3634,N_3815);
nand U5038 (N_5038,N_4179,N_3913);
nor U5039 (N_5039,N_2787,N_3764);
and U5040 (N_5040,N_4957,N_4768);
and U5041 (N_5041,N_2807,N_3819);
nor U5042 (N_5042,N_3126,N_3967);
and U5043 (N_5043,N_4710,N_4310);
and U5044 (N_5044,N_2565,N_4671);
or U5045 (N_5045,N_4311,N_3051);
and U5046 (N_5046,N_4562,N_4240);
and U5047 (N_5047,N_2951,N_3921);
or U5048 (N_5048,N_2705,N_2508);
nor U5049 (N_5049,N_4324,N_4241);
and U5050 (N_5050,N_2804,N_3750);
and U5051 (N_5051,N_2784,N_2683);
and U5052 (N_5052,N_3813,N_2762);
or U5053 (N_5053,N_2976,N_2775);
or U5054 (N_5054,N_2818,N_3210);
nand U5055 (N_5055,N_3970,N_3031);
or U5056 (N_5056,N_3577,N_4471);
or U5057 (N_5057,N_3687,N_3636);
and U5058 (N_5058,N_4199,N_3314);
or U5059 (N_5059,N_4802,N_4016);
nor U5060 (N_5060,N_4764,N_4547);
and U5061 (N_5061,N_4836,N_4840);
and U5062 (N_5062,N_4314,N_3085);
or U5063 (N_5063,N_2922,N_3419);
and U5064 (N_5064,N_4658,N_3584);
and U5065 (N_5065,N_3698,N_3357);
nor U5066 (N_5066,N_2939,N_4295);
nor U5067 (N_5067,N_4358,N_4431);
and U5068 (N_5068,N_4633,N_3517);
nand U5069 (N_5069,N_3403,N_2531);
nor U5070 (N_5070,N_4473,N_4615);
xor U5071 (N_5071,N_3952,N_2831);
nor U5072 (N_5072,N_2962,N_3338);
nand U5073 (N_5073,N_2641,N_3850);
and U5074 (N_5074,N_4742,N_2734);
or U5075 (N_5075,N_4443,N_4154);
nor U5076 (N_5076,N_2603,N_3547);
xor U5077 (N_5077,N_3756,N_4156);
and U5078 (N_5078,N_3623,N_4937);
and U5079 (N_5079,N_2551,N_3765);
nand U5080 (N_5080,N_3509,N_3513);
and U5081 (N_5081,N_2696,N_4481);
and U5082 (N_5082,N_3475,N_4968);
and U5083 (N_5083,N_3653,N_4078);
nand U5084 (N_5084,N_2830,N_4076);
and U5085 (N_5085,N_3744,N_3390);
or U5086 (N_5086,N_3736,N_3591);
nand U5087 (N_5087,N_4498,N_3546);
or U5088 (N_5088,N_4372,N_3905);
nor U5089 (N_5089,N_4999,N_3575);
nand U5090 (N_5090,N_4506,N_3574);
nor U5091 (N_5091,N_3460,N_3199);
or U5092 (N_5092,N_4023,N_4721);
nor U5093 (N_5093,N_3725,N_3416);
nor U5094 (N_5094,N_2644,N_4341);
nor U5095 (N_5095,N_4756,N_4083);
and U5096 (N_5096,N_3873,N_4720);
or U5097 (N_5097,N_3483,N_4149);
and U5098 (N_5098,N_4420,N_3649);
and U5099 (N_5099,N_4128,N_3222);
or U5100 (N_5100,N_2869,N_4987);
nand U5101 (N_5101,N_2526,N_3068);
nand U5102 (N_5102,N_3105,N_4531);
nor U5103 (N_5103,N_2957,N_4360);
or U5104 (N_5104,N_2952,N_3762);
nand U5105 (N_5105,N_4278,N_2796);
or U5106 (N_5106,N_3614,N_3758);
or U5107 (N_5107,N_4159,N_3511);
or U5108 (N_5108,N_4981,N_4713);
and U5109 (N_5109,N_2991,N_4660);
nor U5110 (N_5110,N_4307,N_3735);
or U5111 (N_5111,N_3543,N_4090);
nand U5112 (N_5112,N_3919,N_3134);
nor U5113 (N_5113,N_3333,N_3971);
nor U5114 (N_5114,N_4490,N_4670);
nor U5115 (N_5115,N_3122,N_4799);
nand U5116 (N_5116,N_4034,N_3185);
or U5117 (N_5117,N_2662,N_2695);
nand U5118 (N_5118,N_4487,N_3337);
or U5119 (N_5119,N_3766,N_2623);
nor U5120 (N_5120,N_3072,N_4189);
nand U5121 (N_5121,N_3718,N_4938);
nand U5122 (N_5122,N_3035,N_2988);
and U5123 (N_5123,N_4218,N_3354);
nor U5124 (N_5124,N_4061,N_3731);
and U5125 (N_5125,N_4349,N_4913);
and U5126 (N_5126,N_2766,N_4326);
and U5127 (N_5127,N_3515,N_3722);
xor U5128 (N_5128,N_3070,N_2670);
or U5129 (N_5129,N_4375,N_2640);
nand U5130 (N_5130,N_3128,N_4219);
nor U5131 (N_5131,N_3121,N_4681);
nor U5132 (N_5132,N_2534,N_3352);
and U5133 (N_5133,N_4874,N_4781);
nand U5134 (N_5134,N_3046,N_3530);
nor U5135 (N_5135,N_4141,N_4109);
or U5136 (N_5136,N_4252,N_2607);
and U5137 (N_5137,N_2965,N_3429);
or U5138 (N_5138,N_3748,N_2995);
nor U5139 (N_5139,N_3805,N_4458);
nand U5140 (N_5140,N_4108,N_3422);
nor U5141 (N_5141,N_2652,N_2944);
nor U5142 (N_5142,N_3441,N_2715);
nor U5143 (N_5143,N_4440,N_4955);
or U5144 (N_5144,N_2763,N_2559);
nor U5145 (N_5145,N_4889,N_3379);
nand U5146 (N_5146,N_4530,N_4791);
nand U5147 (N_5147,N_4551,N_4075);
nor U5148 (N_5148,N_4350,N_4488);
and U5149 (N_5149,N_3440,N_4235);
and U5150 (N_5150,N_3524,N_2890);
and U5151 (N_5151,N_3037,N_3545);
nand U5152 (N_5152,N_4146,N_2554);
and U5153 (N_5153,N_3418,N_4323);
or U5154 (N_5154,N_4185,N_3217);
and U5155 (N_5155,N_3172,N_4804);
or U5156 (N_5156,N_3137,N_3025);
and U5157 (N_5157,N_4208,N_3902);
nand U5158 (N_5158,N_3116,N_3969);
and U5159 (N_5159,N_3709,N_4648);
nand U5160 (N_5160,N_4242,N_4160);
nor U5161 (N_5161,N_4514,N_4279);
and U5162 (N_5162,N_2798,N_3657);
or U5163 (N_5163,N_3620,N_3627);
nand U5164 (N_5164,N_4413,N_3784);
and U5165 (N_5165,N_3983,N_3360);
and U5166 (N_5166,N_4707,N_3401);
nand U5167 (N_5167,N_3339,N_3048);
and U5168 (N_5168,N_4205,N_4948);
and U5169 (N_5169,N_4294,N_4539);
and U5170 (N_5170,N_4665,N_3270);
and U5171 (N_5171,N_3716,N_3562);
nand U5172 (N_5172,N_4113,N_2797);
or U5173 (N_5173,N_4784,N_4446);
and U5174 (N_5174,N_4745,N_4120);
or U5175 (N_5175,N_3256,N_3892);
xor U5176 (N_5176,N_2916,N_2870);
xor U5177 (N_5177,N_3526,N_3186);
nand U5178 (N_5178,N_4591,N_4053);
or U5179 (N_5179,N_4359,N_2675);
and U5180 (N_5180,N_4903,N_4818);
nand U5181 (N_5181,N_2679,N_3277);
nand U5182 (N_5182,N_3573,N_3606);
nor U5183 (N_5183,N_2823,N_2989);
or U5184 (N_5184,N_3950,N_3468);
nor U5185 (N_5185,N_2799,N_3166);
nand U5186 (N_5186,N_4717,N_4673);
and U5187 (N_5187,N_4123,N_4521);
and U5188 (N_5188,N_3005,N_4563);
nand U5189 (N_5189,N_4610,N_3294);
nand U5190 (N_5190,N_4543,N_3908);
and U5191 (N_5191,N_4398,N_3041);
or U5192 (N_5192,N_3009,N_4317);
or U5193 (N_5193,N_3073,N_2758);
nand U5194 (N_5194,N_2538,N_4942);
nor U5195 (N_5195,N_4368,N_2584);
and U5196 (N_5196,N_3130,N_4489);
nor U5197 (N_5197,N_3943,N_4693);
nand U5198 (N_5198,N_2953,N_3664);
or U5199 (N_5199,N_4139,N_3164);
nor U5200 (N_5200,N_4203,N_3303);
nand U5201 (N_5201,N_3020,N_2616);
nand U5202 (N_5202,N_3922,N_4478);
nor U5203 (N_5203,N_4599,N_2615);
or U5204 (N_5204,N_4366,N_3506);
nor U5205 (N_5205,N_2691,N_2637);
nand U5206 (N_5206,N_4831,N_3274);
nand U5207 (N_5207,N_3486,N_4698);
nand U5208 (N_5208,N_4211,N_4391);
nor U5209 (N_5209,N_2707,N_3114);
and U5210 (N_5210,N_3733,N_2908);
and U5211 (N_5211,N_3925,N_4724);
nor U5212 (N_5212,N_2808,N_2658);
nor U5213 (N_5213,N_3848,N_3481);
or U5214 (N_5214,N_4003,N_2813);
or U5215 (N_5215,N_3436,N_4722);
nand U5216 (N_5216,N_2923,N_4608);
or U5217 (N_5217,N_2896,N_3686);
nor U5218 (N_5218,N_4404,N_3696);
nand U5219 (N_5219,N_2879,N_2848);
and U5220 (N_5220,N_3890,N_3102);
nand U5221 (N_5221,N_4603,N_4168);
nand U5222 (N_5222,N_3231,N_3299);
or U5223 (N_5223,N_2913,N_4151);
nand U5224 (N_5224,N_3537,N_3125);
nor U5225 (N_5225,N_3615,N_3196);
or U5226 (N_5226,N_3998,N_4223);
nand U5227 (N_5227,N_3098,N_2669);
nor U5228 (N_5228,N_4465,N_4825);
nand U5229 (N_5229,N_4259,N_4546);
and U5230 (N_5230,N_4354,N_4523);
nor U5231 (N_5231,N_3449,N_3342);
nor U5232 (N_5232,N_2732,N_4320);
nor U5233 (N_5233,N_4773,N_3302);
or U5234 (N_5234,N_3236,N_3531);
or U5235 (N_5235,N_4340,N_4632);
and U5236 (N_5236,N_3221,N_4965);
nor U5237 (N_5237,N_3000,N_3180);
nor U5238 (N_5238,N_3508,N_2532);
and U5239 (N_5239,N_4056,N_2912);
or U5240 (N_5240,N_3893,N_3592);
nand U5241 (N_5241,N_3789,N_3938);
nor U5242 (N_5242,N_3737,N_3229);
nor U5243 (N_5243,N_3611,N_3714);
or U5244 (N_5244,N_4272,N_3108);
nand U5245 (N_5245,N_4424,N_4196);
and U5246 (N_5246,N_4244,N_3152);
or U5247 (N_5247,N_3927,N_2588);
and U5248 (N_5248,N_4650,N_2979);
or U5249 (N_5249,N_4654,N_3228);
or U5250 (N_5250,N_4726,N_2780);
xnor U5251 (N_5251,N_2751,N_4678);
nand U5252 (N_5252,N_3979,N_4807);
and U5253 (N_5253,N_3064,N_4923);
or U5254 (N_5254,N_3684,N_3366);
nand U5255 (N_5255,N_3851,N_2997);
nand U5256 (N_5256,N_3055,N_4866);
nand U5257 (N_5257,N_3344,N_3183);
nor U5258 (N_5258,N_3845,N_2873);
nor U5259 (N_5259,N_3995,N_2714);
and U5260 (N_5260,N_4985,N_2558);
or U5261 (N_5261,N_3630,N_3668);
or U5262 (N_5262,N_4518,N_3476);
nand U5263 (N_5263,N_3167,N_3456);
or U5264 (N_5264,N_3891,N_3008);
or U5265 (N_5265,N_2517,N_4653);
or U5266 (N_5266,N_3527,N_3960);
xnor U5267 (N_5267,N_2578,N_4017);
nor U5268 (N_5268,N_3580,N_4050);
nor U5269 (N_5269,N_3127,N_3631);
xnor U5270 (N_5270,N_3715,N_4125);
nor U5271 (N_5271,N_4191,N_3225);
nor U5272 (N_5272,N_4902,N_4730);
and U5273 (N_5273,N_3864,N_4007);
nor U5274 (N_5274,N_2598,N_4322);
nor U5275 (N_5275,N_4561,N_4793);
nand U5276 (N_5276,N_4672,N_4262);
xnor U5277 (N_5277,N_3856,N_3291);
nand U5278 (N_5278,N_4253,N_4345);
nor U5279 (N_5279,N_4117,N_3054);
nor U5280 (N_5280,N_4150,N_4997);
or U5281 (N_5281,N_2501,N_4312);
nor U5282 (N_5282,N_3305,N_3753);
or U5283 (N_5283,N_4695,N_3457);
or U5284 (N_5284,N_3141,N_3712);
nor U5285 (N_5285,N_2746,N_3024);
nand U5286 (N_5286,N_3151,N_3191);
nor U5287 (N_5287,N_3906,N_3143);
or U5288 (N_5288,N_4961,N_4361);
nor U5289 (N_5289,N_3802,N_3334);
and U5290 (N_5290,N_3651,N_3029);
nor U5291 (N_5291,N_3405,N_3315);
nor U5292 (N_5292,N_4402,N_2838);
and U5293 (N_5293,N_4735,N_3555);
or U5294 (N_5294,N_4765,N_2778);
or U5295 (N_5295,N_3233,N_3285);
nand U5296 (N_5296,N_3490,N_2561);
or U5297 (N_5297,N_4288,N_2841);
and U5298 (N_5298,N_2900,N_4048);
or U5299 (N_5299,N_3470,N_4060);
nand U5300 (N_5300,N_4459,N_4925);
or U5301 (N_5301,N_4347,N_4969);
nand U5302 (N_5302,N_4767,N_3540);
nand U5303 (N_5303,N_3706,N_2595);
nand U5304 (N_5304,N_2614,N_4798);
or U5305 (N_5305,N_3044,N_4777);
or U5306 (N_5306,N_4455,N_3017);
nor U5307 (N_5307,N_4754,N_2604);
nor U5308 (N_5308,N_4417,N_3188);
or U5309 (N_5309,N_3855,N_4757);
nand U5310 (N_5310,N_2833,N_4963);
nor U5311 (N_5311,N_3050,N_3487);
or U5312 (N_5312,N_4855,N_3309);
and U5313 (N_5313,N_3239,N_4265);
or U5314 (N_5314,N_4033,N_3433);
nand U5315 (N_5315,N_4983,N_4231);
or U5316 (N_5316,N_3947,N_3713);
and U5317 (N_5317,N_3259,N_2925);
nor U5318 (N_5318,N_2990,N_3688);
nand U5319 (N_5319,N_4255,N_2710);
and U5320 (N_5320,N_4581,N_3417);
and U5321 (N_5321,N_4096,N_4275);
and U5322 (N_5322,N_2546,N_4504);
and U5323 (N_5323,N_3570,N_2506);
or U5324 (N_5324,N_2993,N_2648);
nand U5325 (N_5325,N_4058,N_3830);
xnor U5326 (N_5326,N_2918,N_4163);
and U5327 (N_5327,N_4609,N_3432);
nor U5328 (N_5328,N_2627,N_3198);
or U5329 (N_5329,N_2949,N_3984);
or U5330 (N_5330,N_2694,N_3058);
nor U5331 (N_5331,N_4727,N_4484);
or U5332 (N_5332,N_2967,N_3811);
nor U5333 (N_5333,N_4032,N_3598);
nand U5334 (N_5334,N_4718,N_3625);
nor U5335 (N_5335,N_4881,N_3139);
nand U5336 (N_5336,N_2996,N_4512);
or U5337 (N_5337,N_2826,N_4332);
nand U5338 (N_5338,N_4316,N_2649);
and U5339 (N_5339,N_3884,N_3640);
or U5340 (N_5340,N_3226,N_2779);
nand U5341 (N_5341,N_3205,N_3187);
or U5342 (N_5342,N_4899,N_4351);
xor U5343 (N_5343,N_2851,N_4477);
or U5344 (N_5344,N_3341,N_3140);
or U5345 (N_5345,N_4100,N_3887);
and U5346 (N_5346,N_3768,N_4662);
nand U5347 (N_5347,N_3535,N_2803);
nand U5348 (N_5348,N_2864,N_2946);
or U5349 (N_5349,N_4140,N_3158);
nor U5350 (N_5350,N_4427,N_2629);
or U5351 (N_5351,N_4770,N_3792);
nand U5352 (N_5352,N_2611,N_2660);
nor U5353 (N_5353,N_4451,N_4254);
or U5354 (N_5354,N_2937,N_3437);
nand U5355 (N_5355,N_3292,N_4532);
nor U5356 (N_5356,N_4553,N_3103);
nand U5357 (N_5357,N_4811,N_4579);
nand U5358 (N_5358,N_2825,N_2866);
xor U5359 (N_5359,N_2688,N_2597);
nand U5360 (N_5360,N_4841,N_3556);
nand U5361 (N_5361,N_2843,N_2619);
nor U5362 (N_5362,N_3988,N_4469);
and U5363 (N_5363,N_3451,N_3942);
or U5364 (N_5364,N_2736,N_2786);
or U5365 (N_5365,N_2885,N_4444);
or U5366 (N_5366,N_3016,N_3473);
or U5367 (N_5367,N_4751,N_3425);
nor U5368 (N_5368,N_3557,N_3377);
or U5369 (N_5369,N_4256,N_4495);
or U5370 (N_5370,N_3107,N_3328);
and U5371 (N_5371,N_4456,N_4021);
xnor U5372 (N_5372,N_4950,N_3915);
and U5373 (N_5373,N_3773,N_4704);
or U5374 (N_5374,N_4094,N_2567);
nor U5375 (N_5375,N_4575,N_3175);
nor U5376 (N_5376,N_3464,N_4143);
or U5377 (N_5377,N_4769,N_3797);
or U5378 (N_5378,N_2522,N_2661);
or U5379 (N_5379,N_3312,N_3383);
and U5380 (N_5380,N_3230,N_2840);
or U5381 (N_5381,N_4858,N_4434);
nor U5382 (N_5382,N_4908,N_3525);
and U5383 (N_5383,N_3790,N_3710);
or U5384 (N_5384,N_2739,N_3154);
or U5385 (N_5385,N_4812,N_4181);
xnor U5386 (N_5386,N_3522,N_3002);
or U5387 (N_5387,N_4264,N_3497);
nand U5388 (N_5388,N_3385,N_3280);
or U5389 (N_5389,N_2950,N_4921);
and U5390 (N_5390,N_4386,N_3565);
nor U5391 (N_5391,N_2577,N_4865);
nand U5392 (N_5392,N_4257,N_4849);
and U5393 (N_5393,N_3963,N_3301);
nand U5394 (N_5394,N_2579,N_4709);
or U5395 (N_5395,N_3430,N_2545);
nor U5396 (N_5396,N_3959,N_2543);
or U5397 (N_5397,N_4343,N_3694);
and U5398 (N_5398,N_4584,N_4302);
nand U5399 (N_5399,N_2789,N_4862);
and U5400 (N_5400,N_3160,N_4043);
and U5401 (N_5401,N_2897,N_3348);
nor U5402 (N_5402,N_4336,N_3491);
nor U5403 (N_5403,N_3268,N_4732);
nor U5404 (N_5404,N_3153,N_4492);
and U5405 (N_5405,N_3992,N_4001);
or U5406 (N_5406,N_4321,N_4663);
or U5407 (N_5407,N_3289,N_3184);
or U5408 (N_5408,N_4127,N_3656);
xor U5409 (N_5409,N_4843,N_4863);
or U5410 (N_5410,N_4576,N_3082);
or U5411 (N_5411,N_4882,N_4900);
or U5412 (N_5412,N_4623,N_4292);
and U5413 (N_5413,N_3479,N_4984);
nor U5414 (N_5414,N_4099,N_2749);
or U5415 (N_5415,N_3168,N_2956);
nand U5416 (N_5416,N_4565,N_4787);
or U5417 (N_5417,N_3597,N_3837);
nand U5418 (N_5418,N_2972,N_3655);
nor U5419 (N_5419,N_3165,N_4619);
xnor U5420 (N_5420,N_4379,N_3804);
nor U5421 (N_5421,N_4612,N_3071);
nor U5422 (N_5422,N_4683,N_4731);
and U5423 (N_5423,N_2899,N_2664);
and U5424 (N_5424,N_4276,N_2580);
nor U5425 (N_5425,N_4912,N_2819);
and U5426 (N_5426,N_4069,N_3707);
or U5427 (N_5427,N_2617,N_4197);
nand U5428 (N_5428,N_3269,N_2729);
nand U5429 (N_5429,N_3842,N_4801);
and U5430 (N_5430,N_3129,N_3261);
nor U5431 (N_5431,N_2980,N_3662);
xor U5432 (N_5432,N_3548,N_3823);
and U5433 (N_5433,N_3325,N_4946);
nor U5434 (N_5434,N_4119,N_3727);
nor U5435 (N_5435,N_3695,N_4210);
and U5436 (N_5436,N_3982,N_3964);
and U5437 (N_5437,N_4442,N_4233);
or U5438 (N_5438,N_4714,N_3672);
nand U5439 (N_5439,N_4148,N_2788);
and U5440 (N_5440,N_4030,N_3903);
nand U5441 (N_5441,N_3306,N_2504);
nor U5442 (N_5442,N_3881,N_3489);
and U5443 (N_5443,N_3512,N_4212);
nor U5444 (N_5444,N_3788,N_4385);
nor U5445 (N_5445,N_4407,N_4277);
or U5446 (N_5446,N_4982,N_2777);
nor U5447 (N_5447,N_3032,N_3026);
and U5448 (N_5448,N_4228,N_2785);
and U5449 (N_5449,N_4137,N_3414);
nor U5450 (N_5450,N_4848,N_3538);
and U5451 (N_5451,N_2936,N_2893);
or U5452 (N_5452,N_3595,N_4271);
nand U5453 (N_5453,N_4180,N_4826);
nor U5454 (N_5454,N_2791,N_4377);
and U5455 (N_5455,N_4037,N_3931);
nor U5456 (N_5456,N_2839,N_2687);
or U5457 (N_5457,N_4897,N_2735);
or U5458 (N_5458,N_2753,N_3858);
or U5459 (N_5459,N_3358,N_4071);
nand U5460 (N_5460,N_2750,N_4805);
nand U5461 (N_5461,N_4809,N_4187);
xnor U5462 (N_5462,N_2631,N_4669);
nor U5463 (N_5463,N_2906,N_4869);
nand U5464 (N_5464,N_3742,N_4416);
nor U5465 (N_5465,N_4851,N_2511);
and U5466 (N_5466,N_4047,N_3590);
nand U5467 (N_5467,N_3359,N_3373);
xnor U5468 (N_5468,N_3743,N_4186);
nor U5469 (N_5469,N_4059,N_4298);
nand U5470 (N_5470,N_3136,N_4970);
nor U5471 (N_5471,N_2570,N_3307);
nand U5472 (N_5472,N_2700,N_2984);
and U5473 (N_5473,N_4701,N_3260);
nand U5474 (N_5474,N_3104,N_2889);
and U5475 (N_5475,N_4815,N_2608);
or U5476 (N_5476,N_3946,N_4261);
and U5477 (N_5477,N_3571,N_2883);
and U5478 (N_5478,N_3674,N_3587);
or U5479 (N_5479,N_4860,N_4646);
nor U5480 (N_5480,N_4183,N_4640);
or U5481 (N_5481,N_4232,N_4741);
and U5482 (N_5482,N_3398,N_4018);
nand U5483 (N_5483,N_4676,N_3682);
nand U5484 (N_5484,N_2902,N_3423);
or U5485 (N_5485,N_3162,N_2673);
nor U5486 (N_5486,N_4333,N_4328);
and U5487 (N_5487,N_2858,N_4536);
xor U5488 (N_5488,N_3459,N_3639);
and U5489 (N_5489,N_3415,N_3948);
nand U5490 (N_5490,N_3559,N_4064);
nand U5491 (N_5491,N_4833,N_3030);
and U5492 (N_5492,N_2963,N_3628);
nand U5493 (N_5493,N_4266,N_2888);
and U5494 (N_5494,N_4503,N_4789);
nand U5495 (N_5495,N_2709,N_2942);
or U5496 (N_5496,N_4414,N_4480);
and U5497 (N_5497,N_4178,N_4087);
and U5498 (N_5498,N_4423,N_2754);
or U5499 (N_5499,N_2981,N_3397);
and U5500 (N_5500,N_4009,N_4637);
nor U5501 (N_5501,N_3019,N_3004);
and U5502 (N_5502,N_4878,N_3816);
and U5503 (N_5503,N_3897,N_4144);
nor U5504 (N_5504,N_3898,N_2668);
and U5505 (N_5505,N_4817,N_3721);
nor U5506 (N_5506,N_4237,N_4406);
or U5507 (N_5507,N_4457,N_3276);
and U5508 (N_5508,N_4392,N_3643);
and U5509 (N_5509,N_4622,N_3923);
and U5510 (N_5510,N_4935,N_3215);
nand U5511 (N_5511,N_2633,N_4904);
nand U5512 (N_5512,N_2657,N_4572);
nand U5513 (N_5513,N_3518,N_3677);
nor U5514 (N_5514,N_3472,N_3798);
nand U5515 (N_5515,N_4917,N_2549);
nand U5516 (N_5516,N_2663,N_2719);
nand U5517 (N_5517,N_3442,N_3202);
xnor U5518 (N_5518,N_3741,N_3111);
or U5519 (N_5519,N_4558,N_2612);
nor U5520 (N_5520,N_2628,N_3820);
and U5521 (N_5521,N_2795,N_3586);
nor U5522 (N_5522,N_4519,N_2790);
nor U5523 (N_5523,N_3617,N_4367);
nand U5524 (N_5524,N_4410,N_2844);
nor U5525 (N_5525,N_3387,N_4258);
or U5526 (N_5526,N_4157,N_4689);
nand U5527 (N_5527,N_4753,N_4962);
nand U5528 (N_5528,N_3994,N_2971);
nor U5529 (N_5529,N_4967,N_4651);
and U5530 (N_5530,N_2666,N_4898);
nor U5531 (N_5531,N_3945,N_3266);
nor U5532 (N_5532,N_2639,N_3496);
nor U5533 (N_5533,N_4039,N_4004);
xnor U5534 (N_5534,N_2832,N_3859);
nor U5535 (N_5535,N_4454,N_4499);
or U5536 (N_5536,N_4387,N_4290);
or U5537 (N_5537,N_3917,N_3142);
and U5538 (N_5538,N_4887,N_2575);
nand U5539 (N_5539,N_2516,N_2920);
or U5540 (N_5540,N_4854,N_2745);
nor U5541 (N_5541,N_3059,N_2881);
or U5542 (N_5542,N_4062,N_4373);
or U5543 (N_5543,N_3119,N_3282);
and U5544 (N_5544,N_3411,N_3323);
nor U5545 (N_5545,N_3243,N_3389);
nor U5546 (N_5546,N_3723,N_2651);
nand U5547 (N_5547,N_4535,N_4436);
nor U5548 (N_5548,N_4236,N_2593);
and U5549 (N_5549,N_3961,N_2805);
and U5550 (N_5550,N_4374,N_2926);
and U5551 (N_5551,N_4618,N_4652);
and U5552 (N_5552,N_2621,N_2835);
and U5553 (N_5553,N_2806,N_4540);
or U5554 (N_5554,N_4533,N_3138);
or U5555 (N_5555,N_2948,N_3149);
or U5556 (N_5556,N_4998,N_3427);
nand U5557 (N_5557,N_3928,N_3600);
nand U5558 (N_5558,N_2518,N_3090);
nor U5559 (N_5559,N_3870,N_3319);
nor U5560 (N_5560,N_4790,N_4752);
or U5561 (N_5561,N_4542,N_3224);
and U5562 (N_5562,N_4105,N_4174);
or U5563 (N_5563,N_3249,N_4118);
nand U5564 (N_5564,N_4960,N_3351);
nand U5565 (N_5565,N_4549,N_4002);
nand U5566 (N_5566,N_4428,N_3949);
nand U5567 (N_5567,N_4696,N_2672);
or U5568 (N_5568,N_2674,N_4607);
nand U5569 (N_5569,N_4711,N_4835);
nand U5570 (N_5570,N_2853,N_3219);
nand U5571 (N_5571,N_4524,N_4708);
or U5572 (N_5572,N_3212,N_4130);
nand U5573 (N_5573,N_3690,N_4990);
or U5574 (N_5574,N_2653,N_3331);
nand U5575 (N_5575,N_2523,N_4813);
nand U5576 (N_5576,N_2773,N_3083);
xor U5577 (N_5577,N_4461,N_3989);
nor U5578 (N_5578,N_3190,N_3255);
or U5579 (N_5579,N_3680,N_3271);
nor U5580 (N_5580,N_2748,N_4308);
or U5581 (N_5581,N_4422,N_3933);
nor U5582 (N_5582,N_3400,N_2875);
or U5583 (N_5583,N_3593,N_4852);
or U5584 (N_5584,N_4661,N_2690);
nand U5585 (N_5585,N_3067,N_3267);
or U5586 (N_5586,N_4226,N_3378);
or U5587 (N_5587,N_3079,N_3854);
nor U5588 (N_5588,N_3608,N_4508);
nand U5589 (N_5589,N_4613,N_3552);
nand U5590 (N_5590,N_3438,N_3364);
or U5591 (N_5591,N_2836,N_3853);
and U5592 (N_5592,N_3699,N_4074);
and U5593 (N_5593,N_4247,N_2594);
or U5594 (N_5594,N_4986,N_4112);
and U5595 (N_5595,N_3021,N_3754);
nor U5596 (N_5596,N_4621,N_3504);
or U5597 (N_5597,N_3978,N_3569);
or U5598 (N_5598,N_3831,N_4691);
xor U5599 (N_5599,N_3250,N_3076);
nor U5600 (N_5600,N_2528,N_3751);
nor U5601 (N_5601,N_3641,N_4520);
or U5602 (N_5602,N_2973,N_3987);
nor U5603 (N_5603,N_4892,N_4134);
nor U5604 (N_5604,N_2689,N_2966);
nor U5605 (N_5605,N_4274,N_3242);
or U5606 (N_5606,N_4931,N_4376);
nor U5607 (N_5607,N_2684,N_4082);
or U5608 (N_5608,N_4251,N_4055);
and U5609 (N_5609,N_4486,N_4111);
nor U5610 (N_5610,N_4555,N_4433);
or U5611 (N_5611,N_4657,N_4682);
or U5612 (N_5612,N_2929,N_3568);
or U5613 (N_5613,N_2548,N_2850);
or U5614 (N_5614,N_3028,N_2624);
and U5615 (N_5615,N_3145,N_3412);
or U5616 (N_5616,N_3719,N_3607);
and U5617 (N_5617,N_3528,N_3318);
and U5618 (N_5618,N_3332,N_4220);
or U5619 (N_5619,N_2665,N_3624);
and U5620 (N_5620,N_2891,N_2676);
nor U5621 (N_5621,N_3793,N_3874);
nand U5622 (N_5622,N_4225,N_4992);
nor U5623 (N_5623,N_4049,N_4054);
and U5624 (N_5624,N_2904,N_3238);
nand U5625 (N_5625,N_3404,N_4870);
nor U5626 (N_5626,N_2943,N_2605);
and U5627 (N_5627,N_3075,N_2986);
nor U5628 (N_5628,N_3095,N_3818);
nor U5629 (N_5629,N_4537,N_3161);
nor U5630 (N_5630,N_4677,N_2905);
nor U5631 (N_5631,N_2573,N_2898);
nor U5632 (N_5632,N_4951,N_4888);
or U5633 (N_5633,N_2977,N_4808);
nand U5634 (N_5634,N_4783,N_2829);
or U5635 (N_5635,N_2667,N_3036);
nand U5636 (N_5636,N_3394,N_3011);
or U5637 (N_5637,N_3954,N_4124);
and U5638 (N_5638,N_3685,N_4115);
nand U5639 (N_5639,N_4944,N_2978);
or U5640 (N_5640,N_3510,N_2718);
nor U5641 (N_5641,N_2635,N_3013);
or U5642 (N_5642,N_3311,N_3523);
or U5643 (N_5643,N_4856,N_2583);
and U5644 (N_5644,N_3621,N_2730);
or U5645 (N_5645,N_2919,N_3329);
nor U5646 (N_5646,N_4635,N_4859);
or U5647 (N_5647,N_2759,N_4857);
nand U5648 (N_5648,N_2582,N_2861);
nor U5649 (N_5649,N_4569,N_4926);
or U5650 (N_5650,N_2503,N_3739);
and U5651 (N_5651,N_3836,N_4725);
nand U5652 (N_5652,N_2550,N_2562);
nor U5653 (N_5653,N_2761,N_3860);
nor U5654 (N_5654,N_3638,N_3463);
and U5655 (N_5655,N_2638,N_3974);
nand U5656 (N_5656,N_2792,N_2959);
nor U5657 (N_5657,N_2568,N_4129);
nor U5658 (N_5658,N_4505,N_2728);
nor U5659 (N_5659,N_4517,N_4733);
nand U5660 (N_5660,N_2863,N_4327);
or U5661 (N_5661,N_3783,N_4959);
nand U5662 (N_5662,N_2774,N_2500);
or U5663 (N_5663,N_3878,N_4024);
nor U5664 (N_5664,N_4989,N_3700);
nand U5665 (N_5665,N_4873,N_2970);
and U5666 (N_5666,N_4822,N_4624);
nor U5667 (N_5667,N_4605,N_4580);
nand U5668 (N_5668,N_3033,N_3822);
nand U5669 (N_5669,N_4529,N_3388);
or U5670 (N_5670,N_4511,N_4705);
and U5671 (N_5671,N_4647,N_2915);
and U5672 (N_5672,N_4224,N_4089);
and U5673 (N_5673,N_3316,N_2509);
and U5674 (N_5674,N_3247,N_4821);
and U5675 (N_5675,N_2911,N_3336);
or U5676 (N_5676,N_4173,N_4883);
nor U5677 (N_5677,N_4474,N_3534);
nand U5678 (N_5678,N_3101,N_2505);
nand U5679 (N_5679,N_4772,N_3726);
nand U5680 (N_5680,N_3384,N_3730);
and U5681 (N_5681,N_3663,N_3066);
and U5682 (N_5682,N_4541,N_4029);
or U5683 (N_5683,N_2985,N_2969);
nor U5684 (N_5684,N_3894,N_2903);
and U5685 (N_5685,N_4304,N_4114);
nor U5686 (N_5686,N_2994,N_3814);
nand U5687 (N_5687,N_4245,N_3391);
nand U5688 (N_5688,N_4066,N_4877);
nand U5689 (N_5689,N_4463,N_3374);
or U5690 (N_5690,N_4107,N_4846);
nand U5691 (N_5691,N_3012,N_4890);
and U5692 (N_5692,N_2693,N_3431);
nand U5693 (N_5693,N_3616,N_3769);
or U5694 (N_5694,N_2723,N_3023);
and U5695 (N_5695,N_4092,N_4806);
and U5696 (N_5696,N_3482,N_4507);
and U5697 (N_5697,N_3827,N_2630);
xor U5698 (N_5698,N_4794,N_4052);
and U5699 (N_5699,N_3576,N_3421);
nor U5700 (N_5700,N_4132,N_4943);
nor U5701 (N_5701,N_2574,N_4248);
nand U5702 (N_5702,N_4842,N_4631);
or U5703 (N_5703,N_4911,N_3193);
or U5704 (N_5704,N_4106,N_4356);
and U5705 (N_5705,N_2656,N_4371);
nand U5706 (N_5706,N_3532,N_2907);
nor U5707 (N_5707,N_3581,N_4036);
nand U5708 (N_5708,N_3734,N_4102);
and U5709 (N_5709,N_4980,N_3356);
and U5710 (N_5710,N_3194,N_3899);
nand U5711 (N_5711,N_4552,N_3958);
nand U5712 (N_5712,N_4973,N_4166);
and U5713 (N_5713,N_3455,N_3375);
and U5714 (N_5714,N_4346,N_4194);
nor U5715 (N_5715,N_4920,N_4636);
nand U5716 (N_5716,N_2968,N_2521);
or U5717 (N_5717,N_3567,N_2770);
nand U5718 (N_5718,N_3133,N_4067);
nand U5719 (N_5719,N_4198,N_3977);
or U5720 (N_5720,N_3843,N_2556);
or U5721 (N_5721,N_2650,N_3022);
or U5722 (N_5722,N_2782,N_2744);
nor U5723 (N_5723,N_4079,N_3757);
nand U5724 (N_5724,N_3604,N_2880);
nand U5725 (N_5725,N_3560,N_4318);
and U5726 (N_5726,N_3287,N_4778);
and U5727 (N_5727,N_3087,N_4755);
or U5728 (N_5728,N_4357,N_2544);
or U5729 (N_5729,N_4135,N_4837);
nor U5730 (N_5730,N_4260,N_4467);
nand U5731 (N_5731,N_3370,N_3780);
or U5732 (N_5732,N_4483,N_2852);
and U5733 (N_5733,N_3665,N_3539);
and U5734 (N_5734,N_4595,N_2731);
and U5735 (N_5735,N_4872,N_4656);
or U5736 (N_5736,N_3924,N_4250);
nor U5737 (N_5737,N_4996,N_3610);
xnor U5738 (N_5738,N_3340,N_4639);
nor U5739 (N_5739,N_3078,N_2757);
nor U5740 (N_5740,N_2768,N_2682);
and U5741 (N_5741,N_2874,N_2620);
or U5742 (N_5742,N_4641,N_2576);
nor U5743 (N_5743,N_2960,N_3056);
or U5744 (N_5744,N_3500,N_3632);
nand U5745 (N_5745,N_3711,N_2917);
nand U5746 (N_5746,N_3561,N_4085);
or U5747 (N_5747,N_3918,N_4844);
nor U5748 (N_5748,N_3106,N_4161);
and U5749 (N_5749,N_3637,N_2824);
xnor U5750 (N_5750,N_2701,N_2846);
and U5751 (N_5751,N_2625,N_4091);
or U5752 (N_5752,N_3135,N_4974);
or U5753 (N_5753,N_3439,N_2820);
nand U5754 (N_5754,N_4093,N_2585);
nor U5755 (N_5755,N_3812,N_4234);
nor U5756 (N_5756,N_3791,N_3003);
nor U5757 (N_5757,N_3395,N_2828);
nand U5758 (N_5758,N_3738,N_4666);
nand U5759 (N_5759,N_3443,N_4723);
nor U5760 (N_5760,N_4147,N_2586);
nand U5761 (N_5761,N_3262,N_2814);
nor U5762 (N_5762,N_2961,N_3112);
or U5763 (N_5763,N_4325,N_4988);
nor U5764 (N_5764,N_4249,N_4476);
nand U5765 (N_5765,N_3355,N_3650);
or U5766 (N_5766,N_4918,N_4209);
nor U5767 (N_5767,N_3264,N_4577);
or U5768 (N_5768,N_3626,N_3669);
nand U5769 (N_5769,N_4330,N_3825);
and U5770 (N_5770,N_2941,N_3227);
or U5771 (N_5771,N_3092,N_3801);
nor U5772 (N_5772,N_2632,N_4411);
nor U5773 (N_5773,N_4894,N_4588);
nand U5774 (N_5774,N_4044,N_4940);
nand U5775 (N_5775,N_3888,N_2865);
and U5776 (N_5776,N_3728,N_2933);
nand U5777 (N_5777,N_3179,N_3503);
or U5778 (N_5778,N_4516,N_2622);
nand U5779 (N_5779,N_3755,N_2747);
and U5780 (N_5780,N_4932,N_4070);
nand U5781 (N_5781,N_3246,N_3644);
nor U5782 (N_5782,N_4399,N_4293);
or U5783 (N_5783,N_3096,N_3296);
and U5784 (N_5784,N_3350,N_4206);
nand U5785 (N_5785,N_4281,N_4626);
nand U5786 (N_5786,N_3880,N_4401);
or U5787 (N_5787,N_4885,N_3089);
or U5788 (N_5788,N_4616,N_4828);
or U5789 (N_5789,N_3049,N_2983);
nor U5790 (N_5790,N_4570,N_4785);
or U5791 (N_5791,N_3675,N_3434);
and U5792 (N_5792,N_4644,N_4684);
and U5793 (N_5793,N_2533,N_4627);
nand U5794 (N_5794,N_4832,N_3466);
and U5795 (N_5795,N_4782,N_3424);
nor U5796 (N_5796,N_3392,N_3579);
or U5797 (N_5797,N_4405,N_2564);
nand U5798 (N_5798,N_3216,N_4025);
nand U5799 (N_5799,N_2581,N_4246);
nand U5800 (N_5800,N_3697,N_4421);
nand U5801 (N_5801,N_4338,N_3683);
nand U5802 (N_5802,N_3501,N_4081);
or U5803 (N_5803,N_4133,N_4045);
or U5804 (N_5804,N_3251,N_3297);
and U5805 (N_5805,N_4762,N_3985);
nand U5806 (N_5806,N_3951,N_3907);
or U5807 (N_5807,N_2886,N_3321);
or U5808 (N_5808,N_4396,N_3912);
nor U5809 (N_5809,N_3671,N_3803);
nand U5810 (N_5810,N_3746,N_4930);
nor U5811 (N_5811,N_3324,N_3045);
or U5812 (N_5812,N_3454,N_3155);
or U5813 (N_5813,N_4522,N_3794);
nand U5814 (N_5814,N_3148,N_4435);
nand U5815 (N_5815,N_3069,N_3467);
or U5816 (N_5816,N_2793,N_4214);
nor U5817 (N_5817,N_3189,N_4664);
or U5818 (N_5818,N_4006,N_4700);
nor U5819 (N_5819,N_3173,N_3605);
xnor U5820 (N_5820,N_2815,N_4152);
nand U5821 (N_5821,N_4839,N_3113);
or U5822 (N_5822,N_4450,N_4393);
or U5823 (N_5823,N_4868,N_3159);
nand U5824 (N_5824,N_3458,N_3968);
nand U5825 (N_5825,N_4491,N_4269);
or U5826 (N_5826,N_3882,N_4000);
and U5827 (N_5827,N_4065,N_3939);
nand U5828 (N_5828,N_4838,N_3551);
nor U5829 (N_5829,N_3806,N_4534);
and U5830 (N_5830,N_2932,N_3745);
and U5831 (N_5831,N_3629,N_3676);
or U5832 (N_5832,N_4509,N_3386);
and U5833 (N_5833,N_4780,N_3673);
nor U5834 (N_5834,N_3875,N_4419);
and U5835 (N_5835,N_4496,N_4786);
or U5836 (N_5836,N_4706,N_3040);
or U5837 (N_5837,N_4907,N_3776);
or U5838 (N_5838,N_4395,N_4008);
and U5839 (N_5839,N_3900,N_3647);
xnor U5840 (N_5840,N_4638,N_4747);
and U5841 (N_5841,N_3275,N_4121);
or U5842 (N_5842,N_4589,N_3957);
and U5843 (N_5843,N_2547,N_2887);
or U5844 (N_5844,N_3578,N_2877);
or U5845 (N_5845,N_3484,N_2884);
xnor U5846 (N_5846,N_3237,N_4412);
nor U5847 (N_5847,N_2636,N_4287);
or U5848 (N_5848,N_3123,N_4510);
or U5849 (N_5849,N_4680,N_4038);
nor U5850 (N_5850,N_2542,N_4861);
or U5851 (N_5851,N_4788,N_3223);
and U5852 (N_5852,N_4192,N_4131);
or U5853 (N_5853,N_4335,N_3176);
or U5854 (N_5854,N_4389,N_3871);
nor U5855 (N_5855,N_3828,N_2643);
nor U5856 (N_5856,N_4750,N_3322);
and U5857 (N_5857,N_3514,N_4567);
and U5858 (N_5858,N_3502,N_3399);
nand U5859 (N_5859,N_4922,N_4464);
xor U5860 (N_5860,N_3781,N_3826);
or U5861 (N_5861,N_3485,N_4797);
nor U5862 (N_5862,N_4545,N_2741);
nand U5863 (N_5863,N_4441,N_3209);
and U5864 (N_5864,N_2854,N_4901);
nand U5865 (N_5865,N_3146,N_3053);
or U5866 (N_5866,N_3885,N_3681);
nand U5867 (N_5867,N_3235,N_4329);
and U5868 (N_5868,N_2697,N_4353);
or U5869 (N_5869,N_4602,N_4686);
nand U5870 (N_5870,N_2706,N_2671);
nand U5871 (N_5871,N_4739,N_3426);
or U5872 (N_5872,N_4884,N_2760);
and U5873 (N_5873,N_2618,N_3298);
xor U5874 (N_5874,N_4667,N_4447);
nand U5875 (N_5875,N_4437,N_3435);
or U5876 (N_5876,N_4285,N_2992);
nor U5877 (N_5877,N_3785,N_3926);
nand U5878 (N_5878,N_4426,N_4614);
nand U5879 (N_5879,N_4557,N_4810);
and U5880 (N_5880,N_4175,N_4560);
or U5881 (N_5881,N_3810,N_3494);
or U5882 (N_5882,N_4014,N_4497);
or U5883 (N_5883,N_4564,N_4263);
nand U5884 (N_5884,N_4771,N_3174);
and U5885 (N_5885,N_4956,N_4734);
or U5886 (N_5886,N_2592,N_3886);
nand U5887 (N_5887,N_4694,N_3014);
nor U5888 (N_5888,N_3808,N_4544);
and U5889 (N_5889,N_3807,N_3038);
or U5890 (N_5890,N_3006,N_2982);
nand U5891 (N_5891,N_4649,N_4460);
or U5892 (N_5892,N_3505,N_3367);
and U5893 (N_5893,N_3081,N_3218);
nand U5894 (N_5894,N_2553,N_4697);
nand U5895 (N_5895,N_4462,N_4594);
or U5896 (N_5896,N_2999,N_3461);
nand U5897 (N_5897,N_3027,N_2871);
and U5898 (N_5898,N_4229,N_2512);
or U5899 (N_5899,N_3177,N_2601);
or U5900 (N_5900,N_4703,N_3667);
nor U5901 (N_5901,N_4712,N_4795);
or U5902 (N_5902,N_4086,N_2764);
nand U5903 (N_5903,N_2724,N_4296);
nand U5904 (N_5904,N_4600,N_3533);
and U5905 (N_5905,N_3761,N_2927);
or U5906 (N_5906,N_3368,N_4363);
and U5907 (N_5907,N_4743,N_2572);
and U5908 (N_5908,N_3195,N_2827);
or U5909 (N_5909,N_2536,N_3834);
and U5910 (N_5910,N_3865,N_2716);
nor U5911 (N_5911,N_3214,N_3263);
nand U5912 (N_5912,N_3200,N_3965);
nand U5913 (N_5913,N_4101,N_3795);
nand U5914 (N_5914,N_2599,N_3594);
nand U5915 (N_5915,N_2711,N_3920);
nand U5916 (N_5916,N_2708,N_3622);
or U5917 (N_5917,N_4606,N_4073);
nand U5918 (N_5918,N_3763,N_3660);
nand U5919 (N_5919,N_2699,N_4914);
and U5920 (N_5920,N_4850,N_2742);
and U5921 (N_5921,N_4403,N_4953);
or U5922 (N_5922,N_3062,N_4827);
and U5923 (N_5923,N_3310,N_2563);
or U5924 (N_5924,N_4515,N_3124);
or U5925 (N_5925,N_4630,N_2955);
or U5926 (N_5926,N_4313,N_4068);
or U5927 (N_5927,N_4936,N_2540);
nor U5928 (N_5928,N_3770,N_3646);
nor U5929 (N_5929,N_4418,N_4593);
and U5930 (N_5930,N_4339,N_3245);
and U5931 (N_5931,N_3253,N_3407);
xnor U5932 (N_5932,N_3077,N_4601);
or U5933 (N_5933,N_3829,N_4500);
nand U5934 (N_5934,N_2811,N_3290);
and U5935 (N_5935,N_4692,N_2680);
and U5936 (N_5936,N_4331,N_3052);
and U5937 (N_5937,N_4909,N_3536);
nor U5938 (N_5938,N_2849,N_3839);
nor U5939 (N_5939,N_3599,N_4525);
nor U5940 (N_5940,N_3043,N_4800);
nand U5941 (N_5941,N_2659,N_2743);
nand U5942 (N_5942,N_3371,N_4216);
nand U5943 (N_5943,N_4015,N_2600);
or U5944 (N_5944,N_3840,N_3717);
nand U5945 (N_5945,N_4432,N_3393);
nor U5946 (N_5946,N_4871,N_3589);
and U5947 (N_5947,N_4548,N_3973);
nand U5948 (N_5948,N_3477,N_3240);
and U5949 (N_5949,N_3705,N_3940);
nand U5950 (N_5950,N_4775,N_3896);
and U5951 (N_5951,N_4759,N_3846);
nor U5952 (N_5952,N_4027,N_3642);
or U5953 (N_5953,N_3381,N_3413);
and U5954 (N_5954,N_3499,N_4952);
or U5955 (N_5955,N_3990,N_3849);
or U5956 (N_5956,N_3633,N_4204);
nor U5957 (N_5957,N_4315,N_2756);
or U5958 (N_5958,N_4172,N_3445);
nor U5959 (N_5959,N_2801,N_4719);
or U5960 (N_5960,N_2613,N_4088);
nand U5961 (N_5961,N_3010,N_2514);
nor U5962 (N_5962,N_4063,N_3320);
or U5963 (N_5963,N_2507,N_3777);
nor U5964 (N_5964,N_3935,N_2776);
and U5965 (N_5965,N_2587,N_3446);
and U5966 (N_5966,N_2998,N_3861);
or U5967 (N_5967,N_3937,N_4687);
nand U5968 (N_5968,N_4300,N_4598);
xor U5969 (N_5969,N_4126,N_3474);
nor U5970 (N_5970,N_4365,N_3999);
and U5971 (N_5971,N_4217,N_4819);
and U5972 (N_5972,N_4554,N_4738);
and U5973 (N_5973,N_3163,N_2610);
xnor U5974 (N_5974,N_2609,N_2539);
nand U5975 (N_5975,N_3361,N_3063);
nor U5976 (N_5976,N_4880,N_2857);
nor U5977 (N_5977,N_3244,N_4939);
or U5978 (N_5978,N_4494,N_4162);
xor U5979 (N_5979,N_4084,N_3678);
or U5980 (N_5980,N_2525,N_4910);
nor U5981 (N_5981,N_2938,N_3838);
nor U5982 (N_5982,N_4142,N_4947);
and U5983 (N_5983,N_2859,N_2921);
nor U5984 (N_5984,N_4280,N_3207);
or U5985 (N_5985,N_4803,N_4655);
nor U5986 (N_5986,N_2721,N_2738);
and U5987 (N_5987,N_4201,N_4267);
or U5988 (N_5988,N_2876,N_3347);
and U5989 (N_5989,N_3691,N_4748);
and U5990 (N_5990,N_4452,N_4763);
and U5991 (N_5991,N_2590,N_4239);
nor U5992 (N_5992,N_3799,N_4620);
nand U5993 (N_5993,N_4282,N_3585);
nor U5994 (N_5994,N_4927,N_4227);
nor U5995 (N_5995,N_2520,N_3821);
or U5996 (N_5996,N_3057,N_4746);
xnor U5997 (N_5997,N_4526,N_4243);
and U5998 (N_5998,N_4834,N_4690);
nor U5999 (N_5999,N_4028,N_4824);
nor U6000 (N_6000,N_3349,N_4400);
or U6001 (N_6001,N_4195,N_2975);
nand U6002 (N_6002,N_4306,N_3293);
and U6003 (N_6003,N_4369,N_2821);
or U6004 (N_6004,N_2781,N_3857);
nor U6005 (N_6005,N_3879,N_4976);
nand U6006 (N_6006,N_4042,N_3909);
and U6007 (N_6007,N_4915,N_2606);
nor U6008 (N_6008,N_4238,N_3679);
or U6009 (N_6009,N_4136,N_3720);
nand U6010 (N_6010,N_2589,N_3042);
and U6011 (N_6011,N_4268,N_3094);
and U6012 (N_6012,N_3786,N_3824);
nor U6013 (N_6013,N_3091,N_2530);
or U6014 (N_6014,N_4213,N_4845);
nand U6015 (N_6015,N_3991,N_4057);
or U6016 (N_6016,N_3345,N_4991);
nor U6017 (N_6017,N_3428,N_4774);
nor U6018 (N_6018,N_3914,N_3529);
nand U6019 (N_6019,N_2677,N_4929);
or U6020 (N_6020,N_3471,N_2524);
or U6021 (N_6021,N_4954,N_4378);
nand U6022 (N_6022,N_3981,N_2722);
nand U6023 (N_6023,N_4971,N_4022);
nor U6024 (N_6024,N_3213,N_3618);
and U6025 (N_6025,N_4475,N_3335);
or U6026 (N_6026,N_4668,N_4013);
and U6027 (N_6027,N_4415,N_3704);
and U6028 (N_6028,N_4736,N_4051);
and U6029 (N_6029,N_3117,N_3110);
nor U6030 (N_6030,N_2847,N_4628);
nand U6031 (N_6031,N_4221,N_4040);
nor U6032 (N_6032,N_4097,N_2954);
and U6033 (N_6033,N_4573,N_2591);
xor U6034 (N_6034,N_3034,N_4528);
nand U6035 (N_6035,N_4674,N_3901);
and U6036 (N_6036,N_4729,N_4309);
nand U6037 (N_6037,N_3876,N_4383);
and U6038 (N_6038,N_4171,N_3182);
or U6039 (N_6039,N_4905,N_3278);
and U6040 (N_6040,N_2519,N_2845);
and U6041 (N_6041,N_3689,N_2535);
nor U6042 (N_6042,N_4979,N_3724);
nand U6043 (N_6043,N_4005,N_3362);
and U6044 (N_6044,N_4158,N_4011);
nand U6045 (N_6045,N_3779,N_3284);
nand U6046 (N_6046,N_4876,N_4513);
or U6047 (N_6047,N_4758,N_3353);
or U6048 (N_6048,N_4699,N_3832);
nand U6049 (N_6049,N_3097,N_4592);
and U6050 (N_6050,N_4184,N_4820);
xor U6051 (N_6051,N_3376,N_3934);
nand U6052 (N_6052,N_3941,N_3452);
nand U6053 (N_6053,N_3966,N_3774);
nor U6054 (N_6054,N_3767,N_3654);
nor U6055 (N_6055,N_3178,N_3115);
or U6056 (N_6056,N_2704,N_4919);
or U6057 (N_6057,N_4019,N_2855);
nor U6058 (N_6058,N_3420,N_3099);
nand U6059 (N_6059,N_3782,N_2596);
and U6060 (N_6060,N_3100,N_4384);
nand U6061 (N_6061,N_3564,N_3498);
nand U6062 (N_6062,N_4104,N_4430);
nand U6063 (N_6063,N_3613,N_2862);
xnor U6064 (N_6064,N_2794,N_3208);
and U6065 (N_6065,N_4041,N_4388);
nand U6066 (N_6066,N_3809,N_3204);
nand U6067 (N_6067,N_2810,N_3996);
nand U6068 (N_6068,N_3147,N_2626);
nand U6069 (N_6069,N_4145,N_2940);
and U6070 (N_6070,N_2882,N_4167);
nand U6071 (N_6071,N_3889,N_2713);
nor U6072 (N_6072,N_4169,N_4429);
nor U6073 (N_6073,N_3862,N_3619);
or U6074 (N_6074,N_3465,N_4153);
nand U6075 (N_6075,N_3732,N_4978);
nand U6076 (N_6076,N_3553,N_4425);
and U6077 (N_6077,N_3544,N_3516);
and U6078 (N_6078,N_2737,N_4906);
or U6079 (N_6079,N_3169,N_4766);
nor U6080 (N_6080,N_2513,N_3936);
or U6081 (N_6081,N_2634,N_3883);
or U6082 (N_6082,N_3541,N_4737);
and U6083 (N_6083,N_4994,N_4924);
nor U6084 (N_6084,N_3283,N_4853);
xor U6085 (N_6085,N_3060,N_4122);
nor U6086 (N_6086,N_4586,N_4867);
nor U6087 (N_6087,N_3847,N_4559);
and U6088 (N_6088,N_4303,N_3652);
nand U6089 (N_6089,N_3488,N_2717);
and U6090 (N_6090,N_4342,N_4977);
and U6091 (N_6091,N_3747,N_2726);
xor U6092 (N_6092,N_4188,N_3833);
or U6093 (N_6093,N_3932,N_3603);
and U6094 (N_6094,N_4370,N_4604);
and U6095 (N_6095,N_3693,N_3975);
nand U6096 (N_6096,N_4816,N_4964);
or U6097 (N_6097,N_4449,N_2771);
or U6098 (N_6098,N_3760,N_2860);
or U6099 (N_6099,N_4611,N_3495);
nor U6100 (N_6100,N_4297,N_2515);
nor U6101 (N_6101,N_3740,N_3602);
nand U6102 (N_6102,N_3156,N_2725);
nand U6103 (N_6103,N_3273,N_3272);
and U6104 (N_6104,N_3796,N_2720);
nand U6105 (N_6105,N_4193,N_4688);
or U6106 (N_6106,N_3248,N_4291);
and U6107 (N_6107,N_4590,N_4409);
nand U6108 (N_6108,N_3462,N_4796);
or U6109 (N_6109,N_3197,N_4740);
and U6110 (N_6110,N_2537,N_3120);
or U6111 (N_6111,N_4155,N_3093);
nor U6112 (N_6112,N_2655,N_4896);
nand U6113 (N_6113,N_4164,N_2837);
nand U6114 (N_6114,N_3480,N_2529);
or U6115 (N_6115,N_4891,N_4270);
nand U6116 (N_6116,N_4397,N_2924);
or U6117 (N_6117,N_4685,N_2654);
nor U6118 (N_6118,N_3232,N_2834);
nand U6119 (N_6119,N_2727,N_2945);
or U6120 (N_6120,N_4348,N_2769);
nand U6121 (N_6121,N_3956,N_4138);
or U6122 (N_6122,N_4596,N_3286);
and U6123 (N_6123,N_2712,N_4634);
nor U6124 (N_6124,N_4702,N_3252);
nor U6125 (N_6125,N_2552,N_3007);
nand U6126 (N_6126,N_3729,N_2987);
nand U6127 (N_6127,N_3408,N_4928);
nand U6128 (N_6128,N_3150,N_3308);
and U6129 (N_6129,N_2681,N_3171);
nor U6130 (N_6130,N_2557,N_3911);
nor U6131 (N_6131,N_3444,N_3997);
or U6132 (N_6132,N_4941,N_4886);
nand U6133 (N_6133,N_2867,N_3542);
or U6134 (N_6134,N_3929,N_4642);
nand U6135 (N_6135,N_4046,N_3507);
and U6136 (N_6136,N_4582,N_3372);
nand U6137 (N_6137,N_2642,N_4381);
xnor U6138 (N_6138,N_3493,N_3288);
nor U6139 (N_6139,N_3787,N_3869);
or U6140 (N_6140,N_4098,N_3396);
or U6141 (N_6141,N_3211,N_4744);
and U6142 (N_6142,N_3550,N_3549);
nand U6143 (N_6143,N_3118,N_3666);
nor U6144 (N_6144,N_4625,N_3086);
or U6145 (N_6145,N_4715,N_4438);
and U6146 (N_6146,N_4020,N_2901);
nor U6147 (N_6147,N_4103,N_3583);
or U6148 (N_6148,N_4408,N_3453);
or U6149 (N_6149,N_4895,N_4289);
nand U6150 (N_6150,N_3955,N_4566);
and U6151 (N_6151,N_3061,N_4485);
or U6152 (N_6152,N_2812,N_3203);
nand U6153 (N_6153,N_2733,N_4556);
or U6154 (N_6154,N_3295,N_4273);
or U6155 (N_6155,N_3317,N_3778);
nand U6156 (N_6156,N_4170,N_3157);
or U6157 (N_6157,N_4202,N_2931);
or U6158 (N_6158,N_3759,N_2686);
nand U6159 (N_6159,N_2930,N_3749);
or U6160 (N_6160,N_4077,N_3670);
and U6161 (N_6161,N_3402,N_4470);
nor U6162 (N_6162,N_4829,N_4337);
or U6163 (N_6163,N_2692,N_3326);
nand U6164 (N_6164,N_4394,N_4026);
or U6165 (N_6165,N_3835,N_2934);
nor U6166 (N_6166,N_2678,N_4679);
and U6167 (N_6167,N_3868,N_3201);
nand U6168 (N_6168,N_4355,N_2783);
or U6169 (N_6169,N_2502,N_3863);
and U6170 (N_6170,N_4364,N_3080);
or U6171 (N_6171,N_2974,N_3775);
and U6172 (N_6172,N_3447,N_4305);
nor U6173 (N_6173,N_4286,N_3904);
nor U6174 (N_6174,N_3612,N_2878);
and U6175 (N_6175,N_3944,N_3469);
and U6176 (N_6176,N_3867,N_2646);
and U6177 (N_6177,N_3877,N_4362);
and U6178 (N_6178,N_2928,N_4501);
or U6179 (N_6179,N_3363,N_3300);
nor U6180 (N_6180,N_2817,N_4453);
and U6181 (N_6181,N_3448,N_3703);
and U6182 (N_6182,N_3084,N_4165);
nor U6183 (N_6183,N_3131,N_4035);
nand U6184 (N_6184,N_3817,N_3572);
and U6185 (N_6185,N_3659,N_3409);
or U6186 (N_6186,N_4993,N_4728);
nand U6187 (N_6187,N_3866,N_4583);
xnor U6188 (N_6188,N_4945,N_3872);
or U6189 (N_6189,N_4776,N_3450);
nor U6190 (N_6190,N_4493,N_2822);
and U6191 (N_6191,N_3144,N_2767);
and U6192 (N_6192,N_3645,N_4761);
nor U6193 (N_6193,N_3980,N_4792);
nor U6194 (N_6194,N_2752,N_2802);
and U6195 (N_6195,N_3234,N_2868);
or U6196 (N_6196,N_4031,N_3279);
and U6197 (N_6197,N_3181,N_4675);
and U6198 (N_6198,N_2527,N_2800);
or U6199 (N_6199,N_2510,N_4472);
nor U6200 (N_6200,N_2560,N_4958);
and U6201 (N_6201,N_3519,N_4934);
or U6202 (N_6202,N_3771,N_4659);
or U6203 (N_6203,N_3661,N_2569);
xnor U6204 (N_6204,N_4527,N_4847);
nand U6205 (N_6205,N_2566,N_3313);
nor U6206 (N_6206,N_4597,N_3343);
and U6207 (N_6207,N_4382,N_3254);
nand U6208 (N_6208,N_2935,N_3170);
or U6209 (N_6209,N_4893,N_4482);
nand U6210 (N_6210,N_3601,N_3916);
nand U6211 (N_6211,N_4380,N_4568);
nor U6212 (N_6212,N_2816,N_3192);
and U6213 (N_6213,N_2842,N_4095);
nand U6214 (N_6214,N_3844,N_2647);
or U6215 (N_6215,N_4749,N_3993);
and U6216 (N_6216,N_3109,N_4010);
nand U6217 (N_6217,N_4448,N_4468);
and U6218 (N_6218,N_3382,N_3281);
or U6219 (N_6219,N_3304,N_3018);
nor U6220 (N_6220,N_2685,N_2755);
nor U6221 (N_6221,N_2872,N_3986);
and U6222 (N_6222,N_4466,N_4779);
or U6223 (N_6223,N_4645,N_3065);
nand U6224 (N_6224,N_4176,N_3953);
and U6225 (N_6225,N_2892,N_3752);
nand U6226 (N_6226,N_4617,N_3708);
nand U6227 (N_6227,N_3406,N_3132);
and U6228 (N_6228,N_2772,N_2958);
and U6229 (N_6229,N_3410,N_3346);
nand U6230 (N_6230,N_4571,N_3206);
or U6231 (N_6231,N_2910,N_2909);
nor U6232 (N_6232,N_4830,N_4319);
nor U6233 (N_6233,N_2740,N_3369);
nor U6234 (N_6234,N_4334,N_4879);
and U6235 (N_6235,N_4864,N_2555);
and U6236 (N_6236,N_2809,N_4814);
and U6237 (N_6237,N_3047,N_3852);
and U6238 (N_6238,N_4390,N_4182);
or U6239 (N_6239,N_4222,N_3478);
nor U6240 (N_6240,N_4283,N_3520);
nand U6241 (N_6241,N_3588,N_2894);
nand U6242 (N_6242,N_4080,N_4875);
nand U6243 (N_6243,N_4995,N_3492);
or U6244 (N_6244,N_4933,N_2703);
and U6245 (N_6245,N_4352,N_3930);
and U6246 (N_6246,N_4823,N_4643);
nor U6247 (N_6247,N_3772,N_3554);
or U6248 (N_6248,N_3658,N_4975);
nand U6249 (N_6249,N_4585,N_2698);
and U6250 (N_6250,N_3302,N_2501);
nor U6251 (N_6251,N_4923,N_4728);
nor U6252 (N_6252,N_3168,N_4625);
and U6253 (N_6253,N_3850,N_2700);
nor U6254 (N_6254,N_2667,N_4556);
or U6255 (N_6255,N_2628,N_2572);
nand U6256 (N_6256,N_3604,N_3483);
nor U6257 (N_6257,N_2833,N_2595);
or U6258 (N_6258,N_3970,N_3715);
nand U6259 (N_6259,N_4688,N_4903);
or U6260 (N_6260,N_4218,N_4474);
or U6261 (N_6261,N_4437,N_3583);
nor U6262 (N_6262,N_2680,N_3242);
xnor U6263 (N_6263,N_2709,N_4885);
nand U6264 (N_6264,N_4311,N_2980);
nand U6265 (N_6265,N_4030,N_4229);
nor U6266 (N_6266,N_3562,N_2854);
and U6267 (N_6267,N_2591,N_3115);
xnor U6268 (N_6268,N_4830,N_4895);
and U6269 (N_6269,N_2547,N_4496);
nor U6270 (N_6270,N_4544,N_4569);
or U6271 (N_6271,N_4887,N_4213);
nor U6272 (N_6272,N_4432,N_4454);
and U6273 (N_6273,N_3446,N_3099);
xor U6274 (N_6274,N_3602,N_4820);
nand U6275 (N_6275,N_3599,N_3817);
nor U6276 (N_6276,N_4017,N_2622);
and U6277 (N_6277,N_4897,N_4119);
nand U6278 (N_6278,N_4860,N_4164);
or U6279 (N_6279,N_3451,N_3827);
nand U6280 (N_6280,N_4393,N_2856);
nor U6281 (N_6281,N_4577,N_2636);
nor U6282 (N_6282,N_4698,N_3631);
and U6283 (N_6283,N_4379,N_4171);
or U6284 (N_6284,N_4438,N_3488);
or U6285 (N_6285,N_3772,N_4449);
and U6286 (N_6286,N_3721,N_4077);
or U6287 (N_6287,N_3377,N_3805);
and U6288 (N_6288,N_4652,N_2630);
nor U6289 (N_6289,N_3037,N_3014);
and U6290 (N_6290,N_2506,N_3162);
nor U6291 (N_6291,N_3615,N_2864);
and U6292 (N_6292,N_4076,N_3309);
xnor U6293 (N_6293,N_4850,N_3173);
nand U6294 (N_6294,N_2684,N_4968);
nand U6295 (N_6295,N_3659,N_4728);
nor U6296 (N_6296,N_3106,N_4098);
nor U6297 (N_6297,N_4493,N_4905);
and U6298 (N_6298,N_4683,N_2747);
or U6299 (N_6299,N_3647,N_3671);
and U6300 (N_6300,N_4937,N_4705);
and U6301 (N_6301,N_4974,N_4469);
and U6302 (N_6302,N_3540,N_2506);
xor U6303 (N_6303,N_3986,N_4594);
nor U6304 (N_6304,N_3273,N_3248);
nor U6305 (N_6305,N_3438,N_3454);
or U6306 (N_6306,N_4551,N_3822);
or U6307 (N_6307,N_4128,N_2789);
nand U6308 (N_6308,N_4458,N_3628);
or U6309 (N_6309,N_4051,N_4238);
nor U6310 (N_6310,N_4563,N_2957);
nor U6311 (N_6311,N_3830,N_3640);
nand U6312 (N_6312,N_2553,N_4432);
and U6313 (N_6313,N_4833,N_4753);
and U6314 (N_6314,N_4506,N_3087);
or U6315 (N_6315,N_3670,N_4911);
or U6316 (N_6316,N_2785,N_4317);
nor U6317 (N_6317,N_4183,N_3441);
nand U6318 (N_6318,N_4887,N_3764);
or U6319 (N_6319,N_2589,N_4868);
nor U6320 (N_6320,N_4026,N_4670);
nor U6321 (N_6321,N_4626,N_4881);
nand U6322 (N_6322,N_2563,N_3662);
or U6323 (N_6323,N_4080,N_2893);
nand U6324 (N_6324,N_4453,N_2757);
or U6325 (N_6325,N_2683,N_2678);
nor U6326 (N_6326,N_3442,N_2531);
or U6327 (N_6327,N_3701,N_3454);
nand U6328 (N_6328,N_4403,N_3816);
nor U6329 (N_6329,N_4048,N_2561);
or U6330 (N_6330,N_3615,N_3730);
or U6331 (N_6331,N_4265,N_4389);
nor U6332 (N_6332,N_3546,N_3381);
nand U6333 (N_6333,N_4009,N_2524);
nor U6334 (N_6334,N_4180,N_3608);
or U6335 (N_6335,N_4896,N_3885);
nand U6336 (N_6336,N_2832,N_4711);
and U6337 (N_6337,N_3954,N_3474);
nor U6338 (N_6338,N_3560,N_3755);
nor U6339 (N_6339,N_4840,N_4481);
nor U6340 (N_6340,N_3435,N_4145);
or U6341 (N_6341,N_4287,N_3313);
nor U6342 (N_6342,N_3046,N_4329);
or U6343 (N_6343,N_4323,N_4875);
xnor U6344 (N_6344,N_2837,N_4857);
or U6345 (N_6345,N_3637,N_3813);
and U6346 (N_6346,N_4223,N_2751);
nand U6347 (N_6347,N_2574,N_4825);
nand U6348 (N_6348,N_4584,N_2860);
or U6349 (N_6349,N_3102,N_4457);
xor U6350 (N_6350,N_4877,N_3262);
or U6351 (N_6351,N_4526,N_3956);
nand U6352 (N_6352,N_2545,N_4468);
or U6353 (N_6353,N_2730,N_2588);
or U6354 (N_6354,N_4187,N_3317);
nor U6355 (N_6355,N_4803,N_3601);
and U6356 (N_6356,N_3993,N_2983);
nand U6357 (N_6357,N_3763,N_2560);
nand U6358 (N_6358,N_4442,N_3849);
or U6359 (N_6359,N_3479,N_3469);
nand U6360 (N_6360,N_3471,N_4198);
or U6361 (N_6361,N_4233,N_3267);
or U6362 (N_6362,N_3025,N_4424);
or U6363 (N_6363,N_2933,N_3635);
and U6364 (N_6364,N_3641,N_4917);
and U6365 (N_6365,N_4651,N_3543);
and U6366 (N_6366,N_4050,N_4150);
nor U6367 (N_6367,N_4129,N_4134);
nand U6368 (N_6368,N_4063,N_3685);
nand U6369 (N_6369,N_2963,N_4634);
and U6370 (N_6370,N_3042,N_4904);
nor U6371 (N_6371,N_3432,N_3671);
nor U6372 (N_6372,N_3030,N_2522);
or U6373 (N_6373,N_4051,N_2562);
and U6374 (N_6374,N_3471,N_4461);
and U6375 (N_6375,N_4483,N_3464);
and U6376 (N_6376,N_3687,N_3316);
nor U6377 (N_6377,N_3844,N_2968);
nor U6378 (N_6378,N_3986,N_4614);
nand U6379 (N_6379,N_3217,N_3473);
nand U6380 (N_6380,N_2787,N_4676);
nor U6381 (N_6381,N_2641,N_3635);
or U6382 (N_6382,N_4440,N_3663);
or U6383 (N_6383,N_4163,N_3163);
or U6384 (N_6384,N_4220,N_2728);
nand U6385 (N_6385,N_3368,N_2569);
nor U6386 (N_6386,N_3556,N_3230);
and U6387 (N_6387,N_4892,N_4944);
or U6388 (N_6388,N_4611,N_2761);
and U6389 (N_6389,N_2591,N_4283);
nor U6390 (N_6390,N_4472,N_4705);
nand U6391 (N_6391,N_3579,N_3554);
and U6392 (N_6392,N_2501,N_4997);
and U6393 (N_6393,N_4054,N_3492);
nor U6394 (N_6394,N_4079,N_3396);
and U6395 (N_6395,N_4432,N_3173);
or U6396 (N_6396,N_4400,N_3737);
or U6397 (N_6397,N_2853,N_4639);
nor U6398 (N_6398,N_3194,N_4213);
nand U6399 (N_6399,N_4731,N_3392);
or U6400 (N_6400,N_4611,N_2589);
and U6401 (N_6401,N_3010,N_3911);
nor U6402 (N_6402,N_4684,N_2686);
or U6403 (N_6403,N_3555,N_2855);
or U6404 (N_6404,N_3206,N_2995);
and U6405 (N_6405,N_4085,N_3165);
or U6406 (N_6406,N_4561,N_3274);
xnor U6407 (N_6407,N_3825,N_3710);
nand U6408 (N_6408,N_4811,N_2567);
nor U6409 (N_6409,N_3019,N_3268);
nand U6410 (N_6410,N_2778,N_4353);
or U6411 (N_6411,N_4307,N_2886);
nor U6412 (N_6412,N_2937,N_2774);
nand U6413 (N_6413,N_2819,N_3397);
nor U6414 (N_6414,N_2895,N_4165);
nand U6415 (N_6415,N_3500,N_2639);
and U6416 (N_6416,N_2706,N_3384);
nor U6417 (N_6417,N_2858,N_3862);
xor U6418 (N_6418,N_3753,N_4002);
nor U6419 (N_6419,N_4398,N_2950);
xnor U6420 (N_6420,N_3851,N_4662);
xnor U6421 (N_6421,N_2830,N_4562);
and U6422 (N_6422,N_4972,N_4911);
or U6423 (N_6423,N_4313,N_2531);
xor U6424 (N_6424,N_4941,N_4284);
nand U6425 (N_6425,N_4118,N_2704);
nand U6426 (N_6426,N_3322,N_2596);
nor U6427 (N_6427,N_4187,N_3157);
and U6428 (N_6428,N_3930,N_4900);
and U6429 (N_6429,N_2717,N_3293);
nand U6430 (N_6430,N_3977,N_4029);
nand U6431 (N_6431,N_4313,N_3529);
nor U6432 (N_6432,N_3993,N_4998);
and U6433 (N_6433,N_2615,N_3157);
nand U6434 (N_6434,N_4932,N_3983);
nor U6435 (N_6435,N_4081,N_3423);
nand U6436 (N_6436,N_3721,N_3172);
and U6437 (N_6437,N_4988,N_4938);
nor U6438 (N_6438,N_3954,N_3208);
nor U6439 (N_6439,N_2870,N_3259);
or U6440 (N_6440,N_4734,N_2978);
nand U6441 (N_6441,N_3203,N_4645);
nand U6442 (N_6442,N_3077,N_3082);
nor U6443 (N_6443,N_4519,N_4749);
or U6444 (N_6444,N_3172,N_4207);
nand U6445 (N_6445,N_3391,N_3579);
or U6446 (N_6446,N_2738,N_3040);
and U6447 (N_6447,N_3602,N_4964);
xor U6448 (N_6448,N_2728,N_3401);
or U6449 (N_6449,N_4299,N_4426);
nor U6450 (N_6450,N_4302,N_2899);
nor U6451 (N_6451,N_3976,N_3778);
nor U6452 (N_6452,N_4920,N_3925);
and U6453 (N_6453,N_4288,N_3525);
nand U6454 (N_6454,N_3159,N_3295);
nor U6455 (N_6455,N_4141,N_4369);
nor U6456 (N_6456,N_4307,N_2960);
nand U6457 (N_6457,N_2966,N_4917);
or U6458 (N_6458,N_2939,N_4824);
nor U6459 (N_6459,N_3428,N_3018);
or U6460 (N_6460,N_3929,N_2749);
or U6461 (N_6461,N_2850,N_2960);
or U6462 (N_6462,N_4518,N_3102);
or U6463 (N_6463,N_3811,N_3651);
nand U6464 (N_6464,N_4805,N_3930);
nor U6465 (N_6465,N_3858,N_2976);
or U6466 (N_6466,N_4389,N_3768);
nand U6467 (N_6467,N_4884,N_4503);
nor U6468 (N_6468,N_2813,N_3437);
or U6469 (N_6469,N_3373,N_3690);
nand U6470 (N_6470,N_3836,N_3413);
nand U6471 (N_6471,N_4831,N_2943);
nor U6472 (N_6472,N_3154,N_3766);
and U6473 (N_6473,N_3762,N_2872);
nor U6474 (N_6474,N_4454,N_3279);
and U6475 (N_6475,N_3293,N_4021);
nor U6476 (N_6476,N_2609,N_4105);
nor U6477 (N_6477,N_3935,N_3864);
nor U6478 (N_6478,N_4393,N_3150);
or U6479 (N_6479,N_4386,N_3297);
or U6480 (N_6480,N_2650,N_3200);
nand U6481 (N_6481,N_4353,N_4077);
and U6482 (N_6482,N_4567,N_2956);
or U6483 (N_6483,N_4644,N_2991);
nor U6484 (N_6484,N_4487,N_3731);
nor U6485 (N_6485,N_2680,N_3556);
and U6486 (N_6486,N_4972,N_2656);
or U6487 (N_6487,N_2976,N_3670);
nand U6488 (N_6488,N_4671,N_3745);
nor U6489 (N_6489,N_3512,N_3184);
nand U6490 (N_6490,N_2725,N_2873);
and U6491 (N_6491,N_4301,N_4025);
or U6492 (N_6492,N_3911,N_4674);
and U6493 (N_6493,N_4454,N_3610);
and U6494 (N_6494,N_2673,N_4511);
or U6495 (N_6495,N_2910,N_4233);
nand U6496 (N_6496,N_3203,N_3047);
xor U6497 (N_6497,N_4694,N_4156);
nor U6498 (N_6498,N_2641,N_4572);
nand U6499 (N_6499,N_2950,N_3191);
or U6500 (N_6500,N_3839,N_3360);
and U6501 (N_6501,N_3092,N_3880);
nand U6502 (N_6502,N_3227,N_4039);
nand U6503 (N_6503,N_4614,N_4891);
nand U6504 (N_6504,N_4855,N_4293);
or U6505 (N_6505,N_4474,N_4720);
nand U6506 (N_6506,N_4131,N_4959);
and U6507 (N_6507,N_2775,N_2801);
or U6508 (N_6508,N_2770,N_3308);
or U6509 (N_6509,N_4676,N_3733);
nor U6510 (N_6510,N_3826,N_4129);
xnor U6511 (N_6511,N_2586,N_4551);
or U6512 (N_6512,N_3616,N_3914);
nand U6513 (N_6513,N_4274,N_4896);
and U6514 (N_6514,N_3450,N_4894);
and U6515 (N_6515,N_3767,N_4623);
and U6516 (N_6516,N_2672,N_2648);
nand U6517 (N_6517,N_4229,N_4852);
and U6518 (N_6518,N_3988,N_3007);
nor U6519 (N_6519,N_4824,N_2521);
and U6520 (N_6520,N_3040,N_3674);
and U6521 (N_6521,N_2776,N_4788);
nand U6522 (N_6522,N_2853,N_3829);
nand U6523 (N_6523,N_4413,N_3226);
and U6524 (N_6524,N_4876,N_4704);
nand U6525 (N_6525,N_3815,N_4710);
nand U6526 (N_6526,N_3617,N_3592);
nand U6527 (N_6527,N_4500,N_2689);
nand U6528 (N_6528,N_3932,N_4126);
nor U6529 (N_6529,N_4654,N_4294);
nor U6530 (N_6530,N_3808,N_2810);
nand U6531 (N_6531,N_3947,N_3439);
nor U6532 (N_6532,N_3526,N_2505);
nor U6533 (N_6533,N_3209,N_3918);
or U6534 (N_6534,N_3366,N_4651);
or U6535 (N_6535,N_2687,N_4103);
nand U6536 (N_6536,N_3521,N_4561);
nand U6537 (N_6537,N_4638,N_3651);
or U6538 (N_6538,N_4415,N_2587);
nand U6539 (N_6539,N_3887,N_3895);
or U6540 (N_6540,N_3672,N_4643);
or U6541 (N_6541,N_3712,N_4021);
nand U6542 (N_6542,N_2873,N_4538);
and U6543 (N_6543,N_4590,N_4027);
nand U6544 (N_6544,N_3881,N_3936);
nor U6545 (N_6545,N_2768,N_4856);
and U6546 (N_6546,N_4032,N_3792);
and U6547 (N_6547,N_4763,N_3221);
nor U6548 (N_6548,N_4117,N_4150);
or U6549 (N_6549,N_3839,N_4305);
and U6550 (N_6550,N_4498,N_4853);
nand U6551 (N_6551,N_4387,N_2892);
or U6552 (N_6552,N_3331,N_4430);
xor U6553 (N_6553,N_2954,N_3103);
or U6554 (N_6554,N_4539,N_3663);
and U6555 (N_6555,N_2905,N_4305);
and U6556 (N_6556,N_4867,N_3088);
or U6557 (N_6557,N_4151,N_3385);
and U6558 (N_6558,N_4049,N_3037);
nor U6559 (N_6559,N_3581,N_4523);
nand U6560 (N_6560,N_4753,N_2642);
and U6561 (N_6561,N_3425,N_2585);
or U6562 (N_6562,N_3904,N_3392);
xor U6563 (N_6563,N_4659,N_2517);
or U6564 (N_6564,N_4846,N_3041);
or U6565 (N_6565,N_3479,N_3277);
nand U6566 (N_6566,N_4264,N_4289);
xor U6567 (N_6567,N_3204,N_2659);
or U6568 (N_6568,N_2765,N_3591);
or U6569 (N_6569,N_4079,N_2859);
and U6570 (N_6570,N_3859,N_3651);
or U6571 (N_6571,N_2559,N_3481);
or U6572 (N_6572,N_2572,N_4725);
or U6573 (N_6573,N_3201,N_3458);
and U6574 (N_6574,N_3532,N_3134);
or U6575 (N_6575,N_3090,N_4509);
or U6576 (N_6576,N_3524,N_4187);
and U6577 (N_6577,N_3602,N_3381);
nor U6578 (N_6578,N_3496,N_3143);
nand U6579 (N_6579,N_4339,N_2691);
or U6580 (N_6580,N_3006,N_4299);
and U6581 (N_6581,N_3533,N_4579);
nand U6582 (N_6582,N_4723,N_3865);
or U6583 (N_6583,N_4228,N_2614);
or U6584 (N_6584,N_4401,N_3289);
nand U6585 (N_6585,N_3461,N_4103);
nand U6586 (N_6586,N_4042,N_4770);
nand U6587 (N_6587,N_2763,N_2830);
and U6588 (N_6588,N_3144,N_2614);
and U6589 (N_6589,N_3501,N_4657);
nor U6590 (N_6590,N_3561,N_3821);
nor U6591 (N_6591,N_2724,N_4228);
xor U6592 (N_6592,N_3333,N_3055);
or U6593 (N_6593,N_4876,N_4690);
or U6594 (N_6594,N_3906,N_4260);
and U6595 (N_6595,N_4244,N_4869);
nor U6596 (N_6596,N_4720,N_4789);
nor U6597 (N_6597,N_3499,N_2687);
or U6598 (N_6598,N_2977,N_3957);
nor U6599 (N_6599,N_4359,N_2902);
xor U6600 (N_6600,N_4435,N_3665);
and U6601 (N_6601,N_3923,N_2694);
nand U6602 (N_6602,N_2931,N_3448);
and U6603 (N_6603,N_3294,N_4179);
nand U6604 (N_6604,N_3964,N_3773);
and U6605 (N_6605,N_2982,N_4963);
and U6606 (N_6606,N_4765,N_3802);
and U6607 (N_6607,N_2667,N_4368);
or U6608 (N_6608,N_3892,N_4413);
nor U6609 (N_6609,N_3497,N_3606);
or U6610 (N_6610,N_4021,N_3733);
nor U6611 (N_6611,N_3824,N_3328);
nor U6612 (N_6612,N_3998,N_4485);
or U6613 (N_6613,N_3369,N_3660);
or U6614 (N_6614,N_4659,N_4294);
and U6615 (N_6615,N_3453,N_2609);
nor U6616 (N_6616,N_3060,N_3019);
xor U6617 (N_6617,N_2865,N_3834);
or U6618 (N_6618,N_3763,N_4624);
nand U6619 (N_6619,N_2542,N_4613);
nand U6620 (N_6620,N_4119,N_3656);
nand U6621 (N_6621,N_3669,N_4671);
or U6622 (N_6622,N_3054,N_4276);
nand U6623 (N_6623,N_2641,N_4651);
or U6624 (N_6624,N_4811,N_4458);
nor U6625 (N_6625,N_2897,N_2849);
and U6626 (N_6626,N_3183,N_4639);
xor U6627 (N_6627,N_3475,N_3631);
nand U6628 (N_6628,N_4206,N_4990);
nor U6629 (N_6629,N_4468,N_4944);
nor U6630 (N_6630,N_4155,N_3528);
and U6631 (N_6631,N_4766,N_3136);
and U6632 (N_6632,N_3822,N_3306);
nor U6633 (N_6633,N_4153,N_2698);
nor U6634 (N_6634,N_2994,N_4419);
and U6635 (N_6635,N_4354,N_3981);
nor U6636 (N_6636,N_4193,N_3875);
or U6637 (N_6637,N_4406,N_2808);
nor U6638 (N_6638,N_3315,N_2699);
or U6639 (N_6639,N_4816,N_4464);
nand U6640 (N_6640,N_2948,N_3238);
and U6641 (N_6641,N_4850,N_3233);
nor U6642 (N_6642,N_3661,N_4607);
nand U6643 (N_6643,N_4368,N_3590);
or U6644 (N_6644,N_3108,N_4932);
nand U6645 (N_6645,N_2736,N_4323);
nand U6646 (N_6646,N_4047,N_2728);
and U6647 (N_6647,N_3474,N_3815);
nand U6648 (N_6648,N_3211,N_4555);
nand U6649 (N_6649,N_3447,N_2844);
nor U6650 (N_6650,N_4375,N_4290);
and U6651 (N_6651,N_3482,N_3833);
nor U6652 (N_6652,N_4806,N_4655);
nand U6653 (N_6653,N_4206,N_4309);
and U6654 (N_6654,N_4005,N_4099);
nand U6655 (N_6655,N_4621,N_4668);
xnor U6656 (N_6656,N_3581,N_3099);
nor U6657 (N_6657,N_3395,N_3419);
nor U6658 (N_6658,N_3638,N_3202);
or U6659 (N_6659,N_3628,N_2952);
nand U6660 (N_6660,N_4789,N_4748);
or U6661 (N_6661,N_2739,N_2569);
nor U6662 (N_6662,N_4993,N_4147);
or U6663 (N_6663,N_4588,N_3787);
nor U6664 (N_6664,N_4008,N_2829);
or U6665 (N_6665,N_2651,N_3095);
nor U6666 (N_6666,N_3426,N_4426);
and U6667 (N_6667,N_2624,N_4915);
or U6668 (N_6668,N_3997,N_2541);
nor U6669 (N_6669,N_3238,N_3885);
nand U6670 (N_6670,N_2799,N_2873);
and U6671 (N_6671,N_3388,N_4784);
nor U6672 (N_6672,N_2705,N_4292);
nor U6673 (N_6673,N_3847,N_3240);
or U6674 (N_6674,N_3736,N_4048);
and U6675 (N_6675,N_2860,N_4034);
nor U6676 (N_6676,N_3315,N_4341);
and U6677 (N_6677,N_4130,N_4626);
nor U6678 (N_6678,N_3699,N_4855);
or U6679 (N_6679,N_2995,N_4730);
nand U6680 (N_6680,N_4696,N_4232);
nand U6681 (N_6681,N_2583,N_4792);
nand U6682 (N_6682,N_2624,N_3542);
nand U6683 (N_6683,N_4477,N_4657);
or U6684 (N_6684,N_3705,N_3359);
nand U6685 (N_6685,N_3850,N_4127);
nand U6686 (N_6686,N_2624,N_2891);
nand U6687 (N_6687,N_4130,N_2560);
or U6688 (N_6688,N_4881,N_4914);
and U6689 (N_6689,N_4216,N_2627);
or U6690 (N_6690,N_3996,N_4121);
nand U6691 (N_6691,N_3074,N_4226);
nor U6692 (N_6692,N_3006,N_3463);
nor U6693 (N_6693,N_4352,N_3001);
and U6694 (N_6694,N_3049,N_4139);
and U6695 (N_6695,N_4063,N_2688);
and U6696 (N_6696,N_2518,N_4880);
or U6697 (N_6697,N_4520,N_3266);
nor U6698 (N_6698,N_2711,N_3482);
nand U6699 (N_6699,N_3765,N_3714);
or U6700 (N_6700,N_4111,N_3689);
and U6701 (N_6701,N_4610,N_4407);
nand U6702 (N_6702,N_3717,N_3405);
nor U6703 (N_6703,N_2984,N_2911);
nand U6704 (N_6704,N_4678,N_4223);
or U6705 (N_6705,N_4328,N_3308);
nand U6706 (N_6706,N_3776,N_2577);
xor U6707 (N_6707,N_4203,N_4310);
or U6708 (N_6708,N_3048,N_3744);
or U6709 (N_6709,N_2524,N_4880);
nor U6710 (N_6710,N_4111,N_2867);
or U6711 (N_6711,N_3783,N_4025);
nor U6712 (N_6712,N_3692,N_4153);
nand U6713 (N_6713,N_4582,N_4186);
nor U6714 (N_6714,N_3831,N_4578);
nor U6715 (N_6715,N_4663,N_4598);
and U6716 (N_6716,N_4936,N_2667);
or U6717 (N_6717,N_3592,N_3164);
xnor U6718 (N_6718,N_4595,N_2882);
nor U6719 (N_6719,N_4056,N_2833);
and U6720 (N_6720,N_2833,N_4186);
or U6721 (N_6721,N_4510,N_4795);
xor U6722 (N_6722,N_4920,N_3832);
or U6723 (N_6723,N_4627,N_4060);
nand U6724 (N_6724,N_3333,N_3876);
nor U6725 (N_6725,N_3660,N_3405);
and U6726 (N_6726,N_3261,N_3140);
or U6727 (N_6727,N_3195,N_4046);
nand U6728 (N_6728,N_3079,N_4419);
nor U6729 (N_6729,N_3265,N_3172);
and U6730 (N_6730,N_3513,N_3506);
nor U6731 (N_6731,N_2735,N_4978);
or U6732 (N_6732,N_3555,N_3010);
nand U6733 (N_6733,N_3783,N_4467);
and U6734 (N_6734,N_4088,N_4202);
and U6735 (N_6735,N_4050,N_2989);
and U6736 (N_6736,N_4721,N_3419);
nand U6737 (N_6737,N_3467,N_3473);
or U6738 (N_6738,N_2644,N_4676);
and U6739 (N_6739,N_4181,N_2527);
xnor U6740 (N_6740,N_3769,N_4645);
nor U6741 (N_6741,N_4515,N_4350);
nor U6742 (N_6742,N_3915,N_3545);
nor U6743 (N_6743,N_4393,N_2948);
or U6744 (N_6744,N_4612,N_3157);
nand U6745 (N_6745,N_4317,N_3911);
and U6746 (N_6746,N_4795,N_4146);
and U6747 (N_6747,N_3347,N_2687);
nor U6748 (N_6748,N_4132,N_4261);
and U6749 (N_6749,N_3036,N_4174);
and U6750 (N_6750,N_2849,N_4635);
and U6751 (N_6751,N_3446,N_4578);
and U6752 (N_6752,N_4639,N_4651);
and U6753 (N_6753,N_4794,N_2928);
or U6754 (N_6754,N_3970,N_2643);
and U6755 (N_6755,N_4984,N_3473);
nand U6756 (N_6756,N_3647,N_3663);
nand U6757 (N_6757,N_3283,N_2684);
nor U6758 (N_6758,N_4416,N_3163);
or U6759 (N_6759,N_4288,N_4785);
or U6760 (N_6760,N_3207,N_4094);
and U6761 (N_6761,N_4678,N_4702);
and U6762 (N_6762,N_3567,N_2500);
nand U6763 (N_6763,N_3406,N_2639);
and U6764 (N_6764,N_4690,N_3741);
nor U6765 (N_6765,N_2944,N_4308);
or U6766 (N_6766,N_4192,N_2543);
and U6767 (N_6767,N_2795,N_4911);
or U6768 (N_6768,N_4444,N_4339);
or U6769 (N_6769,N_3646,N_3299);
and U6770 (N_6770,N_4214,N_4492);
nand U6771 (N_6771,N_3816,N_2794);
nor U6772 (N_6772,N_4686,N_3455);
nand U6773 (N_6773,N_4177,N_2956);
nor U6774 (N_6774,N_3860,N_3734);
nand U6775 (N_6775,N_3656,N_4141);
nor U6776 (N_6776,N_4947,N_4135);
or U6777 (N_6777,N_4149,N_3153);
and U6778 (N_6778,N_2983,N_3166);
and U6779 (N_6779,N_2855,N_2592);
and U6780 (N_6780,N_4262,N_3581);
nor U6781 (N_6781,N_3310,N_3216);
nand U6782 (N_6782,N_4100,N_4130);
and U6783 (N_6783,N_3361,N_3714);
nand U6784 (N_6784,N_2986,N_4753);
or U6785 (N_6785,N_2865,N_3426);
and U6786 (N_6786,N_4743,N_3307);
and U6787 (N_6787,N_3927,N_2999);
or U6788 (N_6788,N_4668,N_3599);
nand U6789 (N_6789,N_3852,N_3257);
and U6790 (N_6790,N_2555,N_3008);
and U6791 (N_6791,N_3932,N_3180);
nor U6792 (N_6792,N_4265,N_2662);
and U6793 (N_6793,N_4458,N_4385);
nor U6794 (N_6794,N_3735,N_2544);
or U6795 (N_6795,N_4413,N_2699);
or U6796 (N_6796,N_4619,N_2565);
nand U6797 (N_6797,N_4523,N_3752);
and U6798 (N_6798,N_3246,N_4019);
nor U6799 (N_6799,N_4184,N_2675);
and U6800 (N_6800,N_2847,N_3972);
or U6801 (N_6801,N_3664,N_4262);
and U6802 (N_6802,N_3435,N_3894);
and U6803 (N_6803,N_3953,N_2602);
nor U6804 (N_6804,N_3173,N_4329);
and U6805 (N_6805,N_4288,N_4421);
nand U6806 (N_6806,N_3343,N_4048);
nand U6807 (N_6807,N_3803,N_3084);
or U6808 (N_6808,N_4804,N_3067);
nor U6809 (N_6809,N_3359,N_3297);
nor U6810 (N_6810,N_4202,N_4336);
or U6811 (N_6811,N_4206,N_2660);
nor U6812 (N_6812,N_3388,N_2592);
and U6813 (N_6813,N_3679,N_2655);
and U6814 (N_6814,N_4502,N_2898);
and U6815 (N_6815,N_2787,N_3936);
xnor U6816 (N_6816,N_4792,N_3589);
and U6817 (N_6817,N_4051,N_3577);
nand U6818 (N_6818,N_4766,N_4294);
nand U6819 (N_6819,N_2750,N_3581);
nor U6820 (N_6820,N_4745,N_3138);
nand U6821 (N_6821,N_3667,N_2539);
or U6822 (N_6822,N_4198,N_3031);
xor U6823 (N_6823,N_2923,N_3362);
nor U6824 (N_6824,N_2793,N_3368);
nor U6825 (N_6825,N_3621,N_3516);
nor U6826 (N_6826,N_3689,N_3344);
nor U6827 (N_6827,N_2988,N_4096);
or U6828 (N_6828,N_4268,N_4123);
nor U6829 (N_6829,N_3078,N_2655);
nor U6830 (N_6830,N_3393,N_2653);
nand U6831 (N_6831,N_3116,N_3445);
or U6832 (N_6832,N_3784,N_2849);
nor U6833 (N_6833,N_3607,N_4399);
nand U6834 (N_6834,N_2718,N_4833);
nor U6835 (N_6835,N_3387,N_3757);
or U6836 (N_6836,N_2757,N_2808);
nand U6837 (N_6837,N_2960,N_4633);
nand U6838 (N_6838,N_2572,N_3683);
nand U6839 (N_6839,N_3408,N_4559);
or U6840 (N_6840,N_2935,N_4042);
or U6841 (N_6841,N_2703,N_3931);
nand U6842 (N_6842,N_2559,N_3172);
and U6843 (N_6843,N_4686,N_2848);
and U6844 (N_6844,N_3429,N_2888);
or U6845 (N_6845,N_2959,N_3777);
and U6846 (N_6846,N_4812,N_4539);
or U6847 (N_6847,N_3819,N_4992);
and U6848 (N_6848,N_3980,N_2578);
or U6849 (N_6849,N_4192,N_3236);
nor U6850 (N_6850,N_3708,N_3485);
nor U6851 (N_6851,N_4189,N_4792);
or U6852 (N_6852,N_3766,N_3786);
nand U6853 (N_6853,N_3990,N_3601);
nor U6854 (N_6854,N_3914,N_3199);
nand U6855 (N_6855,N_4596,N_2508);
xor U6856 (N_6856,N_4191,N_3907);
nand U6857 (N_6857,N_2930,N_3757);
xor U6858 (N_6858,N_4850,N_3262);
and U6859 (N_6859,N_4142,N_3257);
xor U6860 (N_6860,N_4252,N_3950);
or U6861 (N_6861,N_4606,N_2955);
nor U6862 (N_6862,N_3223,N_2973);
nor U6863 (N_6863,N_3962,N_3908);
or U6864 (N_6864,N_2785,N_4933);
nand U6865 (N_6865,N_2507,N_4783);
nor U6866 (N_6866,N_3858,N_4743);
or U6867 (N_6867,N_2587,N_3161);
xnor U6868 (N_6868,N_2757,N_3292);
and U6869 (N_6869,N_4725,N_4730);
nand U6870 (N_6870,N_2572,N_3419);
nor U6871 (N_6871,N_3006,N_3103);
and U6872 (N_6872,N_4461,N_3429);
nand U6873 (N_6873,N_4840,N_3846);
and U6874 (N_6874,N_3263,N_2557);
or U6875 (N_6875,N_3649,N_2598);
nor U6876 (N_6876,N_3268,N_4343);
and U6877 (N_6877,N_4926,N_4925);
nor U6878 (N_6878,N_3065,N_4846);
or U6879 (N_6879,N_3160,N_4400);
and U6880 (N_6880,N_2960,N_3901);
or U6881 (N_6881,N_4882,N_4529);
and U6882 (N_6882,N_3868,N_4975);
nand U6883 (N_6883,N_4168,N_4625);
or U6884 (N_6884,N_4615,N_3895);
and U6885 (N_6885,N_4351,N_4065);
or U6886 (N_6886,N_3973,N_2588);
nor U6887 (N_6887,N_3079,N_4018);
nor U6888 (N_6888,N_3332,N_4407);
and U6889 (N_6889,N_4678,N_3254);
or U6890 (N_6890,N_2955,N_4239);
and U6891 (N_6891,N_4080,N_3414);
and U6892 (N_6892,N_4303,N_3604);
and U6893 (N_6893,N_4052,N_3271);
nor U6894 (N_6894,N_2658,N_3964);
nand U6895 (N_6895,N_3584,N_4973);
nor U6896 (N_6896,N_4654,N_4992);
and U6897 (N_6897,N_4413,N_4055);
nor U6898 (N_6898,N_4007,N_2598);
nand U6899 (N_6899,N_2605,N_3450);
nand U6900 (N_6900,N_4739,N_4278);
nor U6901 (N_6901,N_3380,N_3019);
nor U6902 (N_6902,N_2782,N_3902);
or U6903 (N_6903,N_2893,N_4550);
or U6904 (N_6904,N_4556,N_4706);
nor U6905 (N_6905,N_4393,N_3689);
nand U6906 (N_6906,N_3687,N_3372);
and U6907 (N_6907,N_4508,N_3207);
or U6908 (N_6908,N_3081,N_3143);
or U6909 (N_6909,N_3079,N_4730);
xor U6910 (N_6910,N_4592,N_3801);
nand U6911 (N_6911,N_4722,N_3641);
nand U6912 (N_6912,N_4798,N_2683);
and U6913 (N_6913,N_4846,N_3827);
nand U6914 (N_6914,N_3727,N_4600);
nand U6915 (N_6915,N_3587,N_3691);
nor U6916 (N_6916,N_4818,N_4735);
nor U6917 (N_6917,N_4575,N_3820);
and U6918 (N_6918,N_2986,N_3359);
nor U6919 (N_6919,N_2651,N_2923);
and U6920 (N_6920,N_4539,N_4644);
nand U6921 (N_6921,N_3124,N_3272);
nor U6922 (N_6922,N_3066,N_2977);
nor U6923 (N_6923,N_4084,N_4099);
or U6924 (N_6924,N_3135,N_4392);
nor U6925 (N_6925,N_3358,N_4908);
and U6926 (N_6926,N_4495,N_3322);
and U6927 (N_6927,N_3670,N_3897);
nor U6928 (N_6928,N_4146,N_2881);
nand U6929 (N_6929,N_4449,N_3537);
and U6930 (N_6930,N_4978,N_2531);
and U6931 (N_6931,N_3110,N_4044);
nor U6932 (N_6932,N_3841,N_3091);
nand U6933 (N_6933,N_3740,N_4670);
xor U6934 (N_6934,N_4097,N_3659);
or U6935 (N_6935,N_3440,N_2738);
nand U6936 (N_6936,N_2896,N_3790);
nand U6937 (N_6937,N_4131,N_4730);
or U6938 (N_6938,N_2502,N_2978);
nand U6939 (N_6939,N_3284,N_3188);
nand U6940 (N_6940,N_4510,N_4785);
nand U6941 (N_6941,N_2838,N_3129);
and U6942 (N_6942,N_3652,N_2790);
and U6943 (N_6943,N_3134,N_2526);
nor U6944 (N_6944,N_2509,N_3124);
nand U6945 (N_6945,N_4163,N_3483);
or U6946 (N_6946,N_4637,N_3923);
nor U6947 (N_6947,N_2968,N_4028);
or U6948 (N_6948,N_4760,N_3248);
nor U6949 (N_6949,N_3829,N_2952);
or U6950 (N_6950,N_2616,N_4882);
and U6951 (N_6951,N_3983,N_3991);
and U6952 (N_6952,N_4027,N_3099);
nor U6953 (N_6953,N_3897,N_4165);
and U6954 (N_6954,N_3605,N_2704);
nor U6955 (N_6955,N_3942,N_4927);
nor U6956 (N_6956,N_2702,N_4668);
and U6957 (N_6957,N_3531,N_3932);
and U6958 (N_6958,N_3715,N_4201);
nand U6959 (N_6959,N_4489,N_2673);
and U6960 (N_6960,N_3700,N_4974);
nor U6961 (N_6961,N_3548,N_2604);
nand U6962 (N_6962,N_3988,N_3067);
or U6963 (N_6963,N_4850,N_3591);
nor U6964 (N_6964,N_2578,N_3341);
or U6965 (N_6965,N_3271,N_3999);
nor U6966 (N_6966,N_4040,N_4806);
nand U6967 (N_6967,N_4810,N_3237);
nor U6968 (N_6968,N_3652,N_3329);
nand U6969 (N_6969,N_4489,N_4572);
nor U6970 (N_6970,N_4687,N_2536);
or U6971 (N_6971,N_4691,N_4530);
nor U6972 (N_6972,N_2738,N_2768);
nand U6973 (N_6973,N_4452,N_3399);
nor U6974 (N_6974,N_3886,N_2858);
or U6975 (N_6975,N_3247,N_3382);
and U6976 (N_6976,N_4512,N_2873);
or U6977 (N_6977,N_2811,N_3598);
nand U6978 (N_6978,N_4144,N_4165);
or U6979 (N_6979,N_2731,N_3306);
or U6980 (N_6980,N_4349,N_3685);
nand U6981 (N_6981,N_3665,N_4128);
nor U6982 (N_6982,N_4078,N_4247);
or U6983 (N_6983,N_2851,N_4454);
and U6984 (N_6984,N_2587,N_3910);
nand U6985 (N_6985,N_3292,N_4197);
or U6986 (N_6986,N_3540,N_3225);
and U6987 (N_6987,N_4124,N_3682);
or U6988 (N_6988,N_4918,N_4267);
nand U6989 (N_6989,N_3189,N_4844);
xor U6990 (N_6990,N_4593,N_3035);
xor U6991 (N_6991,N_3890,N_4501);
nand U6992 (N_6992,N_4710,N_4080);
and U6993 (N_6993,N_4761,N_4048);
nor U6994 (N_6994,N_3988,N_4750);
or U6995 (N_6995,N_2985,N_4822);
nand U6996 (N_6996,N_2784,N_3760);
nor U6997 (N_6997,N_3456,N_4268);
nand U6998 (N_6998,N_4280,N_3534);
nand U6999 (N_6999,N_2753,N_3706);
nor U7000 (N_7000,N_3439,N_3143);
nor U7001 (N_7001,N_3323,N_4193);
and U7002 (N_7002,N_4831,N_3632);
or U7003 (N_7003,N_3251,N_4132);
and U7004 (N_7004,N_4900,N_4099);
nand U7005 (N_7005,N_3181,N_3194);
nor U7006 (N_7006,N_3146,N_2505);
and U7007 (N_7007,N_4262,N_4911);
nor U7008 (N_7008,N_3303,N_3428);
nand U7009 (N_7009,N_3627,N_4928);
nand U7010 (N_7010,N_2609,N_3511);
or U7011 (N_7011,N_3105,N_4759);
and U7012 (N_7012,N_2971,N_2532);
nand U7013 (N_7013,N_4514,N_4234);
and U7014 (N_7014,N_2844,N_3622);
or U7015 (N_7015,N_3920,N_4925);
nor U7016 (N_7016,N_4716,N_4400);
nand U7017 (N_7017,N_3587,N_3586);
or U7018 (N_7018,N_4055,N_2540);
and U7019 (N_7019,N_2705,N_4988);
xor U7020 (N_7020,N_4894,N_4345);
and U7021 (N_7021,N_3328,N_3232);
and U7022 (N_7022,N_2792,N_4338);
nor U7023 (N_7023,N_3601,N_2974);
nand U7024 (N_7024,N_2524,N_3110);
and U7025 (N_7025,N_3664,N_4099);
nand U7026 (N_7026,N_2542,N_3025);
nor U7027 (N_7027,N_4869,N_3993);
nor U7028 (N_7028,N_3919,N_4738);
nor U7029 (N_7029,N_3110,N_4556);
and U7030 (N_7030,N_2645,N_2994);
and U7031 (N_7031,N_4569,N_3135);
and U7032 (N_7032,N_4551,N_4579);
and U7033 (N_7033,N_4078,N_3596);
or U7034 (N_7034,N_4989,N_4461);
and U7035 (N_7035,N_4105,N_3648);
nand U7036 (N_7036,N_3644,N_4609);
or U7037 (N_7037,N_4331,N_3445);
and U7038 (N_7038,N_3026,N_3235);
and U7039 (N_7039,N_4436,N_4999);
nand U7040 (N_7040,N_2829,N_4933);
xnor U7041 (N_7041,N_4056,N_3214);
or U7042 (N_7042,N_2682,N_3960);
nor U7043 (N_7043,N_3925,N_4368);
xor U7044 (N_7044,N_4840,N_4005);
and U7045 (N_7045,N_3888,N_4058);
xnor U7046 (N_7046,N_4146,N_4525);
and U7047 (N_7047,N_3826,N_4363);
nor U7048 (N_7048,N_3888,N_3167);
or U7049 (N_7049,N_4070,N_4864);
and U7050 (N_7050,N_3313,N_4706);
or U7051 (N_7051,N_2733,N_3898);
and U7052 (N_7052,N_4623,N_4750);
nand U7053 (N_7053,N_4825,N_3728);
nand U7054 (N_7054,N_4552,N_3811);
nand U7055 (N_7055,N_4126,N_2967);
nand U7056 (N_7056,N_3879,N_3271);
nand U7057 (N_7057,N_4555,N_3943);
and U7058 (N_7058,N_4693,N_3566);
nor U7059 (N_7059,N_4557,N_3820);
or U7060 (N_7060,N_4095,N_4716);
nand U7061 (N_7061,N_3280,N_4792);
nor U7062 (N_7062,N_3399,N_3402);
and U7063 (N_7063,N_3441,N_4635);
nor U7064 (N_7064,N_4575,N_4231);
nor U7065 (N_7065,N_4866,N_2862);
nand U7066 (N_7066,N_2583,N_4320);
and U7067 (N_7067,N_3703,N_2559);
and U7068 (N_7068,N_4404,N_3300);
nand U7069 (N_7069,N_4471,N_3289);
or U7070 (N_7070,N_4661,N_4374);
and U7071 (N_7071,N_4495,N_4328);
or U7072 (N_7072,N_3869,N_4038);
and U7073 (N_7073,N_4406,N_3355);
nor U7074 (N_7074,N_3324,N_4730);
and U7075 (N_7075,N_2662,N_2824);
nor U7076 (N_7076,N_4689,N_4734);
and U7077 (N_7077,N_3002,N_3042);
and U7078 (N_7078,N_3352,N_3861);
and U7079 (N_7079,N_4635,N_4950);
and U7080 (N_7080,N_4364,N_2798);
and U7081 (N_7081,N_3430,N_3260);
nor U7082 (N_7082,N_3906,N_4078);
nor U7083 (N_7083,N_4547,N_3590);
xor U7084 (N_7084,N_4710,N_4436);
nand U7085 (N_7085,N_4872,N_2796);
and U7086 (N_7086,N_2963,N_3356);
nand U7087 (N_7087,N_3696,N_3814);
or U7088 (N_7088,N_3450,N_4352);
and U7089 (N_7089,N_2796,N_2587);
or U7090 (N_7090,N_3552,N_3541);
or U7091 (N_7091,N_4937,N_4869);
nor U7092 (N_7092,N_2723,N_3970);
nor U7093 (N_7093,N_4090,N_2929);
nor U7094 (N_7094,N_3082,N_3465);
and U7095 (N_7095,N_2534,N_4185);
nand U7096 (N_7096,N_4495,N_3509);
and U7097 (N_7097,N_3369,N_3461);
xnor U7098 (N_7098,N_4017,N_3650);
or U7099 (N_7099,N_2540,N_3862);
or U7100 (N_7100,N_2814,N_2666);
nand U7101 (N_7101,N_4100,N_3482);
and U7102 (N_7102,N_4533,N_2651);
nor U7103 (N_7103,N_4105,N_3207);
and U7104 (N_7104,N_4564,N_3268);
or U7105 (N_7105,N_4812,N_4797);
and U7106 (N_7106,N_4373,N_3495);
nand U7107 (N_7107,N_2517,N_3600);
nor U7108 (N_7108,N_3168,N_4543);
or U7109 (N_7109,N_2587,N_3251);
nand U7110 (N_7110,N_3019,N_3402);
and U7111 (N_7111,N_2924,N_3442);
nor U7112 (N_7112,N_2726,N_3295);
nor U7113 (N_7113,N_2921,N_3187);
nor U7114 (N_7114,N_4113,N_4244);
xor U7115 (N_7115,N_3800,N_3224);
nor U7116 (N_7116,N_4022,N_3758);
or U7117 (N_7117,N_3227,N_4827);
nor U7118 (N_7118,N_3749,N_2859);
nand U7119 (N_7119,N_2586,N_4860);
and U7120 (N_7120,N_4320,N_3828);
nand U7121 (N_7121,N_4251,N_3148);
and U7122 (N_7122,N_4728,N_2547);
or U7123 (N_7123,N_4749,N_3057);
nor U7124 (N_7124,N_2827,N_4647);
or U7125 (N_7125,N_4047,N_4391);
or U7126 (N_7126,N_3731,N_4430);
or U7127 (N_7127,N_4842,N_2633);
and U7128 (N_7128,N_3904,N_4685);
nand U7129 (N_7129,N_3615,N_3111);
nor U7130 (N_7130,N_3948,N_4428);
and U7131 (N_7131,N_2735,N_2711);
or U7132 (N_7132,N_3807,N_3344);
nor U7133 (N_7133,N_4373,N_4152);
xnor U7134 (N_7134,N_2761,N_2996);
nor U7135 (N_7135,N_2941,N_4362);
nor U7136 (N_7136,N_2730,N_2902);
and U7137 (N_7137,N_4562,N_3540);
nand U7138 (N_7138,N_4322,N_3943);
and U7139 (N_7139,N_4757,N_2866);
and U7140 (N_7140,N_3683,N_3576);
nand U7141 (N_7141,N_4538,N_4244);
and U7142 (N_7142,N_2942,N_3408);
and U7143 (N_7143,N_3513,N_3436);
nor U7144 (N_7144,N_3240,N_4712);
nor U7145 (N_7145,N_3291,N_2845);
or U7146 (N_7146,N_2665,N_3661);
nor U7147 (N_7147,N_4264,N_3098);
or U7148 (N_7148,N_2965,N_3616);
and U7149 (N_7149,N_3933,N_2844);
and U7150 (N_7150,N_3233,N_3553);
nand U7151 (N_7151,N_3689,N_3083);
and U7152 (N_7152,N_3929,N_3539);
and U7153 (N_7153,N_3112,N_4663);
or U7154 (N_7154,N_3741,N_2584);
nand U7155 (N_7155,N_2938,N_3310);
or U7156 (N_7156,N_4374,N_3538);
nand U7157 (N_7157,N_4014,N_4723);
nor U7158 (N_7158,N_4187,N_2641);
nor U7159 (N_7159,N_3600,N_3750);
and U7160 (N_7160,N_3213,N_3637);
nand U7161 (N_7161,N_4526,N_3073);
or U7162 (N_7162,N_2551,N_4337);
or U7163 (N_7163,N_3970,N_2661);
nand U7164 (N_7164,N_4702,N_3154);
or U7165 (N_7165,N_3201,N_4008);
nand U7166 (N_7166,N_4009,N_4202);
nand U7167 (N_7167,N_4854,N_2650);
or U7168 (N_7168,N_4280,N_4902);
or U7169 (N_7169,N_3679,N_2680);
and U7170 (N_7170,N_3662,N_4928);
nand U7171 (N_7171,N_3955,N_3318);
or U7172 (N_7172,N_3323,N_4395);
or U7173 (N_7173,N_3029,N_3207);
nor U7174 (N_7174,N_3297,N_4279);
and U7175 (N_7175,N_2583,N_2835);
or U7176 (N_7176,N_2642,N_2896);
nor U7177 (N_7177,N_4119,N_4515);
or U7178 (N_7178,N_2741,N_3056);
or U7179 (N_7179,N_2885,N_2612);
or U7180 (N_7180,N_3648,N_4206);
and U7181 (N_7181,N_3094,N_3157);
and U7182 (N_7182,N_3227,N_4096);
or U7183 (N_7183,N_4203,N_3803);
xnor U7184 (N_7184,N_4373,N_3176);
or U7185 (N_7185,N_2572,N_4388);
and U7186 (N_7186,N_4747,N_4141);
nor U7187 (N_7187,N_2935,N_3789);
nand U7188 (N_7188,N_4305,N_4117);
nand U7189 (N_7189,N_3973,N_4041);
nand U7190 (N_7190,N_4447,N_4028);
nand U7191 (N_7191,N_3284,N_3307);
nand U7192 (N_7192,N_3085,N_4591);
and U7193 (N_7193,N_3410,N_3465);
and U7194 (N_7194,N_3003,N_2748);
and U7195 (N_7195,N_2818,N_3799);
or U7196 (N_7196,N_4697,N_2690);
and U7197 (N_7197,N_4921,N_4625);
and U7198 (N_7198,N_3670,N_3832);
or U7199 (N_7199,N_4404,N_3970);
nor U7200 (N_7200,N_3039,N_2537);
nand U7201 (N_7201,N_3940,N_2520);
nor U7202 (N_7202,N_4902,N_3356);
nor U7203 (N_7203,N_3516,N_3611);
or U7204 (N_7204,N_4729,N_4279);
nor U7205 (N_7205,N_3264,N_4037);
and U7206 (N_7206,N_2642,N_4229);
xnor U7207 (N_7207,N_4196,N_4214);
xor U7208 (N_7208,N_4762,N_3909);
nor U7209 (N_7209,N_3294,N_4934);
and U7210 (N_7210,N_3246,N_4879);
nor U7211 (N_7211,N_2795,N_4816);
and U7212 (N_7212,N_2617,N_3477);
or U7213 (N_7213,N_3432,N_4993);
nand U7214 (N_7214,N_2517,N_4776);
and U7215 (N_7215,N_3345,N_2824);
or U7216 (N_7216,N_3820,N_2900);
nor U7217 (N_7217,N_4495,N_3976);
or U7218 (N_7218,N_2531,N_2672);
nand U7219 (N_7219,N_4332,N_4249);
or U7220 (N_7220,N_3336,N_3621);
nand U7221 (N_7221,N_4409,N_3294);
nand U7222 (N_7222,N_4360,N_3156);
and U7223 (N_7223,N_4056,N_3190);
nand U7224 (N_7224,N_3391,N_4591);
nand U7225 (N_7225,N_4826,N_2605);
nand U7226 (N_7226,N_3914,N_4771);
nor U7227 (N_7227,N_4225,N_3936);
and U7228 (N_7228,N_2767,N_3796);
and U7229 (N_7229,N_4915,N_4969);
and U7230 (N_7230,N_3123,N_3956);
xnor U7231 (N_7231,N_2521,N_4626);
nand U7232 (N_7232,N_3953,N_2513);
nor U7233 (N_7233,N_4421,N_4389);
and U7234 (N_7234,N_4438,N_2614);
or U7235 (N_7235,N_3536,N_4586);
and U7236 (N_7236,N_3630,N_4989);
and U7237 (N_7237,N_4916,N_2921);
or U7238 (N_7238,N_3335,N_3968);
or U7239 (N_7239,N_2784,N_2672);
nand U7240 (N_7240,N_4164,N_2914);
nor U7241 (N_7241,N_4516,N_3654);
or U7242 (N_7242,N_3958,N_3288);
and U7243 (N_7243,N_2964,N_4305);
or U7244 (N_7244,N_3464,N_2838);
nand U7245 (N_7245,N_3043,N_4899);
nor U7246 (N_7246,N_3815,N_4031);
nand U7247 (N_7247,N_4989,N_4565);
nor U7248 (N_7248,N_2901,N_3110);
or U7249 (N_7249,N_3101,N_3695);
or U7250 (N_7250,N_3994,N_4272);
nand U7251 (N_7251,N_4571,N_3741);
nand U7252 (N_7252,N_2718,N_2949);
nor U7253 (N_7253,N_4760,N_3650);
nor U7254 (N_7254,N_3816,N_3543);
nor U7255 (N_7255,N_4286,N_3761);
and U7256 (N_7256,N_3999,N_3718);
and U7257 (N_7257,N_4228,N_3397);
and U7258 (N_7258,N_3417,N_3198);
and U7259 (N_7259,N_3210,N_3217);
nand U7260 (N_7260,N_2573,N_2822);
or U7261 (N_7261,N_3251,N_3392);
or U7262 (N_7262,N_3087,N_4201);
nor U7263 (N_7263,N_2798,N_3922);
nand U7264 (N_7264,N_3494,N_4976);
nand U7265 (N_7265,N_4293,N_4353);
and U7266 (N_7266,N_3344,N_3663);
and U7267 (N_7267,N_2916,N_2912);
nand U7268 (N_7268,N_3566,N_3692);
or U7269 (N_7269,N_4452,N_4511);
nor U7270 (N_7270,N_4488,N_3626);
nand U7271 (N_7271,N_4169,N_4267);
or U7272 (N_7272,N_3672,N_3772);
nand U7273 (N_7273,N_3125,N_3765);
or U7274 (N_7274,N_3576,N_4650);
nor U7275 (N_7275,N_2805,N_3955);
nor U7276 (N_7276,N_4217,N_2662);
or U7277 (N_7277,N_2753,N_4889);
nor U7278 (N_7278,N_3236,N_3109);
nor U7279 (N_7279,N_3207,N_4861);
or U7280 (N_7280,N_3547,N_3928);
or U7281 (N_7281,N_3307,N_2554);
and U7282 (N_7282,N_4042,N_3888);
nor U7283 (N_7283,N_4881,N_3051);
and U7284 (N_7284,N_4246,N_2541);
and U7285 (N_7285,N_3382,N_2886);
nor U7286 (N_7286,N_3583,N_3851);
and U7287 (N_7287,N_3198,N_3694);
nor U7288 (N_7288,N_3597,N_3897);
or U7289 (N_7289,N_2831,N_3516);
nor U7290 (N_7290,N_3692,N_3229);
or U7291 (N_7291,N_4731,N_4013);
nor U7292 (N_7292,N_3277,N_4818);
and U7293 (N_7293,N_3958,N_4139);
or U7294 (N_7294,N_2919,N_3352);
or U7295 (N_7295,N_2612,N_4284);
or U7296 (N_7296,N_3116,N_4994);
or U7297 (N_7297,N_3088,N_4727);
and U7298 (N_7298,N_3837,N_3013);
nor U7299 (N_7299,N_4820,N_2678);
or U7300 (N_7300,N_3913,N_4206);
nor U7301 (N_7301,N_3271,N_4529);
nor U7302 (N_7302,N_3058,N_3097);
nor U7303 (N_7303,N_3514,N_2582);
or U7304 (N_7304,N_4979,N_4420);
nor U7305 (N_7305,N_3732,N_3357);
nand U7306 (N_7306,N_4324,N_3640);
nor U7307 (N_7307,N_4958,N_4492);
or U7308 (N_7308,N_3213,N_4147);
or U7309 (N_7309,N_2782,N_4256);
nand U7310 (N_7310,N_4322,N_3017);
nand U7311 (N_7311,N_4075,N_4987);
and U7312 (N_7312,N_4802,N_3775);
and U7313 (N_7313,N_3366,N_2710);
nor U7314 (N_7314,N_2913,N_4133);
nor U7315 (N_7315,N_3705,N_2972);
and U7316 (N_7316,N_3538,N_3357);
xnor U7317 (N_7317,N_3415,N_4872);
nor U7318 (N_7318,N_3493,N_2961);
nor U7319 (N_7319,N_4602,N_3787);
xnor U7320 (N_7320,N_3392,N_4028);
nor U7321 (N_7321,N_2715,N_3675);
xnor U7322 (N_7322,N_2774,N_4612);
nor U7323 (N_7323,N_2786,N_3470);
and U7324 (N_7324,N_4554,N_4842);
and U7325 (N_7325,N_4275,N_3419);
nand U7326 (N_7326,N_4314,N_4683);
nand U7327 (N_7327,N_4704,N_4622);
and U7328 (N_7328,N_3181,N_4618);
xor U7329 (N_7329,N_3212,N_3053);
or U7330 (N_7330,N_3594,N_2632);
nor U7331 (N_7331,N_4717,N_3867);
nand U7332 (N_7332,N_4236,N_3373);
or U7333 (N_7333,N_3961,N_4623);
nand U7334 (N_7334,N_4394,N_3739);
nand U7335 (N_7335,N_4407,N_3845);
nand U7336 (N_7336,N_4016,N_4819);
nand U7337 (N_7337,N_4902,N_2818);
and U7338 (N_7338,N_4245,N_4717);
or U7339 (N_7339,N_2631,N_2993);
or U7340 (N_7340,N_3984,N_3319);
nor U7341 (N_7341,N_2739,N_2517);
nor U7342 (N_7342,N_4560,N_3274);
nor U7343 (N_7343,N_3427,N_3638);
nor U7344 (N_7344,N_3128,N_4451);
nor U7345 (N_7345,N_2572,N_4488);
and U7346 (N_7346,N_3468,N_3289);
nor U7347 (N_7347,N_2586,N_2567);
or U7348 (N_7348,N_3142,N_3462);
nand U7349 (N_7349,N_4776,N_3493);
or U7350 (N_7350,N_2621,N_3481);
and U7351 (N_7351,N_3194,N_4906);
nor U7352 (N_7352,N_4744,N_3765);
or U7353 (N_7353,N_3310,N_4230);
nand U7354 (N_7354,N_2883,N_4322);
and U7355 (N_7355,N_4714,N_3945);
or U7356 (N_7356,N_3621,N_3125);
nor U7357 (N_7357,N_2896,N_2742);
nor U7358 (N_7358,N_3137,N_4723);
and U7359 (N_7359,N_4257,N_4141);
or U7360 (N_7360,N_3277,N_3395);
nor U7361 (N_7361,N_4887,N_3756);
nand U7362 (N_7362,N_4738,N_2518);
or U7363 (N_7363,N_4136,N_4411);
and U7364 (N_7364,N_4874,N_2556);
or U7365 (N_7365,N_4934,N_2908);
nand U7366 (N_7366,N_4211,N_4596);
or U7367 (N_7367,N_3598,N_3605);
and U7368 (N_7368,N_3148,N_2737);
or U7369 (N_7369,N_3649,N_3633);
nand U7370 (N_7370,N_2722,N_3498);
or U7371 (N_7371,N_3385,N_4656);
and U7372 (N_7372,N_3373,N_4539);
nand U7373 (N_7373,N_4561,N_3364);
nand U7374 (N_7374,N_4567,N_2999);
and U7375 (N_7375,N_2628,N_4556);
nand U7376 (N_7376,N_2941,N_2717);
or U7377 (N_7377,N_4676,N_4872);
and U7378 (N_7378,N_3372,N_3079);
nor U7379 (N_7379,N_4024,N_4063);
and U7380 (N_7380,N_2771,N_3065);
or U7381 (N_7381,N_4056,N_4833);
or U7382 (N_7382,N_3842,N_3123);
or U7383 (N_7383,N_3363,N_4294);
nor U7384 (N_7384,N_3738,N_4988);
nor U7385 (N_7385,N_3611,N_4044);
nor U7386 (N_7386,N_4343,N_4817);
or U7387 (N_7387,N_2677,N_3691);
nor U7388 (N_7388,N_3239,N_3937);
or U7389 (N_7389,N_4337,N_2787);
nor U7390 (N_7390,N_2761,N_3004);
nor U7391 (N_7391,N_3602,N_4230);
or U7392 (N_7392,N_4032,N_2797);
nand U7393 (N_7393,N_4052,N_4678);
nor U7394 (N_7394,N_4864,N_3606);
nor U7395 (N_7395,N_3469,N_4119);
and U7396 (N_7396,N_3863,N_2947);
xor U7397 (N_7397,N_3410,N_4974);
or U7398 (N_7398,N_3257,N_4718);
or U7399 (N_7399,N_4117,N_2594);
or U7400 (N_7400,N_3182,N_3570);
nand U7401 (N_7401,N_2786,N_3680);
nand U7402 (N_7402,N_2879,N_4661);
and U7403 (N_7403,N_4755,N_3036);
nor U7404 (N_7404,N_2585,N_4981);
or U7405 (N_7405,N_4522,N_4965);
nor U7406 (N_7406,N_3944,N_2767);
and U7407 (N_7407,N_4218,N_4523);
nor U7408 (N_7408,N_2541,N_2711);
and U7409 (N_7409,N_3936,N_2847);
nor U7410 (N_7410,N_4068,N_3523);
xnor U7411 (N_7411,N_4248,N_3169);
and U7412 (N_7412,N_4043,N_2844);
or U7413 (N_7413,N_2833,N_4247);
nor U7414 (N_7414,N_3095,N_4587);
and U7415 (N_7415,N_4691,N_4500);
and U7416 (N_7416,N_3442,N_3194);
nor U7417 (N_7417,N_4495,N_4317);
or U7418 (N_7418,N_3348,N_3063);
nor U7419 (N_7419,N_2506,N_2721);
and U7420 (N_7420,N_2821,N_3073);
or U7421 (N_7421,N_4704,N_2816);
xnor U7422 (N_7422,N_4671,N_4336);
and U7423 (N_7423,N_3018,N_4523);
and U7424 (N_7424,N_3652,N_2932);
or U7425 (N_7425,N_3016,N_4494);
or U7426 (N_7426,N_2686,N_2665);
nor U7427 (N_7427,N_4038,N_2525);
nor U7428 (N_7428,N_3399,N_3806);
nand U7429 (N_7429,N_3476,N_4860);
nand U7430 (N_7430,N_4205,N_3880);
or U7431 (N_7431,N_3485,N_4310);
or U7432 (N_7432,N_2614,N_4790);
nor U7433 (N_7433,N_3851,N_3081);
xnor U7434 (N_7434,N_3556,N_3731);
or U7435 (N_7435,N_3325,N_2966);
nand U7436 (N_7436,N_2838,N_4827);
xor U7437 (N_7437,N_4535,N_3638);
or U7438 (N_7438,N_3915,N_2710);
nand U7439 (N_7439,N_4287,N_4244);
or U7440 (N_7440,N_2534,N_2591);
nand U7441 (N_7441,N_2768,N_4012);
nand U7442 (N_7442,N_4185,N_4883);
nand U7443 (N_7443,N_3240,N_3179);
nand U7444 (N_7444,N_3245,N_3702);
nor U7445 (N_7445,N_4364,N_4235);
nor U7446 (N_7446,N_4896,N_3622);
nand U7447 (N_7447,N_4658,N_3895);
or U7448 (N_7448,N_3288,N_3840);
nand U7449 (N_7449,N_2922,N_3946);
and U7450 (N_7450,N_4048,N_4295);
and U7451 (N_7451,N_4098,N_3773);
nor U7452 (N_7452,N_3666,N_4471);
or U7453 (N_7453,N_4672,N_4196);
nand U7454 (N_7454,N_4113,N_3921);
and U7455 (N_7455,N_4351,N_2932);
nand U7456 (N_7456,N_3476,N_3106);
nor U7457 (N_7457,N_4752,N_2824);
or U7458 (N_7458,N_3526,N_3607);
nand U7459 (N_7459,N_3895,N_4112);
nor U7460 (N_7460,N_4041,N_4819);
or U7461 (N_7461,N_3534,N_3617);
nor U7462 (N_7462,N_2578,N_4826);
and U7463 (N_7463,N_4932,N_3865);
or U7464 (N_7464,N_4547,N_3254);
nand U7465 (N_7465,N_3296,N_4749);
or U7466 (N_7466,N_4060,N_2638);
nor U7467 (N_7467,N_3230,N_4338);
nand U7468 (N_7468,N_2796,N_2605);
or U7469 (N_7469,N_2713,N_2649);
nor U7470 (N_7470,N_3635,N_4590);
or U7471 (N_7471,N_3299,N_3785);
nand U7472 (N_7472,N_4015,N_4758);
or U7473 (N_7473,N_2551,N_2915);
nor U7474 (N_7474,N_3328,N_3888);
and U7475 (N_7475,N_4365,N_3488);
or U7476 (N_7476,N_4292,N_3317);
nor U7477 (N_7477,N_2751,N_3744);
or U7478 (N_7478,N_4548,N_2745);
xor U7479 (N_7479,N_3630,N_2981);
nor U7480 (N_7480,N_4490,N_2652);
nor U7481 (N_7481,N_3493,N_2578);
or U7482 (N_7482,N_3300,N_2860);
nor U7483 (N_7483,N_3487,N_4751);
and U7484 (N_7484,N_4064,N_4265);
nor U7485 (N_7485,N_4646,N_4997);
and U7486 (N_7486,N_3565,N_3321);
nor U7487 (N_7487,N_4949,N_2742);
or U7488 (N_7488,N_3707,N_4254);
nor U7489 (N_7489,N_2535,N_3568);
nor U7490 (N_7490,N_3835,N_4496);
nand U7491 (N_7491,N_4757,N_2566);
nor U7492 (N_7492,N_4176,N_3268);
or U7493 (N_7493,N_4310,N_3482);
nand U7494 (N_7494,N_2893,N_4487);
nor U7495 (N_7495,N_3125,N_4895);
and U7496 (N_7496,N_2602,N_3080);
and U7497 (N_7497,N_4318,N_3856);
or U7498 (N_7498,N_4766,N_3744);
nand U7499 (N_7499,N_4861,N_4678);
nand U7500 (N_7500,N_6547,N_6112);
nor U7501 (N_7501,N_7209,N_6932);
or U7502 (N_7502,N_6132,N_5667);
nand U7503 (N_7503,N_5367,N_5266);
nor U7504 (N_7504,N_7484,N_5985);
xnor U7505 (N_7505,N_6472,N_5861);
nor U7506 (N_7506,N_5601,N_7411);
and U7507 (N_7507,N_5345,N_6442);
and U7508 (N_7508,N_5475,N_6619);
nor U7509 (N_7509,N_5876,N_7111);
nand U7510 (N_7510,N_6174,N_6155);
nor U7511 (N_7511,N_6435,N_5725);
nor U7512 (N_7512,N_5798,N_5931);
and U7513 (N_7513,N_5585,N_5776);
and U7514 (N_7514,N_7454,N_5070);
or U7515 (N_7515,N_5171,N_5088);
nor U7516 (N_7516,N_5384,N_6072);
nor U7517 (N_7517,N_6454,N_6613);
nand U7518 (N_7518,N_6737,N_7308);
or U7519 (N_7519,N_5193,N_5594);
and U7520 (N_7520,N_6245,N_5028);
nor U7521 (N_7521,N_7362,N_5421);
nand U7522 (N_7522,N_7207,N_7139);
nor U7523 (N_7523,N_7155,N_5174);
nand U7524 (N_7524,N_5838,N_6432);
and U7525 (N_7525,N_7266,N_6556);
nor U7526 (N_7526,N_7168,N_7007);
nor U7527 (N_7527,N_7045,N_5511);
nand U7528 (N_7528,N_6934,N_6709);
nand U7529 (N_7529,N_6525,N_5325);
nand U7530 (N_7530,N_5790,N_6942);
and U7531 (N_7531,N_7493,N_7414);
nand U7532 (N_7532,N_5843,N_6748);
nor U7533 (N_7533,N_6597,N_6551);
nand U7534 (N_7534,N_5259,N_5900);
nand U7535 (N_7535,N_5600,N_6183);
or U7536 (N_7536,N_6289,N_6608);
nor U7537 (N_7537,N_5117,N_6614);
nand U7538 (N_7538,N_5777,N_6032);
and U7539 (N_7539,N_6874,N_6450);
and U7540 (N_7540,N_5015,N_7393);
xor U7541 (N_7541,N_6688,N_6424);
nand U7542 (N_7542,N_5632,N_5265);
nor U7543 (N_7543,N_5057,N_6728);
nand U7544 (N_7544,N_7284,N_5822);
or U7545 (N_7545,N_5290,N_6052);
or U7546 (N_7546,N_6576,N_6136);
nor U7547 (N_7547,N_5401,N_5033);
and U7548 (N_7548,N_7213,N_7018);
or U7549 (N_7549,N_6171,N_5187);
or U7550 (N_7550,N_5394,N_6740);
nand U7551 (N_7551,N_5574,N_6528);
and U7552 (N_7552,N_6234,N_5727);
and U7553 (N_7553,N_6128,N_6115);
or U7554 (N_7554,N_6485,N_5014);
nor U7555 (N_7555,N_6302,N_6683);
and U7556 (N_7556,N_6900,N_6014);
nor U7557 (N_7557,N_7053,N_6227);
xnor U7558 (N_7558,N_6361,N_7200);
and U7559 (N_7559,N_6904,N_5583);
nor U7560 (N_7560,N_5506,N_7442);
and U7561 (N_7561,N_5832,N_6458);
xor U7562 (N_7562,N_5796,N_5521);
and U7563 (N_7563,N_6671,N_5605);
nor U7564 (N_7564,N_5108,N_5185);
or U7565 (N_7565,N_6789,N_7447);
nor U7566 (N_7566,N_6827,N_6020);
and U7567 (N_7567,N_5126,N_6978);
and U7568 (N_7568,N_5502,N_7022);
nand U7569 (N_7569,N_6639,N_5012);
and U7570 (N_7570,N_5955,N_6263);
nor U7571 (N_7571,N_7378,N_6929);
and U7572 (N_7572,N_6856,N_6955);
or U7573 (N_7573,N_6021,N_6345);
and U7574 (N_7574,N_7314,N_6566);
and U7575 (N_7575,N_5525,N_6714);
or U7576 (N_7576,N_7462,N_5633);
or U7577 (N_7577,N_6684,N_6393);
nand U7578 (N_7578,N_5204,N_7352);
nor U7579 (N_7579,N_7142,N_5535);
or U7580 (N_7580,N_6785,N_7028);
nand U7581 (N_7581,N_7216,N_7010);
and U7582 (N_7582,N_6126,N_5486);
nor U7583 (N_7583,N_6501,N_6122);
nor U7584 (N_7584,N_6775,N_6086);
and U7585 (N_7585,N_5903,N_5986);
and U7586 (N_7586,N_6570,N_6178);
or U7587 (N_7587,N_5348,N_5901);
nor U7588 (N_7588,N_5139,N_5013);
xor U7589 (N_7589,N_6506,N_5806);
nand U7590 (N_7590,N_5041,N_5217);
nor U7591 (N_7591,N_6217,N_6793);
nor U7592 (N_7592,N_5571,N_5695);
nor U7593 (N_7593,N_5299,N_5890);
and U7594 (N_7594,N_5899,N_7012);
or U7595 (N_7595,N_6726,N_5462);
and U7596 (N_7596,N_5690,N_5984);
xnor U7597 (N_7597,N_5336,N_7339);
nand U7598 (N_7598,N_6257,N_6080);
or U7599 (N_7599,N_5485,N_6776);
nor U7600 (N_7600,N_6814,N_5177);
nand U7601 (N_7601,N_5040,N_6412);
and U7602 (N_7602,N_6866,N_6716);
nor U7603 (N_7603,N_5522,N_6865);
nand U7604 (N_7604,N_5891,N_6455);
xnor U7605 (N_7605,N_6228,N_6969);
nor U7606 (N_7606,N_6146,N_6009);
or U7607 (N_7607,N_5868,N_5073);
and U7608 (N_7608,N_6137,N_5815);
or U7609 (N_7609,N_7077,N_5849);
nor U7610 (N_7610,N_5879,N_5907);
nand U7611 (N_7611,N_7354,N_5129);
or U7612 (N_7612,N_5377,N_6784);
and U7613 (N_7613,N_5779,N_6144);
and U7614 (N_7614,N_6078,N_7319);
and U7615 (N_7615,N_7477,N_7452);
or U7616 (N_7616,N_6051,N_7222);
and U7617 (N_7617,N_6885,N_6670);
and U7618 (N_7618,N_5264,N_7181);
or U7619 (N_7619,N_7166,N_6733);
and U7620 (N_7620,N_7305,N_5051);
nor U7621 (N_7621,N_7151,N_6591);
nor U7622 (N_7622,N_6180,N_6882);
xor U7623 (N_7623,N_5614,N_5215);
and U7624 (N_7624,N_5742,N_5023);
nand U7625 (N_7625,N_6621,N_6190);
nor U7626 (N_7626,N_6140,N_6148);
nand U7627 (N_7627,N_7287,N_6894);
or U7628 (N_7628,N_5257,N_6075);
or U7629 (N_7629,N_5454,N_6836);
nor U7630 (N_7630,N_7434,N_5686);
and U7631 (N_7631,N_7456,N_5653);
and U7632 (N_7632,N_6496,N_5946);
and U7633 (N_7633,N_5789,N_5195);
nor U7634 (N_7634,N_5893,N_5419);
or U7635 (N_7635,N_7299,N_6895);
or U7636 (N_7636,N_6016,N_5810);
nor U7637 (N_7637,N_5763,N_7293);
or U7638 (N_7638,N_7383,N_5182);
and U7639 (N_7639,N_6598,N_6618);
nand U7640 (N_7640,N_6440,N_6892);
nand U7641 (N_7641,N_5697,N_7480);
or U7642 (N_7642,N_6799,N_7020);
nor U7643 (N_7643,N_6518,N_5562);
or U7644 (N_7644,N_5364,N_6073);
nor U7645 (N_7645,N_6792,N_5460);
or U7646 (N_7646,N_7095,N_6915);
nor U7647 (N_7647,N_5563,N_5709);
and U7648 (N_7648,N_6364,N_6077);
xnor U7649 (N_7649,N_7224,N_6341);
nand U7650 (N_7650,N_5423,N_7476);
or U7651 (N_7651,N_5229,N_5038);
or U7652 (N_7652,N_5496,N_6153);
or U7653 (N_7653,N_5218,N_7451);
or U7654 (N_7654,N_6157,N_5479);
nand U7655 (N_7655,N_5524,N_7165);
or U7656 (N_7656,N_7085,N_6891);
and U7657 (N_7657,N_7130,N_6004);
xor U7658 (N_7658,N_5196,N_5778);
and U7659 (N_7659,N_7372,N_6713);
and U7660 (N_7660,N_6343,N_6531);
or U7661 (N_7661,N_6034,N_5314);
nand U7662 (N_7662,N_5783,N_6253);
nand U7663 (N_7663,N_6430,N_5162);
nor U7664 (N_7664,N_5567,N_7178);
nand U7665 (N_7665,N_7078,N_6383);
or U7666 (N_7666,N_7114,N_5349);
nand U7667 (N_7667,N_5378,N_5466);
and U7668 (N_7668,N_6273,N_5141);
and U7669 (N_7669,N_5565,N_5184);
and U7670 (N_7670,N_6757,N_5268);
and U7671 (N_7671,N_6730,N_5029);
nor U7672 (N_7672,N_5211,N_6269);
nor U7673 (N_7673,N_6589,N_7171);
and U7674 (N_7674,N_6351,N_6681);
and U7675 (N_7675,N_6585,N_7107);
or U7676 (N_7676,N_6759,N_6316);
and U7677 (N_7677,N_6642,N_5197);
or U7678 (N_7678,N_6668,N_6047);
nand U7679 (N_7679,N_5555,N_7282);
and U7680 (N_7680,N_6965,N_7080);
nand U7681 (N_7681,N_6087,N_6348);
nor U7682 (N_7682,N_6150,N_6657);
or U7683 (N_7683,N_7251,N_7286);
and U7684 (N_7684,N_5785,N_6067);
nor U7685 (N_7685,N_5214,N_5878);
and U7686 (N_7686,N_5602,N_7348);
nand U7687 (N_7687,N_6797,N_5663);
nand U7688 (N_7688,N_6888,N_6504);
nand U7689 (N_7689,N_6622,N_5249);
or U7690 (N_7690,N_6222,N_7479);
and U7691 (N_7691,N_6049,N_6221);
nand U7692 (N_7692,N_5247,N_6065);
or U7693 (N_7693,N_6421,N_5716);
or U7694 (N_7694,N_7071,N_5880);
nor U7695 (N_7695,N_6444,N_7277);
xnor U7696 (N_7696,N_7360,N_5156);
or U7697 (N_7697,N_6590,N_5418);
nor U7698 (N_7698,N_5176,N_5144);
nor U7699 (N_7699,N_5279,N_5202);
nor U7700 (N_7700,N_6286,N_6391);
and U7701 (N_7701,N_7265,N_7220);
nand U7702 (N_7702,N_5309,N_6889);
nor U7703 (N_7703,N_7173,N_6807);
nand U7704 (N_7704,N_6166,N_6863);
nor U7705 (N_7705,N_6000,N_5760);
nand U7706 (N_7706,N_5769,N_6337);
and U7707 (N_7707,N_7132,N_5085);
or U7708 (N_7708,N_6098,N_7000);
nor U7709 (N_7709,N_7249,N_6970);
nand U7710 (N_7710,N_6327,N_5032);
nand U7711 (N_7711,N_6883,N_6469);
nor U7712 (N_7712,N_5794,N_5019);
or U7713 (N_7713,N_5701,N_6947);
nand U7714 (N_7714,N_7444,N_6609);
nand U7715 (N_7715,N_6890,N_7250);
and U7716 (N_7716,N_7194,N_6854);
nand U7717 (N_7717,N_6511,N_5328);
nand U7718 (N_7718,N_6887,N_5379);
nor U7719 (N_7719,N_6372,N_5362);
nor U7720 (N_7720,N_5741,N_7258);
nor U7721 (N_7721,N_5427,N_6464);
nor U7722 (N_7722,N_5956,N_5319);
or U7723 (N_7723,N_5960,N_5864);
nor U7724 (N_7724,N_6411,N_6489);
or U7725 (N_7725,N_5619,N_5683);
nand U7726 (N_7726,N_6959,N_5731);
and U7727 (N_7727,N_7407,N_6321);
and U7728 (N_7728,N_5618,N_5114);
xor U7729 (N_7729,N_5747,N_5710);
or U7730 (N_7730,N_5316,N_6624);
and U7731 (N_7731,N_6279,N_6937);
nand U7732 (N_7732,N_5078,N_5753);
nor U7733 (N_7733,N_5161,N_5456);
and U7734 (N_7734,N_6040,N_5133);
and U7735 (N_7735,N_5884,N_5160);
and U7736 (N_7736,N_5464,N_6979);
xnor U7737 (N_7737,N_5234,N_6599);
nand U7738 (N_7738,N_5493,N_5998);
or U7739 (N_7739,N_5227,N_7149);
or U7740 (N_7740,N_6405,N_6886);
nand U7741 (N_7741,N_7366,N_6186);
nand U7742 (N_7742,N_6848,N_6207);
xor U7743 (N_7743,N_5654,N_5772);
nand U7744 (N_7744,N_6028,N_6724);
nand U7745 (N_7745,N_7323,N_6416);
and U7746 (N_7746,N_7404,N_5729);
nor U7747 (N_7747,N_5132,N_5065);
xnor U7748 (N_7748,N_5323,N_7494);
or U7749 (N_7749,N_6772,N_6998);
nand U7750 (N_7750,N_5322,N_5934);
or U7751 (N_7751,N_5576,N_5557);
and U7752 (N_7752,N_6818,N_6451);
nand U7753 (N_7753,N_6024,N_5483);
and U7754 (N_7754,N_7295,N_5067);
nor U7755 (N_7755,N_5154,N_6135);
or U7756 (N_7756,N_6203,N_6656);
nand U7757 (N_7757,N_5383,N_5340);
and U7758 (N_7758,N_7312,N_5341);
nor U7759 (N_7759,N_6164,N_5347);
nor U7760 (N_7760,N_5768,N_5665);
xnor U7761 (N_7761,N_6304,N_5406);
or U7762 (N_7762,N_5079,N_6230);
nor U7763 (N_7763,N_6169,N_5397);
nand U7764 (N_7764,N_6353,N_6441);
or U7765 (N_7765,N_6445,N_6834);
nand U7766 (N_7766,N_5577,N_5915);
and U7767 (N_7767,N_7310,N_5740);
nand U7768 (N_7768,N_6971,N_5312);
nand U7769 (N_7769,N_5700,N_5017);
nor U7770 (N_7770,N_6843,N_7497);
or U7771 (N_7771,N_5681,N_6798);
and U7772 (N_7772,N_6840,N_5063);
nor U7773 (N_7773,N_6689,N_5310);
or U7774 (N_7774,N_5646,N_6587);
or U7775 (N_7775,N_5035,N_5009);
nor U7776 (N_7776,N_7488,N_6539);
and U7777 (N_7777,N_6543,N_7174);
and U7778 (N_7778,N_7357,N_5625);
nand U7779 (N_7779,N_6338,N_5242);
nand U7780 (N_7780,N_6344,N_5339);
or U7781 (N_7781,N_6389,N_6336);
and U7782 (N_7782,N_6196,N_7438);
or U7783 (N_7783,N_6787,N_7384);
or U7784 (N_7784,N_7154,N_5717);
nand U7785 (N_7785,N_5267,N_5307);
and U7786 (N_7786,N_6362,N_7375);
or U7787 (N_7787,N_5912,N_5958);
nor U7788 (N_7788,N_6243,N_5640);
and U7789 (N_7789,N_6368,N_7108);
nor U7790 (N_7790,N_5398,N_7070);
nor U7791 (N_7791,N_5848,N_5027);
nand U7792 (N_7792,N_5430,N_5395);
nor U7793 (N_7793,N_5925,N_5820);
nor U7794 (N_7794,N_6452,N_6363);
nand U7795 (N_7795,N_5068,N_6860);
nor U7796 (N_7796,N_5020,N_7148);
and U7797 (N_7797,N_5685,N_7487);
nand U7798 (N_7798,N_5945,N_6718);
nand U7799 (N_7799,N_6750,N_5536);
nand U7800 (N_7800,N_5969,N_7387);
or U7801 (N_7801,N_5971,N_5363);
nor U7802 (N_7802,N_5721,N_6881);
or U7803 (N_7803,N_5745,N_6120);
nand U7804 (N_7804,N_6084,N_6410);
or U7805 (N_7805,N_7292,N_5107);
nand U7806 (N_7806,N_6862,N_5671);
nand U7807 (N_7807,N_6177,N_5509);
nand U7808 (N_7808,N_6679,N_5369);
or U7809 (N_7809,N_6864,N_6513);
or U7810 (N_7810,N_6633,N_5575);
nand U7811 (N_7811,N_6777,N_6572);
nand U7812 (N_7812,N_7096,N_6015);
and U7813 (N_7813,N_5277,N_5262);
or U7814 (N_7814,N_5181,N_5865);
nor U7815 (N_7815,N_5629,N_6082);
or U7816 (N_7816,N_6023,N_5389);
or U7817 (N_7817,N_5857,N_5591);
nor U7818 (N_7818,N_6479,N_5291);
nor U7819 (N_7819,N_6191,N_5708);
and U7820 (N_7820,N_6571,N_6054);
nand U7821 (N_7821,N_5300,N_5411);
nor U7822 (N_7822,N_5975,N_5459);
nor U7823 (N_7823,N_7233,N_7072);
and U7824 (N_7824,N_7042,N_5113);
nand U7825 (N_7825,N_5495,N_6541);
or U7826 (N_7826,N_6267,N_5443);
nor U7827 (N_7827,N_5138,N_5816);
nor U7828 (N_7828,N_6744,N_5782);
nor U7829 (N_7829,N_7202,N_5302);
nor U7830 (N_7830,N_6434,N_6575);
and U7831 (N_7831,N_6595,N_6488);
or U7832 (N_7832,N_7331,N_6703);
or U7833 (N_7833,N_6503,N_7495);
and U7834 (N_7834,N_6992,N_6475);
nand U7835 (N_7835,N_6826,N_6089);
nand U7836 (N_7836,N_6216,N_5544);
and U7837 (N_7837,N_7099,N_5935);
nor U7838 (N_7838,N_7486,N_6235);
nor U7839 (N_7839,N_5659,N_6813);
nand U7840 (N_7840,N_6559,N_5026);
nor U7841 (N_7841,N_5110,N_6630);
and U7842 (N_7842,N_5194,N_6507);
nor U7843 (N_7843,N_5201,N_5586);
or U7844 (N_7844,N_5598,N_6154);
nand U7845 (N_7845,N_5151,N_6844);
nor U7846 (N_7846,N_6335,N_5839);
and U7847 (N_7847,N_7361,N_7203);
nand U7848 (N_7848,N_6181,N_6463);
or U7849 (N_7849,N_7120,N_6113);
xor U7850 (N_7850,N_7026,N_6162);
nand U7851 (N_7851,N_5281,N_5549);
or U7852 (N_7852,N_7433,N_5538);
nor U7853 (N_7853,N_6781,N_6402);
nand U7854 (N_7854,N_5829,N_5966);
nor U7855 (N_7855,N_6495,N_7098);
and U7856 (N_7856,N_5246,N_6097);
and U7857 (N_7857,N_5042,N_6940);
or U7858 (N_7858,N_7380,N_5593);
and U7859 (N_7859,N_5803,N_5682);
or U7860 (N_7860,N_5792,N_7059);
nand U7861 (N_7861,N_5254,N_6175);
or U7862 (N_7862,N_6653,N_6524);
nand U7863 (N_7863,N_6346,N_7272);
or U7864 (N_7864,N_6373,N_5979);
nand U7865 (N_7865,N_5916,N_5275);
nand U7866 (N_7866,N_6011,N_6583);
nor U7867 (N_7867,N_7167,N_5370);
nand U7868 (N_7868,N_6426,N_7214);
nand U7869 (N_7869,N_6991,N_6008);
nor U7870 (N_7870,N_7090,N_6050);
nor U7871 (N_7871,N_7419,N_6557);
nand U7872 (N_7872,N_5136,N_6106);
or U7873 (N_7873,N_6334,N_6006);
nand U7874 (N_7874,N_6835,N_5569);
nor U7875 (N_7875,N_6658,N_5872);
nor U7876 (N_7876,N_5301,N_6220);
nor U7877 (N_7877,N_5664,N_5705);
or U7878 (N_7878,N_5095,N_6069);
nand U7879 (N_7879,N_6938,N_5445);
and U7880 (N_7880,N_6332,N_5457);
and U7881 (N_7881,N_7417,N_7135);
nand U7882 (N_7882,N_6219,N_5351);
nand U7883 (N_7883,N_6107,N_6977);
nand U7884 (N_7884,N_5712,N_7112);
and U7885 (N_7885,N_6118,N_7313);
or U7886 (N_7886,N_5512,N_6218);
nor U7887 (N_7887,N_5327,N_6306);
and U7888 (N_7888,N_5905,N_5155);
nand U7889 (N_7889,N_7037,N_5974);
nor U7890 (N_7890,N_5675,N_5589);
and U7891 (N_7891,N_6825,N_6755);
and U7892 (N_7892,N_5091,N_7475);
nand U7893 (N_7893,N_6857,N_7239);
or U7894 (N_7894,N_6710,N_7386);
and U7895 (N_7895,N_6105,N_5076);
and U7896 (N_7896,N_5561,N_5163);
or U7897 (N_7897,N_6916,N_5635);
or U7898 (N_7898,N_5179,N_5098);
and U7899 (N_7899,N_6339,N_6261);
or U7900 (N_7900,N_6030,N_5170);
and U7901 (N_7901,N_5510,N_6176);
nor U7902 (N_7902,N_6382,N_6920);
and U7903 (N_7903,N_7236,N_5104);
nor U7904 (N_7904,N_6486,N_6918);
nor U7905 (N_7905,N_6094,N_7153);
or U7906 (N_7906,N_5744,N_5944);
nand U7907 (N_7907,N_6909,N_5947);
and U7908 (N_7908,N_6873,N_5866);
nand U7909 (N_7909,N_5704,N_5435);
and U7910 (N_7910,N_6751,N_6201);
nand U7911 (N_7911,N_7358,N_5166);
nand U7912 (N_7912,N_5750,N_5333);
and U7913 (N_7913,N_5147,N_6664);
nor U7914 (N_7914,N_5770,N_5845);
nand U7915 (N_7915,N_5836,N_6019);
nand U7916 (N_7916,N_5018,N_6643);
nor U7917 (N_7917,N_6252,N_5455);
xnor U7918 (N_7918,N_6747,N_6326);
xnor U7919 (N_7919,N_7186,N_5178);
nor U7920 (N_7920,N_5968,N_6439);
nor U7921 (N_7921,N_6872,N_7482);
and U7922 (N_7922,N_5550,N_7334);
nand U7923 (N_7923,N_6982,N_6665);
nand U7924 (N_7924,N_6384,N_5438);
or U7925 (N_7925,N_5006,N_6025);
or U7926 (N_7926,N_7470,N_6617);
nand U7927 (N_7927,N_6502,N_6957);
and U7928 (N_7928,N_5818,N_7322);
and U7929 (N_7929,N_5092,N_6946);
and U7930 (N_7930,N_6563,N_5978);
xnor U7931 (N_7931,N_6552,N_7269);
and U7932 (N_7932,N_6397,N_6066);
or U7933 (N_7933,N_6579,N_5054);
and U7934 (N_7934,N_6232,N_5189);
and U7935 (N_7935,N_6483,N_6482);
or U7936 (N_7936,N_5928,N_5396);
nor U7937 (N_7937,N_5261,N_6480);
or U7938 (N_7938,N_5066,N_5977);
or U7939 (N_7939,N_7371,N_5733);
nor U7940 (N_7940,N_6824,N_6989);
nand U7941 (N_7941,N_5658,N_7136);
nor U7942 (N_7942,N_6884,N_6810);
and U7943 (N_7943,N_6685,N_6871);
and U7944 (N_7944,N_6233,N_7427);
nor U7945 (N_7945,N_6677,N_6379);
nor U7946 (N_7946,N_6448,N_6593);
and U7947 (N_7947,N_6627,N_5850);
and U7948 (N_7948,N_6055,N_5560);
and U7949 (N_7949,N_5424,N_5758);
nor U7950 (N_7950,N_6868,N_7049);
or U7951 (N_7951,N_6509,N_5127);
or U7952 (N_7952,N_7471,N_5096);
nand U7953 (N_7953,N_5273,N_5539);
nand U7954 (N_7954,N_5530,N_7160);
nor U7955 (N_7955,N_6206,N_5886);
nand U7956 (N_7956,N_6095,N_5167);
and U7957 (N_7957,N_6804,N_5375);
or U7958 (N_7958,N_7014,N_5817);
nor U7959 (N_7959,N_7164,N_5883);
or U7960 (N_7960,N_7058,N_5390);
and U7961 (N_7961,N_6644,N_7156);
nand U7962 (N_7962,N_5973,N_6628);
nor U7963 (N_7963,N_6330,N_6297);
nor U7964 (N_7964,N_6375,N_6779);
nor U7965 (N_7965,N_5222,N_5804);
or U7966 (N_7966,N_5405,N_5657);
and U7967 (N_7967,N_7003,N_6377);
nor U7968 (N_7968,N_5149,N_5531);
nand U7969 (N_7969,N_5951,N_6902);
nand U7970 (N_7970,N_7123,N_6702);
or U7971 (N_7971,N_7011,N_7232);
or U7972 (N_7972,N_7199,N_5072);
or U7973 (N_7973,N_7143,N_6851);
and U7974 (N_7974,N_7126,N_6522);
or U7975 (N_7975,N_5797,N_5329);
and U7976 (N_7976,N_5617,N_5702);
nor U7977 (N_7977,N_7385,N_5809);
or U7978 (N_7978,N_6365,N_6961);
or U7979 (N_7979,N_6953,N_6163);
or U7980 (N_7980,N_6035,N_7290);
or U7981 (N_7981,N_7455,N_6223);
or U7982 (N_7982,N_5526,N_5621);
xor U7983 (N_7983,N_6521,N_5735);
or U7984 (N_7984,N_5650,N_6298);
and U7985 (N_7985,N_6548,N_5337);
nand U7986 (N_7986,N_5453,N_7103);
nor U7987 (N_7987,N_7190,N_7106);
and U7988 (N_7988,N_5942,N_6093);
or U7989 (N_7989,N_6114,N_5208);
nand U7990 (N_7990,N_6542,N_6540);
and U7991 (N_7991,N_5458,N_5192);
and U7992 (N_7992,N_7446,N_5644);
and U7993 (N_7993,N_7006,N_6360);
or U7994 (N_7994,N_7278,N_7240);
nand U7995 (N_7995,N_6830,N_7465);
and U7996 (N_7996,N_7219,N_5612);
or U7997 (N_7997,N_5615,N_6285);
and U7998 (N_7998,N_5941,N_6271);
nor U7999 (N_7999,N_6749,N_7122);
nand U8000 (N_8000,N_6960,N_5542);
nor U8001 (N_8001,N_6879,N_5995);
and U8002 (N_8002,N_5470,N_5082);
nand U8003 (N_8003,N_5775,N_7188);
and U8004 (N_8004,N_7307,N_6631);
nor U8005 (N_8005,N_5909,N_5767);
nor U8006 (N_8006,N_5793,N_5230);
nor U8007 (N_8007,N_5965,N_5580);
nor U8008 (N_8008,N_6948,N_6912);
nor U8009 (N_8009,N_5256,N_6817);
and U8010 (N_8010,N_6395,N_6529);
or U8011 (N_8011,N_6850,N_7034);
nor U8012 (N_8012,N_5497,N_5186);
or U8013 (N_8013,N_5637,N_5308);
or U8014 (N_8014,N_5121,N_6041);
and U8015 (N_8015,N_6701,N_5354);
or U8016 (N_8016,N_6038,N_6241);
nand U8017 (N_8017,N_5673,N_6964);
nor U8018 (N_8018,N_6131,N_6380);
nand U8019 (N_8019,N_5918,N_6493);
nor U8020 (N_8020,N_6068,N_6574);
or U8021 (N_8021,N_5624,N_6853);
nand U8022 (N_8022,N_6142,N_6457);
nand U8023 (N_8023,N_5570,N_5010);
or U8024 (N_8024,N_7302,N_6231);
or U8025 (N_8025,N_6340,N_6841);
nor U8026 (N_8026,N_6141,N_5688);
nor U8027 (N_8027,N_5294,N_7056);
and U8028 (N_8028,N_6182,N_7469);
and U8029 (N_8029,N_7088,N_6250);
nand U8030 (N_8030,N_5606,N_5226);
nor U8031 (N_8031,N_5216,N_5800);
and U8032 (N_8032,N_6043,N_7397);
and U8033 (N_8033,N_7311,N_7309);
nor U8034 (N_8034,N_6355,N_5344);
nand U8035 (N_8035,N_7430,N_7032);
and U8036 (N_8036,N_6037,N_5711);
xor U8037 (N_8037,N_5235,N_5558);
or U8038 (N_8038,N_6605,N_6545);
or U8039 (N_8039,N_6108,N_7066);
nor U8040 (N_8040,N_5296,N_6461);
or U8041 (N_8041,N_6046,N_6378);
nor U8042 (N_8042,N_6708,N_6277);
and U8043 (N_8043,N_5691,N_6637);
or U8044 (N_8044,N_7218,N_5655);
or U8045 (N_8045,N_6530,N_5255);
or U8046 (N_8046,N_5599,N_5287);
nor U8047 (N_8047,N_6712,N_6691);
and U8048 (N_8048,N_5620,N_6763);
nor U8049 (N_8049,N_5492,N_7015);
nor U8050 (N_8050,N_6705,N_5751);
nand U8051 (N_8051,N_5209,N_6870);
and U8052 (N_8052,N_5660,N_5158);
and U8053 (N_8053,N_5393,N_5780);
or U8054 (N_8054,N_6550,N_5225);
nor U8055 (N_8055,N_6767,N_6564);
nor U8056 (N_8056,N_6420,N_5446);
nand U8057 (N_8057,N_6822,N_5616);
and U8058 (N_8058,N_5908,N_5252);
nand U8059 (N_8059,N_5873,N_6013);
nand U8060 (N_8060,N_6765,N_5061);
nor U8061 (N_8061,N_7030,N_5205);
nor U8062 (N_8062,N_7445,N_6719);
xnor U8063 (N_8063,N_5648,N_6956);
nand U8064 (N_8064,N_6022,N_7115);
and U8065 (N_8065,N_6453,N_5146);
and U8066 (N_8066,N_6007,N_5272);
nor U8067 (N_8067,N_5168,N_6369);
nand U8068 (N_8068,N_7341,N_6214);
and U8069 (N_8069,N_7198,N_5894);
nand U8070 (N_8070,N_5371,N_7033);
and U8071 (N_8071,N_6031,N_5374);
nor U8072 (N_8072,N_5703,N_6833);
nand U8073 (N_8073,N_5676,N_6845);
or U8074 (N_8074,N_6534,N_5840);
or U8075 (N_8075,N_5052,N_7279);
and U8076 (N_8076,N_6515,N_5352);
nand U8077 (N_8077,N_6739,N_6582);
and U8078 (N_8078,N_7343,N_6695);
or U8079 (N_8079,N_7353,N_7416);
nor U8080 (N_8080,N_7345,N_7196);
nor U8081 (N_8081,N_7390,N_7382);
nand U8082 (N_8082,N_6700,N_5611);
nand U8083 (N_8083,N_6264,N_5784);
or U8084 (N_8084,N_7089,N_6994);
nor U8085 (N_8085,N_7467,N_6492);
nor U8086 (N_8086,N_6949,N_6721);
nor U8087 (N_8087,N_6311,N_6997);
or U8088 (N_8088,N_6735,N_5157);
nand U8089 (N_8089,N_6896,N_6560);
or U8090 (N_8090,N_7074,N_7255);
and U8091 (N_8091,N_6910,N_5100);
and U8092 (N_8092,N_5720,N_5021);
and U8093 (N_8093,N_6972,N_6456);
nor U8094 (N_8094,N_5172,N_5433);
xnor U8095 (N_8095,N_5855,N_6919);
nor U8096 (N_8096,N_6433,N_6152);
nand U8097 (N_8097,N_7254,N_7137);
and U8098 (N_8098,N_7288,N_5922);
nand U8099 (N_8099,N_7350,N_5140);
nand U8100 (N_8100,N_6537,N_7206);
and U8101 (N_8101,N_6010,N_6422);
nand U8102 (N_8102,N_5699,N_7466);
nand U8103 (N_8103,N_6027,N_7276);
or U8104 (N_8104,N_7253,N_5752);
nand U8105 (N_8105,N_5604,N_6811);
nor U8106 (N_8106,N_5221,N_6720);
and U8107 (N_8107,N_6427,N_5271);
xnor U8108 (N_8108,N_5932,N_6562);
and U8109 (N_8109,N_5641,N_7197);
and U8110 (N_8110,N_7027,N_6309);
nand U8111 (N_8111,N_7440,N_5358);
or U8112 (N_8112,N_6669,N_6715);
nor U8113 (N_8113,N_7225,N_6057);
nand U8114 (N_8114,N_6985,N_5191);
nor U8115 (N_8115,N_7415,N_6838);
nor U8116 (N_8116,N_6053,N_7285);
and U8117 (N_8117,N_6808,N_6859);
or U8118 (N_8118,N_6632,N_5484);
and U8119 (N_8119,N_6239,N_6510);
nand U8120 (N_8120,N_5963,N_5305);
xor U8121 (N_8121,N_5097,N_5439);
or U8122 (N_8122,N_7363,N_5833);
and U8123 (N_8123,N_6119,N_6403);
nand U8124 (N_8124,N_6192,N_6244);
or U8125 (N_8125,N_6357,N_5353);
nor U8126 (N_8126,N_6717,N_6476);
and U8127 (N_8127,N_5102,N_6125);
nand U8128 (N_8128,N_5831,N_6242);
nor U8129 (N_8129,N_5387,N_6847);
or U8130 (N_8130,N_5837,N_5578);
nand U8131 (N_8131,N_6268,N_5360);
xor U8132 (N_8132,N_6276,N_5638);
nor U8133 (N_8133,N_5870,N_7187);
nand U8134 (N_8134,N_7210,N_7035);
and U8135 (N_8135,N_6408,N_6921);
nor U8136 (N_8136,N_5283,N_5297);
nand U8137 (N_8137,N_6935,N_7324);
nor U8138 (N_8138,N_7459,N_5643);
and U8139 (N_8139,N_6208,N_5355);
nand U8140 (N_8140,N_6307,N_6990);
nor U8141 (N_8141,N_6036,N_6711);
nor U8142 (N_8142,N_7125,N_5826);
and U8143 (N_8143,N_5888,N_5622);
nor U8144 (N_8144,N_5579,N_7398);
or U8145 (N_8145,N_6736,N_5869);
or U8146 (N_8146,N_6158,N_5004);
and U8147 (N_8147,N_7159,N_7468);
nor U8148 (N_8148,N_5746,N_5278);
nand U8149 (N_8149,N_5630,N_7039);
nand U8150 (N_8150,N_7140,N_6165);
and U8151 (N_8151,N_6555,N_5748);
nor U8152 (N_8152,N_5248,N_5295);
or U8153 (N_8153,N_5519,N_5814);
or U8154 (N_8154,N_5434,N_7483);
nor U8155 (N_8155,N_5011,N_5949);
or U8156 (N_8156,N_5811,N_5060);
and U8157 (N_8157,N_7163,N_6805);
nand U8158 (N_8158,N_5437,N_6867);
and U8159 (N_8159,N_5304,N_5771);
nand U8160 (N_8160,N_7391,N_5694);
or U8161 (N_8161,N_7379,N_7422);
and U8162 (N_8162,N_5967,N_7432);
xor U8163 (N_8163,N_5083,N_6819);
nor U8164 (N_8164,N_6666,N_6565);
nor U8165 (N_8165,N_5180,N_5603);
nand U8166 (N_8166,N_6473,N_6317);
nand U8167 (N_8167,N_5623,N_5842);
nand U8168 (N_8168,N_6400,N_6446);
nand U8169 (N_8169,N_5101,N_6468);
nor U8170 (N_8170,N_6104,N_7489);
nor U8171 (N_8171,N_6652,N_6913);
and U8172 (N_8172,N_6930,N_6324);
or U8173 (N_8173,N_6029,N_5416);
nand U8174 (N_8174,N_7273,N_6923);
nor U8175 (N_8175,N_5053,N_6392);
nor U8176 (N_8176,N_6523,N_5609);
nor U8177 (N_8177,N_5584,N_5099);
or U8178 (N_8178,N_7231,N_6746);
or U8179 (N_8179,N_6266,N_7421);
or U8180 (N_8180,N_6295,N_5568);
nand U8181 (N_8181,N_5749,N_5989);
nor U8182 (N_8182,N_5386,N_7291);
or U8183 (N_8183,N_6941,N_5726);
nor U8184 (N_8184,N_6088,N_7406);
nand U8185 (N_8185,N_5799,N_6404);
nor U8186 (N_8186,N_7212,N_7117);
or U8187 (N_8187,N_5718,N_7062);
and U8188 (N_8188,N_6417,N_5921);
nor U8189 (N_8189,N_5541,N_6625);
and U8190 (N_8190,N_7374,N_7412);
nor U8191 (N_8191,N_6839,N_5980);
or U8192 (N_8192,N_5429,N_7145);
and U8193 (N_8193,N_5902,N_7044);
and U8194 (N_8194,N_5366,N_6880);
or U8195 (N_8195,N_6636,N_5413);
nor U8196 (N_8196,N_6358,N_6320);
nor U8197 (N_8197,N_7113,N_7144);
or U8198 (N_8198,N_7370,N_6151);
and U8199 (N_8199,N_7388,N_6117);
or U8200 (N_8200,N_7150,N_5851);
and U8201 (N_8201,N_7025,N_7458);
or U8202 (N_8202,N_7315,N_6209);
nor U8203 (N_8203,N_6202,N_6260);
nand U8204 (N_8204,N_6976,N_7109);
or U8205 (N_8205,N_5730,N_6161);
and U8206 (N_8206,N_5213,N_6933);
nand U8207 (N_8207,N_6293,N_7264);
nor U8208 (N_8208,N_6837,N_5263);
nand U8209 (N_8209,N_6823,N_6532);
or U8210 (N_8210,N_5206,N_6706);
nand U8211 (N_8211,N_7443,N_5030);
or U8212 (N_8212,N_5403,N_5835);
and U8213 (N_8213,N_6629,N_5228);
nand U8214 (N_8214,N_7141,N_5677);
and U8215 (N_8215,N_6980,N_5473);
or U8216 (N_8216,N_6497,N_6224);
or U8217 (N_8217,N_5852,N_7128);
nor U8218 (N_8218,N_7031,N_5813);
and U8219 (N_8219,N_7102,N_7275);
nand U8220 (N_8220,N_6690,N_5169);
nor U8221 (N_8221,N_6752,N_5338);
nor U8222 (N_8222,N_6988,N_5008);
nor U8223 (N_8223,N_7208,N_5148);
nand U8224 (N_8224,N_6581,N_6725);
or U8225 (N_8225,N_6623,N_6527);
and U8226 (N_8226,N_6663,N_6696);
nand U8227 (N_8227,N_6995,N_5334);
nor U8228 (N_8228,N_7263,N_5128);
and U8229 (N_8229,N_5513,N_5919);
or U8230 (N_8230,N_5001,N_5361);
and U8231 (N_8231,N_5159,N_6963);
or U8232 (N_8232,N_6438,N_5517);
and U8233 (N_8233,N_6213,N_5950);
or U8234 (N_8234,N_5668,N_5410);
or U8235 (N_8235,N_6794,N_7189);
and U8236 (N_8236,N_7496,N_5346);
xor U8237 (N_8237,N_6436,N_7262);
xnor U8238 (N_8238,N_5914,N_7069);
or U8239 (N_8239,N_5972,N_7118);
and U8240 (N_8240,N_6931,N_5592);
nand U8241 (N_8241,N_6655,N_5634);
or U8242 (N_8242,N_7227,N_7230);
or U8243 (N_8243,N_5670,N_6179);
nand U8244 (N_8244,N_5490,N_5996);
nor U8245 (N_8245,N_7040,N_7369);
and U8246 (N_8246,N_5581,N_7175);
and U8247 (N_8247,N_6660,N_6167);
nor U8248 (N_8248,N_6760,N_6620);
or U8249 (N_8249,N_5286,N_5527);
nor U8250 (N_8250,N_7172,N_5626);
nand U8251 (N_8251,N_6399,N_7110);
or U8252 (N_8252,N_5573,N_7211);
nand U8253 (N_8253,N_7296,N_6409);
or U8254 (N_8254,N_5910,N_5392);
nand U8255 (N_8255,N_7351,N_5895);
xor U8256 (N_8256,N_5719,N_6134);
or U8257 (N_8257,N_5723,N_5844);
and U8258 (N_8258,N_5432,N_5188);
nor U8259 (N_8259,N_6648,N_7435);
or U8260 (N_8260,N_5987,N_5442);
nor U8261 (N_8261,N_5824,N_5476);
nand U8262 (N_8262,N_5382,N_5468);
and U8263 (N_8263,N_6901,N_6429);
nand U8264 (N_8264,N_7436,N_6237);
and U8265 (N_8265,N_6795,N_6333);
or U8266 (N_8266,N_6893,N_5090);
nor U8267 (N_8267,N_6875,N_5559);
nand U8268 (N_8268,N_5808,N_7063);
nand U8269 (N_8269,N_5523,N_6908);
nand U8270 (N_8270,N_6606,N_6536);
and U8271 (N_8271,N_7185,N_6225);
xnor U8272 (N_8272,N_5871,N_5858);
nand U8273 (N_8273,N_5465,N_6246);
nor U8274 (N_8274,N_6090,N_7229);
and U8275 (N_8275,N_5022,N_5086);
nor U8276 (N_8276,N_7223,N_6983);
and U8277 (N_8277,N_7437,N_7381);
nand U8278 (N_8278,N_6505,N_6096);
nor U8279 (N_8279,N_7064,N_6698);
nor U8280 (N_8280,N_5518,N_5472);
and U8281 (N_8281,N_5662,N_6160);
nand U8282 (N_8282,N_6519,N_6514);
nand U8283 (N_8283,N_6758,N_5791);
and U8284 (N_8284,N_7023,N_5207);
and U8285 (N_8285,N_5756,N_6602);
or U8286 (N_8286,N_6170,N_6741);
nand U8287 (N_8287,N_5610,N_5724);
nand U8288 (N_8288,N_5292,N_7068);
nand U8289 (N_8289,N_6903,N_5933);
nand U8290 (N_8290,N_6147,N_5331);
xor U8291 (N_8291,N_6756,N_6588);
or U8292 (N_8292,N_6265,N_6676);
or U8293 (N_8293,N_6694,N_5269);
or U8294 (N_8294,N_6301,N_6491);
nor U8295 (N_8295,N_5540,N_6431);
nand U8296 (N_8296,N_6388,N_7330);
nand U8297 (N_8297,N_5130,N_7036);
nand U8298 (N_8298,N_6459,N_5515);
and U8299 (N_8299,N_6962,N_6396);
or U8300 (N_8300,N_6626,N_5467);
nand U8301 (N_8301,N_6842,N_5425);
and U8302 (N_8302,N_5786,N_7338);
and U8303 (N_8303,N_5448,N_5031);
nor U8304 (N_8304,N_5280,N_5200);
nor U8305 (N_8305,N_5080,N_6471);
xnor U8306 (N_8306,N_6356,N_5881);
nor U8307 (N_8307,N_5145,N_6194);
nand U8308 (N_8308,N_7043,N_5330);
nor U8309 (N_8309,N_6314,N_5317);
and U8310 (N_8310,N_5957,N_5111);
nor U8311 (N_8311,N_5651,N_5997);
or U8312 (N_8312,N_5422,N_6993);
or U8313 (N_8313,N_5093,N_6966);
nand U8314 (N_8314,N_6820,N_6484);
and U8315 (N_8315,N_6443,N_5722);
and U8316 (N_8316,N_7177,N_7048);
xnor U8317 (N_8317,N_7337,N_6584);
and U8318 (N_8318,N_7008,N_7481);
or U8319 (N_8319,N_5503,N_7226);
and U8320 (N_8320,N_5084,N_5183);
nand U8321 (N_8321,N_5123,N_6204);
nor U8322 (N_8322,N_5830,N_6638);
xnor U8323 (N_8323,N_6423,N_6470);
or U8324 (N_8324,N_5533,N_7054);
and U8325 (N_8325,N_6743,N_5119);
nand U8326 (N_8326,N_6272,N_5048);
nand U8327 (N_8327,N_7401,N_7002);
or U8328 (N_8328,N_5058,N_6354);
nor U8329 (N_8329,N_7420,N_6615);
nor U8330 (N_8330,N_5692,N_5463);
or U8331 (N_8331,N_7424,N_5135);
and U8332 (N_8332,N_6554,N_5471);
nor U8333 (N_8333,N_5120,N_6258);
and U8334 (N_8334,N_5415,N_6349);
or U8335 (N_8335,N_6791,N_7215);
and U8336 (N_8336,N_6828,N_5190);
and U8337 (N_8337,N_7013,N_6248);
nand U8338 (N_8338,N_6083,N_7134);
nor U8339 (N_8339,N_5923,N_5757);
nand U8340 (N_8340,N_6437,N_5034);
or U8341 (N_8341,N_6924,N_5631);
or U8342 (N_8342,N_5553,N_7234);
nand U8343 (N_8343,N_6291,N_6133);
nand U8344 (N_8344,N_6342,N_5270);
and U8345 (N_8345,N_6282,N_6290);
nand U8346 (N_8346,N_7133,N_7057);
nor U8347 (N_8347,N_7248,N_6414);
nor U8348 (N_8348,N_6764,N_7492);
nand U8349 (N_8349,N_6081,N_5002);
nor U8350 (N_8350,N_5828,N_6952);
or U8351 (N_8351,N_5827,N_5684);
nand U8352 (N_8352,N_7423,N_6193);
or U8353 (N_8353,N_5003,N_5514);
nor U8354 (N_8354,N_5094,N_7389);
nand U8355 (N_8355,N_6060,N_7408);
or U8356 (N_8356,N_5059,N_5628);
nor U8357 (N_8357,N_5669,N_5696);
nand U8358 (N_8358,N_5488,N_5500);
or U8359 (N_8359,N_7298,N_7376);
or U8360 (N_8360,N_6371,N_6498);
and U8361 (N_8361,N_5399,N_5081);
xor U8362 (N_8362,N_5781,N_7152);
nor U8363 (N_8363,N_6103,N_6898);
nand U8364 (N_8364,N_5765,N_6634);
and U8365 (N_8365,N_5388,N_7426);
or U8366 (N_8366,N_7086,N_7146);
nand U8367 (N_8367,N_6048,N_5877);
or U8368 (N_8368,N_6481,N_7256);
and U8369 (N_8369,N_5046,N_7016);
or U8370 (N_8370,N_5687,N_7346);
nor U8371 (N_8371,N_6168,N_6899);
or U8372 (N_8372,N_7499,N_6659);
nand U8373 (N_8373,N_6325,N_7183);
nand U8374 (N_8374,N_6003,N_6544);
nor U8375 (N_8375,N_7019,N_5150);
and U8376 (N_8376,N_6145,N_7359);
nand U8377 (N_8377,N_6200,N_6753);
or U8378 (N_8378,N_5943,N_6056);
nor U8379 (N_8379,N_5841,N_5854);
or U8380 (N_8380,N_5821,N_6329);
nand U8381 (N_8381,N_7448,N_7243);
and U8382 (N_8382,N_6922,N_7405);
nand U8383 (N_8383,N_6517,N_5036);
nor U8384 (N_8384,N_7100,N_6796);
nor U8385 (N_8385,N_7349,N_6549);
and U8386 (N_8386,N_6680,N_6205);
nand U8387 (N_8387,N_6768,N_5245);
or U8388 (N_8388,N_6968,N_6951);
nand U8389 (N_8389,N_6877,N_7268);
nor U8390 (N_8390,N_5994,N_5045);
and U8391 (N_8391,N_6350,N_5556);
nand U8392 (N_8392,N_6533,N_7367);
nand U8393 (N_8393,N_6678,N_7326);
nor U8394 (N_8394,N_6731,N_6447);
nand U8395 (N_8395,N_6033,N_5954);
nand U8396 (N_8396,N_5885,N_7169);
nor U8397 (N_8397,N_6478,N_5450);
or U8398 (N_8398,N_5734,N_5381);
and U8399 (N_8399,N_6367,N_5049);
and U8400 (N_8400,N_6385,N_7176);
nor U8401 (N_8401,N_5649,N_5913);
and U8402 (N_8402,N_5608,N_6771);
and U8403 (N_8403,N_5532,N_5889);
nor U8404 (N_8404,N_5755,N_5250);
nor U8405 (N_8405,N_6769,N_5417);
nand U8406 (N_8406,N_7180,N_6526);
nor U8407 (N_8407,N_6370,N_5543);
nor U8408 (N_8408,N_5860,N_6211);
and U8409 (N_8409,N_6308,N_5385);
nor U8410 (N_8410,N_5489,N_5005);
and U8411 (N_8411,N_6262,N_6926);
or U8412 (N_8412,N_5444,N_6071);
nand U8413 (N_8413,N_7347,N_7394);
nor U8414 (N_8414,N_7038,N_5983);
and U8415 (N_8415,N_6100,N_7046);
nor U8416 (N_8416,N_7335,N_6640);
or U8417 (N_8417,N_6780,N_6778);
nand U8418 (N_8418,N_5738,N_5807);
nand U8419 (N_8419,N_5306,N_6546);
nor U8420 (N_8420,N_5498,N_7373);
and U8421 (N_8421,N_5552,N_6062);
nor U8422 (N_8422,N_5118,N_6195);
or U8423 (N_8423,N_6292,N_5537);
and U8424 (N_8424,N_5115,N_5212);
or U8425 (N_8425,N_6109,N_5874);
nor U8426 (N_8426,N_7336,N_6288);
or U8427 (N_8427,N_5481,N_6199);
nand U8428 (N_8428,N_5203,N_7247);
and U8429 (N_8429,N_5282,N_7260);
or U8430 (N_8430,N_5103,N_7318);
or U8431 (N_8431,N_5258,N_5693);
nand U8432 (N_8432,N_6079,N_5238);
or U8433 (N_8433,N_5474,N_5766);
and U8434 (N_8434,N_5359,N_6462);
nand U8435 (N_8435,N_7195,N_5999);
and U8436 (N_8436,N_6661,N_6376);
nor U8437 (N_8437,N_5551,N_5303);
nand U8438 (N_8438,N_7083,N_7365);
nand U8439 (N_8439,N_6858,N_6592);
or U8440 (N_8440,N_6322,N_6812);
nor U8441 (N_8441,N_5856,N_7097);
nor U8442 (N_8442,N_6359,N_6984);
nand U8443 (N_8443,N_6945,N_7303);
and U8444 (N_8444,N_6635,N_7238);
or U8445 (N_8445,N_6313,N_7441);
or U8446 (N_8446,N_7131,N_5402);
nor U8447 (N_8447,N_5368,N_6328);
or U8448 (N_8448,N_6465,N_6074);
nand U8449 (N_8449,N_5970,N_7170);
or U8450 (N_8450,N_5825,N_6287);
nor U8451 (N_8451,N_6284,N_5240);
and U8452 (N_8452,N_7091,N_6914);
or U8453 (N_8453,N_6352,N_6573);
or U8454 (N_8454,N_7105,N_5823);
nand U8455 (N_8455,N_7368,N_7409);
and U8456 (N_8456,N_5939,N_6732);
or U8457 (N_8457,N_6905,N_5534);
nand U8458 (N_8458,N_6197,N_6236);
or U8459 (N_8459,N_5089,N_6654);
or U8460 (N_8460,N_5636,N_5590);
and U8461 (N_8461,N_7325,N_7270);
and U8462 (N_8462,N_5288,N_5365);
and U8463 (N_8463,N_6604,N_7127);
nand U8464 (N_8464,N_5233,N_7320);
xnor U8465 (N_8465,N_5408,N_5882);
xor U8466 (N_8466,N_5787,N_6607);
or U8467 (N_8467,N_6927,N_6981);
nor U8468 (N_8468,N_5656,N_5689);
nand U8469 (N_8469,N_5477,N_5284);
or U8470 (N_8470,N_7184,N_5896);
nor U8471 (N_8471,N_6723,N_5025);
and U8472 (N_8472,N_6662,N_6401);
nor U8473 (N_8473,N_5122,N_6058);
nor U8474 (N_8474,N_5920,N_6936);
or U8475 (N_8475,N_5834,N_7050);
nand U8476 (N_8476,N_6861,N_5324);
or U8477 (N_8477,N_5953,N_6801);
nor U8478 (N_8478,N_6672,N_5627);
and U8479 (N_8479,N_5074,N_6296);
and U8480 (N_8480,N_5431,N_7129);
nor U8481 (N_8481,N_6975,N_7428);
nand U8482 (N_8482,N_5607,N_7104);
or U8483 (N_8483,N_5243,N_7274);
nor U8484 (N_8484,N_7392,N_5639);
and U8485 (N_8485,N_6939,N_5321);
nor U8486 (N_8486,N_7271,N_6254);
and U8487 (N_8487,N_5528,N_5805);
or U8488 (N_8488,N_6413,N_6907);
nor U8489 (N_8489,N_5237,N_6173);
nor U8490 (N_8490,N_5441,N_7065);
nor U8491 (N_8491,N_5482,N_6829);
xnor U8492 (N_8492,N_6734,N_6110);
and U8493 (N_8493,N_5478,N_7179);
or U8494 (N_8494,N_6596,N_6832);
nor U8495 (N_8495,N_5142,N_6210);
nor U8496 (N_8496,N_5759,N_6123);
and U8497 (N_8497,N_7124,N_7079);
or U8498 (N_8498,N_7364,N_5315);
and U8499 (N_8499,N_5926,N_6419);
xor U8500 (N_8500,N_5862,N_5911);
and U8501 (N_8501,N_7067,N_5311);
and U8502 (N_8502,N_5924,N_7004);
and U8503 (N_8503,N_6070,N_5887);
or U8504 (N_8504,N_6762,N_6121);
and U8505 (N_8505,N_5480,N_5736);
nor U8506 (N_8506,N_6831,N_5773);
and U8507 (N_8507,N_7498,N_6215);
nor U8508 (N_8508,N_7162,N_7242);
nor U8509 (N_8509,N_6586,N_5047);
nor U8510 (N_8510,N_5961,N_5892);
nor U8511 (N_8511,N_5761,N_7425);
nand U8512 (N_8512,N_6143,N_6911);
or U8513 (N_8513,N_6774,N_5173);
nand U8514 (N_8514,N_7439,N_5137);
and U8515 (N_8515,N_5859,N_6092);
or U8516 (N_8516,N_6986,N_6925);
nor U8517 (N_8517,N_7075,N_6578);
nand U8518 (N_8518,N_7147,N_6770);
nand U8519 (N_8519,N_6973,N_5039);
nand U8520 (N_8520,N_7052,N_5508);
nand U8521 (N_8521,N_7205,N_7457);
nand U8522 (N_8522,N_7342,N_7400);
and U8523 (N_8523,N_6682,N_7192);
nand U8524 (N_8524,N_6042,N_6855);
nor U8525 (N_8525,N_6259,N_5743);
and U8526 (N_8526,N_7431,N_7460);
nand U8527 (N_8527,N_5276,N_5373);
nand U8528 (N_8528,N_6226,N_6649);
and U8529 (N_8529,N_6693,N_5545);
and U8530 (N_8530,N_5491,N_5679);
or U8531 (N_8531,N_7017,N_6305);
or U8532 (N_8532,N_7355,N_7138);
nor U8533 (N_8533,N_5596,N_5988);
nand U8534 (N_8534,N_7491,N_5062);
nor U8535 (N_8535,N_5075,N_6766);
nand U8536 (N_8536,N_6650,N_6569);
and U8537 (N_8537,N_6646,N_6538);
or U8538 (N_8538,N_7121,N_6577);
or U8539 (N_8539,N_6647,N_7267);
and U8540 (N_8540,N_5407,N_6603);
nand U8541 (N_8541,N_7084,N_6139);
nor U8542 (N_8542,N_7082,N_5647);
or U8543 (N_8543,N_6600,N_6494);
nor U8544 (N_8544,N_5447,N_6407);
nor U8545 (N_8545,N_5056,N_5802);
nor U8546 (N_8546,N_5666,N_6044);
nor U8547 (N_8547,N_6699,N_7060);
nand U8548 (N_8548,N_7093,N_5964);
and U8549 (N_8549,N_5461,N_6782);
or U8550 (N_8550,N_6783,N_5376);
and U8551 (N_8551,N_5164,N_5112);
and U8552 (N_8552,N_6869,N_5993);
nand U8553 (N_8553,N_5426,N_5595);
or U8554 (N_8554,N_7450,N_7402);
nor U8555 (N_8555,N_6102,N_5210);
xor U8556 (N_8556,N_7304,N_5546);
nand U8557 (N_8557,N_6127,N_6773);
and U8558 (N_8558,N_5064,N_5897);
or U8559 (N_8559,N_7029,N_5754);
or U8560 (N_8560,N_6788,N_5927);
and U8561 (N_8561,N_5812,N_5318);
or U8562 (N_8562,N_6466,N_5713);
or U8563 (N_8563,N_7009,N_5529);
nor U8564 (N_8564,N_5391,N_6745);
nand U8565 (N_8565,N_5853,N_6347);
nor U8566 (N_8566,N_6806,N_6722);
and U8567 (N_8567,N_6821,N_5409);
nor U8568 (N_8568,N_6516,N_5244);
or U8569 (N_8569,N_5285,N_6394);
or U8570 (N_8570,N_5335,N_5116);
nor U8571 (N_8571,N_6188,N_5232);
nand U8572 (N_8572,N_5105,N_5452);
nor U8573 (N_8573,N_5572,N_7116);
nor U8574 (N_8574,N_5343,N_5494);
nor U8575 (N_8575,N_5332,N_7413);
or U8576 (N_8576,N_5420,N_6803);
and U8577 (N_8577,N_5774,N_7395);
or U8578 (N_8578,N_6673,N_6012);
and U8579 (N_8579,N_5982,N_6124);
and U8580 (N_8580,N_7101,N_5106);
or U8581 (N_8581,N_7257,N_5449);
or U8582 (N_8582,N_6026,N_5298);
and U8583 (N_8583,N_6185,N_7280);
or U8584 (N_8584,N_6366,N_6001);
and U8585 (N_8585,N_6101,N_6487);
or U8586 (N_8586,N_5231,N_5372);
nor U8587 (N_8587,N_6601,N_5732);
nor U8588 (N_8588,N_5847,N_6816);
and U8589 (N_8589,N_5412,N_6310);
or U8590 (N_8590,N_5801,N_7061);
nand U8591 (N_8591,N_6508,N_6315);
and U8592 (N_8592,N_5795,N_6686);
and U8593 (N_8593,N_7478,N_5940);
xnor U8594 (N_8594,N_5175,N_5505);
and U8595 (N_8595,N_6172,N_5788);
nor U8596 (N_8596,N_6374,N_7463);
nand U8597 (N_8597,N_7055,N_5069);
or U8598 (N_8598,N_7005,N_5739);
or U8599 (N_8599,N_5936,N_7332);
or U8600 (N_8600,N_6610,N_7294);
or U8601 (N_8601,N_6063,N_5326);
nand U8602 (N_8602,N_5554,N_6386);
nand U8603 (N_8603,N_6727,N_7041);
nand U8604 (N_8604,N_7237,N_5016);
or U8605 (N_8605,N_7301,N_5976);
nor U8606 (N_8606,N_5962,N_6064);
nand U8607 (N_8607,N_5597,N_5224);
and U8608 (N_8608,N_7087,N_7157);
nor U8609 (N_8609,N_7252,N_5404);
nor U8610 (N_8610,N_5320,N_7356);
nor U8611 (N_8611,N_7399,N_5499);
and U8612 (N_8612,N_5645,N_6802);
and U8613 (N_8613,N_6247,N_6212);
nand U8614 (N_8614,N_6256,N_5507);
or U8615 (N_8615,N_6697,N_6418);
or U8616 (N_8616,N_5044,N_6553);
xor U8617 (N_8617,N_5071,N_6312);
and U8618 (N_8618,N_6729,N_6300);
nand U8619 (N_8619,N_5929,N_6499);
or U8620 (N_8620,N_7193,N_5680);
or U8621 (N_8621,N_5737,N_6967);
and U8622 (N_8622,N_7321,N_7228);
and U8623 (N_8623,N_7329,N_7418);
or U8624 (N_8624,N_6943,N_5904);
nand U8625 (N_8625,N_5706,N_6754);
or U8626 (N_8626,N_5152,N_6099);
and U8627 (N_8627,N_6687,N_5674);
nor U8628 (N_8628,N_7001,N_5260);
or U8629 (N_8629,N_6594,N_5863);
or U8630 (N_8630,N_5587,N_5728);
nor U8631 (N_8631,N_5350,N_6240);
or U8632 (N_8632,N_5125,N_6274);
nand U8633 (N_8633,N_6189,N_5055);
and U8634 (N_8634,N_5357,N_6130);
nor U8635 (N_8635,N_5134,N_5077);
nand U8636 (N_8636,N_7340,N_5043);
nor U8637 (N_8637,N_7317,N_6815);
and U8638 (N_8638,N_6876,N_6299);
nand U8639 (N_8639,N_6159,N_6490);
and U8640 (N_8640,N_6275,N_5516);
or U8641 (N_8641,N_6738,N_6800);
or U8642 (N_8642,N_6129,N_6704);
and U8643 (N_8643,N_6005,N_7449);
and U8644 (N_8644,N_5678,N_6283);
or U8645 (N_8645,N_7024,N_5990);
nor U8646 (N_8646,N_6667,N_6255);
and U8647 (N_8647,N_7327,N_5707);
or U8648 (N_8648,N_5661,N_6568);
nor U8649 (N_8649,N_5440,N_5938);
nor U8650 (N_8650,N_6675,N_6002);
nand U8651 (N_8651,N_6580,N_7306);
nand U8652 (N_8652,N_5153,N_7403);
nor U8653 (N_8653,N_6425,N_5867);
nand U8654 (N_8654,N_7051,N_6318);
and U8655 (N_8655,N_7081,N_6928);
and U8656 (N_8656,N_6999,N_6742);
and U8657 (N_8657,N_5220,N_5948);
nand U8658 (N_8658,N_7204,N_6707);
nand U8659 (N_8659,N_6116,N_5251);
nand U8660 (N_8660,N_5652,N_6987);
and U8661 (N_8661,N_7191,N_5582);
nand U8662 (N_8662,N_6852,N_7281);
or U8663 (N_8663,N_6849,N_6561);
nor U8664 (N_8664,N_7473,N_6198);
and U8665 (N_8665,N_7047,N_7259);
nor U8666 (N_8666,N_6474,N_6039);
nand U8667 (N_8667,N_6460,N_5547);
nor U8668 (N_8668,N_7235,N_5548);
nor U8669 (N_8669,N_5356,N_6906);
nor U8670 (N_8670,N_5875,N_6428);
or U8671 (N_8671,N_5050,N_6645);
and U8672 (N_8672,N_6467,N_6651);
nor U8673 (N_8673,N_5898,N_7297);
or U8674 (N_8674,N_6381,N_5672);
xor U8675 (N_8675,N_7461,N_6398);
and U8676 (N_8676,N_6280,N_5143);
or U8677 (N_8677,N_6612,N_6944);
and U8678 (N_8678,N_6512,N_6846);
nand U8679 (N_8679,N_7289,N_6878);
and U8680 (N_8680,N_5642,N_5991);
nor U8681 (N_8681,N_6017,N_7344);
nand U8682 (N_8682,N_7094,N_6149);
nor U8683 (N_8683,N_6156,N_5109);
or U8684 (N_8684,N_6323,N_6786);
or U8685 (N_8685,N_6281,N_7021);
nor U8686 (N_8686,N_5917,N_7073);
or U8687 (N_8687,N_7316,N_5436);
xnor U8688 (N_8688,N_7429,N_7283);
nand U8689 (N_8689,N_5564,N_5236);
and U8690 (N_8690,N_6138,N_6692);
or U8691 (N_8691,N_7092,N_7410);
and U8692 (N_8692,N_6567,N_5131);
or U8693 (N_8693,N_6390,N_7453);
and U8694 (N_8694,N_6958,N_5239);
nand U8695 (N_8695,N_6249,N_5698);
or U8696 (N_8696,N_5380,N_5293);
and U8697 (N_8697,N_5520,N_6294);
or U8698 (N_8698,N_6415,N_7464);
nand U8699 (N_8699,N_6076,N_6061);
nor U8700 (N_8700,N_7333,N_5007);
or U8701 (N_8701,N_5198,N_5274);
and U8702 (N_8702,N_5613,N_5715);
and U8703 (N_8703,N_7241,N_7076);
nand U8704 (N_8704,N_6954,N_7377);
or U8705 (N_8705,N_6059,N_6319);
nor U8706 (N_8706,N_5764,N_7261);
or U8707 (N_8707,N_6238,N_6406);
and U8708 (N_8708,N_6761,N_5024);
nor U8709 (N_8709,N_5819,N_6520);
or U8710 (N_8710,N_6558,N_6045);
or U8711 (N_8711,N_7158,N_5165);
and U8712 (N_8712,N_6996,N_7396);
and U8713 (N_8713,N_5199,N_7474);
or U8714 (N_8714,N_6229,N_5037);
xnor U8715 (N_8715,N_6091,N_6270);
or U8716 (N_8716,N_6917,N_6500);
and U8717 (N_8717,N_6184,N_5762);
nand U8718 (N_8718,N_6085,N_5487);
nand U8719 (N_8719,N_6897,N_5469);
nor U8720 (N_8720,N_6974,N_5959);
nor U8721 (N_8721,N_6674,N_7182);
nor U8722 (N_8722,N_5400,N_6111);
nor U8723 (N_8723,N_5714,N_6535);
nor U8724 (N_8724,N_5428,N_6809);
or U8725 (N_8725,N_7221,N_7245);
nand U8726 (N_8726,N_7217,N_5846);
nor U8727 (N_8727,N_5124,N_5930);
or U8728 (N_8728,N_5087,N_7244);
nor U8729 (N_8729,N_6950,N_5289);
and U8730 (N_8730,N_5937,N_6790);
or U8731 (N_8731,N_6616,N_5313);
and U8732 (N_8732,N_5000,N_7246);
nand U8733 (N_8733,N_6387,N_6477);
nand U8734 (N_8734,N_6331,N_6278);
nand U8735 (N_8735,N_5342,N_5219);
and U8736 (N_8736,N_5414,N_6303);
and U8737 (N_8737,N_5952,N_5588);
nor U8738 (N_8738,N_6449,N_5501);
and U8739 (N_8739,N_6611,N_6251);
nor U8740 (N_8740,N_6641,N_7472);
nor U8741 (N_8741,N_5981,N_7201);
xnor U8742 (N_8742,N_5566,N_7119);
nand U8743 (N_8743,N_5504,N_5241);
nand U8744 (N_8744,N_6018,N_5253);
nand U8745 (N_8745,N_5906,N_5223);
and U8746 (N_8746,N_7485,N_5992);
nor U8747 (N_8747,N_7161,N_5451);
xor U8748 (N_8748,N_7300,N_7490);
nor U8749 (N_8749,N_7328,N_6187);
nor U8750 (N_8750,N_7224,N_6146);
and U8751 (N_8751,N_6609,N_6636);
and U8752 (N_8752,N_5176,N_5575);
or U8753 (N_8753,N_6260,N_6480);
xor U8754 (N_8754,N_6377,N_7028);
nor U8755 (N_8755,N_6730,N_6675);
nand U8756 (N_8756,N_7026,N_5501);
nor U8757 (N_8757,N_5599,N_6561);
or U8758 (N_8758,N_6219,N_7166);
nor U8759 (N_8759,N_5172,N_7485);
and U8760 (N_8760,N_6289,N_6780);
nand U8761 (N_8761,N_7429,N_5139);
or U8762 (N_8762,N_7059,N_6454);
and U8763 (N_8763,N_7136,N_7296);
xor U8764 (N_8764,N_6938,N_6111);
or U8765 (N_8765,N_6185,N_6444);
and U8766 (N_8766,N_6509,N_6077);
nor U8767 (N_8767,N_5816,N_6798);
or U8768 (N_8768,N_7302,N_5181);
nand U8769 (N_8769,N_5506,N_6880);
xor U8770 (N_8770,N_5732,N_6240);
or U8771 (N_8771,N_5212,N_6912);
nor U8772 (N_8772,N_5818,N_6147);
nor U8773 (N_8773,N_6533,N_6733);
or U8774 (N_8774,N_5004,N_5157);
or U8775 (N_8775,N_7246,N_6256);
or U8776 (N_8776,N_6726,N_5030);
nor U8777 (N_8777,N_6431,N_7192);
and U8778 (N_8778,N_6077,N_7277);
nor U8779 (N_8779,N_5693,N_5157);
nor U8780 (N_8780,N_6502,N_6733);
nand U8781 (N_8781,N_6006,N_6323);
or U8782 (N_8782,N_5815,N_6406);
nand U8783 (N_8783,N_7322,N_6610);
nand U8784 (N_8784,N_6890,N_7494);
xor U8785 (N_8785,N_7462,N_6672);
xnor U8786 (N_8786,N_6001,N_6258);
and U8787 (N_8787,N_6295,N_6657);
nor U8788 (N_8788,N_6441,N_7108);
and U8789 (N_8789,N_5668,N_5276);
xnor U8790 (N_8790,N_5931,N_6629);
nor U8791 (N_8791,N_7046,N_7402);
nor U8792 (N_8792,N_7122,N_7101);
xor U8793 (N_8793,N_5077,N_6336);
nor U8794 (N_8794,N_7242,N_6777);
or U8795 (N_8795,N_6885,N_6616);
and U8796 (N_8796,N_6373,N_7304);
nor U8797 (N_8797,N_7441,N_6638);
and U8798 (N_8798,N_5791,N_6385);
nor U8799 (N_8799,N_6496,N_5524);
and U8800 (N_8800,N_7169,N_5851);
nor U8801 (N_8801,N_6096,N_6790);
nor U8802 (N_8802,N_6026,N_6107);
nor U8803 (N_8803,N_5601,N_5575);
nor U8804 (N_8804,N_6187,N_5440);
or U8805 (N_8805,N_5809,N_6510);
and U8806 (N_8806,N_5693,N_5589);
nand U8807 (N_8807,N_7355,N_6318);
nand U8808 (N_8808,N_5285,N_5386);
nand U8809 (N_8809,N_7085,N_7430);
nand U8810 (N_8810,N_6157,N_5737);
nand U8811 (N_8811,N_7208,N_7239);
or U8812 (N_8812,N_5759,N_5157);
or U8813 (N_8813,N_5500,N_5720);
or U8814 (N_8814,N_5281,N_6431);
nor U8815 (N_8815,N_6579,N_7243);
or U8816 (N_8816,N_5458,N_6331);
nor U8817 (N_8817,N_5713,N_5252);
and U8818 (N_8818,N_7476,N_5231);
nor U8819 (N_8819,N_6551,N_6615);
or U8820 (N_8820,N_7032,N_6427);
and U8821 (N_8821,N_6822,N_7176);
nor U8822 (N_8822,N_5896,N_5094);
xor U8823 (N_8823,N_6383,N_7175);
and U8824 (N_8824,N_5529,N_7192);
and U8825 (N_8825,N_5310,N_6473);
and U8826 (N_8826,N_5271,N_6666);
and U8827 (N_8827,N_7077,N_6289);
and U8828 (N_8828,N_5378,N_5577);
and U8829 (N_8829,N_5974,N_7086);
or U8830 (N_8830,N_5299,N_6225);
or U8831 (N_8831,N_5997,N_7178);
nor U8832 (N_8832,N_6438,N_5053);
nand U8833 (N_8833,N_6801,N_7488);
or U8834 (N_8834,N_6959,N_5127);
nor U8835 (N_8835,N_5364,N_6721);
nand U8836 (N_8836,N_5651,N_7446);
and U8837 (N_8837,N_6910,N_5296);
nor U8838 (N_8838,N_5598,N_5012);
nor U8839 (N_8839,N_6739,N_7446);
nand U8840 (N_8840,N_5334,N_7050);
nor U8841 (N_8841,N_5591,N_5248);
xor U8842 (N_8842,N_6531,N_7186);
nand U8843 (N_8843,N_6133,N_6248);
and U8844 (N_8844,N_6662,N_5188);
or U8845 (N_8845,N_5489,N_5388);
nand U8846 (N_8846,N_5765,N_6034);
or U8847 (N_8847,N_5146,N_5226);
nor U8848 (N_8848,N_7474,N_5126);
nand U8849 (N_8849,N_6679,N_5704);
nor U8850 (N_8850,N_5513,N_5632);
or U8851 (N_8851,N_5060,N_5596);
nor U8852 (N_8852,N_5595,N_6968);
and U8853 (N_8853,N_7438,N_6816);
nand U8854 (N_8854,N_6065,N_5072);
or U8855 (N_8855,N_5208,N_6327);
and U8856 (N_8856,N_5639,N_5404);
or U8857 (N_8857,N_6989,N_5484);
nand U8858 (N_8858,N_5376,N_6231);
or U8859 (N_8859,N_6700,N_5152);
and U8860 (N_8860,N_5111,N_6936);
nand U8861 (N_8861,N_6900,N_5182);
or U8862 (N_8862,N_5968,N_5022);
or U8863 (N_8863,N_5558,N_6303);
and U8864 (N_8864,N_7241,N_7385);
nor U8865 (N_8865,N_6080,N_7093);
or U8866 (N_8866,N_7270,N_5036);
and U8867 (N_8867,N_5163,N_6815);
nor U8868 (N_8868,N_6570,N_5678);
or U8869 (N_8869,N_6983,N_5148);
and U8870 (N_8870,N_6497,N_5793);
nor U8871 (N_8871,N_5530,N_5747);
and U8872 (N_8872,N_6338,N_6972);
or U8873 (N_8873,N_5097,N_7449);
or U8874 (N_8874,N_6234,N_5390);
nand U8875 (N_8875,N_6786,N_5786);
nor U8876 (N_8876,N_6473,N_6286);
and U8877 (N_8877,N_6223,N_6200);
or U8878 (N_8878,N_5299,N_5217);
and U8879 (N_8879,N_5459,N_7318);
nor U8880 (N_8880,N_6200,N_6987);
nand U8881 (N_8881,N_6852,N_5450);
and U8882 (N_8882,N_6741,N_6644);
nand U8883 (N_8883,N_5790,N_7269);
nand U8884 (N_8884,N_5961,N_6801);
nor U8885 (N_8885,N_6836,N_6028);
or U8886 (N_8886,N_5079,N_5171);
nor U8887 (N_8887,N_6225,N_5094);
nand U8888 (N_8888,N_6799,N_6175);
and U8889 (N_8889,N_7026,N_6149);
nor U8890 (N_8890,N_6621,N_6614);
nor U8891 (N_8891,N_7290,N_6432);
xor U8892 (N_8892,N_7192,N_5073);
and U8893 (N_8893,N_5861,N_5945);
and U8894 (N_8894,N_5440,N_6260);
or U8895 (N_8895,N_5424,N_6117);
nor U8896 (N_8896,N_5348,N_6789);
or U8897 (N_8897,N_6958,N_6376);
and U8898 (N_8898,N_5361,N_6731);
nor U8899 (N_8899,N_7262,N_5800);
and U8900 (N_8900,N_5772,N_6473);
and U8901 (N_8901,N_6616,N_7170);
and U8902 (N_8902,N_5122,N_6658);
nand U8903 (N_8903,N_6517,N_7324);
nor U8904 (N_8904,N_5802,N_5308);
nor U8905 (N_8905,N_6309,N_7195);
nor U8906 (N_8906,N_5270,N_6373);
nor U8907 (N_8907,N_6784,N_5706);
nand U8908 (N_8908,N_6333,N_6361);
and U8909 (N_8909,N_5409,N_6800);
nor U8910 (N_8910,N_5785,N_5070);
or U8911 (N_8911,N_5593,N_7019);
nand U8912 (N_8912,N_6828,N_6004);
nand U8913 (N_8913,N_5926,N_6917);
or U8914 (N_8914,N_5648,N_7444);
and U8915 (N_8915,N_5295,N_6874);
nand U8916 (N_8916,N_6183,N_5776);
or U8917 (N_8917,N_6888,N_6979);
nor U8918 (N_8918,N_5120,N_5797);
nor U8919 (N_8919,N_6288,N_5304);
or U8920 (N_8920,N_7220,N_6785);
and U8921 (N_8921,N_7319,N_6766);
nand U8922 (N_8922,N_6185,N_6263);
nor U8923 (N_8923,N_7432,N_7132);
nand U8924 (N_8924,N_5065,N_6838);
or U8925 (N_8925,N_7175,N_6066);
or U8926 (N_8926,N_5704,N_6942);
nor U8927 (N_8927,N_5806,N_5720);
and U8928 (N_8928,N_6973,N_5708);
nand U8929 (N_8929,N_5040,N_5864);
and U8930 (N_8930,N_6634,N_5656);
nor U8931 (N_8931,N_7411,N_6962);
nor U8932 (N_8932,N_6445,N_5627);
or U8933 (N_8933,N_6913,N_7410);
nand U8934 (N_8934,N_6836,N_5073);
and U8935 (N_8935,N_7421,N_6046);
or U8936 (N_8936,N_5029,N_5203);
nand U8937 (N_8937,N_5144,N_5754);
and U8938 (N_8938,N_5926,N_6529);
and U8939 (N_8939,N_7426,N_6145);
nand U8940 (N_8940,N_6017,N_6872);
and U8941 (N_8941,N_5270,N_7292);
nor U8942 (N_8942,N_6589,N_5064);
or U8943 (N_8943,N_7476,N_6035);
nand U8944 (N_8944,N_5218,N_6506);
or U8945 (N_8945,N_7035,N_6419);
or U8946 (N_8946,N_6703,N_7100);
nor U8947 (N_8947,N_6879,N_7031);
nand U8948 (N_8948,N_5723,N_5495);
nor U8949 (N_8949,N_6656,N_5141);
or U8950 (N_8950,N_7482,N_5648);
nor U8951 (N_8951,N_5345,N_5386);
nand U8952 (N_8952,N_5333,N_5635);
and U8953 (N_8953,N_5850,N_5124);
and U8954 (N_8954,N_5783,N_5471);
and U8955 (N_8955,N_5404,N_7143);
nor U8956 (N_8956,N_5372,N_6167);
nor U8957 (N_8957,N_5453,N_6438);
and U8958 (N_8958,N_6914,N_7196);
or U8959 (N_8959,N_7102,N_5106);
nor U8960 (N_8960,N_6667,N_7337);
nor U8961 (N_8961,N_5620,N_5683);
nand U8962 (N_8962,N_5532,N_6115);
nand U8963 (N_8963,N_6168,N_5091);
nand U8964 (N_8964,N_6442,N_5986);
nand U8965 (N_8965,N_6506,N_6050);
nand U8966 (N_8966,N_6484,N_7233);
or U8967 (N_8967,N_6323,N_5728);
nand U8968 (N_8968,N_5483,N_7248);
nand U8969 (N_8969,N_5009,N_7139);
or U8970 (N_8970,N_7472,N_5155);
or U8971 (N_8971,N_6292,N_6249);
nor U8972 (N_8972,N_5928,N_5618);
and U8973 (N_8973,N_5249,N_7319);
xnor U8974 (N_8974,N_5791,N_5954);
or U8975 (N_8975,N_5595,N_5592);
and U8976 (N_8976,N_6857,N_6441);
nor U8977 (N_8977,N_5403,N_5613);
or U8978 (N_8978,N_5575,N_6763);
nor U8979 (N_8979,N_7369,N_6338);
nor U8980 (N_8980,N_5117,N_5590);
and U8981 (N_8981,N_5013,N_5292);
xor U8982 (N_8982,N_6625,N_5392);
nor U8983 (N_8983,N_6563,N_7063);
nand U8984 (N_8984,N_5163,N_7284);
nor U8985 (N_8985,N_5820,N_5983);
nand U8986 (N_8986,N_5196,N_5453);
and U8987 (N_8987,N_6407,N_5792);
or U8988 (N_8988,N_5008,N_6361);
nand U8989 (N_8989,N_7130,N_7077);
nand U8990 (N_8990,N_7087,N_6749);
and U8991 (N_8991,N_5338,N_5251);
nor U8992 (N_8992,N_5067,N_7131);
or U8993 (N_8993,N_5973,N_6707);
nand U8994 (N_8994,N_6108,N_6744);
nor U8995 (N_8995,N_5348,N_7286);
nand U8996 (N_8996,N_5894,N_5715);
and U8997 (N_8997,N_6130,N_6902);
or U8998 (N_8998,N_7051,N_6967);
nor U8999 (N_8999,N_6314,N_5463);
nor U9000 (N_9000,N_5599,N_5238);
nor U9001 (N_9001,N_5157,N_6201);
xnor U9002 (N_9002,N_5021,N_6209);
xor U9003 (N_9003,N_5719,N_7475);
nor U9004 (N_9004,N_6416,N_7141);
and U9005 (N_9005,N_6072,N_5375);
nand U9006 (N_9006,N_5964,N_6221);
nand U9007 (N_9007,N_6334,N_7055);
and U9008 (N_9008,N_6653,N_6527);
or U9009 (N_9009,N_6451,N_5525);
or U9010 (N_9010,N_5059,N_6118);
and U9011 (N_9011,N_6717,N_7328);
and U9012 (N_9012,N_5001,N_5077);
and U9013 (N_9013,N_5862,N_6011);
and U9014 (N_9014,N_6525,N_6466);
nand U9015 (N_9015,N_6480,N_6339);
nand U9016 (N_9016,N_7246,N_5970);
nand U9017 (N_9017,N_5798,N_7285);
nand U9018 (N_9018,N_7037,N_5881);
and U9019 (N_9019,N_5520,N_6349);
or U9020 (N_9020,N_5415,N_6402);
and U9021 (N_9021,N_5713,N_6829);
and U9022 (N_9022,N_5876,N_5171);
and U9023 (N_9023,N_5890,N_6150);
nand U9024 (N_9024,N_7393,N_7472);
nor U9025 (N_9025,N_5489,N_5569);
nand U9026 (N_9026,N_5028,N_5606);
xor U9027 (N_9027,N_5157,N_6489);
and U9028 (N_9028,N_6600,N_5100);
nor U9029 (N_9029,N_6492,N_7322);
and U9030 (N_9030,N_5321,N_5156);
and U9031 (N_9031,N_6974,N_6289);
and U9032 (N_9032,N_5200,N_5605);
nand U9033 (N_9033,N_5741,N_5543);
nand U9034 (N_9034,N_7245,N_6907);
and U9035 (N_9035,N_5132,N_5759);
or U9036 (N_9036,N_5370,N_5358);
and U9037 (N_9037,N_5942,N_7281);
or U9038 (N_9038,N_5057,N_7271);
or U9039 (N_9039,N_6741,N_6429);
and U9040 (N_9040,N_5357,N_6022);
or U9041 (N_9041,N_5346,N_6352);
or U9042 (N_9042,N_6809,N_5688);
or U9043 (N_9043,N_5128,N_5501);
or U9044 (N_9044,N_6640,N_6046);
and U9045 (N_9045,N_7274,N_5879);
xnor U9046 (N_9046,N_7146,N_6546);
or U9047 (N_9047,N_7428,N_6659);
nor U9048 (N_9048,N_6563,N_6729);
nand U9049 (N_9049,N_5033,N_7000);
nand U9050 (N_9050,N_5103,N_7281);
nor U9051 (N_9051,N_5115,N_5375);
nand U9052 (N_9052,N_6001,N_6389);
nand U9053 (N_9053,N_6979,N_7448);
nand U9054 (N_9054,N_6299,N_6846);
nor U9055 (N_9055,N_7162,N_5153);
and U9056 (N_9056,N_6490,N_5527);
or U9057 (N_9057,N_6597,N_6150);
or U9058 (N_9058,N_7328,N_5245);
nand U9059 (N_9059,N_6108,N_5390);
nand U9060 (N_9060,N_5177,N_5434);
nor U9061 (N_9061,N_5191,N_6374);
or U9062 (N_9062,N_5831,N_6497);
nand U9063 (N_9063,N_6394,N_6639);
nand U9064 (N_9064,N_6060,N_7021);
and U9065 (N_9065,N_5795,N_5995);
nand U9066 (N_9066,N_7268,N_5906);
or U9067 (N_9067,N_5002,N_5684);
and U9068 (N_9068,N_6429,N_5849);
nand U9069 (N_9069,N_7160,N_7422);
and U9070 (N_9070,N_6826,N_7302);
nor U9071 (N_9071,N_6947,N_5502);
or U9072 (N_9072,N_6612,N_7126);
and U9073 (N_9073,N_5958,N_5115);
or U9074 (N_9074,N_6103,N_6160);
nand U9075 (N_9075,N_6263,N_6620);
or U9076 (N_9076,N_7065,N_6590);
and U9077 (N_9077,N_7037,N_7158);
and U9078 (N_9078,N_5392,N_5882);
nor U9079 (N_9079,N_5899,N_5931);
nand U9080 (N_9080,N_5894,N_6583);
nor U9081 (N_9081,N_5960,N_6181);
or U9082 (N_9082,N_6034,N_6036);
nor U9083 (N_9083,N_7440,N_7211);
nor U9084 (N_9084,N_7256,N_6256);
nand U9085 (N_9085,N_6182,N_6157);
and U9086 (N_9086,N_5115,N_7137);
or U9087 (N_9087,N_5169,N_5549);
and U9088 (N_9088,N_5399,N_6453);
nor U9089 (N_9089,N_6992,N_5688);
and U9090 (N_9090,N_5125,N_5015);
nor U9091 (N_9091,N_6667,N_5837);
or U9092 (N_9092,N_5240,N_5152);
and U9093 (N_9093,N_7262,N_5986);
and U9094 (N_9094,N_5696,N_6769);
or U9095 (N_9095,N_7390,N_6079);
nand U9096 (N_9096,N_7289,N_5333);
nand U9097 (N_9097,N_7436,N_5455);
or U9098 (N_9098,N_7466,N_6585);
and U9099 (N_9099,N_5181,N_5727);
or U9100 (N_9100,N_6950,N_5178);
or U9101 (N_9101,N_6352,N_7269);
nor U9102 (N_9102,N_5682,N_7251);
and U9103 (N_9103,N_5706,N_6190);
or U9104 (N_9104,N_6768,N_6058);
nand U9105 (N_9105,N_6346,N_6243);
or U9106 (N_9106,N_5305,N_5098);
or U9107 (N_9107,N_6479,N_7464);
or U9108 (N_9108,N_5880,N_7167);
nand U9109 (N_9109,N_6952,N_7426);
nor U9110 (N_9110,N_5190,N_5947);
nor U9111 (N_9111,N_7387,N_6073);
or U9112 (N_9112,N_6153,N_7251);
nand U9113 (N_9113,N_5903,N_5384);
nand U9114 (N_9114,N_6975,N_6452);
and U9115 (N_9115,N_6211,N_6475);
nor U9116 (N_9116,N_6377,N_6460);
and U9117 (N_9117,N_6927,N_6597);
nor U9118 (N_9118,N_7222,N_6735);
or U9119 (N_9119,N_5063,N_5917);
or U9120 (N_9120,N_6323,N_6788);
and U9121 (N_9121,N_7105,N_6430);
nand U9122 (N_9122,N_5586,N_6718);
nor U9123 (N_9123,N_6076,N_5427);
nor U9124 (N_9124,N_7104,N_6219);
or U9125 (N_9125,N_7465,N_5857);
nor U9126 (N_9126,N_7407,N_5319);
or U9127 (N_9127,N_6131,N_5886);
and U9128 (N_9128,N_7180,N_5314);
nor U9129 (N_9129,N_5034,N_6123);
and U9130 (N_9130,N_5171,N_7327);
nand U9131 (N_9131,N_5026,N_6602);
or U9132 (N_9132,N_5434,N_6285);
nand U9133 (N_9133,N_5580,N_6359);
and U9134 (N_9134,N_7466,N_7266);
nand U9135 (N_9135,N_6741,N_6716);
nand U9136 (N_9136,N_5468,N_6673);
and U9137 (N_9137,N_7441,N_6142);
nand U9138 (N_9138,N_5551,N_6528);
and U9139 (N_9139,N_6783,N_5151);
xor U9140 (N_9140,N_6450,N_6321);
or U9141 (N_9141,N_6326,N_7473);
and U9142 (N_9142,N_6842,N_5670);
nand U9143 (N_9143,N_5933,N_7077);
or U9144 (N_9144,N_5137,N_6985);
or U9145 (N_9145,N_6033,N_6794);
nand U9146 (N_9146,N_6707,N_5580);
or U9147 (N_9147,N_5379,N_6588);
nand U9148 (N_9148,N_7426,N_6053);
and U9149 (N_9149,N_7179,N_5842);
nor U9150 (N_9150,N_5787,N_7061);
nand U9151 (N_9151,N_6572,N_7126);
or U9152 (N_9152,N_7492,N_5832);
nor U9153 (N_9153,N_5251,N_5295);
or U9154 (N_9154,N_6544,N_6942);
and U9155 (N_9155,N_5247,N_5861);
and U9156 (N_9156,N_5276,N_6645);
nand U9157 (N_9157,N_6548,N_5855);
nand U9158 (N_9158,N_6245,N_7314);
nand U9159 (N_9159,N_5832,N_7131);
nand U9160 (N_9160,N_5785,N_7038);
or U9161 (N_9161,N_7371,N_7329);
nand U9162 (N_9162,N_5044,N_6650);
nor U9163 (N_9163,N_5176,N_6835);
nor U9164 (N_9164,N_6904,N_6427);
and U9165 (N_9165,N_5401,N_5202);
and U9166 (N_9166,N_5189,N_7412);
or U9167 (N_9167,N_5199,N_7265);
and U9168 (N_9168,N_6241,N_5628);
and U9169 (N_9169,N_6110,N_5332);
or U9170 (N_9170,N_5954,N_6866);
nand U9171 (N_9171,N_5580,N_5963);
or U9172 (N_9172,N_7428,N_7496);
or U9173 (N_9173,N_5102,N_5701);
nor U9174 (N_9174,N_6587,N_6406);
nor U9175 (N_9175,N_5838,N_6554);
or U9176 (N_9176,N_5157,N_7064);
and U9177 (N_9177,N_5170,N_7263);
nor U9178 (N_9178,N_5112,N_6773);
nand U9179 (N_9179,N_6657,N_5355);
and U9180 (N_9180,N_6049,N_6584);
or U9181 (N_9181,N_5243,N_5629);
nand U9182 (N_9182,N_6671,N_5942);
nand U9183 (N_9183,N_5413,N_5606);
and U9184 (N_9184,N_5744,N_6917);
or U9185 (N_9185,N_5329,N_6685);
or U9186 (N_9186,N_5068,N_7350);
or U9187 (N_9187,N_6493,N_5890);
xnor U9188 (N_9188,N_6211,N_5377);
nor U9189 (N_9189,N_6258,N_7184);
nand U9190 (N_9190,N_7175,N_5723);
nand U9191 (N_9191,N_5953,N_6802);
nand U9192 (N_9192,N_6582,N_6901);
and U9193 (N_9193,N_6186,N_5972);
nand U9194 (N_9194,N_6919,N_5515);
and U9195 (N_9195,N_5274,N_7339);
nor U9196 (N_9196,N_7158,N_6342);
nor U9197 (N_9197,N_6699,N_7098);
nand U9198 (N_9198,N_6450,N_6782);
nand U9199 (N_9199,N_6855,N_5379);
nand U9200 (N_9200,N_5018,N_6741);
nor U9201 (N_9201,N_6211,N_5872);
nand U9202 (N_9202,N_7121,N_5249);
or U9203 (N_9203,N_7432,N_7170);
or U9204 (N_9204,N_5484,N_6227);
nor U9205 (N_9205,N_6715,N_6402);
and U9206 (N_9206,N_7443,N_5430);
nand U9207 (N_9207,N_5243,N_5214);
and U9208 (N_9208,N_6225,N_5355);
and U9209 (N_9209,N_7034,N_5101);
xnor U9210 (N_9210,N_6468,N_5971);
and U9211 (N_9211,N_5380,N_6448);
or U9212 (N_9212,N_6419,N_7105);
or U9213 (N_9213,N_6414,N_6776);
and U9214 (N_9214,N_5220,N_5603);
nand U9215 (N_9215,N_5741,N_7149);
and U9216 (N_9216,N_6412,N_5728);
or U9217 (N_9217,N_5115,N_5882);
nor U9218 (N_9218,N_5061,N_7281);
nor U9219 (N_9219,N_5102,N_6652);
or U9220 (N_9220,N_5095,N_6585);
nand U9221 (N_9221,N_6405,N_7182);
nand U9222 (N_9222,N_5585,N_6240);
nand U9223 (N_9223,N_6773,N_5965);
and U9224 (N_9224,N_6678,N_5312);
or U9225 (N_9225,N_7287,N_6764);
nor U9226 (N_9226,N_6807,N_5481);
and U9227 (N_9227,N_7335,N_5557);
and U9228 (N_9228,N_5694,N_7450);
nand U9229 (N_9229,N_5247,N_6340);
or U9230 (N_9230,N_5428,N_5210);
nand U9231 (N_9231,N_7001,N_5283);
nand U9232 (N_9232,N_7234,N_5648);
and U9233 (N_9233,N_5890,N_5305);
and U9234 (N_9234,N_6676,N_6492);
xor U9235 (N_9235,N_6851,N_5417);
nand U9236 (N_9236,N_6690,N_7150);
xor U9237 (N_9237,N_5905,N_5289);
or U9238 (N_9238,N_7365,N_7406);
nand U9239 (N_9239,N_5468,N_6185);
nor U9240 (N_9240,N_5496,N_6648);
and U9241 (N_9241,N_5861,N_6212);
and U9242 (N_9242,N_6375,N_6028);
nand U9243 (N_9243,N_6128,N_5973);
or U9244 (N_9244,N_6202,N_6514);
nand U9245 (N_9245,N_5041,N_6538);
nand U9246 (N_9246,N_7043,N_5939);
nand U9247 (N_9247,N_5606,N_5398);
and U9248 (N_9248,N_5873,N_6189);
and U9249 (N_9249,N_6115,N_6135);
nor U9250 (N_9250,N_5400,N_5159);
and U9251 (N_9251,N_6349,N_7116);
nand U9252 (N_9252,N_7008,N_7205);
and U9253 (N_9253,N_6858,N_5932);
and U9254 (N_9254,N_6316,N_6081);
or U9255 (N_9255,N_5522,N_5666);
and U9256 (N_9256,N_6103,N_7090);
nor U9257 (N_9257,N_6720,N_7414);
nand U9258 (N_9258,N_6602,N_7231);
nor U9259 (N_9259,N_6981,N_7025);
nand U9260 (N_9260,N_6896,N_6315);
or U9261 (N_9261,N_6337,N_6657);
or U9262 (N_9262,N_5288,N_7245);
nor U9263 (N_9263,N_5097,N_6165);
and U9264 (N_9264,N_5745,N_7190);
nor U9265 (N_9265,N_5896,N_6064);
nor U9266 (N_9266,N_7408,N_6845);
or U9267 (N_9267,N_7023,N_7448);
nor U9268 (N_9268,N_6060,N_6947);
nand U9269 (N_9269,N_5272,N_5923);
nor U9270 (N_9270,N_6507,N_5782);
nand U9271 (N_9271,N_6813,N_7465);
or U9272 (N_9272,N_7182,N_6309);
nor U9273 (N_9273,N_7324,N_6591);
and U9274 (N_9274,N_5305,N_6575);
and U9275 (N_9275,N_5571,N_6400);
nor U9276 (N_9276,N_5406,N_5420);
and U9277 (N_9277,N_5634,N_5984);
nor U9278 (N_9278,N_6038,N_6843);
nand U9279 (N_9279,N_5409,N_6459);
nand U9280 (N_9280,N_5501,N_6981);
nor U9281 (N_9281,N_5160,N_7218);
nand U9282 (N_9282,N_6574,N_6185);
nor U9283 (N_9283,N_6036,N_6148);
and U9284 (N_9284,N_6339,N_6508);
or U9285 (N_9285,N_5918,N_6459);
or U9286 (N_9286,N_6913,N_6995);
and U9287 (N_9287,N_6763,N_5901);
or U9288 (N_9288,N_7234,N_6906);
nand U9289 (N_9289,N_5078,N_5153);
and U9290 (N_9290,N_5598,N_5031);
and U9291 (N_9291,N_5577,N_6646);
and U9292 (N_9292,N_5758,N_6715);
nand U9293 (N_9293,N_6713,N_6746);
nor U9294 (N_9294,N_5710,N_5664);
nand U9295 (N_9295,N_5214,N_6125);
xor U9296 (N_9296,N_6278,N_5374);
or U9297 (N_9297,N_5213,N_7477);
or U9298 (N_9298,N_5450,N_5407);
xor U9299 (N_9299,N_7110,N_5135);
nor U9300 (N_9300,N_5029,N_7178);
or U9301 (N_9301,N_6193,N_6964);
xnor U9302 (N_9302,N_6249,N_7354);
nor U9303 (N_9303,N_6403,N_7083);
and U9304 (N_9304,N_6822,N_7083);
and U9305 (N_9305,N_7180,N_7303);
nand U9306 (N_9306,N_5114,N_6368);
xnor U9307 (N_9307,N_7124,N_7237);
nor U9308 (N_9308,N_5207,N_6750);
or U9309 (N_9309,N_7130,N_7414);
nand U9310 (N_9310,N_5863,N_5696);
and U9311 (N_9311,N_7121,N_5282);
nor U9312 (N_9312,N_6156,N_7166);
nor U9313 (N_9313,N_5788,N_6496);
nor U9314 (N_9314,N_7482,N_6138);
or U9315 (N_9315,N_5613,N_6559);
and U9316 (N_9316,N_5005,N_6960);
or U9317 (N_9317,N_7231,N_5662);
xnor U9318 (N_9318,N_6486,N_6123);
or U9319 (N_9319,N_6665,N_5607);
and U9320 (N_9320,N_5800,N_5397);
nor U9321 (N_9321,N_7049,N_6511);
or U9322 (N_9322,N_5205,N_6661);
or U9323 (N_9323,N_7152,N_7113);
nand U9324 (N_9324,N_7298,N_6255);
nor U9325 (N_9325,N_7256,N_7041);
nand U9326 (N_9326,N_6878,N_6100);
nor U9327 (N_9327,N_6820,N_6997);
nor U9328 (N_9328,N_6144,N_5961);
nor U9329 (N_9329,N_7436,N_5728);
or U9330 (N_9330,N_5374,N_7373);
nor U9331 (N_9331,N_6582,N_5874);
nand U9332 (N_9332,N_5789,N_7442);
or U9333 (N_9333,N_5780,N_5054);
nor U9334 (N_9334,N_6072,N_6647);
xnor U9335 (N_9335,N_5003,N_6506);
nand U9336 (N_9336,N_5574,N_5887);
or U9337 (N_9337,N_5309,N_6013);
nor U9338 (N_9338,N_5061,N_6095);
nand U9339 (N_9339,N_7065,N_5425);
and U9340 (N_9340,N_6343,N_6717);
nand U9341 (N_9341,N_6108,N_5885);
or U9342 (N_9342,N_5072,N_6089);
nand U9343 (N_9343,N_5315,N_6571);
nor U9344 (N_9344,N_5007,N_7011);
nor U9345 (N_9345,N_6389,N_5799);
nand U9346 (N_9346,N_7174,N_7128);
or U9347 (N_9347,N_6409,N_5437);
and U9348 (N_9348,N_7490,N_6769);
nand U9349 (N_9349,N_5627,N_5913);
nand U9350 (N_9350,N_6620,N_5205);
nand U9351 (N_9351,N_7232,N_6112);
nor U9352 (N_9352,N_5345,N_7327);
nand U9353 (N_9353,N_6599,N_6359);
and U9354 (N_9354,N_5402,N_6605);
nor U9355 (N_9355,N_5176,N_7436);
or U9356 (N_9356,N_6540,N_5469);
nand U9357 (N_9357,N_6203,N_6575);
or U9358 (N_9358,N_7129,N_5961);
or U9359 (N_9359,N_5083,N_6205);
and U9360 (N_9360,N_5907,N_6471);
nand U9361 (N_9361,N_5286,N_6698);
nor U9362 (N_9362,N_6298,N_6005);
nor U9363 (N_9363,N_6598,N_6501);
or U9364 (N_9364,N_5558,N_5940);
nand U9365 (N_9365,N_6062,N_7006);
or U9366 (N_9366,N_5332,N_6513);
nor U9367 (N_9367,N_6038,N_5772);
nand U9368 (N_9368,N_5648,N_5862);
nor U9369 (N_9369,N_5184,N_5651);
nor U9370 (N_9370,N_5563,N_5565);
or U9371 (N_9371,N_5562,N_6843);
nor U9372 (N_9372,N_5986,N_6478);
nand U9373 (N_9373,N_5204,N_6528);
and U9374 (N_9374,N_5037,N_5610);
nor U9375 (N_9375,N_5080,N_5124);
or U9376 (N_9376,N_5571,N_6939);
nand U9377 (N_9377,N_7225,N_7421);
nand U9378 (N_9378,N_7334,N_5549);
nand U9379 (N_9379,N_5638,N_6667);
nand U9380 (N_9380,N_6296,N_6366);
nor U9381 (N_9381,N_5501,N_5161);
or U9382 (N_9382,N_5737,N_5459);
nor U9383 (N_9383,N_7458,N_5793);
nand U9384 (N_9384,N_6533,N_6351);
or U9385 (N_9385,N_6101,N_7184);
and U9386 (N_9386,N_6147,N_6945);
nor U9387 (N_9387,N_5976,N_5885);
nor U9388 (N_9388,N_5130,N_5782);
or U9389 (N_9389,N_7249,N_7263);
nor U9390 (N_9390,N_7132,N_5708);
nand U9391 (N_9391,N_6516,N_6684);
nor U9392 (N_9392,N_5807,N_6461);
and U9393 (N_9393,N_6613,N_5400);
nand U9394 (N_9394,N_6036,N_5580);
or U9395 (N_9395,N_6543,N_5109);
and U9396 (N_9396,N_6934,N_5466);
nand U9397 (N_9397,N_6977,N_6446);
and U9398 (N_9398,N_7053,N_6206);
and U9399 (N_9399,N_6365,N_7213);
or U9400 (N_9400,N_6157,N_7249);
nand U9401 (N_9401,N_6748,N_6680);
nand U9402 (N_9402,N_5536,N_7350);
nor U9403 (N_9403,N_5014,N_6819);
nand U9404 (N_9404,N_5673,N_5715);
nor U9405 (N_9405,N_5207,N_5121);
or U9406 (N_9406,N_7496,N_7042);
or U9407 (N_9407,N_6054,N_6604);
and U9408 (N_9408,N_6865,N_5037);
or U9409 (N_9409,N_6560,N_5205);
xor U9410 (N_9410,N_6615,N_5976);
and U9411 (N_9411,N_6321,N_7143);
and U9412 (N_9412,N_5543,N_5463);
and U9413 (N_9413,N_6409,N_6879);
nand U9414 (N_9414,N_6030,N_6204);
and U9415 (N_9415,N_6400,N_6804);
nor U9416 (N_9416,N_7022,N_7261);
or U9417 (N_9417,N_6843,N_5584);
or U9418 (N_9418,N_7156,N_5838);
and U9419 (N_9419,N_6171,N_6968);
nand U9420 (N_9420,N_5992,N_5283);
and U9421 (N_9421,N_5401,N_5374);
nand U9422 (N_9422,N_6307,N_6162);
nand U9423 (N_9423,N_6089,N_6623);
nor U9424 (N_9424,N_6693,N_6337);
nand U9425 (N_9425,N_6181,N_5400);
or U9426 (N_9426,N_6193,N_6055);
and U9427 (N_9427,N_6089,N_5924);
or U9428 (N_9428,N_5611,N_5292);
nand U9429 (N_9429,N_5407,N_6998);
or U9430 (N_9430,N_6065,N_6040);
or U9431 (N_9431,N_7467,N_6115);
nand U9432 (N_9432,N_5141,N_5183);
nor U9433 (N_9433,N_6211,N_5623);
nor U9434 (N_9434,N_5519,N_6839);
or U9435 (N_9435,N_5994,N_6382);
nor U9436 (N_9436,N_6874,N_5485);
nor U9437 (N_9437,N_5899,N_6949);
or U9438 (N_9438,N_5298,N_5717);
or U9439 (N_9439,N_7225,N_6149);
nand U9440 (N_9440,N_5813,N_5390);
nor U9441 (N_9441,N_5894,N_6312);
xnor U9442 (N_9442,N_6726,N_7255);
or U9443 (N_9443,N_5607,N_7385);
nand U9444 (N_9444,N_6837,N_6669);
and U9445 (N_9445,N_5210,N_6372);
nand U9446 (N_9446,N_5167,N_5618);
nand U9447 (N_9447,N_5392,N_6996);
nor U9448 (N_9448,N_7208,N_5260);
and U9449 (N_9449,N_6802,N_6248);
or U9450 (N_9450,N_7384,N_5538);
or U9451 (N_9451,N_5593,N_6345);
and U9452 (N_9452,N_6714,N_6799);
nor U9453 (N_9453,N_6170,N_5650);
nor U9454 (N_9454,N_5631,N_7312);
nand U9455 (N_9455,N_6893,N_6913);
nor U9456 (N_9456,N_6844,N_6522);
nand U9457 (N_9457,N_6438,N_6815);
nor U9458 (N_9458,N_5293,N_5913);
nor U9459 (N_9459,N_6585,N_6557);
nand U9460 (N_9460,N_6438,N_6782);
nand U9461 (N_9461,N_7363,N_6130);
nor U9462 (N_9462,N_5658,N_5868);
nor U9463 (N_9463,N_5656,N_6423);
or U9464 (N_9464,N_5095,N_6561);
and U9465 (N_9465,N_5149,N_5892);
and U9466 (N_9466,N_5599,N_5113);
and U9467 (N_9467,N_5892,N_7417);
nand U9468 (N_9468,N_6129,N_5643);
nor U9469 (N_9469,N_6688,N_5576);
nand U9470 (N_9470,N_6761,N_7008);
or U9471 (N_9471,N_7196,N_5986);
nor U9472 (N_9472,N_5248,N_5330);
nand U9473 (N_9473,N_6108,N_5416);
nand U9474 (N_9474,N_6886,N_5850);
or U9475 (N_9475,N_6016,N_5896);
and U9476 (N_9476,N_7468,N_5204);
and U9477 (N_9477,N_6703,N_5667);
xor U9478 (N_9478,N_5568,N_6751);
or U9479 (N_9479,N_5055,N_7238);
nor U9480 (N_9480,N_6483,N_5995);
or U9481 (N_9481,N_5648,N_7135);
xnor U9482 (N_9482,N_5296,N_6558);
nand U9483 (N_9483,N_7254,N_6362);
nand U9484 (N_9484,N_5154,N_7369);
nand U9485 (N_9485,N_7119,N_6329);
nand U9486 (N_9486,N_7349,N_5914);
nand U9487 (N_9487,N_5386,N_6871);
nor U9488 (N_9488,N_6534,N_6885);
or U9489 (N_9489,N_6478,N_6861);
or U9490 (N_9490,N_5200,N_6487);
nand U9491 (N_9491,N_6164,N_7208);
and U9492 (N_9492,N_6997,N_5232);
nor U9493 (N_9493,N_5033,N_6651);
or U9494 (N_9494,N_6362,N_6730);
and U9495 (N_9495,N_5566,N_5122);
nor U9496 (N_9496,N_5446,N_5902);
nand U9497 (N_9497,N_6446,N_6935);
and U9498 (N_9498,N_6405,N_5302);
or U9499 (N_9499,N_6047,N_6841);
or U9500 (N_9500,N_7139,N_7433);
and U9501 (N_9501,N_6723,N_5759);
or U9502 (N_9502,N_5696,N_6836);
or U9503 (N_9503,N_6193,N_7434);
nand U9504 (N_9504,N_7427,N_7119);
nor U9505 (N_9505,N_6082,N_6323);
or U9506 (N_9506,N_6257,N_5079);
and U9507 (N_9507,N_7100,N_7241);
xor U9508 (N_9508,N_5006,N_6931);
nand U9509 (N_9509,N_6141,N_7023);
nand U9510 (N_9510,N_7075,N_5633);
and U9511 (N_9511,N_6421,N_6712);
nand U9512 (N_9512,N_6432,N_6019);
nand U9513 (N_9513,N_6042,N_5439);
or U9514 (N_9514,N_6388,N_6862);
nand U9515 (N_9515,N_5938,N_5321);
nand U9516 (N_9516,N_7095,N_7090);
nand U9517 (N_9517,N_7076,N_5521);
nor U9518 (N_9518,N_5361,N_7100);
or U9519 (N_9519,N_5826,N_5230);
and U9520 (N_9520,N_7170,N_5202);
or U9521 (N_9521,N_5250,N_5199);
and U9522 (N_9522,N_5598,N_6663);
or U9523 (N_9523,N_7271,N_5328);
and U9524 (N_9524,N_6308,N_5937);
and U9525 (N_9525,N_6293,N_6472);
and U9526 (N_9526,N_7109,N_7031);
or U9527 (N_9527,N_5871,N_7210);
nor U9528 (N_9528,N_5387,N_6947);
nor U9529 (N_9529,N_5634,N_6815);
nand U9530 (N_9530,N_7427,N_5510);
nor U9531 (N_9531,N_6943,N_6631);
nor U9532 (N_9532,N_5044,N_6387);
nor U9533 (N_9533,N_5871,N_5437);
or U9534 (N_9534,N_5625,N_7099);
nor U9535 (N_9535,N_5650,N_6968);
nor U9536 (N_9536,N_6281,N_6487);
nor U9537 (N_9537,N_6944,N_5582);
or U9538 (N_9538,N_6572,N_6913);
or U9539 (N_9539,N_5938,N_5705);
nor U9540 (N_9540,N_7345,N_5573);
nor U9541 (N_9541,N_5936,N_5565);
nor U9542 (N_9542,N_6682,N_6000);
nor U9543 (N_9543,N_5760,N_6846);
nand U9544 (N_9544,N_5523,N_7460);
and U9545 (N_9545,N_5032,N_6401);
nor U9546 (N_9546,N_7233,N_5269);
or U9547 (N_9547,N_5027,N_6488);
nand U9548 (N_9548,N_6261,N_7341);
nand U9549 (N_9549,N_5311,N_6712);
nor U9550 (N_9550,N_6672,N_5358);
and U9551 (N_9551,N_5084,N_6384);
xnor U9552 (N_9552,N_6191,N_6366);
nand U9553 (N_9553,N_5551,N_6769);
or U9554 (N_9554,N_5924,N_7488);
nor U9555 (N_9555,N_5244,N_5755);
or U9556 (N_9556,N_7073,N_5148);
or U9557 (N_9557,N_6393,N_6852);
nand U9558 (N_9558,N_5534,N_6595);
or U9559 (N_9559,N_5125,N_6431);
nand U9560 (N_9560,N_6465,N_6322);
or U9561 (N_9561,N_7144,N_6770);
nor U9562 (N_9562,N_5953,N_5613);
nor U9563 (N_9563,N_5924,N_7325);
nand U9564 (N_9564,N_6622,N_5337);
and U9565 (N_9565,N_6811,N_6368);
or U9566 (N_9566,N_6858,N_6365);
or U9567 (N_9567,N_6893,N_6798);
or U9568 (N_9568,N_6261,N_6321);
and U9569 (N_9569,N_5686,N_5543);
nand U9570 (N_9570,N_7233,N_6793);
nand U9571 (N_9571,N_5329,N_6809);
xnor U9572 (N_9572,N_5971,N_5775);
nand U9573 (N_9573,N_5749,N_6603);
and U9574 (N_9574,N_7232,N_5161);
nor U9575 (N_9575,N_5247,N_5046);
or U9576 (N_9576,N_5378,N_6657);
and U9577 (N_9577,N_7445,N_7116);
and U9578 (N_9578,N_7410,N_7083);
and U9579 (N_9579,N_5677,N_5895);
or U9580 (N_9580,N_6663,N_5332);
nand U9581 (N_9581,N_6154,N_5169);
nor U9582 (N_9582,N_6519,N_5879);
or U9583 (N_9583,N_6208,N_6897);
or U9584 (N_9584,N_7340,N_6343);
or U9585 (N_9585,N_6719,N_6861);
or U9586 (N_9586,N_7157,N_7273);
xor U9587 (N_9587,N_7127,N_6998);
nor U9588 (N_9588,N_7003,N_5696);
and U9589 (N_9589,N_6986,N_7342);
nor U9590 (N_9590,N_6685,N_6134);
nand U9591 (N_9591,N_6269,N_5422);
xor U9592 (N_9592,N_6439,N_7159);
nor U9593 (N_9593,N_7011,N_5921);
xor U9594 (N_9594,N_6483,N_5738);
or U9595 (N_9595,N_6509,N_5397);
nor U9596 (N_9596,N_6415,N_7027);
or U9597 (N_9597,N_6936,N_6016);
and U9598 (N_9598,N_5303,N_6920);
nand U9599 (N_9599,N_5471,N_6917);
nand U9600 (N_9600,N_5640,N_6722);
and U9601 (N_9601,N_7129,N_5272);
xnor U9602 (N_9602,N_5978,N_6861);
nor U9603 (N_9603,N_5674,N_7264);
and U9604 (N_9604,N_5260,N_6948);
nor U9605 (N_9605,N_5000,N_5673);
nor U9606 (N_9606,N_6250,N_6835);
nand U9607 (N_9607,N_5138,N_6093);
and U9608 (N_9608,N_6091,N_7456);
nand U9609 (N_9609,N_5362,N_6860);
nand U9610 (N_9610,N_5649,N_5127);
and U9611 (N_9611,N_7441,N_6584);
nor U9612 (N_9612,N_5878,N_6487);
or U9613 (N_9613,N_6106,N_5472);
xor U9614 (N_9614,N_6663,N_7414);
nand U9615 (N_9615,N_5688,N_7426);
and U9616 (N_9616,N_5927,N_5575);
nor U9617 (N_9617,N_5519,N_7093);
or U9618 (N_9618,N_7481,N_5814);
and U9619 (N_9619,N_7151,N_7099);
nand U9620 (N_9620,N_6422,N_5792);
nand U9621 (N_9621,N_7444,N_6776);
or U9622 (N_9622,N_5637,N_5560);
nand U9623 (N_9623,N_5654,N_7341);
and U9624 (N_9624,N_5233,N_5072);
nor U9625 (N_9625,N_7367,N_6432);
and U9626 (N_9626,N_5166,N_6560);
nand U9627 (N_9627,N_6589,N_5473);
xnor U9628 (N_9628,N_5190,N_6546);
nor U9629 (N_9629,N_5411,N_5965);
nor U9630 (N_9630,N_5696,N_5745);
and U9631 (N_9631,N_7423,N_5787);
nand U9632 (N_9632,N_7382,N_5898);
or U9633 (N_9633,N_6248,N_6700);
nand U9634 (N_9634,N_5776,N_5616);
or U9635 (N_9635,N_5330,N_6133);
and U9636 (N_9636,N_5582,N_7168);
and U9637 (N_9637,N_5254,N_6665);
or U9638 (N_9638,N_6463,N_5566);
nor U9639 (N_9639,N_6051,N_6806);
nand U9640 (N_9640,N_6902,N_6168);
nor U9641 (N_9641,N_6924,N_6190);
nor U9642 (N_9642,N_7368,N_7108);
nor U9643 (N_9643,N_7291,N_5103);
nor U9644 (N_9644,N_7480,N_5375);
nor U9645 (N_9645,N_7475,N_6170);
and U9646 (N_9646,N_5469,N_6543);
nand U9647 (N_9647,N_6853,N_7049);
nand U9648 (N_9648,N_7228,N_6995);
or U9649 (N_9649,N_7497,N_6233);
xnor U9650 (N_9650,N_6128,N_7204);
nor U9651 (N_9651,N_5674,N_7085);
and U9652 (N_9652,N_5773,N_6334);
nand U9653 (N_9653,N_6725,N_6770);
nand U9654 (N_9654,N_6276,N_5614);
nand U9655 (N_9655,N_7307,N_5856);
or U9656 (N_9656,N_5061,N_6712);
nand U9657 (N_9657,N_6601,N_6996);
and U9658 (N_9658,N_6309,N_7405);
nor U9659 (N_9659,N_6812,N_5993);
and U9660 (N_9660,N_6335,N_7471);
or U9661 (N_9661,N_5505,N_5464);
or U9662 (N_9662,N_7186,N_6969);
or U9663 (N_9663,N_6310,N_5737);
nand U9664 (N_9664,N_7482,N_5697);
nor U9665 (N_9665,N_7322,N_5397);
or U9666 (N_9666,N_5214,N_5876);
nor U9667 (N_9667,N_6143,N_6671);
xnor U9668 (N_9668,N_5978,N_7317);
and U9669 (N_9669,N_5312,N_6257);
or U9670 (N_9670,N_6207,N_7393);
nor U9671 (N_9671,N_5782,N_7446);
nor U9672 (N_9672,N_6073,N_5412);
and U9673 (N_9673,N_6332,N_7281);
nor U9674 (N_9674,N_5564,N_5292);
or U9675 (N_9675,N_5214,N_5317);
nor U9676 (N_9676,N_6074,N_6387);
nand U9677 (N_9677,N_6368,N_7131);
and U9678 (N_9678,N_6749,N_5760);
and U9679 (N_9679,N_7029,N_7277);
or U9680 (N_9680,N_6069,N_7043);
or U9681 (N_9681,N_6160,N_5671);
and U9682 (N_9682,N_7171,N_5988);
nor U9683 (N_9683,N_5730,N_5701);
and U9684 (N_9684,N_6415,N_5267);
nand U9685 (N_9685,N_5691,N_6352);
nand U9686 (N_9686,N_6227,N_5457);
nor U9687 (N_9687,N_5170,N_5720);
nand U9688 (N_9688,N_5551,N_5325);
nor U9689 (N_9689,N_5496,N_5429);
nand U9690 (N_9690,N_5734,N_6410);
nor U9691 (N_9691,N_6033,N_6514);
nand U9692 (N_9692,N_5484,N_5927);
nor U9693 (N_9693,N_5113,N_6998);
xnor U9694 (N_9694,N_6076,N_7157);
nand U9695 (N_9695,N_6285,N_6998);
nor U9696 (N_9696,N_6253,N_6855);
and U9697 (N_9697,N_5692,N_7096);
or U9698 (N_9698,N_5047,N_5817);
or U9699 (N_9699,N_7135,N_6412);
and U9700 (N_9700,N_5862,N_5216);
nand U9701 (N_9701,N_5015,N_7076);
and U9702 (N_9702,N_7020,N_6768);
xnor U9703 (N_9703,N_5266,N_5007);
xor U9704 (N_9704,N_6597,N_5462);
nor U9705 (N_9705,N_6875,N_5802);
nand U9706 (N_9706,N_7150,N_7230);
or U9707 (N_9707,N_6418,N_6856);
and U9708 (N_9708,N_6789,N_5873);
or U9709 (N_9709,N_5976,N_7072);
or U9710 (N_9710,N_7253,N_5730);
xor U9711 (N_9711,N_6233,N_5935);
or U9712 (N_9712,N_6417,N_5279);
nor U9713 (N_9713,N_6425,N_5826);
or U9714 (N_9714,N_7384,N_5055);
nand U9715 (N_9715,N_5200,N_5803);
nand U9716 (N_9716,N_7142,N_6815);
and U9717 (N_9717,N_6190,N_5108);
or U9718 (N_9718,N_7146,N_6455);
xor U9719 (N_9719,N_7308,N_7433);
and U9720 (N_9720,N_6298,N_6062);
nor U9721 (N_9721,N_5075,N_5917);
and U9722 (N_9722,N_6117,N_5414);
xnor U9723 (N_9723,N_6140,N_5417);
or U9724 (N_9724,N_5381,N_5074);
or U9725 (N_9725,N_6426,N_6805);
xor U9726 (N_9726,N_6809,N_6927);
xnor U9727 (N_9727,N_6993,N_7193);
nand U9728 (N_9728,N_6462,N_6772);
nand U9729 (N_9729,N_6424,N_6113);
and U9730 (N_9730,N_6749,N_5042);
nor U9731 (N_9731,N_6730,N_6789);
or U9732 (N_9732,N_6179,N_5701);
or U9733 (N_9733,N_5108,N_5953);
nand U9734 (N_9734,N_5819,N_6886);
and U9735 (N_9735,N_5895,N_7201);
nand U9736 (N_9736,N_7465,N_6068);
nand U9737 (N_9737,N_5867,N_5144);
and U9738 (N_9738,N_6933,N_7240);
nor U9739 (N_9739,N_7084,N_6733);
and U9740 (N_9740,N_5394,N_5027);
nand U9741 (N_9741,N_5115,N_6895);
nor U9742 (N_9742,N_7170,N_5417);
or U9743 (N_9743,N_6278,N_5771);
or U9744 (N_9744,N_5065,N_5452);
xor U9745 (N_9745,N_6685,N_5047);
or U9746 (N_9746,N_5587,N_6355);
or U9747 (N_9747,N_5004,N_6321);
or U9748 (N_9748,N_5429,N_6352);
nand U9749 (N_9749,N_5940,N_7150);
or U9750 (N_9750,N_6975,N_5825);
and U9751 (N_9751,N_5613,N_5831);
nand U9752 (N_9752,N_5380,N_6017);
xnor U9753 (N_9753,N_6006,N_6750);
nand U9754 (N_9754,N_5452,N_5074);
or U9755 (N_9755,N_6493,N_7363);
nand U9756 (N_9756,N_7463,N_6660);
nor U9757 (N_9757,N_6535,N_5409);
nand U9758 (N_9758,N_6927,N_6228);
nand U9759 (N_9759,N_7418,N_5705);
and U9760 (N_9760,N_7475,N_6773);
or U9761 (N_9761,N_5565,N_5808);
or U9762 (N_9762,N_5159,N_5860);
or U9763 (N_9763,N_5283,N_5036);
or U9764 (N_9764,N_5967,N_6270);
nor U9765 (N_9765,N_6916,N_7442);
or U9766 (N_9766,N_7252,N_7304);
nor U9767 (N_9767,N_6386,N_5237);
and U9768 (N_9768,N_5665,N_5078);
or U9769 (N_9769,N_6181,N_5961);
or U9770 (N_9770,N_5171,N_5413);
xnor U9771 (N_9771,N_7398,N_7137);
nand U9772 (N_9772,N_6517,N_6743);
nand U9773 (N_9773,N_6837,N_5550);
or U9774 (N_9774,N_5174,N_7300);
nand U9775 (N_9775,N_5304,N_7354);
nor U9776 (N_9776,N_7008,N_5849);
nand U9777 (N_9777,N_5810,N_6439);
and U9778 (N_9778,N_5438,N_6812);
or U9779 (N_9779,N_7177,N_6948);
nand U9780 (N_9780,N_6573,N_6478);
xnor U9781 (N_9781,N_6890,N_5167);
and U9782 (N_9782,N_7317,N_6992);
and U9783 (N_9783,N_6215,N_6307);
nor U9784 (N_9784,N_5200,N_5708);
nor U9785 (N_9785,N_6970,N_5111);
nand U9786 (N_9786,N_6803,N_6327);
or U9787 (N_9787,N_6133,N_6462);
or U9788 (N_9788,N_7178,N_5497);
or U9789 (N_9789,N_7437,N_6781);
or U9790 (N_9790,N_7495,N_6158);
nor U9791 (N_9791,N_5610,N_5395);
nor U9792 (N_9792,N_7234,N_5102);
nand U9793 (N_9793,N_5664,N_6216);
or U9794 (N_9794,N_7354,N_7273);
nor U9795 (N_9795,N_5478,N_5491);
nand U9796 (N_9796,N_6399,N_5035);
and U9797 (N_9797,N_7169,N_6191);
nor U9798 (N_9798,N_7176,N_5463);
nand U9799 (N_9799,N_5442,N_5282);
nor U9800 (N_9800,N_5399,N_7267);
nand U9801 (N_9801,N_6015,N_7061);
nand U9802 (N_9802,N_5604,N_5016);
nor U9803 (N_9803,N_7476,N_5758);
nor U9804 (N_9804,N_5905,N_6312);
and U9805 (N_9805,N_6908,N_5481);
or U9806 (N_9806,N_5147,N_6343);
xnor U9807 (N_9807,N_5611,N_5610);
nand U9808 (N_9808,N_6577,N_5509);
or U9809 (N_9809,N_6196,N_6864);
nand U9810 (N_9810,N_5798,N_7058);
nor U9811 (N_9811,N_6878,N_5545);
nor U9812 (N_9812,N_7134,N_6137);
nand U9813 (N_9813,N_7156,N_7180);
and U9814 (N_9814,N_5443,N_6766);
nand U9815 (N_9815,N_6041,N_7028);
nand U9816 (N_9816,N_7355,N_6403);
nand U9817 (N_9817,N_7481,N_5793);
or U9818 (N_9818,N_5685,N_6897);
nand U9819 (N_9819,N_6559,N_5755);
nand U9820 (N_9820,N_6046,N_6433);
and U9821 (N_9821,N_5618,N_5729);
nor U9822 (N_9822,N_7121,N_5235);
nor U9823 (N_9823,N_7464,N_7080);
nand U9824 (N_9824,N_5164,N_7336);
or U9825 (N_9825,N_7438,N_5328);
or U9826 (N_9826,N_6558,N_6553);
or U9827 (N_9827,N_5226,N_5143);
nor U9828 (N_9828,N_6932,N_6609);
and U9829 (N_9829,N_6353,N_7365);
or U9830 (N_9830,N_5783,N_5393);
nor U9831 (N_9831,N_7106,N_5167);
nand U9832 (N_9832,N_6877,N_5279);
xor U9833 (N_9833,N_6771,N_6981);
xor U9834 (N_9834,N_5199,N_5217);
or U9835 (N_9835,N_5110,N_5483);
or U9836 (N_9836,N_5220,N_5942);
or U9837 (N_9837,N_7396,N_6572);
or U9838 (N_9838,N_6367,N_5445);
xnor U9839 (N_9839,N_5086,N_5010);
nor U9840 (N_9840,N_5868,N_5543);
or U9841 (N_9841,N_5767,N_7025);
nor U9842 (N_9842,N_5304,N_6236);
nand U9843 (N_9843,N_6430,N_6222);
nand U9844 (N_9844,N_6677,N_6091);
and U9845 (N_9845,N_5283,N_6577);
or U9846 (N_9846,N_7419,N_7479);
nand U9847 (N_9847,N_6636,N_7124);
and U9848 (N_9848,N_5430,N_5010);
nor U9849 (N_9849,N_5355,N_6848);
or U9850 (N_9850,N_5535,N_6221);
nor U9851 (N_9851,N_7167,N_7414);
and U9852 (N_9852,N_7477,N_5915);
nor U9853 (N_9853,N_6585,N_7479);
nand U9854 (N_9854,N_7272,N_5166);
xnor U9855 (N_9855,N_5922,N_7083);
or U9856 (N_9856,N_7094,N_5214);
nor U9857 (N_9857,N_6363,N_6991);
nand U9858 (N_9858,N_6717,N_6888);
and U9859 (N_9859,N_6014,N_5342);
nor U9860 (N_9860,N_5519,N_6493);
nand U9861 (N_9861,N_7397,N_7037);
nor U9862 (N_9862,N_7131,N_5687);
and U9863 (N_9863,N_6476,N_7233);
and U9864 (N_9864,N_5837,N_6636);
nor U9865 (N_9865,N_5595,N_6280);
nand U9866 (N_9866,N_5337,N_7031);
or U9867 (N_9867,N_5811,N_5857);
nor U9868 (N_9868,N_6755,N_5552);
and U9869 (N_9869,N_6418,N_7052);
nor U9870 (N_9870,N_7275,N_6388);
xnor U9871 (N_9871,N_5461,N_6082);
nand U9872 (N_9872,N_6460,N_5425);
nor U9873 (N_9873,N_5493,N_5573);
or U9874 (N_9874,N_6558,N_7481);
and U9875 (N_9875,N_6967,N_7086);
and U9876 (N_9876,N_5529,N_6389);
and U9877 (N_9877,N_6076,N_6078);
nor U9878 (N_9878,N_6094,N_7279);
nand U9879 (N_9879,N_5250,N_5408);
or U9880 (N_9880,N_6774,N_5067);
xnor U9881 (N_9881,N_5257,N_5144);
or U9882 (N_9882,N_6163,N_5205);
or U9883 (N_9883,N_6106,N_6550);
and U9884 (N_9884,N_6050,N_5135);
nand U9885 (N_9885,N_7104,N_6054);
or U9886 (N_9886,N_6659,N_5468);
and U9887 (N_9887,N_7348,N_6662);
nand U9888 (N_9888,N_6101,N_5751);
nor U9889 (N_9889,N_7358,N_7407);
nand U9890 (N_9890,N_7389,N_7290);
nand U9891 (N_9891,N_6542,N_5736);
nand U9892 (N_9892,N_5050,N_5078);
nand U9893 (N_9893,N_6698,N_7205);
nor U9894 (N_9894,N_6951,N_5590);
xor U9895 (N_9895,N_5287,N_5370);
nand U9896 (N_9896,N_5643,N_5985);
or U9897 (N_9897,N_6145,N_5854);
nand U9898 (N_9898,N_6508,N_5295);
nand U9899 (N_9899,N_5917,N_5235);
and U9900 (N_9900,N_5401,N_5519);
or U9901 (N_9901,N_7310,N_5481);
or U9902 (N_9902,N_6240,N_6967);
nor U9903 (N_9903,N_5353,N_5843);
and U9904 (N_9904,N_5770,N_5521);
nand U9905 (N_9905,N_7005,N_5689);
or U9906 (N_9906,N_5116,N_5521);
or U9907 (N_9907,N_5715,N_7390);
or U9908 (N_9908,N_5011,N_7044);
and U9909 (N_9909,N_6645,N_7089);
or U9910 (N_9910,N_7379,N_6156);
or U9911 (N_9911,N_6324,N_5677);
and U9912 (N_9912,N_6695,N_6304);
nand U9913 (N_9913,N_5091,N_5420);
and U9914 (N_9914,N_7462,N_7082);
and U9915 (N_9915,N_7168,N_7446);
or U9916 (N_9916,N_7250,N_6872);
nand U9917 (N_9917,N_6636,N_7109);
nand U9918 (N_9918,N_5562,N_5775);
or U9919 (N_9919,N_5685,N_6774);
or U9920 (N_9920,N_7279,N_6553);
nor U9921 (N_9921,N_7164,N_5905);
or U9922 (N_9922,N_7488,N_6275);
nor U9923 (N_9923,N_6323,N_5876);
nand U9924 (N_9924,N_7151,N_6048);
or U9925 (N_9925,N_5332,N_6306);
nor U9926 (N_9926,N_5634,N_5565);
or U9927 (N_9927,N_6124,N_7445);
and U9928 (N_9928,N_5603,N_6091);
nand U9929 (N_9929,N_6743,N_6531);
nor U9930 (N_9930,N_7165,N_6667);
nor U9931 (N_9931,N_5887,N_5661);
nor U9932 (N_9932,N_5153,N_5590);
or U9933 (N_9933,N_7305,N_7298);
and U9934 (N_9934,N_6054,N_6359);
nor U9935 (N_9935,N_6265,N_7333);
or U9936 (N_9936,N_5284,N_5157);
and U9937 (N_9937,N_7043,N_6165);
nor U9938 (N_9938,N_7471,N_5192);
nor U9939 (N_9939,N_5928,N_5054);
nor U9940 (N_9940,N_5770,N_5234);
nand U9941 (N_9941,N_6656,N_5915);
and U9942 (N_9942,N_5440,N_5666);
or U9943 (N_9943,N_6780,N_6118);
or U9944 (N_9944,N_6326,N_5030);
nand U9945 (N_9945,N_6903,N_6460);
or U9946 (N_9946,N_7181,N_7148);
nand U9947 (N_9947,N_6334,N_5710);
or U9948 (N_9948,N_6413,N_5393);
nor U9949 (N_9949,N_6620,N_6888);
nor U9950 (N_9950,N_6049,N_5052);
or U9951 (N_9951,N_6757,N_7464);
nor U9952 (N_9952,N_6791,N_5357);
or U9953 (N_9953,N_5801,N_5434);
nor U9954 (N_9954,N_6933,N_6890);
and U9955 (N_9955,N_5210,N_6569);
nor U9956 (N_9956,N_5958,N_6122);
and U9957 (N_9957,N_6844,N_6712);
nor U9958 (N_9958,N_5751,N_6365);
or U9959 (N_9959,N_7498,N_6232);
or U9960 (N_9960,N_6423,N_7014);
or U9961 (N_9961,N_5329,N_5281);
and U9962 (N_9962,N_6775,N_6628);
nand U9963 (N_9963,N_6575,N_5421);
nor U9964 (N_9964,N_5862,N_7043);
nand U9965 (N_9965,N_5698,N_7156);
nor U9966 (N_9966,N_5293,N_6265);
nor U9967 (N_9967,N_6337,N_7188);
nor U9968 (N_9968,N_7035,N_6951);
and U9969 (N_9969,N_5125,N_6397);
and U9970 (N_9970,N_7358,N_6691);
or U9971 (N_9971,N_6672,N_6714);
nor U9972 (N_9972,N_5678,N_6085);
nor U9973 (N_9973,N_6445,N_5129);
nor U9974 (N_9974,N_6019,N_5698);
and U9975 (N_9975,N_5914,N_5970);
nand U9976 (N_9976,N_5930,N_5348);
nand U9977 (N_9977,N_6095,N_6816);
nor U9978 (N_9978,N_7461,N_7027);
nor U9979 (N_9979,N_7185,N_7012);
and U9980 (N_9980,N_5405,N_7461);
nor U9981 (N_9981,N_6937,N_6302);
and U9982 (N_9982,N_7026,N_5857);
nand U9983 (N_9983,N_6894,N_5528);
or U9984 (N_9984,N_5772,N_5948);
nand U9985 (N_9985,N_6170,N_6038);
nand U9986 (N_9986,N_7082,N_6912);
or U9987 (N_9987,N_6840,N_5118);
nor U9988 (N_9988,N_7406,N_5734);
nor U9989 (N_9989,N_6139,N_6826);
nand U9990 (N_9990,N_7118,N_6367);
or U9991 (N_9991,N_5275,N_5661);
and U9992 (N_9992,N_6427,N_5093);
or U9993 (N_9993,N_6638,N_5434);
nor U9994 (N_9994,N_5788,N_5365);
nor U9995 (N_9995,N_6352,N_6768);
and U9996 (N_9996,N_6346,N_5899);
and U9997 (N_9997,N_5820,N_6225);
nand U9998 (N_9998,N_6982,N_5427);
nor U9999 (N_9999,N_7407,N_5653);
nand UO_0 (O_0,N_9951,N_8291);
nand UO_1 (O_1,N_9708,N_8882);
nand UO_2 (O_2,N_7730,N_8085);
and UO_3 (O_3,N_9537,N_9794);
nor UO_4 (O_4,N_9825,N_7552);
and UO_5 (O_5,N_9745,N_8825);
or UO_6 (O_6,N_8601,N_7922);
or UO_7 (O_7,N_9229,N_8005);
nor UO_8 (O_8,N_7896,N_8096);
or UO_9 (O_9,N_8612,N_8669);
or UO_10 (O_10,N_8387,N_8023);
or UO_11 (O_11,N_8801,N_8166);
or UO_12 (O_12,N_9432,N_9602);
nor UO_13 (O_13,N_8804,N_8087);
nand UO_14 (O_14,N_9230,N_8870);
or UO_15 (O_15,N_7527,N_8433);
or UO_16 (O_16,N_8182,N_8131);
nor UO_17 (O_17,N_9726,N_8768);
xor UO_18 (O_18,N_7990,N_8875);
and UO_19 (O_19,N_8216,N_8456);
and UO_20 (O_20,N_7688,N_8396);
or UO_21 (O_21,N_8385,N_9623);
nor UO_22 (O_22,N_9577,N_9416);
nor UO_23 (O_23,N_8064,N_9682);
or UO_24 (O_24,N_9600,N_7947);
or UO_25 (O_25,N_9518,N_7856);
nor UO_26 (O_26,N_8996,N_8472);
xor UO_27 (O_27,N_7549,N_7544);
nand UO_28 (O_28,N_8817,N_8880);
nor UO_29 (O_29,N_9816,N_8213);
nor UO_30 (O_30,N_8530,N_9281);
and UO_31 (O_31,N_9985,N_7735);
nor UO_32 (O_32,N_8859,N_7720);
or UO_33 (O_33,N_7818,N_9860);
xnor UO_34 (O_34,N_9197,N_8294);
and UO_35 (O_35,N_8717,N_8307);
or UO_36 (O_36,N_9504,N_7602);
and UO_37 (O_37,N_9711,N_7944);
nor UO_38 (O_38,N_9851,N_9071);
and UO_39 (O_39,N_8537,N_7873);
nor UO_40 (O_40,N_9942,N_9909);
nor UO_41 (O_41,N_9944,N_8247);
and UO_42 (O_42,N_8257,N_7752);
nor UO_43 (O_43,N_8561,N_8262);
nor UO_44 (O_44,N_8480,N_7572);
nor UO_45 (O_45,N_9929,N_7807);
nor UO_46 (O_46,N_8376,N_8624);
or UO_47 (O_47,N_8107,N_9172);
and UO_48 (O_48,N_7661,N_9262);
nor UO_49 (O_49,N_8366,N_9439);
nor UO_50 (O_50,N_7874,N_9332);
or UO_51 (O_51,N_8125,N_7779);
and UO_52 (O_52,N_9468,N_9203);
nor UO_53 (O_53,N_9486,N_7765);
xnor UO_54 (O_54,N_8532,N_8957);
or UO_55 (O_55,N_8050,N_7576);
and UO_56 (O_56,N_8409,N_8414);
nor UO_57 (O_57,N_9303,N_9645);
nor UO_58 (O_58,N_8716,N_9192);
and UO_59 (O_59,N_9383,N_8094);
nand UO_60 (O_60,N_7728,N_9307);
and UO_61 (O_61,N_8171,N_7995);
or UO_62 (O_62,N_9924,N_8721);
and UO_63 (O_63,N_9419,N_9854);
and UO_64 (O_64,N_7609,N_9263);
or UO_65 (O_65,N_7813,N_7789);
and UO_66 (O_66,N_8205,N_7969);
nor UO_67 (O_67,N_7895,N_9343);
nor UO_68 (O_68,N_9939,N_7855);
or UO_69 (O_69,N_8685,N_8489);
or UO_70 (O_70,N_9215,N_8885);
nand UO_71 (O_71,N_8299,N_9019);
nor UO_72 (O_72,N_9817,N_9260);
or UO_73 (O_73,N_7999,N_8623);
nand UO_74 (O_74,N_8097,N_9901);
nand UO_75 (O_75,N_8117,N_8128);
or UO_76 (O_76,N_7601,N_9920);
and UO_77 (O_77,N_7748,N_9231);
or UO_78 (O_78,N_7757,N_9448);
nand UO_79 (O_79,N_7773,N_8405);
or UO_80 (O_80,N_9484,N_9082);
nor UO_81 (O_81,N_9357,N_8520);
xor UO_82 (O_82,N_8713,N_8983);
and UO_83 (O_83,N_7968,N_9361);
nand UO_84 (O_84,N_9405,N_8383);
nor UO_85 (O_85,N_9898,N_7580);
and UO_86 (O_86,N_9717,N_9005);
nand UO_87 (O_87,N_8587,N_9927);
nor UO_88 (O_88,N_7745,N_9747);
or UO_89 (O_89,N_8941,N_8554);
nor UO_90 (O_90,N_8726,N_7917);
nor UO_91 (O_91,N_7866,N_9770);
or UO_92 (O_92,N_9107,N_9205);
nand UO_93 (O_93,N_7673,N_7579);
and UO_94 (O_94,N_8905,N_8673);
nor UO_95 (O_95,N_8608,N_8364);
and UO_96 (O_96,N_9850,N_8846);
nor UO_97 (O_97,N_9266,N_9769);
xnor UO_98 (O_98,N_9295,N_8045);
nor UO_99 (O_99,N_8206,N_8279);
and UO_100 (O_100,N_8080,N_9418);
and UO_101 (O_101,N_8931,N_9715);
nand UO_102 (O_102,N_8938,N_9812);
nor UO_103 (O_103,N_8700,N_8703);
nor UO_104 (O_104,N_8656,N_9237);
nand UO_105 (O_105,N_9204,N_9591);
and UO_106 (O_106,N_9589,N_8598);
nor UO_107 (O_107,N_8120,N_8487);
nor UO_108 (O_108,N_7829,N_9169);
or UO_109 (O_109,N_8872,N_7702);
xor UO_110 (O_110,N_7657,N_8900);
nor UO_111 (O_111,N_8347,N_8536);
nor UO_112 (O_112,N_9114,N_7827);
nor UO_113 (O_113,N_9248,N_8785);
or UO_114 (O_114,N_7506,N_9056);
nand UO_115 (O_115,N_7791,N_7704);
nand UO_116 (O_116,N_7690,N_7772);
nor UO_117 (O_117,N_7908,N_8670);
or UO_118 (O_118,N_8403,N_8625);
or UO_119 (O_119,N_8004,N_8814);
and UO_120 (O_120,N_7509,N_9883);
or UO_121 (O_121,N_8044,N_7986);
or UO_122 (O_122,N_7965,N_8515);
nand UO_123 (O_123,N_8394,N_8193);
and UO_124 (O_124,N_8769,N_7733);
nor UO_125 (O_125,N_7905,N_7758);
nand UO_126 (O_126,N_7897,N_9157);
or UO_127 (O_127,N_8180,N_8651);
or UO_128 (O_128,N_8548,N_8633);
nor UO_129 (O_129,N_8642,N_9786);
nand UO_130 (O_130,N_8968,N_8657);
nor UO_131 (O_131,N_8783,N_8209);
xnor UO_132 (O_132,N_8372,N_9138);
and UO_133 (O_133,N_7822,N_8643);
and UO_134 (O_134,N_8820,N_8511);
or UO_135 (O_135,N_8920,N_7608);
nand UO_136 (O_136,N_9167,N_8384);
xor UO_137 (O_137,N_9836,N_9534);
nor UO_138 (O_138,N_8415,N_8610);
and UO_139 (O_139,N_9321,N_8142);
or UO_140 (O_140,N_7635,N_9364);
or UO_141 (O_141,N_8184,N_8545);
nand UO_142 (O_142,N_9308,N_8252);
nor UO_143 (O_143,N_7899,N_9703);
nor UO_144 (O_144,N_8140,N_9346);
nor UO_145 (O_145,N_7597,N_8778);
and UO_146 (O_146,N_9811,N_9838);
nand UO_147 (O_147,N_7668,N_9906);
nand UO_148 (O_148,N_8422,N_8162);
or UO_149 (O_149,N_8151,N_9656);
nor UO_150 (O_150,N_9273,N_8571);
and UO_151 (O_151,N_8639,N_8179);
nand UO_152 (O_152,N_9585,N_9800);
and UO_153 (O_153,N_9543,N_8637);
or UO_154 (O_154,N_9669,N_8310);
or UO_155 (O_155,N_7877,N_9970);
and UO_156 (O_156,N_9644,N_7556);
nand UO_157 (O_157,N_9768,N_8831);
and UO_158 (O_158,N_8380,N_9814);
nor UO_159 (O_159,N_9080,N_9158);
and UO_160 (O_160,N_9557,N_9441);
or UO_161 (O_161,N_7639,N_7871);
nand UO_162 (O_162,N_9788,N_9104);
and UO_163 (O_163,N_9379,N_8565);
nand UO_164 (O_164,N_9899,N_7981);
or UO_165 (O_165,N_7820,N_8873);
or UO_166 (O_166,N_8283,N_8081);
nand UO_167 (O_167,N_7755,N_8513);
nor UO_168 (O_168,N_9422,N_8326);
and UO_169 (O_169,N_9487,N_9451);
nand UO_170 (O_170,N_9362,N_9784);
or UO_171 (O_171,N_8190,N_8771);
and UO_172 (O_172,N_9617,N_8406);
or UO_173 (O_173,N_9210,N_8455);
and UO_174 (O_174,N_9724,N_8517);
nand UO_175 (O_175,N_9756,N_8744);
nand UO_176 (O_176,N_9828,N_9201);
and UO_177 (O_177,N_7562,N_9615);
nand UO_178 (O_178,N_7536,N_8926);
or UO_179 (O_179,N_9185,N_9036);
nand UO_180 (O_180,N_9221,N_8784);
or UO_181 (O_181,N_9672,N_9098);
or UO_182 (O_182,N_8998,N_9957);
and UO_183 (O_183,N_9922,N_9493);
nand UO_184 (O_184,N_9896,N_9029);
and UO_185 (O_185,N_9601,N_8187);
and UO_186 (O_186,N_8779,N_9731);
nor UO_187 (O_187,N_7614,N_8711);
xnor UO_188 (O_188,N_7727,N_9502);
and UO_189 (O_189,N_9755,N_9519);
nand UO_190 (O_190,N_9734,N_9241);
or UO_191 (O_191,N_8139,N_9884);
nand UO_192 (O_192,N_9253,N_9966);
or UO_193 (O_193,N_7988,N_7526);
nor UO_194 (O_194,N_9533,N_9477);
xnor UO_195 (O_195,N_7846,N_8352);
xor UO_196 (O_196,N_9729,N_7564);
nor UO_197 (O_197,N_9514,N_8071);
nand UO_198 (O_198,N_8550,N_9633);
nor UO_199 (O_199,N_7975,N_7776);
and UO_200 (O_200,N_8292,N_8954);
nor UO_201 (O_201,N_8172,N_9127);
or UO_202 (O_202,N_9956,N_7978);
and UO_203 (O_203,N_8330,N_9753);
or UO_204 (O_204,N_7522,N_8696);
and UO_205 (O_205,N_9099,N_7849);
nor UO_206 (O_206,N_9511,N_9730);
xnor UO_207 (O_207,N_9181,N_8258);
nor UO_208 (O_208,N_7740,N_8278);
or UO_209 (O_209,N_8516,N_9044);
nand UO_210 (O_210,N_8564,N_8523);
and UO_211 (O_211,N_9213,N_8393);
nand UO_212 (O_212,N_9949,N_8723);
and UO_213 (O_213,N_8966,N_8095);
nand UO_214 (O_214,N_8890,N_9987);
or UO_215 (O_215,N_8596,N_9277);
and UO_216 (O_216,N_8178,N_9718);
and UO_217 (O_217,N_8073,N_8776);
nand UO_218 (O_218,N_9495,N_8246);
or UO_219 (O_219,N_9870,N_9251);
or UO_220 (O_220,N_7598,N_9491);
or UO_221 (O_221,N_8566,N_8359);
nand UO_222 (O_222,N_9936,N_7606);
or UO_223 (O_223,N_8597,N_9604);
and UO_224 (O_224,N_8593,N_9696);
or UO_225 (O_225,N_9848,N_7955);
nand UO_226 (O_226,N_8975,N_8982);
and UO_227 (O_227,N_8930,N_7670);
nor UO_228 (O_228,N_8275,N_9077);
nand UO_229 (O_229,N_9049,N_9837);
or UO_230 (O_230,N_9023,N_9928);
nor UO_231 (O_231,N_8582,N_7898);
nand UO_232 (O_232,N_9530,N_9396);
and UO_233 (O_233,N_7594,N_9444);
nor UO_234 (O_234,N_9286,N_9888);
nor UO_235 (O_235,N_8604,N_8256);
xor UO_236 (O_236,N_7911,N_8945);
and UO_237 (O_237,N_7587,N_9395);
nor UO_238 (O_238,N_9829,N_8600);
and UO_239 (O_239,N_8646,N_8719);
nor UO_240 (O_240,N_9186,N_9775);
and UO_241 (O_241,N_9677,N_7920);
and UO_242 (O_242,N_8039,N_9638);
nand UO_243 (O_243,N_9568,N_9259);
nand UO_244 (O_244,N_9905,N_7555);
nor UO_245 (O_245,N_8411,N_8958);
nor UO_246 (O_246,N_8104,N_9655);
nor UO_247 (O_247,N_8847,N_8068);
nor UO_248 (O_248,N_7739,N_9805);
or UO_249 (O_249,N_9710,N_9844);
nand UO_250 (O_250,N_8892,N_9914);
nand UO_251 (O_251,N_8720,N_9121);
and UO_252 (O_252,N_7810,N_8743);
nor UO_253 (O_253,N_8022,N_9834);
nand UO_254 (O_254,N_9574,N_9762);
nand UO_255 (O_255,N_7656,N_8132);
nor UO_256 (O_256,N_9761,N_9686);
or UO_257 (O_257,N_8250,N_8148);
or UO_258 (O_258,N_7956,N_9426);
or UO_259 (O_259,N_9129,N_8533);
or UO_260 (O_260,N_9522,N_7630);
or UO_261 (O_261,N_9060,N_9141);
or UO_262 (O_262,N_7714,N_9429);
and UO_263 (O_263,N_7962,N_8876);
or UO_264 (O_264,N_9527,N_7516);
nor UO_265 (O_265,N_8976,N_8955);
nand UO_266 (O_266,N_9421,N_8447);
nor UO_267 (O_267,N_9973,N_9627);
nor UO_268 (O_268,N_8186,N_9058);
nor UO_269 (O_269,N_8099,N_8581);
or UO_270 (O_270,N_9685,N_9605);
nor UO_271 (O_271,N_8621,N_9050);
or UO_272 (O_272,N_9620,N_9801);
nand UO_273 (O_273,N_8553,N_7531);
and UO_274 (O_274,N_9390,N_7761);
or UO_275 (O_275,N_7811,N_9716);
or UO_276 (O_276,N_8869,N_9320);
or UO_277 (O_277,N_9055,N_8054);
nor UO_278 (O_278,N_8706,N_9063);
nor UO_279 (O_279,N_8198,N_8122);
or UO_280 (O_280,N_9120,N_8842);
or UO_281 (O_281,N_9930,N_9199);
nor UO_282 (O_282,N_8344,N_9692);
nand UO_283 (O_283,N_8340,N_8135);
nand UO_284 (O_284,N_8204,N_7759);
and UO_285 (O_285,N_8217,N_7993);
or UO_286 (O_286,N_8038,N_9274);
or UO_287 (O_287,N_9759,N_8464);
nand UO_288 (O_288,N_9030,N_8276);
and UO_289 (O_289,N_8630,N_9806);
nor UO_290 (O_290,N_7775,N_9802);
nand UO_291 (O_291,N_7629,N_9482);
xor UO_292 (O_292,N_7798,N_9960);
nand UO_293 (O_293,N_8650,N_9641);
and UO_294 (O_294,N_9465,N_9123);
or UO_295 (O_295,N_7880,N_9146);
or UO_296 (O_296,N_9377,N_9271);
nand UO_297 (O_297,N_8261,N_9431);
nor UO_298 (O_298,N_9306,N_9176);
and UO_299 (O_299,N_9846,N_9112);
nor UO_300 (O_300,N_8745,N_8302);
and UO_301 (O_301,N_9469,N_9526);
nor UO_302 (O_302,N_8987,N_8838);
and UO_303 (O_303,N_9485,N_7838);
or UO_304 (O_304,N_9833,N_8255);
nand UO_305 (O_305,N_8751,N_9516);
nor UO_306 (O_306,N_7738,N_9116);
nand UO_307 (O_307,N_9918,N_7510);
and UO_308 (O_308,N_8884,N_9551);
and UO_309 (O_309,N_9272,N_9689);
or UO_310 (O_310,N_9865,N_9025);
and UO_311 (O_311,N_8683,N_8453);
or UO_312 (O_312,N_8948,N_9318);
nand UO_313 (O_313,N_9868,N_8089);
nand UO_314 (O_314,N_8407,N_7860);
or UO_315 (O_315,N_8871,N_9174);
nand UO_316 (O_316,N_7966,N_7957);
nand UO_317 (O_317,N_8021,N_8688);
nand UO_318 (O_318,N_9773,N_8568);
nand UO_319 (O_319,N_8260,N_8615);
and UO_320 (O_320,N_9965,N_9570);
and UO_321 (O_321,N_9268,N_8234);
or UO_322 (O_322,N_8188,N_7857);
nor UO_323 (O_323,N_7613,N_8300);
nand UO_324 (O_324,N_8781,N_9643);
nand UO_325 (O_325,N_7709,N_8508);
nor UO_326 (O_326,N_8853,N_7655);
or UO_327 (O_327,N_8944,N_8210);
and UO_328 (O_328,N_9592,N_8609);
nor UO_329 (O_329,N_8037,N_7972);
nor UO_330 (O_330,N_8857,N_7611);
nand UO_331 (O_331,N_7731,N_9256);
nor UO_332 (O_332,N_8828,N_7650);
or UO_333 (O_333,N_8663,N_7582);
and UO_334 (O_334,N_8457,N_8585);
or UO_335 (O_335,N_8592,N_9911);
nor UO_336 (O_336,N_7677,N_8752);
and UO_337 (O_337,N_9351,N_7753);
nor UO_338 (O_338,N_8059,N_8235);
nand UO_339 (O_339,N_8413,N_8689);
nand UO_340 (O_340,N_8271,N_9872);
xnor UO_341 (O_341,N_8556,N_8429);
or UO_342 (O_342,N_8273,N_9249);
and UO_343 (O_343,N_8959,N_7959);
or UO_344 (O_344,N_9879,N_8787);
and UO_345 (O_345,N_9744,N_7692);
or UO_346 (O_346,N_9581,N_7826);
nor UO_347 (O_347,N_8167,N_8978);
and UO_348 (O_348,N_7924,N_7561);
nor UO_349 (O_349,N_9874,N_8607);
nand UO_350 (O_350,N_7754,N_8728);
and UO_351 (O_351,N_9573,N_8789);
and UO_352 (O_352,N_7628,N_8896);
and UO_353 (O_353,N_8452,N_8077);
nor UO_354 (O_354,N_8908,N_8780);
nand UO_355 (O_355,N_8061,N_9582);
nand UO_356 (O_356,N_9776,N_9206);
nor UO_357 (O_357,N_8546,N_8067);
nor UO_358 (O_358,N_9414,N_9635);
xnor UO_359 (O_359,N_9629,N_7521);
or UO_360 (O_360,N_8694,N_8439);
and UO_361 (O_361,N_7648,N_8488);
and UO_362 (O_362,N_8986,N_8351);
or UO_363 (O_363,N_8834,N_9086);
nor UO_364 (O_364,N_8334,N_8019);
and UO_365 (O_365,N_7676,N_9932);
nor UO_366 (O_366,N_9375,N_7770);
nand UO_367 (O_367,N_8569,N_9663);
nor UO_368 (O_368,N_8109,N_8686);
nor UO_369 (O_369,N_9136,N_8704);
or UO_370 (O_370,N_7919,N_9191);
or UO_371 (O_371,N_9391,N_7742);
and UO_372 (O_372,N_8988,N_7963);
nor UO_373 (O_373,N_7964,N_9139);
nand UO_374 (O_374,N_9075,N_8041);
nor UO_375 (O_375,N_8648,N_9064);
or UO_376 (O_376,N_9190,N_9069);
xor UO_377 (O_377,N_9549,N_9178);
and UO_378 (O_378,N_9137,N_7557);
nor UO_379 (O_379,N_7584,N_8309);
or UO_380 (O_380,N_8124,N_8365);
nor UO_381 (O_381,N_9472,N_7710);
nand UO_382 (O_382,N_9247,N_7891);
nor UO_383 (O_383,N_9880,N_8977);
or UO_384 (O_384,N_8692,N_7513);
nand UO_385 (O_385,N_9532,N_8211);
or UO_386 (O_386,N_9611,N_7799);
nand UO_387 (O_387,N_9741,N_7788);
or UO_388 (O_388,N_9925,N_9344);
and UO_389 (O_389,N_8417,N_9316);
and UO_390 (O_390,N_8829,N_9388);
nand UO_391 (O_391,N_8355,N_9873);
nor UO_392 (O_392,N_7713,N_9087);
or UO_393 (O_393,N_9445,N_9242);
or UO_394 (O_394,N_9842,N_9946);
nand UO_395 (O_395,N_8503,N_8850);
and UO_396 (O_396,N_7583,N_7687);
or UO_397 (O_397,N_9588,N_9859);
nor UO_398 (O_398,N_7669,N_9435);
nor UO_399 (O_399,N_9983,N_7563);
nand UO_400 (O_400,N_8268,N_8232);
or UO_401 (O_401,N_8123,N_8191);
or UO_402 (O_402,N_7746,N_8865);
nor UO_403 (O_403,N_9180,N_8697);
or UO_404 (O_404,N_7722,N_8725);
nor UO_405 (O_405,N_9891,N_8408);
nor UO_406 (O_406,N_8315,N_7851);
and UO_407 (O_407,N_9733,N_9820);
or UO_408 (O_408,N_9521,N_8181);
nor UO_409 (O_409,N_9841,N_7543);
or UO_410 (O_410,N_9774,N_7945);
nor UO_411 (O_411,N_8377,N_9073);
nor UO_412 (O_412,N_7693,N_9035);
and UO_413 (O_413,N_8014,N_9803);
nor UO_414 (O_414,N_9590,N_8765);
nor UO_415 (O_415,N_8567,N_7662);
and UO_416 (O_416,N_7703,N_7892);
xor UO_417 (O_417,N_9554,N_8588);
and UO_418 (O_418,N_8519,N_9683);
nor UO_419 (O_419,N_9542,N_8177);
nand UO_420 (O_420,N_8962,N_8301);
xnor UO_421 (O_421,N_9131,N_7520);
nor UO_422 (O_422,N_9291,N_9651);
nand UO_423 (O_423,N_7805,N_9397);
nand UO_424 (O_424,N_7689,N_9488);
nor UO_425 (O_425,N_8888,N_8318);
nor UO_426 (O_426,N_9171,N_7502);
nand UO_427 (O_427,N_8845,N_9561);
xor UO_428 (O_428,N_8620,N_8492);
or UO_429 (O_429,N_9566,N_7640);
xor UO_430 (O_430,N_9010,N_8494);
or UO_431 (O_431,N_8985,N_8722);
or UO_432 (O_432,N_8999,N_9048);
nor UO_433 (O_433,N_7645,N_8507);
nand UO_434 (O_434,N_8086,N_9338);
and UO_435 (O_435,N_9311,N_8467);
nand UO_436 (O_436,N_8251,N_7607);
xor UO_437 (O_437,N_9789,N_9154);
nand UO_438 (O_438,N_8940,N_9017);
and UO_439 (O_439,N_9456,N_9309);
or UO_440 (O_440,N_9606,N_8707);
or UO_441 (O_441,N_7812,N_9553);
and UO_442 (O_442,N_9470,N_9151);
or UO_443 (O_443,N_7801,N_9302);
and UO_444 (O_444,N_9305,N_9989);
nand UO_445 (O_445,N_8329,N_9093);
or UO_446 (O_446,N_9219,N_9312);
and UO_447 (O_447,N_8879,N_8390);
nor UO_448 (O_448,N_9567,N_9618);
and UO_449 (O_449,N_8018,N_8868);
and UO_450 (O_450,N_8430,N_8052);
and UO_451 (O_451,N_8062,N_8265);
and UO_452 (O_452,N_7828,N_9406);
nand UO_453 (O_453,N_9360,N_8736);
nand UO_454 (O_454,N_9424,N_9953);
or UO_455 (O_455,N_7989,N_7793);
and UO_456 (O_456,N_9895,N_9184);
or UO_457 (O_457,N_8136,N_7567);
nand UO_458 (O_458,N_7715,N_9436);
nand UO_459 (O_459,N_8638,N_7647);
nor UO_460 (O_460,N_8147,N_8227);
and UO_461 (O_461,N_9150,N_9506);
nand UO_462 (O_462,N_9818,N_8809);
and UO_463 (O_463,N_9373,N_9548);
nand UO_464 (O_464,N_9646,N_8036);
nand UO_465 (O_465,N_9125,N_9727);
nand UO_466 (O_466,N_8233,N_7603);
nand UO_467 (O_467,N_8027,N_9287);
nor UO_468 (O_468,N_9649,N_8155);
or UO_469 (O_469,N_8647,N_8916);
nor UO_470 (O_470,N_9298,N_8306);
and UO_471 (O_471,N_8731,N_9857);
and UO_472 (O_472,N_8427,N_9474);
nand UO_473 (O_473,N_7699,N_9684);
nor UO_474 (O_474,N_9317,N_8950);
nand UO_475 (O_475,N_7681,N_9547);
or UO_476 (O_476,N_9688,N_8195);
or UO_477 (O_477,N_7953,N_9937);
nor UO_478 (O_478,N_8426,N_9155);
or UO_479 (O_479,N_7800,N_8043);
nand UO_480 (O_480,N_7833,N_8629);
or UO_481 (O_481,N_9001,N_9780);
and UO_482 (O_482,N_9849,N_9562);
nand UO_483 (O_483,N_8346,N_8370);
nor UO_484 (O_484,N_9265,N_9033);
nor UO_485 (O_485,N_9257,N_9376);
and UO_486 (O_486,N_7633,N_8715);
nand UO_487 (O_487,N_8048,N_8678);
nand UO_488 (O_488,N_9763,N_9997);
nor UO_489 (O_489,N_9349,N_9301);
nand UO_490 (O_490,N_7631,N_9027);
nand UO_491 (O_491,N_8102,N_9402);
xor UO_492 (O_492,N_8748,N_7718);
or UO_493 (O_493,N_9804,N_7847);
nor UO_494 (O_494,N_9721,N_9232);
or UO_495 (O_495,N_9153,N_8493);
nand UO_496 (O_496,N_9188,N_7823);
nand UO_497 (O_497,N_9065,N_8145);
nand UO_498 (O_498,N_9853,N_8732);
nand UO_499 (O_499,N_9198,N_8358);
or UO_500 (O_500,N_7553,N_8101);
nor UO_501 (O_501,N_9982,N_7627);
or UO_502 (O_502,N_8058,N_7705);
nand UO_503 (O_503,N_7653,N_8777);
nand UO_504 (O_504,N_8555,N_7534);
nor UO_505 (O_505,N_9143,N_8486);
nand UO_506 (O_506,N_8214,N_7889);
nor UO_507 (O_507,N_9455,N_9382);
nor UO_508 (O_508,N_8574,N_9524);
or UO_509 (O_509,N_8543,N_7641);
nor UO_510 (O_510,N_7806,N_8212);
nor UO_511 (O_511,N_8170,N_8308);
nor UO_512 (O_512,N_9665,N_8682);
or UO_513 (O_513,N_8012,N_9059);
xnor UO_514 (O_514,N_9675,N_7604);
or UO_515 (O_515,N_9785,N_8652);
nor UO_516 (O_516,N_9166,N_8756);
or UO_517 (O_517,N_7983,N_9212);
or UO_518 (O_518,N_7893,N_7696);
nor UO_519 (O_519,N_9520,N_9039);
nand UO_520 (O_520,N_9015,N_9765);
nor UO_521 (O_521,N_7726,N_9326);
nand UO_522 (O_522,N_9464,N_8912);
nand UO_523 (O_523,N_7698,N_7697);
nor UO_524 (O_524,N_7961,N_8603);
nor UO_525 (O_525,N_8946,N_9764);
nor UO_526 (O_526,N_9195,N_8143);
nand UO_527 (O_527,N_9777,N_8911);
nor UO_528 (O_528,N_8443,N_8510);
nand UO_529 (O_529,N_9680,N_9179);
or UO_530 (O_530,N_9479,N_9862);
or UO_531 (O_531,N_8671,N_8267);
nand UO_532 (O_532,N_9845,N_9117);
nand UO_533 (O_533,N_9378,N_7783);
nor UO_534 (O_534,N_8542,N_9637);
or UO_535 (O_535,N_7814,N_7803);
nor UO_536 (O_536,N_8356,N_9324);
or UO_537 (O_537,N_8730,N_8812);
nand UO_538 (O_538,N_9616,N_8606);
and UO_539 (O_539,N_7907,N_9132);
nor UO_540 (O_540,N_9494,N_8848);
nor UO_541 (O_541,N_8434,N_8254);
or UO_542 (O_542,N_8797,N_8450);
or UO_543 (O_543,N_8465,N_7998);
and UO_544 (O_544,N_7625,N_8491);
nor UO_545 (O_545,N_8514,N_7537);
and UO_546 (O_546,N_9245,N_7712);
nor UO_547 (O_547,N_7862,N_9450);
or UO_548 (O_548,N_8599,N_8796);
and UO_549 (O_549,N_9827,N_9668);
nor UO_550 (O_550,N_8851,N_9356);
nand UO_551 (O_551,N_9160,N_7948);
xor UO_552 (O_552,N_7570,N_7790);
or UO_553 (O_553,N_8821,N_7987);
and UO_554 (O_554,N_9003,N_7683);
or UO_555 (O_555,N_8734,N_8981);
nor UO_556 (O_556,N_8074,N_8617);
and UO_557 (O_557,N_9403,N_8887);
nand UO_558 (O_558,N_9740,N_9975);
nand UO_559 (O_559,N_7724,N_7763);
or UO_560 (O_560,N_9948,N_8460);
nor UO_561 (O_561,N_7646,N_9639);
nand UO_562 (O_562,N_7589,N_9447);
nor UO_563 (O_563,N_8325,N_9043);
nor UO_564 (O_564,N_8215,N_9512);
nor UO_565 (O_565,N_9124,N_9187);
or UO_566 (O_566,N_9754,N_8013);
nor UO_567 (O_567,N_8055,N_9342);
and UO_568 (O_568,N_8655,N_9847);
or UO_569 (O_569,N_7508,N_8904);
nor UO_570 (O_570,N_7588,N_8057);
or UO_571 (O_571,N_9270,N_7910);
and UO_572 (O_572,N_9294,N_9076);
and UO_573 (O_573,N_7929,N_9018);
nand UO_574 (O_574,N_7660,N_8541);
nand UO_575 (O_575,N_8010,N_8007);
or UO_576 (O_576,N_9284,N_9791);
nand UO_577 (O_577,N_9950,N_9892);
or UO_578 (O_578,N_8339,N_9224);
nor UO_579 (O_579,N_7706,N_7926);
nor UO_580 (O_580,N_8738,N_7734);
and UO_581 (O_581,N_8627,N_8197);
nor UO_582 (O_582,N_8425,N_8906);
or UO_583 (O_583,N_8535,N_9409);
nor UO_584 (O_584,N_8584,N_8967);
or UO_585 (O_585,N_7787,N_9938);
xnor UO_586 (O_586,N_8333,N_8379);
or UO_587 (O_587,N_9810,N_8551);
and UO_588 (O_588,N_8644,N_7565);
and UO_589 (O_589,N_9037,N_8219);
or UO_590 (O_590,N_8051,N_7994);
nor UO_591 (O_591,N_8544,N_8762);
or UO_592 (O_592,N_8994,N_9159);
or UO_593 (O_593,N_8654,N_9333);
nor UO_594 (O_594,N_7869,N_8238);
xnor UO_595 (O_595,N_9239,N_8091);
nand UO_596 (O_596,N_8805,N_7723);
or UO_597 (O_597,N_9217,N_9995);
and UO_598 (O_598,N_7512,N_7915);
nand UO_599 (O_599,N_9743,N_8361);
nand UO_600 (O_600,N_9134,N_7736);
nand UO_601 (O_601,N_8808,N_7585);
nor UO_602 (O_602,N_7744,N_8531);
or UO_603 (O_603,N_8923,N_7780);
and UO_604 (O_604,N_9130,N_8935);
or UO_605 (O_605,N_8118,N_8224);
nand UO_606 (O_606,N_9809,N_8223);
or UO_607 (O_607,N_9913,N_9958);
and UO_608 (O_608,N_9650,N_9430);
and UO_609 (O_609,N_8286,N_8645);
nand UO_610 (O_610,N_8521,N_8322);
and UO_611 (O_611,N_7934,N_9128);
or UO_612 (O_612,N_9452,N_9067);
or UO_613 (O_613,N_9757,N_9921);
nor UO_614 (O_614,N_9334,N_9923);
and UO_615 (O_615,N_9040,N_8589);
and UO_616 (O_616,N_8910,N_7651);
nor UO_617 (O_617,N_9622,N_9489);
nand UO_618 (O_618,N_9787,N_8733);
nor UO_619 (O_619,N_8203,N_9283);
nor UO_620 (O_620,N_8056,N_8973);
nand UO_621 (O_621,N_8028,N_8437);
nor UO_622 (O_622,N_7747,N_8702);
and UO_623 (O_623,N_9002,N_9483);
and UO_624 (O_624,N_8474,N_7741);
and UO_625 (O_625,N_7938,N_9564);
and UO_626 (O_626,N_9563,N_7865);
or UO_627 (O_627,N_8207,N_7560);
nand UO_628 (O_628,N_9149,N_9168);
or UO_629 (O_629,N_9575,N_7928);
nor UO_630 (O_630,N_7909,N_9540);
or UO_631 (O_631,N_8354,N_7550);
nand UO_632 (O_632,N_8183,N_7782);
nand UO_633 (O_633,N_8909,N_8786);
or UO_634 (O_634,N_7804,N_7936);
nand UO_635 (O_635,N_9636,N_7619);
and UO_636 (O_636,N_7605,N_8463);
or UO_637 (O_637,N_8628,N_7636);
nand UO_638 (O_638,N_9678,N_7528);
nor UO_639 (O_639,N_8595,N_8758);
or UO_640 (O_640,N_8807,N_9410);
and UO_641 (O_641,N_9824,N_9440);
nor UO_642 (O_642,N_8939,N_8154);
nor UO_643 (O_643,N_9194,N_7675);
or UO_644 (O_644,N_9140,N_9999);
and UO_645 (O_645,N_7599,N_9476);
and UO_646 (O_646,N_9061,N_8176);
nand UO_647 (O_647,N_9313,N_9855);
and UO_648 (O_648,N_7686,N_8806);
or UO_649 (O_649,N_8591,N_8894);
or UO_650 (O_650,N_9051,N_9631);
or UO_651 (O_651,N_7882,N_9238);
nand UO_652 (O_652,N_9742,N_8070);
or UO_653 (O_653,N_8843,N_9471);
nand UO_654 (O_654,N_8932,N_9832);
nor UO_655 (O_655,N_8381,N_9091);
nand UO_656 (O_656,N_8083,N_8701);
nor UO_657 (O_657,N_8032,N_8189);
and UO_658 (O_658,N_9016,N_8559);
or UO_659 (O_659,N_8008,N_9503);
nor UO_660 (O_660,N_8483,N_8304);
xnor UO_661 (O_661,N_9529,N_9613);
or UO_662 (O_662,N_9458,N_7749);
and UO_663 (O_663,N_9461,N_9882);
nand UO_664 (O_664,N_7548,N_8353);
or UO_665 (O_665,N_8740,N_8727);
nand UO_666 (O_666,N_8490,N_7885);
or UO_667 (O_667,N_8914,N_9728);
and UO_668 (O_668,N_8895,N_7795);
xnor UO_669 (O_669,N_8698,N_9941);
or UO_670 (O_670,N_8680,N_8440);
and UO_671 (O_671,N_7518,N_8201);
and UO_672 (O_672,N_9808,N_9867);
or UO_673 (O_673,N_9449,N_9752);
nand UO_674 (O_674,N_9234,N_9135);
xor UO_675 (O_675,N_9760,N_8378);
nand UO_676 (O_676,N_9693,N_8391);
nand UO_677 (O_677,N_8759,N_8813);
or UO_678 (O_678,N_8270,N_9009);
nor UO_679 (O_679,N_9915,N_7778);
and UO_680 (O_680,N_8192,N_9988);
or UO_681 (O_681,N_8127,N_9007);
nand UO_682 (O_682,N_9586,N_9235);
or UO_683 (O_683,N_8739,N_9423);
or UO_684 (O_684,N_9399,N_7767);
nor UO_685 (O_685,N_8774,N_7875);
or UO_686 (O_686,N_9113,N_9657);
nand UO_687 (O_687,N_7511,N_9671);
nand UO_688 (O_688,N_9681,N_7887);
or UO_689 (O_689,N_8435,N_7836);
and UO_690 (O_690,N_8382,N_9304);
nand UO_691 (O_691,N_9697,N_8679);
nand UO_692 (O_692,N_9142,N_7716);
nor UO_693 (O_693,N_8907,N_7996);
nand UO_694 (O_694,N_9374,N_9370);
or UO_695 (O_695,N_9193,N_9443);
or UO_696 (O_696,N_8836,N_9583);
or UO_697 (O_697,N_9517,N_8431);
nor UO_698 (O_698,N_9706,N_9336);
nor UO_699 (O_699,N_7950,N_9442);
or UO_700 (O_700,N_9793,N_9595);
nor UO_701 (O_701,N_9408,N_9830);
and UO_702 (O_702,N_8861,N_9767);
nand UO_703 (O_703,N_7612,N_8712);
nand UO_704 (O_704,N_8709,N_9106);
and UO_705 (O_705,N_8919,N_9823);
xnor UO_706 (O_706,N_8921,N_8862);
and UO_707 (O_707,N_8296,N_9216);
nand UO_708 (O_708,N_8763,N_7667);
xnor UO_709 (O_709,N_8485,N_8735);
nand UO_710 (O_710,N_9699,N_8332);
nor UO_711 (O_711,N_8622,N_7638);
and UO_712 (O_712,N_8672,N_8891);
xnor UO_713 (O_713,N_7593,N_8991);
nor UO_714 (O_714,N_8134,N_7643);
nor UO_715 (O_715,N_7774,N_8667);
and UO_716 (O_716,N_7575,N_9425);
nand UO_717 (O_717,N_9739,N_8802);
or UO_718 (O_718,N_8934,N_9108);
nor UO_719 (O_719,N_9782,N_9790);
and UO_720 (O_720,N_8832,N_8269);
nor UO_721 (O_721,N_9746,N_9090);
or UO_722 (O_722,N_7824,N_9890);
xor UO_723 (O_723,N_7695,N_8795);
nand UO_724 (O_724,N_7618,N_9621);
nand UO_725 (O_725,N_7751,N_9569);
xor UO_726 (O_726,N_8199,N_9492);
nand UO_727 (O_727,N_9042,N_9713);
nand UO_728 (O_728,N_9969,N_7532);
and UO_729 (O_729,N_9398,N_7595);
or UO_730 (O_730,N_7750,N_9314);
nand UO_731 (O_731,N_7756,N_8965);
nor UO_732 (O_732,N_8423,N_8448);
and UO_733 (O_733,N_9772,N_8964);
nand UO_734 (O_734,N_8578,N_9714);
nor UO_735 (O_735,N_8063,N_8560);
xnor UO_736 (O_736,N_9544,N_8974);
and UO_737 (O_737,N_9057,N_9630);
or UO_738 (O_738,N_9546,N_7921);
nand UO_739 (O_739,N_8860,N_8505);
and UO_740 (O_740,N_8881,N_9392);
or UO_741 (O_741,N_7615,N_8146);
nand UO_742 (O_742,N_9500,N_7590);
or UO_743 (O_743,N_9246,N_9348);
or UO_744 (O_744,N_7923,N_7644);
and UO_745 (O_745,N_9990,N_8775);
nand UO_746 (O_746,N_8342,N_8137);
or UO_747 (O_747,N_8684,N_9558);
and UO_748 (O_748,N_7725,N_7578);
or UO_749 (O_749,N_9735,N_8158);
nand UO_750 (O_750,N_8886,N_8150);
nor UO_751 (O_751,N_8690,N_8116);
and UO_752 (O_752,N_8153,N_8371);
nor UO_753 (O_753,N_8320,N_7517);
nor UO_754 (O_754,N_9866,N_8653);
or UO_755 (O_755,N_9719,N_9325);
and UO_756 (O_756,N_9165,N_7664);
and UO_757 (O_757,N_9282,N_7566);
nor UO_758 (O_758,N_9779,N_8328);
nor UO_759 (O_759,N_9156,N_8710);
and UO_760 (O_760,N_7623,N_8169);
or UO_761 (O_761,N_8000,N_9466);
or UO_762 (O_762,N_9148,N_9371);
or UO_763 (O_763,N_7935,N_7682);
nand UO_764 (O_764,N_8253,N_9144);
or UO_765 (O_765,N_9240,N_8373);
or UO_766 (O_766,N_9664,N_8816);
or UO_767 (O_767,N_9353,N_7515);
or UO_768 (O_768,N_7901,N_7982);
or UO_769 (O_769,N_7977,N_7886);
and UO_770 (O_770,N_9624,N_9227);
nand UO_771 (O_771,N_8220,N_9598);
nand UO_772 (O_772,N_8827,N_8277);
nor UO_773 (O_773,N_9118,N_8695);
nor UO_774 (O_774,N_9661,N_9475);
nor UO_775 (O_775,N_8174,N_7816);
nor UO_776 (O_776,N_9288,N_7837);
nor UO_777 (O_777,N_8144,N_8445);
or UO_778 (O_778,N_9096,N_8236);
and UO_779 (O_779,N_9667,N_8826);
nor UO_780 (O_780,N_9541,N_8266);
or UO_781 (O_781,N_7610,N_9078);
nand UO_782 (O_782,N_8011,N_7551);
nand UO_783 (O_783,N_9454,N_7954);
nor UO_784 (O_784,N_8025,N_7864);
nor UO_785 (O_785,N_8496,N_9831);
nand UO_786 (O_786,N_8518,N_9815);
nor UO_787 (O_787,N_9034,N_8993);
and UO_788 (O_788,N_9264,N_9102);
or UO_789 (O_789,N_9612,N_9014);
nor UO_790 (O_790,N_8937,N_8092);
and UO_791 (O_791,N_8943,N_9659);
nor UO_792 (O_792,N_8149,N_8248);
nand UO_793 (O_793,N_8078,N_7985);
nand UO_794 (O_794,N_7949,N_7830);
or UO_795 (O_795,N_7622,N_9878);
and UO_796 (O_796,N_8075,N_9434);
or UO_797 (O_797,N_9826,N_9947);
and UO_798 (O_798,N_7839,N_8482);
nor UO_799 (O_799,N_9597,N_7659);
or UO_800 (O_800,N_7967,N_8992);
xnor UO_801 (O_801,N_7867,N_9839);
or UO_802 (O_802,N_9457,N_8458);
and UO_803 (O_803,N_9296,N_8337);
nand UO_804 (O_804,N_9381,N_9467);
or UO_805 (O_805,N_8449,N_7571);
xor UO_806 (O_806,N_8311,N_9275);
and UO_807 (O_807,N_8297,N_9323);
nand UO_808 (O_808,N_8105,N_9365);
nand UO_809 (O_809,N_7649,N_9648);
nor UO_810 (O_810,N_8009,N_8228);
and UO_811 (O_811,N_7809,N_8082);
or UO_812 (O_812,N_9712,N_7694);
or UO_813 (O_813,N_8616,N_9004);
or UO_814 (O_814,N_8708,N_7852);
nor UO_815 (O_815,N_7854,N_8026);
nor UO_816 (O_816,N_8761,N_9189);
nand UO_817 (O_817,N_8350,N_8126);
nor UO_818 (O_818,N_9653,N_9501);
nand UO_819 (O_819,N_8687,N_9032);
nand UO_820 (O_820,N_7797,N_8579);
or UO_821 (O_821,N_9945,N_8298);
or UO_822 (O_822,N_9555,N_9289);
nor UO_823 (O_823,N_8156,N_8951);
or UO_824 (O_824,N_9182,N_8522);
and UO_825 (O_825,N_7815,N_8461);
and UO_826 (O_826,N_8030,N_8173);
nor UO_827 (O_827,N_8913,N_7933);
nor UO_828 (O_828,N_8338,N_8098);
nand UO_829 (O_829,N_9175,N_8242);
or UO_830 (O_830,N_9647,N_9977);
nand UO_831 (O_831,N_9347,N_9766);
or UO_832 (O_832,N_8249,N_9781);
nand UO_833 (O_833,N_8524,N_9819);
nor UO_834 (O_834,N_8395,N_8470);
or UO_835 (O_835,N_9394,N_8035);
or UO_836 (O_836,N_7503,N_8336);
and UO_837 (O_837,N_9991,N_9749);
nand UO_838 (O_838,N_8840,N_9907);
nor UO_839 (O_839,N_8130,N_9299);
and UO_840 (O_840,N_8858,N_9407);
or UO_841 (O_841,N_9164,N_7973);
and UO_842 (O_842,N_7762,N_9835);
nor UO_843 (O_843,N_8090,N_9545);
or UO_844 (O_844,N_8066,N_8397);
or UO_845 (O_845,N_8855,N_7658);
and UO_846 (O_846,N_9046,N_9876);
nand UO_847 (O_847,N_9607,N_9700);
and UO_848 (O_848,N_8053,N_7771);
or UO_849 (O_849,N_8844,N_8229);
nor UO_850 (O_850,N_8626,N_7671);
nor UO_851 (O_851,N_9783,N_8674);
and UO_852 (O_852,N_8558,N_8925);
nor UO_853 (O_853,N_9100,N_8466);
and UO_854 (O_854,N_7834,N_7700);
or UO_855 (O_855,N_8874,N_7796);
nor UO_856 (O_856,N_8196,N_8401);
nor UO_857 (O_857,N_9209,N_7760);
nand UO_858 (O_858,N_7541,N_8997);
nor UO_859 (O_859,N_7971,N_9572);
nor UO_860 (O_860,N_9389,N_9798);
nor UO_861 (O_861,N_8575,N_8803);
and UO_862 (O_862,N_8676,N_9690);
or UO_863 (O_863,N_8108,N_7624);
nor UO_864 (O_864,N_7904,N_9085);
nand UO_865 (O_865,N_9459,N_8363);
or UO_866 (O_866,N_7547,N_8611);
nand UO_867 (O_867,N_8016,N_8161);
nand UO_868 (O_868,N_7592,N_9608);
nor UO_869 (O_869,N_8446,N_8525);
nor UO_870 (O_870,N_9935,N_9980);
nand UO_871 (O_871,N_9674,N_9111);
xnor UO_872 (O_872,N_9225,N_8632);
and UO_873 (O_873,N_8289,N_9968);
nand UO_874 (O_874,N_8295,N_9183);
nand UO_875 (O_875,N_9428,N_9673);
nand UO_876 (O_876,N_8631,N_8226);
and UO_877 (O_877,N_8854,N_9877);
nor UO_878 (O_878,N_9119,N_8138);
nor UO_879 (O_879,N_8001,N_8580);
and UO_880 (O_880,N_9662,N_7766);
nand UO_881 (O_881,N_8400,N_8552);
nor UO_882 (O_882,N_9052,N_8741);
nor UO_883 (O_883,N_9709,N_9088);
nor UO_884 (O_884,N_8788,N_9535);
nor UO_885 (O_885,N_9964,N_8280);
or UO_886 (O_886,N_7863,N_8319);
nand UO_887 (O_887,N_8031,N_7581);
or UO_888 (O_888,N_8175,N_9628);
and UO_889 (O_889,N_8810,N_8024);
and UO_890 (O_890,N_8952,N_9322);
or UO_891 (O_891,N_9267,N_8367);
nand UO_892 (O_892,N_8478,N_8824);
nand UO_893 (O_893,N_8990,N_9910);
nor UO_894 (O_894,N_7729,N_8794);
nand UO_895 (O_895,N_9609,N_9358);
nor UO_896 (O_896,N_9579,N_7708);
nor UO_897 (O_897,N_7545,N_8034);
nor UO_898 (O_898,N_8047,N_7930);
or UO_899 (O_899,N_8049,N_8924);
nor UO_900 (O_900,N_9993,N_8953);
nand UO_901 (O_901,N_8970,N_9698);
nand UO_902 (O_902,N_8613,N_8691);
and UO_903 (O_903,N_8115,N_7616);
nor UO_904 (O_904,N_8245,N_8866);
nor UO_905 (O_905,N_7927,N_9881);
and UO_906 (O_906,N_9736,N_7840);
or UO_907 (O_907,N_8263,N_8194);
and UO_908 (O_908,N_8042,N_9070);
nor UO_909 (O_909,N_8017,N_7654);
and UO_910 (O_910,N_9147,N_7984);
nor UO_911 (O_911,N_7784,N_9578);
nand UO_912 (O_912,N_9222,N_7832);
or UO_913 (O_913,N_9252,N_8903);
and UO_914 (O_914,N_7769,N_8321);
nand UO_915 (O_915,N_8856,N_9840);
nand UO_916 (O_916,N_8852,N_9380);
nand UO_917 (O_917,N_9115,N_8121);
xnor UO_918 (O_918,N_8509,N_9571);
or UO_919 (O_919,N_9843,N_7672);
and UO_920 (O_920,N_8576,N_9632);
or UO_921 (O_921,N_8562,N_8015);
or UO_922 (O_922,N_9603,N_9510);
and UO_923 (O_923,N_8772,N_9053);
or UO_924 (O_924,N_9041,N_9079);
nand UO_925 (O_925,N_9072,N_9329);
or UO_926 (O_926,N_8661,N_8040);
nand UO_927 (O_927,N_8428,N_9886);
and UO_928 (O_928,N_7952,N_9640);
nand UO_929 (O_929,N_9550,N_8971);
nand UO_930 (O_930,N_9523,N_9387);
or UO_931 (O_931,N_8241,N_9254);
nor UO_932 (O_932,N_9795,N_8416);
nor UO_933 (O_933,N_8399,N_8995);
nor UO_934 (O_934,N_9054,N_9109);
and UO_935 (O_935,N_8100,N_9226);
nand UO_936 (O_936,N_8767,N_8164);
nor UO_937 (O_937,N_9292,N_8512);
nor UO_938 (O_938,N_8502,N_8244);
and UO_939 (O_939,N_8020,N_8936);
or UO_940 (O_940,N_9473,N_8335);
nand UO_941 (O_941,N_8424,N_9634);
and UO_942 (O_942,N_8152,N_9177);
nand UO_943 (O_943,N_9152,N_8918);
nand UO_944 (O_944,N_9038,N_9196);
nor UO_945 (O_945,N_7674,N_8662);
nor UO_946 (O_946,N_9207,N_7960);
nand UO_947 (O_947,N_8605,N_9330);
and UO_948 (O_948,N_7884,N_9276);
nor UO_949 (O_949,N_8583,N_9097);
or UO_950 (O_950,N_8369,N_7523);
nand UO_951 (O_951,N_9011,N_7573);
nor UO_952 (O_952,N_8471,N_8343);
nor UO_953 (O_953,N_7902,N_9748);
xor UO_954 (O_954,N_8818,N_9300);
and UO_955 (O_955,N_8477,N_9625);
nand UO_956 (O_956,N_8112,N_9885);
nor UO_957 (O_957,N_7504,N_7974);
nor UO_958 (O_958,N_9103,N_9170);
and UO_959 (O_959,N_8305,N_7942);
nor UO_960 (O_960,N_8165,N_8185);
nand UO_961 (O_961,N_9089,N_9508);
and UO_962 (O_962,N_8497,N_9707);
or UO_963 (O_963,N_7717,N_8374);
nor UO_964 (O_964,N_8281,N_8729);
nor UO_965 (O_965,N_8362,N_9695);
nor UO_966 (O_966,N_9463,N_8718);
and UO_967 (O_967,N_9926,N_9412);
or UO_968 (O_968,N_8590,N_8345);
nor UO_969 (O_969,N_8504,N_8527);
or UO_970 (O_970,N_9228,N_8773);
nand UO_971 (O_971,N_7701,N_9654);
nor UO_972 (O_972,N_7843,N_8822);
nand UO_973 (O_973,N_8481,N_9723);
nand UO_974 (O_974,N_7600,N_8929);
or UO_975 (O_975,N_8274,N_9509);
nor UO_976 (O_976,N_9243,N_9062);
nand UO_977 (O_977,N_7666,N_7617);
and UO_978 (O_978,N_9433,N_8231);
nand UO_979 (O_979,N_9525,N_9660);
nor UO_980 (O_980,N_9912,N_9000);
nor UO_981 (O_981,N_9319,N_7684);
and UO_982 (O_982,N_9110,N_8799);
or UO_983 (O_983,N_8119,N_9369);
nor UO_984 (O_984,N_9539,N_7937);
and UO_985 (O_985,N_8666,N_9404);
nor UO_986 (O_986,N_8418,N_7861);
nand UO_987 (O_987,N_8259,N_7743);
nor UO_988 (O_988,N_9101,N_8577);
nor UO_989 (O_989,N_8141,N_8084);
or UO_990 (O_990,N_8901,N_9704);
nor UO_991 (O_991,N_8705,N_9919);
nor UO_992 (O_992,N_9352,N_8324);
and UO_993 (O_993,N_9725,N_9214);
or UO_994 (O_994,N_9796,N_9813);
nand UO_995 (O_995,N_9994,N_8357);
or UO_996 (O_996,N_7870,N_7879);
and UO_997 (O_997,N_9978,N_9218);
nor UO_998 (O_998,N_7546,N_9385);
nor UO_999 (O_999,N_9900,N_9856);
nor UO_1000 (O_1000,N_8290,N_9255);
nand UO_1001 (O_1001,N_7844,N_7903);
nand UO_1002 (O_1002,N_8168,N_7842);
nand UO_1003 (O_1003,N_7825,N_8157);
nand UO_1004 (O_1004,N_7652,N_7707);
nand UO_1005 (O_1005,N_9280,N_8451);
nand UO_1006 (O_1006,N_7958,N_7914);
nor UO_1007 (O_1007,N_8398,N_7764);
nand UO_1008 (O_1008,N_8902,N_9220);
nor UO_1009 (O_1009,N_9327,N_9496);
and UO_1010 (O_1010,N_9074,N_9961);
xnor UO_1011 (O_1011,N_8635,N_8833);
nand UO_1012 (O_1012,N_8570,N_7685);
or UO_1013 (O_1013,N_9642,N_8839);
nand UO_1014 (O_1014,N_8547,N_7781);
nor UO_1015 (O_1015,N_9490,N_7568);
or UO_1016 (O_1016,N_8819,N_9963);
nor UO_1017 (O_1017,N_8288,N_8113);
nand UO_1018 (O_1018,N_8243,N_9341);
nor UO_1019 (O_1019,N_9498,N_8475);
nand UO_1020 (O_1020,N_7848,N_8984);
nor UO_1021 (O_1021,N_8837,N_8421);
and UO_1022 (O_1022,N_8586,N_9536);
nand UO_1023 (O_1023,N_7737,N_9852);
and UO_1024 (O_1024,N_9453,N_9161);
or UO_1025 (O_1025,N_9875,N_8835);
and UO_1026 (O_1026,N_9460,N_9580);
nand UO_1027 (O_1027,N_9427,N_9887);
nor UO_1028 (O_1028,N_9335,N_8668);
or UO_1029 (O_1029,N_8724,N_8314);
nor UO_1030 (O_1030,N_8420,N_7890);
or UO_1031 (O_1031,N_9691,N_9384);
nand UO_1032 (O_1032,N_8549,N_8602);
nand UO_1033 (O_1033,N_9513,N_7637);
or UO_1034 (O_1034,N_8557,N_8877);
nor UO_1035 (O_1035,N_8757,N_9821);
nand UO_1036 (O_1036,N_7538,N_8441);
or UO_1037 (O_1037,N_9799,N_8658);
and UO_1038 (O_1038,N_8539,N_8506);
nand UO_1039 (O_1039,N_9163,N_8240);
and UO_1040 (O_1040,N_7500,N_8699);
and UO_1041 (O_1041,N_7872,N_8412);
or UO_1042 (O_1042,N_7626,N_9933);
nand UO_1043 (O_1043,N_8468,N_8360);
or UO_1044 (O_1044,N_8636,N_8915);
nor UO_1045 (O_1045,N_9986,N_8163);
and UO_1046 (O_1046,N_8980,N_7680);
nand UO_1047 (O_1047,N_8714,N_8160);
nand UO_1048 (O_1048,N_9261,N_9732);
or UO_1049 (O_1049,N_8867,N_9587);
and UO_1050 (O_1050,N_9894,N_9386);
nor UO_1051 (O_1051,N_7711,N_9967);
xor UO_1052 (O_1052,N_8331,N_8029);
or UO_1053 (O_1053,N_8681,N_9438);
nor UO_1054 (O_1054,N_7997,N_7992);
nand UO_1055 (O_1055,N_9021,N_9702);
or UO_1056 (O_1056,N_9145,N_9626);
nor UO_1057 (O_1057,N_9092,N_8764);
and UO_1058 (O_1058,N_9269,N_9497);
nor UO_1059 (O_1059,N_9081,N_7786);
and UO_1060 (O_1060,N_7913,N_8079);
and UO_1061 (O_1061,N_7819,N_7539);
or UO_1062 (O_1062,N_9208,N_8664);
nor UO_1063 (O_1063,N_9955,N_8928);
or UO_1064 (O_1064,N_9008,N_9417);
or UO_1065 (O_1065,N_9792,N_7946);
nand UO_1066 (O_1066,N_9596,N_8815);
nand UO_1067 (O_1067,N_9652,N_9552);
or UO_1068 (O_1068,N_7501,N_7632);
nor UO_1069 (O_1069,N_8264,N_8114);
nor UO_1070 (O_1070,N_7507,N_8284);
nand UO_1071 (O_1071,N_8285,N_9904);
nor UO_1072 (O_1072,N_9917,N_9258);
nand UO_1073 (O_1073,N_7525,N_8221);
or UO_1074 (O_1074,N_8327,N_8969);
nor UO_1075 (O_1075,N_8386,N_9908);
nand UO_1076 (O_1076,N_8133,N_9737);
or UO_1077 (O_1077,N_7530,N_8462);
or UO_1078 (O_1078,N_9236,N_7943);
nand UO_1079 (O_1079,N_7868,N_7951);
and UO_1080 (O_1080,N_7835,N_8432);
xnor UO_1081 (O_1081,N_8823,N_9952);
or UO_1082 (O_1082,N_8282,N_8649);
nand UO_1083 (O_1083,N_9446,N_9614);
and UO_1084 (O_1084,N_9293,N_9676);
and UO_1085 (O_1085,N_8793,N_9858);
nor UO_1086 (O_1086,N_8534,N_7894);
nor UO_1087 (O_1087,N_8942,N_9666);
nand UO_1088 (O_1088,N_8754,N_9462);
and UO_1089 (O_1089,N_7991,N_9863);
or UO_1090 (O_1090,N_7970,N_8791);
nor UO_1091 (O_1091,N_9974,N_9971);
nor UO_1092 (O_1092,N_8272,N_8563);
nor UO_1093 (O_1093,N_8956,N_8349);
or UO_1094 (O_1094,N_9133,N_8972);
and UO_1095 (O_1095,N_7569,N_7721);
nand UO_1096 (O_1096,N_9619,N_8883);
nor UO_1097 (O_1097,N_9954,N_9670);
and UO_1098 (O_1098,N_7792,N_8573);
nor UO_1099 (O_1099,N_8800,N_9105);
nand UO_1100 (O_1100,N_9565,N_9751);
xor UO_1101 (O_1101,N_9505,N_9705);
nand UO_1102 (O_1102,N_9931,N_8402);
and UO_1103 (O_1103,N_8798,N_9420);
and UO_1104 (O_1104,N_8619,N_8476);
nor UO_1105 (O_1105,N_9771,N_9013);
nor UO_1106 (O_1106,N_9094,N_7540);
and UO_1107 (O_1107,N_7912,N_7931);
or UO_1108 (O_1108,N_9415,N_8454);
nand UO_1109 (O_1109,N_7529,N_7679);
nand UO_1110 (O_1110,N_8960,N_7505);
or UO_1111 (O_1111,N_8989,N_9331);
nor UO_1112 (O_1112,N_7918,N_8618);
or UO_1113 (O_1113,N_8947,N_9822);
nor UO_1114 (O_1114,N_7939,N_8529);
nand UO_1115 (O_1115,N_8659,N_9916);
or UO_1116 (O_1116,N_8046,N_9401);
or UO_1117 (O_1117,N_9028,N_8864);
or UO_1118 (O_1118,N_8442,N_8747);
nand UO_1119 (O_1119,N_9400,N_8317);
nand UO_1120 (O_1120,N_8693,N_8979);
nor UO_1121 (O_1121,N_7768,N_9722);
nand UO_1122 (O_1122,N_8312,N_8863);
nand UO_1123 (O_1123,N_7634,N_8495);
or UO_1124 (O_1124,N_9593,N_9340);
nor UO_1125 (O_1125,N_9531,N_9372);
or UO_1126 (O_1126,N_8760,N_7524);
and UO_1127 (O_1127,N_9095,N_7785);
and UO_1128 (O_1128,N_9022,N_7841);
and UO_1129 (O_1129,N_8484,N_9031);
and UO_1130 (O_1130,N_9162,N_8368);
nand UO_1131 (O_1131,N_8841,N_7808);
nand UO_1132 (O_1132,N_9972,N_9807);
and UO_1133 (O_1133,N_9599,N_9515);
or UO_1134 (O_1134,N_8341,N_8830);
nand UO_1135 (O_1135,N_9024,N_8766);
or UO_1136 (O_1136,N_9437,N_8675);
and UO_1137 (O_1137,N_9934,N_7853);
nor UO_1138 (O_1138,N_9084,N_8849);
and UO_1139 (O_1139,N_8222,N_9687);
nor UO_1140 (O_1140,N_8750,N_9202);
and UO_1141 (O_1141,N_8753,N_8917);
and UO_1142 (O_1142,N_8933,N_8660);
and UO_1143 (O_1143,N_7858,N_9962);
nor UO_1144 (O_1144,N_7906,N_8770);
or UO_1145 (O_1145,N_7596,N_9200);
or UO_1146 (O_1146,N_8961,N_8093);
nand UO_1147 (O_1147,N_9278,N_9006);
nand UO_1148 (O_1148,N_9244,N_9337);
nor UO_1149 (O_1149,N_7642,N_9122);
nand UO_1150 (O_1150,N_7979,N_9368);
nand UO_1151 (O_1151,N_8790,N_8111);
nor UO_1152 (O_1152,N_8893,N_8293);
nor UO_1153 (O_1153,N_8225,N_9594);
nand UO_1154 (O_1154,N_7577,N_7976);
or UO_1155 (O_1155,N_8076,N_8528);
nor UO_1156 (O_1156,N_9083,N_9992);
or UO_1157 (O_1157,N_9758,N_9984);
or UO_1158 (O_1158,N_7691,N_9750);
and UO_1159 (O_1159,N_8375,N_8202);
or UO_1160 (O_1160,N_9233,N_9211);
nor UO_1161 (O_1161,N_8963,N_8538);
nand UO_1162 (O_1162,N_7817,N_7831);
nand UO_1163 (O_1163,N_7663,N_8348);
or UO_1164 (O_1164,N_7732,N_9026);
or UO_1165 (O_1165,N_7665,N_8889);
or UO_1166 (O_1166,N_9310,N_9797);
nor UO_1167 (O_1167,N_7554,N_7533);
or UO_1168 (O_1168,N_8419,N_8949);
nor UO_1169 (O_1169,N_9778,N_9499);
and UO_1170 (O_1170,N_9943,N_7900);
xor UO_1171 (O_1171,N_8749,N_9959);
nor UO_1172 (O_1172,N_8069,N_7932);
xnor UO_1173 (O_1173,N_7542,N_8316);
and UO_1174 (O_1174,N_9480,N_9066);
or UO_1175 (O_1175,N_7881,N_8614);
or UO_1176 (O_1176,N_9976,N_7519);
and UO_1177 (O_1177,N_7586,N_9560);
and UO_1178 (O_1178,N_9559,N_8594);
or UO_1179 (O_1179,N_8677,N_9528);
and UO_1180 (O_1180,N_9285,N_7883);
nand UO_1181 (O_1181,N_8792,N_8898);
nor UO_1182 (O_1182,N_8323,N_8033);
or UO_1183 (O_1183,N_8878,N_9889);
and UO_1184 (O_1184,N_8469,N_7940);
or UO_1185 (O_1185,N_9020,N_9701);
xnor UO_1186 (O_1186,N_9411,N_8388);
and UO_1187 (O_1187,N_7850,N_9350);
nand UO_1188 (O_1188,N_7845,N_7876);
and UO_1189 (O_1189,N_8410,N_8239);
nor UO_1190 (O_1190,N_9871,N_9940);
nand UO_1191 (O_1191,N_9367,N_8072);
nor UO_1192 (O_1192,N_9413,N_7941);
nand UO_1193 (O_1193,N_9861,N_8404);
or UO_1194 (O_1194,N_7535,N_9047);
nor UO_1195 (O_1195,N_9478,N_8498);
and UO_1196 (O_1196,N_8746,N_9393);
nand UO_1197 (O_1197,N_8473,N_8811);
nand UO_1198 (O_1198,N_9359,N_9996);
nor UO_1199 (O_1199,N_8006,N_9481);
and UO_1200 (O_1200,N_8103,N_8444);
nor UO_1201 (O_1201,N_8640,N_9355);
nand UO_1202 (O_1202,N_9538,N_7794);
xnor UO_1203 (O_1203,N_9173,N_8572);
or UO_1204 (O_1204,N_8002,N_8500);
xor UO_1205 (O_1205,N_8501,N_8200);
and UO_1206 (O_1206,N_7574,N_9068);
nor UO_1207 (O_1207,N_9979,N_7620);
and UO_1208 (O_1208,N_9610,N_9363);
nand UO_1209 (O_1209,N_7621,N_9738);
or UO_1210 (O_1210,N_8499,N_9720);
nor UO_1211 (O_1211,N_9045,N_8927);
nor UO_1212 (O_1212,N_8313,N_9290);
and UO_1213 (O_1213,N_9893,N_8459);
nand UO_1214 (O_1214,N_8088,N_7514);
and UO_1215 (O_1215,N_7925,N_9869);
nor UO_1216 (O_1216,N_9297,N_8897);
nand UO_1217 (O_1217,N_8230,N_8782);
and UO_1218 (O_1218,N_9998,N_8237);
nor UO_1219 (O_1219,N_9315,N_9658);
nor UO_1220 (O_1220,N_7878,N_9679);
nand UO_1221 (O_1221,N_8208,N_7859);
nor UO_1222 (O_1222,N_8540,N_8106);
and UO_1223 (O_1223,N_7558,N_8899);
and UO_1224 (O_1224,N_9345,N_7980);
nor UO_1225 (O_1225,N_8129,N_7916);
or UO_1226 (O_1226,N_9584,N_9279);
nand UO_1227 (O_1227,N_9366,N_9012);
nor UO_1228 (O_1228,N_7777,N_9507);
and UO_1229 (O_1229,N_7559,N_8110);
or UO_1230 (O_1230,N_9576,N_7802);
nor UO_1231 (O_1231,N_8303,N_8065);
or UO_1232 (O_1232,N_9354,N_8003);
nand UO_1233 (O_1233,N_8737,N_9126);
nor UO_1234 (O_1234,N_8526,N_9250);
or UO_1235 (O_1235,N_9694,N_9556);
nor UO_1236 (O_1236,N_8665,N_9981);
or UO_1237 (O_1237,N_8479,N_8436);
and UO_1238 (O_1238,N_7591,N_7821);
and UO_1239 (O_1239,N_9328,N_8922);
or UO_1240 (O_1240,N_9339,N_9903);
or UO_1241 (O_1241,N_8060,N_8742);
nand UO_1242 (O_1242,N_9223,N_8287);
nor UO_1243 (O_1243,N_8641,N_8634);
nand UO_1244 (O_1244,N_8392,N_8755);
nand UO_1245 (O_1245,N_7888,N_9902);
nor UO_1246 (O_1246,N_7719,N_8438);
and UO_1247 (O_1247,N_8389,N_9864);
nor UO_1248 (O_1248,N_8159,N_7678);
and UO_1249 (O_1249,N_9897,N_8218);
nor UO_1250 (O_1250,N_7575,N_8842);
or UO_1251 (O_1251,N_9043,N_9352);
or UO_1252 (O_1252,N_8674,N_8044);
nor UO_1253 (O_1253,N_7701,N_7613);
nor UO_1254 (O_1254,N_9007,N_7936);
nand UO_1255 (O_1255,N_7703,N_7908);
nor UO_1256 (O_1256,N_9535,N_8715);
or UO_1257 (O_1257,N_9435,N_7972);
and UO_1258 (O_1258,N_8242,N_8541);
nor UO_1259 (O_1259,N_8478,N_9031);
nand UO_1260 (O_1260,N_8937,N_9991);
or UO_1261 (O_1261,N_7537,N_9025);
or UO_1262 (O_1262,N_8406,N_8097);
nand UO_1263 (O_1263,N_7828,N_7816);
and UO_1264 (O_1264,N_9164,N_8241);
or UO_1265 (O_1265,N_8293,N_9802);
nand UO_1266 (O_1266,N_8875,N_7703);
nand UO_1267 (O_1267,N_9390,N_9734);
nor UO_1268 (O_1268,N_9778,N_9639);
and UO_1269 (O_1269,N_9573,N_9860);
nor UO_1270 (O_1270,N_8318,N_7884);
nand UO_1271 (O_1271,N_8005,N_9261);
and UO_1272 (O_1272,N_9185,N_8120);
or UO_1273 (O_1273,N_7751,N_8274);
and UO_1274 (O_1274,N_8008,N_9521);
nand UO_1275 (O_1275,N_9276,N_9571);
or UO_1276 (O_1276,N_9844,N_8217);
and UO_1277 (O_1277,N_9245,N_9241);
nor UO_1278 (O_1278,N_7930,N_8194);
nand UO_1279 (O_1279,N_7512,N_9158);
nor UO_1280 (O_1280,N_8907,N_9956);
nor UO_1281 (O_1281,N_9961,N_9953);
nor UO_1282 (O_1282,N_7539,N_8676);
nand UO_1283 (O_1283,N_9431,N_9073);
nor UO_1284 (O_1284,N_8647,N_9004);
nor UO_1285 (O_1285,N_8184,N_8994);
or UO_1286 (O_1286,N_8981,N_8081);
or UO_1287 (O_1287,N_8442,N_8735);
nor UO_1288 (O_1288,N_7779,N_8563);
or UO_1289 (O_1289,N_8552,N_9035);
or UO_1290 (O_1290,N_8189,N_7975);
or UO_1291 (O_1291,N_8576,N_7885);
or UO_1292 (O_1292,N_7979,N_9907);
nor UO_1293 (O_1293,N_9589,N_7584);
or UO_1294 (O_1294,N_8931,N_8989);
xnor UO_1295 (O_1295,N_9124,N_9546);
and UO_1296 (O_1296,N_8338,N_8410);
nand UO_1297 (O_1297,N_7588,N_8216);
or UO_1298 (O_1298,N_8053,N_8967);
and UO_1299 (O_1299,N_8808,N_8145);
and UO_1300 (O_1300,N_8071,N_8963);
nand UO_1301 (O_1301,N_9934,N_7510);
nor UO_1302 (O_1302,N_8757,N_9430);
or UO_1303 (O_1303,N_8698,N_7818);
or UO_1304 (O_1304,N_9743,N_8791);
nand UO_1305 (O_1305,N_8443,N_7829);
and UO_1306 (O_1306,N_9614,N_8169);
or UO_1307 (O_1307,N_8921,N_9800);
and UO_1308 (O_1308,N_8229,N_8798);
and UO_1309 (O_1309,N_8468,N_7740);
nand UO_1310 (O_1310,N_9756,N_8555);
nand UO_1311 (O_1311,N_9650,N_8407);
nand UO_1312 (O_1312,N_8463,N_9772);
or UO_1313 (O_1313,N_8899,N_8609);
nor UO_1314 (O_1314,N_9263,N_9352);
and UO_1315 (O_1315,N_7866,N_7521);
nand UO_1316 (O_1316,N_9866,N_9197);
or UO_1317 (O_1317,N_9956,N_8642);
nand UO_1318 (O_1318,N_8882,N_9755);
nand UO_1319 (O_1319,N_9469,N_8772);
or UO_1320 (O_1320,N_8143,N_7597);
nand UO_1321 (O_1321,N_9048,N_9383);
nand UO_1322 (O_1322,N_9467,N_7968);
and UO_1323 (O_1323,N_8319,N_9968);
or UO_1324 (O_1324,N_9268,N_8250);
and UO_1325 (O_1325,N_8578,N_9100);
and UO_1326 (O_1326,N_7592,N_8913);
or UO_1327 (O_1327,N_8746,N_8003);
nor UO_1328 (O_1328,N_8678,N_8388);
and UO_1329 (O_1329,N_8428,N_8476);
nor UO_1330 (O_1330,N_9679,N_8932);
nand UO_1331 (O_1331,N_7856,N_9356);
and UO_1332 (O_1332,N_9687,N_8383);
nor UO_1333 (O_1333,N_8840,N_9979);
or UO_1334 (O_1334,N_9060,N_8306);
and UO_1335 (O_1335,N_8332,N_8859);
or UO_1336 (O_1336,N_9400,N_8242);
nand UO_1337 (O_1337,N_9149,N_9245);
or UO_1338 (O_1338,N_9775,N_8544);
nor UO_1339 (O_1339,N_8776,N_8550);
or UO_1340 (O_1340,N_9880,N_9162);
nand UO_1341 (O_1341,N_7824,N_8032);
nor UO_1342 (O_1342,N_8147,N_7892);
nand UO_1343 (O_1343,N_9014,N_7812);
or UO_1344 (O_1344,N_8024,N_8174);
nand UO_1345 (O_1345,N_8254,N_9376);
or UO_1346 (O_1346,N_7642,N_7706);
and UO_1347 (O_1347,N_8471,N_9859);
or UO_1348 (O_1348,N_8365,N_9603);
nor UO_1349 (O_1349,N_8626,N_7525);
or UO_1350 (O_1350,N_8279,N_8848);
nand UO_1351 (O_1351,N_9539,N_9664);
or UO_1352 (O_1352,N_7568,N_8388);
nor UO_1353 (O_1353,N_8862,N_8934);
or UO_1354 (O_1354,N_8293,N_8309);
and UO_1355 (O_1355,N_8399,N_8852);
and UO_1356 (O_1356,N_8612,N_7833);
nor UO_1357 (O_1357,N_9186,N_8745);
nand UO_1358 (O_1358,N_8896,N_9718);
and UO_1359 (O_1359,N_7651,N_9770);
nand UO_1360 (O_1360,N_9300,N_8707);
nand UO_1361 (O_1361,N_8704,N_9344);
nor UO_1362 (O_1362,N_8196,N_9304);
and UO_1363 (O_1363,N_8018,N_7882);
or UO_1364 (O_1364,N_8211,N_9015);
nand UO_1365 (O_1365,N_9155,N_8229);
nand UO_1366 (O_1366,N_8228,N_8167);
nand UO_1367 (O_1367,N_9925,N_9578);
nand UO_1368 (O_1368,N_7544,N_7538);
nor UO_1369 (O_1369,N_9255,N_7667);
nor UO_1370 (O_1370,N_8676,N_7874);
nor UO_1371 (O_1371,N_9479,N_9789);
nand UO_1372 (O_1372,N_9477,N_9356);
nand UO_1373 (O_1373,N_9451,N_8103);
and UO_1374 (O_1374,N_8730,N_9395);
nand UO_1375 (O_1375,N_7574,N_7962);
nand UO_1376 (O_1376,N_9713,N_7619);
nand UO_1377 (O_1377,N_8796,N_7533);
nand UO_1378 (O_1378,N_8126,N_9646);
nor UO_1379 (O_1379,N_8207,N_7659);
nand UO_1380 (O_1380,N_8142,N_8754);
nand UO_1381 (O_1381,N_8974,N_8630);
or UO_1382 (O_1382,N_8159,N_8847);
nor UO_1383 (O_1383,N_8602,N_9104);
or UO_1384 (O_1384,N_9199,N_9000);
nand UO_1385 (O_1385,N_8299,N_8129);
or UO_1386 (O_1386,N_8934,N_8218);
or UO_1387 (O_1387,N_9298,N_9047);
and UO_1388 (O_1388,N_7595,N_8242);
nand UO_1389 (O_1389,N_7699,N_7758);
or UO_1390 (O_1390,N_8868,N_8479);
nor UO_1391 (O_1391,N_8488,N_8565);
and UO_1392 (O_1392,N_8709,N_9239);
nor UO_1393 (O_1393,N_9348,N_9113);
nand UO_1394 (O_1394,N_9235,N_9253);
and UO_1395 (O_1395,N_8466,N_9651);
nand UO_1396 (O_1396,N_9987,N_8571);
xor UO_1397 (O_1397,N_8146,N_9026);
nor UO_1398 (O_1398,N_9989,N_8346);
and UO_1399 (O_1399,N_8588,N_9532);
nand UO_1400 (O_1400,N_8417,N_9073);
and UO_1401 (O_1401,N_9989,N_9452);
and UO_1402 (O_1402,N_7870,N_9140);
and UO_1403 (O_1403,N_8507,N_8568);
or UO_1404 (O_1404,N_9209,N_8401);
and UO_1405 (O_1405,N_9919,N_8133);
nand UO_1406 (O_1406,N_8801,N_7814);
nor UO_1407 (O_1407,N_8019,N_8394);
nand UO_1408 (O_1408,N_8856,N_9339);
and UO_1409 (O_1409,N_9616,N_8210);
and UO_1410 (O_1410,N_9015,N_9221);
or UO_1411 (O_1411,N_9022,N_9228);
nor UO_1412 (O_1412,N_7903,N_9775);
and UO_1413 (O_1413,N_7962,N_9323);
nand UO_1414 (O_1414,N_8166,N_9331);
nor UO_1415 (O_1415,N_8367,N_9078);
and UO_1416 (O_1416,N_9072,N_9189);
and UO_1417 (O_1417,N_7899,N_7878);
nor UO_1418 (O_1418,N_8517,N_9508);
nor UO_1419 (O_1419,N_8081,N_9813);
nor UO_1420 (O_1420,N_8706,N_8898);
nand UO_1421 (O_1421,N_8408,N_8426);
nor UO_1422 (O_1422,N_9380,N_8596);
nand UO_1423 (O_1423,N_8871,N_8172);
and UO_1424 (O_1424,N_7737,N_9650);
or UO_1425 (O_1425,N_7598,N_9239);
nand UO_1426 (O_1426,N_8496,N_8350);
nand UO_1427 (O_1427,N_8390,N_8597);
xnor UO_1428 (O_1428,N_9972,N_8432);
nor UO_1429 (O_1429,N_7997,N_8201);
nand UO_1430 (O_1430,N_8800,N_7593);
or UO_1431 (O_1431,N_9972,N_9506);
or UO_1432 (O_1432,N_8727,N_9427);
or UO_1433 (O_1433,N_8812,N_9917);
and UO_1434 (O_1434,N_7651,N_9667);
nor UO_1435 (O_1435,N_7933,N_8367);
nand UO_1436 (O_1436,N_8248,N_8688);
nand UO_1437 (O_1437,N_8612,N_9235);
nor UO_1438 (O_1438,N_9161,N_7685);
nand UO_1439 (O_1439,N_9914,N_9253);
nand UO_1440 (O_1440,N_9552,N_7761);
nand UO_1441 (O_1441,N_8748,N_7919);
and UO_1442 (O_1442,N_8179,N_8449);
nand UO_1443 (O_1443,N_8396,N_9856);
and UO_1444 (O_1444,N_7757,N_9388);
and UO_1445 (O_1445,N_8618,N_9779);
nor UO_1446 (O_1446,N_9605,N_9158);
and UO_1447 (O_1447,N_9957,N_8545);
or UO_1448 (O_1448,N_8766,N_9409);
or UO_1449 (O_1449,N_8282,N_7864);
and UO_1450 (O_1450,N_9997,N_8201);
or UO_1451 (O_1451,N_7703,N_7683);
or UO_1452 (O_1452,N_8014,N_8491);
nor UO_1453 (O_1453,N_8497,N_9910);
or UO_1454 (O_1454,N_8393,N_8199);
nor UO_1455 (O_1455,N_9395,N_8563);
nand UO_1456 (O_1456,N_7512,N_9347);
nor UO_1457 (O_1457,N_9339,N_8819);
and UO_1458 (O_1458,N_9300,N_8937);
nand UO_1459 (O_1459,N_9513,N_9895);
and UO_1460 (O_1460,N_7858,N_9916);
and UO_1461 (O_1461,N_8820,N_9641);
or UO_1462 (O_1462,N_8236,N_9303);
or UO_1463 (O_1463,N_8786,N_8999);
and UO_1464 (O_1464,N_7525,N_9103);
and UO_1465 (O_1465,N_8215,N_8000);
and UO_1466 (O_1466,N_8118,N_9698);
nor UO_1467 (O_1467,N_8467,N_7542);
xor UO_1468 (O_1468,N_9863,N_8184);
nand UO_1469 (O_1469,N_9541,N_8055);
or UO_1470 (O_1470,N_8434,N_8922);
or UO_1471 (O_1471,N_9985,N_8588);
nand UO_1472 (O_1472,N_9895,N_7948);
nor UO_1473 (O_1473,N_8746,N_7848);
nor UO_1474 (O_1474,N_8506,N_8705);
nand UO_1475 (O_1475,N_9725,N_9106);
nor UO_1476 (O_1476,N_9488,N_7639);
nand UO_1477 (O_1477,N_8876,N_7923);
nand UO_1478 (O_1478,N_7979,N_8405);
nand UO_1479 (O_1479,N_9890,N_9892);
xnor UO_1480 (O_1480,N_8414,N_9800);
xnor UO_1481 (O_1481,N_9916,N_9522);
and UO_1482 (O_1482,N_9358,N_7509);
xnor UO_1483 (O_1483,N_8275,N_9090);
and UO_1484 (O_1484,N_9437,N_8153);
xor UO_1485 (O_1485,N_9367,N_9383);
or UO_1486 (O_1486,N_9568,N_7812);
nor UO_1487 (O_1487,N_9451,N_8392);
and UO_1488 (O_1488,N_7882,N_9652);
and UO_1489 (O_1489,N_9811,N_8510);
nor UO_1490 (O_1490,N_9366,N_8446);
nand UO_1491 (O_1491,N_8196,N_8169);
nor UO_1492 (O_1492,N_7513,N_8389);
nand UO_1493 (O_1493,N_9085,N_9200);
nand UO_1494 (O_1494,N_9129,N_8058);
or UO_1495 (O_1495,N_9888,N_9569);
nor UO_1496 (O_1496,N_9942,N_9902);
nor UO_1497 (O_1497,N_8280,N_8844);
nor UO_1498 (O_1498,N_8484,N_9166);
xor UO_1499 (O_1499,N_7935,N_8433);
endmodule