module basic_5000_50000_5000_10_levels_10xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,In_3000,In_3001,In_3002,In_3003,In_3004,In_3005,In_3006,In_3007,In_3008,In_3009,In_3010,In_3011,In_3012,In_3013,In_3014,In_3015,In_3016,In_3017,In_3018,In_3019,In_3020,In_3021,In_3022,In_3023,In_3024,In_3025,In_3026,In_3027,In_3028,In_3029,In_3030,In_3031,In_3032,In_3033,In_3034,In_3035,In_3036,In_3037,In_3038,In_3039,In_3040,In_3041,In_3042,In_3043,In_3044,In_3045,In_3046,In_3047,In_3048,In_3049,In_3050,In_3051,In_3052,In_3053,In_3054,In_3055,In_3056,In_3057,In_3058,In_3059,In_3060,In_3061,In_3062,In_3063,In_3064,In_3065,In_3066,In_3067,In_3068,In_3069,In_3070,In_3071,In_3072,In_3073,In_3074,In_3075,In_3076,In_3077,In_3078,In_3079,In_3080,In_3081,In_3082,In_3083,In_3084,In_3085,In_3086,In_3087,In_3088,In_3089,In_3090,In_3091,In_3092,In_3093,In_3094,In_3095,In_3096,In_3097,In_3098,In_3099,In_3100,In_3101,In_3102,In_3103,In_3104,In_3105,In_3106,In_3107,In_3108,In_3109,In_3110,In_3111,In_3112,In_3113,In_3114,In_3115,In_3116,In_3117,In_3118,In_3119,In_3120,In_3121,In_3122,In_3123,In_3124,In_3125,In_3126,In_3127,In_3128,In_3129,In_3130,In_3131,In_3132,In_3133,In_3134,In_3135,In_3136,In_3137,In_3138,In_3139,In_3140,In_3141,In_3142,In_3143,In_3144,In_3145,In_3146,In_3147,In_3148,In_3149,In_3150,In_3151,In_3152,In_3153,In_3154,In_3155,In_3156,In_3157,In_3158,In_3159,In_3160,In_3161,In_3162,In_3163,In_3164,In_3165,In_3166,In_3167,In_3168,In_3169,In_3170,In_3171,In_3172,In_3173,In_3174,In_3175,In_3176,In_3177,In_3178,In_3179,In_3180,In_3181,In_3182,In_3183,In_3184,In_3185,In_3186,In_3187,In_3188,In_3189,In_3190,In_3191,In_3192,In_3193,In_3194,In_3195,In_3196,In_3197,In_3198,In_3199,In_3200,In_3201,In_3202,In_3203,In_3204,In_3205,In_3206,In_3207,In_3208,In_3209,In_3210,In_3211,In_3212,In_3213,In_3214,In_3215,In_3216,In_3217,In_3218,In_3219,In_3220,In_3221,In_3222,In_3223,In_3224,In_3225,In_3226,In_3227,In_3228,In_3229,In_3230,In_3231,In_3232,In_3233,In_3234,In_3235,In_3236,In_3237,In_3238,In_3239,In_3240,In_3241,In_3242,In_3243,In_3244,In_3245,In_3246,In_3247,In_3248,In_3249,In_3250,In_3251,In_3252,In_3253,In_3254,In_3255,In_3256,In_3257,In_3258,In_3259,In_3260,In_3261,In_3262,In_3263,In_3264,In_3265,In_3266,In_3267,In_3268,In_3269,In_3270,In_3271,In_3272,In_3273,In_3274,In_3275,In_3276,In_3277,In_3278,In_3279,In_3280,In_3281,In_3282,In_3283,In_3284,In_3285,In_3286,In_3287,In_3288,In_3289,In_3290,In_3291,In_3292,In_3293,In_3294,In_3295,In_3296,In_3297,In_3298,In_3299,In_3300,In_3301,In_3302,In_3303,In_3304,In_3305,In_3306,In_3307,In_3308,In_3309,In_3310,In_3311,In_3312,In_3313,In_3314,In_3315,In_3316,In_3317,In_3318,In_3319,In_3320,In_3321,In_3322,In_3323,In_3324,In_3325,In_3326,In_3327,In_3328,In_3329,In_3330,In_3331,In_3332,In_3333,In_3334,In_3335,In_3336,In_3337,In_3338,In_3339,In_3340,In_3341,In_3342,In_3343,In_3344,In_3345,In_3346,In_3347,In_3348,In_3349,In_3350,In_3351,In_3352,In_3353,In_3354,In_3355,In_3356,In_3357,In_3358,In_3359,In_3360,In_3361,In_3362,In_3363,In_3364,In_3365,In_3366,In_3367,In_3368,In_3369,In_3370,In_3371,In_3372,In_3373,In_3374,In_3375,In_3376,In_3377,In_3378,In_3379,In_3380,In_3381,In_3382,In_3383,In_3384,In_3385,In_3386,In_3387,In_3388,In_3389,In_3390,In_3391,In_3392,In_3393,In_3394,In_3395,In_3396,In_3397,In_3398,In_3399,In_3400,In_3401,In_3402,In_3403,In_3404,In_3405,In_3406,In_3407,In_3408,In_3409,In_3410,In_3411,In_3412,In_3413,In_3414,In_3415,In_3416,In_3417,In_3418,In_3419,In_3420,In_3421,In_3422,In_3423,In_3424,In_3425,In_3426,In_3427,In_3428,In_3429,In_3430,In_3431,In_3432,In_3433,In_3434,In_3435,In_3436,In_3437,In_3438,In_3439,In_3440,In_3441,In_3442,In_3443,In_3444,In_3445,In_3446,In_3447,In_3448,In_3449,In_3450,In_3451,In_3452,In_3453,In_3454,In_3455,In_3456,In_3457,In_3458,In_3459,In_3460,In_3461,In_3462,In_3463,In_3464,In_3465,In_3466,In_3467,In_3468,In_3469,In_3470,In_3471,In_3472,In_3473,In_3474,In_3475,In_3476,In_3477,In_3478,In_3479,In_3480,In_3481,In_3482,In_3483,In_3484,In_3485,In_3486,In_3487,In_3488,In_3489,In_3490,In_3491,In_3492,In_3493,In_3494,In_3495,In_3496,In_3497,In_3498,In_3499,In_3500,In_3501,In_3502,In_3503,In_3504,In_3505,In_3506,In_3507,In_3508,In_3509,In_3510,In_3511,In_3512,In_3513,In_3514,In_3515,In_3516,In_3517,In_3518,In_3519,In_3520,In_3521,In_3522,In_3523,In_3524,In_3525,In_3526,In_3527,In_3528,In_3529,In_3530,In_3531,In_3532,In_3533,In_3534,In_3535,In_3536,In_3537,In_3538,In_3539,In_3540,In_3541,In_3542,In_3543,In_3544,In_3545,In_3546,In_3547,In_3548,In_3549,In_3550,In_3551,In_3552,In_3553,In_3554,In_3555,In_3556,In_3557,In_3558,In_3559,In_3560,In_3561,In_3562,In_3563,In_3564,In_3565,In_3566,In_3567,In_3568,In_3569,In_3570,In_3571,In_3572,In_3573,In_3574,In_3575,In_3576,In_3577,In_3578,In_3579,In_3580,In_3581,In_3582,In_3583,In_3584,In_3585,In_3586,In_3587,In_3588,In_3589,In_3590,In_3591,In_3592,In_3593,In_3594,In_3595,In_3596,In_3597,In_3598,In_3599,In_3600,In_3601,In_3602,In_3603,In_3604,In_3605,In_3606,In_3607,In_3608,In_3609,In_3610,In_3611,In_3612,In_3613,In_3614,In_3615,In_3616,In_3617,In_3618,In_3619,In_3620,In_3621,In_3622,In_3623,In_3624,In_3625,In_3626,In_3627,In_3628,In_3629,In_3630,In_3631,In_3632,In_3633,In_3634,In_3635,In_3636,In_3637,In_3638,In_3639,In_3640,In_3641,In_3642,In_3643,In_3644,In_3645,In_3646,In_3647,In_3648,In_3649,In_3650,In_3651,In_3652,In_3653,In_3654,In_3655,In_3656,In_3657,In_3658,In_3659,In_3660,In_3661,In_3662,In_3663,In_3664,In_3665,In_3666,In_3667,In_3668,In_3669,In_3670,In_3671,In_3672,In_3673,In_3674,In_3675,In_3676,In_3677,In_3678,In_3679,In_3680,In_3681,In_3682,In_3683,In_3684,In_3685,In_3686,In_3687,In_3688,In_3689,In_3690,In_3691,In_3692,In_3693,In_3694,In_3695,In_3696,In_3697,In_3698,In_3699,In_3700,In_3701,In_3702,In_3703,In_3704,In_3705,In_3706,In_3707,In_3708,In_3709,In_3710,In_3711,In_3712,In_3713,In_3714,In_3715,In_3716,In_3717,In_3718,In_3719,In_3720,In_3721,In_3722,In_3723,In_3724,In_3725,In_3726,In_3727,In_3728,In_3729,In_3730,In_3731,In_3732,In_3733,In_3734,In_3735,In_3736,In_3737,In_3738,In_3739,In_3740,In_3741,In_3742,In_3743,In_3744,In_3745,In_3746,In_3747,In_3748,In_3749,In_3750,In_3751,In_3752,In_3753,In_3754,In_3755,In_3756,In_3757,In_3758,In_3759,In_3760,In_3761,In_3762,In_3763,In_3764,In_3765,In_3766,In_3767,In_3768,In_3769,In_3770,In_3771,In_3772,In_3773,In_3774,In_3775,In_3776,In_3777,In_3778,In_3779,In_3780,In_3781,In_3782,In_3783,In_3784,In_3785,In_3786,In_3787,In_3788,In_3789,In_3790,In_3791,In_3792,In_3793,In_3794,In_3795,In_3796,In_3797,In_3798,In_3799,In_3800,In_3801,In_3802,In_3803,In_3804,In_3805,In_3806,In_3807,In_3808,In_3809,In_3810,In_3811,In_3812,In_3813,In_3814,In_3815,In_3816,In_3817,In_3818,In_3819,In_3820,In_3821,In_3822,In_3823,In_3824,In_3825,In_3826,In_3827,In_3828,In_3829,In_3830,In_3831,In_3832,In_3833,In_3834,In_3835,In_3836,In_3837,In_3838,In_3839,In_3840,In_3841,In_3842,In_3843,In_3844,In_3845,In_3846,In_3847,In_3848,In_3849,In_3850,In_3851,In_3852,In_3853,In_3854,In_3855,In_3856,In_3857,In_3858,In_3859,In_3860,In_3861,In_3862,In_3863,In_3864,In_3865,In_3866,In_3867,In_3868,In_3869,In_3870,In_3871,In_3872,In_3873,In_3874,In_3875,In_3876,In_3877,In_3878,In_3879,In_3880,In_3881,In_3882,In_3883,In_3884,In_3885,In_3886,In_3887,In_3888,In_3889,In_3890,In_3891,In_3892,In_3893,In_3894,In_3895,In_3896,In_3897,In_3898,In_3899,In_3900,In_3901,In_3902,In_3903,In_3904,In_3905,In_3906,In_3907,In_3908,In_3909,In_3910,In_3911,In_3912,In_3913,In_3914,In_3915,In_3916,In_3917,In_3918,In_3919,In_3920,In_3921,In_3922,In_3923,In_3924,In_3925,In_3926,In_3927,In_3928,In_3929,In_3930,In_3931,In_3932,In_3933,In_3934,In_3935,In_3936,In_3937,In_3938,In_3939,In_3940,In_3941,In_3942,In_3943,In_3944,In_3945,In_3946,In_3947,In_3948,In_3949,In_3950,In_3951,In_3952,In_3953,In_3954,In_3955,In_3956,In_3957,In_3958,In_3959,In_3960,In_3961,In_3962,In_3963,In_3964,In_3965,In_3966,In_3967,In_3968,In_3969,In_3970,In_3971,In_3972,In_3973,In_3974,In_3975,In_3976,In_3977,In_3978,In_3979,In_3980,In_3981,In_3982,In_3983,In_3984,In_3985,In_3986,In_3987,In_3988,In_3989,In_3990,In_3991,In_3992,In_3993,In_3994,In_3995,In_3996,In_3997,In_3998,In_3999,In_4000,In_4001,In_4002,In_4003,In_4004,In_4005,In_4006,In_4007,In_4008,In_4009,In_4010,In_4011,In_4012,In_4013,In_4014,In_4015,In_4016,In_4017,In_4018,In_4019,In_4020,In_4021,In_4022,In_4023,In_4024,In_4025,In_4026,In_4027,In_4028,In_4029,In_4030,In_4031,In_4032,In_4033,In_4034,In_4035,In_4036,In_4037,In_4038,In_4039,In_4040,In_4041,In_4042,In_4043,In_4044,In_4045,In_4046,In_4047,In_4048,In_4049,In_4050,In_4051,In_4052,In_4053,In_4054,In_4055,In_4056,In_4057,In_4058,In_4059,In_4060,In_4061,In_4062,In_4063,In_4064,In_4065,In_4066,In_4067,In_4068,In_4069,In_4070,In_4071,In_4072,In_4073,In_4074,In_4075,In_4076,In_4077,In_4078,In_4079,In_4080,In_4081,In_4082,In_4083,In_4084,In_4085,In_4086,In_4087,In_4088,In_4089,In_4090,In_4091,In_4092,In_4093,In_4094,In_4095,In_4096,In_4097,In_4098,In_4099,In_4100,In_4101,In_4102,In_4103,In_4104,In_4105,In_4106,In_4107,In_4108,In_4109,In_4110,In_4111,In_4112,In_4113,In_4114,In_4115,In_4116,In_4117,In_4118,In_4119,In_4120,In_4121,In_4122,In_4123,In_4124,In_4125,In_4126,In_4127,In_4128,In_4129,In_4130,In_4131,In_4132,In_4133,In_4134,In_4135,In_4136,In_4137,In_4138,In_4139,In_4140,In_4141,In_4142,In_4143,In_4144,In_4145,In_4146,In_4147,In_4148,In_4149,In_4150,In_4151,In_4152,In_4153,In_4154,In_4155,In_4156,In_4157,In_4158,In_4159,In_4160,In_4161,In_4162,In_4163,In_4164,In_4165,In_4166,In_4167,In_4168,In_4169,In_4170,In_4171,In_4172,In_4173,In_4174,In_4175,In_4176,In_4177,In_4178,In_4179,In_4180,In_4181,In_4182,In_4183,In_4184,In_4185,In_4186,In_4187,In_4188,In_4189,In_4190,In_4191,In_4192,In_4193,In_4194,In_4195,In_4196,In_4197,In_4198,In_4199,In_4200,In_4201,In_4202,In_4203,In_4204,In_4205,In_4206,In_4207,In_4208,In_4209,In_4210,In_4211,In_4212,In_4213,In_4214,In_4215,In_4216,In_4217,In_4218,In_4219,In_4220,In_4221,In_4222,In_4223,In_4224,In_4225,In_4226,In_4227,In_4228,In_4229,In_4230,In_4231,In_4232,In_4233,In_4234,In_4235,In_4236,In_4237,In_4238,In_4239,In_4240,In_4241,In_4242,In_4243,In_4244,In_4245,In_4246,In_4247,In_4248,In_4249,In_4250,In_4251,In_4252,In_4253,In_4254,In_4255,In_4256,In_4257,In_4258,In_4259,In_4260,In_4261,In_4262,In_4263,In_4264,In_4265,In_4266,In_4267,In_4268,In_4269,In_4270,In_4271,In_4272,In_4273,In_4274,In_4275,In_4276,In_4277,In_4278,In_4279,In_4280,In_4281,In_4282,In_4283,In_4284,In_4285,In_4286,In_4287,In_4288,In_4289,In_4290,In_4291,In_4292,In_4293,In_4294,In_4295,In_4296,In_4297,In_4298,In_4299,In_4300,In_4301,In_4302,In_4303,In_4304,In_4305,In_4306,In_4307,In_4308,In_4309,In_4310,In_4311,In_4312,In_4313,In_4314,In_4315,In_4316,In_4317,In_4318,In_4319,In_4320,In_4321,In_4322,In_4323,In_4324,In_4325,In_4326,In_4327,In_4328,In_4329,In_4330,In_4331,In_4332,In_4333,In_4334,In_4335,In_4336,In_4337,In_4338,In_4339,In_4340,In_4341,In_4342,In_4343,In_4344,In_4345,In_4346,In_4347,In_4348,In_4349,In_4350,In_4351,In_4352,In_4353,In_4354,In_4355,In_4356,In_4357,In_4358,In_4359,In_4360,In_4361,In_4362,In_4363,In_4364,In_4365,In_4366,In_4367,In_4368,In_4369,In_4370,In_4371,In_4372,In_4373,In_4374,In_4375,In_4376,In_4377,In_4378,In_4379,In_4380,In_4381,In_4382,In_4383,In_4384,In_4385,In_4386,In_4387,In_4388,In_4389,In_4390,In_4391,In_4392,In_4393,In_4394,In_4395,In_4396,In_4397,In_4398,In_4399,In_4400,In_4401,In_4402,In_4403,In_4404,In_4405,In_4406,In_4407,In_4408,In_4409,In_4410,In_4411,In_4412,In_4413,In_4414,In_4415,In_4416,In_4417,In_4418,In_4419,In_4420,In_4421,In_4422,In_4423,In_4424,In_4425,In_4426,In_4427,In_4428,In_4429,In_4430,In_4431,In_4432,In_4433,In_4434,In_4435,In_4436,In_4437,In_4438,In_4439,In_4440,In_4441,In_4442,In_4443,In_4444,In_4445,In_4446,In_4447,In_4448,In_4449,In_4450,In_4451,In_4452,In_4453,In_4454,In_4455,In_4456,In_4457,In_4458,In_4459,In_4460,In_4461,In_4462,In_4463,In_4464,In_4465,In_4466,In_4467,In_4468,In_4469,In_4470,In_4471,In_4472,In_4473,In_4474,In_4475,In_4476,In_4477,In_4478,In_4479,In_4480,In_4481,In_4482,In_4483,In_4484,In_4485,In_4486,In_4487,In_4488,In_4489,In_4490,In_4491,In_4492,In_4493,In_4494,In_4495,In_4496,In_4497,In_4498,In_4499,In_4500,In_4501,In_4502,In_4503,In_4504,In_4505,In_4506,In_4507,In_4508,In_4509,In_4510,In_4511,In_4512,In_4513,In_4514,In_4515,In_4516,In_4517,In_4518,In_4519,In_4520,In_4521,In_4522,In_4523,In_4524,In_4525,In_4526,In_4527,In_4528,In_4529,In_4530,In_4531,In_4532,In_4533,In_4534,In_4535,In_4536,In_4537,In_4538,In_4539,In_4540,In_4541,In_4542,In_4543,In_4544,In_4545,In_4546,In_4547,In_4548,In_4549,In_4550,In_4551,In_4552,In_4553,In_4554,In_4555,In_4556,In_4557,In_4558,In_4559,In_4560,In_4561,In_4562,In_4563,In_4564,In_4565,In_4566,In_4567,In_4568,In_4569,In_4570,In_4571,In_4572,In_4573,In_4574,In_4575,In_4576,In_4577,In_4578,In_4579,In_4580,In_4581,In_4582,In_4583,In_4584,In_4585,In_4586,In_4587,In_4588,In_4589,In_4590,In_4591,In_4592,In_4593,In_4594,In_4595,In_4596,In_4597,In_4598,In_4599,In_4600,In_4601,In_4602,In_4603,In_4604,In_4605,In_4606,In_4607,In_4608,In_4609,In_4610,In_4611,In_4612,In_4613,In_4614,In_4615,In_4616,In_4617,In_4618,In_4619,In_4620,In_4621,In_4622,In_4623,In_4624,In_4625,In_4626,In_4627,In_4628,In_4629,In_4630,In_4631,In_4632,In_4633,In_4634,In_4635,In_4636,In_4637,In_4638,In_4639,In_4640,In_4641,In_4642,In_4643,In_4644,In_4645,In_4646,In_4647,In_4648,In_4649,In_4650,In_4651,In_4652,In_4653,In_4654,In_4655,In_4656,In_4657,In_4658,In_4659,In_4660,In_4661,In_4662,In_4663,In_4664,In_4665,In_4666,In_4667,In_4668,In_4669,In_4670,In_4671,In_4672,In_4673,In_4674,In_4675,In_4676,In_4677,In_4678,In_4679,In_4680,In_4681,In_4682,In_4683,In_4684,In_4685,In_4686,In_4687,In_4688,In_4689,In_4690,In_4691,In_4692,In_4693,In_4694,In_4695,In_4696,In_4697,In_4698,In_4699,In_4700,In_4701,In_4702,In_4703,In_4704,In_4705,In_4706,In_4707,In_4708,In_4709,In_4710,In_4711,In_4712,In_4713,In_4714,In_4715,In_4716,In_4717,In_4718,In_4719,In_4720,In_4721,In_4722,In_4723,In_4724,In_4725,In_4726,In_4727,In_4728,In_4729,In_4730,In_4731,In_4732,In_4733,In_4734,In_4735,In_4736,In_4737,In_4738,In_4739,In_4740,In_4741,In_4742,In_4743,In_4744,In_4745,In_4746,In_4747,In_4748,In_4749,In_4750,In_4751,In_4752,In_4753,In_4754,In_4755,In_4756,In_4757,In_4758,In_4759,In_4760,In_4761,In_4762,In_4763,In_4764,In_4765,In_4766,In_4767,In_4768,In_4769,In_4770,In_4771,In_4772,In_4773,In_4774,In_4775,In_4776,In_4777,In_4778,In_4779,In_4780,In_4781,In_4782,In_4783,In_4784,In_4785,In_4786,In_4787,In_4788,In_4789,In_4790,In_4791,In_4792,In_4793,In_4794,In_4795,In_4796,In_4797,In_4798,In_4799,In_4800,In_4801,In_4802,In_4803,In_4804,In_4805,In_4806,In_4807,In_4808,In_4809,In_4810,In_4811,In_4812,In_4813,In_4814,In_4815,In_4816,In_4817,In_4818,In_4819,In_4820,In_4821,In_4822,In_4823,In_4824,In_4825,In_4826,In_4827,In_4828,In_4829,In_4830,In_4831,In_4832,In_4833,In_4834,In_4835,In_4836,In_4837,In_4838,In_4839,In_4840,In_4841,In_4842,In_4843,In_4844,In_4845,In_4846,In_4847,In_4848,In_4849,In_4850,In_4851,In_4852,In_4853,In_4854,In_4855,In_4856,In_4857,In_4858,In_4859,In_4860,In_4861,In_4862,In_4863,In_4864,In_4865,In_4866,In_4867,In_4868,In_4869,In_4870,In_4871,In_4872,In_4873,In_4874,In_4875,In_4876,In_4877,In_4878,In_4879,In_4880,In_4881,In_4882,In_4883,In_4884,In_4885,In_4886,In_4887,In_4888,In_4889,In_4890,In_4891,In_4892,In_4893,In_4894,In_4895,In_4896,In_4897,In_4898,In_4899,In_4900,In_4901,In_4902,In_4903,In_4904,In_4905,In_4906,In_4907,In_4908,In_4909,In_4910,In_4911,In_4912,In_4913,In_4914,In_4915,In_4916,In_4917,In_4918,In_4919,In_4920,In_4921,In_4922,In_4923,In_4924,In_4925,In_4926,In_4927,In_4928,In_4929,In_4930,In_4931,In_4932,In_4933,In_4934,In_4935,In_4936,In_4937,In_4938,In_4939,In_4940,In_4941,In_4942,In_4943,In_4944,In_4945,In_4946,In_4947,In_4948,In_4949,In_4950,In_4951,In_4952,In_4953,In_4954,In_4955,In_4956,In_4957,In_4958,In_4959,In_4960,In_4961,In_4962,In_4963,In_4964,In_4965,In_4966,In_4967,In_4968,In_4969,In_4970,In_4971,In_4972,In_4973,In_4974,In_4975,In_4976,In_4977,In_4978,In_4979,In_4980,In_4981,In_4982,In_4983,In_4984,In_4985,In_4986,In_4987,In_4988,In_4989,In_4990,In_4991,In_4992,In_4993,In_4994,In_4995,In_4996,In_4997,In_4998,In_4999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499,O_3500,O_3501,O_3502,O_3503,O_3504,O_3505,O_3506,O_3507,O_3508,O_3509,O_3510,O_3511,O_3512,O_3513,O_3514,O_3515,O_3516,O_3517,O_3518,O_3519,O_3520,O_3521,O_3522,O_3523,O_3524,O_3525,O_3526,O_3527,O_3528,O_3529,O_3530,O_3531,O_3532,O_3533,O_3534,O_3535,O_3536,O_3537,O_3538,O_3539,O_3540,O_3541,O_3542,O_3543,O_3544,O_3545,O_3546,O_3547,O_3548,O_3549,O_3550,O_3551,O_3552,O_3553,O_3554,O_3555,O_3556,O_3557,O_3558,O_3559,O_3560,O_3561,O_3562,O_3563,O_3564,O_3565,O_3566,O_3567,O_3568,O_3569,O_3570,O_3571,O_3572,O_3573,O_3574,O_3575,O_3576,O_3577,O_3578,O_3579,O_3580,O_3581,O_3582,O_3583,O_3584,O_3585,O_3586,O_3587,O_3588,O_3589,O_3590,O_3591,O_3592,O_3593,O_3594,O_3595,O_3596,O_3597,O_3598,O_3599,O_3600,O_3601,O_3602,O_3603,O_3604,O_3605,O_3606,O_3607,O_3608,O_3609,O_3610,O_3611,O_3612,O_3613,O_3614,O_3615,O_3616,O_3617,O_3618,O_3619,O_3620,O_3621,O_3622,O_3623,O_3624,O_3625,O_3626,O_3627,O_3628,O_3629,O_3630,O_3631,O_3632,O_3633,O_3634,O_3635,O_3636,O_3637,O_3638,O_3639,O_3640,O_3641,O_3642,O_3643,O_3644,O_3645,O_3646,O_3647,O_3648,O_3649,O_3650,O_3651,O_3652,O_3653,O_3654,O_3655,O_3656,O_3657,O_3658,O_3659,O_3660,O_3661,O_3662,O_3663,O_3664,O_3665,O_3666,O_3667,O_3668,O_3669,O_3670,O_3671,O_3672,O_3673,O_3674,O_3675,O_3676,O_3677,O_3678,O_3679,O_3680,O_3681,O_3682,O_3683,O_3684,O_3685,O_3686,O_3687,O_3688,O_3689,O_3690,O_3691,O_3692,O_3693,O_3694,O_3695,O_3696,O_3697,O_3698,O_3699,O_3700,O_3701,O_3702,O_3703,O_3704,O_3705,O_3706,O_3707,O_3708,O_3709,O_3710,O_3711,O_3712,O_3713,O_3714,O_3715,O_3716,O_3717,O_3718,O_3719,O_3720,O_3721,O_3722,O_3723,O_3724,O_3725,O_3726,O_3727,O_3728,O_3729,O_3730,O_3731,O_3732,O_3733,O_3734,O_3735,O_3736,O_3737,O_3738,O_3739,O_3740,O_3741,O_3742,O_3743,O_3744,O_3745,O_3746,O_3747,O_3748,O_3749,O_3750,O_3751,O_3752,O_3753,O_3754,O_3755,O_3756,O_3757,O_3758,O_3759,O_3760,O_3761,O_3762,O_3763,O_3764,O_3765,O_3766,O_3767,O_3768,O_3769,O_3770,O_3771,O_3772,O_3773,O_3774,O_3775,O_3776,O_3777,O_3778,O_3779,O_3780,O_3781,O_3782,O_3783,O_3784,O_3785,O_3786,O_3787,O_3788,O_3789,O_3790,O_3791,O_3792,O_3793,O_3794,O_3795,O_3796,O_3797,O_3798,O_3799,O_3800,O_3801,O_3802,O_3803,O_3804,O_3805,O_3806,O_3807,O_3808,O_3809,O_3810,O_3811,O_3812,O_3813,O_3814,O_3815,O_3816,O_3817,O_3818,O_3819,O_3820,O_3821,O_3822,O_3823,O_3824,O_3825,O_3826,O_3827,O_3828,O_3829,O_3830,O_3831,O_3832,O_3833,O_3834,O_3835,O_3836,O_3837,O_3838,O_3839,O_3840,O_3841,O_3842,O_3843,O_3844,O_3845,O_3846,O_3847,O_3848,O_3849,O_3850,O_3851,O_3852,O_3853,O_3854,O_3855,O_3856,O_3857,O_3858,O_3859,O_3860,O_3861,O_3862,O_3863,O_3864,O_3865,O_3866,O_3867,O_3868,O_3869,O_3870,O_3871,O_3872,O_3873,O_3874,O_3875,O_3876,O_3877,O_3878,O_3879,O_3880,O_3881,O_3882,O_3883,O_3884,O_3885,O_3886,O_3887,O_3888,O_3889,O_3890,O_3891,O_3892,O_3893,O_3894,O_3895,O_3896,O_3897,O_3898,O_3899,O_3900,O_3901,O_3902,O_3903,O_3904,O_3905,O_3906,O_3907,O_3908,O_3909,O_3910,O_3911,O_3912,O_3913,O_3914,O_3915,O_3916,O_3917,O_3918,O_3919,O_3920,O_3921,O_3922,O_3923,O_3924,O_3925,O_3926,O_3927,O_3928,O_3929,O_3930,O_3931,O_3932,O_3933,O_3934,O_3935,O_3936,O_3937,O_3938,O_3939,O_3940,O_3941,O_3942,O_3943,O_3944,O_3945,O_3946,O_3947,O_3948,O_3949,O_3950,O_3951,O_3952,O_3953,O_3954,O_3955,O_3956,O_3957,O_3958,O_3959,O_3960,O_3961,O_3962,O_3963,O_3964,O_3965,O_3966,O_3967,O_3968,O_3969,O_3970,O_3971,O_3972,O_3973,O_3974,O_3975,O_3976,O_3977,O_3978,O_3979,O_3980,O_3981,O_3982,O_3983,O_3984,O_3985,O_3986,O_3987,O_3988,O_3989,O_3990,O_3991,O_3992,O_3993,O_3994,O_3995,O_3996,O_3997,O_3998,O_3999,O_4000,O_4001,O_4002,O_4003,O_4004,O_4005,O_4006,O_4007,O_4008,O_4009,O_4010,O_4011,O_4012,O_4013,O_4014,O_4015,O_4016,O_4017,O_4018,O_4019,O_4020,O_4021,O_4022,O_4023,O_4024,O_4025,O_4026,O_4027,O_4028,O_4029,O_4030,O_4031,O_4032,O_4033,O_4034,O_4035,O_4036,O_4037,O_4038,O_4039,O_4040,O_4041,O_4042,O_4043,O_4044,O_4045,O_4046,O_4047,O_4048,O_4049,O_4050,O_4051,O_4052,O_4053,O_4054,O_4055,O_4056,O_4057,O_4058,O_4059,O_4060,O_4061,O_4062,O_4063,O_4064,O_4065,O_4066,O_4067,O_4068,O_4069,O_4070,O_4071,O_4072,O_4073,O_4074,O_4075,O_4076,O_4077,O_4078,O_4079,O_4080,O_4081,O_4082,O_4083,O_4084,O_4085,O_4086,O_4087,O_4088,O_4089,O_4090,O_4091,O_4092,O_4093,O_4094,O_4095,O_4096,O_4097,O_4098,O_4099,O_4100,O_4101,O_4102,O_4103,O_4104,O_4105,O_4106,O_4107,O_4108,O_4109,O_4110,O_4111,O_4112,O_4113,O_4114,O_4115,O_4116,O_4117,O_4118,O_4119,O_4120,O_4121,O_4122,O_4123,O_4124,O_4125,O_4126,O_4127,O_4128,O_4129,O_4130,O_4131,O_4132,O_4133,O_4134,O_4135,O_4136,O_4137,O_4138,O_4139,O_4140,O_4141,O_4142,O_4143,O_4144,O_4145,O_4146,O_4147,O_4148,O_4149,O_4150,O_4151,O_4152,O_4153,O_4154,O_4155,O_4156,O_4157,O_4158,O_4159,O_4160,O_4161,O_4162,O_4163,O_4164,O_4165,O_4166,O_4167,O_4168,O_4169,O_4170,O_4171,O_4172,O_4173,O_4174,O_4175,O_4176,O_4177,O_4178,O_4179,O_4180,O_4181,O_4182,O_4183,O_4184,O_4185,O_4186,O_4187,O_4188,O_4189,O_4190,O_4191,O_4192,O_4193,O_4194,O_4195,O_4196,O_4197,O_4198,O_4199,O_4200,O_4201,O_4202,O_4203,O_4204,O_4205,O_4206,O_4207,O_4208,O_4209,O_4210,O_4211,O_4212,O_4213,O_4214,O_4215,O_4216,O_4217,O_4218,O_4219,O_4220,O_4221,O_4222,O_4223,O_4224,O_4225,O_4226,O_4227,O_4228,O_4229,O_4230,O_4231,O_4232,O_4233,O_4234,O_4235,O_4236,O_4237,O_4238,O_4239,O_4240,O_4241,O_4242,O_4243,O_4244,O_4245,O_4246,O_4247,O_4248,O_4249,O_4250,O_4251,O_4252,O_4253,O_4254,O_4255,O_4256,O_4257,O_4258,O_4259,O_4260,O_4261,O_4262,O_4263,O_4264,O_4265,O_4266,O_4267,O_4268,O_4269,O_4270,O_4271,O_4272,O_4273,O_4274,O_4275,O_4276,O_4277,O_4278,O_4279,O_4280,O_4281,O_4282,O_4283,O_4284,O_4285,O_4286,O_4287,O_4288,O_4289,O_4290,O_4291,O_4292,O_4293,O_4294,O_4295,O_4296,O_4297,O_4298,O_4299,O_4300,O_4301,O_4302,O_4303,O_4304,O_4305,O_4306,O_4307,O_4308,O_4309,O_4310,O_4311,O_4312,O_4313,O_4314,O_4315,O_4316,O_4317,O_4318,O_4319,O_4320,O_4321,O_4322,O_4323,O_4324,O_4325,O_4326,O_4327,O_4328,O_4329,O_4330,O_4331,O_4332,O_4333,O_4334,O_4335,O_4336,O_4337,O_4338,O_4339,O_4340,O_4341,O_4342,O_4343,O_4344,O_4345,O_4346,O_4347,O_4348,O_4349,O_4350,O_4351,O_4352,O_4353,O_4354,O_4355,O_4356,O_4357,O_4358,O_4359,O_4360,O_4361,O_4362,O_4363,O_4364,O_4365,O_4366,O_4367,O_4368,O_4369,O_4370,O_4371,O_4372,O_4373,O_4374,O_4375,O_4376,O_4377,O_4378,O_4379,O_4380,O_4381,O_4382,O_4383,O_4384,O_4385,O_4386,O_4387,O_4388,O_4389,O_4390,O_4391,O_4392,O_4393,O_4394,O_4395,O_4396,O_4397,O_4398,O_4399,O_4400,O_4401,O_4402,O_4403,O_4404,O_4405,O_4406,O_4407,O_4408,O_4409,O_4410,O_4411,O_4412,O_4413,O_4414,O_4415,O_4416,O_4417,O_4418,O_4419,O_4420,O_4421,O_4422,O_4423,O_4424,O_4425,O_4426,O_4427,O_4428,O_4429,O_4430,O_4431,O_4432,O_4433,O_4434,O_4435,O_4436,O_4437,O_4438,O_4439,O_4440,O_4441,O_4442,O_4443,O_4444,O_4445,O_4446,O_4447,O_4448,O_4449,O_4450,O_4451,O_4452,O_4453,O_4454,O_4455,O_4456,O_4457,O_4458,O_4459,O_4460,O_4461,O_4462,O_4463,O_4464,O_4465,O_4466,O_4467,O_4468,O_4469,O_4470,O_4471,O_4472,O_4473,O_4474,O_4475,O_4476,O_4477,O_4478,O_4479,O_4480,O_4481,O_4482,O_4483,O_4484,O_4485,O_4486,O_4487,O_4488,O_4489,O_4490,O_4491,O_4492,O_4493,O_4494,O_4495,O_4496,O_4497,O_4498,O_4499,O_4500,O_4501,O_4502,O_4503,O_4504,O_4505,O_4506,O_4507,O_4508,O_4509,O_4510,O_4511,O_4512,O_4513,O_4514,O_4515,O_4516,O_4517,O_4518,O_4519,O_4520,O_4521,O_4522,O_4523,O_4524,O_4525,O_4526,O_4527,O_4528,O_4529,O_4530,O_4531,O_4532,O_4533,O_4534,O_4535,O_4536,O_4537,O_4538,O_4539,O_4540,O_4541,O_4542,O_4543,O_4544,O_4545,O_4546,O_4547,O_4548,O_4549,O_4550,O_4551,O_4552,O_4553,O_4554,O_4555,O_4556,O_4557,O_4558,O_4559,O_4560,O_4561,O_4562,O_4563,O_4564,O_4565,O_4566,O_4567,O_4568,O_4569,O_4570,O_4571,O_4572,O_4573,O_4574,O_4575,O_4576,O_4577,O_4578,O_4579,O_4580,O_4581,O_4582,O_4583,O_4584,O_4585,O_4586,O_4587,O_4588,O_4589,O_4590,O_4591,O_4592,O_4593,O_4594,O_4595,O_4596,O_4597,O_4598,O_4599,O_4600,O_4601,O_4602,O_4603,O_4604,O_4605,O_4606,O_4607,O_4608,O_4609,O_4610,O_4611,O_4612,O_4613,O_4614,O_4615,O_4616,O_4617,O_4618,O_4619,O_4620,O_4621,O_4622,O_4623,O_4624,O_4625,O_4626,O_4627,O_4628,O_4629,O_4630,O_4631,O_4632,O_4633,O_4634,O_4635,O_4636,O_4637,O_4638,O_4639,O_4640,O_4641,O_4642,O_4643,O_4644,O_4645,O_4646,O_4647,O_4648,O_4649,O_4650,O_4651,O_4652,O_4653,O_4654,O_4655,O_4656,O_4657,O_4658,O_4659,O_4660,O_4661,O_4662,O_4663,O_4664,O_4665,O_4666,O_4667,O_4668,O_4669,O_4670,O_4671,O_4672,O_4673,O_4674,O_4675,O_4676,O_4677,O_4678,O_4679,O_4680,O_4681,O_4682,O_4683,O_4684,O_4685,O_4686,O_4687,O_4688,O_4689,O_4690,O_4691,O_4692,O_4693,O_4694,O_4695,O_4696,O_4697,O_4698,O_4699,O_4700,O_4701,O_4702,O_4703,O_4704,O_4705,O_4706,O_4707,O_4708,O_4709,O_4710,O_4711,O_4712,O_4713,O_4714,O_4715,O_4716,O_4717,O_4718,O_4719,O_4720,O_4721,O_4722,O_4723,O_4724,O_4725,O_4726,O_4727,O_4728,O_4729,O_4730,O_4731,O_4732,O_4733,O_4734,O_4735,O_4736,O_4737,O_4738,O_4739,O_4740,O_4741,O_4742,O_4743,O_4744,O_4745,O_4746,O_4747,O_4748,O_4749,O_4750,O_4751,O_4752,O_4753,O_4754,O_4755,O_4756,O_4757,O_4758,O_4759,O_4760,O_4761,O_4762,O_4763,O_4764,O_4765,O_4766,O_4767,O_4768,O_4769,O_4770,O_4771,O_4772,O_4773,O_4774,O_4775,O_4776,O_4777,O_4778,O_4779,O_4780,O_4781,O_4782,O_4783,O_4784,O_4785,O_4786,O_4787,O_4788,O_4789,O_4790,O_4791,O_4792,O_4793,O_4794,O_4795,O_4796,O_4797,O_4798,O_4799,O_4800,O_4801,O_4802,O_4803,O_4804,O_4805,O_4806,O_4807,O_4808,O_4809,O_4810,O_4811,O_4812,O_4813,O_4814,O_4815,O_4816,O_4817,O_4818,O_4819,O_4820,O_4821,O_4822,O_4823,O_4824,O_4825,O_4826,O_4827,O_4828,O_4829,O_4830,O_4831,O_4832,O_4833,O_4834,O_4835,O_4836,O_4837,O_4838,O_4839,O_4840,O_4841,O_4842,O_4843,O_4844,O_4845,O_4846,O_4847,O_4848,O_4849,O_4850,O_4851,O_4852,O_4853,O_4854,O_4855,O_4856,O_4857,O_4858,O_4859,O_4860,O_4861,O_4862,O_4863,O_4864,O_4865,O_4866,O_4867,O_4868,O_4869,O_4870,O_4871,O_4872,O_4873,O_4874,O_4875,O_4876,O_4877,O_4878,O_4879,O_4880,O_4881,O_4882,O_4883,O_4884,O_4885,O_4886,O_4887,O_4888,O_4889,O_4890,O_4891,O_4892,O_4893,O_4894,O_4895,O_4896,O_4897,O_4898,O_4899,O_4900,O_4901,O_4902,O_4903,O_4904,O_4905,O_4906,O_4907,O_4908,O_4909,O_4910,O_4911,O_4912,O_4913,O_4914,O_4915,O_4916,O_4917,O_4918,O_4919,O_4920,O_4921,O_4922,O_4923,O_4924,O_4925,O_4926,O_4927,O_4928,O_4929,O_4930,O_4931,O_4932,O_4933,O_4934,O_4935,O_4936,O_4937,O_4938,O_4939,O_4940,O_4941,O_4942,O_4943,O_4944,O_4945,O_4946,O_4947,O_4948,O_4949,O_4950,O_4951,O_4952,O_4953,O_4954,O_4955,O_4956,O_4957,O_4958,O_4959,O_4960,O_4961,O_4962,O_4963,O_4964,O_4965,O_4966,O_4967,O_4968,O_4969,O_4970,O_4971,O_4972,O_4973,O_4974,O_4975,O_4976,O_4977,O_4978,O_4979,O_4980,O_4981,O_4982,O_4983,O_4984,O_4985,O_4986,O_4987,O_4988,O_4989,O_4990,O_4991,O_4992,O_4993,O_4994,O_4995,O_4996,O_4997,O_4998,O_4999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999,N_30000,N_30001,N_30002,N_30003,N_30004,N_30005,N_30006,N_30007,N_30008,N_30009,N_30010,N_30011,N_30012,N_30013,N_30014,N_30015,N_30016,N_30017,N_30018,N_30019,N_30020,N_30021,N_30022,N_30023,N_30024,N_30025,N_30026,N_30027,N_30028,N_30029,N_30030,N_30031,N_30032,N_30033,N_30034,N_30035,N_30036,N_30037,N_30038,N_30039,N_30040,N_30041,N_30042,N_30043,N_30044,N_30045,N_30046,N_30047,N_30048,N_30049,N_30050,N_30051,N_30052,N_30053,N_30054,N_30055,N_30056,N_30057,N_30058,N_30059,N_30060,N_30061,N_30062,N_30063,N_30064,N_30065,N_30066,N_30067,N_30068,N_30069,N_30070,N_30071,N_30072,N_30073,N_30074,N_30075,N_30076,N_30077,N_30078,N_30079,N_30080,N_30081,N_30082,N_30083,N_30084,N_30085,N_30086,N_30087,N_30088,N_30089,N_30090,N_30091,N_30092,N_30093,N_30094,N_30095,N_30096,N_30097,N_30098,N_30099,N_30100,N_30101,N_30102,N_30103,N_30104,N_30105,N_30106,N_30107,N_30108,N_30109,N_30110,N_30111,N_30112,N_30113,N_30114,N_30115,N_30116,N_30117,N_30118,N_30119,N_30120,N_30121,N_30122,N_30123,N_30124,N_30125,N_30126,N_30127,N_30128,N_30129,N_30130,N_30131,N_30132,N_30133,N_30134,N_30135,N_30136,N_30137,N_30138,N_30139,N_30140,N_30141,N_30142,N_30143,N_30144,N_30145,N_30146,N_30147,N_30148,N_30149,N_30150,N_30151,N_30152,N_30153,N_30154,N_30155,N_30156,N_30157,N_30158,N_30159,N_30160,N_30161,N_30162,N_30163,N_30164,N_30165,N_30166,N_30167,N_30168,N_30169,N_30170,N_30171,N_30172,N_30173,N_30174,N_30175,N_30176,N_30177,N_30178,N_30179,N_30180,N_30181,N_30182,N_30183,N_30184,N_30185,N_30186,N_30187,N_30188,N_30189,N_30190,N_30191,N_30192,N_30193,N_30194,N_30195,N_30196,N_30197,N_30198,N_30199,N_30200,N_30201,N_30202,N_30203,N_30204,N_30205,N_30206,N_30207,N_30208,N_30209,N_30210,N_30211,N_30212,N_30213,N_30214,N_30215,N_30216,N_30217,N_30218,N_30219,N_30220,N_30221,N_30222,N_30223,N_30224,N_30225,N_30226,N_30227,N_30228,N_30229,N_30230,N_30231,N_30232,N_30233,N_30234,N_30235,N_30236,N_30237,N_30238,N_30239,N_30240,N_30241,N_30242,N_30243,N_30244,N_30245,N_30246,N_30247,N_30248,N_30249,N_30250,N_30251,N_30252,N_30253,N_30254,N_30255,N_30256,N_30257,N_30258,N_30259,N_30260,N_30261,N_30262,N_30263,N_30264,N_30265,N_30266,N_30267,N_30268,N_30269,N_30270,N_30271,N_30272,N_30273,N_30274,N_30275,N_30276,N_30277,N_30278,N_30279,N_30280,N_30281,N_30282,N_30283,N_30284,N_30285,N_30286,N_30287,N_30288,N_30289,N_30290,N_30291,N_30292,N_30293,N_30294,N_30295,N_30296,N_30297,N_30298,N_30299,N_30300,N_30301,N_30302,N_30303,N_30304,N_30305,N_30306,N_30307,N_30308,N_30309,N_30310,N_30311,N_30312,N_30313,N_30314,N_30315,N_30316,N_30317,N_30318,N_30319,N_30320,N_30321,N_30322,N_30323,N_30324,N_30325,N_30326,N_30327,N_30328,N_30329,N_30330,N_30331,N_30332,N_30333,N_30334,N_30335,N_30336,N_30337,N_30338,N_30339,N_30340,N_30341,N_30342,N_30343,N_30344,N_30345,N_30346,N_30347,N_30348,N_30349,N_30350,N_30351,N_30352,N_30353,N_30354,N_30355,N_30356,N_30357,N_30358,N_30359,N_30360,N_30361,N_30362,N_30363,N_30364,N_30365,N_30366,N_30367,N_30368,N_30369,N_30370,N_30371,N_30372,N_30373,N_30374,N_30375,N_30376,N_30377,N_30378,N_30379,N_30380,N_30381,N_30382,N_30383,N_30384,N_30385,N_30386,N_30387,N_30388,N_30389,N_30390,N_30391,N_30392,N_30393,N_30394,N_30395,N_30396,N_30397,N_30398,N_30399,N_30400,N_30401,N_30402,N_30403,N_30404,N_30405,N_30406,N_30407,N_30408,N_30409,N_30410,N_30411,N_30412,N_30413,N_30414,N_30415,N_30416,N_30417,N_30418,N_30419,N_30420,N_30421,N_30422,N_30423,N_30424,N_30425,N_30426,N_30427,N_30428,N_30429,N_30430,N_30431,N_30432,N_30433,N_30434,N_30435,N_30436,N_30437,N_30438,N_30439,N_30440,N_30441,N_30442,N_30443,N_30444,N_30445,N_30446,N_30447,N_30448,N_30449,N_30450,N_30451,N_30452,N_30453,N_30454,N_30455,N_30456,N_30457,N_30458,N_30459,N_30460,N_30461,N_30462,N_30463,N_30464,N_30465,N_30466,N_30467,N_30468,N_30469,N_30470,N_30471,N_30472,N_30473,N_30474,N_30475,N_30476,N_30477,N_30478,N_30479,N_30480,N_30481,N_30482,N_30483,N_30484,N_30485,N_30486,N_30487,N_30488,N_30489,N_30490,N_30491,N_30492,N_30493,N_30494,N_30495,N_30496,N_30497,N_30498,N_30499,N_30500,N_30501,N_30502,N_30503,N_30504,N_30505,N_30506,N_30507,N_30508,N_30509,N_30510,N_30511,N_30512,N_30513,N_30514,N_30515,N_30516,N_30517,N_30518,N_30519,N_30520,N_30521,N_30522,N_30523,N_30524,N_30525,N_30526,N_30527,N_30528,N_30529,N_30530,N_30531,N_30532,N_30533,N_30534,N_30535,N_30536,N_30537,N_30538,N_30539,N_30540,N_30541,N_30542,N_30543,N_30544,N_30545,N_30546,N_30547,N_30548,N_30549,N_30550,N_30551,N_30552,N_30553,N_30554,N_30555,N_30556,N_30557,N_30558,N_30559,N_30560,N_30561,N_30562,N_30563,N_30564,N_30565,N_30566,N_30567,N_30568,N_30569,N_30570,N_30571,N_30572,N_30573,N_30574,N_30575,N_30576,N_30577,N_30578,N_30579,N_30580,N_30581,N_30582,N_30583,N_30584,N_30585,N_30586,N_30587,N_30588,N_30589,N_30590,N_30591,N_30592,N_30593,N_30594,N_30595,N_30596,N_30597,N_30598,N_30599,N_30600,N_30601,N_30602,N_30603,N_30604,N_30605,N_30606,N_30607,N_30608,N_30609,N_30610,N_30611,N_30612,N_30613,N_30614,N_30615,N_30616,N_30617,N_30618,N_30619,N_30620,N_30621,N_30622,N_30623,N_30624,N_30625,N_30626,N_30627,N_30628,N_30629,N_30630,N_30631,N_30632,N_30633,N_30634,N_30635,N_30636,N_30637,N_30638,N_30639,N_30640,N_30641,N_30642,N_30643,N_30644,N_30645,N_30646,N_30647,N_30648,N_30649,N_30650,N_30651,N_30652,N_30653,N_30654,N_30655,N_30656,N_30657,N_30658,N_30659,N_30660,N_30661,N_30662,N_30663,N_30664,N_30665,N_30666,N_30667,N_30668,N_30669,N_30670,N_30671,N_30672,N_30673,N_30674,N_30675,N_30676,N_30677,N_30678,N_30679,N_30680,N_30681,N_30682,N_30683,N_30684,N_30685,N_30686,N_30687,N_30688,N_30689,N_30690,N_30691,N_30692,N_30693,N_30694,N_30695,N_30696,N_30697,N_30698,N_30699,N_30700,N_30701,N_30702,N_30703,N_30704,N_30705,N_30706,N_30707,N_30708,N_30709,N_30710,N_30711,N_30712,N_30713,N_30714,N_30715,N_30716,N_30717,N_30718,N_30719,N_30720,N_30721,N_30722,N_30723,N_30724,N_30725,N_30726,N_30727,N_30728,N_30729,N_30730,N_30731,N_30732,N_30733,N_30734,N_30735,N_30736,N_30737,N_30738,N_30739,N_30740,N_30741,N_30742,N_30743,N_30744,N_30745,N_30746,N_30747,N_30748,N_30749,N_30750,N_30751,N_30752,N_30753,N_30754,N_30755,N_30756,N_30757,N_30758,N_30759,N_30760,N_30761,N_30762,N_30763,N_30764,N_30765,N_30766,N_30767,N_30768,N_30769,N_30770,N_30771,N_30772,N_30773,N_30774,N_30775,N_30776,N_30777,N_30778,N_30779,N_30780,N_30781,N_30782,N_30783,N_30784,N_30785,N_30786,N_30787,N_30788,N_30789,N_30790,N_30791,N_30792,N_30793,N_30794,N_30795,N_30796,N_30797,N_30798,N_30799,N_30800,N_30801,N_30802,N_30803,N_30804,N_30805,N_30806,N_30807,N_30808,N_30809,N_30810,N_30811,N_30812,N_30813,N_30814,N_30815,N_30816,N_30817,N_30818,N_30819,N_30820,N_30821,N_30822,N_30823,N_30824,N_30825,N_30826,N_30827,N_30828,N_30829,N_30830,N_30831,N_30832,N_30833,N_30834,N_30835,N_30836,N_30837,N_30838,N_30839,N_30840,N_30841,N_30842,N_30843,N_30844,N_30845,N_30846,N_30847,N_30848,N_30849,N_30850,N_30851,N_30852,N_30853,N_30854,N_30855,N_30856,N_30857,N_30858,N_30859,N_30860,N_30861,N_30862,N_30863,N_30864,N_30865,N_30866,N_30867,N_30868,N_30869,N_30870,N_30871,N_30872,N_30873,N_30874,N_30875,N_30876,N_30877,N_30878,N_30879,N_30880,N_30881,N_30882,N_30883,N_30884,N_30885,N_30886,N_30887,N_30888,N_30889,N_30890,N_30891,N_30892,N_30893,N_30894,N_30895,N_30896,N_30897,N_30898,N_30899,N_30900,N_30901,N_30902,N_30903,N_30904,N_30905,N_30906,N_30907,N_30908,N_30909,N_30910,N_30911,N_30912,N_30913,N_30914,N_30915,N_30916,N_30917,N_30918,N_30919,N_30920,N_30921,N_30922,N_30923,N_30924,N_30925,N_30926,N_30927,N_30928,N_30929,N_30930,N_30931,N_30932,N_30933,N_30934,N_30935,N_30936,N_30937,N_30938,N_30939,N_30940,N_30941,N_30942,N_30943,N_30944,N_30945,N_30946,N_30947,N_30948,N_30949,N_30950,N_30951,N_30952,N_30953,N_30954,N_30955,N_30956,N_30957,N_30958,N_30959,N_30960,N_30961,N_30962,N_30963,N_30964,N_30965,N_30966,N_30967,N_30968,N_30969,N_30970,N_30971,N_30972,N_30973,N_30974,N_30975,N_30976,N_30977,N_30978,N_30979,N_30980,N_30981,N_30982,N_30983,N_30984,N_30985,N_30986,N_30987,N_30988,N_30989,N_30990,N_30991,N_30992,N_30993,N_30994,N_30995,N_30996,N_30997,N_30998,N_30999,N_31000,N_31001,N_31002,N_31003,N_31004,N_31005,N_31006,N_31007,N_31008,N_31009,N_31010,N_31011,N_31012,N_31013,N_31014,N_31015,N_31016,N_31017,N_31018,N_31019,N_31020,N_31021,N_31022,N_31023,N_31024,N_31025,N_31026,N_31027,N_31028,N_31029,N_31030,N_31031,N_31032,N_31033,N_31034,N_31035,N_31036,N_31037,N_31038,N_31039,N_31040,N_31041,N_31042,N_31043,N_31044,N_31045,N_31046,N_31047,N_31048,N_31049,N_31050,N_31051,N_31052,N_31053,N_31054,N_31055,N_31056,N_31057,N_31058,N_31059,N_31060,N_31061,N_31062,N_31063,N_31064,N_31065,N_31066,N_31067,N_31068,N_31069,N_31070,N_31071,N_31072,N_31073,N_31074,N_31075,N_31076,N_31077,N_31078,N_31079,N_31080,N_31081,N_31082,N_31083,N_31084,N_31085,N_31086,N_31087,N_31088,N_31089,N_31090,N_31091,N_31092,N_31093,N_31094,N_31095,N_31096,N_31097,N_31098,N_31099,N_31100,N_31101,N_31102,N_31103,N_31104,N_31105,N_31106,N_31107,N_31108,N_31109,N_31110,N_31111,N_31112,N_31113,N_31114,N_31115,N_31116,N_31117,N_31118,N_31119,N_31120,N_31121,N_31122,N_31123,N_31124,N_31125,N_31126,N_31127,N_31128,N_31129,N_31130,N_31131,N_31132,N_31133,N_31134,N_31135,N_31136,N_31137,N_31138,N_31139,N_31140,N_31141,N_31142,N_31143,N_31144,N_31145,N_31146,N_31147,N_31148,N_31149,N_31150,N_31151,N_31152,N_31153,N_31154,N_31155,N_31156,N_31157,N_31158,N_31159,N_31160,N_31161,N_31162,N_31163,N_31164,N_31165,N_31166,N_31167,N_31168,N_31169,N_31170,N_31171,N_31172,N_31173,N_31174,N_31175,N_31176,N_31177,N_31178,N_31179,N_31180,N_31181,N_31182,N_31183,N_31184,N_31185,N_31186,N_31187,N_31188,N_31189,N_31190,N_31191,N_31192,N_31193,N_31194,N_31195,N_31196,N_31197,N_31198,N_31199,N_31200,N_31201,N_31202,N_31203,N_31204,N_31205,N_31206,N_31207,N_31208,N_31209,N_31210,N_31211,N_31212,N_31213,N_31214,N_31215,N_31216,N_31217,N_31218,N_31219,N_31220,N_31221,N_31222,N_31223,N_31224,N_31225,N_31226,N_31227,N_31228,N_31229,N_31230,N_31231,N_31232,N_31233,N_31234,N_31235,N_31236,N_31237,N_31238,N_31239,N_31240,N_31241,N_31242,N_31243,N_31244,N_31245,N_31246,N_31247,N_31248,N_31249,N_31250,N_31251,N_31252,N_31253,N_31254,N_31255,N_31256,N_31257,N_31258,N_31259,N_31260,N_31261,N_31262,N_31263,N_31264,N_31265,N_31266,N_31267,N_31268,N_31269,N_31270,N_31271,N_31272,N_31273,N_31274,N_31275,N_31276,N_31277,N_31278,N_31279,N_31280,N_31281,N_31282,N_31283,N_31284,N_31285,N_31286,N_31287,N_31288,N_31289,N_31290,N_31291,N_31292,N_31293,N_31294,N_31295,N_31296,N_31297,N_31298,N_31299,N_31300,N_31301,N_31302,N_31303,N_31304,N_31305,N_31306,N_31307,N_31308,N_31309,N_31310,N_31311,N_31312,N_31313,N_31314,N_31315,N_31316,N_31317,N_31318,N_31319,N_31320,N_31321,N_31322,N_31323,N_31324,N_31325,N_31326,N_31327,N_31328,N_31329,N_31330,N_31331,N_31332,N_31333,N_31334,N_31335,N_31336,N_31337,N_31338,N_31339,N_31340,N_31341,N_31342,N_31343,N_31344,N_31345,N_31346,N_31347,N_31348,N_31349,N_31350,N_31351,N_31352,N_31353,N_31354,N_31355,N_31356,N_31357,N_31358,N_31359,N_31360,N_31361,N_31362,N_31363,N_31364,N_31365,N_31366,N_31367,N_31368,N_31369,N_31370,N_31371,N_31372,N_31373,N_31374,N_31375,N_31376,N_31377,N_31378,N_31379,N_31380,N_31381,N_31382,N_31383,N_31384,N_31385,N_31386,N_31387,N_31388,N_31389,N_31390,N_31391,N_31392,N_31393,N_31394,N_31395,N_31396,N_31397,N_31398,N_31399,N_31400,N_31401,N_31402,N_31403,N_31404,N_31405,N_31406,N_31407,N_31408,N_31409,N_31410,N_31411,N_31412,N_31413,N_31414,N_31415,N_31416,N_31417,N_31418,N_31419,N_31420,N_31421,N_31422,N_31423,N_31424,N_31425,N_31426,N_31427,N_31428,N_31429,N_31430,N_31431,N_31432,N_31433,N_31434,N_31435,N_31436,N_31437,N_31438,N_31439,N_31440,N_31441,N_31442,N_31443,N_31444,N_31445,N_31446,N_31447,N_31448,N_31449,N_31450,N_31451,N_31452,N_31453,N_31454,N_31455,N_31456,N_31457,N_31458,N_31459,N_31460,N_31461,N_31462,N_31463,N_31464,N_31465,N_31466,N_31467,N_31468,N_31469,N_31470,N_31471,N_31472,N_31473,N_31474,N_31475,N_31476,N_31477,N_31478,N_31479,N_31480,N_31481,N_31482,N_31483,N_31484,N_31485,N_31486,N_31487,N_31488,N_31489,N_31490,N_31491,N_31492,N_31493,N_31494,N_31495,N_31496,N_31497,N_31498,N_31499,N_31500,N_31501,N_31502,N_31503,N_31504,N_31505,N_31506,N_31507,N_31508,N_31509,N_31510,N_31511,N_31512,N_31513,N_31514,N_31515,N_31516,N_31517,N_31518,N_31519,N_31520,N_31521,N_31522,N_31523,N_31524,N_31525,N_31526,N_31527,N_31528,N_31529,N_31530,N_31531,N_31532,N_31533,N_31534,N_31535,N_31536,N_31537,N_31538,N_31539,N_31540,N_31541,N_31542,N_31543,N_31544,N_31545,N_31546,N_31547,N_31548,N_31549,N_31550,N_31551,N_31552,N_31553,N_31554,N_31555,N_31556,N_31557,N_31558,N_31559,N_31560,N_31561,N_31562,N_31563,N_31564,N_31565,N_31566,N_31567,N_31568,N_31569,N_31570,N_31571,N_31572,N_31573,N_31574,N_31575,N_31576,N_31577,N_31578,N_31579,N_31580,N_31581,N_31582,N_31583,N_31584,N_31585,N_31586,N_31587,N_31588,N_31589,N_31590,N_31591,N_31592,N_31593,N_31594,N_31595,N_31596,N_31597,N_31598,N_31599,N_31600,N_31601,N_31602,N_31603,N_31604,N_31605,N_31606,N_31607,N_31608,N_31609,N_31610,N_31611,N_31612,N_31613,N_31614,N_31615,N_31616,N_31617,N_31618,N_31619,N_31620,N_31621,N_31622,N_31623,N_31624,N_31625,N_31626,N_31627,N_31628,N_31629,N_31630,N_31631,N_31632,N_31633,N_31634,N_31635,N_31636,N_31637,N_31638,N_31639,N_31640,N_31641,N_31642,N_31643,N_31644,N_31645,N_31646,N_31647,N_31648,N_31649,N_31650,N_31651,N_31652,N_31653,N_31654,N_31655,N_31656,N_31657,N_31658,N_31659,N_31660,N_31661,N_31662,N_31663,N_31664,N_31665,N_31666,N_31667,N_31668,N_31669,N_31670,N_31671,N_31672,N_31673,N_31674,N_31675,N_31676,N_31677,N_31678,N_31679,N_31680,N_31681,N_31682,N_31683,N_31684,N_31685,N_31686,N_31687,N_31688,N_31689,N_31690,N_31691,N_31692,N_31693,N_31694,N_31695,N_31696,N_31697,N_31698,N_31699,N_31700,N_31701,N_31702,N_31703,N_31704,N_31705,N_31706,N_31707,N_31708,N_31709,N_31710,N_31711,N_31712,N_31713,N_31714,N_31715,N_31716,N_31717,N_31718,N_31719,N_31720,N_31721,N_31722,N_31723,N_31724,N_31725,N_31726,N_31727,N_31728,N_31729,N_31730,N_31731,N_31732,N_31733,N_31734,N_31735,N_31736,N_31737,N_31738,N_31739,N_31740,N_31741,N_31742,N_31743,N_31744,N_31745,N_31746,N_31747,N_31748,N_31749,N_31750,N_31751,N_31752,N_31753,N_31754,N_31755,N_31756,N_31757,N_31758,N_31759,N_31760,N_31761,N_31762,N_31763,N_31764,N_31765,N_31766,N_31767,N_31768,N_31769,N_31770,N_31771,N_31772,N_31773,N_31774,N_31775,N_31776,N_31777,N_31778,N_31779,N_31780,N_31781,N_31782,N_31783,N_31784,N_31785,N_31786,N_31787,N_31788,N_31789,N_31790,N_31791,N_31792,N_31793,N_31794,N_31795,N_31796,N_31797,N_31798,N_31799,N_31800,N_31801,N_31802,N_31803,N_31804,N_31805,N_31806,N_31807,N_31808,N_31809,N_31810,N_31811,N_31812,N_31813,N_31814,N_31815,N_31816,N_31817,N_31818,N_31819,N_31820,N_31821,N_31822,N_31823,N_31824,N_31825,N_31826,N_31827,N_31828,N_31829,N_31830,N_31831,N_31832,N_31833,N_31834,N_31835,N_31836,N_31837,N_31838,N_31839,N_31840,N_31841,N_31842,N_31843,N_31844,N_31845,N_31846,N_31847,N_31848,N_31849,N_31850,N_31851,N_31852,N_31853,N_31854,N_31855,N_31856,N_31857,N_31858,N_31859,N_31860,N_31861,N_31862,N_31863,N_31864,N_31865,N_31866,N_31867,N_31868,N_31869,N_31870,N_31871,N_31872,N_31873,N_31874,N_31875,N_31876,N_31877,N_31878,N_31879,N_31880,N_31881,N_31882,N_31883,N_31884,N_31885,N_31886,N_31887,N_31888,N_31889,N_31890,N_31891,N_31892,N_31893,N_31894,N_31895,N_31896,N_31897,N_31898,N_31899,N_31900,N_31901,N_31902,N_31903,N_31904,N_31905,N_31906,N_31907,N_31908,N_31909,N_31910,N_31911,N_31912,N_31913,N_31914,N_31915,N_31916,N_31917,N_31918,N_31919,N_31920,N_31921,N_31922,N_31923,N_31924,N_31925,N_31926,N_31927,N_31928,N_31929,N_31930,N_31931,N_31932,N_31933,N_31934,N_31935,N_31936,N_31937,N_31938,N_31939,N_31940,N_31941,N_31942,N_31943,N_31944,N_31945,N_31946,N_31947,N_31948,N_31949,N_31950,N_31951,N_31952,N_31953,N_31954,N_31955,N_31956,N_31957,N_31958,N_31959,N_31960,N_31961,N_31962,N_31963,N_31964,N_31965,N_31966,N_31967,N_31968,N_31969,N_31970,N_31971,N_31972,N_31973,N_31974,N_31975,N_31976,N_31977,N_31978,N_31979,N_31980,N_31981,N_31982,N_31983,N_31984,N_31985,N_31986,N_31987,N_31988,N_31989,N_31990,N_31991,N_31992,N_31993,N_31994,N_31995,N_31996,N_31997,N_31998,N_31999,N_32000,N_32001,N_32002,N_32003,N_32004,N_32005,N_32006,N_32007,N_32008,N_32009,N_32010,N_32011,N_32012,N_32013,N_32014,N_32015,N_32016,N_32017,N_32018,N_32019,N_32020,N_32021,N_32022,N_32023,N_32024,N_32025,N_32026,N_32027,N_32028,N_32029,N_32030,N_32031,N_32032,N_32033,N_32034,N_32035,N_32036,N_32037,N_32038,N_32039,N_32040,N_32041,N_32042,N_32043,N_32044,N_32045,N_32046,N_32047,N_32048,N_32049,N_32050,N_32051,N_32052,N_32053,N_32054,N_32055,N_32056,N_32057,N_32058,N_32059,N_32060,N_32061,N_32062,N_32063,N_32064,N_32065,N_32066,N_32067,N_32068,N_32069,N_32070,N_32071,N_32072,N_32073,N_32074,N_32075,N_32076,N_32077,N_32078,N_32079,N_32080,N_32081,N_32082,N_32083,N_32084,N_32085,N_32086,N_32087,N_32088,N_32089,N_32090,N_32091,N_32092,N_32093,N_32094,N_32095,N_32096,N_32097,N_32098,N_32099,N_32100,N_32101,N_32102,N_32103,N_32104,N_32105,N_32106,N_32107,N_32108,N_32109,N_32110,N_32111,N_32112,N_32113,N_32114,N_32115,N_32116,N_32117,N_32118,N_32119,N_32120,N_32121,N_32122,N_32123,N_32124,N_32125,N_32126,N_32127,N_32128,N_32129,N_32130,N_32131,N_32132,N_32133,N_32134,N_32135,N_32136,N_32137,N_32138,N_32139,N_32140,N_32141,N_32142,N_32143,N_32144,N_32145,N_32146,N_32147,N_32148,N_32149,N_32150,N_32151,N_32152,N_32153,N_32154,N_32155,N_32156,N_32157,N_32158,N_32159,N_32160,N_32161,N_32162,N_32163,N_32164,N_32165,N_32166,N_32167,N_32168,N_32169,N_32170,N_32171,N_32172,N_32173,N_32174,N_32175,N_32176,N_32177,N_32178,N_32179,N_32180,N_32181,N_32182,N_32183,N_32184,N_32185,N_32186,N_32187,N_32188,N_32189,N_32190,N_32191,N_32192,N_32193,N_32194,N_32195,N_32196,N_32197,N_32198,N_32199,N_32200,N_32201,N_32202,N_32203,N_32204,N_32205,N_32206,N_32207,N_32208,N_32209,N_32210,N_32211,N_32212,N_32213,N_32214,N_32215,N_32216,N_32217,N_32218,N_32219,N_32220,N_32221,N_32222,N_32223,N_32224,N_32225,N_32226,N_32227,N_32228,N_32229,N_32230,N_32231,N_32232,N_32233,N_32234,N_32235,N_32236,N_32237,N_32238,N_32239,N_32240,N_32241,N_32242,N_32243,N_32244,N_32245,N_32246,N_32247,N_32248,N_32249,N_32250,N_32251,N_32252,N_32253,N_32254,N_32255,N_32256,N_32257,N_32258,N_32259,N_32260,N_32261,N_32262,N_32263,N_32264,N_32265,N_32266,N_32267,N_32268,N_32269,N_32270,N_32271,N_32272,N_32273,N_32274,N_32275,N_32276,N_32277,N_32278,N_32279,N_32280,N_32281,N_32282,N_32283,N_32284,N_32285,N_32286,N_32287,N_32288,N_32289,N_32290,N_32291,N_32292,N_32293,N_32294,N_32295,N_32296,N_32297,N_32298,N_32299,N_32300,N_32301,N_32302,N_32303,N_32304,N_32305,N_32306,N_32307,N_32308,N_32309,N_32310,N_32311,N_32312,N_32313,N_32314,N_32315,N_32316,N_32317,N_32318,N_32319,N_32320,N_32321,N_32322,N_32323,N_32324,N_32325,N_32326,N_32327,N_32328,N_32329,N_32330,N_32331,N_32332,N_32333,N_32334,N_32335,N_32336,N_32337,N_32338,N_32339,N_32340,N_32341,N_32342,N_32343,N_32344,N_32345,N_32346,N_32347,N_32348,N_32349,N_32350,N_32351,N_32352,N_32353,N_32354,N_32355,N_32356,N_32357,N_32358,N_32359,N_32360,N_32361,N_32362,N_32363,N_32364,N_32365,N_32366,N_32367,N_32368,N_32369,N_32370,N_32371,N_32372,N_32373,N_32374,N_32375,N_32376,N_32377,N_32378,N_32379,N_32380,N_32381,N_32382,N_32383,N_32384,N_32385,N_32386,N_32387,N_32388,N_32389,N_32390,N_32391,N_32392,N_32393,N_32394,N_32395,N_32396,N_32397,N_32398,N_32399,N_32400,N_32401,N_32402,N_32403,N_32404,N_32405,N_32406,N_32407,N_32408,N_32409,N_32410,N_32411,N_32412,N_32413,N_32414,N_32415,N_32416,N_32417,N_32418,N_32419,N_32420,N_32421,N_32422,N_32423,N_32424,N_32425,N_32426,N_32427,N_32428,N_32429,N_32430,N_32431,N_32432,N_32433,N_32434,N_32435,N_32436,N_32437,N_32438,N_32439,N_32440,N_32441,N_32442,N_32443,N_32444,N_32445,N_32446,N_32447,N_32448,N_32449,N_32450,N_32451,N_32452,N_32453,N_32454,N_32455,N_32456,N_32457,N_32458,N_32459,N_32460,N_32461,N_32462,N_32463,N_32464,N_32465,N_32466,N_32467,N_32468,N_32469,N_32470,N_32471,N_32472,N_32473,N_32474,N_32475,N_32476,N_32477,N_32478,N_32479,N_32480,N_32481,N_32482,N_32483,N_32484,N_32485,N_32486,N_32487,N_32488,N_32489,N_32490,N_32491,N_32492,N_32493,N_32494,N_32495,N_32496,N_32497,N_32498,N_32499,N_32500,N_32501,N_32502,N_32503,N_32504,N_32505,N_32506,N_32507,N_32508,N_32509,N_32510,N_32511,N_32512,N_32513,N_32514,N_32515,N_32516,N_32517,N_32518,N_32519,N_32520,N_32521,N_32522,N_32523,N_32524,N_32525,N_32526,N_32527,N_32528,N_32529,N_32530,N_32531,N_32532,N_32533,N_32534,N_32535,N_32536,N_32537,N_32538,N_32539,N_32540,N_32541,N_32542,N_32543,N_32544,N_32545,N_32546,N_32547,N_32548,N_32549,N_32550,N_32551,N_32552,N_32553,N_32554,N_32555,N_32556,N_32557,N_32558,N_32559,N_32560,N_32561,N_32562,N_32563,N_32564,N_32565,N_32566,N_32567,N_32568,N_32569,N_32570,N_32571,N_32572,N_32573,N_32574,N_32575,N_32576,N_32577,N_32578,N_32579,N_32580,N_32581,N_32582,N_32583,N_32584,N_32585,N_32586,N_32587,N_32588,N_32589,N_32590,N_32591,N_32592,N_32593,N_32594,N_32595,N_32596,N_32597,N_32598,N_32599,N_32600,N_32601,N_32602,N_32603,N_32604,N_32605,N_32606,N_32607,N_32608,N_32609,N_32610,N_32611,N_32612,N_32613,N_32614,N_32615,N_32616,N_32617,N_32618,N_32619,N_32620,N_32621,N_32622,N_32623,N_32624,N_32625,N_32626,N_32627,N_32628,N_32629,N_32630,N_32631,N_32632,N_32633,N_32634,N_32635,N_32636,N_32637,N_32638,N_32639,N_32640,N_32641,N_32642,N_32643,N_32644,N_32645,N_32646,N_32647,N_32648,N_32649,N_32650,N_32651,N_32652,N_32653,N_32654,N_32655,N_32656,N_32657,N_32658,N_32659,N_32660,N_32661,N_32662,N_32663,N_32664,N_32665,N_32666,N_32667,N_32668,N_32669,N_32670,N_32671,N_32672,N_32673,N_32674,N_32675,N_32676,N_32677,N_32678,N_32679,N_32680,N_32681,N_32682,N_32683,N_32684,N_32685,N_32686,N_32687,N_32688,N_32689,N_32690,N_32691,N_32692,N_32693,N_32694,N_32695,N_32696,N_32697,N_32698,N_32699,N_32700,N_32701,N_32702,N_32703,N_32704,N_32705,N_32706,N_32707,N_32708,N_32709,N_32710,N_32711,N_32712,N_32713,N_32714,N_32715,N_32716,N_32717,N_32718,N_32719,N_32720,N_32721,N_32722,N_32723,N_32724,N_32725,N_32726,N_32727,N_32728,N_32729,N_32730,N_32731,N_32732,N_32733,N_32734,N_32735,N_32736,N_32737,N_32738,N_32739,N_32740,N_32741,N_32742,N_32743,N_32744,N_32745,N_32746,N_32747,N_32748,N_32749,N_32750,N_32751,N_32752,N_32753,N_32754,N_32755,N_32756,N_32757,N_32758,N_32759,N_32760,N_32761,N_32762,N_32763,N_32764,N_32765,N_32766,N_32767,N_32768,N_32769,N_32770,N_32771,N_32772,N_32773,N_32774,N_32775,N_32776,N_32777,N_32778,N_32779,N_32780,N_32781,N_32782,N_32783,N_32784,N_32785,N_32786,N_32787,N_32788,N_32789,N_32790,N_32791,N_32792,N_32793,N_32794,N_32795,N_32796,N_32797,N_32798,N_32799,N_32800,N_32801,N_32802,N_32803,N_32804,N_32805,N_32806,N_32807,N_32808,N_32809,N_32810,N_32811,N_32812,N_32813,N_32814,N_32815,N_32816,N_32817,N_32818,N_32819,N_32820,N_32821,N_32822,N_32823,N_32824,N_32825,N_32826,N_32827,N_32828,N_32829,N_32830,N_32831,N_32832,N_32833,N_32834,N_32835,N_32836,N_32837,N_32838,N_32839,N_32840,N_32841,N_32842,N_32843,N_32844,N_32845,N_32846,N_32847,N_32848,N_32849,N_32850,N_32851,N_32852,N_32853,N_32854,N_32855,N_32856,N_32857,N_32858,N_32859,N_32860,N_32861,N_32862,N_32863,N_32864,N_32865,N_32866,N_32867,N_32868,N_32869,N_32870,N_32871,N_32872,N_32873,N_32874,N_32875,N_32876,N_32877,N_32878,N_32879,N_32880,N_32881,N_32882,N_32883,N_32884,N_32885,N_32886,N_32887,N_32888,N_32889,N_32890,N_32891,N_32892,N_32893,N_32894,N_32895,N_32896,N_32897,N_32898,N_32899,N_32900,N_32901,N_32902,N_32903,N_32904,N_32905,N_32906,N_32907,N_32908,N_32909,N_32910,N_32911,N_32912,N_32913,N_32914,N_32915,N_32916,N_32917,N_32918,N_32919,N_32920,N_32921,N_32922,N_32923,N_32924,N_32925,N_32926,N_32927,N_32928,N_32929,N_32930,N_32931,N_32932,N_32933,N_32934,N_32935,N_32936,N_32937,N_32938,N_32939,N_32940,N_32941,N_32942,N_32943,N_32944,N_32945,N_32946,N_32947,N_32948,N_32949,N_32950,N_32951,N_32952,N_32953,N_32954,N_32955,N_32956,N_32957,N_32958,N_32959,N_32960,N_32961,N_32962,N_32963,N_32964,N_32965,N_32966,N_32967,N_32968,N_32969,N_32970,N_32971,N_32972,N_32973,N_32974,N_32975,N_32976,N_32977,N_32978,N_32979,N_32980,N_32981,N_32982,N_32983,N_32984,N_32985,N_32986,N_32987,N_32988,N_32989,N_32990,N_32991,N_32992,N_32993,N_32994,N_32995,N_32996,N_32997,N_32998,N_32999,N_33000,N_33001,N_33002,N_33003,N_33004,N_33005,N_33006,N_33007,N_33008,N_33009,N_33010,N_33011,N_33012,N_33013,N_33014,N_33015,N_33016,N_33017,N_33018,N_33019,N_33020,N_33021,N_33022,N_33023,N_33024,N_33025,N_33026,N_33027,N_33028,N_33029,N_33030,N_33031,N_33032,N_33033,N_33034,N_33035,N_33036,N_33037,N_33038,N_33039,N_33040,N_33041,N_33042,N_33043,N_33044,N_33045,N_33046,N_33047,N_33048,N_33049,N_33050,N_33051,N_33052,N_33053,N_33054,N_33055,N_33056,N_33057,N_33058,N_33059,N_33060,N_33061,N_33062,N_33063,N_33064,N_33065,N_33066,N_33067,N_33068,N_33069,N_33070,N_33071,N_33072,N_33073,N_33074,N_33075,N_33076,N_33077,N_33078,N_33079,N_33080,N_33081,N_33082,N_33083,N_33084,N_33085,N_33086,N_33087,N_33088,N_33089,N_33090,N_33091,N_33092,N_33093,N_33094,N_33095,N_33096,N_33097,N_33098,N_33099,N_33100,N_33101,N_33102,N_33103,N_33104,N_33105,N_33106,N_33107,N_33108,N_33109,N_33110,N_33111,N_33112,N_33113,N_33114,N_33115,N_33116,N_33117,N_33118,N_33119,N_33120,N_33121,N_33122,N_33123,N_33124,N_33125,N_33126,N_33127,N_33128,N_33129,N_33130,N_33131,N_33132,N_33133,N_33134,N_33135,N_33136,N_33137,N_33138,N_33139,N_33140,N_33141,N_33142,N_33143,N_33144,N_33145,N_33146,N_33147,N_33148,N_33149,N_33150,N_33151,N_33152,N_33153,N_33154,N_33155,N_33156,N_33157,N_33158,N_33159,N_33160,N_33161,N_33162,N_33163,N_33164,N_33165,N_33166,N_33167,N_33168,N_33169,N_33170,N_33171,N_33172,N_33173,N_33174,N_33175,N_33176,N_33177,N_33178,N_33179,N_33180,N_33181,N_33182,N_33183,N_33184,N_33185,N_33186,N_33187,N_33188,N_33189,N_33190,N_33191,N_33192,N_33193,N_33194,N_33195,N_33196,N_33197,N_33198,N_33199,N_33200,N_33201,N_33202,N_33203,N_33204,N_33205,N_33206,N_33207,N_33208,N_33209,N_33210,N_33211,N_33212,N_33213,N_33214,N_33215,N_33216,N_33217,N_33218,N_33219,N_33220,N_33221,N_33222,N_33223,N_33224,N_33225,N_33226,N_33227,N_33228,N_33229,N_33230,N_33231,N_33232,N_33233,N_33234,N_33235,N_33236,N_33237,N_33238,N_33239,N_33240,N_33241,N_33242,N_33243,N_33244,N_33245,N_33246,N_33247,N_33248,N_33249,N_33250,N_33251,N_33252,N_33253,N_33254,N_33255,N_33256,N_33257,N_33258,N_33259,N_33260,N_33261,N_33262,N_33263,N_33264,N_33265,N_33266,N_33267,N_33268,N_33269,N_33270,N_33271,N_33272,N_33273,N_33274,N_33275,N_33276,N_33277,N_33278,N_33279,N_33280,N_33281,N_33282,N_33283,N_33284,N_33285,N_33286,N_33287,N_33288,N_33289,N_33290,N_33291,N_33292,N_33293,N_33294,N_33295,N_33296,N_33297,N_33298,N_33299,N_33300,N_33301,N_33302,N_33303,N_33304,N_33305,N_33306,N_33307,N_33308,N_33309,N_33310,N_33311,N_33312,N_33313,N_33314,N_33315,N_33316,N_33317,N_33318,N_33319,N_33320,N_33321,N_33322,N_33323,N_33324,N_33325,N_33326,N_33327,N_33328,N_33329,N_33330,N_33331,N_33332,N_33333,N_33334,N_33335,N_33336,N_33337,N_33338,N_33339,N_33340,N_33341,N_33342,N_33343,N_33344,N_33345,N_33346,N_33347,N_33348,N_33349,N_33350,N_33351,N_33352,N_33353,N_33354,N_33355,N_33356,N_33357,N_33358,N_33359,N_33360,N_33361,N_33362,N_33363,N_33364,N_33365,N_33366,N_33367,N_33368,N_33369,N_33370,N_33371,N_33372,N_33373,N_33374,N_33375,N_33376,N_33377,N_33378,N_33379,N_33380,N_33381,N_33382,N_33383,N_33384,N_33385,N_33386,N_33387,N_33388,N_33389,N_33390,N_33391,N_33392,N_33393,N_33394,N_33395,N_33396,N_33397,N_33398,N_33399,N_33400,N_33401,N_33402,N_33403,N_33404,N_33405,N_33406,N_33407,N_33408,N_33409,N_33410,N_33411,N_33412,N_33413,N_33414,N_33415,N_33416,N_33417,N_33418,N_33419,N_33420,N_33421,N_33422,N_33423,N_33424,N_33425,N_33426,N_33427,N_33428,N_33429,N_33430,N_33431,N_33432,N_33433,N_33434,N_33435,N_33436,N_33437,N_33438,N_33439,N_33440,N_33441,N_33442,N_33443,N_33444,N_33445,N_33446,N_33447,N_33448,N_33449,N_33450,N_33451,N_33452,N_33453,N_33454,N_33455,N_33456,N_33457,N_33458,N_33459,N_33460,N_33461,N_33462,N_33463,N_33464,N_33465,N_33466,N_33467,N_33468,N_33469,N_33470,N_33471,N_33472,N_33473,N_33474,N_33475,N_33476,N_33477,N_33478,N_33479,N_33480,N_33481,N_33482,N_33483,N_33484,N_33485,N_33486,N_33487,N_33488,N_33489,N_33490,N_33491,N_33492,N_33493,N_33494,N_33495,N_33496,N_33497,N_33498,N_33499,N_33500,N_33501,N_33502,N_33503,N_33504,N_33505,N_33506,N_33507,N_33508,N_33509,N_33510,N_33511,N_33512,N_33513,N_33514,N_33515,N_33516,N_33517,N_33518,N_33519,N_33520,N_33521,N_33522,N_33523,N_33524,N_33525,N_33526,N_33527,N_33528,N_33529,N_33530,N_33531,N_33532,N_33533,N_33534,N_33535,N_33536,N_33537,N_33538,N_33539,N_33540,N_33541,N_33542,N_33543,N_33544,N_33545,N_33546,N_33547,N_33548,N_33549,N_33550,N_33551,N_33552,N_33553,N_33554,N_33555,N_33556,N_33557,N_33558,N_33559,N_33560,N_33561,N_33562,N_33563,N_33564,N_33565,N_33566,N_33567,N_33568,N_33569,N_33570,N_33571,N_33572,N_33573,N_33574,N_33575,N_33576,N_33577,N_33578,N_33579,N_33580,N_33581,N_33582,N_33583,N_33584,N_33585,N_33586,N_33587,N_33588,N_33589,N_33590,N_33591,N_33592,N_33593,N_33594,N_33595,N_33596,N_33597,N_33598,N_33599,N_33600,N_33601,N_33602,N_33603,N_33604,N_33605,N_33606,N_33607,N_33608,N_33609,N_33610,N_33611,N_33612,N_33613,N_33614,N_33615,N_33616,N_33617,N_33618,N_33619,N_33620,N_33621,N_33622,N_33623,N_33624,N_33625,N_33626,N_33627,N_33628,N_33629,N_33630,N_33631,N_33632,N_33633,N_33634,N_33635,N_33636,N_33637,N_33638,N_33639,N_33640,N_33641,N_33642,N_33643,N_33644,N_33645,N_33646,N_33647,N_33648,N_33649,N_33650,N_33651,N_33652,N_33653,N_33654,N_33655,N_33656,N_33657,N_33658,N_33659,N_33660,N_33661,N_33662,N_33663,N_33664,N_33665,N_33666,N_33667,N_33668,N_33669,N_33670,N_33671,N_33672,N_33673,N_33674,N_33675,N_33676,N_33677,N_33678,N_33679,N_33680,N_33681,N_33682,N_33683,N_33684,N_33685,N_33686,N_33687,N_33688,N_33689,N_33690,N_33691,N_33692,N_33693,N_33694,N_33695,N_33696,N_33697,N_33698,N_33699,N_33700,N_33701,N_33702,N_33703,N_33704,N_33705,N_33706,N_33707,N_33708,N_33709,N_33710,N_33711,N_33712,N_33713,N_33714,N_33715,N_33716,N_33717,N_33718,N_33719,N_33720,N_33721,N_33722,N_33723,N_33724,N_33725,N_33726,N_33727,N_33728,N_33729,N_33730,N_33731,N_33732,N_33733,N_33734,N_33735,N_33736,N_33737,N_33738,N_33739,N_33740,N_33741,N_33742,N_33743,N_33744,N_33745,N_33746,N_33747,N_33748,N_33749,N_33750,N_33751,N_33752,N_33753,N_33754,N_33755,N_33756,N_33757,N_33758,N_33759,N_33760,N_33761,N_33762,N_33763,N_33764,N_33765,N_33766,N_33767,N_33768,N_33769,N_33770,N_33771,N_33772,N_33773,N_33774,N_33775,N_33776,N_33777,N_33778,N_33779,N_33780,N_33781,N_33782,N_33783,N_33784,N_33785,N_33786,N_33787,N_33788,N_33789,N_33790,N_33791,N_33792,N_33793,N_33794,N_33795,N_33796,N_33797,N_33798,N_33799,N_33800,N_33801,N_33802,N_33803,N_33804,N_33805,N_33806,N_33807,N_33808,N_33809,N_33810,N_33811,N_33812,N_33813,N_33814,N_33815,N_33816,N_33817,N_33818,N_33819,N_33820,N_33821,N_33822,N_33823,N_33824,N_33825,N_33826,N_33827,N_33828,N_33829,N_33830,N_33831,N_33832,N_33833,N_33834,N_33835,N_33836,N_33837,N_33838,N_33839,N_33840,N_33841,N_33842,N_33843,N_33844,N_33845,N_33846,N_33847,N_33848,N_33849,N_33850,N_33851,N_33852,N_33853,N_33854,N_33855,N_33856,N_33857,N_33858,N_33859,N_33860,N_33861,N_33862,N_33863,N_33864,N_33865,N_33866,N_33867,N_33868,N_33869,N_33870,N_33871,N_33872,N_33873,N_33874,N_33875,N_33876,N_33877,N_33878,N_33879,N_33880,N_33881,N_33882,N_33883,N_33884,N_33885,N_33886,N_33887,N_33888,N_33889,N_33890,N_33891,N_33892,N_33893,N_33894,N_33895,N_33896,N_33897,N_33898,N_33899,N_33900,N_33901,N_33902,N_33903,N_33904,N_33905,N_33906,N_33907,N_33908,N_33909,N_33910,N_33911,N_33912,N_33913,N_33914,N_33915,N_33916,N_33917,N_33918,N_33919,N_33920,N_33921,N_33922,N_33923,N_33924,N_33925,N_33926,N_33927,N_33928,N_33929,N_33930,N_33931,N_33932,N_33933,N_33934,N_33935,N_33936,N_33937,N_33938,N_33939,N_33940,N_33941,N_33942,N_33943,N_33944,N_33945,N_33946,N_33947,N_33948,N_33949,N_33950,N_33951,N_33952,N_33953,N_33954,N_33955,N_33956,N_33957,N_33958,N_33959,N_33960,N_33961,N_33962,N_33963,N_33964,N_33965,N_33966,N_33967,N_33968,N_33969,N_33970,N_33971,N_33972,N_33973,N_33974,N_33975,N_33976,N_33977,N_33978,N_33979,N_33980,N_33981,N_33982,N_33983,N_33984,N_33985,N_33986,N_33987,N_33988,N_33989,N_33990,N_33991,N_33992,N_33993,N_33994,N_33995,N_33996,N_33997,N_33998,N_33999,N_34000,N_34001,N_34002,N_34003,N_34004,N_34005,N_34006,N_34007,N_34008,N_34009,N_34010,N_34011,N_34012,N_34013,N_34014,N_34015,N_34016,N_34017,N_34018,N_34019,N_34020,N_34021,N_34022,N_34023,N_34024,N_34025,N_34026,N_34027,N_34028,N_34029,N_34030,N_34031,N_34032,N_34033,N_34034,N_34035,N_34036,N_34037,N_34038,N_34039,N_34040,N_34041,N_34042,N_34043,N_34044,N_34045,N_34046,N_34047,N_34048,N_34049,N_34050,N_34051,N_34052,N_34053,N_34054,N_34055,N_34056,N_34057,N_34058,N_34059,N_34060,N_34061,N_34062,N_34063,N_34064,N_34065,N_34066,N_34067,N_34068,N_34069,N_34070,N_34071,N_34072,N_34073,N_34074,N_34075,N_34076,N_34077,N_34078,N_34079,N_34080,N_34081,N_34082,N_34083,N_34084,N_34085,N_34086,N_34087,N_34088,N_34089,N_34090,N_34091,N_34092,N_34093,N_34094,N_34095,N_34096,N_34097,N_34098,N_34099,N_34100,N_34101,N_34102,N_34103,N_34104,N_34105,N_34106,N_34107,N_34108,N_34109,N_34110,N_34111,N_34112,N_34113,N_34114,N_34115,N_34116,N_34117,N_34118,N_34119,N_34120,N_34121,N_34122,N_34123,N_34124,N_34125,N_34126,N_34127,N_34128,N_34129,N_34130,N_34131,N_34132,N_34133,N_34134,N_34135,N_34136,N_34137,N_34138,N_34139,N_34140,N_34141,N_34142,N_34143,N_34144,N_34145,N_34146,N_34147,N_34148,N_34149,N_34150,N_34151,N_34152,N_34153,N_34154,N_34155,N_34156,N_34157,N_34158,N_34159,N_34160,N_34161,N_34162,N_34163,N_34164,N_34165,N_34166,N_34167,N_34168,N_34169,N_34170,N_34171,N_34172,N_34173,N_34174,N_34175,N_34176,N_34177,N_34178,N_34179,N_34180,N_34181,N_34182,N_34183,N_34184,N_34185,N_34186,N_34187,N_34188,N_34189,N_34190,N_34191,N_34192,N_34193,N_34194,N_34195,N_34196,N_34197,N_34198,N_34199,N_34200,N_34201,N_34202,N_34203,N_34204,N_34205,N_34206,N_34207,N_34208,N_34209,N_34210,N_34211,N_34212,N_34213,N_34214,N_34215,N_34216,N_34217,N_34218,N_34219,N_34220,N_34221,N_34222,N_34223,N_34224,N_34225,N_34226,N_34227,N_34228,N_34229,N_34230,N_34231,N_34232,N_34233,N_34234,N_34235,N_34236,N_34237,N_34238,N_34239,N_34240,N_34241,N_34242,N_34243,N_34244,N_34245,N_34246,N_34247,N_34248,N_34249,N_34250,N_34251,N_34252,N_34253,N_34254,N_34255,N_34256,N_34257,N_34258,N_34259,N_34260,N_34261,N_34262,N_34263,N_34264,N_34265,N_34266,N_34267,N_34268,N_34269,N_34270,N_34271,N_34272,N_34273,N_34274,N_34275,N_34276,N_34277,N_34278,N_34279,N_34280,N_34281,N_34282,N_34283,N_34284,N_34285,N_34286,N_34287,N_34288,N_34289,N_34290,N_34291,N_34292,N_34293,N_34294,N_34295,N_34296,N_34297,N_34298,N_34299,N_34300,N_34301,N_34302,N_34303,N_34304,N_34305,N_34306,N_34307,N_34308,N_34309,N_34310,N_34311,N_34312,N_34313,N_34314,N_34315,N_34316,N_34317,N_34318,N_34319,N_34320,N_34321,N_34322,N_34323,N_34324,N_34325,N_34326,N_34327,N_34328,N_34329,N_34330,N_34331,N_34332,N_34333,N_34334,N_34335,N_34336,N_34337,N_34338,N_34339,N_34340,N_34341,N_34342,N_34343,N_34344,N_34345,N_34346,N_34347,N_34348,N_34349,N_34350,N_34351,N_34352,N_34353,N_34354,N_34355,N_34356,N_34357,N_34358,N_34359,N_34360,N_34361,N_34362,N_34363,N_34364,N_34365,N_34366,N_34367,N_34368,N_34369,N_34370,N_34371,N_34372,N_34373,N_34374,N_34375,N_34376,N_34377,N_34378,N_34379,N_34380,N_34381,N_34382,N_34383,N_34384,N_34385,N_34386,N_34387,N_34388,N_34389,N_34390,N_34391,N_34392,N_34393,N_34394,N_34395,N_34396,N_34397,N_34398,N_34399,N_34400,N_34401,N_34402,N_34403,N_34404,N_34405,N_34406,N_34407,N_34408,N_34409,N_34410,N_34411,N_34412,N_34413,N_34414,N_34415,N_34416,N_34417,N_34418,N_34419,N_34420,N_34421,N_34422,N_34423,N_34424,N_34425,N_34426,N_34427,N_34428,N_34429,N_34430,N_34431,N_34432,N_34433,N_34434,N_34435,N_34436,N_34437,N_34438,N_34439,N_34440,N_34441,N_34442,N_34443,N_34444,N_34445,N_34446,N_34447,N_34448,N_34449,N_34450,N_34451,N_34452,N_34453,N_34454,N_34455,N_34456,N_34457,N_34458,N_34459,N_34460,N_34461,N_34462,N_34463,N_34464,N_34465,N_34466,N_34467,N_34468,N_34469,N_34470,N_34471,N_34472,N_34473,N_34474,N_34475,N_34476,N_34477,N_34478,N_34479,N_34480,N_34481,N_34482,N_34483,N_34484,N_34485,N_34486,N_34487,N_34488,N_34489,N_34490,N_34491,N_34492,N_34493,N_34494,N_34495,N_34496,N_34497,N_34498,N_34499,N_34500,N_34501,N_34502,N_34503,N_34504,N_34505,N_34506,N_34507,N_34508,N_34509,N_34510,N_34511,N_34512,N_34513,N_34514,N_34515,N_34516,N_34517,N_34518,N_34519,N_34520,N_34521,N_34522,N_34523,N_34524,N_34525,N_34526,N_34527,N_34528,N_34529,N_34530,N_34531,N_34532,N_34533,N_34534,N_34535,N_34536,N_34537,N_34538,N_34539,N_34540,N_34541,N_34542,N_34543,N_34544,N_34545,N_34546,N_34547,N_34548,N_34549,N_34550,N_34551,N_34552,N_34553,N_34554,N_34555,N_34556,N_34557,N_34558,N_34559,N_34560,N_34561,N_34562,N_34563,N_34564,N_34565,N_34566,N_34567,N_34568,N_34569,N_34570,N_34571,N_34572,N_34573,N_34574,N_34575,N_34576,N_34577,N_34578,N_34579,N_34580,N_34581,N_34582,N_34583,N_34584,N_34585,N_34586,N_34587,N_34588,N_34589,N_34590,N_34591,N_34592,N_34593,N_34594,N_34595,N_34596,N_34597,N_34598,N_34599,N_34600,N_34601,N_34602,N_34603,N_34604,N_34605,N_34606,N_34607,N_34608,N_34609,N_34610,N_34611,N_34612,N_34613,N_34614,N_34615,N_34616,N_34617,N_34618,N_34619,N_34620,N_34621,N_34622,N_34623,N_34624,N_34625,N_34626,N_34627,N_34628,N_34629,N_34630,N_34631,N_34632,N_34633,N_34634,N_34635,N_34636,N_34637,N_34638,N_34639,N_34640,N_34641,N_34642,N_34643,N_34644,N_34645,N_34646,N_34647,N_34648,N_34649,N_34650,N_34651,N_34652,N_34653,N_34654,N_34655,N_34656,N_34657,N_34658,N_34659,N_34660,N_34661,N_34662,N_34663,N_34664,N_34665,N_34666,N_34667,N_34668,N_34669,N_34670,N_34671,N_34672,N_34673,N_34674,N_34675,N_34676,N_34677,N_34678,N_34679,N_34680,N_34681,N_34682,N_34683,N_34684,N_34685,N_34686,N_34687,N_34688,N_34689,N_34690,N_34691,N_34692,N_34693,N_34694,N_34695,N_34696,N_34697,N_34698,N_34699,N_34700,N_34701,N_34702,N_34703,N_34704,N_34705,N_34706,N_34707,N_34708,N_34709,N_34710,N_34711,N_34712,N_34713,N_34714,N_34715,N_34716,N_34717,N_34718,N_34719,N_34720,N_34721,N_34722,N_34723,N_34724,N_34725,N_34726,N_34727,N_34728,N_34729,N_34730,N_34731,N_34732,N_34733,N_34734,N_34735,N_34736,N_34737,N_34738,N_34739,N_34740,N_34741,N_34742,N_34743,N_34744,N_34745,N_34746,N_34747,N_34748,N_34749,N_34750,N_34751,N_34752,N_34753,N_34754,N_34755,N_34756,N_34757,N_34758,N_34759,N_34760,N_34761,N_34762,N_34763,N_34764,N_34765,N_34766,N_34767,N_34768,N_34769,N_34770,N_34771,N_34772,N_34773,N_34774,N_34775,N_34776,N_34777,N_34778,N_34779,N_34780,N_34781,N_34782,N_34783,N_34784,N_34785,N_34786,N_34787,N_34788,N_34789,N_34790,N_34791,N_34792,N_34793,N_34794,N_34795,N_34796,N_34797,N_34798,N_34799,N_34800,N_34801,N_34802,N_34803,N_34804,N_34805,N_34806,N_34807,N_34808,N_34809,N_34810,N_34811,N_34812,N_34813,N_34814,N_34815,N_34816,N_34817,N_34818,N_34819,N_34820,N_34821,N_34822,N_34823,N_34824,N_34825,N_34826,N_34827,N_34828,N_34829,N_34830,N_34831,N_34832,N_34833,N_34834,N_34835,N_34836,N_34837,N_34838,N_34839,N_34840,N_34841,N_34842,N_34843,N_34844,N_34845,N_34846,N_34847,N_34848,N_34849,N_34850,N_34851,N_34852,N_34853,N_34854,N_34855,N_34856,N_34857,N_34858,N_34859,N_34860,N_34861,N_34862,N_34863,N_34864,N_34865,N_34866,N_34867,N_34868,N_34869,N_34870,N_34871,N_34872,N_34873,N_34874,N_34875,N_34876,N_34877,N_34878,N_34879,N_34880,N_34881,N_34882,N_34883,N_34884,N_34885,N_34886,N_34887,N_34888,N_34889,N_34890,N_34891,N_34892,N_34893,N_34894,N_34895,N_34896,N_34897,N_34898,N_34899,N_34900,N_34901,N_34902,N_34903,N_34904,N_34905,N_34906,N_34907,N_34908,N_34909,N_34910,N_34911,N_34912,N_34913,N_34914,N_34915,N_34916,N_34917,N_34918,N_34919,N_34920,N_34921,N_34922,N_34923,N_34924,N_34925,N_34926,N_34927,N_34928,N_34929,N_34930,N_34931,N_34932,N_34933,N_34934,N_34935,N_34936,N_34937,N_34938,N_34939,N_34940,N_34941,N_34942,N_34943,N_34944,N_34945,N_34946,N_34947,N_34948,N_34949,N_34950,N_34951,N_34952,N_34953,N_34954,N_34955,N_34956,N_34957,N_34958,N_34959,N_34960,N_34961,N_34962,N_34963,N_34964,N_34965,N_34966,N_34967,N_34968,N_34969,N_34970,N_34971,N_34972,N_34973,N_34974,N_34975,N_34976,N_34977,N_34978,N_34979,N_34980,N_34981,N_34982,N_34983,N_34984,N_34985,N_34986,N_34987,N_34988,N_34989,N_34990,N_34991,N_34992,N_34993,N_34994,N_34995,N_34996,N_34997,N_34998,N_34999,N_35000,N_35001,N_35002,N_35003,N_35004,N_35005,N_35006,N_35007,N_35008,N_35009,N_35010,N_35011,N_35012,N_35013,N_35014,N_35015,N_35016,N_35017,N_35018,N_35019,N_35020,N_35021,N_35022,N_35023,N_35024,N_35025,N_35026,N_35027,N_35028,N_35029,N_35030,N_35031,N_35032,N_35033,N_35034,N_35035,N_35036,N_35037,N_35038,N_35039,N_35040,N_35041,N_35042,N_35043,N_35044,N_35045,N_35046,N_35047,N_35048,N_35049,N_35050,N_35051,N_35052,N_35053,N_35054,N_35055,N_35056,N_35057,N_35058,N_35059,N_35060,N_35061,N_35062,N_35063,N_35064,N_35065,N_35066,N_35067,N_35068,N_35069,N_35070,N_35071,N_35072,N_35073,N_35074,N_35075,N_35076,N_35077,N_35078,N_35079,N_35080,N_35081,N_35082,N_35083,N_35084,N_35085,N_35086,N_35087,N_35088,N_35089,N_35090,N_35091,N_35092,N_35093,N_35094,N_35095,N_35096,N_35097,N_35098,N_35099,N_35100,N_35101,N_35102,N_35103,N_35104,N_35105,N_35106,N_35107,N_35108,N_35109,N_35110,N_35111,N_35112,N_35113,N_35114,N_35115,N_35116,N_35117,N_35118,N_35119,N_35120,N_35121,N_35122,N_35123,N_35124,N_35125,N_35126,N_35127,N_35128,N_35129,N_35130,N_35131,N_35132,N_35133,N_35134,N_35135,N_35136,N_35137,N_35138,N_35139,N_35140,N_35141,N_35142,N_35143,N_35144,N_35145,N_35146,N_35147,N_35148,N_35149,N_35150,N_35151,N_35152,N_35153,N_35154,N_35155,N_35156,N_35157,N_35158,N_35159,N_35160,N_35161,N_35162,N_35163,N_35164,N_35165,N_35166,N_35167,N_35168,N_35169,N_35170,N_35171,N_35172,N_35173,N_35174,N_35175,N_35176,N_35177,N_35178,N_35179,N_35180,N_35181,N_35182,N_35183,N_35184,N_35185,N_35186,N_35187,N_35188,N_35189,N_35190,N_35191,N_35192,N_35193,N_35194,N_35195,N_35196,N_35197,N_35198,N_35199,N_35200,N_35201,N_35202,N_35203,N_35204,N_35205,N_35206,N_35207,N_35208,N_35209,N_35210,N_35211,N_35212,N_35213,N_35214,N_35215,N_35216,N_35217,N_35218,N_35219,N_35220,N_35221,N_35222,N_35223,N_35224,N_35225,N_35226,N_35227,N_35228,N_35229,N_35230,N_35231,N_35232,N_35233,N_35234,N_35235,N_35236,N_35237,N_35238,N_35239,N_35240,N_35241,N_35242,N_35243,N_35244,N_35245,N_35246,N_35247,N_35248,N_35249,N_35250,N_35251,N_35252,N_35253,N_35254,N_35255,N_35256,N_35257,N_35258,N_35259,N_35260,N_35261,N_35262,N_35263,N_35264,N_35265,N_35266,N_35267,N_35268,N_35269,N_35270,N_35271,N_35272,N_35273,N_35274,N_35275,N_35276,N_35277,N_35278,N_35279,N_35280,N_35281,N_35282,N_35283,N_35284,N_35285,N_35286,N_35287,N_35288,N_35289,N_35290,N_35291,N_35292,N_35293,N_35294,N_35295,N_35296,N_35297,N_35298,N_35299,N_35300,N_35301,N_35302,N_35303,N_35304,N_35305,N_35306,N_35307,N_35308,N_35309,N_35310,N_35311,N_35312,N_35313,N_35314,N_35315,N_35316,N_35317,N_35318,N_35319,N_35320,N_35321,N_35322,N_35323,N_35324,N_35325,N_35326,N_35327,N_35328,N_35329,N_35330,N_35331,N_35332,N_35333,N_35334,N_35335,N_35336,N_35337,N_35338,N_35339,N_35340,N_35341,N_35342,N_35343,N_35344,N_35345,N_35346,N_35347,N_35348,N_35349,N_35350,N_35351,N_35352,N_35353,N_35354,N_35355,N_35356,N_35357,N_35358,N_35359,N_35360,N_35361,N_35362,N_35363,N_35364,N_35365,N_35366,N_35367,N_35368,N_35369,N_35370,N_35371,N_35372,N_35373,N_35374,N_35375,N_35376,N_35377,N_35378,N_35379,N_35380,N_35381,N_35382,N_35383,N_35384,N_35385,N_35386,N_35387,N_35388,N_35389,N_35390,N_35391,N_35392,N_35393,N_35394,N_35395,N_35396,N_35397,N_35398,N_35399,N_35400,N_35401,N_35402,N_35403,N_35404,N_35405,N_35406,N_35407,N_35408,N_35409,N_35410,N_35411,N_35412,N_35413,N_35414,N_35415,N_35416,N_35417,N_35418,N_35419,N_35420,N_35421,N_35422,N_35423,N_35424,N_35425,N_35426,N_35427,N_35428,N_35429,N_35430,N_35431,N_35432,N_35433,N_35434,N_35435,N_35436,N_35437,N_35438,N_35439,N_35440,N_35441,N_35442,N_35443,N_35444,N_35445,N_35446,N_35447,N_35448,N_35449,N_35450,N_35451,N_35452,N_35453,N_35454,N_35455,N_35456,N_35457,N_35458,N_35459,N_35460,N_35461,N_35462,N_35463,N_35464,N_35465,N_35466,N_35467,N_35468,N_35469,N_35470,N_35471,N_35472,N_35473,N_35474,N_35475,N_35476,N_35477,N_35478,N_35479,N_35480,N_35481,N_35482,N_35483,N_35484,N_35485,N_35486,N_35487,N_35488,N_35489,N_35490,N_35491,N_35492,N_35493,N_35494,N_35495,N_35496,N_35497,N_35498,N_35499,N_35500,N_35501,N_35502,N_35503,N_35504,N_35505,N_35506,N_35507,N_35508,N_35509,N_35510,N_35511,N_35512,N_35513,N_35514,N_35515,N_35516,N_35517,N_35518,N_35519,N_35520,N_35521,N_35522,N_35523,N_35524,N_35525,N_35526,N_35527,N_35528,N_35529,N_35530,N_35531,N_35532,N_35533,N_35534,N_35535,N_35536,N_35537,N_35538,N_35539,N_35540,N_35541,N_35542,N_35543,N_35544,N_35545,N_35546,N_35547,N_35548,N_35549,N_35550,N_35551,N_35552,N_35553,N_35554,N_35555,N_35556,N_35557,N_35558,N_35559,N_35560,N_35561,N_35562,N_35563,N_35564,N_35565,N_35566,N_35567,N_35568,N_35569,N_35570,N_35571,N_35572,N_35573,N_35574,N_35575,N_35576,N_35577,N_35578,N_35579,N_35580,N_35581,N_35582,N_35583,N_35584,N_35585,N_35586,N_35587,N_35588,N_35589,N_35590,N_35591,N_35592,N_35593,N_35594,N_35595,N_35596,N_35597,N_35598,N_35599,N_35600,N_35601,N_35602,N_35603,N_35604,N_35605,N_35606,N_35607,N_35608,N_35609,N_35610,N_35611,N_35612,N_35613,N_35614,N_35615,N_35616,N_35617,N_35618,N_35619,N_35620,N_35621,N_35622,N_35623,N_35624,N_35625,N_35626,N_35627,N_35628,N_35629,N_35630,N_35631,N_35632,N_35633,N_35634,N_35635,N_35636,N_35637,N_35638,N_35639,N_35640,N_35641,N_35642,N_35643,N_35644,N_35645,N_35646,N_35647,N_35648,N_35649,N_35650,N_35651,N_35652,N_35653,N_35654,N_35655,N_35656,N_35657,N_35658,N_35659,N_35660,N_35661,N_35662,N_35663,N_35664,N_35665,N_35666,N_35667,N_35668,N_35669,N_35670,N_35671,N_35672,N_35673,N_35674,N_35675,N_35676,N_35677,N_35678,N_35679,N_35680,N_35681,N_35682,N_35683,N_35684,N_35685,N_35686,N_35687,N_35688,N_35689,N_35690,N_35691,N_35692,N_35693,N_35694,N_35695,N_35696,N_35697,N_35698,N_35699,N_35700,N_35701,N_35702,N_35703,N_35704,N_35705,N_35706,N_35707,N_35708,N_35709,N_35710,N_35711,N_35712,N_35713,N_35714,N_35715,N_35716,N_35717,N_35718,N_35719,N_35720,N_35721,N_35722,N_35723,N_35724,N_35725,N_35726,N_35727,N_35728,N_35729,N_35730,N_35731,N_35732,N_35733,N_35734,N_35735,N_35736,N_35737,N_35738,N_35739,N_35740,N_35741,N_35742,N_35743,N_35744,N_35745,N_35746,N_35747,N_35748,N_35749,N_35750,N_35751,N_35752,N_35753,N_35754,N_35755,N_35756,N_35757,N_35758,N_35759,N_35760,N_35761,N_35762,N_35763,N_35764,N_35765,N_35766,N_35767,N_35768,N_35769,N_35770,N_35771,N_35772,N_35773,N_35774,N_35775,N_35776,N_35777,N_35778,N_35779,N_35780,N_35781,N_35782,N_35783,N_35784,N_35785,N_35786,N_35787,N_35788,N_35789,N_35790,N_35791,N_35792,N_35793,N_35794,N_35795,N_35796,N_35797,N_35798,N_35799,N_35800,N_35801,N_35802,N_35803,N_35804,N_35805,N_35806,N_35807,N_35808,N_35809,N_35810,N_35811,N_35812,N_35813,N_35814,N_35815,N_35816,N_35817,N_35818,N_35819,N_35820,N_35821,N_35822,N_35823,N_35824,N_35825,N_35826,N_35827,N_35828,N_35829,N_35830,N_35831,N_35832,N_35833,N_35834,N_35835,N_35836,N_35837,N_35838,N_35839,N_35840,N_35841,N_35842,N_35843,N_35844,N_35845,N_35846,N_35847,N_35848,N_35849,N_35850,N_35851,N_35852,N_35853,N_35854,N_35855,N_35856,N_35857,N_35858,N_35859,N_35860,N_35861,N_35862,N_35863,N_35864,N_35865,N_35866,N_35867,N_35868,N_35869,N_35870,N_35871,N_35872,N_35873,N_35874,N_35875,N_35876,N_35877,N_35878,N_35879,N_35880,N_35881,N_35882,N_35883,N_35884,N_35885,N_35886,N_35887,N_35888,N_35889,N_35890,N_35891,N_35892,N_35893,N_35894,N_35895,N_35896,N_35897,N_35898,N_35899,N_35900,N_35901,N_35902,N_35903,N_35904,N_35905,N_35906,N_35907,N_35908,N_35909,N_35910,N_35911,N_35912,N_35913,N_35914,N_35915,N_35916,N_35917,N_35918,N_35919,N_35920,N_35921,N_35922,N_35923,N_35924,N_35925,N_35926,N_35927,N_35928,N_35929,N_35930,N_35931,N_35932,N_35933,N_35934,N_35935,N_35936,N_35937,N_35938,N_35939,N_35940,N_35941,N_35942,N_35943,N_35944,N_35945,N_35946,N_35947,N_35948,N_35949,N_35950,N_35951,N_35952,N_35953,N_35954,N_35955,N_35956,N_35957,N_35958,N_35959,N_35960,N_35961,N_35962,N_35963,N_35964,N_35965,N_35966,N_35967,N_35968,N_35969,N_35970,N_35971,N_35972,N_35973,N_35974,N_35975,N_35976,N_35977,N_35978,N_35979,N_35980,N_35981,N_35982,N_35983,N_35984,N_35985,N_35986,N_35987,N_35988,N_35989,N_35990,N_35991,N_35992,N_35993,N_35994,N_35995,N_35996,N_35997,N_35998,N_35999,N_36000,N_36001,N_36002,N_36003,N_36004,N_36005,N_36006,N_36007,N_36008,N_36009,N_36010,N_36011,N_36012,N_36013,N_36014,N_36015,N_36016,N_36017,N_36018,N_36019,N_36020,N_36021,N_36022,N_36023,N_36024,N_36025,N_36026,N_36027,N_36028,N_36029,N_36030,N_36031,N_36032,N_36033,N_36034,N_36035,N_36036,N_36037,N_36038,N_36039,N_36040,N_36041,N_36042,N_36043,N_36044,N_36045,N_36046,N_36047,N_36048,N_36049,N_36050,N_36051,N_36052,N_36053,N_36054,N_36055,N_36056,N_36057,N_36058,N_36059,N_36060,N_36061,N_36062,N_36063,N_36064,N_36065,N_36066,N_36067,N_36068,N_36069,N_36070,N_36071,N_36072,N_36073,N_36074,N_36075,N_36076,N_36077,N_36078,N_36079,N_36080,N_36081,N_36082,N_36083,N_36084,N_36085,N_36086,N_36087,N_36088,N_36089,N_36090,N_36091,N_36092,N_36093,N_36094,N_36095,N_36096,N_36097,N_36098,N_36099,N_36100,N_36101,N_36102,N_36103,N_36104,N_36105,N_36106,N_36107,N_36108,N_36109,N_36110,N_36111,N_36112,N_36113,N_36114,N_36115,N_36116,N_36117,N_36118,N_36119,N_36120,N_36121,N_36122,N_36123,N_36124,N_36125,N_36126,N_36127,N_36128,N_36129,N_36130,N_36131,N_36132,N_36133,N_36134,N_36135,N_36136,N_36137,N_36138,N_36139,N_36140,N_36141,N_36142,N_36143,N_36144,N_36145,N_36146,N_36147,N_36148,N_36149,N_36150,N_36151,N_36152,N_36153,N_36154,N_36155,N_36156,N_36157,N_36158,N_36159,N_36160,N_36161,N_36162,N_36163,N_36164,N_36165,N_36166,N_36167,N_36168,N_36169,N_36170,N_36171,N_36172,N_36173,N_36174,N_36175,N_36176,N_36177,N_36178,N_36179,N_36180,N_36181,N_36182,N_36183,N_36184,N_36185,N_36186,N_36187,N_36188,N_36189,N_36190,N_36191,N_36192,N_36193,N_36194,N_36195,N_36196,N_36197,N_36198,N_36199,N_36200,N_36201,N_36202,N_36203,N_36204,N_36205,N_36206,N_36207,N_36208,N_36209,N_36210,N_36211,N_36212,N_36213,N_36214,N_36215,N_36216,N_36217,N_36218,N_36219,N_36220,N_36221,N_36222,N_36223,N_36224,N_36225,N_36226,N_36227,N_36228,N_36229,N_36230,N_36231,N_36232,N_36233,N_36234,N_36235,N_36236,N_36237,N_36238,N_36239,N_36240,N_36241,N_36242,N_36243,N_36244,N_36245,N_36246,N_36247,N_36248,N_36249,N_36250,N_36251,N_36252,N_36253,N_36254,N_36255,N_36256,N_36257,N_36258,N_36259,N_36260,N_36261,N_36262,N_36263,N_36264,N_36265,N_36266,N_36267,N_36268,N_36269,N_36270,N_36271,N_36272,N_36273,N_36274,N_36275,N_36276,N_36277,N_36278,N_36279,N_36280,N_36281,N_36282,N_36283,N_36284,N_36285,N_36286,N_36287,N_36288,N_36289,N_36290,N_36291,N_36292,N_36293,N_36294,N_36295,N_36296,N_36297,N_36298,N_36299,N_36300,N_36301,N_36302,N_36303,N_36304,N_36305,N_36306,N_36307,N_36308,N_36309,N_36310,N_36311,N_36312,N_36313,N_36314,N_36315,N_36316,N_36317,N_36318,N_36319,N_36320,N_36321,N_36322,N_36323,N_36324,N_36325,N_36326,N_36327,N_36328,N_36329,N_36330,N_36331,N_36332,N_36333,N_36334,N_36335,N_36336,N_36337,N_36338,N_36339,N_36340,N_36341,N_36342,N_36343,N_36344,N_36345,N_36346,N_36347,N_36348,N_36349,N_36350,N_36351,N_36352,N_36353,N_36354,N_36355,N_36356,N_36357,N_36358,N_36359,N_36360,N_36361,N_36362,N_36363,N_36364,N_36365,N_36366,N_36367,N_36368,N_36369,N_36370,N_36371,N_36372,N_36373,N_36374,N_36375,N_36376,N_36377,N_36378,N_36379,N_36380,N_36381,N_36382,N_36383,N_36384,N_36385,N_36386,N_36387,N_36388,N_36389,N_36390,N_36391,N_36392,N_36393,N_36394,N_36395,N_36396,N_36397,N_36398,N_36399,N_36400,N_36401,N_36402,N_36403,N_36404,N_36405,N_36406,N_36407,N_36408,N_36409,N_36410,N_36411,N_36412,N_36413,N_36414,N_36415,N_36416,N_36417,N_36418,N_36419,N_36420,N_36421,N_36422,N_36423,N_36424,N_36425,N_36426,N_36427,N_36428,N_36429,N_36430,N_36431,N_36432,N_36433,N_36434,N_36435,N_36436,N_36437,N_36438,N_36439,N_36440,N_36441,N_36442,N_36443,N_36444,N_36445,N_36446,N_36447,N_36448,N_36449,N_36450,N_36451,N_36452,N_36453,N_36454,N_36455,N_36456,N_36457,N_36458,N_36459,N_36460,N_36461,N_36462,N_36463,N_36464,N_36465,N_36466,N_36467,N_36468,N_36469,N_36470,N_36471,N_36472,N_36473,N_36474,N_36475,N_36476,N_36477,N_36478,N_36479,N_36480,N_36481,N_36482,N_36483,N_36484,N_36485,N_36486,N_36487,N_36488,N_36489,N_36490,N_36491,N_36492,N_36493,N_36494,N_36495,N_36496,N_36497,N_36498,N_36499,N_36500,N_36501,N_36502,N_36503,N_36504,N_36505,N_36506,N_36507,N_36508,N_36509,N_36510,N_36511,N_36512,N_36513,N_36514,N_36515,N_36516,N_36517,N_36518,N_36519,N_36520,N_36521,N_36522,N_36523,N_36524,N_36525,N_36526,N_36527,N_36528,N_36529,N_36530,N_36531,N_36532,N_36533,N_36534,N_36535,N_36536,N_36537,N_36538,N_36539,N_36540,N_36541,N_36542,N_36543,N_36544,N_36545,N_36546,N_36547,N_36548,N_36549,N_36550,N_36551,N_36552,N_36553,N_36554,N_36555,N_36556,N_36557,N_36558,N_36559,N_36560,N_36561,N_36562,N_36563,N_36564,N_36565,N_36566,N_36567,N_36568,N_36569,N_36570,N_36571,N_36572,N_36573,N_36574,N_36575,N_36576,N_36577,N_36578,N_36579,N_36580,N_36581,N_36582,N_36583,N_36584,N_36585,N_36586,N_36587,N_36588,N_36589,N_36590,N_36591,N_36592,N_36593,N_36594,N_36595,N_36596,N_36597,N_36598,N_36599,N_36600,N_36601,N_36602,N_36603,N_36604,N_36605,N_36606,N_36607,N_36608,N_36609,N_36610,N_36611,N_36612,N_36613,N_36614,N_36615,N_36616,N_36617,N_36618,N_36619,N_36620,N_36621,N_36622,N_36623,N_36624,N_36625,N_36626,N_36627,N_36628,N_36629,N_36630,N_36631,N_36632,N_36633,N_36634,N_36635,N_36636,N_36637,N_36638,N_36639,N_36640,N_36641,N_36642,N_36643,N_36644,N_36645,N_36646,N_36647,N_36648,N_36649,N_36650,N_36651,N_36652,N_36653,N_36654,N_36655,N_36656,N_36657,N_36658,N_36659,N_36660,N_36661,N_36662,N_36663,N_36664,N_36665,N_36666,N_36667,N_36668,N_36669,N_36670,N_36671,N_36672,N_36673,N_36674,N_36675,N_36676,N_36677,N_36678,N_36679,N_36680,N_36681,N_36682,N_36683,N_36684,N_36685,N_36686,N_36687,N_36688,N_36689,N_36690,N_36691,N_36692,N_36693,N_36694,N_36695,N_36696,N_36697,N_36698,N_36699,N_36700,N_36701,N_36702,N_36703,N_36704,N_36705,N_36706,N_36707,N_36708,N_36709,N_36710,N_36711,N_36712,N_36713,N_36714,N_36715,N_36716,N_36717,N_36718,N_36719,N_36720,N_36721,N_36722,N_36723,N_36724,N_36725,N_36726,N_36727,N_36728,N_36729,N_36730,N_36731,N_36732,N_36733,N_36734,N_36735,N_36736,N_36737,N_36738,N_36739,N_36740,N_36741,N_36742,N_36743,N_36744,N_36745,N_36746,N_36747,N_36748,N_36749,N_36750,N_36751,N_36752,N_36753,N_36754,N_36755,N_36756,N_36757,N_36758,N_36759,N_36760,N_36761,N_36762,N_36763,N_36764,N_36765,N_36766,N_36767,N_36768,N_36769,N_36770,N_36771,N_36772,N_36773,N_36774,N_36775,N_36776,N_36777,N_36778,N_36779,N_36780,N_36781,N_36782,N_36783,N_36784,N_36785,N_36786,N_36787,N_36788,N_36789,N_36790,N_36791,N_36792,N_36793,N_36794,N_36795,N_36796,N_36797,N_36798,N_36799,N_36800,N_36801,N_36802,N_36803,N_36804,N_36805,N_36806,N_36807,N_36808,N_36809,N_36810,N_36811,N_36812,N_36813,N_36814,N_36815,N_36816,N_36817,N_36818,N_36819,N_36820,N_36821,N_36822,N_36823,N_36824,N_36825,N_36826,N_36827,N_36828,N_36829,N_36830,N_36831,N_36832,N_36833,N_36834,N_36835,N_36836,N_36837,N_36838,N_36839,N_36840,N_36841,N_36842,N_36843,N_36844,N_36845,N_36846,N_36847,N_36848,N_36849,N_36850,N_36851,N_36852,N_36853,N_36854,N_36855,N_36856,N_36857,N_36858,N_36859,N_36860,N_36861,N_36862,N_36863,N_36864,N_36865,N_36866,N_36867,N_36868,N_36869,N_36870,N_36871,N_36872,N_36873,N_36874,N_36875,N_36876,N_36877,N_36878,N_36879,N_36880,N_36881,N_36882,N_36883,N_36884,N_36885,N_36886,N_36887,N_36888,N_36889,N_36890,N_36891,N_36892,N_36893,N_36894,N_36895,N_36896,N_36897,N_36898,N_36899,N_36900,N_36901,N_36902,N_36903,N_36904,N_36905,N_36906,N_36907,N_36908,N_36909,N_36910,N_36911,N_36912,N_36913,N_36914,N_36915,N_36916,N_36917,N_36918,N_36919,N_36920,N_36921,N_36922,N_36923,N_36924,N_36925,N_36926,N_36927,N_36928,N_36929,N_36930,N_36931,N_36932,N_36933,N_36934,N_36935,N_36936,N_36937,N_36938,N_36939,N_36940,N_36941,N_36942,N_36943,N_36944,N_36945,N_36946,N_36947,N_36948,N_36949,N_36950,N_36951,N_36952,N_36953,N_36954,N_36955,N_36956,N_36957,N_36958,N_36959,N_36960,N_36961,N_36962,N_36963,N_36964,N_36965,N_36966,N_36967,N_36968,N_36969,N_36970,N_36971,N_36972,N_36973,N_36974,N_36975,N_36976,N_36977,N_36978,N_36979,N_36980,N_36981,N_36982,N_36983,N_36984,N_36985,N_36986,N_36987,N_36988,N_36989,N_36990,N_36991,N_36992,N_36993,N_36994,N_36995,N_36996,N_36997,N_36998,N_36999,N_37000,N_37001,N_37002,N_37003,N_37004,N_37005,N_37006,N_37007,N_37008,N_37009,N_37010,N_37011,N_37012,N_37013,N_37014,N_37015,N_37016,N_37017,N_37018,N_37019,N_37020,N_37021,N_37022,N_37023,N_37024,N_37025,N_37026,N_37027,N_37028,N_37029,N_37030,N_37031,N_37032,N_37033,N_37034,N_37035,N_37036,N_37037,N_37038,N_37039,N_37040,N_37041,N_37042,N_37043,N_37044,N_37045,N_37046,N_37047,N_37048,N_37049,N_37050,N_37051,N_37052,N_37053,N_37054,N_37055,N_37056,N_37057,N_37058,N_37059,N_37060,N_37061,N_37062,N_37063,N_37064,N_37065,N_37066,N_37067,N_37068,N_37069,N_37070,N_37071,N_37072,N_37073,N_37074,N_37075,N_37076,N_37077,N_37078,N_37079,N_37080,N_37081,N_37082,N_37083,N_37084,N_37085,N_37086,N_37087,N_37088,N_37089,N_37090,N_37091,N_37092,N_37093,N_37094,N_37095,N_37096,N_37097,N_37098,N_37099,N_37100,N_37101,N_37102,N_37103,N_37104,N_37105,N_37106,N_37107,N_37108,N_37109,N_37110,N_37111,N_37112,N_37113,N_37114,N_37115,N_37116,N_37117,N_37118,N_37119,N_37120,N_37121,N_37122,N_37123,N_37124,N_37125,N_37126,N_37127,N_37128,N_37129,N_37130,N_37131,N_37132,N_37133,N_37134,N_37135,N_37136,N_37137,N_37138,N_37139,N_37140,N_37141,N_37142,N_37143,N_37144,N_37145,N_37146,N_37147,N_37148,N_37149,N_37150,N_37151,N_37152,N_37153,N_37154,N_37155,N_37156,N_37157,N_37158,N_37159,N_37160,N_37161,N_37162,N_37163,N_37164,N_37165,N_37166,N_37167,N_37168,N_37169,N_37170,N_37171,N_37172,N_37173,N_37174,N_37175,N_37176,N_37177,N_37178,N_37179,N_37180,N_37181,N_37182,N_37183,N_37184,N_37185,N_37186,N_37187,N_37188,N_37189,N_37190,N_37191,N_37192,N_37193,N_37194,N_37195,N_37196,N_37197,N_37198,N_37199,N_37200,N_37201,N_37202,N_37203,N_37204,N_37205,N_37206,N_37207,N_37208,N_37209,N_37210,N_37211,N_37212,N_37213,N_37214,N_37215,N_37216,N_37217,N_37218,N_37219,N_37220,N_37221,N_37222,N_37223,N_37224,N_37225,N_37226,N_37227,N_37228,N_37229,N_37230,N_37231,N_37232,N_37233,N_37234,N_37235,N_37236,N_37237,N_37238,N_37239,N_37240,N_37241,N_37242,N_37243,N_37244,N_37245,N_37246,N_37247,N_37248,N_37249,N_37250,N_37251,N_37252,N_37253,N_37254,N_37255,N_37256,N_37257,N_37258,N_37259,N_37260,N_37261,N_37262,N_37263,N_37264,N_37265,N_37266,N_37267,N_37268,N_37269,N_37270,N_37271,N_37272,N_37273,N_37274,N_37275,N_37276,N_37277,N_37278,N_37279,N_37280,N_37281,N_37282,N_37283,N_37284,N_37285,N_37286,N_37287,N_37288,N_37289,N_37290,N_37291,N_37292,N_37293,N_37294,N_37295,N_37296,N_37297,N_37298,N_37299,N_37300,N_37301,N_37302,N_37303,N_37304,N_37305,N_37306,N_37307,N_37308,N_37309,N_37310,N_37311,N_37312,N_37313,N_37314,N_37315,N_37316,N_37317,N_37318,N_37319,N_37320,N_37321,N_37322,N_37323,N_37324,N_37325,N_37326,N_37327,N_37328,N_37329,N_37330,N_37331,N_37332,N_37333,N_37334,N_37335,N_37336,N_37337,N_37338,N_37339,N_37340,N_37341,N_37342,N_37343,N_37344,N_37345,N_37346,N_37347,N_37348,N_37349,N_37350,N_37351,N_37352,N_37353,N_37354,N_37355,N_37356,N_37357,N_37358,N_37359,N_37360,N_37361,N_37362,N_37363,N_37364,N_37365,N_37366,N_37367,N_37368,N_37369,N_37370,N_37371,N_37372,N_37373,N_37374,N_37375,N_37376,N_37377,N_37378,N_37379,N_37380,N_37381,N_37382,N_37383,N_37384,N_37385,N_37386,N_37387,N_37388,N_37389,N_37390,N_37391,N_37392,N_37393,N_37394,N_37395,N_37396,N_37397,N_37398,N_37399,N_37400,N_37401,N_37402,N_37403,N_37404,N_37405,N_37406,N_37407,N_37408,N_37409,N_37410,N_37411,N_37412,N_37413,N_37414,N_37415,N_37416,N_37417,N_37418,N_37419,N_37420,N_37421,N_37422,N_37423,N_37424,N_37425,N_37426,N_37427,N_37428,N_37429,N_37430,N_37431,N_37432,N_37433,N_37434,N_37435,N_37436,N_37437,N_37438,N_37439,N_37440,N_37441,N_37442,N_37443,N_37444,N_37445,N_37446,N_37447,N_37448,N_37449,N_37450,N_37451,N_37452,N_37453,N_37454,N_37455,N_37456,N_37457,N_37458,N_37459,N_37460,N_37461,N_37462,N_37463,N_37464,N_37465,N_37466,N_37467,N_37468,N_37469,N_37470,N_37471,N_37472,N_37473,N_37474,N_37475,N_37476,N_37477,N_37478,N_37479,N_37480,N_37481,N_37482,N_37483,N_37484,N_37485,N_37486,N_37487,N_37488,N_37489,N_37490,N_37491,N_37492,N_37493,N_37494,N_37495,N_37496,N_37497,N_37498,N_37499,N_37500,N_37501,N_37502,N_37503,N_37504,N_37505,N_37506,N_37507,N_37508,N_37509,N_37510,N_37511,N_37512,N_37513,N_37514,N_37515,N_37516,N_37517,N_37518,N_37519,N_37520,N_37521,N_37522,N_37523,N_37524,N_37525,N_37526,N_37527,N_37528,N_37529,N_37530,N_37531,N_37532,N_37533,N_37534,N_37535,N_37536,N_37537,N_37538,N_37539,N_37540,N_37541,N_37542,N_37543,N_37544,N_37545,N_37546,N_37547,N_37548,N_37549,N_37550,N_37551,N_37552,N_37553,N_37554,N_37555,N_37556,N_37557,N_37558,N_37559,N_37560,N_37561,N_37562,N_37563,N_37564,N_37565,N_37566,N_37567,N_37568,N_37569,N_37570,N_37571,N_37572,N_37573,N_37574,N_37575,N_37576,N_37577,N_37578,N_37579,N_37580,N_37581,N_37582,N_37583,N_37584,N_37585,N_37586,N_37587,N_37588,N_37589,N_37590,N_37591,N_37592,N_37593,N_37594,N_37595,N_37596,N_37597,N_37598,N_37599,N_37600,N_37601,N_37602,N_37603,N_37604,N_37605,N_37606,N_37607,N_37608,N_37609,N_37610,N_37611,N_37612,N_37613,N_37614,N_37615,N_37616,N_37617,N_37618,N_37619,N_37620,N_37621,N_37622,N_37623,N_37624,N_37625,N_37626,N_37627,N_37628,N_37629,N_37630,N_37631,N_37632,N_37633,N_37634,N_37635,N_37636,N_37637,N_37638,N_37639,N_37640,N_37641,N_37642,N_37643,N_37644,N_37645,N_37646,N_37647,N_37648,N_37649,N_37650,N_37651,N_37652,N_37653,N_37654,N_37655,N_37656,N_37657,N_37658,N_37659,N_37660,N_37661,N_37662,N_37663,N_37664,N_37665,N_37666,N_37667,N_37668,N_37669,N_37670,N_37671,N_37672,N_37673,N_37674,N_37675,N_37676,N_37677,N_37678,N_37679,N_37680,N_37681,N_37682,N_37683,N_37684,N_37685,N_37686,N_37687,N_37688,N_37689,N_37690,N_37691,N_37692,N_37693,N_37694,N_37695,N_37696,N_37697,N_37698,N_37699,N_37700,N_37701,N_37702,N_37703,N_37704,N_37705,N_37706,N_37707,N_37708,N_37709,N_37710,N_37711,N_37712,N_37713,N_37714,N_37715,N_37716,N_37717,N_37718,N_37719,N_37720,N_37721,N_37722,N_37723,N_37724,N_37725,N_37726,N_37727,N_37728,N_37729,N_37730,N_37731,N_37732,N_37733,N_37734,N_37735,N_37736,N_37737,N_37738,N_37739,N_37740,N_37741,N_37742,N_37743,N_37744,N_37745,N_37746,N_37747,N_37748,N_37749,N_37750,N_37751,N_37752,N_37753,N_37754,N_37755,N_37756,N_37757,N_37758,N_37759,N_37760,N_37761,N_37762,N_37763,N_37764,N_37765,N_37766,N_37767,N_37768,N_37769,N_37770,N_37771,N_37772,N_37773,N_37774,N_37775,N_37776,N_37777,N_37778,N_37779,N_37780,N_37781,N_37782,N_37783,N_37784,N_37785,N_37786,N_37787,N_37788,N_37789,N_37790,N_37791,N_37792,N_37793,N_37794,N_37795,N_37796,N_37797,N_37798,N_37799,N_37800,N_37801,N_37802,N_37803,N_37804,N_37805,N_37806,N_37807,N_37808,N_37809,N_37810,N_37811,N_37812,N_37813,N_37814,N_37815,N_37816,N_37817,N_37818,N_37819,N_37820,N_37821,N_37822,N_37823,N_37824,N_37825,N_37826,N_37827,N_37828,N_37829,N_37830,N_37831,N_37832,N_37833,N_37834,N_37835,N_37836,N_37837,N_37838,N_37839,N_37840,N_37841,N_37842,N_37843,N_37844,N_37845,N_37846,N_37847,N_37848,N_37849,N_37850,N_37851,N_37852,N_37853,N_37854,N_37855,N_37856,N_37857,N_37858,N_37859,N_37860,N_37861,N_37862,N_37863,N_37864,N_37865,N_37866,N_37867,N_37868,N_37869,N_37870,N_37871,N_37872,N_37873,N_37874,N_37875,N_37876,N_37877,N_37878,N_37879,N_37880,N_37881,N_37882,N_37883,N_37884,N_37885,N_37886,N_37887,N_37888,N_37889,N_37890,N_37891,N_37892,N_37893,N_37894,N_37895,N_37896,N_37897,N_37898,N_37899,N_37900,N_37901,N_37902,N_37903,N_37904,N_37905,N_37906,N_37907,N_37908,N_37909,N_37910,N_37911,N_37912,N_37913,N_37914,N_37915,N_37916,N_37917,N_37918,N_37919,N_37920,N_37921,N_37922,N_37923,N_37924,N_37925,N_37926,N_37927,N_37928,N_37929,N_37930,N_37931,N_37932,N_37933,N_37934,N_37935,N_37936,N_37937,N_37938,N_37939,N_37940,N_37941,N_37942,N_37943,N_37944,N_37945,N_37946,N_37947,N_37948,N_37949,N_37950,N_37951,N_37952,N_37953,N_37954,N_37955,N_37956,N_37957,N_37958,N_37959,N_37960,N_37961,N_37962,N_37963,N_37964,N_37965,N_37966,N_37967,N_37968,N_37969,N_37970,N_37971,N_37972,N_37973,N_37974,N_37975,N_37976,N_37977,N_37978,N_37979,N_37980,N_37981,N_37982,N_37983,N_37984,N_37985,N_37986,N_37987,N_37988,N_37989,N_37990,N_37991,N_37992,N_37993,N_37994,N_37995,N_37996,N_37997,N_37998,N_37999,N_38000,N_38001,N_38002,N_38003,N_38004,N_38005,N_38006,N_38007,N_38008,N_38009,N_38010,N_38011,N_38012,N_38013,N_38014,N_38015,N_38016,N_38017,N_38018,N_38019,N_38020,N_38021,N_38022,N_38023,N_38024,N_38025,N_38026,N_38027,N_38028,N_38029,N_38030,N_38031,N_38032,N_38033,N_38034,N_38035,N_38036,N_38037,N_38038,N_38039,N_38040,N_38041,N_38042,N_38043,N_38044,N_38045,N_38046,N_38047,N_38048,N_38049,N_38050,N_38051,N_38052,N_38053,N_38054,N_38055,N_38056,N_38057,N_38058,N_38059,N_38060,N_38061,N_38062,N_38063,N_38064,N_38065,N_38066,N_38067,N_38068,N_38069,N_38070,N_38071,N_38072,N_38073,N_38074,N_38075,N_38076,N_38077,N_38078,N_38079,N_38080,N_38081,N_38082,N_38083,N_38084,N_38085,N_38086,N_38087,N_38088,N_38089,N_38090,N_38091,N_38092,N_38093,N_38094,N_38095,N_38096,N_38097,N_38098,N_38099,N_38100,N_38101,N_38102,N_38103,N_38104,N_38105,N_38106,N_38107,N_38108,N_38109,N_38110,N_38111,N_38112,N_38113,N_38114,N_38115,N_38116,N_38117,N_38118,N_38119,N_38120,N_38121,N_38122,N_38123,N_38124,N_38125,N_38126,N_38127,N_38128,N_38129,N_38130,N_38131,N_38132,N_38133,N_38134,N_38135,N_38136,N_38137,N_38138,N_38139,N_38140,N_38141,N_38142,N_38143,N_38144,N_38145,N_38146,N_38147,N_38148,N_38149,N_38150,N_38151,N_38152,N_38153,N_38154,N_38155,N_38156,N_38157,N_38158,N_38159,N_38160,N_38161,N_38162,N_38163,N_38164,N_38165,N_38166,N_38167,N_38168,N_38169,N_38170,N_38171,N_38172,N_38173,N_38174,N_38175,N_38176,N_38177,N_38178,N_38179,N_38180,N_38181,N_38182,N_38183,N_38184,N_38185,N_38186,N_38187,N_38188,N_38189,N_38190,N_38191,N_38192,N_38193,N_38194,N_38195,N_38196,N_38197,N_38198,N_38199,N_38200,N_38201,N_38202,N_38203,N_38204,N_38205,N_38206,N_38207,N_38208,N_38209,N_38210,N_38211,N_38212,N_38213,N_38214,N_38215,N_38216,N_38217,N_38218,N_38219,N_38220,N_38221,N_38222,N_38223,N_38224,N_38225,N_38226,N_38227,N_38228,N_38229,N_38230,N_38231,N_38232,N_38233,N_38234,N_38235,N_38236,N_38237,N_38238,N_38239,N_38240,N_38241,N_38242,N_38243,N_38244,N_38245,N_38246,N_38247,N_38248,N_38249,N_38250,N_38251,N_38252,N_38253,N_38254,N_38255,N_38256,N_38257,N_38258,N_38259,N_38260,N_38261,N_38262,N_38263,N_38264,N_38265,N_38266,N_38267,N_38268,N_38269,N_38270,N_38271,N_38272,N_38273,N_38274,N_38275,N_38276,N_38277,N_38278,N_38279,N_38280,N_38281,N_38282,N_38283,N_38284,N_38285,N_38286,N_38287,N_38288,N_38289,N_38290,N_38291,N_38292,N_38293,N_38294,N_38295,N_38296,N_38297,N_38298,N_38299,N_38300,N_38301,N_38302,N_38303,N_38304,N_38305,N_38306,N_38307,N_38308,N_38309,N_38310,N_38311,N_38312,N_38313,N_38314,N_38315,N_38316,N_38317,N_38318,N_38319,N_38320,N_38321,N_38322,N_38323,N_38324,N_38325,N_38326,N_38327,N_38328,N_38329,N_38330,N_38331,N_38332,N_38333,N_38334,N_38335,N_38336,N_38337,N_38338,N_38339,N_38340,N_38341,N_38342,N_38343,N_38344,N_38345,N_38346,N_38347,N_38348,N_38349,N_38350,N_38351,N_38352,N_38353,N_38354,N_38355,N_38356,N_38357,N_38358,N_38359,N_38360,N_38361,N_38362,N_38363,N_38364,N_38365,N_38366,N_38367,N_38368,N_38369,N_38370,N_38371,N_38372,N_38373,N_38374,N_38375,N_38376,N_38377,N_38378,N_38379,N_38380,N_38381,N_38382,N_38383,N_38384,N_38385,N_38386,N_38387,N_38388,N_38389,N_38390,N_38391,N_38392,N_38393,N_38394,N_38395,N_38396,N_38397,N_38398,N_38399,N_38400,N_38401,N_38402,N_38403,N_38404,N_38405,N_38406,N_38407,N_38408,N_38409,N_38410,N_38411,N_38412,N_38413,N_38414,N_38415,N_38416,N_38417,N_38418,N_38419,N_38420,N_38421,N_38422,N_38423,N_38424,N_38425,N_38426,N_38427,N_38428,N_38429,N_38430,N_38431,N_38432,N_38433,N_38434,N_38435,N_38436,N_38437,N_38438,N_38439,N_38440,N_38441,N_38442,N_38443,N_38444,N_38445,N_38446,N_38447,N_38448,N_38449,N_38450,N_38451,N_38452,N_38453,N_38454,N_38455,N_38456,N_38457,N_38458,N_38459,N_38460,N_38461,N_38462,N_38463,N_38464,N_38465,N_38466,N_38467,N_38468,N_38469,N_38470,N_38471,N_38472,N_38473,N_38474,N_38475,N_38476,N_38477,N_38478,N_38479,N_38480,N_38481,N_38482,N_38483,N_38484,N_38485,N_38486,N_38487,N_38488,N_38489,N_38490,N_38491,N_38492,N_38493,N_38494,N_38495,N_38496,N_38497,N_38498,N_38499,N_38500,N_38501,N_38502,N_38503,N_38504,N_38505,N_38506,N_38507,N_38508,N_38509,N_38510,N_38511,N_38512,N_38513,N_38514,N_38515,N_38516,N_38517,N_38518,N_38519,N_38520,N_38521,N_38522,N_38523,N_38524,N_38525,N_38526,N_38527,N_38528,N_38529,N_38530,N_38531,N_38532,N_38533,N_38534,N_38535,N_38536,N_38537,N_38538,N_38539,N_38540,N_38541,N_38542,N_38543,N_38544,N_38545,N_38546,N_38547,N_38548,N_38549,N_38550,N_38551,N_38552,N_38553,N_38554,N_38555,N_38556,N_38557,N_38558,N_38559,N_38560,N_38561,N_38562,N_38563,N_38564,N_38565,N_38566,N_38567,N_38568,N_38569,N_38570,N_38571,N_38572,N_38573,N_38574,N_38575,N_38576,N_38577,N_38578,N_38579,N_38580,N_38581,N_38582,N_38583,N_38584,N_38585,N_38586,N_38587,N_38588,N_38589,N_38590,N_38591,N_38592,N_38593,N_38594,N_38595,N_38596,N_38597,N_38598,N_38599,N_38600,N_38601,N_38602,N_38603,N_38604,N_38605,N_38606,N_38607,N_38608,N_38609,N_38610,N_38611,N_38612,N_38613,N_38614,N_38615,N_38616,N_38617,N_38618,N_38619,N_38620,N_38621,N_38622,N_38623,N_38624,N_38625,N_38626,N_38627,N_38628,N_38629,N_38630,N_38631,N_38632,N_38633,N_38634,N_38635,N_38636,N_38637,N_38638,N_38639,N_38640,N_38641,N_38642,N_38643,N_38644,N_38645,N_38646,N_38647,N_38648,N_38649,N_38650,N_38651,N_38652,N_38653,N_38654,N_38655,N_38656,N_38657,N_38658,N_38659,N_38660,N_38661,N_38662,N_38663,N_38664,N_38665,N_38666,N_38667,N_38668,N_38669,N_38670,N_38671,N_38672,N_38673,N_38674,N_38675,N_38676,N_38677,N_38678,N_38679,N_38680,N_38681,N_38682,N_38683,N_38684,N_38685,N_38686,N_38687,N_38688,N_38689,N_38690,N_38691,N_38692,N_38693,N_38694,N_38695,N_38696,N_38697,N_38698,N_38699,N_38700,N_38701,N_38702,N_38703,N_38704,N_38705,N_38706,N_38707,N_38708,N_38709,N_38710,N_38711,N_38712,N_38713,N_38714,N_38715,N_38716,N_38717,N_38718,N_38719,N_38720,N_38721,N_38722,N_38723,N_38724,N_38725,N_38726,N_38727,N_38728,N_38729,N_38730,N_38731,N_38732,N_38733,N_38734,N_38735,N_38736,N_38737,N_38738,N_38739,N_38740,N_38741,N_38742,N_38743,N_38744,N_38745,N_38746,N_38747,N_38748,N_38749,N_38750,N_38751,N_38752,N_38753,N_38754,N_38755,N_38756,N_38757,N_38758,N_38759,N_38760,N_38761,N_38762,N_38763,N_38764,N_38765,N_38766,N_38767,N_38768,N_38769,N_38770,N_38771,N_38772,N_38773,N_38774,N_38775,N_38776,N_38777,N_38778,N_38779,N_38780,N_38781,N_38782,N_38783,N_38784,N_38785,N_38786,N_38787,N_38788,N_38789,N_38790,N_38791,N_38792,N_38793,N_38794,N_38795,N_38796,N_38797,N_38798,N_38799,N_38800,N_38801,N_38802,N_38803,N_38804,N_38805,N_38806,N_38807,N_38808,N_38809,N_38810,N_38811,N_38812,N_38813,N_38814,N_38815,N_38816,N_38817,N_38818,N_38819,N_38820,N_38821,N_38822,N_38823,N_38824,N_38825,N_38826,N_38827,N_38828,N_38829,N_38830,N_38831,N_38832,N_38833,N_38834,N_38835,N_38836,N_38837,N_38838,N_38839,N_38840,N_38841,N_38842,N_38843,N_38844,N_38845,N_38846,N_38847,N_38848,N_38849,N_38850,N_38851,N_38852,N_38853,N_38854,N_38855,N_38856,N_38857,N_38858,N_38859,N_38860,N_38861,N_38862,N_38863,N_38864,N_38865,N_38866,N_38867,N_38868,N_38869,N_38870,N_38871,N_38872,N_38873,N_38874,N_38875,N_38876,N_38877,N_38878,N_38879,N_38880,N_38881,N_38882,N_38883,N_38884,N_38885,N_38886,N_38887,N_38888,N_38889,N_38890,N_38891,N_38892,N_38893,N_38894,N_38895,N_38896,N_38897,N_38898,N_38899,N_38900,N_38901,N_38902,N_38903,N_38904,N_38905,N_38906,N_38907,N_38908,N_38909,N_38910,N_38911,N_38912,N_38913,N_38914,N_38915,N_38916,N_38917,N_38918,N_38919,N_38920,N_38921,N_38922,N_38923,N_38924,N_38925,N_38926,N_38927,N_38928,N_38929,N_38930,N_38931,N_38932,N_38933,N_38934,N_38935,N_38936,N_38937,N_38938,N_38939,N_38940,N_38941,N_38942,N_38943,N_38944,N_38945,N_38946,N_38947,N_38948,N_38949,N_38950,N_38951,N_38952,N_38953,N_38954,N_38955,N_38956,N_38957,N_38958,N_38959,N_38960,N_38961,N_38962,N_38963,N_38964,N_38965,N_38966,N_38967,N_38968,N_38969,N_38970,N_38971,N_38972,N_38973,N_38974,N_38975,N_38976,N_38977,N_38978,N_38979,N_38980,N_38981,N_38982,N_38983,N_38984,N_38985,N_38986,N_38987,N_38988,N_38989,N_38990,N_38991,N_38992,N_38993,N_38994,N_38995,N_38996,N_38997,N_38998,N_38999,N_39000,N_39001,N_39002,N_39003,N_39004,N_39005,N_39006,N_39007,N_39008,N_39009,N_39010,N_39011,N_39012,N_39013,N_39014,N_39015,N_39016,N_39017,N_39018,N_39019,N_39020,N_39021,N_39022,N_39023,N_39024,N_39025,N_39026,N_39027,N_39028,N_39029,N_39030,N_39031,N_39032,N_39033,N_39034,N_39035,N_39036,N_39037,N_39038,N_39039,N_39040,N_39041,N_39042,N_39043,N_39044,N_39045,N_39046,N_39047,N_39048,N_39049,N_39050,N_39051,N_39052,N_39053,N_39054,N_39055,N_39056,N_39057,N_39058,N_39059,N_39060,N_39061,N_39062,N_39063,N_39064,N_39065,N_39066,N_39067,N_39068,N_39069,N_39070,N_39071,N_39072,N_39073,N_39074,N_39075,N_39076,N_39077,N_39078,N_39079,N_39080,N_39081,N_39082,N_39083,N_39084,N_39085,N_39086,N_39087,N_39088,N_39089,N_39090,N_39091,N_39092,N_39093,N_39094,N_39095,N_39096,N_39097,N_39098,N_39099,N_39100,N_39101,N_39102,N_39103,N_39104,N_39105,N_39106,N_39107,N_39108,N_39109,N_39110,N_39111,N_39112,N_39113,N_39114,N_39115,N_39116,N_39117,N_39118,N_39119,N_39120,N_39121,N_39122,N_39123,N_39124,N_39125,N_39126,N_39127,N_39128,N_39129,N_39130,N_39131,N_39132,N_39133,N_39134,N_39135,N_39136,N_39137,N_39138,N_39139,N_39140,N_39141,N_39142,N_39143,N_39144,N_39145,N_39146,N_39147,N_39148,N_39149,N_39150,N_39151,N_39152,N_39153,N_39154,N_39155,N_39156,N_39157,N_39158,N_39159,N_39160,N_39161,N_39162,N_39163,N_39164,N_39165,N_39166,N_39167,N_39168,N_39169,N_39170,N_39171,N_39172,N_39173,N_39174,N_39175,N_39176,N_39177,N_39178,N_39179,N_39180,N_39181,N_39182,N_39183,N_39184,N_39185,N_39186,N_39187,N_39188,N_39189,N_39190,N_39191,N_39192,N_39193,N_39194,N_39195,N_39196,N_39197,N_39198,N_39199,N_39200,N_39201,N_39202,N_39203,N_39204,N_39205,N_39206,N_39207,N_39208,N_39209,N_39210,N_39211,N_39212,N_39213,N_39214,N_39215,N_39216,N_39217,N_39218,N_39219,N_39220,N_39221,N_39222,N_39223,N_39224,N_39225,N_39226,N_39227,N_39228,N_39229,N_39230,N_39231,N_39232,N_39233,N_39234,N_39235,N_39236,N_39237,N_39238,N_39239,N_39240,N_39241,N_39242,N_39243,N_39244,N_39245,N_39246,N_39247,N_39248,N_39249,N_39250,N_39251,N_39252,N_39253,N_39254,N_39255,N_39256,N_39257,N_39258,N_39259,N_39260,N_39261,N_39262,N_39263,N_39264,N_39265,N_39266,N_39267,N_39268,N_39269,N_39270,N_39271,N_39272,N_39273,N_39274,N_39275,N_39276,N_39277,N_39278,N_39279,N_39280,N_39281,N_39282,N_39283,N_39284,N_39285,N_39286,N_39287,N_39288,N_39289,N_39290,N_39291,N_39292,N_39293,N_39294,N_39295,N_39296,N_39297,N_39298,N_39299,N_39300,N_39301,N_39302,N_39303,N_39304,N_39305,N_39306,N_39307,N_39308,N_39309,N_39310,N_39311,N_39312,N_39313,N_39314,N_39315,N_39316,N_39317,N_39318,N_39319,N_39320,N_39321,N_39322,N_39323,N_39324,N_39325,N_39326,N_39327,N_39328,N_39329,N_39330,N_39331,N_39332,N_39333,N_39334,N_39335,N_39336,N_39337,N_39338,N_39339,N_39340,N_39341,N_39342,N_39343,N_39344,N_39345,N_39346,N_39347,N_39348,N_39349,N_39350,N_39351,N_39352,N_39353,N_39354,N_39355,N_39356,N_39357,N_39358,N_39359,N_39360,N_39361,N_39362,N_39363,N_39364,N_39365,N_39366,N_39367,N_39368,N_39369,N_39370,N_39371,N_39372,N_39373,N_39374,N_39375,N_39376,N_39377,N_39378,N_39379,N_39380,N_39381,N_39382,N_39383,N_39384,N_39385,N_39386,N_39387,N_39388,N_39389,N_39390,N_39391,N_39392,N_39393,N_39394,N_39395,N_39396,N_39397,N_39398,N_39399,N_39400,N_39401,N_39402,N_39403,N_39404,N_39405,N_39406,N_39407,N_39408,N_39409,N_39410,N_39411,N_39412,N_39413,N_39414,N_39415,N_39416,N_39417,N_39418,N_39419,N_39420,N_39421,N_39422,N_39423,N_39424,N_39425,N_39426,N_39427,N_39428,N_39429,N_39430,N_39431,N_39432,N_39433,N_39434,N_39435,N_39436,N_39437,N_39438,N_39439,N_39440,N_39441,N_39442,N_39443,N_39444,N_39445,N_39446,N_39447,N_39448,N_39449,N_39450,N_39451,N_39452,N_39453,N_39454,N_39455,N_39456,N_39457,N_39458,N_39459,N_39460,N_39461,N_39462,N_39463,N_39464,N_39465,N_39466,N_39467,N_39468,N_39469,N_39470,N_39471,N_39472,N_39473,N_39474,N_39475,N_39476,N_39477,N_39478,N_39479,N_39480,N_39481,N_39482,N_39483,N_39484,N_39485,N_39486,N_39487,N_39488,N_39489,N_39490,N_39491,N_39492,N_39493,N_39494,N_39495,N_39496,N_39497,N_39498,N_39499,N_39500,N_39501,N_39502,N_39503,N_39504,N_39505,N_39506,N_39507,N_39508,N_39509,N_39510,N_39511,N_39512,N_39513,N_39514,N_39515,N_39516,N_39517,N_39518,N_39519,N_39520,N_39521,N_39522,N_39523,N_39524,N_39525,N_39526,N_39527,N_39528,N_39529,N_39530,N_39531,N_39532,N_39533,N_39534,N_39535,N_39536,N_39537,N_39538,N_39539,N_39540,N_39541,N_39542,N_39543,N_39544,N_39545,N_39546,N_39547,N_39548,N_39549,N_39550,N_39551,N_39552,N_39553,N_39554,N_39555,N_39556,N_39557,N_39558,N_39559,N_39560,N_39561,N_39562,N_39563,N_39564,N_39565,N_39566,N_39567,N_39568,N_39569,N_39570,N_39571,N_39572,N_39573,N_39574,N_39575,N_39576,N_39577,N_39578,N_39579,N_39580,N_39581,N_39582,N_39583,N_39584,N_39585,N_39586,N_39587,N_39588,N_39589,N_39590,N_39591,N_39592,N_39593,N_39594,N_39595,N_39596,N_39597,N_39598,N_39599,N_39600,N_39601,N_39602,N_39603,N_39604,N_39605,N_39606,N_39607,N_39608,N_39609,N_39610,N_39611,N_39612,N_39613,N_39614,N_39615,N_39616,N_39617,N_39618,N_39619,N_39620,N_39621,N_39622,N_39623,N_39624,N_39625,N_39626,N_39627,N_39628,N_39629,N_39630,N_39631,N_39632,N_39633,N_39634,N_39635,N_39636,N_39637,N_39638,N_39639,N_39640,N_39641,N_39642,N_39643,N_39644,N_39645,N_39646,N_39647,N_39648,N_39649,N_39650,N_39651,N_39652,N_39653,N_39654,N_39655,N_39656,N_39657,N_39658,N_39659,N_39660,N_39661,N_39662,N_39663,N_39664,N_39665,N_39666,N_39667,N_39668,N_39669,N_39670,N_39671,N_39672,N_39673,N_39674,N_39675,N_39676,N_39677,N_39678,N_39679,N_39680,N_39681,N_39682,N_39683,N_39684,N_39685,N_39686,N_39687,N_39688,N_39689,N_39690,N_39691,N_39692,N_39693,N_39694,N_39695,N_39696,N_39697,N_39698,N_39699,N_39700,N_39701,N_39702,N_39703,N_39704,N_39705,N_39706,N_39707,N_39708,N_39709,N_39710,N_39711,N_39712,N_39713,N_39714,N_39715,N_39716,N_39717,N_39718,N_39719,N_39720,N_39721,N_39722,N_39723,N_39724,N_39725,N_39726,N_39727,N_39728,N_39729,N_39730,N_39731,N_39732,N_39733,N_39734,N_39735,N_39736,N_39737,N_39738,N_39739,N_39740,N_39741,N_39742,N_39743,N_39744,N_39745,N_39746,N_39747,N_39748,N_39749,N_39750,N_39751,N_39752,N_39753,N_39754,N_39755,N_39756,N_39757,N_39758,N_39759,N_39760,N_39761,N_39762,N_39763,N_39764,N_39765,N_39766,N_39767,N_39768,N_39769,N_39770,N_39771,N_39772,N_39773,N_39774,N_39775,N_39776,N_39777,N_39778,N_39779,N_39780,N_39781,N_39782,N_39783,N_39784,N_39785,N_39786,N_39787,N_39788,N_39789,N_39790,N_39791,N_39792,N_39793,N_39794,N_39795,N_39796,N_39797,N_39798,N_39799,N_39800,N_39801,N_39802,N_39803,N_39804,N_39805,N_39806,N_39807,N_39808,N_39809,N_39810,N_39811,N_39812,N_39813,N_39814,N_39815,N_39816,N_39817,N_39818,N_39819,N_39820,N_39821,N_39822,N_39823,N_39824,N_39825,N_39826,N_39827,N_39828,N_39829,N_39830,N_39831,N_39832,N_39833,N_39834,N_39835,N_39836,N_39837,N_39838,N_39839,N_39840,N_39841,N_39842,N_39843,N_39844,N_39845,N_39846,N_39847,N_39848,N_39849,N_39850,N_39851,N_39852,N_39853,N_39854,N_39855,N_39856,N_39857,N_39858,N_39859,N_39860,N_39861,N_39862,N_39863,N_39864,N_39865,N_39866,N_39867,N_39868,N_39869,N_39870,N_39871,N_39872,N_39873,N_39874,N_39875,N_39876,N_39877,N_39878,N_39879,N_39880,N_39881,N_39882,N_39883,N_39884,N_39885,N_39886,N_39887,N_39888,N_39889,N_39890,N_39891,N_39892,N_39893,N_39894,N_39895,N_39896,N_39897,N_39898,N_39899,N_39900,N_39901,N_39902,N_39903,N_39904,N_39905,N_39906,N_39907,N_39908,N_39909,N_39910,N_39911,N_39912,N_39913,N_39914,N_39915,N_39916,N_39917,N_39918,N_39919,N_39920,N_39921,N_39922,N_39923,N_39924,N_39925,N_39926,N_39927,N_39928,N_39929,N_39930,N_39931,N_39932,N_39933,N_39934,N_39935,N_39936,N_39937,N_39938,N_39939,N_39940,N_39941,N_39942,N_39943,N_39944,N_39945,N_39946,N_39947,N_39948,N_39949,N_39950,N_39951,N_39952,N_39953,N_39954,N_39955,N_39956,N_39957,N_39958,N_39959,N_39960,N_39961,N_39962,N_39963,N_39964,N_39965,N_39966,N_39967,N_39968,N_39969,N_39970,N_39971,N_39972,N_39973,N_39974,N_39975,N_39976,N_39977,N_39978,N_39979,N_39980,N_39981,N_39982,N_39983,N_39984,N_39985,N_39986,N_39987,N_39988,N_39989,N_39990,N_39991,N_39992,N_39993,N_39994,N_39995,N_39996,N_39997,N_39998,N_39999,N_40000,N_40001,N_40002,N_40003,N_40004,N_40005,N_40006,N_40007,N_40008,N_40009,N_40010,N_40011,N_40012,N_40013,N_40014,N_40015,N_40016,N_40017,N_40018,N_40019,N_40020,N_40021,N_40022,N_40023,N_40024,N_40025,N_40026,N_40027,N_40028,N_40029,N_40030,N_40031,N_40032,N_40033,N_40034,N_40035,N_40036,N_40037,N_40038,N_40039,N_40040,N_40041,N_40042,N_40043,N_40044,N_40045,N_40046,N_40047,N_40048,N_40049,N_40050,N_40051,N_40052,N_40053,N_40054,N_40055,N_40056,N_40057,N_40058,N_40059,N_40060,N_40061,N_40062,N_40063,N_40064,N_40065,N_40066,N_40067,N_40068,N_40069,N_40070,N_40071,N_40072,N_40073,N_40074,N_40075,N_40076,N_40077,N_40078,N_40079,N_40080,N_40081,N_40082,N_40083,N_40084,N_40085,N_40086,N_40087,N_40088,N_40089,N_40090,N_40091,N_40092,N_40093,N_40094,N_40095,N_40096,N_40097,N_40098,N_40099,N_40100,N_40101,N_40102,N_40103,N_40104,N_40105,N_40106,N_40107,N_40108,N_40109,N_40110,N_40111,N_40112,N_40113,N_40114,N_40115,N_40116,N_40117,N_40118,N_40119,N_40120,N_40121,N_40122,N_40123,N_40124,N_40125,N_40126,N_40127,N_40128,N_40129,N_40130,N_40131,N_40132,N_40133,N_40134,N_40135,N_40136,N_40137,N_40138,N_40139,N_40140,N_40141,N_40142,N_40143,N_40144,N_40145,N_40146,N_40147,N_40148,N_40149,N_40150,N_40151,N_40152,N_40153,N_40154,N_40155,N_40156,N_40157,N_40158,N_40159,N_40160,N_40161,N_40162,N_40163,N_40164,N_40165,N_40166,N_40167,N_40168,N_40169,N_40170,N_40171,N_40172,N_40173,N_40174,N_40175,N_40176,N_40177,N_40178,N_40179,N_40180,N_40181,N_40182,N_40183,N_40184,N_40185,N_40186,N_40187,N_40188,N_40189,N_40190,N_40191,N_40192,N_40193,N_40194,N_40195,N_40196,N_40197,N_40198,N_40199,N_40200,N_40201,N_40202,N_40203,N_40204,N_40205,N_40206,N_40207,N_40208,N_40209,N_40210,N_40211,N_40212,N_40213,N_40214,N_40215,N_40216,N_40217,N_40218,N_40219,N_40220,N_40221,N_40222,N_40223,N_40224,N_40225,N_40226,N_40227,N_40228,N_40229,N_40230,N_40231,N_40232,N_40233,N_40234,N_40235,N_40236,N_40237,N_40238,N_40239,N_40240,N_40241,N_40242,N_40243,N_40244,N_40245,N_40246,N_40247,N_40248,N_40249,N_40250,N_40251,N_40252,N_40253,N_40254,N_40255,N_40256,N_40257,N_40258,N_40259,N_40260,N_40261,N_40262,N_40263,N_40264,N_40265,N_40266,N_40267,N_40268,N_40269,N_40270,N_40271,N_40272,N_40273,N_40274,N_40275,N_40276,N_40277,N_40278,N_40279,N_40280,N_40281,N_40282,N_40283,N_40284,N_40285,N_40286,N_40287,N_40288,N_40289,N_40290,N_40291,N_40292,N_40293,N_40294,N_40295,N_40296,N_40297,N_40298,N_40299,N_40300,N_40301,N_40302,N_40303,N_40304,N_40305,N_40306,N_40307,N_40308,N_40309,N_40310,N_40311,N_40312,N_40313,N_40314,N_40315,N_40316,N_40317,N_40318,N_40319,N_40320,N_40321,N_40322,N_40323,N_40324,N_40325,N_40326,N_40327,N_40328,N_40329,N_40330,N_40331,N_40332,N_40333,N_40334,N_40335,N_40336,N_40337,N_40338,N_40339,N_40340,N_40341,N_40342,N_40343,N_40344,N_40345,N_40346,N_40347,N_40348,N_40349,N_40350,N_40351,N_40352,N_40353,N_40354,N_40355,N_40356,N_40357,N_40358,N_40359,N_40360,N_40361,N_40362,N_40363,N_40364,N_40365,N_40366,N_40367,N_40368,N_40369,N_40370,N_40371,N_40372,N_40373,N_40374,N_40375,N_40376,N_40377,N_40378,N_40379,N_40380,N_40381,N_40382,N_40383,N_40384,N_40385,N_40386,N_40387,N_40388,N_40389,N_40390,N_40391,N_40392,N_40393,N_40394,N_40395,N_40396,N_40397,N_40398,N_40399,N_40400,N_40401,N_40402,N_40403,N_40404,N_40405,N_40406,N_40407,N_40408,N_40409,N_40410,N_40411,N_40412,N_40413,N_40414,N_40415,N_40416,N_40417,N_40418,N_40419,N_40420,N_40421,N_40422,N_40423,N_40424,N_40425,N_40426,N_40427,N_40428,N_40429,N_40430,N_40431,N_40432,N_40433,N_40434,N_40435,N_40436,N_40437,N_40438,N_40439,N_40440,N_40441,N_40442,N_40443,N_40444,N_40445,N_40446,N_40447,N_40448,N_40449,N_40450,N_40451,N_40452,N_40453,N_40454,N_40455,N_40456,N_40457,N_40458,N_40459,N_40460,N_40461,N_40462,N_40463,N_40464,N_40465,N_40466,N_40467,N_40468,N_40469,N_40470,N_40471,N_40472,N_40473,N_40474,N_40475,N_40476,N_40477,N_40478,N_40479,N_40480,N_40481,N_40482,N_40483,N_40484,N_40485,N_40486,N_40487,N_40488,N_40489,N_40490,N_40491,N_40492,N_40493,N_40494,N_40495,N_40496,N_40497,N_40498,N_40499,N_40500,N_40501,N_40502,N_40503,N_40504,N_40505,N_40506,N_40507,N_40508,N_40509,N_40510,N_40511,N_40512,N_40513,N_40514,N_40515,N_40516,N_40517,N_40518,N_40519,N_40520,N_40521,N_40522,N_40523,N_40524,N_40525,N_40526,N_40527,N_40528,N_40529,N_40530,N_40531,N_40532,N_40533,N_40534,N_40535,N_40536,N_40537,N_40538,N_40539,N_40540,N_40541,N_40542,N_40543,N_40544,N_40545,N_40546,N_40547,N_40548,N_40549,N_40550,N_40551,N_40552,N_40553,N_40554,N_40555,N_40556,N_40557,N_40558,N_40559,N_40560,N_40561,N_40562,N_40563,N_40564,N_40565,N_40566,N_40567,N_40568,N_40569,N_40570,N_40571,N_40572,N_40573,N_40574,N_40575,N_40576,N_40577,N_40578,N_40579,N_40580,N_40581,N_40582,N_40583,N_40584,N_40585,N_40586,N_40587,N_40588,N_40589,N_40590,N_40591,N_40592,N_40593,N_40594,N_40595,N_40596,N_40597,N_40598,N_40599,N_40600,N_40601,N_40602,N_40603,N_40604,N_40605,N_40606,N_40607,N_40608,N_40609,N_40610,N_40611,N_40612,N_40613,N_40614,N_40615,N_40616,N_40617,N_40618,N_40619,N_40620,N_40621,N_40622,N_40623,N_40624,N_40625,N_40626,N_40627,N_40628,N_40629,N_40630,N_40631,N_40632,N_40633,N_40634,N_40635,N_40636,N_40637,N_40638,N_40639,N_40640,N_40641,N_40642,N_40643,N_40644,N_40645,N_40646,N_40647,N_40648,N_40649,N_40650,N_40651,N_40652,N_40653,N_40654,N_40655,N_40656,N_40657,N_40658,N_40659,N_40660,N_40661,N_40662,N_40663,N_40664,N_40665,N_40666,N_40667,N_40668,N_40669,N_40670,N_40671,N_40672,N_40673,N_40674,N_40675,N_40676,N_40677,N_40678,N_40679,N_40680,N_40681,N_40682,N_40683,N_40684,N_40685,N_40686,N_40687,N_40688,N_40689,N_40690,N_40691,N_40692,N_40693,N_40694,N_40695,N_40696,N_40697,N_40698,N_40699,N_40700,N_40701,N_40702,N_40703,N_40704,N_40705,N_40706,N_40707,N_40708,N_40709,N_40710,N_40711,N_40712,N_40713,N_40714,N_40715,N_40716,N_40717,N_40718,N_40719,N_40720,N_40721,N_40722,N_40723,N_40724,N_40725,N_40726,N_40727,N_40728,N_40729,N_40730,N_40731,N_40732,N_40733,N_40734,N_40735,N_40736,N_40737,N_40738,N_40739,N_40740,N_40741,N_40742,N_40743,N_40744,N_40745,N_40746,N_40747,N_40748,N_40749,N_40750,N_40751,N_40752,N_40753,N_40754,N_40755,N_40756,N_40757,N_40758,N_40759,N_40760,N_40761,N_40762,N_40763,N_40764,N_40765,N_40766,N_40767,N_40768,N_40769,N_40770,N_40771,N_40772,N_40773,N_40774,N_40775,N_40776,N_40777,N_40778,N_40779,N_40780,N_40781,N_40782,N_40783,N_40784,N_40785,N_40786,N_40787,N_40788,N_40789,N_40790,N_40791,N_40792,N_40793,N_40794,N_40795,N_40796,N_40797,N_40798,N_40799,N_40800,N_40801,N_40802,N_40803,N_40804,N_40805,N_40806,N_40807,N_40808,N_40809,N_40810,N_40811,N_40812,N_40813,N_40814,N_40815,N_40816,N_40817,N_40818,N_40819,N_40820,N_40821,N_40822,N_40823,N_40824,N_40825,N_40826,N_40827,N_40828,N_40829,N_40830,N_40831,N_40832,N_40833,N_40834,N_40835,N_40836,N_40837,N_40838,N_40839,N_40840,N_40841,N_40842,N_40843,N_40844,N_40845,N_40846,N_40847,N_40848,N_40849,N_40850,N_40851,N_40852,N_40853,N_40854,N_40855,N_40856,N_40857,N_40858,N_40859,N_40860,N_40861,N_40862,N_40863,N_40864,N_40865,N_40866,N_40867,N_40868,N_40869,N_40870,N_40871,N_40872,N_40873,N_40874,N_40875,N_40876,N_40877,N_40878,N_40879,N_40880,N_40881,N_40882,N_40883,N_40884,N_40885,N_40886,N_40887,N_40888,N_40889,N_40890,N_40891,N_40892,N_40893,N_40894,N_40895,N_40896,N_40897,N_40898,N_40899,N_40900,N_40901,N_40902,N_40903,N_40904,N_40905,N_40906,N_40907,N_40908,N_40909,N_40910,N_40911,N_40912,N_40913,N_40914,N_40915,N_40916,N_40917,N_40918,N_40919,N_40920,N_40921,N_40922,N_40923,N_40924,N_40925,N_40926,N_40927,N_40928,N_40929,N_40930,N_40931,N_40932,N_40933,N_40934,N_40935,N_40936,N_40937,N_40938,N_40939,N_40940,N_40941,N_40942,N_40943,N_40944,N_40945,N_40946,N_40947,N_40948,N_40949,N_40950,N_40951,N_40952,N_40953,N_40954,N_40955,N_40956,N_40957,N_40958,N_40959,N_40960,N_40961,N_40962,N_40963,N_40964,N_40965,N_40966,N_40967,N_40968,N_40969,N_40970,N_40971,N_40972,N_40973,N_40974,N_40975,N_40976,N_40977,N_40978,N_40979,N_40980,N_40981,N_40982,N_40983,N_40984,N_40985,N_40986,N_40987,N_40988,N_40989,N_40990,N_40991,N_40992,N_40993,N_40994,N_40995,N_40996,N_40997,N_40998,N_40999,N_41000,N_41001,N_41002,N_41003,N_41004,N_41005,N_41006,N_41007,N_41008,N_41009,N_41010,N_41011,N_41012,N_41013,N_41014,N_41015,N_41016,N_41017,N_41018,N_41019,N_41020,N_41021,N_41022,N_41023,N_41024,N_41025,N_41026,N_41027,N_41028,N_41029,N_41030,N_41031,N_41032,N_41033,N_41034,N_41035,N_41036,N_41037,N_41038,N_41039,N_41040,N_41041,N_41042,N_41043,N_41044,N_41045,N_41046,N_41047,N_41048,N_41049,N_41050,N_41051,N_41052,N_41053,N_41054,N_41055,N_41056,N_41057,N_41058,N_41059,N_41060,N_41061,N_41062,N_41063,N_41064,N_41065,N_41066,N_41067,N_41068,N_41069,N_41070,N_41071,N_41072,N_41073,N_41074,N_41075,N_41076,N_41077,N_41078,N_41079,N_41080,N_41081,N_41082,N_41083,N_41084,N_41085,N_41086,N_41087,N_41088,N_41089,N_41090,N_41091,N_41092,N_41093,N_41094,N_41095,N_41096,N_41097,N_41098,N_41099,N_41100,N_41101,N_41102,N_41103,N_41104,N_41105,N_41106,N_41107,N_41108,N_41109,N_41110,N_41111,N_41112,N_41113,N_41114,N_41115,N_41116,N_41117,N_41118,N_41119,N_41120,N_41121,N_41122,N_41123,N_41124,N_41125,N_41126,N_41127,N_41128,N_41129,N_41130,N_41131,N_41132,N_41133,N_41134,N_41135,N_41136,N_41137,N_41138,N_41139,N_41140,N_41141,N_41142,N_41143,N_41144,N_41145,N_41146,N_41147,N_41148,N_41149,N_41150,N_41151,N_41152,N_41153,N_41154,N_41155,N_41156,N_41157,N_41158,N_41159,N_41160,N_41161,N_41162,N_41163,N_41164,N_41165,N_41166,N_41167,N_41168,N_41169,N_41170,N_41171,N_41172,N_41173,N_41174,N_41175,N_41176,N_41177,N_41178,N_41179,N_41180,N_41181,N_41182,N_41183,N_41184,N_41185,N_41186,N_41187,N_41188,N_41189,N_41190,N_41191,N_41192,N_41193,N_41194,N_41195,N_41196,N_41197,N_41198,N_41199,N_41200,N_41201,N_41202,N_41203,N_41204,N_41205,N_41206,N_41207,N_41208,N_41209,N_41210,N_41211,N_41212,N_41213,N_41214,N_41215,N_41216,N_41217,N_41218,N_41219,N_41220,N_41221,N_41222,N_41223,N_41224,N_41225,N_41226,N_41227,N_41228,N_41229,N_41230,N_41231,N_41232,N_41233,N_41234,N_41235,N_41236,N_41237,N_41238,N_41239,N_41240,N_41241,N_41242,N_41243,N_41244,N_41245,N_41246,N_41247,N_41248,N_41249,N_41250,N_41251,N_41252,N_41253,N_41254,N_41255,N_41256,N_41257,N_41258,N_41259,N_41260,N_41261,N_41262,N_41263,N_41264,N_41265,N_41266,N_41267,N_41268,N_41269,N_41270,N_41271,N_41272,N_41273,N_41274,N_41275,N_41276,N_41277,N_41278,N_41279,N_41280,N_41281,N_41282,N_41283,N_41284,N_41285,N_41286,N_41287,N_41288,N_41289,N_41290,N_41291,N_41292,N_41293,N_41294,N_41295,N_41296,N_41297,N_41298,N_41299,N_41300,N_41301,N_41302,N_41303,N_41304,N_41305,N_41306,N_41307,N_41308,N_41309,N_41310,N_41311,N_41312,N_41313,N_41314,N_41315,N_41316,N_41317,N_41318,N_41319,N_41320,N_41321,N_41322,N_41323,N_41324,N_41325,N_41326,N_41327,N_41328,N_41329,N_41330,N_41331,N_41332,N_41333,N_41334,N_41335,N_41336,N_41337,N_41338,N_41339,N_41340,N_41341,N_41342,N_41343,N_41344,N_41345,N_41346,N_41347,N_41348,N_41349,N_41350,N_41351,N_41352,N_41353,N_41354,N_41355,N_41356,N_41357,N_41358,N_41359,N_41360,N_41361,N_41362,N_41363,N_41364,N_41365,N_41366,N_41367,N_41368,N_41369,N_41370,N_41371,N_41372,N_41373,N_41374,N_41375,N_41376,N_41377,N_41378,N_41379,N_41380,N_41381,N_41382,N_41383,N_41384,N_41385,N_41386,N_41387,N_41388,N_41389,N_41390,N_41391,N_41392,N_41393,N_41394,N_41395,N_41396,N_41397,N_41398,N_41399,N_41400,N_41401,N_41402,N_41403,N_41404,N_41405,N_41406,N_41407,N_41408,N_41409,N_41410,N_41411,N_41412,N_41413,N_41414,N_41415,N_41416,N_41417,N_41418,N_41419,N_41420,N_41421,N_41422,N_41423,N_41424,N_41425,N_41426,N_41427,N_41428,N_41429,N_41430,N_41431,N_41432,N_41433,N_41434,N_41435,N_41436,N_41437,N_41438,N_41439,N_41440,N_41441,N_41442,N_41443,N_41444,N_41445,N_41446,N_41447,N_41448,N_41449,N_41450,N_41451,N_41452,N_41453,N_41454,N_41455,N_41456,N_41457,N_41458,N_41459,N_41460,N_41461,N_41462,N_41463,N_41464,N_41465,N_41466,N_41467,N_41468,N_41469,N_41470,N_41471,N_41472,N_41473,N_41474,N_41475,N_41476,N_41477,N_41478,N_41479,N_41480,N_41481,N_41482,N_41483,N_41484,N_41485,N_41486,N_41487,N_41488,N_41489,N_41490,N_41491,N_41492,N_41493,N_41494,N_41495,N_41496,N_41497,N_41498,N_41499,N_41500,N_41501,N_41502,N_41503,N_41504,N_41505,N_41506,N_41507,N_41508,N_41509,N_41510,N_41511,N_41512,N_41513,N_41514,N_41515,N_41516,N_41517,N_41518,N_41519,N_41520,N_41521,N_41522,N_41523,N_41524,N_41525,N_41526,N_41527,N_41528,N_41529,N_41530,N_41531,N_41532,N_41533,N_41534,N_41535,N_41536,N_41537,N_41538,N_41539,N_41540,N_41541,N_41542,N_41543,N_41544,N_41545,N_41546,N_41547,N_41548,N_41549,N_41550,N_41551,N_41552,N_41553,N_41554,N_41555,N_41556,N_41557,N_41558,N_41559,N_41560,N_41561,N_41562,N_41563,N_41564,N_41565,N_41566,N_41567,N_41568,N_41569,N_41570,N_41571,N_41572,N_41573,N_41574,N_41575,N_41576,N_41577,N_41578,N_41579,N_41580,N_41581,N_41582,N_41583,N_41584,N_41585,N_41586,N_41587,N_41588,N_41589,N_41590,N_41591,N_41592,N_41593,N_41594,N_41595,N_41596,N_41597,N_41598,N_41599,N_41600,N_41601,N_41602,N_41603,N_41604,N_41605,N_41606,N_41607,N_41608,N_41609,N_41610,N_41611,N_41612,N_41613,N_41614,N_41615,N_41616,N_41617,N_41618,N_41619,N_41620,N_41621,N_41622,N_41623,N_41624,N_41625,N_41626,N_41627,N_41628,N_41629,N_41630,N_41631,N_41632,N_41633,N_41634,N_41635,N_41636,N_41637,N_41638,N_41639,N_41640,N_41641,N_41642,N_41643,N_41644,N_41645,N_41646,N_41647,N_41648,N_41649,N_41650,N_41651,N_41652,N_41653,N_41654,N_41655,N_41656,N_41657,N_41658,N_41659,N_41660,N_41661,N_41662,N_41663,N_41664,N_41665,N_41666,N_41667,N_41668,N_41669,N_41670,N_41671,N_41672,N_41673,N_41674,N_41675,N_41676,N_41677,N_41678,N_41679,N_41680,N_41681,N_41682,N_41683,N_41684,N_41685,N_41686,N_41687,N_41688,N_41689,N_41690,N_41691,N_41692,N_41693,N_41694,N_41695,N_41696,N_41697,N_41698,N_41699,N_41700,N_41701,N_41702,N_41703,N_41704,N_41705,N_41706,N_41707,N_41708,N_41709,N_41710,N_41711,N_41712,N_41713,N_41714,N_41715,N_41716,N_41717,N_41718,N_41719,N_41720,N_41721,N_41722,N_41723,N_41724,N_41725,N_41726,N_41727,N_41728,N_41729,N_41730,N_41731,N_41732,N_41733,N_41734,N_41735,N_41736,N_41737,N_41738,N_41739,N_41740,N_41741,N_41742,N_41743,N_41744,N_41745,N_41746,N_41747,N_41748,N_41749,N_41750,N_41751,N_41752,N_41753,N_41754,N_41755,N_41756,N_41757,N_41758,N_41759,N_41760,N_41761,N_41762,N_41763,N_41764,N_41765,N_41766,N_41767,N_41768,N_41769,N_41770,N_41771,N_41772,N_41773,N_41774,N_41775,N_41776,N_41777,N_41778,N_41779,N_41780,N_41781,N_41782,N_41783,N_41784,N_41785,N_41786,N_41787,N_41788,N_41789,N_41790,N_41791,N_41792,N_41793,N_41794,N_41795,N_41796,N_41797,N_41798,N_41799,N_41800,N_41801,N_41802,N_41803,N_41804,N_41805,N_41806,N_41807,N_41808,N_41809,N_41810,N_41811,N_41812,N_41813,N_41814,N_41815,N_41816,N_41817,N_41818,N_41819,N_41820,N_41821,N_41822,N_41823,N_41824,N_41825,N_41826,N_41827,N_41828,N_41829,N_41830,N_41831,N_41832,N_41833,N_41834,N_41835,N_41836,N_41837,N_41838,N_41839,N_41840,N_41841,N_41842,N_41843,N_41844,N_41845,N_41846,N_41847,N_41848,N_41849,N_41850,N_41851,N_41852,N_41853,N_41854,N_41855,N_41856,N_41857,N_41858,N_41859,N_41860,N_41861,N_41862,N_41863,N_41864,N_41865,N_41866,N_41867,N_41868,N_41869,N_41870,N_41871,N_41872,N_41873,N_41874,N_41875,N_41876,N_41877,N_41878,N_41879,N_41880,N_41881,N_41882,N_41883,N_41884,N_41885,N_41886,N_41887,N_41888,N_41889,N_41890,N_41891,N_41892,N_41893,N_41894,N_41895,N_41896,N_41897,N_41898,N_41899,N_41900,N_41901,N_41902,N_41903,N_41904,N_41905,N_41906,N_41907,N_41908,N_41909,N_41910,N_41911,N_41912,N_41913,N_41914,N_41915,N_41916,N_41917,N_41918,N_41919,N_41920,N_41921,N_41922,N_41923,N_41924,N_41925,N_41926,N_41927,N_41928,N_41929,N_41930,N_41931,N_41932,N_41933,N_41934,N_41935,N_41936,N_41937,N_41938,N_41939,N_41940,N_41941,N_41942,N_41943,N_41944,N_41945,N_41946,N_41947,N_41948,N_41949,N_41950,N_41951,N_41952,N_41953,N_41954,N_41955,N_41956,N_41957,N_41958,N_41959,N_41960,N_41961,N_41962,N_41963,N_41964,N_41965,N_41966,N_41967,N_41968,N_41969,N_41970,N_41971,N_41972,N_41973,N_41974,N_41975,N_41976,N_41977,N_41978,N_41979,N_41980,N_41981,N_41982,N_41983,N_41984,N_41985,N_41986,N_41987,N_41988,N_41989,N_41990,N_41991,N_41992,N_41993,N_41994,N_41995,N_41996,N_41997,N_41998,N_41999,N_42000,N_42001,N_42002,N_42003,N_42004,N_42005,N_42006,N_42007,N_42008,N_42009,N_42010,N_42011,N_42012,N_42013,N_42014,N_42015,N_42016,N_42017,N_42018,N_42019,N_42020,N_42021,N_42022,N_42023,N_42024,N_42025,N_42026,N_42027,N_42028,N_42029,N_42030,N_42031,N_42032,N_42033,N_42034,N_42035,N_42036,N_42037,N_42038,N_42039,N_42040,N_42041,N_42042,N_42043,N_42044,N_42045,N_42046,N_42047,N_42048,N_42049,N_42050,N_42051,N_42052,N_42053,N_42054,N_42055,N_42056,N_42057,N_42058,N_42059,N_42060,N_42061,N_42062,N_42063,N_42064,N_42065,N_42066,N_42067,N_42068,N_42069,N_42070,N_42071,N_42072,N_42073,N_42074,N_42075,N_42076,N_42077,N_42078,N_42079,N_42080,N_42081,N_42082,N_42083,N_42084,N_42085,N_42086,N_42087,N_42088,N_42089,N_42090,N_42091,N_42092,N_42093,N_42094,N_42095,N_42096,N_42097,N_42098,N_42099,N_42100,N_42101,N_42102,N_42103,N_42104,N_42105,N_42106,N_42107,N_42108,N_42109,N_42110,N_42111,N_42112,N_42113,N_42114,N_42115,N_42116,N_42117,N_42118,N_42119,N_42120,N_42121,N_42122,N_42123,N_42124,N_42125,N_42126,N_42127,N_42128,N_42129,N_42130,N_42131,N_42132,N_42133,N_42134,N_42135,N_42136,N_42137,N_42138,N_42139,N_42140,N_42141,N_42142,N_42143,N_42144,N_42145,N_42146,N_42147,N_42148,N_42149,N_42150,N_42151,N_42152,N_42153,N_42154,N_42155,N_42156,N_42157,N_42158,N_42159,N_42160,N_42161,N_42162,N_42163,N_42164,N_42165,N_42166,N_42167,N_42168,N_42169,N_42170,N_42171,N_42172,N_42173,N_42174,N_42175,N_42176,N_42177,N_42178,N_42179,N_42180,N_42181,N_42182,N_42183,N_42184,N_42185,N_42186,N_42187,N_42188,N_42189,N_42190,N_42191,N_42192,N_42193,N_42194,N_42195,N_42196,N_42197,N_42198,N_42199,N_42200,N_42201,N_42202,N_42203,N_42204,N_42205,N_42206,N_42207,N_42208,N_42209,N_42210,N_42211,N_42212,N_42213,N_42214,N_42215,N_42216,N_42217,N_42218,N_42219,N_42220,N_42221,N_42222,N_42223,N_42224,N_42225,N_42226,N_42227,N_42228,N_42229,N_42230,N_42231,N_42232,N_42233,N_42234,N_42235,N_42236,N_42237,N_42238,N_42239,N_42240,N_42241,N_42242,N_42243,N_42244,N_42245,N_42246,N_42247,N_42248,N_42249,N_42250,N_42251,N_42252,N_42253,N_42254,N_42255,N_42256,N_42257,N_42258,N_42259,N_42260,N_42261,N_42262,N_42263,N_42264,N_42265,N_42266,N_42267,N_42268,N_42269,N_42270,N_42271,N_42272,N_42273,N_42274,N_42275,N_42276,N_42277,N_42278,N_42279,N_42280,N_42281,N_42282,N_42283,N_42284,N_42285,N_42286,N_42287,N_42288,N_42289,N_42290,N_42291,N_42292,N_42293,N_42294,N_42295,N_42296,N_42297,N_42298,N_42299,N_42300,N_42301,N_42302,N_42303,N_42304,N_42305,N_42306,N_42307,N_42308,N_42309,N_42310,N_42311,N_42312,N_42313,N_42314,N_42315,N_42316,N_42317,N_42318,N_42319,N_42320,N_42321,N_42322,N_42323,N_42324,N_42325,N_42326,N_42327,N_42328,N_42329,N_42330,N_42331,N_42332,N_42333,N_42334,N_42335,N_42336,N_42337,N_42338,N_42339,N_42340,N_42341,N_42342,N_42343,N_42344,N_42345,N_42346,N_42347,N_42348,N_42349,N_42350,N_42351,N_42352,N_42353,N_42354,N_42355,N_42356,N_42357,N_42358,N_42359,N_42360,N_42361,N_42362,N_42363,N_42364,N_42365,N_42366,N_42367,N_42368,N_42369,N_42370,N_42371,N_42372,N_42373,N_42374,N_42375,N_42376,N_42377,N_42378,N_42379,N_42380,N_42381,N_42382,N_42383,N_42384,N_42385,N_42386,N_42387,N_42388,N_42389,N_42390,N_42391,N_42392,N_42393,N_42394,N_42395,N_42396,N_42397,N_42398,N_42399,N_42400,N_42401,N_42402,N_42403,N_42404,N_42405,N_42406,N_42407,N_42408,N_42409,N_42410,N_42411,N_42412,N_42413,N_42414,N_42415,N_42416,N_42417,N_42418,N_42419,N_42420,N_42421,N_42422,N_42423,N_42424,N_42425,N_42426,N_42427,N_42428,N_42429,N_42430,N_42431,N_42432,N_42433,N_42434,N_42435,N_42436,N_42437,N_42438,N_42439,N_42440,N_42441,N_42442,N_42443,N_42444,N_42445,N_42446,N_42447,N_42448,N_42449,N_42450,N_42451,N_42452,N_42453,N_42454,N_42455,N_42456,N_42457,N_42458,N_42459,N_42460,N_42461,N_42462,N_42463,N_42464,N_42465,N_42466,N_42467,N_42468,N_42469,N_42470,N_42471,N_42472,N_42473,N_42474,N_42475,N_42476,N_42477,N_42478,N_42479,N_42480,N_42481,N_42482,N_42483,N_42484,N_42485,N_42486,N_42487,N_42488,N_42489,N_42490,N_42491,N_42492,N_42493,N_42494,N_42495,N_42496,N_42497,N_42498,N_42499,N_42500,N_42501,N_42502,N_42503,N_42504,N_42505,N_42506,N_42507,N_42508,N_42509,N_42510,N_42511,N_42512,N_42513,N_42514,N_42515,N_42516,N_42517,N_42518,N_42519,N_42520,N_42521,N_42522,N_42523,N_42524,N_42525,N_42526,N_42527,N_42528,N_42529,N_42530,N_42531,N_42532,N_42533,N_42534,N_42535,N_42536,N_42537,N_42538,N_42539,N_42540,N_42541,N_42542,N_42543,N_42544,N_42545,N_42546,N_42547,N_42548,N_42549,N_42550,N_42551,N_42552,N_42553,N_42554,N_42555,N_42556,N_42557,N_42558,N_42559,N_42560,N_42561,N_42562,N_42563,N_42564,N_42565,N_42566,N_42567,N_42568,N_42569,N_42570,N_42571,N_42572,N_42573,N_42574,N_42575,N_42576,N_42577,N_42578,N_42579,N_42580,N_42581,N_42582,N_42583,N_42584,N_42585,N_42586,N_42587,N_42588,N_42589,N_42590,N_42591,N_42592,N_42593,N_42594,N_42595,N_42596,N_42597,N_42598,N_42599,N_42600,N_42601,N_42602,N_42603,N_42604,N_42605,N_42606,N_42607,N_42608,N_42609,N_42610,N_42611,N_42612,N_42613,N_42614,N_42615,N_42616,N_42617,N_42618,N_42619,N_42620,N_42621,N_42622,N_42623,N_42624,N_42625,N_42626,N_42627,N_42628,N_42629,N_42630,N_42631,N_42632,N_42633,N_42634,N_42635,N_42636,N_42637,N_42638,N_42639,N_42640,N_42641,N_42642,N_42643,N_42644,N_42645,N_42646,N_42647,N_42648,N_42649,N_42650,N_42651,N_42652,N_42653,N_42654,N_42655,N_42656,N_42657,N_42658,N_42659,N_42660,N_42661,N_42662,N_42663,N_42664,N_42665,N_42666,N_42667,N_42668,N_42669,N_42670,N_42671,N_42672,N_42673,N_42674,N_42675,N_42676,N_42677,N_42678,N_42679,N_42680,N_42681,N_42682,N_42683,N_42684,N_42685,N_42686,N_42687,N_42688,N_42689,N_42690,N_42691,N_42692,N_42693,N_42694,N_42695,N_42696,N_42697,N_42698,N_42699,N_42700,N_42701,N_42702,N_42703,N_42704,N_42705,N_42706,N_42707,N_42708,N_42709,N_42710,N_42711,N_42712,N_42713,N_42714,N_42715,N_42716,N_42717,N_42718,N_42719,N_42720,N_42721,N_42722,N_42723,N_42724,N_42725,N_42726,N_42727,N_42728,N_42729,N_42730,N_42731,N_42732,N_42733,N_42734,N_42735,N_42736,N_42737,N_42738,N_42739,N_42740,N_42741,N_42742,N_42743,N_42744,N_42745,N_42746,N_42747,N_42748,N_42749,N_42750,N_42751,N_42752,N_42753,N_42754,N_42755,N_42756,N_42757,N_42758,N_42759,N_42760,N_42761,N_42762,N_42763,N_42764,N_42765,N_42766,N_42767,N_42768,N_42769,N_42770,N_42771,N_42772,N_42773,N_42774,N_42775,N_42776,N_42777,N_42778,N_42779,N_42780,N_42781,N_42782,N_42783,N_42784,N_42785,N_42786,N_42787,N_42788,N_42789,N_42790,N_42791,N_42792,N_42793,N_42794,N_42795,N_42796,N_42797,N_42798,N_42799,N_42800,N_42801,N_42802,N_42803,N_42804,N_42805,N_42806,N_42807,N_42808,N_42809,N_42810,N_42811,N_42812,N_42813,N_42814,N_42815,N_42816,N_42817,N_42818,N_42819,N_42820,N_42821,N_42822,N_42823,N_42824,N_42825,N_42826,N_42827,N_42828,N_42829,N_42830,N_42831,N_42832,N_42833,N_42834,N_42835,N_42836,N_42837,N_42838,N_42839,N_42840,N_42841,N_42842,N_42843,N_42844,N_42845,N_42846,N_42847,N_42848,N_42849,N_42850,N_42851,N_42852,N_42853,N_42854,N_42855,N_42856,N_42857,N_42858,N_42859,N_42860,N_42861,N_42862,N_42863,N_42864,N_42865,N_42866,N_42867,N_42868,N_42869,N_42870,N_42871,N_42872,N_42873,N_42874,N_42875,N_42876,N_42877,N_42878,N_42879,N_42880,N_42881,N_42882,N_42883,N_42884,N_42885,N_42886,N_42887,N_42888,N_42889,N_42890,N_42891,N_42892,N_42893,N_42894,N_42895,N_42896,N_42897,N_42898,N_42899,N_42900,N_42901,N_42902,N_42903,N_42904,N_42905,N_42906,N_42907,N_42908,N_42909,N_42910,N_42911,N_42912,N_42913,N_42914,N_42915,N_42916,N_42917,N_42918,N_42919,N_42920,N_42921,N_42922,N_42923,N_42924,N_42925,N_42926,N_42927,N_42928,N_42929,N_42930,N_42931,N_42932,N_42933,N_42934,N_42935,N_42936,N_42937,N_42938,N_42939,N_42940,N_42941,N_42942,N_42943,N_42944,N_42945,N_42946,N_42947,N_42948,N_42949,N_42950,N_42951,N_42952,N_42953,N_42954,N_42955,N_42956,N_42957,N_42958,N_42959,N_42960,N_42961,N_42962,N_42963,N_42964,N_42965,N_42966,N_42967,N_42968,N_42969,N_42970,N_42971,N_42972,N_42973,N_42974,N_42975,N_42976,N_42977,N_42978,N_42979,N_42980,N_42981,N_42982,N_42983,N_42984,N_42985,N_42986,N_42987,N_42988,N_42989,N_42990,N_42991,N_42992,N_42993,N_42994,N_42995,N_42996,N_42997,N_42998,N_42999,N_43000,N_43001,N_43002,N_43003,N_43004,N_43005,N_43006,N_43007,N_43008,N_43009,N_43010,N_43011,N_43012,N_43013,N_43014,N_43015,N_43016,N_43017,N_43018,N_43019,N_43020,N_43021,N_43022,N_43023,N_43024,N_43025,N_43026,N_43027,N_43028,N_43029,N_43030,N_43031,N_43032,N_43033,N_43034,N_43035,N_43036,N_43037,N_43038,N_43039,N_43040,N_43041,N_43042,N_43043,N_43044,N_43045,N_43046,N_43047,N_43048,N_43049,N_43050,N_43051,N_43052,N_43053,N_43054,N_43055,N_43056,N_43057,N_43058,N_43059,N_43060,N_43061,N_43062,N_43063,N_43064,N_43065,N_43066,N_43067,N_43068,N_43069,N_43070,N_43071,N_43072,N_43073,N_43074,N_43075,N_43076,N_43077,N_43078,N_43079,N_43080,N_43081,N_43082,N_43083,N_43084,N_43085,N_43086,N_43087,N_43088,N_43089,N_43090,N_43091,N_43092,N_43093,N_43094,N_43095,N_43096,N_43097,N_43098,N_43099,N_43100,N_43101,N_43102,N_43103,N_43104,N_43105,N_43106,N_43107,N_43108,N_43109,N_43110,N_43111,N_43112,N_43113,N_43114,N_43115,N_43116,N_43117,N_43118,N_43119,N_43120,N_43121,N_43122,N_43123,N_43124,N_43125,N_43126,N_43127,N_43128,N_43129,N_43130,N_43131,N_43132,N_43133,N_43134,N_43135,N_43136,N_43137,N_43138,N_43139,N_43140,N_43141,N_43142,N_43143,N_43144,N_43145,N_43146,N_43147,N_43148,N_43149,N_43150,N_43151,N_43152,N_43153,N_43154,N_43155,N_43156,N_43157,N_43158,N_43159,N_43160,N_43161,N_43162,N_43163,N_43164,N_43165,N_43166,N_43167,N_43168,N_43169,N_43170,N_43171,N_43172,N_43173,N_43174,N_43175,N_43176,N_43177,N_43178,N_43179,N_43180,N_43181,N_43182,N_43183,N_43184,N_43185,N_43186,N_43187,N_43188,N_43189,N_43190,N_43191,N_43192,N_43193,N_43194,N_43195,N_43196,N_43197,N_43198,N_43199,N_43200,N_43201,N_43202,N_43203,N_43204,N_43205,N_43206,N_43207,N_43208,N_43209,N_43210,N_43211,N_43212,N_43213,N_43214,N_43215,N_43216,N_43217,N_43218,N_43219,N_43220,N_43221,N_43222,N_43223,N_43224,N_43225,N_43226,N_43227,N_43228,N_43229,N_43230,N_43231,N_43232,N_43233,N_43234,N_43235,N_43236,N_43237,N_43238,N_43239,N_43240,N_43241,N_43242,N_43243,N_43244,N_43245,N_43246,N_43247,N_43248,N_43249,N_43250,N_43251,N_43252,N_43253,N_43254,N_43255,N_43256,N_43257,N_43258,N_43259,N_43260,N_43261,N_43262,N_43263,N_43264,N_43265,N_43266,N_43267,N_43268,N_43269,N_43270,N_43271,N_43272,N_43273,N_43274,N_43275,N_43276,N_43277,N_43278,N_43279,N_43280,N_43281,N_43282,N_43283,N_43284,N_43285,N_43286,N_43287,N_43288,N_43289,N_43290,N_43291,N_43292,N_43293,N_43294,N_43295,N_43296,N_43297,N_43298,N_43299,N_43300,N_43301,N_43302,N_43303,N_43304,N_43305,N_43306,N_43307,N_43308,N_43309,N_43310,N_43311,N_43312,N_43313,N_43314,N_43315,N_43316,N_43317,N_43318,N_43319,N_43320,N_43321,N_43322,N_43323,N_43324,N_43325,N_43326,N_43327,N_43328,N_43329,N_43330,N_43331,N_43332,N_43333,N_43334,N_43335,N_43336,N_43337,N_43338,N_43339,N_43340,N_43341,N_43342,N_43343,N_43344,N_43345,N_43346,N_43347,N_43348,N_43349,N_43350,N_43351,N_43352,N_43353,N_43354,N_43355,N_43356,N_43357,N_43358,N_43359,N_43360,N_43361,N_43362,N_43363,N_43364,N_43365,N_43366,N_43367,N_43368,N_43369,N_43370,N_43371,N_43372,N_43373,N_43374,N_43375,N_43376,N_43377,N_43378,N_43379,N_43380,N_43381,N_43382,N_43383,N_43384,N_43385,N_43386,N_43387,N_43388,N_43389,N_43390,N_43391,N_43392,N_43393,N_43394,N_43395,N_43396,N_43397,N_43398,N_43399,N_43400,N_43401,N_43402,N_43403,N_43404,N_43405,N_43406,N_43407,N_43408,N_43409,N_43410,N_43411,N_43412,N_43413,N_43414,N_43415,N_43416,N_43417,N_43418,N_43419,N_43420,N_43421,N_43422,N_43423,N_43424,N_43425,N_43426,N_43427,N_43428,N_43429,N_43430,N_43431,N_43432,N_43433,N_43434,N_43435,N_43436,N_43437,N_43438,N_43439,N_43440,N_43441,N_43442,N_43443,N_43444,N_43445,N_43446,N_43447,N_43448,N_43449,N_43450,N_43451,N_43452,N_43453,N_43454,N_43455,N_43456,N_43457,N_43458,N_43459,N_43460,N_43461,N_43462,N_43463,N_43464,N_43465,N_43466,N_43467,N_43468,N_43469,N_43470,N_43471,N_43472,N_43473,N_43474,N_43475,N_43476,N_43477,N_43478,N_43479,N_43480,N_43481,N_43482,N_43483,N_43484,N_43485,N_43486,N_43487,N_43488,N_43489,N_43490,N_43491,N_43492,N_43493,N_43494,N_43495,N_43496,N_43497,N_43498,N_43499,N_43500,N_43501,N_43502,N_43503,N_43504,N_43505,N_43506,N_43507,N_43508,N_43509,N_43510,N_43511,N_43512,N_43513,N_43514,N_43515,N_43516,N_43517,N_43518,N_43519,N_43520,N_43521,N_43522,N_43523,N_43524,N_43525,N_43526,N_43527,N_43528,N_43529,N_43530,N_43531,N_43532,N_43533,N_43534,N_43535,N_43536,N_43537,N_43538,N_43539,N_43540,N_43541,N_43542,N_43543,N_43544,N_43545,N_43546,N_43547,N_43548,N_43549,N_43550,N_43551,N_43552,N_43553,N_43554,N_43555,N_43556,N_43557,N_43558,N_43559,N_43560,N_43561,N_43562,N_43563,N_43564,N_43565,N_43566,N_43567,N_43568,N_43569,N_43570,N_43571,N_43572,N_43573,N_43574,N_43575,N_43576,N_43577,N_43578,N_43579,N_43580,N_43581,N_43582,N_43583,N_43584,N_43585,N_43586,N_43587,N_43588,N_43589,N_43590,N_43591,N_43592,N_43593,N_43594,N_43595,N_43596,N_43597,N_43598,N_43599,N_43600,N_43601,N_43602,N_43603,N_43604,N_43605,N_43606,N_43607,N_43608,N_43609,N_43610,N_43611,N_43612,N_43613,N_43614,N_43615,N_43616,N_43617,N_43618,N_43619,N_43620,N_43621,N_43622,N_43623,N_43624,N_43625,N_43626,N_43627,N_43628,N_43629,N_43630,N_43631,N_43632,N_43633,N_43634,N_43635,N_43636,N_43637,N_43638,N_43639,N_43640,N_43641,N_43642,N_43643,N_43644,N_43645,N_43646,N_43647,N_43648,N_43649,N_43650,N_43651,N_43652,N_43653,N_43654,N_43655,N_43656,N_43657,N_43658,N_43659,N_43660,N_43661,N_43662,N_43663,N_43664,N_43665,N_43666,N_43667,N_43668,N_43669,N_43670,N_43671,N_43672,N_43673,N_43674,N_43675,N_43676,N_43677,N_43678,N_43679,N_43680,N_43681,N_43682,N_43683,N_43684,N_43685,N_43686,N_43687,N_43688,N_43689,N_43690,N_43691,N_43692,N_43693,N_43694,N_43695,N_43696,N_43697,N_43698,N_43699,N_43700,N_43701,N_43702,N_43703,N_43704,N_43705,N_43706,N_43707,N_43708,N_43709,N_43710,N_43711,N_43712,N_43713,N_43714,N_43715,N_43716,N_43717,N_43718,N_43719,N_43720,N_43721,N_43722,N_43723,N_43724,N_43725,N_43726,N_43727,N_43728,N_43729,N_43730,N_43731,N_43732,N_43733,N_43734,N_43735,N_43736,N_43737,N_43738,N_43739,N_43740,N_43741,N_43742,N_43743,N_43744,N_43745,N_43746,N_43747,N_43748,N_43749,N_43750,N_43751,N_43752,N_43753,N_43754,N_43755,N_43756,N_43757,N_43758,N_43759,N_43760,N_43761,N_43762,N_43763,N_43764,N_43765,N_43766,N_43767,N_43768,N_43769,N_43770,N_43771,N_43772,N_43773,N_43774,N_43775,N_43776,N_43777,N_43778,N_43779,N_43780,N_43781,N_43782,N_43783,N_43784,N_43785,N_43786,N_43787,N_43788,N_43789,N_43790,N_43791,N_43792,N_43793,N_43794,N_43795,N_43796,N_43797,N_43798,N_43799,N_43800,N_43801,N_43802,N_43803,N_43804,N_43805,N_43806,N_43807,N_43808,N_43809,N_43810,N_43811,N_43812,N_43813,N_43814,N_43815,N_43816,N_43817,N_43818,N_43819,N_43820,N_43821,N_43822,N_43823,N_43824,N_43825,N_43826,N_43827,N_43828,N_43829,N_43830,N_43831,N_43832,N_43833,N_43834,N_43835,N_43836,N_43837,N_43838,N_43839,N_43840,N_43841,N_43842,N_43843,N_43844,N_43845,N_43846,N_43847,N_43848,N_43849,N_43850,N_43851,N_43852,N_43853,N_43854,N_43855,N_43856,N_43857,N_43858,N_43859,N_43860,N_43861,N_43862,N_43863,N_43864,N_43865,N_43866,N_43867,N_43868,N_43869,N_43870,N_43871,N_43872,N_43873,N_43874,N_43875,N_43876,N_43877,N_43878,N_43879,N_43880,N_43881,N_43882,N_43883,N_43884,N_43885,N_43886,N_43887,N_43888,N_43889,N_43890,N_43891,N_43892,N_43893,N_43894,N_43895,N_43896,N_43897,N_43898,N_43899,N_43900,N_43901,N_43902,N_43903,N_43904,N_43905,N_43906,N_43907,N_43908,N_43909,N_43910,N_43911,N_43912,N_43913,N_43914,N_43915,N_43916,N_43917,N_43918,N_43919,N_43920,N_43921,N_43922,N_43923,N_43924,N_43925,N_43926,N_43927,N_43928,N_43929,N_43930,N_43931,N_43932,N_43933,N_43934,N_43935,N_43936,N_43937,N_43938,N_43939,N_43940,N_43941,N_43942,N_43943,N_43944,N_43945,N_43946,N_43947,N_43948,N_43949,N_43950,N_43951,N_43952,N_43953,N_43954,N_43955,N_43956,N_43957,N_43958,N_43959,N_43960,N_43961,N_43962,N_43963,N_43964,N_43965,N_43966,N_43967,N_43968,N_43969,N_43970,N_43971,N_43972,N_43973,N_43974,N_43975,N_43976,N_43977,N_43978,N_43979,N_43980,N_43981,N_43982,N_43983,N_43984,N_43985,N_43986,N_43987,N_43988,N_43989,N_43990,N_43991,N_43992,N_43993,N_43994,N_43995,N_43996,N_43997,N_43998,N_43999,N_44000,N_44001,N_44002,N_44003,N_44004,N_44005,N_44006,N_44007,N_44008,N_44009,N_44010,N_44011,N_44012,N_44013,N_44014,N_44015,N_44016,N_44017,N_44018,N_44019,N_44020,N_44021,N_44022,N_44023,N_44024,N_44025,N_44026,N_44027,N_44028,N_44029,N_44030,N_44031,N_44032,N_44033,N_44034,N_44035,N_44036,N_44037,N_44038,N_44039,N_44040,N_44041,N_44042,N_44043,N_44044,N_44045,N_44046,N_44047,N_44048,N_44049,N_44050,N_44051,N_44052,N_44053,N_44054,N_44055,N_44056,N_44057,N_44058,N_44059,N_44060,N_44061,N_44062,N_44063,N_44064,N_44065,N_44066,N_44067,N_44068,N_44069,N_44070,N_44071,N_44072,N_44073,N_44074,N_44075,N_44076,N_44077,N_44078,N_44079,N_44080,N_44081,N_44082,N_44083,N_44084,N_44085,N_44086,N_44087,N_44088,N_44089,N_44090,N_44091,N_44092,N_44093,N_44094,N_44095,N_44096,N_44097,N_44098,N_44099,N_44100,N_44101,N_44102,N_44103,N_44104,N_44105,N_44106,N_44107,N_44108,N_44109,N_44110,N_44111,N_44112,N_44113,N_44114,N_44115,N_44116,N_44117,N_44118,N_44119,N_44120,N_44121,N_44122,N_44123,N_44124,N_44125,N_44126,N_44127,N_44128,N_44129,N_44130,N_44131,N_44132,N_44133,N_44134,N_44135,N_44136,N_44137,N_44138,N_44139,N_44140,N_44141,N_44142,N_44143,N_44144,N_44145,N_44146,N_44147,N_44148,N_44149,N_44150,N_44151,N_44152,N_44153,N_44154,N_44155,N_44156,N_44157,N_44158,N_44159,N_44160,N_44161,N_44162,N_44163,N_44164,N_44165,N_44166,N_44167,N_44168,N_44169,N_44170,N_44171,N_44172,N_44173,N_44174,N_44175,N_44176,N_44177,N_44178,N_44179,N_44180,N_44181,N_44182,N_44183,N_44184,N_44185,N_44186,N_44187,N_44188,N_44189,N_44190,N_44191,N_44192,N_44193,N_44194,N_44195,N_44196,N_44197,N_44198,N_44199,N_44200,N_44201,N_44202,N_44203,N_44204,N_44205,N_44206,N_44207,N_44208,N_44209,N_44210,N_44211,N_44212,N_44213,N_44214,N_44215,N_44216,N_44217,N_44218,N_44219,N_44220,N_44221,N_44222,N_44223,N_44224,N_44225,N_44226,N_44227,N_44228,N_44229,N_44230,N_44231,N_44232,N_44233,N_44234,N_44235,N_44236,N_44237,N_44238,N_44239,N_44240,N_44241,N_44242,N_44243,N_44244,N_44245,N_44246,N_44247,N_44248,N_44249,N_44250,N_44251,N_44252,N_44253,N_44254,N_44255,N_44256,N_44257,N_44258,N_44259,N_44260,N_44261,N_44262,N_44263,N_44264,N_44265,N_44266,N_44267,N_44268,N_44269,N_44270,N_44271,N_44272,N_44273,N_44274,N_44275,N_44276,N_44277,N_44278,N_44279,N_44280,N_44281,N_44282,N_44283,N_44284,N_44285,N_44286,N_44287,N_44288,N_44289,N_44290,N_44291,N_44292,N_44293,N_44294,N_44295,N_44296,N_44297,N_44298,N_44299,N_44300,N_44301,N_44302,N_44303,N_44304,N_44305,N_44306,N_44307,N_44308,N_44309,N_44310,N_44311,N_44312,N_44313,N_44314,N_44315,N_44316,N_44317,N_44318,N_44319,N_44320,N_44321,N_44322,N_44323,N_44324,N_44325,N_44326,N_44327,N_44328,N_44329,N_44330,N_44331,N_44332,N_44333,N_44334,N_44335,N_44336,N_44337,N_44338,N_44339,N_44340,N_44341,N_44342,N_44343,N_44344,N_44345,N_44346,N_44347,N_44348,N_44349,N_44350,N_44351,N_44352,N_44353,N_44354,N_44355,N_44356,N_44357,N_44358,N_44359,N_44360,N_44361,N_44362,N_44363,N_44364,N_44365,N_44366,N_44367,N_44368,N_44369,N_44370,N_44371,N_44372,N_44373,N_44374,N_44375,N_44376,N_44377,N_44378,N_44379,N_44380,N_44381,N_44382,N_44383,N_44384,N_44385,N_44386,N_44387,N_44388,N_44389,N_44390,N_44391,N_44392,N_44393,N_44394,N_44395,N_44396,N_44397,N_44398,N_44399,N_44400,N_44401,N_44402,N_44403,N_44404,N_44405,N_44406,N_44407,N_44408,N_44409,N_44410,N_44411,N_44412,N_44413,N_44414,N_44415,N_44416,N_44417,N_44418,N_44419,N_44420,N_44421,N_44422,N_44423,N_44424,N_44425,N_44426,N_44427,N_44428,N_44429,N_44430,N_44431,N_44432,N_44433,N_44434,N_44435,N_44436,N_44437,N_44438,N_44439,N_44440,N_44441,N_44442,N_44443,N_44444,N_44445,N_44446,N_44447,N_44448,N_44449,N_44450,N_44451,N_44452,N_44453,N_44454,N_44455,N_44456,N_44457,N_44458,N_44459,N_44460,N_44461,N_44462,N_44463,N_44464,N_44465,N_44466,N_44467,N_44468,N_44469,N_44470,N_44471,N_44472,N_44473,N_44474,N_44475,N_44476,N_44477,N_44478,N_44479,N_44480,N_44481,N_44482,N_44483,N_44484,N_44485,N_44486,N_44487,N_44488,N_44489,N_44490,N_44491,N_44492,N_44493,N_44494,N_44495,N_44496,N_44497,N_44498,N_44499,N_44500,N_44501,N_44502,N_44503,N_44504,N_44505,N_44506,N_44507,N_44508,N_44509,N_44510,N_44511,N_44512,N_44513,N_44514,N_44515,N_44516,N_44517,N_44518,N_44519,N_44520,N_44521,N_44522,N_44523,N_44524,N_44525,N_44526,N_44527,N_44528,N_44529,N_44530,N_44531,N_44532,N_44533,N_44534,N_44535,N_44536,N_44537,N_44538,N_44539,N_44540,N_44541,N_44542,N_44543,N_44544,N_44545,N_44546,N_44547,N_44548,N_44549,N_44550,N_44551,N_44552,N_44553,N_44554,N_44555,N_44556,N_44557,N_44558,N_44559,N_44560,N_44561,N_44562,N_44563,N_44564,N_44565,N_44566,N_44567,N_44568,N_44569,N_44570,N_44571,N_44572,N_44573,N_44574,N_44575,N_44576,N_44577,N_44578,N_44579,N_44580,N_44581,N_44582,N_44583,N_44584,N_44585,N_44586,N_44587,N_44588,N_44589,N_44590,N_44591,N_44592,N_44593,N_44594,N_44595,N_44596,N_44597,N_44598,N_44599,N_44600,N_44601,N_44602,N_44603,N_44604,N_44605,N_44606,N_44607,N_44608,N_44609,N_44610,N_44611,N_44612,N_44613,N_44614,N_44615,N_44616,N_44617,N_44618,N_44619,N_44620,N_44621,N_44622,N_44623,N_44624,N_44625,N_44626,N_44627,N_44628,N_44629,N_44630,N_44631,N_44632,N_44633,N_44634,N_44635,N_44636,N_44637,N_44638,N_44639,N_44640,N_44641,N_44642,N_44643,N_44644,N_44645,N_44646,N_44647,N_44648,N_44649,N_44650,N_44651,N_44652,N_44653,N_44654,N_44655,N_44656,N_44657,N_44658,N_44659,N_44660,N_44661,N_44662,N_44663,N_44664,N_44665,N_44666,N_44667,N_44668,N_44669,N_44670,N_44671,N_44672,N_44673,N_44674,N_44675,N_44676,N_44677,N_44678,N_44679,N_44680,N_44681,N_44682,N_44683,N_44684,N_44685,N_44686,N_44687,N_44688,N_44689,N_44690,N_44691,N_44692,N_44693,N_44694,N_44695,N_44696,N_44697,N_44698,N_44699,N_44700,N_44701,N_44702,N_44703,N_44704,N_44705,N_44706,N_44707,N_44708,N_44709,N_44710,N_44711,N_44712,N_44713,N_44714,N_44715,N_44716,N_44717,N_44718,N_44719,N_44720,N_44721,N_44722,N_44723,N_44724,N_44725,N_44726,N_44727,N_44728,N_44729,N_44730,N_44731,N_44732,N_44733,N_44734,N_44735,N_44736,N_44737,N_44738,N_44739,N_44740,N_44741,N_44742,N_44743,N_44744,N_44745,N_44746,N_44747,N_44748,N_44749,N_44750,N_44751,N_44752,N_44753,N_44754,N_44755,N_44756,N_44757,N_44758,N_44759,N_44760,N_44761,N_44762,N_44763,N_44764,N_44765,N_44766,N_44767,N_44768,N_44769,N_44770,N_44771,N_44772,N_44773,N_44774,N_44775,N_44776,N_44777,N_44778,N_44779,N_44780,N_44781,N_44782,N_44783,N_44784,N_44785,N_44786,N_44787,N_44788,N_44789,N_44790,N_44791,N_44792,N_44793,N_44794,N_44795,N_44796,N_44797,N_44798,N_44799,N_44800,N_44801,N_44802,N_44803,N_44804,N_44805,N_44806,N_44807,N_44808,N_44809,N_44810,N_44811,N_44812,N_44813,N_44814,N_44815,N_44816,N_44817,N_44818,N_44819,N_44820,N_44821,N_44822,N_44823,N_44824,N_44825,N_44826,N_44827,N_44828,N_44829,N_44830,N_44831,N_44832,N_44833,N_44834,N_44835,N_44836,N_44837,N_44838,N_44839,N_44840,N_44841,N_44842,N_44843,N_44844,N_44845,N_44846,N_44847,N_44848,N_44849,N_44850,N_44851,N_44852,N_44853,N_44854,N_44855,N_44856,N_44857,N_44858,N_44859,N_44860,N_44861,N_44862,N_44863,N_44864,N_44865,N_44866,N_44867,N_44868,N_44869,N_44870,N_44871,N_44872,N_44873,N_44874,N_44875,N_44876,N_44877,N_44878,N_44879,N_44880,N_44881,N_44882,N_44883,N_44884,N_44885,N_44886,N_44887,N_44888,N_44889,N_44890,N_44891,N_44892,N_44893,N_44894,N_44895,N_44896,N_44897,N_44898,N_44899,N_44900,N_44901,N_44902,N_44903,N_44904,N_44905,N_44906,N_44907,N_44908,N_44909,N_44910,N_44911,N_44912,N_44913,N_44914,N_44915,N_44916,N_44917,N_44918,N_44919,N_44920,N_44921,N_44922,N_44923,N_44924,N_44925,N_44926,N_44927,N_44928,N_44929,N_44930,N_44931,N_44932,N_44933,N_44934,N_44935,N_44936,N_44937,N_44938,N_44939,N_44940,N_44941,N_44942,N_44943,N_44944,N_44945,N_44946,N_44947,N_44948,N_44949,N_44950,N_44951,N_44952,N_44953,N_44954,N_44955,N_44956,N_44957,N_44958,N_44959,N_44960,N_44961,N_44962,N_44963,N_44964,N_44965,N_44966,N_44967,N_44968,N_44969,N_44970,N_44971,N_44972,N_44973,N_44974,N_44975,N_44976,N_44977,N_44978,N_44979,N_44980,N_44981,N_44982,N_44983,N_44984,N_44985,N_44986,N_44987,N_44988,N_44989,N_44990,N_44991,N_44992,N_44993,N_44994,N_44995,N_44996,N_44997,N_44998,N_44999,N_45000,N_45001,N_45002,N_45003,N_45004,N_45005,N_45006,N_45007,N_45008,N_45009,N_45010,N_45011,N_45012,N_45013,N_45014,N_45015,N_45016,N_45017,N_45018,N_45019,N_45020,N_45021,N_45022,N_45023,N_45024,N_45025,N_45026,N_45027,N_45028,N_45029,N_45030,N_45031,N_45032,N_45033,N_45034,N_45035,N_45036,N_45037,N_45038,N_45039,N_45040,N_45041,N_45042,N_45043,N_45044,N_45045,N_45046,N_45047,N_45048,N_45049,N_45050,N_45051,N_45052,N_45053,N_45054,N_45055,N_45056,N_45057,N_45058,N_45059,N_45060,N_45061,N_45062,N_45063,N_45064,N_45065,N_45066,N_45067,N_45068,N_45069,N_45070,N_45071,N_45072,N_45073,N_45074,N_45075,N_45076,N_45077,N_45078,N_45079,N_45080,N_45081,N_45082,N_45083,N_45084,N_45085,N_45086,N_45087,N_45088,N_45089,N_45090,N_45091,N_45092,N_45093,N_45094,N_45095,N_45096,N_45097,N_45098,N_45099,N_45100,N_45101,N_45102,N_45103,N_45104,N_45105,N_45106,N_45107,N_45108,N_45109,N_45110,N_45111,N_45112,N_45113,N_45114,N_45115,N_45116,N_45117,N_45118,N_45119,N_45120,N_45121,N_45122,N_45123,N_45124,N_45125,N_45126,N_45127,N_45128,N_45129,N_45130,N_45131,N_45132,N_45133,N_45134,N_45135,N_45136,N_45137,N_45138,N_45139,N_45140,N_45141,N_45142,N_45143,N_45144,N_45145,N_45146,N_45147,N_45148,N_45149,N_45150,N_45151,N_45152,N_45153,N_45154,N_45155,N_45156,N_45157,N_45158,N_45159,N_45160,N_45161,N_45162,N_45163,N_45164,N_45165,N_45166,N_45167,N_45168,N_45169,N_45170,N_45171,N_45172,N_45173,N_45174,N_45175,N_45176,N_45177,N_45178,N_45179,N_45180,N_45181,N_45182,N_45183,N_45184,N_45185,N_45186,N_45187,N_45188,N_45189,N_45190,N_45191,N_45192,N_45193,N_45194,N_45195,N_45196,N_45197,N_45198,N_45199,N_45200,N_45201,N_45202,N_45203,N_45204,N_45205,N_45206,N_45207,N_45208,N_45209,N_45210,N_45211,N_45212,N_45213,N_45214,N_45215,N_45216,N_45217,N_45218,N_45219,N_45220,N_45221,N_45222,N_45223,N_45224,N_45225,N_45226,N_45227,N_45228,N_45229,N_45230,N_45231,N_45232,N_45233,N_45234,N_45235,N_45236,N_45237,N_45238,N_45239,N_45240,N_45241,N_45242,N_45243,N_45244,N_45245,N_45246,N_45247,N_45248,N_45249,N_45250,N_45251,N_45252,N_45253,N_45254,N_45255,N_45256,N_45257,N_45258,N_45259,N_45260,N_45261,N_45262,N_45263,N_45264,N_45265,N_45266,N_45267,N_45268,N_45269,N_45270,N_45271,N_45272,N_45273,N_45274,N_45275,N_45276,N_45277,N_45278,N_45279,N_45280,N_45281,N_45282,N_45283,N_45284,N_45285,N_45286,N_45287,N_45288,N_45289,N_45290,N_45291,N_45292,N_45293,N_45294,N_45295,N_45296,N_45297,N_45298,N_45299,N_45300,N_45301,N_45302,N_45303,N_45304,N_45305,N_45306,N_45307,N_45308,N_45309,N_45310,N_45311,N_45312,N_45313,N_45314,N_45315,N_45316,N_45317,N_45318,N_45319,N_45320,N_45321,N_45322,N_45323,N_45324,N_45325,N_45326,N_45327,N_45328,N_45329,N_45330,N_45331,N_45332,N_45333,N_45334,N_45335,N_45336,N_45337,N_45338,N_45339,N_45340,N_45341,N_45342,N_45343,N_45344,N_45345,N_45346,N_45347,N_45348,N_45349,N_45350,N_45351,N_45352,N_45353,N_45354,N_45355,N_45356,N_45357,N_45358,N_45359,N_45360,N_45361,N_45362,N_45363,N_45364,N_45365,N_45366,N_45367,N_45368,N_45369,N_45370,N_45371,N_45372,N_45373,N_45374,N_45375,N_45376,N_45377,N_45378,N_45379,N_45380,N_45381,N_45382,N_45383,N_45384,N_45385,N_45386,N_45387,N_45388,N_45389,N_45390,N_45391,N_45392,N_45393,N_45394,N_45395,N_45396,N_45397,N_45398,N_45399,N_45400,N_45401,N_45402,N_45403,N_45404,N_45405,N_45406,N_45407,N_45408,N_45409,N_45410,N_45411,N_45412,N_45413,N_45414,N_45415,N_45416,N_45417,N_45418,N_45419,N_45420,N_45421,N_45422,N_45423,N_45424,N_45425,N_45426,N_45427,N_45428,N_45429,N_45430,N_45431,N_45432,N_45433,N_45434,N_45435,N_45436,N_45437,N_45438,N_45439,N_45440,N_45441,N_45442,N_45443,N_45444,N_45445,N_45446,N_45447,N_45448,N_45449,N_45450,N_45451,N_45452,N_45453,N_45454,N_45455,N_45456,N_45457,N_45458,N_45459,N_45460,N_45461,N_45462,N_45463,N_45464,N_45465,N_45466,N_45467,N_45468,N_45469,N_45470,N_45471,N_45472,N_45473,N_45474,N_45475,N_45476,N_45477,N_45478,N_45479,N_45480,N_45481,N_45482,N_45483,N_45484,N_45485,N_45486,N_45487,N_45488,N_45489,N_45490,N_45491,N_45492,N_45493,N_45494,N_45495,N_45496,N_45497,N_45498,N_45499,N_45500,N_45501,N_45502,N_45503,N_45504,N_45505,N_45506,N_45507,N_45508,N_45509,N_45510,N_45511,N_45512,N_45513,N_45514,N_45515,N_45516,N_45517,N_45518,N_45519,N_45520,N_45521,N_45522,N_45523,N_45524,N_45525,N_45526,N_45527,N_45528,N_45529,N_45530,N_45531,N_45532,N_45533,N_45534,N_45535,N_45536,N_45537,N_45538,N_45539,N_45540,N_45541,N_45542,N_45543,N_45544,N_45545,N_45546,N_45547,N_45548,N_45549,N_45550,N_45551,N_45552,N_45553,N_45554,N_45555,N_45556,N_45557,N_45558,N_45559,N_45560,N_45561,N_45562,N_45563,N_45564,N_45565,N_45566,N_45567,N_45568,N_45569,N_45570,N_45571,N_45572,N_45573,N_45574,N_45575,N_45576,N_45577,N_45578,N_45579,N_45580,N_45581,N_45582,N_45583,N_45584,N_45585,N_45586,N_45587,N_45588,N_45589,N_45590,N_45591,N_45592,N_45593,N_45594,N_45595,N_45596,N_45597,N_45598,N_45599,N_45600,N_45601,N_45602,N_45603,N_45604,N_45605,N_45606,N_45607,N_45608,N_45609,N_45610,N_45611,N_45612,N_45613,N_45614,N_45615,N_45616,N_45617,N_45618,N_45619,N_45620,N_45621,N_45622,N_45623,N_45624,N_45625,N_45626,N_45627,N_45628,N_45629,N_45630,N_45631,N_45632,N_45633,N_45634,N_45635,N_45636,N_45637,N_45638,N_45639,N_45640,N_45641,N_45642,N_45643,N_45644,N_45645,N_45646,N_45647,N_45648,N_45649,N_45650,N_45651,N_45652,N_45653,N_45654,N_45655,N_45656,N_45657,N_45658,N_45659,N_45660,N_45661,N_45662,N_45663,N_45664,N_45665,N_45666,N_45667,N_45668,N_45669,N_45670,N_45671,N_45672,N_45673,N_45674,N_45675,N_45676,N_45677,N_45678,N_45679,N_45680,N_45681,N_45682,N_45683,N_45684,N_45685,N_45686,N_45687,N_45688,N_45689,N_45690,N_45691,N_45692,N_45693,N_45694,N_45695,N_45696,N_45697,N_45698,N_45699,N_45700,N_45701,N_45702,N_45703,N_45704,N_45705,N_45706,N_45707,N_45708,N_45709,N_45710,N_45711,N_45712,N_45713,N_45714,N_45715,N_45716,N_45717,N_45718,N_45719,N_45720,N_45721,N_45722,N_45723,N_45724,N_45725,N_45726,N_45727,N_45728,N_45729,N_45730,N_45731,N_45732,N_45733,N_45734,N_45735,N_45736,N_45737,N_45738,N_45739,N_45740,N_45741,N_45742,N_45743,N_45744,N_45745,N_45746,N_45747,N_45748,N_45749,N_45750,N_45751,N_45752,N_45753,N_45754,N_45755,N_45756,N_45757,N_45758,N_45759,N_45760,N_45761,N_45762,N_45763,N_45764,N_45765,N_45766,N_45767,N_45768,N_45769,N_45770,N_45771,N_45772,N_45773,N_45774,N_45775,N_45776,N_45777,N_45778,N_45779,N_45780,N_45781,N_45782,N_45783,N_45784,N_45785,N_45786,N_45787,N_45788,N_45789,N_45790,N_45791,N_45792,N_45793,N_45794,N_45795,N_45796,N_45797,N_45798,N_45799,N_45800,N_45801,N_45802,N_45803,N_45804,N_45805,N_45806,N_45807,N_45808,N_45809,N_45810,N_45811,N_45812,N_45813,N_45814,N_45815,N_45816,N_45817,N_45818,N_45819,N_45820,N_45821,N_45822,N_45823,N_45824,N_45825,N_45826,N_45827,N_45828,N_45829,N_45830,N_45831,N_45832,N_45833,N_45834,N_45835,N_45836,N_45837,N_45838,N_45839,N_45840,N_45841,N_45842,N_45843,N_45844,N_45845,N_45846,N_45847,N_45848,N_45849,N_45850,N_45851,N_45852,N_45853,N_45854,N_45855,N_45856,N_45857,N_45858,N_45859,N_45860,N_45861,N_45862,N_45863,N_45864,N_45865,N_45866,N_45867,N_45868,N_45869,N_45870,N_45871,N_45872,N_45873,N_45874,N_45875,N_45876,N_45877,N_45878,N_45879,N_45880,N_45881,N_45882,N_45883,N_45884,N_45885,N_45886,N_45887,N_45888,N_45889,N_45890,N_45891,N_45892,N_45893,N_45894,N_45895,N_45896,N_45897,N_45898,N_45899,N_45900,N_45901,N_45902,N_45903,N_45904,N_45905,N_45906,N_45907,N_45908,N_45909,N_45910,N_45911,N_45912,N_45913,N_45914,N_45915,N_45916,N_45917,N_45918,N_45919,N_45920,N_45921,N_45922,N_45923,N_45924,N_45925,N_45926,N_45927,N_45928,N_45929,N_45930,N_45931,N_45932,N_45933,N_45934,N_45935,N_45936,N_45937,N_45938,N_45939,N_45940,N_45941,N_45942,N_45943,N_45944,N_45945,N_45946,N_45947,N_45948,N_45949,N_45950,N_45951,N_45952,N_45953,N_45954,N_45955,N_45956,N_45957,N_45958,N_45959,N_45960,N_45961,N_45962,N_45963,N_45964,N_45965,N_45966,N_45967,N_45968,N_45969,N_45970,N_45971,N_45972,N_45973,N_45974,N_45975,N_45976,N_45977,N_45978,N_45979,N_45980,N_45981,N_45982,N_45983,N_45984,N_45985,N_45986,N_45987,N_45988,N_45989,N_45990,N_45991,N_45992,N_45993,N_45994,N_45995,N_45996,N_45997,N_45998,N_45999,N_46000,N_46001,N_46002,N_46003,N_46004,N_46005,N_46006,N_46007,N_46008,N_46009,N_46010,N_46011,N_46012,N_46013,N_46014,N_46015,N_46016,N_46017,N_46018,N_46019,N_46020,N_46021,N_46022,N_46023,N_46024,N_46025,N_46026,N_46027,N_46028,N_46029,N_46030,N_46031,N_46032,N_46033,N_46034,N_46035,N_46036,N_46037,N_46038,N_46039,N_46040,N_46041,N_46042,N_46043,N_46044,N_46045,N_46046,N_46047,N_46048,N_46049,N_46050,N_46051,N_46052,N_46053,N_46054,N_46055,N_46056,N_46057,N_46058,N_46059,N_46060,N_46061,N_46062,N_46063,N_46064,N_46065,N_46066,N_46067,N_46068,N_46069,N_46070,N_46071,N_46072,N_46073,N_46074,N_46075,N_46076,N_46077,N_46078,N_46079,N_46080,N_46081,N_46082,N_46083,N_46084,N_46085,N_46086,N_46087,N_46088,N_46089,N_46090,N_46091,N_46092,N_46093,N_46094,N_46095,N_46096,N_46097,N_46098,N_46099,N_46100,N_46101,N_46102,N_46103,N_46104,N_46105,N_46106,N_46107,N_46108,N_46109,N_46110,N_46111,N_46112,N_46113,N_46114,N_46115,N_46116,N_46117,N_46118,N_46119,N_46120,N_46121,N_46122,N_46123,N_46124,N_46125,N_46126,N_46127,N_46128,N_46129,N_46130,N_46131,N_46132,N_46133,N_46134,N_46135,N_46136,N_46137,N_46138,N_46139,N_46140,N_46141,N_46142,N_46143,N_46144,N_46145,N_46146,N_46147,N_46148,N_46149,N_46150,N_46151,N_46152,N_46153,N_46154,N_46155,N_46156,N_46157,N_46158,N_46159,N_46160,N_46161,N_46162,N_46163,N_46164,N_46165,N_46166,N_46167,N_46168,N_46169,N_46170,N_46171,N_46172,N_46173,N_46174,N_46175,N_46176,N_46177,N_46178,N_46179,N_46180,N_46181,N_46182,N_46183,N_46184,N_46185,N_46186,N_46187,N_46188,N_46189,N_46190,N_46191,N_46192,N_46193,N_46194,N_46195,N_46196,N_46197,N_46198,N_46199,N_46200,N_46201,N_46202,N_46203,N_46204,N_46205,N_46206,N_46207,N_46208,N_46209,N_46210,N_46211,N_46212,N_46213,N_46214,N_46215,N_46216,N_46217,N_46218,N_46219,N_46220,N_46221,N_46222,N_46223,N_46224,N_46225,N_46226,N_46227,N_46228,N_46229,N_46230,N_46231,N_46232,N_46233,N_46234,N_46235,N_46236,N_46237,N_46238,N_46239,N_46240,N_46241,N_46242,N_46243,N_46244,N_46245,N_46246,N_46247,N_46248,N_46249,N_46250,N_46251,N_46252,N_46253,N_46254,N_46255,N_46256,N_46257,N_46258,N_46259,N_46260,N_46261,N_46262,N_46263,N_46264,N_46265,N_46266,N_46267,N_46268,N_46269,N_46270,N_46271,N_46272,N_46273,N_46274,N_46275,N_46276,N_46277,N_46278,N_46279,N_46280,N_46281,N_46282,N_46283,N_46284,N_46285,N_46286,N_46287,N_46288,N_46289,N_46290,N_46291,N_46292,N_46293,N_46294,N_46295,N_46296,N_46297,N_46298,N_46299,N_46300,N_46301,N_46302,N_46303,N_46304,N_46305,N_46306,N_46307,N_46308,N_46309,N_46310,N_46311,N_46312,N_46313,N_46314,N_46315,N_46316,N_46317,N_46318,N_46319,N_46320,N_46321,N_46322,N_46323,N_46324,N_46325,N_46326,N_46327,N_46328,N_46329,N_46330,N_46331,N_46332,N_46333,N_46334,N_46335,N_46336,N_46337,N_46338,N_46339,N_46340,N_46341,N_46342,N_46343,N_46344,N_46345,N_46346,N_46347,N_46348,N_46349,N_46350,N_46351,N_46352,N_46353,N_46354,N_46355,N_46356,N_46357,N_46358,N_46359,N_46360,N_46361,N_46362,N_46363,N_46364,N_46365,N_46366,N_46367,N_46368,N_46369,N_46370,N_46371,N_46372,N_46373,N_46374,N_46375,N_46376,N_46377,N_46378,N_46379,N_46380,N_46381,N_46382,N_46383,N_46384,N_46385,N_46386,N_46387,N_46388,N_46389,N_46390,N_46391,N_46392,N_46393,N_46394,N_46395,N_46396,N_46397,N_46398,N_46399,N_46400,N_46401,N_46402,N_46403,N_46404,N_46405,N_46406,N_46407,N_46408,N_46409,N_46410,N_46411,N_46412,N_46413,N_46414,N_46415,N_46416,N_46417,N_46418,N_46419,N_46420,N_46421,N_46422,N_46423,N_46424,N_46425,N_46426,N_46427,N_46428,N_46429,N_46430,N_46431,N_46432,N_46433,N_46434,N_46435,N_46436,N_46437,N_46438,N_46439,N_46440,N_46441,N_46442,N_46443,N_46444,N_46445,N_46446,N_46447,N_46448,N_46449,N_46450,N_46451,N_46452,N_46453,N_46454,N_46455,N_46456,N_46457,N_46458,N_46459,N_46460,N_46461,N_46462,N_46463,N_46464,N_46465,N_46466,N_46467,N_46468,N_46469,N_46470,N_46471,N_46472,N_46473,N_46474,N_46475,N_46476,N_46477,N_46478,N_46479,N_46480,N_46481,N_46482,N_46483,N_46484,N_46485,N_46486,N_46487,N_46488,N_46489,N_46490,N_46491,N_46492,N_46493,N_46494,N_46495,N_46496,N_46497,N_46498,N_46499,N_46500,N_46501,N_46502,N_46503,N_46504,N_46505,N_46506,N_46507,N_46508,N_46509,N_46510,N_46511,N_46512,N_46513,N_46514,N_46515,N_46516,N_46517,N_46518,N_46519,N_46520,N_46521,N_46522,N_46523,N_46524,N_46525,N_46526,N_46527,N_46528,N_46529,N_46530,N_46531,N_46532,N_46533,N_46534,N_46535,N_46536,N_46537,N_46538,N_46539,N_46540,N_46541,N_46542,N_46543,N_46544,N_46545,N_46546,N_46547,N_46548,N_46549,N_46550,N_46551,N_46552,N_46553,N_46554,N_46555,N_46556,N_46557,N_46558,N_46559,N_46560,N_46561,N_46562,N_46563,N_46564,N_46565,N_46566,N_46567,N_46568,N_46569,N_46570,N_46571,N_46572,N_46573,N_46574,N_46575,N_46576,N_46577,N_46578,N_46579,N_46580,N_46581,N_46582,N_46583,N_46584,N_46585,N_46586,N_46587,N_46588,N_46589,N_46590,N_46591,N_46592,N_46593,N_46594,N_46595,N_46596,N_46597,N_46598,N_46599,N_46600,N_46601,N_46602,N_46603,N_46604,N_46605,N_46606,N_46607,N_46608,N_46609,N_46610,N_46611,N_46612,N_46613,N_46614,N_46615,N_46616,N_46617,N_46618,N_46619,N_46620,N_46621,N_46622,N_46623,N_46624,N_46625,N_46626,N_46627,N_46628,N_46629,N_46630,N_46631,N_46632,N_46633,N_46634,N_46635,N_46636,N_46637,N_46638,N_46639,N_46640,N_46641,N_46642,N_46643,N_46644,N_46645,N_46646,N_46647,N_46648,N_46649,N_46650,N_46651,N_46652,N_46653,N_46654,N_46655,N_46656,N_46657,N_46658,N_46659,N_46660,N_46661,N_46662,N_46663,N_46664,N_46665,N_46666,N_46667,N_46668,N_46669,N_46670,N_46671,N_46672,N_46673,N_46674,N_46675,N_46676,N_46677,N_46678,N_46679,N_46680,N_46681,N_46682,N_46683,N_46684,N_46685,N_46686,N_46687,N_46688,N_46689,N_46690,N_46691,N_46692,N_46693,N_46694,N_46695,N_46696,N_46697,N_46698,N_46699,N_46700,N_46701,N_46702,N_46703,N_46704,N_46705,N_46706,N_46707,N_46708,N_46709,N_46710,N_46711,N_46712,N_46713,N_46714,N_46715,N_46716,N_46717,N_46718,N_46719,N_46720,N_46721,N_46722,N_46723,N_46724,N_46725,N_46726,N_46727,N_46728,N_46729,N_46730,N_46731,N_46732,N_46733,N_46734,N_46735,N_46736,N_46737,N_46738,N_46739,N_46740,N_46741,N_46742,N_46743,N_46744,N_46745,N_46746,N_46747,N_46748,N_46749,N_46750,N_46751,N_46752,N_46753,N_46754,N_46755,N_46756,N_46757,N_46758,N_46759,N_46760,N_46761,N_46762,N_46763,N_46764,N_46765,N_46766,N_46767,N_46768,N_46769,N_46770,N_46771,N_46772,N_46773,N_46774,N_46775,N_46776,N_46777,N_46778,N_46779,N_46780,N_46781,N_46782,N_46783,N_46784,N_46785,N_46786,N_46787,N_46788,N_46789,N_46790,N_46791,N_46792,N_46793,N_46794,N_46795,N_46796,N_46797,N_46798,N_46799,N_46800,N_46801,N_46802,N_46803,N_46804,N_46805,N_46806,N_46807,N_46808,N_46809,N_46810,N_46811,N_46812,N_46813,N_46814,N_46815,N_46816,N_46817,N_46818,N_46819,N_46820,N_46821,N_46822,N_46823,N_46824,N_46825,N_46826,N_46827,N_46828,N_46829,N_46830,N_46831,N_46832,N_46833,N_46834,N_46835,N_46836,N_46837,N_46838,N_46839,N_46840,N_46841,N_46842,N_46843,N_46844,N_46845,N_46846,N_46847,N_46848,N_46849,N_46850,N_46851,N_46852,N_46853,N_46854,N_46855,N_46856,N_46857,N_46858,N_46859,N_46860,N_46861,N_46862,N_46863,N_46864,N_46865,N_46866,N_46867,N_46868,N_46869,N_46870,N_46871,N_46872,N_46873,N_46874,N_46875,N_46876,N_46877,N_46878,N_46879,N_46880,N_46881,N_46882,N_46883,N_46884,N_46885,N_46886,N_46887,N_46888,N_46889,N_46890,N_46891,N_46892,N_46893,N_46894,N_46895,N_46896,N_46897,N_46898,N_46899,N_46900,N_46901,N_46902,N_46903,N_46904,N_46905,N_46906,N_46907,N_46908,N_46909,N_46910,N_46911,N_46912,N_46913,N_46914,N_46915,N_46916,N_46917,N_46918,N_46919,N_46920,N_46921,N_46922,N_46923,N_46924,N_46925,N_46926,N_46927,N_46928,N_46929,N_46930,N_46931,N_46932,N_46933,N_46934,N_46935,N_46936,N_46937,N_46938,N_46939,N_46940,N_46941,N_46942,N_46943,N_46944,N_46945,N_46946,N_46947,N_46948,N_46949,N_46950,N_46951,N_46952,N_46953,N_46954,N_46955,N_46956,N_46957,N_46958,N_46959,N_46960,N_46961,N_46962,N_46963,N_46964,N_46965,N_46966,N_46967,N_46968,N_46969,N_46970,N_46971,N_46972,N_46973,N_46974,N_46975,N_46976,N_46977,N_46978,N_46979,N_46980,N_46981,N_46982,N_46983,N_46984,N_46985,N_46986,N_46987,N_46988,N_46989,N_46990,N_46991,N_46992,N_46993,N_46994,N_46995,N_46996,N_46997,N_46998,N_46999,N_47000,N_47001,N_47002,N_47003,N_47004,N_47005,N_47006,N_47007,N_47008,N_47009,N_47010,N_47011,N_47012,N_47013,N_47014,N_47015,N_47016,N_47017,N_47018,N_47019,N_47020,N_47021,N_47022,N_47023,N_47024,N_47025,N_47026,N_47027,N_47028,N_47029,N_47030,N_47031,N_47032,N_47033,N_47034,N_47035,N_47036,N_47037,N_47038,N_47039,N_47040,N_47041,N_47042,N_47043,N_47044,N_47045,N_47046,N_47047,N_47048,N_47049,N_47050,N_47051,N_47052,N_47053,N_47054,N_47055,N_47056,N_47057,N_47058,N_47059,N_47060,N_47061,N_47062,N_47063,N_47064,N_47065,N_47066,N_47067,N_47068,N_47069,N_47070,N_47071,N_47072,N_47073,N_47074,N_47075,N_47076,N_47077,N_47078,N_47079,N_47080,N_47081,N_47082,N_47083,N_47084,N_47085,N_47086,N_47087,N_47088,N_47089,N_47090,N_47091,N_47092,N_47093,N_47094,N_47095,N_47096,N_47097,N_47098,N_47099,N_47100,N_47101,N_47102,N_47103,N_47104,N_47105,N_47106,N_47107,N_47108,N_47109,N_47110,N_47111,N_47112,N_47113,N_47114,N_47115,N_47116,N_47117,N_47118,N_47119,N_47120,N_47121,N_47122,N_47123,N_47124,N_47125,N_47126,N_47127,N_47128,N_47129,N_47130,N_47131,N_47132,N_47133,N_47134,N_47135,N_47136,N_47137,N_47138,N_47139,N_47140,N_47141,N_47142,N_47143,N_47144,N_47145,N_47146,N_47147,N_47148,N_47149,N_47150,N_47151,N_47152,N_47153,N_47154,N_47155,N_47156,N_47157,N_47158,N_47159,N_47160,N_47161,N_47162,N_47163,N_47164,N_47165,N_47166,N_47167,N_47168,N_47169,N_47170,N_47171,N_47172,N_47173,N_47174,N_47175,N_47176,N_47177,N_47178,N_47179,N_47180,N_47181,N_47182,N_47183,N_47184,N_47185,N_47186,N_47187,N_47188,N_47189,N_47190,N_47191,N_47192,N_47193,N_47194,N_47195,N_47196,N_47197,N_47198,N_47199,N_47200,N_47201,N_47202,N_47203,N_47204,N_47205,N_47206,N_47207,N_47208,N_47209,N_47210,N_47211,N_47212,N_47213,N_47214,N_47215,N_47216,N_47217,N_47218,N_47219,N_47220,N_47221,N_47222,N_47223,N_47224,N_47225,N_47226,N_47227,N_47228,N_47229,N_47230,N_47231,N_47232,N_47233,N_47234,N_47235,N_47236,N_47237,N_47238,N_47239,N_47240,N_47241,N_47242,N_47243,N_47244,N_47245,N_47246,N_47247,N_47248,N_47249,N_47250,N_47251,N_47252,N_47253,N_47254,N_47255,N_47256,N_47257,N_47258,N_47259,N_47260,N_47261,N_47262,N_47263,N_47264,N_47265,N_47266,N_47267,N_47268,N_47269,N_47270,N_47271,N_47272,N_47273,N_47274,N_47275,N_47276,N_47277,N_47278,N_47279,N_47280,N_47281,N_47282,N_47283,N_47284,N_47285,N_47286,N_47287,N_47288,N_47289,N_47290,N_47291,N_47292,N_47293,N_47294,N_47295,N_47296,N_47297,N_47298,N_47299,N_47300,N_47301,N_47302,N_47303,N_47304,N_47305,N_47306,N_47307,N_47308,N_47309,N_47310,N_47311,N_47312,N_47313,N_47314,N_47315,N_47316,N_47317,N_47318,N_47319,N_47320,N_47321,N_47322,N_47323,N_47324,N_47325,N_47326,N_47327,N_47328,N_47329,N_47330,N_47331,N_47332,N_47333,N_47334,N_47335,N_47336,N_47337,N_47338,N_47339,N_47340,N_47341,N_47342,N_47343,N_47344,N_47345,N_47346,N_47347,N_47348,N_47349,N_47350,N_47351,N_47352,N_47353,N_47354,N_47355,N_47356,N_47357,N_47358,N_47359,N_47360,N_47361,N_47362,N_47363,N_47364,N_47365,N_47366,N_47367,N_47368,N_47369,N_47370,N_47371,N_47372,N_47373,N_47374,N_47375,N_47376,N_47377,N_47378,N_47379,N_47380,N_47381,N_47382,N_47383,N_47384,N_47385,N_47386,N_47387,N_47388,N_47389,N_47390,N_47391,N_47392,N_47393,N_47394,N_47395,N_47396,N_47397,N_47398,N_47399,N_47400,N_47401,N_47402,N_47403,N_47404,N_47405,N_47406,N_47407,N_47408,N_47409,N_47410,N_47411,N_47412,N_47413,N_47414,N_47415,N_47416,N_47417,N_47418,N_47419,N_47420,N_47421,N_47422,N_47423,N_47424,N_47425,N_47426,N_47427,N_47428,N_47429,N_47430,N_47431,N_47432,N_47433,N_47434,N_47435,N_47436,N_47437,N_47438,N_47439,N_47440,N_47441,N_47442,N_47443,N_47444,N_47445,N_47446,N_47447,N_47448,N_47449,N_47450,N_47451,N_47452,N_47453,N_47454,N_47455,N_47456,N_47457,N_47458,N_47459,N_47460,N_47461,N_47462,N_47463,N_47464,N_47465,N_47466,N_47467,N_47468,N_47469,N_47470,N_47471,N_47472,N_47473,N_47474,N_47475,N_47476,N_47477,N_47478,N_47479,N_47480,N_47481,N_47482,N_47483,N_47484,N_47485,N_47486,N_47487,N_47488,N_47489,N_47490,N_47491,N_47492,N_47493,N_47494,N_47495,N_47496,N_47497,N_47498,N_47499,N_47500,N_47501,N_47502,N_47503,N_47504,N_47505,N_47506,N_47507,N_47508,N_47509,N_47510,N_47511,N_47512,N_47513,N_47514,N_47515,N_47516,N_47517,N_47518,N_47519,N_47520,N_47521,N_47522,N_47523,N_47524,N_47525,N_47526,N_47527,N_47528,N_47529,N_47530,N_47531,N_47532,N_47533,N_47534,N_47535,N_47536,N_47537,N_47538,N_47539,N_47540,N_47541,N_47542,N_47543,N_47544,N_47545,N_47546,N_47547,N_47548,N_47549,N_47550,N_47551,N_47552,N_47553,N_47554,N_47555,N_47556,N_47557,N_47558,N_47559,N_47560,N_47561,N_47562,N_47563,N_47564,N_47565,N_47566,N_47567,N_47568,N_47569,N_47570,N_47571,N_47572,N_47573,N_47574,N_47575,N_47576,N_47577,N_47578,N_47579,N_47580,N_47581,N_47582,N_47583,N_47584,N_47585,N_47586,N_47587,N_47588,N_47589,N_47590,N_47591,N_47592,N_47593,N_47594,N_47595,N_47596,N_47597,N_47598,N_47599,N_47600,N_47601,N_47602,N_47603,N_47604,N_47605,N_47606,N_47607,N_47608,N_47609,N_47610,N_47611,N_47612,N_47613,N_47614,N_47615,N_47616,N_47617,N_47618,N_47619,N_47620,N_47621,N_47622,N_47623,N_47624,N_47625,N_47626,N_47627,N_47628,N_47629,N_47630,N_47631,N_47632,N_47633,N_47634,N_47635,N_47636,N_47637,N_47638,N_47639,N_47640,N_47641,N_47642,N_47643,N_47644,N_47645,N_47646,N_47647,N_47648,N_47649,N_47650,N_47651,N_47652,N_47653,N_47654,N_47655,N_47656,N_47657,N_47658,N_47659,N_47660,N_47661,N_47662,N_47663,N_47664,N_47665,N_47666,N_47667,N_47668,N_47669,N_47670,N_47671,N_47672,N_47673,N_47674,N_47675,N_47676,N_47677,N_47678,N_47679,N_47680,N_47681,N_47682,N_47683,N_47684,N_47685,N_47686,N_47687,N_47688,N_47689,N_47690,N_47691,N_47692,N_47693,N_47694,N_47695,N_47696,N_47697,N_47698,N_47699,N_47700,N_47701,N_47702,N_47703,N_47704,N_47705,N_47706,N_47707,N_47708,N_47709,N_47710,N_47711,N_47712,N_47713,N_47714,N_47715,N_47716,N_47717,N_47718,N_47719,N_47720,N_47721,N_47722,N_47723,N_47724,N_47725,N_47726,N_47727,N_47728,N_47729,N_47730,N_47731,N_47732,N_47733,N_47734,N_47735,N_47736,N_47737,N_47738,N_47739,N_47740,N_47741,N_47742,N_47743,N_47744,N_47745,N_47746,N_47747,N_47748,N_47749,N_47750,N_47751,N_47752,N_47753,N_47754,N_47755,N_47756,N_47757,N_47758,N_47759,N_47760,N_47761,N_47762,N_47763,N_47764,N_47765,N_47766,N_47767,N_47768,N_47769,N_47770,N_47771,N_47772,N_47773,N_47774,N_47775,N_47776,N_47777,N_47778,N_47779,N_47780,N_47781,N_47782,N_47783,N_47784,N_47785,N_47786,N_47787,N_47788,N_47789,N_47790,N_47791,N_47792,N_47793,N_47794,N_47795,N_47796,N_47797,N_47798,N_47799,N_47800,N_47801,N_47802,N_47803,N_47804,N_47805,N_47806,N_47807,N_47808,N_47809,N_47810,N_47811,N_47812,N_47813,N_47814,N_47815,N_47816,N_47817,N_47818,N_47819,N_47820,N_47821,N_47822,N_47823,N_47824,N_47825,N_47826,N_47827,N_47828,N_47829,N_47830,N_47831,N_47832,N_47833,N_47834,N_47835,N_47836,N_47837,N_47838,N_47839,N_47840,N_47841,N_47842,N_47843,N_47844,N_47845,N_47846,N_47847,N_47848,N_47849,N_47850,N_47851,N_47852,N_47853,N_47854,N_47855,N_47856,N_47857,N_47858,N_47859,N_47860,N_47861,N_47862,N_47863,N_47864,N_47865,N_47866,N_47867,N_47868,N_47869,N_47870,N_47871,N_47872,N_47873,N_47874,N_47875,N_47876,N_47877,N_47878,N_47879,N_47880,N_47881,N_47882,N_47883,N_47884,N_47885,N_47886,N_47887,N_47888,N_47889,N_47890,N_47891,N_47892,N_47893,N_47894,N_47895,N_47896,N_47897,N_47898,N_47899,N_47900,N_47901,N_47902,N_47903,N_47904,N_47905,N_47906,N_47907,N_47908,N_47909,N_47910,N_47911,N_47912,N_47913,N_47914,N_47915,N_47916,N_47917,N_47918,N_47919,N_47920,N_47921,N_47922,N_47923,N_47924,N_47925,N_47926,N_47927,N_47928,N_47929,N_47930,N_47931,N_47932,N_47933,N_47934,N_47935,N_47936,N_47937,N_47938,N_47939,N_47940,N_47941,N_47942,N_47943,N_47944,N_47945,N_47946,N_47947,N_47948,N_47949,N_47950,N_47951,N_47952,N_47953,N_47954,N_47955,N_47956,N_47957,N_47958,N_47959,N_47960,N_47961,N_47962,N_47963,N_47964,N_47965,N_47966,N_47967,N_47968,N_47969,N_47970,N_47971,N_47972,N_47973,N_47974,N_47975,N_47976,N_47977,N_47978,N_47979,N_47980,N_47981,N_47982,N_47983,N_47984,N_47985,N_47986,N_47987,N_47988,N_47989,N_47990,N_47991,N_47992,N_47993,N_47994,N_47995,N_47996,N_47997,N_47998,N_47999,N_48000,N_48001,N_48002,N_48003,N_48004,N_48005,N_48006,N_48007,N_48008,N_48009,N_48010,N_48011,N_48012,N_48013,N_48014,N_48015,N_48016,N_48017,N_48018,N_48019,N_48020,N_48021,N_48022,N_48023,N_48024,N_48025,N_48026,N_48027,N_48028,N_48029,N_48030,N_48031,N_48032,N_48033,N_48034,N_48035,N_48036,N_48037,N_48038,N_48039,N_48040,N_48041,N_48042,N_48043,N_48044,N_48045,N_48046,N_48047,N_48048,N_48049,N_48050,N_48051,N_48052,N_48053,N_48054,N_48055,N_48056,N_48057,N_48058,N_48059,N_48060,N_48061,N_48062,N_48063,N_48064,N_48065,N_48066,N_48067,N_48068,N_48069,N_48070,N_48071,N_48072,N_48073,N_48074,N_48075,N_48076,N_48077,N_48078,N_48079,N_48080,N_48081,N_48082,N_48083,N_48084,N_48085,N_48086,N_48087,N_48088,N_48089,N_48090,N_48091,N_48092,N_48093,N_48094,N_48095,N_48096,N_48097,N_48098,N_48099,N_48100,N_48101,N_48102,N_48103,N_48104,N_48105,N_48106,N_48107,N_48108,N_48109,N_48110,N_48111,N_48112,N_48113,N_48114,N_48115,N_48116,N_48117,N_48118,N_48119,N_48120,N_48121,N_48122,N_48123,N_48124,N_48125,N_48126,N_48127,N_48128,N_48129,N_48130,N_48131,N_48132,N_48133,N_48134,N_48135,N_48136,N_48137,N_48138,N_48139,N_48140,N_48141,N_48142,N_48143,N_48144,N_48145,N_48146,N_48147,N_48148,N_48149,N_48150,N_48151,N_48152,N_48153,N_48154,N_48155,N_48156,N_48157,N_48158,N_48159,N_48160,N_48161,N_48162,N_48163,N_48164,N_48165,N_48166,N_48167,N_48168,N_48169,N_48170,N_48171,N_48172,N_48173,N_48174,N_48175,N_48176,N_48177,N_48178,N_48179,N_48180,N_48181,N_48182,N_48183,N_48184,N_48185,N_48186,N_48187,N_48188,N_48189,N_48190,N_48191,N_48192,N_48193,N_48194,N_48195,N_48196,N_48197,N_48198,N_48199,N_48200,N_48201,N_48202,N_48203,N_48204,N_48205,N_48206,N_48207,N_48208,N_48209,N_48210,N_48211,N_48212,N_48213,N_48214,N_48215,N_48216,N_48217,N_48218,N_48219,N_48220,N_48221,N_48222,N_48223,N_48224,N_48225,N_48226,N_48227,N_48228,N_48229,N_48230,N_48231,N_48232,N_48233,N_48234,N_48235,N_48236,N_48237,N_48238,N_48239,N_48240,N_48241,N_48242,N_48243,N_48244,N_48245,N_48246,N_48247,N_48248,N_48249,N_48250,N_48251,N_48252,N_48253,N_48254,N_48255,N_48256,N_48257,N_48258,N_48259,N_48260,N_48261,N_48262,N_48263,N_48264,N_48265,N_48266,N_48267,N_48268,N_48269,N_48270,N_48271,N_48272,N_48273,N_48274,N_48275,N_48276,N_48277,N_48278,N_48279,N_48280,N_48281,N_48282,N_48283,N_48284,N_48285,N_48286,N_48287,N_48288,N_48289,N_48290,N_48291,N_48292,N_48293,N_48294,N_48295,N_48296,N_48297,N_48298,N_48299,N_48300,N_48301,N_48302,N_48303,N_48304,N_48305,N_48306,N_48307,N_48308,N_48309,N_48310,N_48311,N_48312,N_48313,N_48314,N_48315,N_48316,N_48317,N_48318,N_48319,N_48320,N_48321,N_48322,N_48323,N_48324,N_48325,N_48326,N_48327,N_48328,N_48329,N_48330,N_48331,N_48332,N_48333,N_48334,N_48335,N_48336,N_48337,N_48338,N_48339,N_48340,N_48341,N_48342,N_48343,N_48344,N_48345,N_48346,N_48347,N_48348,N_48349,N_48350,N_48351,N_48352,N_48353,N_48354,N_48355,N_48356,N_48357,N_48358,N_48359,N_48360,N_48361,N_48362,N_48363,N_48364,N_48365,N_48366,N_48367,N_48368,N_48369,N_48370,N_48371,N_48372,N_48373,N_48374,N_48375,N_48376,N_48377,N_48378,N_48379,N_48380,N_48381,N_48382,N_48383,N_48384,N_48385,N_48386,N_48387,N_48388,N_48389,N_48390,N_48391,N_48392,N_48393,N_48394,N_48395,N_48396,N_48397,N_48398,N_48399,N_48400,N_48401,N_48402,N_48403,N_48404,N_48405,N_48406,N_48407,N_48408,N_48409,N_48410,N_48411,N_48412,N_48413,N_48414,N_48415,N_48416,N_48417,N_48418,N_48419,N_48420,N_48421,N_48422,N_48423,N_48424,N_48425,N_48426,N_48427,N_48428,N_48429,N_48430,N_48431,N_48432,N_48433,N_48434,N_48435,N_48436,N_48437,N_48438,N_48439,N_48440,N_48441,N_48442,N_48443,N_48444,N_48445,N_48446,N_48447,N_48448,N_48449,N_48450,N_48451,N_48452,N_48453,N_48454,N_48455,N_48456,N_48457,N_48458,N_48459,N_48460,N_48461,N_48462,N_48463,N_48464,N_48465,N_48466,N_48467,N_48468,N_48469,N_48470,N_48471,N_48472,N_48473,N_48474,N_48475,N_48476,N_48477,N_48478,N_48479,N_48480,N_48481,N_48482,N_48483,N_48484,N_48485,N_48486,N_48487,N_48488,N_48489,N_48490,N_48491,N_48492,N_48493,N_48494,N_48495,N_48496,N_48497,N_48498,N_48499,N_48500,N_48501,N_48502,N_48503,N_48504,N_48505,N_48506,N_48507,N_48508,N_48509,N_48510,N_48511,N_48512,N_48513,N_48514,N_48515,N_48516,N_48517,N_48518,N_48519,N_48520,N_48521,N_48522,N_48523,N_48524,N_48525,N_48526,N_48527,N_48528,N_48529,N_48530,N_48531,N_48532,N_48533,N_48534,N_48535,N_48536,N_48537,N_48538,N_48539,N_48540,N_48541,N_48542,N_48543,N_48544,N_48545,N_48546,N_48547,N_48548,N_48549,N_48550,N_48551,N_48552,N_48553,N_48554,N_48555,N_48556,N_48557,N_48558,N_48559,N_48560,N_48561,N_48562,N_48563,N_48564,N_48565,N_48566,N_48567,N_48568,N_48569,N_48570,N_48571,N_48572,N_48573,N_48574,N_48575,N_48576,N_48577,N_48578,N_48579,N_48580,N_48581,N_48582,N_48583,N_48584,N_48585,N_48586,N_48587,N_48588,N_48589,N_48590,N_48591,N_48592,N_48593,N_48594,N_48595,N_48596,N_48597,N_48598,N_48599,N_48600,N_48601,N_48602,N_48603,N_48604,N_48605,N_48606,N_48607,N_48608,N_48609,N_48610,N_48611,N_48612,N_48613,N_48614,N_48615,N_48616,N_48617,N_48618,N_48619,N_48620,N_48621,N_48622,N_48623,N_48624,N_48625,N_48626,N_48627,N_48628,N_48629,N_48630,N_48631,N_48632,N_48633,N_48634,N_48635,N_48636,N_48637,N_48638,N_48639,N_48640,N_48641,N_48642,N_48643,N_48644,N_48645,N_48646,N_48647,N_48648,N_48649,N_48650,N_48651,N_48652,N_48653,N_48654,N_48655,N_48656,N_48657,N_48658,N_48659,N_48660,N_48661,N_48662,N_48663,N_48664,N_48665,N_48666,N_48667,N_48668,N_48669,N_48670,N_48671,N_48672,N_48673,N_48674,N_48675,N_48676,N_48677,N_48678,N_48679,N_48680,N_48681,N_48682,N_48683,N_48684,N_48685,N_48686,N_48687,N_48688,N_48689,N_48690,N_48691,N_48692,N_48693,N_48694,N_48695,N_48696,N_48697,N_48698,N_48699,N_48700,N_48701,N_48702,N_48703,N_48704,N_48705,N_48706,N_48707,N_48708,N_48709,N_48710,N_48711,N_48712,N_48713,N_48714,N_48715,N_48716,N_48717,N_48718,N_48719,N_48720,N_48721,N_48722,N_48723,N_48724,N_48725,N_48726,N_48727,N_48728,N_48729,N_48730,N_48731,N_48732,N_48733,N_48734,N_48735,N_48736,N_48737,N_48738,N_48739,N_48740,N_48741,N_48742,N_48743,N_48744,N_48745,N_48746,N_48747,N_48748,N_48749,N_48750,N_48751,N_48752,N_48753,N_48754,N_48755,N_48756,N_48757,N_48758,N_48759,N_48760,N_48761,N_48762,N_48763,N_48764,N_48765,N_48766,N_48767,N_48768,N_48769,N_48770,N_48771,N_48772,N_48773,N_48774,N_48775,N_48776,N_48777,N_48778,N_48779,N_48780,N_48781,N_48782,N_48783,N_48784,N_48785,N_48786,N_48787,N_48788,N_48789,N_48790,N_48791,N_48792,N_48793,N_48794,N_48795,N_48796,N_48797,N_48798,N_48799,N_48800,N_48801,N_48802,N_48803,N_48804,N_48805,N_48806,N_48807,N_48808,N_48809,N_48810,N_48811,N_48812,N_48813,N_48814,N_48815,N_48816,N_48817,N_48818,N_48819,N_48820,N_48821,N_48822,N_48823,N_48824,N_48825,N_48826,N_48827,N_48828,N_48829,N_48830,N_48831,N_48832,N_48833,N_48834,N_48835,N_48836,N_48837,N_48838,N_48839,N_48840,N_48841,N_48842,N_48843,N_48844,N_48845,N_48846,N_48847,N_48848,N_48849,N_48850,N_48851,N_48852,N_48853,N_48854,N_48855,N_48856,N_48857,N_48858,N_48859,N_48860,N_48861,N_48862,N_48863,N_48864,N_48865,N_48866,N_48867,N_48868,N_48869,N_48870,N_48871,N_48872,N_48873,N_48874,N_48875,N_48876,N_48877,N_48878,N_48879,N_48880,N_48881,N_48882,N_48883,N_48884,N_48885,N_48886,N_48887,N_48888,N_48889,N_48890,N_48891,N_48892,N_48893,N_48894,N_48895,N_48896,N_48897,N_48898,N_48899,N_48900,N_48901,N_48902,N_48903,N_48904,N_48905,N_48906,N_48907,N_48908,N_48909,N_48910,N_48911,N_48912,N_48913,N_48914,N_48915,N_48916,N_48917,N_48918,N_48919,N_48920,N_48921,N_48922,N_48923,N_48924,N_48925,N_48926,N_48927,N_48928,N_48929,N_48930,N_48931,N_48932,N_48933,N_48934,N_48935,N_48936,N_48937,N_48938,N_48939,N_48940,N_48941,N_48942,N_48943,N_48944,N_48945,N_48946,N_48947,N_48948,N_48949,N_48950,N_48951,N_48952,N_48953,N_48954,N_48955,N_48956,N_48957,N_48958,N_48959,N_48960,N_48961,N_48962,N_48963,N_48964,N_48965,N_48966,N_48967,N_48968,N_48969,N_48970,N_48971,N_48972,N_48973,N_48974,N_48975,N_48976,N_48977,N_48978,N_48979,N_48980,N_48981,N_48982,N_48983,N_48984,N_48985,N_48986,N_48987,N_48988,N_48989,N_48990,N_48991,N_48992,N_48993,N_48994,N_48995,N_48996,N_48997,N_48998,N_48999,N_49000,N_49001,N_49002,N_49003,N_49004,N_49005,N_49006,N_49007,N_49008,N_49009,N_49010,N_49011,N_49012,N_49013,N_49014,N_49015,N_49016,N_49017,N_49018,N_49019,N_49020,N_49021,N_49022,N_49023,N_49024,N_49025,N_49026,N_49027,N_49028,N_49029,N_49030,N_49031,N_49032,N_49033,N_49034,N_49035,N_49036,N_49037,N_49038,N_49039,N_49040,N_49041,N_49042,N_49043,N_49044,N_49045,N_49046,N_49047,N_49048,N_49049,N_49050,N_49051,N_49052,N_49053,N_49054,N_49055,N_49056,N_49057,N_49058,N_49059,N_49060,N_49061,N_49062,N_49063,N_49064,N_49065,N_49066,N_49067,N_49068,N_49069,N_49070,N_49071,N_49072,N_49073,N_49074,N_49075,N_49076,N_49077,N_49078,N_49079,N_49080,N_49081,N_49082,N_49083,N_49084,N_49085,N_49086,N_49087,N_49088,N_49089,N_49090,N_49091,N_49092,N_49093,N_49094,N_49095,N_49096,N_49097,N_49098,N_49099,N_49100,N_49101,N_49102,N_49103,N_49104,N_49105,N_49106,N_49107,N_49108,N_49109,N_49110,N_49111,N_49112,N_49113,N_49114,N_49115,N_49116,N_49117,N_49118,N_49119,N_49120,N_49121,N_49122,N_49123,N_49124,N_49125,N_49126,N_49127,N_49128,N_49129,N_49130,N_49131,N_49132,N_49133,N_49134,N_49135,N_49136,N_49137,N_49138,N_49139,N_49140,N_49141,N_49142,N_49143,N_49144,N_49145,N_49146,N_49147,N_49148,N_49149,N_49150,N_49151,N_49152,N_49153,N_49154,N_49155,N_49156,N_49157,N_49158,N_49159,N_49160,N_49161,N_49162,N_49163,N_49164,N_49165,N_49166,N_49167,N_49168,N_49169,N_49170,N_49171,N_49172,N_49173,N_49174,N_49175,N_49176,N_49177,N_49178,N_49179,N_49180,N_49181,N_49182,N_49183,N_49184,N_49185,N_49186,N_49187,N_49188,N_49189,N_49190,N_49191,N_49192,N_49193,N_49194,N_49195,N_49196,N_49197,N_49198,N_49199,N_49200,N_49201,N_49202,N_49203,N_49204,N_49205,N_49206,N_49207,N_49208,N_49209,N_49210,N_49211,N_49212,N_49213,N_49214,N_49215,N_49216,N_49217,N_49218,N_49219,N_49220,N_49221,N_49222,N_49223,N_49224,N_49225,N_49226,N_49227,N_49228,N_49229,N_49230,N_49231,N_49232,N_49233,N_49234,N_49235,N_49236,N_49237,N_49238,N_49239,N_49240,N_49241,N_49242,N_49243,N_49244,N_49245,N_49246,N_49247,N_49248,N_49249,N_49250,N_49251,N_49252,N_49253,N_49254,N_49255,N_49256,N_49257,N_49258,N_49259,N_49260,N_49261,N_49262,N_49263,N_49264,N_49265,N_49266,N_49267,N_49268,N_49269,N_49270,N_49271,N_49272,N_49273,N_49274,N_49275,N_49276,N_49277,N_49278,N_49279,N_49280,N_49281,N_49282,N_49283,N_49284,N_49285,N_49286,N_49287,N_49288,N_49289,N_49290,N_49291,N_49292,N_49293,N_49294,N_49295,N_49296,N_49297,N_49298,N_49299,N_49300,N_49301,N_49302,N_49303,N_49304,N_49305,N_49306,N_49307,N_49308,N_49309,N_49310,N_49311,N_49312,N_49313,N_49314,N_49315,N_49316,N_49317,N_49318,N_49319,N_49320,N_49321,N_49322,N_49323,N_49324,N_49325,N_49326,N_49327,N_49328,N_49329,N_49330,N_49331,N_49332,N_49333,N_49334,N_49335,N_49336,N_49337,N_49338,N_49339,N_49340,N_49341,N_49342,N_49343,N_49344,N_49345,N_49346,N_49347,N_49348,N_49349,N_49350,N_49351,N_49352,N_49353,N_49354,N_49355,N_49356,N_49357,N_49358,N_49359,N_49360,N_49361,N_49362,N_49363,N_49364,N_49365,N_49366,N_49367,N_49368,N_49369,N_49370,N_49371,N_49372,N_49373,N_49374,N_49375,N_49376,N_49377,N_49378,N_49379,N_49380,N_49381,N_49382,N_49383,N_49384,N_49385,N_49386,N_49387,N_49388,N_49389,N_49390,N_49391,N_49392,N_49393,N_49394,N_49395,N_49396,N_49397,N_49398,N_49399,N_49400,N_49401,N_49402,N_49403,N_49404,N_49405,N_49406,N_49407,N_49408,N_49409,N_49410,N_49411,N_49412,N_49413,N_49414,N_49415,N_49416,N_49417,N_49418,N_49419,N_49420,N_49421,N_49422,N_49423,N_49424,N_49425,N_49426,N_49427,N_49428,N_49429,N_49430,N_49431,N_49432,N_49433,N_49434,N_49435,N_49436,N_49437,N_49438,N_49439,N_49440,N_49441,N_49442,N_49443,N_49444,N_49445,N_49446,N_49447,N_49448,N_49449,N_49450,N_49451,N_49452,N_49453,N_49454,N_49455,N_49456,N_49457,N_49458,N_49459,N_49460,N_49461,N_49462,N_49463,N_49464,N_49465,N_49466,N_49467,N_49468,N_49469,N_49470,N_49471,N_49472,N_49473,N_49474,N_49475,N_49476,N_49477,N_49478,N_49479,N_49480,N_49481,N_49482,N_49483,N_49484,N_49485,N_49486,N_49487,N_49488,N_49489,N_49490,N_49491,N_49492,N_49493,N_49494,N_49495,N_49496,N_49497,N_49498,N_49499,N_49500,N_49501,N_49502,N_49503,N_49504,N_49505,N_49506,N_49507,N_49508,N_49509,N_49510,N_49511,N_49512,N_49513,N_49514,N_49515,N_49516,N_49517,N_49518,N_49519,N_49520,N_49521,N_49522,N_49523,N_49524,N_49525,N_49526,N_49527,N_49528,N_49529,N_49530,N_49531,N_49532,N_49533,N_49534,N_49535,N_49536,N_49537,N_49538,N_49539,N_49540,N_49541,N_49542,N_49543,N_49544,N_49545,N_49546,N_49547,N_49548,N_49549,N_49550,N_49551,N_49552,N_49553,N_49554,N_49555,N_49556,N_49557,N_49558,N_49559,N_49560,N_49561,N_49562,N_49563,N_49564,N_49565,N_49566,N_49567,N_49568,N_49569,N_49570,N_49571,N_49572,N_49573,N_49574,N_49575,N_49576,N_49577,N_49578,N_49579,N_49580,N_49581,N_49582,N_49583,N_49584,N_49585,N_49586,N_49587,N_49588,N_49589,N_49590,N_49591,N_49592,N_49593,N_49594,N_49595,N_49596,N_49597,N_49598,N_49599,N_49600,N_49601,N_49602,N_49603,N_49604,N_49605,N_49606,N_49607,N_49608,N_49609,N_49610,N_49611,N_49612,N_49613,N_49614,N_49615,N_49616,N_49617,N_49618,N_49619,N_49620,N_49621,N_49622,N_49623,N_49624,N_49625,N_49626,N_49627,N_49628,N_49629,N_49630,N_49631,N_49632,N_49633,N_49634,N_49635,N_49636,N_49637,N_49638,N_49639,N_49640,N_49641,N_49642,N_49643,N_49644,N_49645,N_49646,N_49647,N_49648,N_49649,N_49650,N_49651,N_49652,N_49653,N_49654,N_49655,N_49656,N_49657,N_49658,N_49659,N_49660,N_49661,N_49662,N_49663,N_49664,N_49665,N_49666,N_49667,N_49668,N_49669,N_49670,N_49671,N_49672,N_49673,N_49674,N_49675,N_49676,N_49677,N_49678,N_49679,N_49680,N_49681,N_49682,N_49683,N_49684,N_49685,N_49686,N_49687,N_49688,N_49689,N_49690,N_49691,N_49692,N_49693,N_49694,N_49695,N_49696,N_49697,N_49698,N_49699,N_49700,N_49701,N_49702,N_49703,N_49704,N_49705,N_49706,N_49707,N_49708,N_49709,N_49710,N_49711,N_49712,N_49713,N_49714,N_49715,N_49716,N_49717,N_49718,N_49719,N_49720,N_49721,N_49722,N_49723,N_49724,N_49725,N_49726,N_49727,N_49728,N_49729,N_49730,N_49731,N_49732,N_49733,N_49734,N_49735,N_49736,N_49737,N_49738,N_49739,N_49740,N_49741,N_49742,N_49743,N_49744,N_49745,N_49746,N_49747,N_49748,N_49749,N_49750,N_49751,N_49752,N_49753,N_49754,N_49755,N_49756,N_49757,N_49758,N_49759,N_49760,N_49761,N_49762,N_49763,N_49764,N_49765,N_49766,N_49767,N_49768,N_49769,N_49770,N_49771,N_49772,N_49773,N_49774,N_49775,N_49776,N_49777,N_49778,N_49779,N_49780,N_49781,N_49782,N_49783,N_49784,N_49785,N_49786,N_49787,N_49788,N_49789,N_49790,N_49791,N_49792,N_49793,N_49794,N_49795,N_49796,N_49797,N_49798,N_49799,N_49800,N_49801,N_49802,N_49803,N_49804,N_49805,N_49806,N_49807,N_49808,N_49809,N_49810,N_49811,N_49812,N_49813,N_49814,N_49815,N_49816,N_49817,N_49818,N_49819,N_49820,N_49821,N_49822,N_49823,N_49824,N_49825,N_49826,N_49827,N_49828,N_49829,N_49830,N_49831,N_49832,N_49833,N_49834,N_49835,N_49836,N_49837,N_49838,N_49839,N_49840,N_49841,N_49842,N_49843,N_49844,N_49845,N_49846,N_49847,N_49848,N_49849,N_49850,N_49851,N_49852,N_49853,N_49854,N_49855,N_49856,N_49857,N_49858,N_49859,N_49860,N_49861,N_49862,N_49863,N_49864,N_49865,N_49866,N_49867,N_49868,N_49869,N_49870,N_49871,N_49872,N_49873,N_49874,N_49875,N_49876,N_49877,N_49878,N_49879,N_49880,N_49881,N_49882,N_49883,N_49884,N_49885,N_49886,N_49887,N_49888,N_49889,N_49890,N_49891,N_49892,N_49893,N_49894,N_49895,N_49896,N_49897,N_49898,N_49899,N_49900,N_49901,N_49902,N_49903,N_49904,N_49905,N_49906,N_49907,N_49908,N_49909,N_49910,N_49911,N_49912,N_49913,N_49914,N_49915,N_49916,N_49917,N_49918,N_49919,N_49920,N_49921,N_49922,N_49923,N_49924,N_49925,N_49926,N_49927,N_49928,N_49929,N_49930,N_49931,N_49932,N_49933,N_49934,N_49935,N_49936,N_49937,N_49938,N_49939,N_49940,N_49941,N_49942,N_49943,N_49944,N_49945,N_49946,N_49947,N_49948,N_49949,N_49950,N_49951,N_49952,N_49953,N_49954,N_49955,N_49956,N_49957,N_49958,N_49959,N_49960,N_49961,N_49962,N_49963,N_49964,N_49965,N_49966,N_49967,N_49968,N_49969,N_49970,N_49971,N_49972,N_49973,N_49974,N_49975,N_49976,N_49977,N_49978,N_49979,N_49980,N_49981,N_49982,N_49983,N_49984,N_49985,N_49986,N_49987,N_49988,N_49989,N_49990,N_49991,N_49992,N_49993,N_49994,N_49995,N_49996,N_49997,N_49998,N_49999;
and U0 (N_0,In_4185,In_2968);
or U1 (N_1,In_724,In_459);
nor U2 (N_2,In_2460,In_2953);
or U3 (N_3,In_3015,In_615);
nand U4 (N_4,In_403,In_3656);
nor U5 (N_5,In_3781,In_4632);
and U6 (N_6,In_984,In_1941);
nand U7 (N_7,In_2045,In_2513);
and U8 (N_8,In_2334,In_1580);
and U9 (N_9,In_4746,In_4515);
xnor U10 (N_10,In_3988,In_460);
or U11 (N_11,In_4701,In_1294);
xnor U12 (N_12,In_3976,In_3624);
or U13 (N_13,In_2634,In_4647);
nor U14 (N_14,In_1692,In_1991);
xor U15 (N_15,In_4600,In_3148);
and U16 (N_16,In_2618,In_3554);
nor U17 (N_17,In_2866,In_256);
xor U18 (N_18,In_3128,In_4865);
and U19 (N_19,In_4931,In_1851);
xnor U20 (N_20,In_3182,In_3357);
nor U21 (N_21,In_2889,In_660);
and U22 (N_22,In_1940,In_827);
nor U23 (N_23,In_3707,In_423);
nor U24 (N_24,In_1373,In_4445);
nor U25 (N_25,In_2369,In_1368);
nor U26 (N_26,In_2496,In_174);
and U27 (N_27,In_2498,In_1952);
nand U28 (N_28,In_4683,In_1737);
or U29 (N_29,In_364,In_1367);
or U30 (N_30,In_2570,In_4689);
nand U31 (N_31,In_539,In_437);
nor U32 (N_32,In_4012,In_1839);
nor U33 (N_33,In_4978,In_1116);
xnor U34 (N_34,In_2022,In_2550);
nor U35 (N_35,In_2954,In_156);
xnor U36 (N_36,In_3939,In_3219);
or U37 (N_37,In_3599,In_753);
and U38 (N_38,In_428,In_2907);
xor U39 (N_39,In_2972,In_2210);
nand U40 (N_40,In_2764,In_3441);
xor U41 (N_41,In_1127,In_166);
nand U42 (N_42,In_4203,In_3226);
or U43 (N_43,In_4700,In_1460);
xnor U44 (N_44,In_4707,In_508);
nor U45 (N_45,In_3870,In_2152);
nand U46 (N_46,In_2287,In_749);
xor U47 (N_47,In_3686,In_4432);
nor U48 (N_48,In_3388,In_783);
xor U49 (N_49,In_1789,In_34);
nor U50 (N_50,In_3542,In_2707);
and U51 (N_51,In_3437,In_3551);
nand U52 (N_52,In_1233,In_4208);
or U53 (N_53,In_1485,In_1240);
xor U54 (N_54,In_4688,In_3106);
or U55 (N_55,In_3984,In_348);
nand U56 (N_56,In_128,In_163);
nand U57 (N_57,In_4182,In_347);
nand U58 (N_58,In_3623,In_2259);
nand U59 (N_59,In_3242,In_2232);
nand U60 (N_60,In_439,In_4564);
and U61 (N_61,In_2184,In_932);
xor U62 (N_62,In_4528,In_1708);
nand U63 (N_63,In_4177,In_4684);
xnor U64 (N_64,In_3941,In_1497);
and U65 (N_65,In_2733,In_1750);
or U66 (N_66,In_1339,In_4811);
xor U67 (N_67,In_3125,In_3943);
and U68 (N_68,In_2816,In_1615);
or U69 (N_69,In_4205,In_1535);
nor U70 (N_70,In_612,In_4840);
nand U71 (N_71,In_1985,In_398);
nand U72 (N_72,In_414,In_297);
nand U73 (N_73,In_2857,In_4072);
xor U74 (N_74,In_4704,In_1584);
and U75 (N_75,In_4249,In_2731);
or U76 (N_76,In_4738,In_671);
xnor U77 (N_77,In_1515,In_3848);
xor U78 (N_78,In_3229,In_746);
nand U79 (N_79,In_3638,In_4856);
nor U80 (N_80,In_4215,In_4863);
or U81 (N_81,In_3466,In_1380);
or U82 (N_82,In_4385,In_3213);
nor U83 (N_83,In_2141,In_4725);
xnor U84 (N_84,In_2019,In_3833);
nor U85 (N_85,In_3865,In_4345);
nand U86 (N_86,In_421,In_3123);
xor U87 (N_87,In_2162,In_4122);
xnor U88 (N_88,In_4771,In_2047);
and U89 (N_89,In_4229,In_422);
xnor U90 (N_90,In_1138,In_2769);
or U91 (N_91,In_4923,In_3922);
xnor U92 (N_92,In_2678,In_828);
or U93 (N_93,In_3491,In_4278);
xor U94 (N_94,In_1014,In_602);
nor U95 (N_95,In_3626,In_4536);
nand U96 (N_96,In_2121,In_2712);
nand U97 (N_97,In_2868,In_2400);
nand U98 (N_98,In_3692,In_103);
nand U99 (N_99,In_3012,In_2796);
nor U100 (N_100,In_1434,In_583);
nor U101 (N_101,In_3897,In_4641);
nand U102 (N_102,In_3187,In_2831);
and U103 (N_103,In_4845,In_4464);
nand U104 (N_104,In_3379,In_3178);
and U105 (N_105,In_914,In_4286);
and U106 (N_106,In_3001,In_194);
or U107 (N_107,In_4498,In_4921);
nand U108 (N_108,In_1664,In_2684);
nand U109 (N_109,In_2113,In_3141);
and U110 (N_110,In_1933,In_2252);
xnor U111 (N_111,In_2685,In_4376);
nand U112 (N_112,In_1490,In_4189);
and U113 (N_113,In_2814,In_3817);
xor U114 (N_114,In_430,In_3749);
nor U115 (N_115,In_2066,In_3492);
and U116 (N_116,In_3728,In_1243);
xor U117 (N_117,In_807,In_4158);
nand U118 (N_118,In_3206,In_906);
xnor U119 (N_119,In_1528,In_779);
nor U120 (N_120,In_1844,In_3667);
xnor U121 (N_121,In_1634,In_186);
nor U122 (N_122,In_2027,In_3700);
nor U123 (N_123,In_2402,In_3470);
nor U124 (N_124,In_3025,In_418);
or U125 (N_125,In_112,In_3895);
or U126 (N_126,In_1854,In_164);
xnor U127 (N_127,In_3806,In_1140);
nand U128 (N_128,In_3612,In_1047);
or U129 (N_129,In_1922,In_406);
xor U130 (N_130,In_3344,In_4344);
xnor U131 (N_131,In_1308,In_4932);
nand U132 (N_132,In_3261,In_4724);
nor U133 (N_133,In_2134,In_1471);
nor U134 (N_134,In_4057,In_4369);
nand U135 (N_135,In_505,In_2671);
xor U136 (N_136,In_3006,In_4567);
xnor U137 (N_137,In_2319,In_4802);
and U138 (N_138,In_3854,In_744);
nor U139 (N_139,In_3300,In_2782);
or U140 (N_140,In_4956,In_4324);
xor U141 (N_141,In_4669,In_2625);
or U142 (N_142,In_3360,In_642);
and U143 (N_143,In_1147,In_3868);
nor U144 (N_144,In_4220,In_3037);
or U145 (N_145,In_3654,In_2490);
or U146 (N_146,In_2603,In_1075);
nand U147 (N_147,In_699,In_2263);
nand U148 (N_148,In_1421,In_1216);
nor U149 (N_149,In_3752,In_2269);
nand U150 (N_150,In_2414,In_2412);
and U151 (N_151,In_2147,In_159);
nor U152 (N_152,In_3113,In_4413);
nand U153 (N_153,In_1804,In_716);
or U154 (N_154,In_1365,In_1028);
nor U155 (N_155,In_4470,In_1377);
nand U156 (N_156,In_1801,In_4611);
nand U157 (N_157,In_4092,In_3999);
nand U158 (N_158,In_805,In_2331);
and U159 (N_159,In_2196,In_148);
and U160 (N_160,In_3812,In_647);
xnor U161 (N_161,In_4473,In_2254);
and U162 (N_162,In_2897,In_2051);
or U163 (N_163,In_4251,In_1561);
nand U164 (N_164,In_4965,In_1627);
nand U165 (N_165,In_3191,In_104);
nand U166 (N_166,In_3475,In_1565);
and U167 (N_167,In_2918,In_2621);
nor U168 (N_168,In_1224,In_4588);
xor U169 (N_169,In_443,In_1864);
nand U170 (N_170,In_538,In_2140);
nand U171 (N_171,In_84,In_2489);
and U172 (N_172,In_1836,In_20);
or U173 (N_173,In_54,In_2619);
nor U174 (N_174,In_489,In_1967);
or U175 (N_175,In_1694,In_482);
xnor U176 (N_176,In_494,In_1752);
xnor U177 (N_177,In_4101,In_2075);
xor U178 (N_178,In_1576,In_2574);
nand U179 (N_179,In_1180,In_2748);
nand U180 (N_180,In_132,In_1206);
or U181 (N_181,In_1329,In_1792);
nor U182 (N_182,In_4513,In_1472);
nand U183 (N_183,In_2710,In_2435);
nand U184 (N_184,In_2899,In_3056);
nand U185 (N_185,In_1374,In_1894);
nor U186 (N_186,In_2662,In_4420);
or U187 (N_187,In_4495,In_2393);
nand U188 (N_188,In_1437,In_576);
xnor U189 (N_189,In_574,In_2175);
and U190 (N_190,In_2370,In_763);
and U191 (N_191,In_4703,In_2491);
and U192 (N_192,In_1908,In_288);
or U193 (N_193,In_3019,In_4397);
or U194 (N_194,In_3851,In_1770);
and U195 (N_195,In_4407,In_2554);
or U196 (N_196,In_4361,In_4363);
or U197 (N_197,In_2193,In_215);
nor U198 (N_198,In_4099,In_973);
nor U199 (N_199,In_4633,In_2647);
nand U200 (N_200,In_4031,In_1262);
nor U201 (N_201,In_3741,In_3940);
nor U202 (N_202,In_455,In_3615);
xor U203 (N_203,In_1409,In_2220);
and U204 (N_204,In_227,In_449);
nand U205 (N_205,In_2026,In_1823);
nor U206 (N_206,In_4418,In_672);
nand U207 (N_207,In_1959,In_834);
xor U208 (N_208,In_4757,In_442);
nor U209 (N_209,In_1719,In_3232);
xor U210 (N_210,In_4793,In_361);
nand U211 (N_211,In_870,In_1977);
xnor U212 (N_212,In_704,In_2653);
and U213 (N_213,In_1614,In_4890);
nor U214 (N_214,In_2589,In_2841);
xnor U215 (N_215,In_2089,In_498);
nand U216 (N_216,In_120,In_1872);
nor U217 (N_217,In_1878,In_670);
nor U218 (N_218,In_2883,In_2119);
nand U219 (N_219,In_2326,In_1779);
and U220 (N_220,In_935,In_1379);
or U221 (N_221,In_526,In_2601);
nor U222 (N_222,In_1404,In_199);
and U223 (N_223,In_1364,In_3899);
nand U224 (N_224,In_4779,In_2573);
nand U225 (N_225,In_4997,In_654);
and U226 (N_226,In_734,In_3131);
and U227 (N_227,In_2273,In_4843);
nand U228 (N_228,In_4422,In_2327);
xnor U229 (N_229,In_2071,In_1623);
nand U230 (N_230,In_3644,In_1524);
nor U231 (N_231,In_3453,In_2955);
nor U232 (N_232,In_4283,In_3162);
nor U233 (N_233,In_3565,In_4850);
and U234 (N_234,In_295,In_2424);
and U235 (N_235,In_2768,In_4103);
and U236 (N_236,In_907,In_3152);
and U237 (N_237,In_2833,In_982);
or U238 (N_238,In_3507,In_1103);
xor U239 (N_239,In_3714,In_2068);
xnor U240 (N_240,In_519,In_393);
and U241 (N_241,In_3304,In_2276);
and U242 (N_242,In_441,In_335);
xor U243 (N_243,In_3456,In_1755);
nor U244 (N_244,In_3795,In_762);
nand U245 (N_245,In_3964,In_4770);
nor U246 (N_246,In_999,In_1514);
xor U247 (N_247,In_1414,In_444);
nor U248 (N_248,In_1451,In_930);
and U249 (N_249,In_3350,In_4673);
and U250 (N_250,In_629,In_3704);
xor U251 (N_251,In_3991,In_878);
and U252 (N_252,In_4062,In_2996);
xor U253 (N_253,In_456,In_1467);
xor U254 (N_254,In_4194,In_4810);
nand U255 (N_255,In_3282,In_2957);
nand U256 (N_256,In_1903,In_4783);
nor U257 (N_257,In_3007,In_2994);
xnor U258 (N_258,In_3605,In_1154);
nor U259 (N_259,In_1825,In_1884);
nor U260 (N_260,In_91,In_2317);
and U261 (N_261,In_1696,In_2668);
xnor U262 (N_262,In_1182,In_4058);
or U263 (N_263,In_3077,In_1678);
nor U264 (N_264,In_1793,In_1929);
nor U265 (N_265,In_1670,In_1137);
or U266 (N_266,In_980,In_176);
and U267 (N_267,In_369,In_2679);
nand U268 (N_268,In_302,In_170);
nor U269 (N_269,In_4957,In_2443);
nand U270 (N_270,In_3670,In_2239);
or U271 (N_271,In_185,In_3078);
and U272 (N_272,In_4225,In_4553);
nand U273 (N_273,In_946,In_44);
xnor U274 (N_274,In_3249,In_1122);
nand U275 (N_275,In_4264,In_2545);
or U276 (N_276,In_3035,In_2851);
nor U277 (N_277,In_2258,In_3495);
or U278 (N_278,In_693,In_1695);
and U279 (N_279,In_2484,In_2480);
or U280 (N_280,In_808,In_3850);
or U281 (N_281,In_2038,In_3591);
and U282 (N_282,In_960,In_2342);
nor U283 (N_283,In_1178,In_3387);
nor U284 (N_284,In_3169,In_3746);
and U285 (N_285,In_3032,In_3712);
and U286 (N_286,In_2368,In_1295);
nor U287 (N_287,In_820,In_3643);
xnor U288 (N_288,In_540,In_531);
or U289 (N_289,In_4670,In_1229);
xnor U290 (N_290,In_3235,In_3133);
xnor U291 (N_291,In_2860,In_184);
or U292 (N_292,In_4410,In_899);
xnor U293 (N_293,In_4444,In_1263);
xnor U294 (N_294,In_2818,In_2632);
or U295 (N_295,In_651,In_511);
or U296 (N_296,In_1051,In_2219);
or U297 (N_297,In_2810,In_4557);
and U298 (N_298,In_240,In_995);
nand U299 (N_299,In_3585,In_2537);
xor U300 (N_300,In_445,In_1799);
nand U301 (N_301,In_2927,In_4254);
and U302 (N_302,In_1305,In_2962);
xnor U303 (N_303,In_1320,In_547);
nor U304 (N_304,In_1860,In_2770);
or U305 (N_305,In_1539,In_1759);
or U306 (N_306,In_3651,In_4574);
xor U307 (N_307,In_1435,In_835);
nor U308 (N_308,In_3188,In_4467);
nand U309 (N_309,In_2846,In_1119);
nor U310 (N_310,In_3708,In_3950);
nor U311 (N_311,In_3804,In_3505);
xor U312 (N_312,In_909,In_3655);
or U313 (N_313,In_126,In_3693);
nor U314 (N_314,In_3675,In_1077);
and U315 (N_315,In_4443,In_1598);
and U316 (N_316,In_96,In_2813);
nor U317 (N_317,In_4596,In_4181);
nor U318 (N_318,In_3230,In_4535);
or U319 (N_319,In_3218,In_3183);
or U320 (N_320,In_56,In_3364);
xnor U321 (N_321,In_3333,In_1310);
nor U322 (N_322,In_1301,In_688);
or U323 (N_323,In_429,In_3535);
nand U324 (N_324,In_2997,In_4760);
and U325 (N_325,In_4450,In_3962);
and U326 (N_326,In_1344,In_3457);
and U327 (N_327,In_1474,In_3005);
or U328 (N_328,In_1511,In_1470);
nor U329 (N_329,In_2881,In_2898);
nor U330 (N_330,In_1403,In_4869);
xor U331 (N_331,In_3914,In_1742);
and U332 (N_332,In_1441,In_1660);
or U333 (N_333,In_1275,In_4506);
xnor U334 (N_334,In_4942,In_3260);
nor U335 (N_335,In_2516,In_789);
or U336 (N_336,In_2624,In_4726);
nor U337 (N_337,In_3496,In_2627);
nor U338 (N_338,In_1297,In_4275);
nand U339 (N_339,In_1427,In_1601);
nor U340 (N_340,In_1955,In_4392);
nor U341 (N_341,In_4824,In_462);
nand U342 (N_342,In_849,In_61);
or U343 (N_343,In_2974,In_2885);
or U344 (N_344,In_992,In_3657);
and U345 (N_345,In_2434,In_3292);
or U346 (N_346,In_1384,In_4402);
nand U347 (N_347,In_4690,In_2597);
xor U348 (N_348,In_1285,In_2576);
nor U349 (N_349,In_3144,In_3583);
and U350 (N_350,In_3010,In_4077);
nand U351 (N_351,In_4301,In_1251);
xnor U352 (N_352,In_2155,In_3061);
nor U353 (N_353,In_4417,In_1444);
or U354 (N_354,In_4984,In_2674);
and U355 (N_355,In_1419,In_507);
or U356 (N_356,In_3761,In_2947);
xor U357 (N_357,In_4065,In_2329);
and U358 (N_358,In_2541,In_4868);
and U359 (N_359,In_1984,In_2732);
and U360 (N_360,In_719,In_4538);
xnor U361 (N_361,In_3805,In_3444);
nor U362 (N_362,In_345,In_1768);
and U363 (N_363,In_273,In_2064);
nand U364 (N_364,In_1287,In_1070);
and U365 (N_365,In_2111,In_4591);
and U366 (N_366,In_69,In_1944);
nor U367 (N_367,In_1817,In_1537);
xor U368 (N_368,In_4861,In_2514);
xnor U369 (N_369,In_3823,In_3048);
and U370 (N_370,In_720,In_2893);
and U371 (N_371,In_892,In_3103);
xor U372 (N_372,In_1311,In_4149);
or U373 (N_373,In_1304,In_1389);
nor U374 (N_374,In_4826,In_2950);
or U375 (N_375,In_1350,In_4728);
nor U376 (N_376,In_1832,In_1267);
xor U377 (N_377,In_3070,In_3951);
nand U378 (N_378,In_3872,In_3190);
nor U379 (N_379,In_4736,In_3952);
nand U380 (N_380,In_2408,In_291);
xnor U381 (N_381,In_2998,In_3278);
nor U382 (N_382,In_614,In_424);
xnor U383 (N_383,In_4960,In_937);
or U384 (N_384,In_178,In_3954);
xor U385 (N_385,In_200,In_2804);
and U386 (N_386,In_3995,In_2316);
and U387 (N_387,In_1885,In_1754);
nand U388 (N_388,In_1290,In_31);
nand U389 (N_389,In_2224,In_3446);
and U390 (N_390,In_3448,In_4814);
nor U391 (N_391,In_4572,In_2355);
xnor U392 (N_392,In_1084,In_1299);
nand U393 (N_393,In_3729,In_4291);
nand U394 (N_394,In_1574,In_4664);
or U395 (N_395,In_79,In_1778);
nor U396 (N_396,In_2696,In_4339);
xor U397 (N_397,In_1605,In_3987);
xor U398 (N_398,In_2808,In_3073);
and U399 (N_399,In_64,In_1230);
nand U400 (N_400,In_2956,In_635);
and U401 (N_401,In_2807,In_3794);
xor U402 (N_402,In_1982,In_4035);
nor U403 (N_403,In_4382,In_4516);
nor U404 (N_404,In_4132,In_4964);
and U405 (N_405,In_1644,In_945);
nor U406 (N_406,In_2803,In_709);
and U407 (N_407,In_142,In_3632);
or U408 (N_408,In_1087,In_2633);
nor U409 (N_409,In_2659,In_2345);
nand U410 (N_410,In_2636,In_4328);
nor U411 (N_411,In_3407,In_1276);
xor U412 (N_412,In_4549,In_1689);
or U413 (N_413,In_4243,In_3273);
and U414 (N_414,In_2418,In_4457);
nor U415 (N_415,In_3210,In_4579);
or U416 (N_416,In_1433,In_1432);
xor U417 (N_417,In_2381,In_4815);
xnor U418 (N_418,In_4419,In_131);
and U419 (N_419,In_29,In_1741);
and U420 (N_420,In_543,In_3297);
nor U421 (N_421,In_845,In_4927);
xnor U422 (N_422,In_1966,In_2250);
nand U423 (N_423,In_3465,In_1248);
or U424 (N_424,In_2291,In_3135);
xnor U425 (N_425,In_4014,In_1082);
nor U426 (N_426,In_3394,In_4082);
xnor U427 (N_427,In_4095,In_1930);
and U428 (N_428,In_2308,In_3140);
or U429 (N_429,In_4855,In_1499);
nand U430 (N_430,In_2971,In_2604);
and U431 (N_431,In_3658,In_3181);
or U432 (N_432,In_1593,In_2153);
or U433 (N_433,In_4431,In_4166);
or U434 (N_434,In_3075,In_1237);
nor U435 (N_435,In_3620,In_3497);
and U436 (N_436,In_4270,In_2073);
nor U437 (N_437,In_3842,In_3563);
xnor U438 (N_438,In_1239,In_4755);
nand U439 (N_439,In_384,In_448);
and U440 (N_440,In_708,In_2858);
nor U441 (N_441,In_3532,In_3919);
xnor U442 (N_442,In_2044,In_4556);
nand U443 (N_443,In_4234,In_2900);
nor U444 (N_444,In_366,In_28);
nor U445 (N_445,In_4847,In_4034);
nand U446 (N_446,In_375,In_1023);
nor U447 (N_447,In_410,In_2970);
and U448 (N_448,In_1926,In_4491);
and U449 (N_449,In_242,In_3502);
xnor U450 (N_450,In_3664,In_4232);
or U451 (N_451,In_4066,In_817);
and U452 (N_452,In_1091,In_263);
xor U453 (N_453,In_3485,In_2669);
nand U454 (N_454,In_1193,In_3362);
or U455 (N_455,In_864,In_3322);
or U456 (N_456,In_1585,In_1699);
xnor U457 (N_457,In_515,In_4844);
or U458 (N_458,In_898,In_451);
nor U459 (N_459,In_210,In_4590);
nor U460 (N_460,In_1181,In_3861);
nand U461 (N_461,In_745,In_1079);
xnor U462 (N_462,In_1645,In_1351);
xnor U463 (N_463,In_4317,In_2020);
nor U464 (N_464,In_3438,In_90);
nor U465 (N_465,In_2060,In_2741);
or U466 (N_466,In_4562,In_490);
xnor U467 (N_467,In_3528,In_3262);
nand U468 (N_468,In_3713,In_4056);
xnor U469 (N_469,In_2493,In_1993);
and U470 (N_470,In_3004,In_3736);
and U471 (N_471,In_4086,In_4722);
nor U472 (N_472,In_3718,In_1066);
xnor U473 (N_473,In_2778,In_4304);
or U474 (N_474,In_2447,In_2419);
xor U475 (N_475,In_791,In_1402);
nor U476 (N_476,In_4052,In_2407);
xor U477 (N_477,In_3594,In_1508);
nor U478 (N_478,In_1292,In_1577);
xor U479 (N_479,In_3246,In_4380);
xnor U480 (N_480,In_4827,In_3556);
nor U481 (N_481,In_1949,In_1717);
and U482 (N_482,In_3404,In_1709);
xor U483 (N_483,In_136,In_2088);
and U484 (N_484,In_3942,In_4872);
xnor U485 (N_485,In_117,In_3482);
and U486 (N_486,In_1981,In_1022);
and U487 (N_487,In_4218,In_4260);
xnor U488 (N_488,In_4860,In_3617);
xnor U489 (N_489,In_4262,In_3710);
xnor U490 (N_490,In_601,In_4348);
or U491 (N_491,In_4616,In_3808);
or U492 (N_492,In_1814,In_1834);
nand U493 (N_493,In_3701,In_1527);
or U494 (N_494,In_2783,In_4871);
or U495 (N_495,In_4873,In_471);
and U496 (N_496,In_3649,In_2445);
or U497 (N_497,In_885,In_739);
nor U498 (N_498,In_2297,In_3274);
and U499 (N_499,In_4112,In_2660);
and U500 (N_500,In_2018,In_50);
nand U501 (N_501,In_2450,In_3602);
or U502 (N_502,In_4575,In_2914);
nand U503 (N_503,In_4250,In_4028);
xor U504 (N_504,In_532,In_1064);
or U505 (N_505,In_1357,In_3562);
or U506 (N_506,In_2122,In_3857);
nand U507 (N_507,In_3824,In_3014);
xor U508 (N_508,In_4364,In_1667);
or U509 (N_509,In_3399,In_2951);
or U510 (N_510,In_1995,In_931);
xor U511 (N_511,In_4175,In_432);
nand U512 (N_512,In_4321,In_4106);
and U513 (N_513,In_1277,In_2840);
nand U514 (N_514,In_4456,In_3918);
and U515 (N_515,In_360,In_2495);
and U516 (N_516,In_4682,In_3568);
or U517 (N_517,In_2178,In_683);
xor U518 (N_518,In_580,In_3199);
nand U519 (N_519,In_3411,In_81);
nor U520 (N_520,In_1706,In_188);
and U521 (N_521,In_4825,In_2622);
nand U522 (N_522,In_4258,In_2417);
nor U523 (N_523,In_2924,In_3405);
and U524 (N_524,In_1319,In_2195);
nor U525 (N_525,In_1252,In_3785);
nor U526 (N_526,In_3621,In_801);
and U527 (N_527,In_294,In_2845);
or U528 (N_528,In_32,In_607);
nand U529 (N_529,In_2440,In_3880);
xnor U530 (N_530,In_4210,In_3307);
and U531 (N_531,In_3454,In_3782);
and U532 (N_532,In_2009,In_2231);
and U533 (N_533,In_21,In_963);
nand U534 (N_534,In_66,In_3247);
nor U535 (N_535,In_1716,In_1788);
xnor U536 (N_536,In_67,In_4206);
xnor U537 (N_537,In_1431,In_3634);
nor U538 (N_538,In_2582,In_2166);
or U539 (N_539,In_3050,In_2307);
xor U540 (N_540,In_1591,In_1938);
nor U541 (N_541,In_998,In_4652);
nor U542 (N_542,In_2098,In_1613);
and U543 (N_543,In_4226,In_775);
or U544 (N_544,In_3347,In_4754);
xor U545 (N_545,In_2992,In_477);
nor U546 (N_546,In_3208,In_324);
nor U547 (N_547,In_1543,In_1774);
xnor U548 (N_548,In_1776,In_219);
nor U549 (N_549,In_401,In_3661);
nand U550 (N_550,In_3154,In_2729);
or U551 (N_551,In_4130,In_2799);
or U552 (N_552,In_180,In_2004);
xor U553 (N_553,In_3236,In_3474);
nor U554 (N_554,In_3439,In_1571);
nand U555 (N_555,In_2535,In_4367);
nor U556 (N_556,In_1190,In_4298);
nand U557 (N_557,In_1187,In_157);
and U558 (N_558,In_1225,In_2301);
nor U559 (N_559,In_4809,In_1009);
and U560 (N_560,In_2335,In_2097);
nor U561 (N_561,In_4638,In_4566);
nor U562 (N_562,In_1669,In_4654);
or U563 (N_563,In_1896,In_3600);
and U564 (N_564,In_664,In_3030);
xor U565 (N_565,In_4715,In_1196);
or U566 (N_566,In_3849,In_4714);
or U567 (N_567,In_4667,In_3443);
and U568 (N_568,In_4613,In_1124);
or U569 (N_569,In_1236,In_3088);
nor U570 (N_570,In_3847,In_1383);
nand U571 (N_571,In_4004,In_1712);
xnor U572 (N_572,In_1255,In_2934);
nand U573 (N_573,In_1390,In_4666);
and U574 (N_574,In_961,In_2534);
and U575 (N_575,In_3510,In_2766);
and U576 (N_576,In_652,In_3639);
nand U577 (N_577,In_431,In_4522);
nand U578 (N_578,In_2595,In_4316);
and U579 (N_579,In_2354,In_4539);
xnor U580 (N_580,In_2203,In_2087);
xor U581 (N_581,In_3660,In_3192);
xor U582 (N_582,In_4263,In_1999);
nand U583 (N_583,In_773,In_3319);
nand U584 (N_584,In_1874,In_4903);
xor U585 (N_585,In_3059,In_1200);
or U586 (N_586,In_1399,In_1279);
or U587 (N_587,In_3908,In_3317);
xor U588 (N_588,In_4698,In_4318);
or U589 (N_589,In_59,In_1650);
nand U590 (N_590,In_4389,In_530);
or U591 (N_591,In_3267,In_4694);
nor U592 (N_592,In_3095,In_2518);
nor U593 (N_593,In_705,In_267);
or U594 (N_594,In_2965,In_4374);
nor U595 (N_595,In_465,In_1906);
or U596 (N_596,In_3312,In_4558);
or U597 (N_597,In_593,In_1821);
and U598 (N_598,In_2609,In_2906);
nand U599 (N_599,In_3486,In_3925);
nand U600 (N_600,In_4151,In_1386);
or U601 (N_601,In_4357,In_2118);
nor U602 (N_602,In_556,In_389);
nor U603 (N_603,In_1979,In_4915);
nor U604 (N_604,In_662,In_3888);
xnor U605 (N_605,In_4492,In_2980);
and U606 (N_606,In_2366,In_1141);
xor U607 (N_607,In_611,In_3597);
nand U608 (N_608,In_4646,In_3250);
xnor U609 (N_609,In_2229,In_1078);
and U610 (N_610,In_4105,In_3356);
nand U611 (N_611,In_4607,In_2142);
xor U612 (N_612,In_3549,In_528);
or U613 (N_613,In_1641,In_4995);
or U614 (N_614,In_4463,In_3220);
nand U615 (N_615,In_2932,In_3923);
nor U616 (N_616,In_119,In_3687);
xor U617 (N_617,In_3743,In_1455);
nor U618 (N_618,In_3796,In_3158);
and U619 (N_619,In_208,In_1923);
nand U620 (N_620,In_1133,In_1980);
nor U621 (N_621,In_1757,In_3009);
nor U622 (N_622,In_3674,In_1815);
nand U623 (N_623,In_2110,In_1881);
nor U624 (N_624,In_3780,In_182);
xnor U625 (N_625,In_454,In_1965);
or U626 (N_626,In_3207,In_4525);
nand U627 (N_627,In_1232,In_752);
xnor U628 (N_628,In_4716,In_3268);
nand U629 (N_629,In_4365,In_1188);
nor U630 (N_630,In_1636,In_1157);
and U631 (N_631,In_954,In_3266);
nor U632 (N_632,In_3832,In_2864);
or U633 (N_633,In_3305,In_4113);
xnor U634 (N_634,In_3682,In_3846);
and U635 (N_635,In_391,In_3935);
nand U636 (N_636,In_1487,In_3256);
nor U637 (N_637,In_4547,In_2515);
and U638 (N_638,In_3783,In_3699);
nor U639 (N_639,In_1076,In_4313);
nor U640 (N_640,In_2438,In_2967);
nand U641 (N_641,In_3912,In_3516);
nor U642 (N_642,In_2284,In_204);
xnor U643 (N_643,In_3500,In_841);
or U644 (N_644,In_3552,In_1197);
xor U645 (N_645,In_1827,In_296);
and U646 (N_646,In_3802,In_4299);
or U647 (N_647,In_3413,In_3931);
xnor U648 (N_648,In_1638,In_1665);
or U649 (N_649,In_1686,In_2244);
and U650 (N_650,In_2454,In_2471);
nand U651 (N_651,In_2077,In_2099);
xor U652 (N_652,In_3244,In_2532);
or U653 (N_653,In_2048,In_2538);
xor U654 (N_654,In_1573,In_731);
or U655 (N_655,In_3094,In_903);
and U656 (N_656,In_1207,In_1622);
or U657 (N_657,In_2835,In_632);
xnor U658 (N_658,In_3299,In_503);
and U659 (N_659,In_4453,In_4461);
and U660 (N_660,In_3825,In_3117);
xor U661 (N_661,In_3784,In_2012);
nand U662 (N_662,In_799,In_4628);
nand U663 (N_663,In_95,In_1226);
nand U664 (N_664,In_4595,In_3767);
xnor U665 (N_665,In_3204,In_3598);
or U666 (N_666,In_169,In_2984);
nor U667 (N_667,In_1813,In_4093);
xnor U668 (N_668,In_3170,In_1054);
and U669 (N_669,In_3313,In_4179);
nor U670 (N_670,In_1452,In_481);
or U671 (N_671,In_75,In_2630);
nand U672 (N_672,In_3538,In_4379);
and U673 (N_673,In_3136,In_1408);
xor U674 (N_674,In_2256,In_3519);
nor U675 (N_675,In_856,In_4213);
and U676 (N_676,In_1041,In_4157);
nor U677 (N_677,In_4016,In_3402);
or U678 (N_678,In_1246,In_4900);
xnor U679 (N_679,In_2006,In_4980);
nand U680 (N_680,In_3198,In_1125);
nand U681 (N_681,In_917,In_1385);
or U682 (N_682,In_1596,In_2823);
and U683 (N_683,In_4817,In_1974);
xor U684 (N_684,In_1529,In_2929);
xor U685 (N_685,In_1089,In_4289);
nand U686 (N_686,In_2880,In_3284);
or U687 (N_687,In_3000,In_1996);
xor U688 (N_688,In_2233,In_1810);
xor U689 (N_689,In_49,In_2116);
nand U690 (N_690,In_2797,In_1067);
or U691 (N_691,In_4411,In_1234);
nand U692 (N_692,In_3747,In_4765);
xor U693 (N_693,In_4240,In_2509);
nor U694 (N_694,In_3938,In_93);
xor U695 (N_695,In_3715,In_774);
and U696 (N_696,In_812,In_1599);
nor U697 (N_697,In_1477,In_4368);
nor U698 (N_698,In_3209,In_702);
nor U699 (N_699,In_2266,In_341);
xnor U700 (N_700,In_4929,In_1951);
nor U701 (N_701,In_4474,In_546);
or U702 (N_702,In_1440,In_4776);
or U703 (N_703,In_1146,In_784);
nor U704 (N_704,In_3534,In_3731);
xnor U705 (N_705,In_2035,In_553);
nor U706 (N_706,In_223,In_1521);
nor U707 (N_707,In_474,In_4383);
and U708 (N_708,In_3211,In_3757);
nand U709 (N_709,In_2451,In_3372);
nor U710 (N_710,In_4829,In_1505);
xor U711 (N_711,In_1840,In_2780);
nand U712 (N_712,In_2754,In_1570);
xor U713 (N_713,In_3487,In_3316);
or U714 (N_714,In_694,In_2693);
nor U715 (N_715,In_1506,In_2937);
and U716 (N_716,In_1274,In_1826);
nand U717 (N_717,In_383,In_3156);
nand U718 (N_718,In_2999,In_2942);
and U719 (N_719,In_1562,In_3359);
or U720 (N_720,In_1714,In_2543);
or U721 (N_721,In_4412,In_2396);
or U722 (N_722,In_1978,In_4883);
nand U723 (N_723,In_1381,In_1866);
xor U724 (N_724,In_2727,In_3877);
nand U725 (N_725,In_191,In_312);
nand U726 (N_726,In_2964,In_3459);
and U727 (N_727,In_643,In_2930);
or U728 (N_728,In_3499,In_728);
and U729 (N_729,In_2372,In_2240);
and U730 (N_730,In_4261,In_475);
or U731 (N_731,In_926,In_122);
and U732 (N_732,In_304,In_3341);
xnor U733 (N_733,In_1626,In_3225);
or U734 (N_734,In_4561,In_2165);
nor U735 (N_735,In_308,In_1002);
nor U736 (N_736,In_910,In_3124);
xnor U737 (N_737,In_3115,In_3238);
nand U738 (N_738,In_2548,In_4603);
nor U739 (N_739,In_4405,In_4375);
xnor U740 (N_740,In_129,In_3034);
nand U741 (N_741,In_1865,In_370);
or U742 (N_742,In_840,In_1892);
or U743 (N_743,In_1703,In_2430);
or U744 (N_744,In_4452,In_2170);
xor U745 (N_745,In_1803,In_1135);
nand U746 (N_746,In_3455,In_1671);
nor U747 (N_747,In_55,In_3468);
nor U748 (N_748,In_276,In_3258);
nand U749 (N_749,In_4565,In_4195);
nand U750 (N_750,In_3331,In_2616);
nand U751 (N_751,In_3038,In_1331);
nor U752 (N_752,In_3911,In_4469);
nand U753 (N_753,In_2485,In_3288);
and U754 (N_754,In_53,In_281);
xor U755 (N_755,In_4626,In_1588);
nor U756 (N_756,In_3290,In_4437);
or U757 (N_757,In_747,In_838);
xor U758 (N_758,In_4568,In_3546);
nand U759 (N_759,In_3668,In_4630);
xnor U760 (N_760,In_4734,In_42);
or U761 (N_761,In_4747,In_2935);
nand U762 (N_762,In_1740,In_2631);
and U763 (N_763,In_1007,In_4838);
and U764 (N_764,In_1126,In_4610);
or U765 (N_765,In_4390,In_4219);
and U766 (N_766,In_1540,In_1936);
nor U767 (N_767,In_1453,In_3921);
xor U768 (N_768,In_2686,In_6);
xor U769 (N_769,In_3186,In_4388);
nor U770 (N_770,In_4818,In_1557);
or U771 (N_771,In_2021,In_582);
or U772 (N_772,In_3361,In_814);
and U773 (N_773,In_4172,In_1450);
and U774 (N_774,In_4472,In_4429);
and U775 (N_775,In_1052,In_2245);
and U776 (N_776,In_2730,In_1059);
and U777 (N_777,In_2101,In_750);
nor U778 (N_778,In_894,In_3927);
nand U779 (N_779,In_4239,In_4801);
xnor U780 (N_780,In_3285,In_2805);
or U781 (N_781,In_3759,In_4544);
nor U782 (N_782,In_1131,In_23);
or U783 (N_783,In_3543,In_3397);
nand U784 (N_784,In_2221,In_1044);
or U785 (N_785,In_4191,In_4268);
or U786 (N_786,In_1852,In_320);
xnor U787 (N_787,In_2293,In_3679);
or U788 (N_788,In_1211,In_1532);
and U789 (N_789,In_1531,In_2457);
or U790 (N_790,In_63,In_3122);
and U791 (N_791,In_1478,In_1791);
or U792 (N_792,In_1438,In_1083);
nor U793 (N_793,In_3318,In_327);
nand U794 (N_794,In_3685,In_292);
and U795 (N_795,In_1278,In_2677);
and U796 (N_796,In_4764,In_2560);
nor U797 (N_797,In_2249,In_3092);
xnor U798 (N_798,In_1118,In_2681);
or U799 (N_799,In_4858,In_4233);
nor U800 (N_800,In_3610,In_1533);
nor U801 (N_801,In_510,In_748);
nor U802 (N_802,In_646,In_2201);
nor U803 (N_803,In_1786,In_4920);
and U804 (N_804,In_560,In_1681);
nand U805 (N_805,In_1958,In_1323);
nor U806 (N_806,In_4663,In_4303);
or U807 (N_807,In_4914,In_3147);
xor U808 (N_808,In_3120,In_4851);
xnor U809 (N_809,In_2644,In_4599);
nor U810 (N_810,In_2579,In_2709);
nor U811 (N_811,In_3325,In_3560);
nand U812 (N_812,In_4834,In_4201);
xor U813 (N_813,In_2718,In_951);
or U814 (N_814,In_653,In_1683);
nor U815 (N_815,In_4107,In_2373);
and U816 (N_816,In_550,In_332);
nand U817 (N_817,In_2065,In_1861);
nand U818 (N_818,In_2349,In_3368);
nand U819 (N_819,In_2894,In_3901);
and U820 (N_820,In_2901,In_4394);
and U821 (N_821,In_4211,In_1491);
xnor U822 (N_822,In_4852,In_4819);
or U823 (N_823,In_2013,In_3882);
and U824 (N_824,In_4656,In_1479);
nand U825 (N_825,In_1203,In_3852);
or U826 (N_826,In_1018,In_252);
xor U827 (N_827,In_4737,In_162);
or U828 (N_828,In_3677,In_983);
nand U829 (N_829,In_730,In_1167);
or U830 (N_830,In_4999,In_1546);
nand U831 (N_831,In_4938,In_2699);
nand U832 (N_832,In_2666,In_190);
nand U833 (N_833,In_2452,In_3074);
and U834 (N_834,In_4297,In_1603);
nor U835 (N_835,In_1218,In_3813);
xnor U836 (N_836,In_4735,In_3253);
xnor U837 (N_837,In_1567,In_2304);
nor U838 (N_838,In_803,In_446);
nand U839 (N_839,In_3303,In_1563);
xnor U840 (N_840,In_1202,In_3381);
nand U841 (N_841,In_1300,In_1816);
nand U842 (N_842,In_4416,In_957);
or U843 (N_843,In_2298,In_3172);
nand U844 (N_844,In_101,In_908);
or U845 (N_845,In_16,In_1777);
nor U846 (N_846,In_663,In_1322);
or U847 (N_847,In_3689,In_3650);
and U848 (N_848,In_1281,In_1268);
nor U849 (N_849,In_3203,In_1484);
nand U850 (N_850,In_2983,In_4503);
xor U851 (N_851,In_86,In_108);
and U852 (N_852,In_913,In_2795);
nand U853 (N_853,In_4499,In_4745);
nor U854 (N_854,In_301,In_4127);
xnor U855 (N_855,In_3257,In_1284);
or U856 (N_856,In_4952,In_2849);
nor U857 (N_857,In_4614,In_2197);
xnor U858 (N_858,In_3,In_2076);
or U859 (N_859,In_4391,In_4448);
and U860 (N_860,In_1191,In_4081);
nor U861 (N_861,In_883,In_4050);
xnor U862 (N_862,In_1199,In_977);
nor U863 (N_863,In_516,In_4427);
and U864 (N_864,In_485,In_4622);
or U865 (N_865,In_2157,In_2740);
nand U866 (N_866,In_3047,In_3339);
and U867 (N_867,In_4078,In_2074);
and U868 (N_868,In_346,In_4161);
nor U869 (N_869,In_2989,In_3928);
nand U870 (N_870,In_3862,In_3269);
and U871 (N_871,In_2641,In_4257);
and U872 (N_872,In_3440,In_4486);
and U873 (N_873,In_4803,In_1725);
xnor U874 (N_874,In_1169,In_1021);
nor U875 (N_875,In_4706,In_2150);
or U876 (N_876,In_2188,In_1010);
xor U877 (N_877,In_524,In_4878);
and U878 (N_878,In_665,In_2854);
nor U879 (N_879,In_2590,In_216);
xor U880 (N_880,In_1504,In_2665);
xnor U881 (N_881,In_4337,In_822);
and U882 (N_882,In_2333,In_3609);
nor U883 (N_883,In_4447,In_1227);
and U884 (N_884,In_3473,In_3968);
or U885 (N_885,In_2177,In_4326);
nor U886 (N_886,In_1194,In_4180);
and U887 (N_887,In_189,In_2056);
and U888 (N_888,In_4293,In_2268);
nand U889 (N_889,In_4612,In_3892);
xor U890 (N_890,In_2531,In_3270);
xnor U891 (N_891,In_4020,In_377);
or U892 (N_892,In_855,In_1679);
and U893 (N_893,In_4620,In_4721);
nand U894 (N_894,In_2544,In_1693);
and U895 (N_895,In_2321,In_1520);
and U896 (N_896,In_2761,In_2002);
nand U897 (N_897,In_579,In_4272);
and U898 (N_898,In_3678,In_1656);
nand U899 (N_899,In_3858,In_2243);
and U900 (N_900,In_3458,In_4922);
or U901 (N_901,In_472,In_1038);
and U902 (N_902,In_2923,In_628);
or U903 (N_903,In_4758,In_2525);
or U904 (N_904,In_2340,In_2760);
xnor U905 (N_905,In_1672,In_1889);
and U906 (N_906,In_1136,In_722);
or U907 (N_907,In_2102,In_2209);
nand U908 (N_908,In_259,In_941);
and U909 (N_909,In_4601,In_4292);
or U910 (N_910,In_4529,In_842);
and U911 (N_911,In_3671,In_1035);
nor U912 (N_912,In_2948,In_1700);
xor U913 (N_913,In_3836,In_3595);
and U914 (N_914,In_97,In_135);
nand U915 (N_915,In_1935,In_2226);
nand U916 (N_916,In_548,In_3422);
xnor U917 (N_917,In_1422,In_3275);
nor U918 (N_918,In_2474,In_1818);
nor U919 (N_919,In_956,In_4425);
nand U920 (N_920,In_4512,In_1335);
nor U921 (N_921,In_1727,In_2672);
and U922 (N_922,In_1904,In_1353);
and U923 (N_923,In_4563,In_3200);
nand U924 (N_924,In_4867,In_3084);
nor U925 (N_925,In_1231,In_2842);
nor U926 (N_926,In_3993,In_3581);
xnor U927 (N_927,In_3320,In_1983);
or U928 (N_928,In_2108,In_1711);
xor U929 (N_929,In_2356,In_1819);
or U930 (N_930,In_4573,In_2933);
nand U931 (N_931,In_3100,In_290);
or U932 (N_932,In_71,In_3116);
nand U933 (N_933,In_3653,In_1358);
nor U934 (N_934,In_741,In_2592);
and U935 (N_935,In_979,In_721);
nor U936 (N_936,In_269,In_4586);
xor U937 (N_937,In_3121,In_4152);
or U938 (N_938,In_621,In_2723);
or U939 (N_939,In_2756,In_134);
nor U940 (N_940,In_4329,In_1006);
nand U941 (N_941,In_2427,In_711);
and U942 (N_942,In_3760,In_9);
nand U943 (N_943,In_4908,In_3471);
nor U944 (N_944,In_3579,In_1017);
and U945 (N_945,In_3720,In_4966);
nor U946 (N_946,In_2739,In_4387);
and U947 (N_947,In_3508,In_2583);
and U948 (N_948,In_2456,In_286);
or U949 (N_949,In_1842,In_4333);
xnor U950 (N_950,In_4954,In_958);
xnor U951 (N_951,In_2856,In_3369);
xor U952 (N_952,In_2528,In_994);
nor U953 (N_953,In_3224,In_4805);
nand U954 (N_954,In_3463,In_2374);
xor U955 (N_955,In_850,In_3807);
nand U956 (N_956,In_3835,In_3067);
and U957 (N_957,In_4154,In_2943);
nand U958 (N_958,In_4256,In_1525);
and U959 (N_959,In_2867,In_667);
xor U960 (N_960,In_3881,In_1415);
nor U961 (N_961,In_1213,In_3352);
or U962 (N_962,In_1512,In_3716);
and U963 (N_963,In_1743,In_1732);
xnor U964 (N_964,In_1734,In_880);
and U965 (N_965,In_314,In_2661);
nor U966 (N_966,In_2236,In_3588);
or U967 (N_967,In_2908,In_4904);
or U968 (N_968,In_2553,In_4854);
nand U969 (N_969,In_4864,In_679);
and U970 (N_970,In_407,In_3531);
nand U971 (N_971,In_2828,In_2837);
or U972 (N_972,In_2911,In_3734);
nor U973 (N_973,In_2620,In_3592);
nor U974 (N_974,In_4131,In_666);
or U975 (N_975,In_2106,In_3223);
and U976 (N_976,In_3522,In_4578);
nand U977 (N_977,In_2472,In_923);
or U978 (N_978,In_3280,In_558);
nand U979 (N_979,In_1643,In_1910);
xor U980 (N_980,In_1198,In_2146);
and U981 (N_981,In_220,In_2117);
nor U982 (N_982,In_1654,In_2945);
nor U983 (N_983,In_1476,In_317);
xor U984 (N_984,In_4951,In_1033);
nor U985 (N_985,In_211,In_2237);
and U986 (N_986,In_1361,In_39);
nor U987 (N_987,In_4697,In_1756);
nand U988 (N_988,In_848,In_3335);
nor U989 (N_989,In_3417,In_1048);
nand U990 (N_990,In_1635,In_4773);
nand U991 (N_991,In_3431,In_2593);
xor U992 (N_992,In_1060,In_2336);
nor U993 (N_993,In_567,In_4370);
nor U994 (N_994,In_249,In_525);
xnor U995 (N_995,In_2608,In_4279);
xor U996 (N_996,In_2596,In_4274);
and U997 (N_997,In_1888,In_1046);
nor U998 (N_998,In_326,In_1334);
nor U999 (N_999,In_1212,In_4036);
or U1000 (N_1000,In_342,In_1110);
or U1001 (N_1001,In_229,In_3071);
and U1002 (N_1002,In_1099,In_1713);
nand U1003 (N_1003,In_2431,In_3890);
xnor U1004 (N_1004,In_2687,In_4098);
nor U1005 (N_1005,In_3827,In_1843);
and U1006 (N_1006,In_847,In_2931);
or U1007 (N_1007,In_2829,In_809);
xnor U1008 (N_1008,In_2773,In_2567);
or U1009 (N_1009,In_680,In_1517);
or U1010 (N_1010,In_4523,In_3957);
xnor U1011 (N_1011,In_3251,In_3351);
and U1012 (N_1012,In_867,In_4325);
and U1013 (N_1013,In_2168,In_2218);
or U1014 (N_1014,In_4608,In_4377);
nor U1015 (N_1015,In_787,In_1767);
and U1016 (N_1016,In_1081,In_316);
and U1017 (N_1017,In_3046,In_1129);
or U1018 (N_1018,In_3028,In_4792);
nor U1019 (N_1019,In_279,In_2386);
nand U1020 (N_1020,In_3929,In_3514);
xor U1021 (N_1021,In_780,In_4104);
or U1022 (N_1022,In_3022,In_2486);
or U1023 (N_1023,In_502,In_111);
nand U1024 (N_1024,In_255,In_1065);
or U1025 (N_1025,In_1360,In_2398);
xnor U1026 (N_1026,In_4434,In_4816);
or U1027 (N_1027,In_2526,In_3082);
nand U1028 (N_1028,In_2096,In_3665);
nand U1029 (N_1029,In_4695,In_2230);
nor U1030 (N_1030,In_3604,In_2878);
or U1031 (N_1031,In_2439,In_4332);
nor U1032 (N_1032,In_198,In_4489);
xor U1033 (N_1033,In_2160,In_889);
nor U1034 (N_1034,In_3916,In_2277);
nand U1035 (N_1035,In_2081,In_2991);
xnor U1036 (N_1036,In_916,In_4001);
nand U1037 (N_1037,In_3966,In_777);
and U1038 (N_1038,In_2981,In_3974);
or U1039 (N_1039,In_3432,In_2235);
and U1040 (N_1040,In_3688,In_2859);
xor U1041 (N_1041,In_4436,In_1973);
xnor U1042 (N_1042,In_3314,In_648);
nand U1043 (N_1043,In_4123,In_2041);
nor U1044 (N_1044,In_1425,In_1828);
and U1045 (N_1045,In_1184,In_2305);
xor U1046 (N_1046,In_859,In_2688);
xor U1047 (N_1047,In_768,In_3727);
nor U1048 (N_1048,In_1256,In_1068);
and U1049 (N_1049,In_2185,In_772);
nor U1050 (N_1050,In_2771,In_207);
or U1051 (N_1051,In_2792,In_3419);
or U1052 (N_1052,In_4533,In_2477);
nand U1053 (N_1053,In_3628,In_2135);
xnor U1054 (N_1054,In_890,In_2758);
or U1055 (N_1055,In_3856,In_3031);
xnor U1056 (N_1056,In_1416,In_382);
and U1057 (N_1057,In_1298,In_3323);
nor U1058 (N_1058,In_1812,In_4808);
nor U1059 (N_1059,In_2855,In_1988);
nor U1060 (N_1060,In_2578,In_4774);
xor U1061 (N_1061,In_4199,In_3003);
xnor U1062 (N_1062,In_3547,In_863);
nand U1063 (N_1063,In_3744,In_697);
or U1064 (N_1064,In_2793,In_1346);
nand U1065 (N_1065,In_1418,In_4985);
nor U1066 (N_1066,In_133,In_3342);
and U1067 (N_1067,In_1423,In_2517);
and U1068 (N_1068,In_2658,In_3445);
nand U1069 (N_1069,In_1161,In_1876);
xor U1070 (N_1070,In_4055,In_1436);
and U1071 (N_1071,In_1575,In_3683);
nor U1072 (N_1072,In_1919,In_1375);
nand U1073 (N_1073,In_3042,In_1101);
and U1074 (N_1074,In_3972,In_4276);
xor U1075 (N_1075,In_2324,In_4145);
xnor U1076 (N_1076,In_272,In_415);
nor U1077 (N_1077,In_3754,In_4791);
and U1078 (N_1078,In_434,In_4732);
or U1079 (N_1079,In_2902,In_3326);
or U1080 (N_1080,In_3090,In_4569);
xor U1081 (N_1081,In_1609,In_1223);
nand U1082 (N_1082,In_2192,In_3214);
nor U1083 (N_1083,In_2120,In_1214);
xor U1084 (N_1084,In_785,In_3177);
nand U1085 (N_1085,In_4027,In_4917);
or U1086 (N_1086,In_2191,In_2332);
nor U1087 (N_1087,In_1765,In_1366);
xnor U1088 (N_1088,In_1457,In_2695);
or U1089 (N_1089,In_1109,In_479);
nor U1090 (N_1090,In_78,In_989);
and U1091 (N_1091,In_3309,In_2772);
nand U1092 (N_1092,In_924,In_3751);
and U1093 (N_1093,In_3272,In_2070);
and U1094 (N_1094,In_2819,In_2848);
and U1095 (N_1095,In_2267,In_2341);
nor U1096 (N_1096,In_3329,In_4619);
nand U1097 (N_1097,In_3866,In_2742);
and U1098 (N_1098,In_3348,In_2215);
xnor U1099 (N_1099,In_905,In_4961);
nor U1100 (N_1100,In_4039,In_891);
nand U1101 (N_1101,In_4520,In_996);
or U1102 (N_1102,In_2144,In_116);
nor U1103 (N_1103,In_192,In_3376);
xor U1104 (N_1104,In_2639,In_4605);
nand U1105 (N_1105,In_4979,In_587);
nand U1106 (N_1106,In_3944,In_2607);
xor U1107 (N_1107,In_2314,In_4343);
nor U1108 (N_1108,In_3709,In_4209);
nand U1109 (N_1109,In_1646,In_3332);
xnor U1110 (N_1110,In_4167,In_3932);
nand U1111 (N_1111,In_2265,In_2085);
nor U1112 (N_1112,In_4108,In_1806);
or U1113 (N_1113,In_4570,In_4831);
xnor U1114 (N_1114,In_1549,In_4200);
and U1115 (N_1115,In_2494,In_2757);
and U1116 (N_1116,In_225,In_4711);
and U1117 (N_1117,In_363,In_4691);
xnor U1118 (N_1118,In_4686,In_2556);
and U1119 (N_1119,In_4282,In_1555);
and U1120 (N_1120,In_902,In_3231);
or U1121 (N_1121,In_571,In_3814);
nand U1122 (N_1122,In_1835,In_1004);
nor U1123 (N_1123,In_2648,In_4837);
nor U1124 (N_1124,In_1019,In_645);
nor U1125 (N_1125,In_98,In_1947);
nor U1126 (N_1126,In_764,In_3910);
nand U1127 (N_1127,In_2753,In_1971);
and U1128 (N_1128,In_3179,In_4085);
and U1129 (N_1129,In_3176,In_3662);
and U1130 (N_1130,In_707,In_4799);
nand U1131 (N_1131,In_2575,In_754);
and U1132 (N_1132,In_4901,In_4302);
and U1133 (N_1133,In_2692,In_1674);
nor U1134 (N_1134,In_2212,In_4940);
nor U1135 (N_1135,In_2281,In_3874);
and U1136 (N_1136,In_3906,In_486);
xor U1137 (N_1137,In_2781,In_967);
nor U1138 (N_1138,In_1055,In_300);
nand U1139 (N_1139,In_4948,In_4505);
nor U1140 (N_1140,In_678,In_3801);
and U1141 (N_1141,In_2112,In_2995);
nand U1142 (N_1142,In_3099,In_4640);
and U1143 (N_1143,In_3021,In_514);
xnor U1144 (N_1144,In_2869,In_2690);
nor U1145 (N_1145,In_2542,In_1850);
and U1146 (N_1146,In_3234,In_3985);
nor U1147 (N_1147,In_4885,In_1003);
nor U1148 (N_1148,In_4800,In_2726);
nand U1149 (N_1149,In_2571,In_1990);
or U1150 (N_1150,In_340,In_1302);
or U1151 (N_1151,In_4045,In_512);
xor U1152 (N_1152,In_4159,In_3920);
and U1153 (N_1153,In_4115,In_4192);
or U1154 (N_1154,In_529,In_1773);
or U1155 (N_1155,In_4994,In_1151);
nand U1156 (N_1156,In_2279,In_4739);
nor U1157 (N_1157,In_2361,In_3345);
nand U1158 (N_1158,In_4944,In_2257);
or U1159 (N_1159,In_743,In_3451);
nor U1160 (N_1160,In_146,In_3489);
xnor U1161 (N_1161,In_733,In_4813);
nor U1162 (N_1162,In_4842,In_3434);
nor U1163 (N_1163,In_4018,In_1869);
and U1164 (N_1164,In_2520,In_452);
nand U1165 (N_1165,In_1611,In_2987);
xor U1166 (N_1166,In_492,In_3967);
or U1167 (N_1167,In_2467,In_4598);
or U1168 (N_1168,In_1921,In_4221);
and U1169 (N_1169,In_895,In_3834);
and U1170 (N_1170,In_3603,In_1554);
xor U1171 (N_1171,In_3986,In_2392);
nand U1172 (N_1172,In_88,In_4763);
or U1173 (N_1173,In_3797,In_1498);
nand U1174 (N_1174,In_2861,In_3112);
nand U1175 (N_1175,In_203,In_1446);
or U1176 (N_1176,In_3040,In_160);
or U1177 (N_1177,In_2429,In_1600);
xnor U1178 (N_1178,In_3301,In_38);
and U1179 (N_1179,In_682,In_1495);
xor U1180 (N_1180,In_4120,In_1170);
nor U1181 (N_1181,In_968,In_4710);
or U1182 (N_1182,In_1762,In_876);
nor U1183 (N_1183,In_3252,In_4606);
or U1184 (N_1184,In_4680,In_4111);
nand U1185 (N_1185,In_589,In_2602);
nor U1186 (N_1186,In_3574,In_1094);
xor U1187 (N_1187,In_2216,In_1871);
xor U1188 (N_1188,In_2248,In_4466);
xnor U1189 (N_1189,In_18,In_3798);
xnor U1190 (N_1190,In_4937,In_4592);
nor U1191 (N_1191,In_473,In_3818);
and U1192 (N_1192,In_3393,In_2426);
nor U1193 (N_1193,In_40,In_4781);
xnor U1194 (N_1194,In_76,In_4759);
and U1195 (N_1195,In_2222,In_2717);
nand U1196 (N_1196,In_4355,In_3772);
xor U1197 (N_1197,In_2746,In_970);
nand U1198 (N_1198,In_1056,In_542);
nor U1199 (N_1199,In_729,In_4265);
and U1200 (N_1200,In_2715,In_1286);
nor U1201 (N_1201,In_2029,In_3069);
or U1202 (N_1202,In_3990,In_4285);
or U1203 (N_1203,In_1338,In_2478);
xnor U1204 (N_1204,In_2131,In_1877);
xor U1205 (N_1205,In_3501,In_3477);
or U1206 (N_1206,In_3815,In_2390);
xnor U1207 (N_1207,In_2105,In_2655);
xnor U1208 (N_1208,In_4090,In_603);
xnor U1209 (N_1209,In_2328,In_3786);
or U1210 (N_1210,In_4358,In_3527);
nand U1211 (N_1211,In_3567,In_3645);
or U1212 (N_1212,In_732,In_3118);
nor U1213 (N_1213,In_261,In_3334);
nand U1214 (N_1214,In_2186,In_1333);
xnor U1215 (N_1215,In_2519,In_4857);
nand U1216 (N_1216,In_555,In_1387);
and U1217 (N_1217,In_1820,In_4804);
nand U1218 (N_1218,In_1841,In_3164);
nand U1219 (N_1219,In_2459,In_4047);
or U1220 (N_1220,In_796,In_3913);
nand U1221 (N_1221,In_1217,In_886);
nor U1222 (N_1222,In_1412,In_4362);
or U1223 (N_1223,In_965,In_4821);
nor U1224 (N_1224,In_3997,In_387);
xnor U1225 (N_1225,In_2425,In_1204);
nor U1226 (N_1226,In_1378,In_4373);
or U1227 (N_1227,In_990,In_3091);
xor U1228 (N_1228,In_4409,In_1536);
nor U1229 (N_1229,In_2132,In_3291);
and U1230 (N_1230,In_1970,In_325);
and U1231 (N_1231,In_790,In_4178);
and U1232 (N_1232,In_3051,In_2646);
xnor U1233 (N_1233,In_976,In_4839);
and U1234 (N_1234,In_4017,In_1130);
or U1235 (N_1235,In_1556,In_3536);
nor U1236 (N_1236,In_1221,In_572);
and U1237 (N_1237,In_521,In_2442);
or U1238 (N_1238,In_2205,In_4894);
xnor U1239 (N_1239,In_3726,In_2093);
nand U1240 (N_1240,In_3049,In_1787);
or U1241 (N_1241,In_2270,In_2963);
nand U1242 (N_1242,In_1150,In_4126);
and U1243 (N_1243,In_3601,In_912);
or U1244 (N_1244,In_4637,In_251);
nor U1245 (N_1245,In_265,In_4749);
and U1246 (N_1246,In_2563,In_2437);
nand U1247 (N_1247,In_3461,In_2289);
nor U1248 (N_1248,In_2086,In_2876);
nor U1249 (N_1249,In_378,In_3864);
nand U1250 (N_1250,In_4631,In_3608);
nor U1251 (N_1251,In_3992,In_1748);
xor U1252 (N_1252,In_309,In_4320);
nor U1253 (N_1253,In_2565,In_127);
nor U1254 (N_1254,In_413,In_554);
xnor U1255 (N_1255,In_2312,In_4785);
xnor U1256 (N_1256,In_1011,In_4459);
xor U1257 (N_1257,In_2404,In_22);
nor U1258 (N_1258,In_1359,In_3636);
xnor U1259 (N_1259,In_1220,In_319);
and U1260 (N_1260,In_36,In_1481);
and U1261 (N_1261,In_3571,In_517);
xor U1262 (N_1262,In_964,In_1175);
or U1263 (N_1263,In_575,In_1691);
and U1264 (N_1264,In_4347,In_1659);
nand U1265 (N_1265,In_4743,In_197);
or U1266 (N_1266,In_3011,In_2183);
xnor U1267 (N_1267,In_2049,In_2376);
xnor U1268 (N_1268,In_3607,In_3089);
or U1269 (N_1269,In_4949,In_1975);
nor U1270 (N_1270,In_943,In_3041);
nand U1271 (N_1271,In_2405,In_2551);
xnor U1272 (N_1272,In_3435,In_3174);
or U1273 (N_1273,In_3878,In_1766);
nand U1274 (N_1274,In_4295,In_4230);
nand U1275 (N_1275,In_4496,In_823);
or U1276 (N_1276,In_124,In_1997);
nand U1277 (N_1277,In_2403,In_684);
xor U1278 (N_1278,In_4080,In_4977);
or U1279 (N_1279,In_1492,In_2109);
and U1280 (N_1280,In_778,In_3119);
nand U1281 (N_1281,In_1880,In_991);
xor U1282 (N_1282,In_3484,In_881);
xnor U1283 (N_1283,In_4836,In_4545);
nor U1284 (N_1284,In_4371,In_4797);
nand U1285 (N_1285,In_509,In_2800);
or U1286 (N_1286,In_2359,In_2909);
or U1287 (N_1287,In_4227,In_3855);
nand U1288 (N_1288,In_1875,In_887);
xnor U1289 (N_1289,In_1343,In_594);
and U1290 (N_1290,In_3217,In_1318);
or U1291 (N_1291,In_2180,In_395);
xor U1292 (N_1292,In_260,In_3098);
xor U1293 (N_1293,In_3640,In_2882);
xnor U1294 (N_1294,In_2031,In_1723);
xnor U1295 (N_1295,In_3114,In_1925);
and U1296 (N_1296,In_3548,In_2458);
nand U1297 (N_1297,In_3558,In_3629);
and U1298 (N_1298,In_1080,In_2241);
or U1299 (N_1299,In_187,In_2468);
and U1300 (N_1300,In_1807,In_2133);
and U1301 (N_1301,In_4968,In_1873);
nand U1302 (N_1302,In_1179,In_168);
nor U1303 (N_1303,In_1447,In_3961);
or U1304 (N_1304,In_4346,In_2171);
or U1305 (N_1305,In_4661,In_703);
nor U1306 (N_1306,In_4381,In_4705);
nor U1307 (N_1307,In_4128,In_1426);
or U1308 (N_1308,In_1496,In_2084);
nand U1309 (N_1309,In_2055,In_3883);
nor U1310 (N_1310,In_2453,In_2812);
and U1311 (N_1311,In_115,In_214);
and U1312 (N_1312,In_171,In_2654);
nor U1313 (N_1313,In_3043,In_1648);
xnor U1314 (N_1314,In_107,In_284);
nand U1315 (N_1315,In_4998,In_2960);
and U1316 (N_1316,In_4526,In_4782);
xor U1317 (N_1317,In_2208,In_797);
xnor U1318 (N_1318,In_623,In_4485);
or U1319 (N_1319,In_356,In_3264);
xnor U1320 (N_1320,In_2566,In_4281);
and U1321 (N_1321,In_4571,In_4655);
or U1322 (N_1322,In_634,In_4946);
xor U1323 (N_1323,In_4835,In_4037);
xor U1324 (N_1324,In_1107,In_698);
and U1325 (N_1325,In_2714,In_3168);
and U1326 (N_1326,In_4252,In_4138);
xnor U1327 (N_1327,In_24,In_2286);
and U1328 (N_1328,In_1685,In_3389);
and U1329 (N_1329,In_4162,In_1162);
xor U1330 (N_1330,In_2700,In_2530);
or U1331 (N_1331,In_1106,In_3430);
nor U1332 (N_1332,In_70,In_161);
xnor U1333 (N_1333,In_2919,In_280);
nand U1334 (N_1334,In_2916,In_920);
or U1335 (N_1335,In_3590,In_4196);
or U1336 (N_1336,In_3239,In_2473);
and U1337 (N_1337,In_1488,In_4895);
nor U1338 (N_1338,In_4015,In_4323);
nor U1339 (N_1339,In_4784,In_247);
and U1340 (N_1340,In_4891,In_4849);
or U1341 (N_1341,In_2500,In_4423);
nand U1342 (N_1342,In_1027,In_710);
nor U1343 (N_1343,In_1012,In_2786);
nand U1344 (N_1344,In_2721,In_4581);
nand U1345 (N_1345,In_2052,In_535);
nand U1346 (N_1346,In_4993,In_1328);
xor U1347 (N_1347,In_177,In_1417);
or U1348 (N_1348,In_4216,In_408);
xor U1349 (N_1349,In_2689,In_1159);
xor U1350 (N_1350,In_3512,In_4163);
or U1351 (N_1351,In_3054,In_2822);
nor U1352 (N_1352,In_2561,In_1057);
nor U1353 (N_1353,In_4943,In_350);
nor U1354 (N_1354,In_687,In_877);
nand U1355 (N_1355,In_4787,In_4403);
nand U1356 (N_1356,In_3641,In_759);
nand U1357 (N_1357,In_2154,In_322);
or U1358 (N_1358,In_4148,In_2839);
or U1359 (N_1359,In_3570,In_1480);
xnor U1360 (N_1360,In_3365,In_1956);
nand U1361 (N_1361,In_1473,In_836);
nand U1362 (N_1362,In_3774,In_4541);
xor U1363 (N_1363,In_4083,In_1195);
and U1364 (N_1364,In_1163,In_4546);
or U1365 (N_1365,In_2033,In_4032);
or U1366 (N_1366,In_4033,In_2874);
xor U1367 (N_1367,In_2488,In_1632);
xnor U1368 (N_1368,In_1915,In_2271);
xnor U1369 (N_1369,In_520,In_1735);
xnor U1370 (N_1370,In_833,In_1655);
and U1371 (N_1371,In_2585,In_4990);
nand U1372 (N_1372,In_3254,In_929);
nand U1373 (N_1373,In_278,In_4246);
nand U1374 (N_1374,In_4079,In_2423);
or U1375 (N_1375,In_2504,In_1201);
xor U1376 (N_1376,In_2682,In_4296);
and U1377 (N_1377,In_2722,In_1794);
or U1378 (N_1378,In_1293,In_2214);
or U1379 (N_1379,In_1449,In_3371);
xor U1380 (N_1380,In_2371,In_1142);
nor U1381 (N_1381,In_1036,In_3635);
and U1382 (N_1382,In_3111,In_438);
nand U1383 (N_1383,In_68,In_534);
xnor U1384 (N_1384,In_1758,In_4024);
nor U1385 (N_1385,In_756,In_1690);
nand U1386 (N_1386,In_1918,In_4284);
xor U1387 (N_1387,In_4040,In_1859);
nor U1388 (N_1388,In_140,In_3386);
xnor U1389 (N_1389,In_1553,In_4846);
nand U1390 (N_1390,In_4435,In_2028);
or U1391 (N_1391,In_285,In_3917);
and U1392 (N_1392,In_1891,In_2358);
nand U1393 (N_1393,In_676,In_3421);
nand U1394 (N_1394,In_3194,In_1494);
nor U1395 (N_1395,In_2251,In_4330);
or U1396 (N_1396,In_4356,In_3086);
nor U1397 (N_1397,In_4756,In_2738);
nand U1398 (N_1398,In_3963,In_4953);
or U1399 (N_1399,In_1502,In_1493);
nor U1400 (N_1400,In_1062,In_4887);
and U1401 (N_1401,In_4342,In_3013);
xnor U1402 (N_1402,In_436,In_4334);
nand U1403 (N_1403,In_458,In_4139);
and U1404 (N_1404,In_2683,In_1475);
nor U1405 (N_1405,In_1244,In_2136);
nor U1406 (N_1406,In_2234,In_2850);
or U1407 (N_1407,In_949,In_3063);
or U1408 (N_1408,In_2225,In_1013);
xor U1409 (N_1409,In_686,In_1782);
nor U1410 (N_1410,In_2522,In_857);
or U1411 (N_1411,In_1523,In_3740);
or U1412 (N_1412,In_3673,In_3690);
xor U1413 (N_1413,In_4702,In_619);
and U1414 (N_1414,In_1001,In_4930);
xor U1415 (N_1415,In_2503,In_1612);
or U1416 (N_1416,In_1228,In_2802);
nand U1417 (N_1417,In_3959,In_1617);
nor U1418 (N_1418,In_4963,In_2156);
nand U1419 (N_1419,In_2499,In_655);
nand U1420 (N_1420,In_1587,In_1913);
nand U1421 (N_1421,In_1697,In_399);
nor U1422 (N_1422,In_41,In_2872);
xnor U1423 (N_1423,In_4091,In_271);
nand U1424 (N_1424,In_1849,In_782);
xnor U1425 (N_1425,In_4468,In_270);
xnor U1426 (N_1426,In_3401,In_2759);
nor U1427 (N_1427,In_3076,In_100);
nand U1428 (N_1428,In_3915,In_2569);
nand U1429 (N_1429,In_374,In_2164);
nor U1430 (N_1430,In_987,In_4962);
or U1431 (N_1431,In_2401,In_13);
or U1432 (N_1432,In_695,In_1560);
nand U1433 (N_1433,In_4483,In_3582);
nor U1434 (N_1434,In_882,In_1257);
or U1435 (N_1435,In_4287,In_4424);
and U1436 (N_1436,In_3544,In_245);
nor U1437 (N_1437,In_3093,In_1901);
xor U1438 (N_1438,In_4155,In_1145);
or U1439 (N_1439,In_4589,In_1594);
and U1440 (N_1440,In_2100,In_1074);
or U1441 (N_1441,In_4959,In_2642);
nand U1442 (N_1442,In_3395,In_3066);
or U1443 (N_1443,In_4044,In_3810);
or U1444 (N_1444,In_4897,In_3020);
and U1445 (N_1445,In_1590,In_46);
and U1446 (N_1446,In_1856,In_19);
nor U1447 (N_1447,In_3493,In_3110);
xor U1448 (N_1448,In_933,In_4460);
and U1449 (N_1449,In_1448,In_2137);
xnor U1450 (N_1450,In_1313,In_3479);
nor U1451 (N_1451,In_3189,In_4022);
nor U1452 (N_1452,In_2844,In_3533);
and U1453 (N_1453,In_3907,In_2487);
and U1454 (N_1454,In_3283,In_4651);
xor U1455 (N_1455,In_985,In_2395);
and U1456 (N_1456,In_4621,In_1811);
xnor U1457 (N_1457,In_4510,In_318);
or U1458 (N_1458,In_1829,In_205);
nor U1459 (N_1459,In_4048,In_305);
nand U1460 (N_1460,In_2915,In_4548);
and U1461 (N_1461,In_4958,In_2174);
nand U1462 (N_1462,In_62,In_4479);
and U1463 (N_1463,In_2853,In_4733);
nand U1464 (N_1464,In_3753,In_2242);
xor U1465 (N_1465,In_4070,In_1424);
nor U1466 (N_1466,In_2387,In_3424);
or U1467 (N_1467,In_2865,In_3216);
nor U1468 (N_1468,In_2928,In_2936);
or U1469 (N_1469,In_1558,In_1396);
and U1470 (N_1470,In_1837,In_3971);
nor U1471 (N_1471,In_2704,In_2095);
or U1472 (N_1472,In_175,In_2187);
or U1473 (N_1473,In_400,In_3196);
and U1474 (N_1474,In_3843,In_4170);
nand U1475 (N_1475,In_4870,In_2645);
and U1476 (N_1476,In_2961,In_3142);
nor U1477 (N_1477,In_3138,In_4623);
nor U1478 (N_1478,In_4648,In_3127);
xor U1479 (N_1479,In_1134,In_755);
nor U1480 (N_1480,In_4609,In_4577);
nor U1481 (N_1481,In_2925,In_3416);
nor U1482 (N_1482,In_1538,In_1031);
nor U1483 (N_1483,In_939,In_1833);
nor U1484 (N_1484,In_1153,In_4888);
nand U1485 (N_1485,In_3150,In_37);
xor U1486 (N_1486,In_4933,In_2204);
xnor U1487 (N_1487,In_4696,In_4277);
nand U1488 (N_1488,In_865,In_3002);
nor U1489 (N_1489,In_854,In_4662);
nand U1490 (N_1490,In_2163,In_4615);
nand U1491 (N_1491,In_4076,In_2912);
nand U1492 (N_1492,In_4051,In_4882);
and U1493 (N_1493,In_4121,In_425);
xnor U1494 (N_1494,In_3481,In_829);
nand U1495 (N_1495,In_2294,In_4484);
xnor U1496 (N_1496,In_3221,In_3642);
and U1497 (N_1497,In_3778,In_4237);
or U1498 (N_1498,In_3587,In_315);
nor U1499 (N_1499,In_1937,In_463);
or U1500 (N_1500,In_2557,In_3222);
nand U1501 (N_1501,In_2958,In_30);
nand U1502 (N_1502,In_4635,In_344);
or U1503 (N_1503,In_4438,In_2008);
and U1504 (N_1504,In_149,In_2130);
xor U1505 (N_1505,In_1746,In_1628);
and U1506 (N_1506,In_2895,In_2975);
and U1507 (N_1507,In_2697,In_3442);
or U1508 (N_1508,In_3975,In_1468);
xor U1509 (N_1509,In_4902,In_4398);
nand U1510 (N_1510,In_3770,In_4129);
xor U1511 (N_1511,In_4160,In_1783);
nor U1512 (N_1512,In_2735,In_4207);
nor U1513 (N_1513,In_4150,In_1718);
and U1514 (N_1514,In_2546,In_2862);
nor U1515 (N_1515,In_3902,In_3934);
or U1516 (N_1516,In_2272,In_381);
nand U1517 (N_1517,In_562,In_2315);
xnor U1518 (N_1518,In_581,In_1886);
nor U1519 (N_1519,In_3965,In_1510);
xor U1520 (N_1520,In_4242,In_564);
nor U1521 (N_1521,In_689,In_2202);
and U1522 (N_1522,In_3296,In_3799);
xor U1523 (N_1523,In_4059,In_282);
xor U1524 (N_1524,In_1349,In_4502);
nand U1525 (N_1525,In_3933,In_1454);
or U1526 (N_1526,In_2600,In_1428);
xor U1527 (N_1527,In_1657,In_3068);
or U1528 (N_1528,In_893,In_2656);
and U1529 (N_1529,In_1582,In_3771);
xnor U1530 (N_1530,In_875,In_3363);
xnor U1531 (N_1531,In_4665,In_4007);
nand U1532 (N_1532,In_2990,In_1501);
nor U1533 (N_1533,In_592,In_497);
nand U1534 (N_1534,In_4629,In_2941);
nor U1535 (N_1535,In_4011,In_3622);
and U1536 (N_1536,In_209,In_1998);
nor U1537 (N_1537,In_860,In_4228);
xnor U1538 (N_1538,In_685,In_3777);
and U1539 (N_1539,In_3982,In_4886);
or U1540 (N_1540,In_3948,In_3464);
nor U1541 (N_1541,In_760,In_3773);
or U1542 (N_1542,In_2751,In_4238);
and U1543 (N_1543,In_3977,In_409);
xor U1544 (N_1544,In_3580,In_3669);
or U1545 (N_1545,In_3633,In_2357);
and U1546 (N_1546,In_2432,In_298);
or U1547 (N_1547,In_3367,In_4408);
or U1548 (N_1548,In_1769,In_4480);
nor U1549 (N_1549,In_1604,In_99);
and U1550 (N_1550,In_4290,In_3830);
or U1551 (N_1551,In_3979,In_2179);
and U1552 (N_1552,In_1920,In_1831);
or U1553 (N_1553,In_4197,In_2449);
nand U1554 (N_1554,In_608,In_2533);
nor U1555 (N_1555,In_4786,In_3572);
nor U1556 (N_1556,In_4433,In_2023);
or U1557 (N_1557,In_2223,In_3702);
xor U1558 (N_1558,In_4481,In_2181);
nand U1559 (N_1559,In_1105,In_4428);
nand U1560 (N_1560,In_3625,In_1222);
and U1561 (N_1561,In_4853,In_2383);
and U1562 (N_1562,In_2017,In_993);
or U1563 (N_1563,In_1152,In_536);
and U1564 (N_1564,In_4778,In_484);
xnor U1565 (N_1565,In_2465,In_4393);
xor U1566 (N_1566,In_2295,In_1932);
nor U1567 (N_1567,In_675,In_1461);
nor U1568 (N_1568,In_767,In_493);
xor U1569 (N_1569,In_1898,In_4338);
xor U1570 (N_1570,In_266,In_3659);
or U1571 (N_1571,In_2896,In_500);
xnor U1572 (N_1572,In_1701,In_4639);
nand U1573 (N_1573,In_1954,In_988);
and U1574 (N_1574,In_1744,In_3026);
nand U1575 (N_1575,In_1210,In_2466);
and U1576 (N_1576,In_2079,In_3008);
xnor U1577 (N_1577,In_3377,In_3983);
or U1578 (N_1578,In_4823,In_718);
or U1579 (N_1579,In_735,In_1568);
xor U1580 (N_1580,In_2030,In_3637);
nor U1581 (N_1581,In_866,In_12);
or U1582 (N_1582,In_1250,In_4003);
or U1583 (N_1583,In_2787,In_2884);
and U1584 (N_1584,In_4244,In_2870);
xor U1585 (N_1585,In_60,In_2736);
and U1586 (N_1586,In_1113,In_3876);
or U1587 (N_1587,In_1602,In_3550);
xnor U1588 (N_1588,In_1924,In_2325);
xnor U1589 (N_1589,In_3065,In_1269);
xor U1590 (N_1590,In_1677,In_239);
or U1591 (N_1591,In_1518,In_1731);
or U1592 (N_1592,In_3589,In_4752);
xor U1593 (N_1593,In_3719,In_4171);
nor U1594 (N_1594,In_3859,In_677);
nor U1595 (N_1595,In_2664,In_3691);
or U1596 (N_1596,In_4478,In_925);
xnor U1597 (N_1597,In_4043,In_1513);
xnor U1598 (N_1598,In_1326,In_1189);
or U1599 (N_1599,In_2348,In_2264);
and U1600 (N_1600,In_2584,In_4744);
xnor U1601 (N_1601,In_4266,In_717);
or U1602 (N_1602,In_3766,In_3151);
or U1603 (N_1603,In_3057,In_4143);
nor U1604 (N_1604,In_911,In_3052);
and U1605 (N_1605,In_757,In_1177);
nand U1606 (N_1606,In_3875,In_962);
or U1607 (N_1607,In_4699,In_4102);
xor U1608 (N_1608,In_4761,In_3029);
xnor U1609 (N_1609,In_3509,In_3160);
or U1610 (N_1610,In_2774,In_1724);
nor U1611 (N_1611,In_3081,In_4913);
nand U1612 (N_1612,In_4509,In_238);
nor U1613 (N_1613,In_4687,In_4730);
or U1614 (N_1614,In_3337,In_3540);
nor U1615 (N_1615,In_3279,In_4780);
nor U1616 (N_1616,In_3904,In_3134);
and U1617 (N_1617,In_85,In_1883);
xnor U1618 (N_1618,In_4550,In_3676);
nor U1619 (N_1619,In_3764,In_714);
and U1620 (N_1620,In_2482,In_4624);
xnor U1621 (N_1621,In_1550,In_2815);
or U1622 (N_1622,In_3085,In_4308);
xor U1623 (N_1623,In_4909,In_2651);
nor U1624 (N_1624,In_798,In_3769);
nor U1625 (N_1625,In_4644,In_869);
and U1626 (N_1626,In_2125,In_1025);
and U1627 (N_1627,In_2606,In_1254);
and U1628 (N_1628,In_2339,In_3340);
nand U1629 (N_1629,In_1715,In_1610);
xnor U1630 (N_1630,In_4164,In_4642);
or U1631 (N_1631,In_2072,In_1962);
xnor U1632 (N_1632,In_2979,In_1413);
or U1633 (N_1633,In_1085,In_330);
and U1634 (N_1634,In_2888,In_1589);
nand U1635 (N_1635,In_3392,In_4718);
and U1636 (N_1636,In_3889,In_3523);
and U1637 (N_1637,In_2586,In_4110);
nand U1638 (N_1638,In_4924,In_3779);
xnor U1639 (N_1639,In_3173,In_3289);
or U1640 (N_1640,In_1624,In_936);
nand U1641 (N_1641,In_4449,In_3611);
nor U1642 (N_1642,In_2873,In_862);
nand U1643 (N_1643,In_4991,In_1726);
nand U1644 (N_1644,In_3240,In_3494);
nand U1645 (N_1645,In_4147,In_4010);
and U1646 (N_1646,In_2806,In_362);
or U1647 (N_1647,In_2836,In_4769);
or U1648 (N_1648,In_948,In_3108);
and U1649 (N_1649,In_2344,In_846);
or U1650 (N_1650,In_1185,In_206);
nand U1651 (N_1651,In_2283,In_3163);
xnor U1652 (N_1652,In_4255,In_2428);
xor U1653 (N_1653,In_1489,In_657);
nor U1654 (N_1654,In_3840,In_150);
and U1655 (N_1655,In_2275,In_3358);
and U1656 (N_1656,In_4019,In_2811);
nor U1657 (N_1657,In_4919,In_1144);
and U1658 (N_1658,In_143,In_4584);
nand U1659 (N_1659,In_641,In_333);
nand U1660 (N_1660,In_4807,In_3044);
or U1661 (N_1661,In_2827,In_4880);
or U1662 (N_1662,In_3353,In_2306);
and U1663 (N_1663,In_1629,In_1092);
or U1664 (N_1664,In_4723,In_2078);
nand U1665 (N_1665,In_3705,In_4798);
nor U1666 (N_1666,In_4025,In_3696);
xor U1667 (N_1667,In_2605,In_334);
nand U1668 (N_1668,In_4280,In_3566);
xnor U1669 (N_1669,In_3627,In_2003);
or U1670 (N_1670,In_1315,In_2364);
xnor U1671 (N_1671,In_2059,In_1370);
nand U1672 (N_1672,In_1847,In_1309);
nand U1673 (N_1673,In_4223,In_2378);
nor U1674 (N_1674,In_1382,In_2444);
nor U1675 (N_1675,In_217,In_392);
nor U1676 (N_1676,In_2637,In_3298);
xnor U1677 (N_1677,In_3652,In_1728);
and U1678 (N_1678,In_4981,In_2747);
xnor U1679 (N_1679,In_3723,In_4729);
and U1680 (N_1680,In_4305,In_380);
or U1681 (N_1681,In_2420,In_1327);
and U1682 (N_1682,In_955,In_2703);
nor U1683 (N_1683,In_1401,In_1547);
nor U1684 (N_1684,In_4146,In_4859);
nand U1685 (N_1685,In_1117,In_1219);
nand U1686 (N_1686,In_2673,In_1407);
xnor U1687 (N_1687,In_3557,In_658);
or U1688 (N_1688,In_4719,In_527);
nor U1689 (N_1689,In_3321,In_4190);
or U1690 (N_1690,In_4939,In_3346);
xnor U1691 (N_1691,In_4069,In_2701);
and U1692 (N_1692,In_4748,In_231);
nor U1693 (N_1693,In_1972,In_622);
nand U1694 (N_1694,In_450,In_919);
nor U1695 (N_1695,In_595,In_1355);
or U1696 (N_1696,In_1867,In_1388);
nand U1697 (N_1697,In_141,In_453);
and U1698 (N_1698,In_4907,In_2046);
or U1699 (N_1699,In_3894,In_3366);
or U1700 (N_1700,In_2151,In_4866);
or U1701 (N_1701,In_3811,In_287);
nor U1702 (N_1702,In_2944,In_4008);
and U1703 (N_1703,In_3423,In_2322);
nor U1704 (N_1704,In_4156,In_3327);
nor U1705 (N_1705,In_3143,In_3630);
nand U1706 (N_1706,In_2510,In_1751);
nand U1707 (N_1707,In_4618,In_1939);
nor U1708 (N_1708,In_806,In_661);
or U1709 (N_1709,In_3349,In_2469);
xor U1710 (N_1710,In_4125,In_3831);
and U1711 (N_1711,In_4645,In_3039);
nor U1712 (N_1712,In_4482,In_3027);
nor U1713 (N_1713,In_2940,In_4731);
nand U1714 (N_1714,In_639,In_3820);
nor U1715 (N_1715,In_58,In_3155);
nand U1716 (N_1716,In_1324,In_4235);
or U1717 (N_1717,In_2053,In_3079);
and U1718 (N_1718,In_1362,In_2555);
nor U1719 (N_1719,In_1621,In_1907);
xor U1720 (N_1720,In_3958,In_3476);
xnor U1721 (N_1721,In_1969,In_1397);
and U1722 (N_1722,In_172,In_1307);
or U1723 (N_1723,In_353,In_4273);
nand U1724 (N_1724,In_4889,In_351);
xor U1725 (N_1725,In_2788,In_2698);
nand U1726 (N_1726,In_1156,In_1376);
xor U1727 (N_1727,In_2825,In_3800);
or U1728 (N_1728,In_2090,In_2462);
xnor U1729 (N_1729,In_2879,In_1443);
or U1730 (N_1730,In_2502,In_795);
xor U1731 (N_1731,In_467,In_3511);
nor U1732 (N_1732,In_816,In_4193);
or U1733 (N_1733,In_616,In_2169);
nand U1734 (N_1734,In_701,In_2069);
nand U1735 (N_1735,In_4925,In_427);
nor U1736 (N_1736,In_1802,In_975);
and U1737 (N_1737,In_2615,In_1192);
or U1738 (N_1738,In_2536,In_1945);
and U1739 (N_1739,In_1950,In_3338);
and U1740 (N_1740,In_901,In_4822);
nand U1741 (N_1741,In_2728,In_43);
or U1742 (N_1742,In_2061,In_4976);
nor U1743 (N_1743,In_1961,In_3647);
or U1744 (N_1744,In_2572,In_4340);
and U1745 (N_1745,In_636,In_1862);
xnor U1746 (N_1746,In_354,In_306);
nor U1747 (N_1747,In_3829,In_2891);
or U1748 (N_1748,In_468,In_4524);
or U1749 (N_1749,In_1086,In_596);
or U1750 (N_1750,In_1509,In_2391);
or U1751 (N_1751,In_1398,In_2290);
nor U1752 (N_1752,In_1682,In_2719);
nor U1753 (N_1753,In_3553,In_3765);
xnor U1754 (N_1754,In_4353,In_357);
or U1755 (N_1755,In_4421,In_971);
and U1756 (N_1756,In_928,In_1805);
nand U1757 (N_1757,In_2415,In_4142);
or U1758 (N_1758,In_1095,In_3828);
nor U1759 (N_1759,In_1775,In_758);
nor U1760 (N_1760,In_2198,In_1045);
nand U1761 (N_1761,In_1503,In_1500);
and U1762 (N_1762,In_4335,In_419);
nor U1763 (N_1763,In_3062,In_4987);
or U1764 (N_1764,In_3867,In_83);
nor U1765 (N_1765,In_4247,In_1902);
and U1766 (N_1766,In_339,In_2167);
xor U1767 (N_1767,In_1702,In_2413);
and U1768 (N_1768,In_2725,In_2050);
and U1769 (N_1769,In_329,In_2394);
nor U1770 (N_1770,In_4061,In_3978);
and U1771 (N_1771,In_625,In_1855);
nand U1772 (N_1772,In_2720,In_4527);
xor U1773 (N_1773,In_3412,In_3541);
xor U1774 (N_1774,In_303,In_3869);
or U1775 (N_1775,In_1342,In_794);
nor U1776 (N_1776,In_4777,In_4400);
xor U1777 (N_1777,In_2115,In_1838);
xnor U1778 (N_1778,In_368,In_3517);
or U1779 (N_1779,In_825,In_1661);
xnor U1780 (N_1780,In_1905,In_3271);
xor U1781 (N_1781,In_2952,In_4350);
and U1782 (N_1782,In_3561,In_2042);
and U1783 (N_1783,In_1132,In_1253);
and U1784 (N_1784,In_800,In_2564);
and U1785 (N_1785,In_766,In_4029);
xnor U1786 (N_1786,In_4625,In_1796);
nor U1787 (N_1787,In_2080,In_3593);
xnor U1788 (N_1788,In_3472,In_2966);
or U1789 (N_1789,In_1483,In_1953);
nand U1790 (N_1790,In_3452,In_72);
or U1791 (N_1791,In_4071,In_2379);
and U1792 (N_1792,In_852,In_1899);
nor U1793 (N_1793,In_736,In_151);
nand U1794 (N_1794,In_3281,In_1673);
or U1795 (N_1795,In_195,In_1139);
or U1796 (N_1796,In_1631,In_2913);
nand U1797 (N_1797,In_1039,In_2014);
or U1798 (N_1798,In_3380,In_1870);
nor U1799 (N_1799,In_2508,In_1548);
and U1800 (N_1800,In_1112,In_4971);
and U1801 (N_1801,In_4926,In_1104);
xnor U1802 (N_1802,In_3433,In_258);
or U1803 (N_1803,In_1942,In_1149);
or U1804 (N_1804,In_2724,In_918);
or U1805 (N_1805,In_700,In_896);
xnor U1806 (N_1806,In_4231,In_3537);
and U1807 (N_1807,In_3406,In_1581);
xor U1808 (N_1808,In_3460,In_2172);
or U1809 (N_1809,In_264,In_2483);
nand U1810 (N_1810,In_4309,In_433);
nand U1811 (N_1811,In_3577,In_4396);
nor U1812 (N_1812,In_2384,In_1283);
xor U1813 (N_1813,In_1625,In_1155);
nor U1814 (N_1814,In_4674,In_3478);
nor U1815 (N_1815,In_3695,In_1312);
and U1816 (N_1816,In_2211,In_2005);
nand U1817 (N_1817,In_2785,In_4830);
or U1818 (N_1818,In_268,In_2594);
and U1819 (N_1819,In_1215,In_3201);
nand U1820 (N_1820,In_1249,In_723);
xnor U1821 (N_1821,In_537,In_557);
and U1822 (N_1822,In_3989,In_2200);
xor U1823 (N_1823,In_1395,In_934);
and U1824 (N_1824,In_4877,In_153);
or U1825 (N_1825,In_3060,In_2126);
nor U1826 (N_1826,In_843,In_1652);
and U1827 (N_1827,In_1405,In_349);
nor U1828 (N_1828,In_3555,In_33);
or U1829 (N_1829,In_1482,In_3873);
and U1830 (N_1830,In_3955,In_336);
nor U1831 (N_1831,In_4497,In_1863);
and U1832 (N_1832,In_3722,In_4518);
or U1833 (N_1833,In_1280,In_3755);
and U1834 (N_1834,In_2524,In_3373);
or U1835 (N_1835,In_2128,In_2523);
xor U1836 (N_1836,In_1649,In_4658);
xor U1837 (N_1837,In_461,In_3469);
or U1838 (N_1838,In_2278,In_1063);
or U1839 (N_1839,In_1579,In_4005);
xor U1840 (N_1840,In_2436,In_4187);
or U1841 (N_1841,In_781,In_4559);
or U1842 (N_1842,In_712,In_4259);
and U1843 (N_1843,In_4712,In_1238);
nand U1844 (N_1844,In_3017,In_1158);
nor U1845 (N_1845,In_4879,In_1186);
xor U1846 (N_1846,In_2626,In_2189);
nand U1847 (N_1847,In_1688,In_464);
and U1848 (N_1848,In_57,In_3286);
nor U1849 (N_1849,In_10,In_3559);
and U1850 (N_1850,In_1761,In_1963);
and U1851 (N_1851,In_751,In_3839);
nand U1852 (N_1852,In_1174,In_277);
nand U1853 (N_1853,In_737,In_4992);
and U1854 (N_1854,In_2776,In_1123);
nor U1855 (N_1855,In_321,In_2794);
xnor U1856 (N_1856,In_1764,In_3382);
and U1857 (N_1857,In_1043,In_4311);
or U1858 (N_1858,In_947,In_4972);
xnor U1859 (N_1859,In_4141,In_4186);
or U1860 (N_1860,In_3096,In_110);
nor U1861 (N_1861,In_2497,In_2422);
and U1862 (N_1862,In_3613,In_4176);
nor U1863 (N_1863,In_310,In_627);
xnor U1864 (N_1864,In_1098,In_1394);
or U1865 (N_1865,In_412,In_2892);
or U1866 (N_1866,In_4906,In_3816);
nand U1867 (N_1867,In_3762,In_668);
and U1868 (N_1868,In_1050,In_2629);
or U1869 (N_1869,In_4404,In_2511);
or U1870 (N_1870,In_3276,In_4013);
or U1871 (N_1871,In_1459,In_3171);
nor U1872 (N_1872,In_2643,In_563);
nand U1873 (N_1873,In_244,In_1780);
xnor U1874 (N_1874,In_818,In_690);
nand U1875 (N_1875,In_2247,In_2905);
nand U1876 (N_1876,In_1895,In_2949);
xnor U1877 (N_1877,In_1164,In_4668);
or U1878 (N_1878,In_2562,In_390);
or U1879 (N_1879,In_3998,In_2107);
and U1880 (N_1880,In_3586,In_4352);
or U1881 (N_1881,In_469,In_2129);
nor U1882 (N_1882,In_1745,In_2886);
nand U1883 (N_1883,In_533,In_1347);
and U1884 (N_1884,In_1530,In_2353);
xnor U1885 (N_1885,In_2711,In_1917);
nor U1886 (N_1886,In_2716,In_1356);
or U1887 (N_1887,In_2820,In_2789);
nor U1888 (N_1888,In_713,In_4094);
nand U1889 (N_1889,In_2791,In_2675);
and U1890 (N_1890,In_4881,In_4088);
nand U1891 (N_1891,In_248,In_3539);
xnor U1892 (N_1892,In_1111,In_2507);
and U1893 (N_1893,In_3871,In_289);
xor U1894 (N_1894,In_915,In_4973);
nand U1895 (N_1895,In_2032,In_1072);
or U1896 (N_1896,In_52,In_4659);
nor U1897 (N_1897,In_3265,In_2765);
nand U1898 (N_1898,In_4084,In_234);
or U1899 (N_1899,In_3732,In_202);
nor U1900 (N_1900,In_1858,In_2194);
nor U1901 (N_1901,In_1916,In_1578);
nand U1902 (N_1902,In_212,In_2176);
nand U1903 (N_1903,In_3768,In_541);
nand U1904 (N_1904,In_466,In_959);
nor U1905 (N_1905,In_1128,In_343);
or U1906 (N_1906,In_25,In_1120);
and U1907 (N_1907,In_4671,In_4063);
xnor U1908 (N_1908,In_1960,In_283);
xor U1909 (N_1909,In_4504,In_1668);
nor U1910 (N_1910,In_2330,In_4399);
xor U1911 (N_1911,In_1469,In_832);
xnor U1912 (N_1912,In_2311,In_3787);
nor U1913 (N_1913,In_3569,In_2628);
and U1914 (N_1914,In_3414,In_3844);
nor U1915 (N_1915,In_4713,In_2441);
or U1916 (N_1916,In_2114,In_1208);
and U1917 (N_1917,In_3530,In_1730);
and U1918 (N_1918,In_386,In_1273);
nor U1919 (N_1919,In_2470,In_2852);
and U1920 (N_1920,In_706,In_4693);
or U1921 (N_1921,In_3763,In_610);
nand U1922 (N_1922,In_839,In_631);
or U1923 (N_1923,In_2063,In_3520);
and U1924 (N_1924,In_2617,In_3860);
nand U1925 (N_1925,In_3841,In_2702);
or U1926 (N_1926,In_1037,In_2904);
or U1927 (N_1927,In_3374,In_4075);
nand U1928 (N_1928,In_2763,In_2591);
xnor U1929 (N_1929,In_669,In_4916);
nand U1930 (N_1930,In_830,In_2351);
nor U1931 (N_1931,In_1541,In_1800);
xnor U1932 (N_1932,In_659,In_1445);
nand U1933 (N_1933,In_844,In_35);
or U1934 (N_1934,In_3526,In_3024);
and U1935 (N_1935,In_4401,In_3981);
nor U1936 (N_1936,In_1897,In_145);
or U1937 (N_1937,In_331,In_578);
or U1938 (N_1938,In_2446,In_80);
nand U1939 (N_1939,In_1172,In_4100);
or U1940 (N_1940,In_1143,In_411);
and U1941 (N_1941,In_125,In_4351);
or U1942 (N_1942,In_1176,In_2274);
xnor U1943 (N_1943,In_3243,In_2255);
and U1944 (N_1944,In_3420,In_222);
and U1945 (N_1945,In_3480,In_2667);
xor U1946 (N_1946,In_4936,In_2448);
xor U1947 (N_1947,In_2529,In_4657);
and U1948 (N_1948,In_2346,In_1992);
or U1949 (N_1949,In_2830,In_4893);
and U1950 (N_1950,In_4306,In_2512);
nand U1951 (N_1951,In_2821,In_620);
and U1952 (N_1952,In_1544,In_1647);
or U1953 (N_1953,In_4970,In_1882);
and U1954 (N_1954,In_673,In_2734);
nand U1955 (N_1955,In_1790,In_4006);
and U1956 (N_1956,In_570,In_1148);
or U1957 (N_1957,In_405,In_819);
nor U1958 (N_1958,In_726,In_3721);
nand U1959 (N_1959,In_4672,In_2397);
xor U1960 (N_1960,In_3694,In_4967);
nand U1961 (N_1961,In_4030,In_858);
nand U1962 (N_1962,In_3228,In_246);
or U1963 (N_1963,In_4597,In_4349);
and U1964 (N_1964,In_3616,In_2890);
nor U1965 (N_1965,In_3684,In_1314);
xor U1966 (N_1966,In_2875,In_1486);
and U1967 (N_1967,In_4386,In_3663);
or U1968 (N_1968,In_1034,In_4583);
or U1969 (N_1969,In_173,In_4742);
and U1970 (N_1970,In_952,In_1171);
xnor U1971 (N_1971,In_1330,In_1680);
nor U1972 (N_1972,In_1058,In_3584);
nor U1973 (N_1973,In_1053,In_4955);
nor U1974 (N_1974,In_165,In_1911);
or U1975 (N_1975,In_1830,In_114);
nor U1976 (N_1976,In_3885,In_613);
xnor U1977 (N_1977,In_4000,In_2011);
nor U1978 (N_1978,In_2124,In_496);
and U1979 (N_1979,In_2926,In_457);
nand U1980 (N_1980,In_293,In_1429);
xor U1981 (N_1981,In_3462,In_4678);
or U1982 (N_1982,In_2199,In_4708);
and U1983 (N_1983,In_2973,In_2598);
or U1984 (N_1984,In_1566,In_3409);
xnor U1985 (N_1985,In_262,In_2015);
xnor U1986 (N_1986,In_3776,In_3053);
or U1987 (N_1987,In_3370,In_2985);
or U1988 (N_1988,In_3515,In_2292);
xnor U1989 (N_1989,In_2938,In_3884);
or U1990 (N_1990,In_365,In_873);
nor U1991 (N_1991,In_2246,In_2676);
or U1992 (N_1992,In_1662,In_237);
nand U1993 (N_1993,In_1245,In_1392);
and U1994 (N_1994,In_4222,In_804);
or U1995 (N_1995,In_1720,In_2612);
and U1996 (N_1996,In_5,In_4511);
nor U1997 (N_1997,In_3408,In_3946);
nor U1998 (N_1998,In_3513,In_1606);
nand U1999 (N_1999,In_3739,In_1183);
xor U2000 (N_2000,In_4314,In_2705);
xor U2001 (N_2001,In_228,In_3378);
or U2002 (N_2002,In_2104,In_861);
nor U2003 (N_2003,In_2296,In_4360);
or U2004 (N_2004,In_4521,In_4168);
nor U2005 (N_2005,In_3681,In_4173);
xor U2006 (N_2006,In_2613,In_1096);
or U2007 (N_2007,In_953,In_373);
or U2008 (N_2008,In_1698,In_74);
or U2009 (N_2009,In_2691,In_2549);
xor U2010 (N_2010,In_3936,In_3287);
nand U2011 (N_2011,In_2922,In_47);
or U2012 (N_2012,In_1845,In_3146);
or U2013 (N_2013,In_3792,In_2694);
nor U2014 (N_2014,In_4327,In_4874);
nand U2015 (N_2015,In_491,In_2817);
or U2016 (N_2016,In_4064,In_4514);
and U2017 (N_2017,In_1049,In_1261);
or U2018 (N_2018,In_417,In_2959);
or U2019 (N_2019,In_974,In_696);
nand U2020 (N_2020,In_559,In_978);
nor U2021 (N_2021,In_1809,In_3080);
and U2022 (N_2022,In_1371,In_1943);
or U2023 (N_2023,In_565,In_4555);
or U2024 (N_2024,In_3064,In_600);
nor U2025 (N_2025,In_1957,In_2083);
xor U2026 (N_2026,In_4643,In_379);
and U2027 (N_2027,In_2652,In_545);
or U2028 (N_2028,In_4751,In_4551);
nor U2029 (N_2029,In_2903,In_3575);
xnor U2030 (N_2030,In_2094,In_2016);
or U2031 (N_2031,In_2228,In_1739);
or U2032 (N_2032,In_1456,In_4788);
xor U2033 (N_2033,In_3167,In_2755);
and U2034 (N_2034,In_549,In_14);
nand U2035 (N_2035,In_3614,In_4576);
or U2036 (N_2036,In_4594,In_4487);
nor U2037 (N_2037,In_4241,In_606);
nand U2038 (N_2038,In_257,In_2145);
and U2039 (N_2039,In_2367,In_4988);
xor U2040 (N_2040,In_2479,In_3524);
or U2041 (N_2041,In_3973,In_3996);
or U2042 (N_2042,In_1721,In_4653);
xor U2043 (N_2043,In_3903,In_1);
xnor U2044 (N_2044,In_3241,In_224);
nand U2045 (N_2045,In_2227,In_420);
nand U2046 (N_2046,In_3898,In_4975);
nor U2047 (N_2047,In_4023,In_2416);
nand U2048 (N_2048,In_4775,In_1040);
and U2049 (N_2049,In_3294,In_3969);
and U2050 (N_2050,In_3564,In_77);
or U2051 (N_2051,In_813,In_89);
nand U2052 (N_2052,In_3930,In_1430);
nand U2053 (N_2053,In_2337,In_2623);
nand U2054 (N_2054,In_3033,In_4026);
and U2055 (N_2055,In_4969,In_2285);
xnor U2056 (N_2056,In_1887,In_1015);
nand U2057 (N_2057,In_4768,In_815);
nand U2058 (N_2058,In_2347,In_0);
nor U2059 (N_2059,In_1597,In_3945);
or U2060 (N_2060,In_4507,In_3425);
xor U2061 (N_2061,In_4974,In_4892);
nor U2062 (N_2062,In_1108,In_1633);
nor U2063 (N_2063,In_1569,In_997);
or U2064 (N_2064,In_4677,In_3102);
nand U2065 (N_2065,In_4134,In_201);
xnor U2066 (N_2066,In_196,In_3960);
xnor U2067 (N_2067,In_1102,In_274);
xnor U2068 (N_2068,In_4097,In_584);
nand U2069 (N_2069,In_2043,In_4935);
nor U2070 (N_2070,In_1258,In_1173);
nand U2071 (N_2071,In_1296,In_2745);
and U2072 (N_2072,In_742,In_2);
xnor U2073 (N_2073,In_4947,In_2475);
xor U2074 (N_2074,In_2838,In_4271);
xnor U2075 (N_2075,In_4493,In_3403);
or U2076 (N_2076,In_4124,In_3742);
xor U2077 (N_2077,In_4679,In_4604);
and U2078 (N_2078,In_3738,In_786);
and U2079 (N_2079,In_3666,In_2680);
and U2080 (N_2080,In_2138,In_972);
nand U2081 (N_2081,In_2313,In_1986);
nor U2082 (N_2082,In_193,In_644);
nor U2083 (N_2083,In_4580,In_1071);
xnor U2084 (N_2084,In_1572,In_3970);
nand U2085 (N_2085,In_2037,In_1097);
nand U2086 (N_2086,In_3293,In_904);
nor U2087 (N_2087,In_3498,In_4053);
nor U2088 (N_2088,In_2824,In_2670);
or U2089 (N_2089,In_4137,In_2767);
nand U2090 (N_2090,In_3175,In_4762);
nor U2091 (N_2091,In_1747,In_2380);
or U2092 (N_2092,In_793,In_986);
nand U2093 (N_2093,In_826,In_4294);
nand U2094 (N_2094,In_1463,In_2238);
or U2095 (N_2095,In_4636,In_3926);
or U2096 (N_2096,In_2743,In_1592);
nor U2097 (N_2097,In_2288,In_3521);
nor U2098 (N_2098,In_2784,In_1785);
nand U2099 (N_2099,In_4188,In_2650);
or U2100 (N_2100,In_3506,In_4319);
nor U2101 (N_2101,In_2411,In_3428);
nor U2102 (N_2102,In_4560,In_3227);
xnor U2103 (N_2103,In_311,In_2843);
or U2104 (N_2104,In_1676,In_3606);
and U2105 (N_2105,In_4060,In_3724);
and U2106 (N_2106,In_585,In_650);
xnor U2107 (N_2107,In_1282,In_4627);
or U2108 (N_2108,In_139,In_218);
nor U2109 (N_2109,In_4114,In_3545);
nand U2110 (N_2110,In_1687,In_4475);
xnor U2111 (N_2111,In_4073,In_2067);
and U2112 (N_2112,In_2058,In_2343);
and U2113 (N_2113,In_2501,In_2640);
nor U2114 (N_2114,In_3237,In_2505);
xor U2115 (N_2115,In_637,In_2749);
nor U2116 (N_2116,In_1630,In_1271);
xor U2117 (N_2117,In_831,In_3697);
and U2118 (N_2118,In_3165,In_4833);
xnor U2119 (N_2119,In_26,In_1760);
nor U2120 (N_2120,In_3706,In_3750);
and U2121 (N_2121,In_4501,In_4331);
xor U2122 (N_2122,In_3717,In_2559);
nor U2123 (N_2123,In_3504,In_4458);
xnor U2124 (N_2124,In_3161,In_1710);
and U2125 (N_2125,In_1516,In_2206);
xor U2126 (N_2126,In_4184,In_3483);
xnor U2127 (N_2127,In_3023,In_624);
or U2128 (N_2128,In_2433,In_109);
nand U2129 (N_2129,In_4989,In_3157);
nor U2130 (N_2130,In_1016,In_2832);
and U2131 (N_2131,In_254,In_4582);
nor U2132 (N_2132,In_942,In_3180);
xnor U2133 (N_2133,In_3137,In_1909);
or U2134 (N_2134,In_2920,In_2663);
xnor U2135 (N_2135,In_3863,In_1340);
or U2136 (N_2136,In_2421,In_944);
nor U2137 (N_2137,In_3324,In_3821);
or U2138 (N_2138,In_3775,In_2547);
nor U2139 (N_2139,In_2969,In_2463);
xnor U2140 (N_2140,In_4224,In_2978);
and U2141 (N_2141,In_385,In_118);
or U2142 (N_2142,In_1020,In_2350);
nand U2143 (N_2143,In_1822,In_727);
and U2144 (N_2144,In_1928,In_4794);
nand U2145 (N_2145,In_138,In_167);
or U2146 (N_2146,In_2649,In_4136);
and U2147 (N_2147,In_3212,In_338);
and U2148 (N_2148,In_591,In_4532);
nand U2149 (N_2149,In_154,In_487);
or U2150 (N_2150,In_1763,In_4720);
nand U2151 (N_2151,In_4038,In_3058);
and U2152 (N_2152,In_4928,In_3924);
xor U2153 (N_2153,In_4341,In_3909);
or U2154 (N_2154,In_4709,In_4795);
or U2155 (N_2155,In_2082,In_2036);
nand U2156 (N_2156,In_966,In_2320);
and U2157 (N_2157,In_2752,In_179);
and U2158 (N_2158,In_725,In_2010);
nand U2159 (N_2159,In_4440,In_2338);
nand U2160 (N_2160,In_4789,In_1465);
and U2161 (N_2161,In_51,In_1306);
or U2162 (N_2162,In_2303,In_4530);
nand U2163 (N_2163,In_2527,In_788);
and U2164 (N_2164,In_2539,In_4442);
or U2165 (N_2165,In_3129,In_4508);
nor U2166 (N_2166,In_4537,In_824);
or U2167 (N_2167,In_1666,In_144);
xor U2168 (N_2168,In_4617,In_2713);
and U2169 (N_2169,In_853,In_3295);
or U2170 (N_2170,In_1260,In_4996);
nand U2171 (N_2171,In_2982,In_4543);
nor U2172 (N_2172,In_3879,In_2581);
and U2173 (N_2173,In_3893,In_577);
and U2174 (N_2174,In_1090,In_48);
xor U2175 (N_2175,In_2300,In_11);
nor U2176 (N_2176,In_4534,In_1675);
xnor U2177 (N_2177,In_1808,In_4950);
or U2178 (N_2178,In_2580,In_1653);
and U2179 (N_2179,In_1165,In_3735);
or U2180 (N_2180,In_4054,In_1704);
or U2181 (N_2181,In_2217,In_3730);
nand U2182 (N_2182,In_130,In_3788);
or U2183 (N_2183,In_1893,In_2057);
or U2184 (N_2184,In_588,In_1026);
and U2185 (N_2185,In_1410,In_1166);
nand U2186 (N_2186,In_2744,In_307);
nand U2187 (N_2187,In_2910,In_1291);
nor U2188 (N_2188,In_478,In_4552);
or U2189 (N_2189,In_1458,In_3427);
and U2190 (N_2190,In_4253,In_4165);
or U2191 (N_2191,In_765,In_1341);
and U2192 (N_2192,In_3263,In_183);
nor U2193 (N_2193,In_4876,In_2587);
xor U2194 (N_2194,In_416,In_1000);
and U2195 (N_2195,In_323,In_105);
nand U2196 (N_2196,In_1663,In_4796);
or U2197 (N_2197,In_3793,In_1369);
or U2198 (N_2198,In_4593,In_4414);
nor U2199 (N_2199,In_1857,In_2552);
xnor U2200 (N_2200,In_4740,In_1824);
nand U2201 (N_2201,In_2280,In_3838);
nor U2202 (N_2202,In_3980,In_3525);
or U2203 (N_2203,In_3197,In_2299);
nand U2204 (N_2204,In_2464,In_3826);
and U2205 (N_2205,In_1637,In_4204);
xor U2206 (N_2206,In_3937,In_1586);
and U2207 (N_2207,In_3822,In_3072);
and U2208 (N_2208,In_3215,In_4087);
nand U2209 (N_2209,In_352,In_45);
or U2210 (N_2210,In_3328,In_1235);
or U2211 (N_2211,In_3680,In_3488);
or U2212 (N_2212,In_1205,In_609);
or U2213 (N_2213,In_3809,In_4488);
nor U2214 (N_2214,In_1100,In_488);
nand U2215 (N_2215,In_3055,In_2779);
nand U2216 (N_2216,In_404,In_522);
nor U2217 (N_2217,In_4217,In_1616);
nand U2218 (N_2218,In_2362,In_1620);
nand U2219 (N_2219,In_4174,In_4322);
nand U2220 (N_2220,In_4046,In_1288);
or U2221 (N_2221,In_2318,In_73);
or U2222 (N_2222,In_3384,In_4212);
nor U2223 (N_2223,In_2455,In_1931);
nand U2224 (N_2224,In_3949,In_4426);
nand U2225 (N_2225,In_2887,In_2777);
xnor U2226 (N_2226,In_3819,In_1270);
and U2227 (N_2227,In_2939,In_4806);
xnor U2228 (N_2228,In_871,In_551);
and U2229 (N_2229,In_868,In_4384);
or U2230 (N_2230,In_499,In_4439);
and U2231 (N_2231,In_4366,In_1024);
or U2232 (N_2232,In_158,In_4692);
nor U2233 (N_2233,In_4476,In_4812);
nand U2234 (N_2234,In_691,In_3900);
nor U2235 (N_2235,In_2000,In_4021);
or U2236 (N_2236,In_4727,In_241);
nand U2237 (N_2237,In_837,In_313);
xor U2238 (N_2238,In_2917,In_2775);
nor U2239 (N_2239,In_921,In_3166);
nor U2240 (N_2240,In_3953,In_3248);
and U2241 (N_2241,In_4074,In_4848);
or U2242 (N_2242,In_2762,In_3159);
and U2243 (N_2243,In_4477,In_513);
nor U2244 (N_2244,In_4650,In_1608);
nor U2245 (N_2245,In_4681,In_4540);
or U2246 (N_2246,In_3375,In_3467);
and U2247 (N_2247,In_4531,In_1061);
or U2248 (N_2248,In_2588,In_2834);
or U2249 (N_2249,In_2024,In_376);
nor U2250 (N_2250,In_4067,In_4214);
and U2251 (N_2251,In_1289,In_561);
nand U2252 (N_2252,In_3803,In_2798);
xor U2253 (N_2253,In_1642,In_1317);
xnor U2254 (N_2254,In_1088,In_1684);
nor U2255 (N_2255,In_504,In_2054);
and U2256 (N_2256,In_3202,In_2382);
nor U2257 (N_2257,In_1391,In_4336);
nor U2258 (N_2258,In_4841,In_4009);
nor U2259 (N_2259,In_3450,In_1853);
or U2260 (N_2260,In_470,In_2149);
xnor U2261 (N_2261,In_4096,In_3097);
xnor U2262 (N_2262,In_1442,In_4912);
and U2263 (N_2263,In_4109,In_2127);
nor U2264 (N_2264,In_1242,In_1336);
and U2265 (N_2265,In_2614,In_626);
or U2266 (N_2266,In_3383,In_4685);
and U2267 (N_2267,In_4772,In_2638);
xnor U2268 (N_2268,In_1551,In_1564);
or U2269 (N_2269,In_1400,In_1900);
xnor U2270 (N_2270,In_1640,In_4494);
xnor U2271 (N_2271,In_328,In_1439);
and U2272 (N_2272,In_2363,In_568);
nand U2273 (N_2273,In_3758,In_1303);
or U2274 (N_2274,In_674,In_523);
nor U2275 (N_2275,In_253,In_4982);
nand U2276 (N_2276,In_87,In_371);
nor U2277 (N_2277,In_981,In_1069);
and U2278 (N_2278,In_94,In_821);
or U2279 (N_2279,In_3447,In_3310);
and U2280 (N_2280,In_250,In_2863);
nor U2281 (N_2281,In_1332,In_2123);
nand U2282 (N_2282,In_3490,In_874);
or U2283 (N_2283,In_552,In_181);
xnor U2284 (N_2284,In_3233,In_1462);
nand U2285 (N_2285,In_1542,In_544);
and U2286 (N_2286,In_232,In_3791);
and U2287 (N_2287,In_3631,In_3756);
nand U2288 (N_2288,In_1093,In_4910);
xnor U2289 (N_2289,In_969,In_3036);
and U2290 (N_2290,In_3503,In_604);
or U2291 (N_2291,In_2706,In_17);
nand U2292 (N_2292,In_2506,In_3132);
xnor U2293 (N_2293,In_236,In_3790);
and U2294 (N_2294,In_3415,In_3618);
and U2295 (N_2295,In_1846,In_2461);
nand U2296 (N_2296,In_2310,In_792);
nor U2297 (N_2297,In_1976,In_1964);
nor U2298 (N_2298,In_3994,In_1583);
and U2299 (N_2299,In_1749,In_388);
nand U2300 (N_2300,In_3390,In_4236);
nand U2301 (N_2301,In_1736,In_372);
or U2302 (N_2302,In_3016,In_938);
nor U2303 (N_2303,In_147,In_3354);
or U2304 (N_2304,In_633,In_3745);
nor U2305 (N_2305,In_4133,In_2161);
or U2306 (N_2306,In_1738,In_618);
nand U2307 (N_2307,In_927,In_900);
nor U2308 (N_2308,In_586,In_3596);
nor U2309 (N_2309,In_4828,In_221);
and U2310 (N_2310,In_1264,In_3711);
nand U2311 (N_2311,In_1946,In_888);
xnor U2312 (N_2312,In_4300,In_3311);
xor U2313 (N_2313,In_1522,In_4135);
or U2314 (N_2314,In_3789,In_3896);
nand U2315 (N_2315,In_121,In_1987);
and U2316 (N_2316,In_1890,In_3578);
xor U2317 (N_2317,In_1619,In_922);
nand U2318 (N_2318,In_638,In_506);
and U2319 (N_2319,In_3336,In_2988);
or U2320 (N_2320,In_137,In_2253);
or U2321 (N_2321,In_872,In_4119);
nand U2322 (N_2322,In_1753,In_3355);
xor U2323 (N_2323,In_4490,In_4911);
xor U2324 (N_2324,In_4471,In_4750);
and U2325 (N_2325,In_3429,In_501);
nand U2326 (N_2326,In_3018,In_65);
or U2327 (N_2327,In_3648,In_1914);
nand U2328 (N_2328,In_4153,In_4307);
nor U2329 (N_2329,In_2410,In_2610);
or U2330 (N_2330,In_123,In_2399);
and U2331 (N_2331,In_1879,In_2558);
nor U2332 (N_2332,In_2025,In_4406);
and U2333 (N_2333,In_299,In_15);
or U2334 (N_2334,In_761,In_1168);
or U2335 (N_2335,In_3396,In_1912);
nand U2336 (N_2336,In_640,In_3343);
and U2337 (N_2337,In_3845,In_2708);
xnor U2338 (N_2338,In_2750,In_598);
xor U2339 (N_2339,In_1507,In_4089);
or U2340 (N_2340,In_3529,In_4790);
or U2341 (N_2341,In_1265,In_1354);
xor U2342 (N_2342,In_3703,In_1406);
or U2343 (N_2343,In_4542,In_3410);
nand U2344 (N_2344,In_3400,In_4183);
nand U2345 (N_2345,In_2577,In_2309);
or U2346 (N_2346,In_566,In_3149);
xor U2347 (N_2347,In_2847,In_2388);
xnor U2348 (N_2348,In_4766,In_2385);
xnor U2349 (N_2349,In_4372,In_3905);
and U2350 (N_2350,In_3105,In_483);
nor U2351 (N_2351,In_649,In_1784);
nor U2352 (N_2352,In_2635,In_4945);
and U2353 (N_2353,In_1209,In_397);
and U2354 (N_2354,In_3302,In_2143);
nor U2355 (N_2355,In_3956,In_4202);
and U2356 (N_2356,In_1658,In_1772);
or U2357 (N_2357,In_776,In_4451);
nand U2358 (N_2358,In_2091,In_3891);
and U2359 (N_2359,In_2568,In_3449);
and U2360 (N_2360,In_4002,In_3737);
nand U2361 (N_2361,In_4465,In_1241);
and U2362 (N_2362,In_1008,In_2986);
or U2363 (N_2363,In_3886,In_4446);
nand U2364 (N_2364,In_940,In_2159);
or U2365 (N_2365,In_1595,In_3195);
xnor U2366 (N_2366,In_358,In_106);
nor U2367 (N_2367,In_2521,In_2599);
nand U2368 (N_2368,In_4269,In_4116);
and U2369 (N_2369,In_1363,In_3277);
nor U2370 (N_2370,In_1393,In_3418);
xnor U2371 (N_2371,In_4587,In_359);
and U2372 (N_2372,In_4899,In_3205);
and U2373 (N_2373,In_738,In_2540);
nand U2374 (N_2374,In_2040,In_1030);
or U2375 (N_2375,In_2946,In_1032);
nor U2376 (N_2376,In_4454,In_4117);
nand U2377 (N_2377,In_4675,In_1607);
or U2378 (N_2378,In_4934,In_2737);
and U2379 (N_2379,In_4359,In_4660);
nor U2380 (N_2380,In_2207,In_2389);
and U2381 (N_2381,In_4905,In_394);
xnor U2382 (N_2382,In_4676,In_2993);
and U2383 (N_2383,In_1795,In_1247);
nor U2384 (N_2384,In_155,In_1848);
nor U2385 (N_2385,In_4585,In_4415);
nor U2386 (N_2386,In_275,In_3573);
xor U2387 (N_2387,In_1420,In_630);
nand U2388 (N_2388,In_3391,In_2492);
nand U2389 (N_2389,In_3837,In_4741);
or U2390 (N_2390,In_4862,In_2976);
xnor U2391 (N_2391,In_1968,In_1005);
and U2392 (N_2392,In_2062,In_1639);
nor U2393 (N_2393,In_2007,In_769);
or U2394 (N_2394,In_4455,In_2360);
nand U2395 (N_2395,In_569,In_435);
or U2396 (N_2396,In_950,In_4042);
and U2397 (N_2397,In_1352,In_4169);
or U2398 (N_2398,In_1411,In_7);
nor U2399 (N_2399,In_3101,In_1325);
nand U2400 (N_2400,In_426,In_4354);
nor U2401 (N_2401,In_4248,In_2921);
nand U2402 (N_2402,In_396,In_3308);
and U2403 (N_2403,In_3083,In_4315);
nor U2404 (N_2404,In_2261,In_4140);
nor U2405 (N_2405,In_102,In_617);
or U2406 (N_2406,In_2406,In_2375);
xnor U2407 (N_2407,In_3306,In_4517);
or U2408 (N_2408,In_1345,In_2182);
or U2409 (N_2409,In_152,In_4519);
nor U2410 (N_2410,In_4918,In_3259);
or U2411 (N_2411,In_1464,In_8);
nor U2412 (N_2412,In_4310,In_447);
nand U2413 (N_2413,In_4717,In_233);
or U2414 (N_2414,In_1618,In_2262);
or U2415 (N_2415,In_235,In_1948);
nand U2416 (N_2416,In_2377,In_810);
nor U2417 (N_2417,In_597,In_4462);
xor U2418 (N_2418,In_3315,In_4602);
nand U2419 (N_2419,In_3185,In_1771);
nor U2420 (N_2420,In_113,In_440);
nor U2421 (N_2421,In_3255,In_3245);
nor U2422 (N_2422,In_2657,In_2158);
or U2423 (N_2423,In_3853,In_1781);
xnor U2424 (N_2424,In_771,In_4875);
nor U2425 (N_2425,In_1733,In_1272);
nand U2426 (N_2426,In_2877,In_3045);
nand U2427 (N_2427,In_3646,In_1372);
or U2428 (N_2428,In_884,In_3184);
xnor U2429 (N_2429,In_1337,In_1259);
and U2430 (N_2430,In_1989,In_715);
nor U2431 (N_2431,In_3576,In_2801);
and U2432 (N_2432,In_2282,In_4288);
xnor U2433 (N_2433,In_4068,In_337);
and U2434 (N_2434,In_3087,In_4378);
nand U2435 (N_2435,In_4245,In_2190);
nand U2436 (N_2436,In_1552,In_2352);
or U2437 (N_2437,In_2871,In_2809);
nor U2438 (N_2438,In_2001,In_4634);
or U2439 (N_2439,In_4198,In_4896);
nor U2440 (N_2440,In_2103,In_605);
or U2441 (N_2441,In_1705,In_4649);
xnor U2442 (N_2442,In_802,In_4267);
nand U2443 (N_2443,In_3725,In_3107);
or U2444 (N_2444,In_681,In_3887);
xnor U2445 (N_2445,In_599,In_4430);
and U2446 (N_2446,In_27,In_1266);
xnor U2447 (N_2447,In_2977,In_4767);
xnor U2448 (N_2448,In_3385,In_495);
nand U2449 (N_2449,In_402,In_1160);
nand U2450 (N_2450,In_3193,In_590);
nor U2451 (N_2451,In_1729,In_770);
and U2452 (N_2452,In_3619,In_4049);
or U2453 (N_2453,In_4118,In_2476);
xor U2454 (N_2454,In_3733,In_1707);
nand U2455 (N_2455,In_1559,In_1651);
or U2456 (N_2456,In_851,In_2173);
and U2457 (N_2457,In_4554,In_3109);
or U2458 (N_2458,In_811,In_2611);
nand U2459 (N_2459,In_3398,In_1798);
nor U2460 (N_2460,In_3126,In_1029);
or U2461 (N_2461,In_1994,In_230);
xnor U2462 (N_2462,In_1466,In_2302);
nor U2463 (N_2463,In_2409,In_1545);
or U2464 (N_2464,In_1519,In_1868);
nor U2465 (N_2465,In_4884,In_3130);
nand U2466 (N_2466,In_4144,In_2481);
and U2467 (N_2467,In_518,In_1073);
and U2468 (N_2468,In_1934,In_3947);
nor U2469 (N_2469,In_243,In_4832);
nor U2470 (N_2470,In_1114,In_1797);
and U2471 (N_2471,In_213,In_4941);
and U2472 (N_2472,In_879,In_4312);
or U2473 (N_2473,In_4395,In_4986);
and U2474 (N_2474,In_656,In_1316);
and U2475 (N_2475,In_3139,In_480);
and U2476 (N_2476,In_1722,In_82);
xnor U2477 (N_2477,In_3426,In_3330);
and U2478 (N_2478,In_476,In_4820);
nand U2479 (N_2479,In_3153,In_3104);
nand U2480 (N_2480,In_1121,In_1115);
or U2481 (N_2481,In_2260,In_2148);
and U2482 (N_2482,In_2092,In_1526);
and U2483 (N_2483,In_4983,In_355);
nand U2484 (N_2484,In_226,In_1348);
or U2485 (N_2485,In_692,In_2213);
nor U2486 (N_2486,In_897,In_2826);
nor U2487 (N_2487,In_4753,In_92);
and U2488 (N_2488,In_3145,In_2034);
nor U2489 (N_2489,In_3672,In_4500);
and U2490 (N_2490,In_2790,In_2323);
xor U2491 (N_2491,In_573,In_367);
nor U2492 (N_2492,In_3518,In_4);
and U2493 (N_2493,In_3698,In_3436);
xnor U2494 (N_2494,In_1042,In_2139);
or U2495 (N_2495,In_4041,In_2039);
and U2496 (N_2496,In_2365,In_4898);
nor U2497 (N_2497,In_4441,In_740);
nor U2498 (N_2498,In_1321,In_3748);
xor U2499 (N_2499,In_1534,In_1927);
nor U2500 (N_2500,In_2933,In_4134);
nor U2501 (N_2501,In_4446,In_2471);
or U2502 (N_2502,In_2850,In_1793);
and U2503 (N_2503,In_1091,In_4931);
or U2504 (N_2504,In_596,In_4571);
or U2505 (N_2505,In_956,In_2642);
and U2506 (N_2506,In_933,In_1263);
and U2507 (N_2507,In_4479,In_2533);
or U2508 (N_2508,In_2375,In_764);
and U2509 (N_2509,In_149,In_2701);
or U2510 (N_2510,In_3537,In_911);
and U2511 (N_2511,In_931,In_3036);
or U2512 (N_2512,In_4083,In_2081);
nor U2513 (N_2513,In_2797,In_4995);
and U2514 (N_2514,In_2062,In_3077);
nand U2515 (N_2515,In_351,In_2406);
nor U2516 (N_2516,In_141,In_1014);
and U2517 (N_2517,In_1416,In_1087);
nand U2518 (N_2518,In_656,In_2915);
xnor U2519 (N_2519,In_2447,In_1456);
and U2520 (N_2520,In_1607,In_3460);
nand U2521 (N_2521,In_3947,In_2971);
and U2522 (N_2522,In_2289,In_1383);
xnor U2523 (N_2523,In_2392,In_212);
nand U2524 (N_2524,In_3300,In_2734);
xor U2525 (N_2525,In_424,In_2555);
nand U2526 (N_2526,In_2062,In_3140);
or U2527 (N_2527,In_1352,In_1020);
nor U2528 (N_2528,In_1588,In_4678);
xor U2529 (N_2529,In_112,In_3132);
and U2530 (N_2530,In_504,In_161);
and U2531 (N_2531,In_4844,In_2766);
xor U2532 (N_2532,In_1632,In_4966);
nand U2533 (N_2533,In_1969,In_1333);
or U2534 (N_2534,In_87,In_4343);
nor U2535 (N_2535,In_960,In_3256);
xor U2536 (N_2536,In_907,In_3520);
nor U2537 (N_2537,In_728,In_670);
nor U2538 (N_2538,In_2174,In_2710);
nor U2539 (N_2539,In_4618,In_4169);
nor U2540 (N_2540,In_3996,In_2749);
and U2541 (N_2541,In_1182,In_954);
xor U2542 (N_2542,In_1706,In_3336);
or U2543 (N_2543,In_3253,In_1120);
nand U2544 (N_2544,In_3636,In_2608);
nand U2545 (N_2545,In_1720,In_4398);
nor U2546 (N_2546,In_4704,In_2310);
and U2547 (N_2547,In_1043,In_4788);
xor U2548 (N_2548,In_2133,In_1179);
nor U2549 (N_2549,In_2899,In_3508);
and U2550 (N_2550,In_4693,In_3231);
or U2551 (N_2551,In_4185,In_4647);
nor U2552 (N_2552,In_743,In_1469);
xnor U2553 (N_2553,In_1991,In_4420);
and U2554 (N_2554,In_2847,In_4655);
nor U2555 (N_2555,In_3683,In_724);
nand U2556 (N_2556,In_2614,In_260);
nor U2557 (N_2557,In_2217,In_355);
nand U2558 (N_2558,In_3200,In_4498);
nand U2559 (N_2559,In_485,In_3254);
or U2560 (N_2560,In_4786,In_2741);
or U2561 (N_2561,In_3284,In_227);
nand U2562 (N_2562,In_1069,In_4078);
nand U2563 (N_2563,In_456,In_3114);
nor U2564 (N_2564,In_2167,In_676);
and U2565 (N_2565,In_3191,In_3485);
xor U2566 (N_2566,In_2967,In_2985);
xor U2567 (N_2567,In_580,In_3886);
xnor U2568 (N_2568,In_63,In_3949);
nand U2569 (N_2569,In_13,In_773);
nand U2570 (N_2570,In_4751,In_3506);
xnor U2571 (N_2571,In_4446,In_196);
nor U2572 (N_2572,In_2948,In_1180);
and U2573 (N_2573,In_3526,In_4771);
xnor U2574 (N_2574,In_4630,In_2949);
or U2575 (N_2575,In_944,In_4914);
xor U2576 (N_2576,In_1768,In_23);
and U2577 (N_2577,In_4810,In_1599);
and U2578 (N_2578,In_3876,In_3118);
and U2579 (N_2579,In_3470,In_4103);
and U2580 (N_2580,In_3406,In_137);
nand U2581 (N_2581,In_1976,In_822);
nand U2582 (N_2582,In_3166,In_4199);
or U2583 (N_2583,In_2174,In_1105);
or U2584 (N_2584,In_2575,In_3375);
nor U2585 (N_2585,In_4052,In_4888);
or U2586 (N_2586,In_1501,In_363);
xnor U2587 (N_2587,In_3282,In_73);
or U2588 (N_2588,In_1183,In_3522);
nor U2589 (N_2589,In_3003,In_2920);
nand U2590 (N_2590,In_2720,In_1252);
xnor U2591 (N_2591,In_4090,In_956);
nor U2592 (N_2592,In_2345,In_1537);
and U2593 (N_2593,In_1082,In_476);
xnor U2594 (N_2594,In_1575,In_454);
and U2595 (N_2595,In_4441,In_4128);
and U2596 (N_2596,In_3912,In_4581);
xor U2597 (N_2597,In_1297,In_716);
and U2598 (N_2598,In_949,In_826);
and U2599 (N_2599,In_1035,In_4923);
and U2600 (N_2600,In_2288,In_2371);
nand U2601 (N_2601,In_4467,In_1048);
nor U2602 (N_2602,In_207,In_3746);
xnor U2603 (N_2603,In_4851,In_940);
nand U2604 (N_2604,In_2875,In_3493);
nand U2605 (N_2605,In_4130,In_1496);
nand U2606 (N_2606,In_3770,In_3742);
nand U2607 (N_2607,In_463,In_1042);
nand U2608 (N_2608,In_671,In_775);
xnor U2609 (N_2609,In_674,In_3499);
and U2610 (N_2610,In_3114,In_1960);
or U2611 (N_2611,In_4269,In_3282);
nor U2612 (N_2612,In_2047,In_4709);
xnor U2613 (N_2613,In_724,In_308);
and U2614 (N_2614,In_693,In_1711);
nor U2615 (N_2615,In_2954,In_991);
or U2616 (N_2616,In_2846,In_1315);
and U2617 (N_2617,In_3875,In_748);
nand U2618 (N_2618,In_302,In_2246);
or U2619 (N_2619,In_2544,In_832);
nor U2620 (N_2620,In_2863,In_4878);
xnor U2621 (N_2621,In_3916,In_451);
nand U2622 (N_2622,In_4256,In_4596);
and U2623 (N_2623,In_1846,In_4005);
xnor U2624 (N_2624,In_4257,In_1838);
nor U2625 (N_2625,In_399,In_1756);
nand U2626 (N_2626,In_1791,In_3901);
nor U2627 (N_2627,In_177,In_4369);
nand U2628 (N_2628,In_1435,In_2019);
and U2629 (N_2629,In_900,In_1345);
nor U2630 (N_2630,In_2257,In_4851);
nand U2631 (N_2631,In_2927,In_3014);
xnor U2632 (N_2632,In_918,In_3131);
and U2633 (N_2633,In_511,In_1018);
or U2634 (N_2634,In_3572,In_3543);
nand U2635 (N_2635,In_2100,In_2091);
and U2636 (N_2636,In_2111,In_3157);
nand U2637 (N_2637,In_1312,In_839);
nand U2638 (N_2638,In_2630,In_667);
xnor U2639 (N_2639,In_716,In_843);
and U2640 (N_2640,In_2699,In_1717);
and U2641 (N_2641,In_3880,In_1902);
and U2642 (N_2642,In_2519,In_2980);
xnor U2643 (N_2643,In_4330,In_1522);
nand U2644 (N_2644,In_2887,In_1155);
nor U2645 (N_2645,In_2956,In_1106);
nor U2646 (N_2646,In_4606,In_1789);
nor U2647 (N_2647,In_2323,In_376);
nand U2648 (N_2648,In_818,In_4573);
nand U2649 (N_2649,In_1412,In_3008);
or U2650 (N_2650,In_2694,In_3551);
xnor U2651 (N_2651,In_249,In_2501);
and U2652 (N_2652,In_2697,In_2051);
nor U2653 (N_2653,In_2260,In_3244);
and U2654 (N_2654,In_4483,In_3878);
or U2655 (N_2655,In_3121,In_2085);
nor U2656 (N_2656,In_968,In_4131);
nand U2657 (N_2657,In_4844,In_4573);
or U2658 (N_2658,In_3983,In_2260);
or U2659 (N_2659,In_3347,In_860);
xor U2660 (N_2660,In_702,In_2801);
xnor U2661 (N_2661,In_489,In_4729);
nor U2662 (N_2662,In_2577,In_4103);
nand U2663 (N_2663,In_1689,In_2911);
nor U2664 (N_2664,In_4959,In_1922);
nand U2665 (N_2665,In_2219,In_2131);
nor U2666 (N_2666,In_1672,In_1499);
xnor U2667 (N_2667,In_1185,In_2397);
xnor U2668 (N_2668,In_4033,In_4689);
nor U2669 (N_2669,In_4091,In_3508);
and U2670 (N_2670,In_2828,In_209);
or U2671 (N_2671,In_1495,In_2213);
xnor U2672 (N_2672,In_4722,In_2766);
nand U2673 (N_2673,In_4094,In_2234);
or U2674 (N_2674,In_219,In_1624);
and U2675 (N_2675,In_3606,In_4468);
xnor U2676 (N_2676,In_2508,In_1381);
or U2677 (N_2677,In_980,In_2244);
nand U2678 (N_2678,In_4005,In_1048);
xnor U2679 (N_2679,In_1148,In_4903);
and U2680 (N_2680,In_2518,In_999);
nand U2681 (N_2681,In_4078,In_3440);
nand U2682 (N_2682,In_4549,In_2502);
and U2683 (N_2683,In_4574,In_558);
nor U2684 (N_2684,In_3163,In_4878);
and U2685 (N_2685,In_3239,In_828);
and U2686 (N_2686,In_2916,In_1907);
nor U2687 (N_2687,In_943,In_421);
xor U2688 (N_2688,In_3495,In_2483);
nor U2689 (N_2689,In_554,In_4745);
or U2690 (N_2690,In_134,In_4453);
xor U2691 (N_2691,In_4513,In_280);
xor U2692 (N_2692,In_4446,In_634);
and U2693 (N_2693,In_3249,In_596);
nor U2694 (N_2694,In_1501,In_3543);
nor U2695 (N_2695,In_4011,In_1507);
or U2696 (N_2696,In_3544,In_1921);
nand U2697 (N_2697,In_900,In_3930);
nor U2698 (N_2698,In_1352,In_2898);
nand U2699 (N_2699,In_772,In_4527);
nor U2700 (N_2700,In_4517,In_3647);
nor U2701 (N_2701,In_152,In_3480);
nand U2702 (N_2702,In_279,In_4779);
or U2703 (N_2703,In_1077,In_1827);
or U2704 (N_2704,In_2949,In_3580);
or U2705 (N_2705,In_4897,In_89);
xnor U2706 (N_2706,In_3301,In_865);
xnor U2707 (N_2707,In_4965,In_871);
or U2708 (N_2708,In_179,In_2307);
xnor U2709 (N_2709,In_4767,In_2851);
nor U2710 (N_2710,In_4932,In_4921);
nor U2711 (N_2711,In_3324,In_3706);
and U2712 (N_2712,In_2263,In_4335);
and U2713 (N_2713,In_3839,In_1359);
nand U2714 (N_2714,In_304,In_3951);
nand U2715 (N_2715,In_1348,In_4625);
and U2716 (N_2716,In_366,In_2523);
or U2717 (N_2717,In_768,In_1509);
or U2718 (N_2718,In_1700,In_3092);
nand U2719 (N_2719,In_2175,In_4197);
or U2720 (N_2720,In_3333,In_2364);
nand U2721 (N_2721,In_4723,In_4695);
or U2722 (N_2722,In_3435,In_3515);
xnor U2723 (N_2723,In_4657,In_1376);
and U2724 (N_2724,In_487,In_1501);
nand U2725 (N_2725,In_2041,In_374);
xor U2726 (N_2726,In_2378,In_3652);
or U2727 (N_2727,In_2012,In_3297);
nor U2728 (N_2728,In_3809,In_1934);
xnor U2729 (N_2729,In_1465,In_2744);
or U2730 (N_2730,In_2794,In_205);
or U2731 (N_2731,In_4671,In_4878);
nor U2732 (N_2732,In_4906,In_3886);
xor U2733 (N_2733,In_2970,In_3886);
or U2734 (N_2734,In_1640,In_2097);
xor U2735 (N_2735,In_1352,In_4254);
and U2736 (N_2736,In_2808,In_3781);
and U2737 (N_2737,In_3393,In_476);
xnor U2738 (N_2738,In_4516,In_369);
nand U2739 (N_2739,In_2147,In_3602);
nand U2740 (N_2740,In_694,In_2511);
xnor U2741 (N_2741,In_772,In_3228);
and U2742 (N_2742,In_1926,In_4673);
or U2743 (N_2743,In_3032,In_3367);
xnor U2744 (N_2744,In_2798,In_662);
or U2745 (N_2745,In_4905,In_801);
nand U2746 (N_2746,In_928,In_4293);
xnor U2747 (N_2747,In_4138,In_407);
or U2748 (N_2748,In_1399,In_3354);
or U2749 (N_2749,In_3292,In_823);
and U2750 (N_2750,In_1137,In_3903);
nor U2751 (N_2751,In_2871,In_4060);
nand U2752 (N_2752,In_1619,In_2813);
or U2753 (N_2753,In_4527,In_2868);
and U2754 (N_2754,In_2890,In_3523);
nand U2755 (N_2755,In_2272,In_374);
or U2756 (N_2756,In_834,In_3298);
or U2757 (N_2757,In_2121,In_108);
xor U2758 (N_2758,In_129,In_1630);
and U2759 (N_2759,In_1510,In_1179);
and U2760 (N_2760,In_4336,In_4264);
nor U2761 (N_2761,In_1123,In_1853);
or U2762 (N_2762,In_1143,In_4482);
xor U2763 (N_2763,In_3088,In_2366);
nand U2764 (N_2764,In_3211,In_4928);
or U2765 (N_2765,In_2178,In_2917);
or U2766 (N_2766,In_4784,In_2404);
and U2767 (N_2767,In_2403,In_3145);
or U2768 (N_2768,In_3639,In_3011);
nor U2769 (N_2769,In_4086,In_4732);
xnor U2770 (N_2770,In_4253,In_3600);
or U2771 (N_2771,In_921,In_3619);
or U2772 (N_2772,In_560,In_1776);
and U2773 (N_2773,In_2565,In_1950);
xnor U2774 (N_2774,In_4883,In_984);
nor U2775 (N_2775,In_2850,In_3818);
xor U2776 (N_2776,In_4648,In_3962);
and U2777 (N_2777,In_3761,In_3255);
and U2778 (N_2778,In_4681,In_12);
nor U2779 (N_2779,In_3759,In_2334);
nand U2780 (N_2780,In_2940,In_3548);
nand U2781 (N_2781,In_2181,In_1107);
or U2782 (N_2782,In_560,In_1502);
xnor U2783 (N_2783,In_3986,In_1935);
nor U2784 (N_2784,In_3990,In_905);
nor U2785 (N_2785,In_3840,In_3896);
nor U2786 (N_2786,In_4837,In_2666);
nand U2787 (N_2787,In_869,In_2346);
and U2788 (N_2788,In_2641,In_2875);
nand U2789 (N_2789,In_3952,In_4163);
nor U2790 (N_2790,In_3631,In_1463);
nor U2791 (N_2791,In_1145,In_4169);
xnor U2792 (N_2792,In_3554,In_4686);
or U2793 (N_2793,In_4635,In_52);
or U2794 (N_2794,In_2183,In_1177);
xor U2795 (N_2795,In_383,In_3791);
and U2796 (N_2796,In_1180,In_1265);
nand U2797 (N_2797,In_1952,In_4222);
nor U2798 (N_2798,In_3394,In_3929);
and U2799 (N_2799,In_829,In_1215);
xor U2800 (N_2800,In_403,In_3249);
or U2801 (N_2801,In_1621,In_3965);
or U2802 (N_2802,In_1650,In_4465);
or U2803 (N_2803,In_968,In_3256);
nand U2804 (N_2804,In_844,In_3124);
nor U2805 (N_2805,In_210,In_132);
nand U2806 (N_2806,In_1286,In_566);
nand U2807 (N_2807,In_1076,In_3794);
xor U2808 (N_2808,In_1344,In_3120);
nand U2809 (N_2809,In_2473,In_4858);
nand U2810 (N_2810,In_1014,In_3494);
nand U2811 (N_2811,In_2533,In_2132);
nor U2812 (N_2812,In_4024,In_4160);
or U2813 (N_2813,In_2341,In_3008);
or U2814 (N_2814,In_1635,In_4085);
and U2815 (N_2815,In_3845,In_1620);
xor U2816 (N_2816,In_2105,In_3103);
and U2817 (N_2817,In_2818,In_2975);
nor U2818 (N_2818,In_2405,In_4773);
and U2819 (N_2819,In_770,In_717);
or U2820 (N_2820,In_1762,In_1955);
xnor U2821 (N_2821,In_625,In_3451);
xor U2822 (N_2822,In_2276,In_113);
or U2823 (N_2823,In_4455,In_3468);
xnor U2824 (N_2824,In_4157,In_87);
xnor U2825 (N_2825,In_2136,In_4264);
xnor U2826 (N_2826,In_159,In_1455);
xor U2827 (N_2827,In_369,In_1343);
nand U2828 (N_2828,In_522,In_273);
nor U2829 (N_2829,In_268,In_210);
and U2830 (N_2830,In_2792,In_4122);
nand U2831 (N_2831,In_977,In_3464);
or U2832 (N_2832,In_4542,In_2834);
xnor U2833 (N_2833,In_2876,In_1469);
and U2834 (N_2834,In_1380,In_4426);
nand U2835 (N_2835,In_1513,In_1846);
and U2836 (N_2836,In_1465,In_567);
nor U2837 (N_2837,In_3349,In_3390);
nor U2838 (N_2838,In_4002,In_4551);
nand U2839 (N_2839,In_3260,In_3241);
nand U2840 (N_2840,In_3732,In_3022);
nor U2841 (N_2841,In_2106,In_2466);
xnor U2842 (N_2842,In_3597,In_1667);
xnor U2843 (N_2843,In_3032,In_4814);
xnor U2844 (N_2844,In_3129,In_1080);
xor U2845 (N_2845,In_4139,In_2619);
xor U2846 (N_2846,In_1452,In_269);
or U2847 (N_2847,In_2848,In_3179);
nand U2848 (N_2848,In_122,In_790);
and U2849 (N_2849,In_3879,In_108);
or U2850 (N_2850,In_4675,In_1321);
xor U2851 (N_2851,In_1846,In_3276);
and U2852 (N_2852,In_2937,In_495);
nand U2853 (N_2853,In_564,In_1366);
nor U2854 (N_2854,In_3592,In_2384);
and U2855 (N_2855,In_631,In_738);
nor U2856 (N_2856,In_625,In_1991);
nand U2857 (N_2857,In_4547,In_1518);
xnor U2858 (N_2858,In_1841,In_2805);
nand U2859 (N_2859,In_1013,In_3054);
xnor U2860 (N_2860,In_1085,In_4460);
nor U2861 (N_2861,In_1751,In_1195);
and U2862 (N_2862,In_4509,In_2068);
nand U2863 (N_2863,In_109,In_1192);
nand U2864 (N_2864,In_1833,In_4385);
and U2865 (N_2865,In_2271,In_2746);
and U2866 (N_2866,In_690,In_4254);
xnor U2867 (N_2867,In_1432,In_410);
nor U2868 (N_2868,In_669,In_221);
nand U2869 (N_2869,In_4937,In_4688);
xor U2870 (N_2870,In_4192,In_4213);
or U2871 (N_2871,In_3667,In_712);
nor U2872 (N_2872,In_4484,In_2757);
nor U2873 (N_2873,In_1558,In_982);
nor U2874 (N_2874,In_4232,In_3437);
nor U2875 (N_2875,In_2212,In_829);
nor U2876 (N_2876,In_2179,In_2635);
nand U2877 (N_2877,In_2046,In_598);
nor U2878 (N_2878,In_287,In_3185);
xor U2879 (N_2879,In_2159,In_113);
nor U2880 (N_2880,In_3404,In_472);
nor U2881 (N_2881,In_77,In_2706);
nor U2882 (N_2882,In_2207,In_884);
nand U2883 (N_2883,In_4081,In_4717);
xor U2884 (N_2884,In_753,In_3957);
xor U2885 (N_2885,In_4034,In_3323);
or U2886 (N_2886,In_1045,In_99);
or U2887 (N_2887,In_4174,In_3579);
and U2888 (N_2888,In_1693,In_2395);
or U2889 (N_2889,In_3226,In_4257);
and U2890 (N_2890,In_2604,In_124);
nand U2891 (N_2891,In_313,In_1701);
nor U2892 (N_2892,In_351,In_3285);
and U2893 (N_2893,In_1275,In_1155);
nand U2894 (N_2894,In_1351,In_2686);
nor U2895 (N_2895,In_367,In_204);
xnor U2896 (N_2896,In_3591,In_2744);
and U2897 (N_2897,In_1175,In_853);
nand U2898 (N_2898,In_4436,In_3958);
nand U2899 (N_2899,In_2694,In_500);
nand U2900 (N_2900,In_121,In_2702);
and U2901 (N_2901,In_2420,In_2827);
and U2902 (N_2902,In_4449,In_2299);
xnor U2903 (N_2903,In_4112,In_688);
or U2904 (N_2904,In_3350,In_3883);
or U2905 (N_2905,In_3944,In_4352);
and U2906 (N_2906,In_817,In_4478);
or U2907 (N_2907,In_4790,In_2323);
or U2908 (N_2908,In_4330,In_4450);
nor U2909 (N_2909,In_1005,In_2425);
nor U2910 (N_2910,In_565,In_214);
or U2911 (N_2911,In_1812,In_2402);
nand U2912 (N_2912,In_2243,In_621);
xor U2913 (N_2913,In_1258,In_1071);
nand U2914 (N_2914,In_3443,In_3952);
nor U2915 (N_2915,In_1200,In_1763);
or U2916 (N_2916,In_354,In_2122);
xor U2917 (N_2917,In_2095,In_4098);
and U2918 (N_2918,In_2550,In_4056);
or U2919 (N_2919,In_949,In_3143);
nand U2920 (N_2920,In_119,In_720);
nand U2921 (N_2921,In_1359,In_2397);
nand U2922 (N_2922,In_605,In_596);
nor U2923 (N_2923,In_768,In_4775);
xnor U2924 (N_2924,In_892,In_1750);
and U2925 (N_2925,In_125,In_4407);
and U2926 (N_2926,In_3518,In_3647);
or U2927 (N_2927,In_2424,In_282);
xor U2928 (N_2928,In_1911,In_3361);
or U2929 (N_2929,In_196,In_4349);
nor U2930 (N_2930,In_4289,In_3137);
and U2931 (N_2931,In_1041,In_2513);
or U2932 (N_2932,In_2325,In_3685);
nor U2933 (N_2933,In_3261,In_4599);
nor U2934 (N_2934,In_1921,In_4431);
nor U2935 (N_2935,In_4421,In_179);
nor U2936 (N_2936,In_3630,In_4409);
nor U2937 (N_2937,In_515,In_2311);
or U2938 (N_2938,In_1863,In_3581);
xnor U2939 (N_2939,In_373,In_3778);
nor U2940 (N_2940,In_103,In_1957);
and U2941 (N_2941,In_1528,In_872);
nor U2942 (N_2942,In_108,In_1407);
or U2943 (N_2943,In_2344,In_4760);
nor U2944 (N_2944,In_4416,In_2978);
xnor U2945 (N_2945,In_3343,In_343);
xor U2946 (N_2946,In_4338,In_143);
xor U2947 (N_2947,In_4488,In_3192);
or U2948 (N_2948,In_2253,In_122);
xnor U2949 (N_2949,In_4746,In_2208);
and U2950 (N_2950,In_2792,In_3435);
xnor U2951 (N_2951,In_4990,In_1105);
nor U2952 (N_2952,In_572,In_2528);
and U2953 (N_2953,In_1927,In_1362);
nor U2954 (N_2954,In_2525,In_1112);
nor U2955 (N_2955,In_3106,In_2496);
or U2956 (N_2956,In_255,In_192);
and U2957 (N_2957,In_1170,In_1319);
nor U2958 (N_2958,In_202,In_2544);
and U2959 (N_2959,In_1385,In_8);
nor U2960 (N_2960,In_1638,In_948);
and U2961 (N_2961,In_4899,In_617);
nand U2962 (N_2962,In_2332,In_674);
nor U2963 (N_2963,In_667,In_1728);
and U2964 (N_2964,In_186,In_61);
nand U2965 (N_2965,In_90,In_2601);
nor U2966 (N_2966,In_1599,In_45);
nor U2967 (N_2967,In_958,In_2749);
xor U2968 (N_2968,In_1071,In_4037);
nand U2969 (N_2969,In_3446,In_85);
xnor U2970 (N_2970,In_4955,In_3115);
xor U2971 (N_2971,In_4120,In_2612);
and U2972 (N_2972,In_1197,In_221);
nand U2973 (N_2973,In_4984,In_3025);
nor U2974 (N_2974,In_1228,In_4938);
xnor U2975 (N_2975,In_4802,In_1294);
and U2976 (N_2976,In_71,In_578);
nor U2977 (N_2977,In_2597,In_1321);
or U2978 (N_2978,In_3227,In_293);
xnor U2979 (N_2979,In_1635,In_579);
xnor U2980 (N_2980,In_4056,In_3307);
and U2981 (N_2981,In_2446,In_2905);
xor U2982 (N_2982,In_2251,In_1233);
or U2983 (N_2983,In_2839,In_1667);
and U2984 (N_2984,In_1322,In_1833);
nand U2985 (N_2985,In_1770,In_1654);
and U2986 (N_2986,In_116,In_3998);
xor U2987 (N_2987,In_1939,In_4468);
nor U2988 (N_2988,In_2792,In_1472);
or U2989 (N_2989,In_3099,In_4710);
xnor U2990 (N_2990,In_1526,In_1639);
nand U2991 (N_2991,In_4015,In_2915);
nand U2992 (N_2992,In_3801,In_2045);
or U2993 (N_2993,In_3587,In_2743);
and U2994 (N_2994,In_3644,In_2961);
and U2995 (N_2995,In_3021,In_1303);
xnor U2996 (N_2996,In_3137,In_3316);
xnor U2997 (N_2997,In_3253,In_101);
nor U2998 (N_2998,In_2607,In_1053);
xor U2999 (N_2999,In_4222,In_2518);
and U3000 (N_3000,In_3845,In_3628);
xnor U3001 (N_3001,In_74,In_2346);
nor U3002 (N_3002,In_3026,In_2742);
nand U3003 (N_3003,In_676,In_2563);
and U3004 (N_3004,In_50,In_326);
xnor U3005 (N_3005,In_2177,In_3563);
and U3006 (N_3006,In_1223,In_779);
or U3007 (N_3007,In_746,In_3902);
xnor U3008 (N_3008,In_425,In_4429);
xnor U3009 (N_3009,In_1190,In_795);
and U3010 (N_3010,In_1900,In_3515);
xnor U3011 (N_3011,In_3082,In_2754);
xor U3012 (N_3012,In_3716,In_642);
nor U3013 (N_3013,In_4896,In_3428);
and U3014 (N_3014,In_2995,In_2190);
and U3015 (N_3015,In_109,In_3479);
nand U3016 (N_3016,In_4191,In_1848);
and U3017 (N_3017,In_3189,In_775);
nand U3018 (N_3018,In_4156,In_4853);
and U3019 (N_3019,In_3665,In_1281);
or U3020 (N_3020,In_3034,In_4270);
nand U3021 (N_3021,In_35,In_3000);
xor U3022 (N_3022,In_1437,In_3223);
and U3023 (N_3023,In_617,In_3835);
or U3024 (N_3024,In_3469,In_4110);
or U3025 (N_3025,In_3648,In_2617);
and U3026 (N_3026,In_3746,In_3826);
xor U3027 (N_3027,In_1340,In_3833);
xnor U3028 (N_3028,In_4180,In_2462);
nor U3029 (N_3029,In_3667,In_295);
and U3030 (N_3030,In_1918,In_4458);
or U3031 (N_3031,In_3062,In_2212);
and U3032 (N_3032,In_1721,In_1190);
nor U3033 (N_3033,In_946,In_4598);
nand U3034 (N_3034,In_1332,In_1757);
or U3035 (N_3035,In_3149,In_4931);
nand U3036 (N_3036,In_4874,In_2290);
nand U3037 (N_3037,In_840,In_4914);
and U3038 (N_3038,In_2463,In_917);
and U3039 (N_3039,In_1056,In_2103);
and U3040 (N_3040,In_147,In_3764);
and U3041 (N_3041,In_3967,In_4702);
or U3042 (N_3042,In_4533,In_4885);
nor U3043 (N_3043,In_652,In_1313);
nor U3044 (N_3044,In_1685,In_1293);
or U3045 (N_3045,In_1093,In_898);
and U3046 (N_3046,In_4528,In_4626);
and U3047 (N_3047,In_3124,In_493);
and U3048 (N_3048,In_2084,In_3595);
nor U3049 (N_3049,In_3159,In_1456);
nor U3050 (N_3050,In_2526,In_1527);
or U3051 (N_3051,In_1646,In_2590);
or U3052 (N_3052,In_1901,In_4600);
nor U3053 (N_3053,In_3277,In_362);
nor U3054 (N_3054,In_475,In_3857);
nand U3055 (N_3055,In_1988,In_3431);
nor U3056 (N_3056,In_4408,In_2169);
and U3057 (N_3057,In_3196,In_2774);
xor U3058 (N_3058,In_4025,In_3458);
or U3059 (N_3059,In_483,In_2823);
nand U3060 (N_3060,In_42,In_4999);
nor U3061 (N_3061,In_819,In_3220);
xnor U3062 (N_3062,In_3262,In_4220);
xnor U3063 (N_3063,In_622,In_86);
or U3064 (N_3064,In_2560,In_1135);
xnor U3065 (N_3065,In_2004,In_82);
nand U3066 (N_3066,In_416,In_739);
or U3067 (N_3067,In_1341,In_2262);
xnor U3068 (N_3068,In_2984,In_3279);
xor U3069 (N_3069,In_4486,In_829);
nor U3070 (N_3070,In_4715,In_1178);
and U3071 (N_3071,In_4496,In_618);
nand U3072 (N_3072,In_3097,In_3860);
nor U3073 (N_3073,In_751,In_1099);
xnor U3074 (N_3074,In_1739,In_3443);
and U3075 (N_3075,In_3497,In_3894);
xnor U3076 (N_3076,In_4755,In_2163);
nor U3077 (N_3077,In_4638,In_952);
nor U3078 (N_3078,In_1706,In_149);
nand U3079 (N_3079,In_4836,In_833);
nor U3080 (N_3080,In_2225,In_2254);
or U3081 (N_3081,In_3199,In_4214);
nor U3082 (N_3082,In_550,In_2848);
and U3083 (N_3083,In_490,In_3261);
xnor U3084 (N_3084,In_4309,In_4489);
and U3085 (N_3085,In_4208,In_4803);
nand U3086 (N_3086,In_3568,In_1877);
and U3087 (N_3087,In_1184,In_774);
nor U3088 (N_3088,In_4682,In_3663);
and U3089 (N_3089,In_2877,In_234);
nand U3090 (N_3090,In_3565,In_4599);
or U3091 (N_3091,In_1605,In_607);
nor U3092 (N_3092,In_3208,In_4086);
xnor U3093 (N_3093,In_351,In_353);
and U3094 (N_3094,In_2049,In_1719);
nand U3095 (N_3095,In_3059,In_4454);
or U3096 (N_3096,In_4880,In_123);
or U3097 (N_3097,In_2666,In_3787);
xnor U3098 (N_3098,In_1799,In_1512);
xor U3099 (N_3099,In_1716,In_4585);
nand U3100 (N_3100,In_4471,In_910);
nand U3101 (N_3101,In_4013,In_3596);
nand U3102 (N_3102,In_4791,In_3304);
or U3103 (N_3103,In_624,In_1769);
nand U3104 (N_3104,In_4750,In_3761);
nand U3105 (N_3105,In_4225,In_4258);
or U3106 (N_3106,In_169,In_1992);
nand U3107 (N_3107,In_4764,In_3280);
xor U3108 (N_3108,In_3863,In_17);
and U3109 (N_3109,In_3273,In_2445);
and U3110 (N_3110,In_2135,In_4848);
nand U3111 (N_3111,In_2035,In_3838);
or U3112 (N_3112,In_955,In_2802);
xnor U3113 (N_3113,In_1746,In_4720);
and U3114 (N_3114,In_3474,In_563);
and U3115 (N_3115,In_2631,In_429);
or U3116 (N_3116,In_818,In_4727);
and U3117 (N_3117,In_1304,In_3582);
and U3118 (N_3118,In_1984,In_4220);
and U3119 (N_3119,In_4880,In_606);
xnor U3120 (N_3120,In_2624,In_74);
nor U3121 (N_3121,In_1719,In_4396);
nand U3122 (N_3122,In_2973,In_3625);
nor U3123 (N_3123,In_1722,In_1733);
xor U3124 (N_3124,In_3138,In_3241);
nand U3125 (N_3125,In_2545,In_3359);
or U3126 (N_3126,In_858,In_2499);
nor U3127 (N_3127,In_2874,In_225);
and U3128 (N_3128,In_3427,In_3621);
nor U3129 (N_3129,In_3412,In_3040);
nand U3130 (N_3130,In_2016,In_513);
nand U3131 (N_3131,In_4751,In_292);
and U3132 (N_3132,In_585,In_3920);
nor U3133 (N_3133,In_1349,In_2599);
nor U3134 (N_3134,In_3603,In_4836);
and U3135 (N_3135,In_4436,In_3586);
and U3136 (N_3136,In_3872,In_4362);
nand U3137 (N_3137,In_769,In_3792);
xor U3138 (N_3138,In_2137,In_24);
or U3139 (N_3139,In_4436,In_4434);
or U3140 (N_3140,In_4739,In_3629);
nand U3141 (N_3141,In_327,In_742);
nand U3142 (N_3142,In_4228,In_2443);
nor U3143 (N_3143,In_535,In_625);
xnor U3144 (N_3144,In_1015,In_1641);
nand U3145 (N_3145,In_3447,In_2189);
nor U3146 (N_3146,In_288,In_244);
or U3147 (N_3147,In_348,In_40);
and U3148 (N_3148,In_3649,In_10);
nor U3149 (N_3149,In_1945,In_2384);
or U3150 (N_3150,In_3139,In_4662);
xor U3151 (N_3151,In_3771,In_1212);
nor U3152 (N_3152,In_1769,In_2345);
nor U3153 (N_3153,In_326,In_4256);
xor U3154 (N_3154,In_3780,In_893);
or U3155 (N_3155,In_3056,In_3965);
nor U3156 (N_3156,In_2484,In_3358);
xnor U3157 (N_3157,In_2519,In_4010);
nand U3158 (N_3158,In_2250,In_1872);
xor U3159 (N_3159,In_1668,In_2572);
and U3160 (N_3160,In_4815,In_3688);
xnor U3161 (N_3161,In_2511,In_2233);
nor U3162 (N_3162,In_3070,In_3106);
nor U3163 (N_3163,In_281,In_2356);
or U3164 (N_3164,In_4138,In_386);
xnor U3165 (N_3165,In_1970,In_4659);
or U3166 (N_3166,In_2110,In_3032);
nand U3167 (N_3167,In_3555,In_4127);
nand U3168 (N_3168,In_4821,In_3157);
nor U3169 (N_3169,In_757,In_2449);
and U3170 (N_3170,In_1542,In_1870);
and U3171 (N_3171,In_4666,In_3730);
nor U3172 (N_3172,In_624,In_2846);
nor U3173 (N_3173,In_418,In_2659);
xnor U3174 (N_3174,In_1496,In_1488);
or U3175 (N_3175,In_3558,In_900);
nand U3176 (N_3176,In_4445,In_3855);
or U3177 (N_3177,In_4637,In_3801);
nor U3178 (N_3178,In_1231,In_4264);
nand U3179 (N_3179,In_4843,In_2754);
and U3180 (N_3180,In_1381,In_3148);
and U3181 (N_3181,In_4584,In_746);
nand U3182 (N_3182,In_3496,In_3021);
xnor U3183 (N_3183,In_374,In_2403);
nor U3184 (N_3184,In_2700,In_4748);
xor U3185 (N_3185,In_4930,In_2014);
nor U3186 (N_3186,In_3118,In_1239);
nand U3187 (N_3187,In_3981,In_2521);
or U3188 (N_3188,In_2522,In_4145);
and U3189 (N_3189,In_2167,In_1256);
nor U3190 (N_3190,In_4906,In_3542);
or U3191 (N_3191,In_674,In_1842);
or U3192 (N_3192,In_2106,In_4935);
nor U3193 (N_3193,In_1388,In_3167);
xnor U3194 (N_3194,In_397,In_3130);
and U3195 (N_3195,In_4240,In_4096);
nor U3196 (N_3196,In_1177,In_4186);
or U3197 (N_3197,In_2695,In_3272);
and U3198 (N_3198,In_1359,In_414);
nor U3199 (N_3199,In_3122,In_4245);
nand U3200 (N_3200,In_4910,In_947);
or U3201 (N_3201,In_4557,In_2699);
xor U3202 (N_3202,In_1527,In_3765);
or U3203 (N_3203,In_2875,In_2332);
or U3204 (N_3204,In_4098,In_2703);
xnor U3205 (N_3205,In_1760,In_4052);
xnor U3206 (N_3206,In_4149,In_943);
nand U3207 (N_3207,In_3008,In_3403);
nor U3208 (N_3208,In_1126,In_3189);
nor U3209 (N_3209,In_1283,In_1504);
xnor U3210 (N_3210,In_3989,In_1883);
and U3211 (N_3211,In_3147,In_2060);
xnor U3212 (N_3212,In_1130,In_2257);
or U3213 (N_3213,In_4670,In_1308);
nand U3214 (N_3214,In_2575,In_3705);
nor U3215 (N_3215,In_3685,In_799);
or U3216 (N_3216,In_4652,In_4850);
xnor U3217 (N_3217,In_4306,In_649);
nor U3218 (N_3218,In_3353,In_1989);
nand U3219 (N_3219,In_4233,In_4349);
nand U3220 (N_3220,In_3957,In_2461);
nand U3221 (N_3221,In_4141,In_3233);
or U3222 (N_3222,In_3125,In_4445);
and U3223 (N_3223,In_4709,In_2650);
and U3224 (N_3224,In_686,In_2336);
xnor U3225 (N_3225,In_107,In_4341);
and U3226 (N_3226,In_4782,In_3523);
nand U3227 (N_3227,In_4298,In_664);
nand U3228 (N_3228,In_3132,In_1834);
nand U3229 (N_3229,In_3643,In_1426);
nand U3230 (N_3230,In_2144,In_3449);
nand U3231 (N_3231,In_3334,In_1278);
nand U3232 (N_3232,In_466,In_2412);
or U3233 (N_3233,In_41,In_1372);
or U3234 (N_3234,In_2350,In_381);
or U3235 (N_3235,In_3506,In_3617);
and U3236 (N_3236,In_4342,In_191);
and U3237 (N_3237,In_4723,In_1722);
xnor U3238 (N_3238,In_2500,In_1326);
nand U3239 (N_3239,In_2504,In_2148);
nand U3240 (N_3240,In_3306,In_2206);
or U3241 (N_3241,In_2233,In_224);
nand U3242 (N_3242,In_1624,In_4213);
or U3243 (N_3243,In_3590,In_150);
nor U3244 (N_3244,In_2069,In_4063);
nor U3245 (N_3245,In_2410,In_1550);
or U3246 (N_3246,In_1761,In_4855);
or U3247 (N_3247,In_4900,In_4458);
or U3248 (N_3248,In_2124,In_1149);
nand U3249 (N_3249,In_4528,In_2610);
and U3250 (N_3250,In_4524,In_2964);
nand U3251 (N_3251,In_1456,In_3323);
nand U3252 (N_3252,In_267,In_3068);
xor U3253 (N_3253,In_1482,In_4114);
nand U3254 (N_3254,In_3139,In_1226);
nand U3255 (N_3255,In_2573,In_4720);
or U3256 (N_3256,In_3006,In_2917);
or U3257 (N_3257,In_2026,In_999);
or U3258 (N_3258,In_3483,In_1051);
nand U3259 (N_3259,In_2162,In_105);
xor U3260 (N_3260,In_1606,In_3620);
xor U3261 (N_3261,In_860,In_2989);
xnor U3262 (N_3262,In_668,In_1940);
nand U3263 (N_3263,In_54,In_601);
or U3264 (N_3264,In_3445,In_4082);
nor U3265 (N_3265,In_2099,In_4446);
and U3266 (N_3266,In_2436,In_1832);
and U3267 (N_3267,In_2330,In_3350);
nand U3268 (N_3268,In_993,In_3690);
or U3269 (N_3269,In_3411,In_2624);
xor U3270 (N_3270,In_4677,In_3182);
or U3271 (N_3271,In_2689,In_3941);
nor U3272 (N_3272,In_61,In_2478);
nand U3273 (N_3273,In_350,In_3643);
nand U3274 (N_3274,In_4803,In_4502);
and U3275 (N_3275,In_4843,In_8);
xnor U3276 (N_3276,In_3994,In_1912);
nand U3277 (N_3277,In_2621,In_1169);
xnor U3278 (N_3278,In_4419,In_417);
xor U3279 (N_3279,In_4712,In_3409);
nand U3280 (N_3280,In_3008,In_1024);
nor U3281 (N_3281,In_370,In_4407);
nor U3282 (N_3282,In_4894,In_2708);
nand U3283 (N_3283,In_4940,In_2541);
and U3284 (N_3284,In_1590,In_2682);
xnor U3285 (N_3285,In_3392,In_4472);
or U3286 (N_3286,In_2339,In_4183);
or U3287 (N_3287,In_4050,In_1862);
nand U3288 (N_3288,In_3276,In_4203);
nor U3289 (N_3289,In_4165,In_408);
or U3290 (N_3290,In_2288,In_4996);
nand U3291 (N_3291,In_2148,In_12);
nand U3292 (N_3292,In_844,In_4591);
and U3293 (N_3293,In_3536,In_3725);
or U3294 (N_3294,In_4785,In_1464);
and U3295 (N_3295,In_3546,In_2930);
nand U3296 (N_3296,In_2413,In_3956);
and U3297 (N_3297,In_2640,In_2903);
nor U3298 (N_3298,In_799,In_2292);
nor U3299 (N_3299,In_2061,In_2539);
or U3300 (N_3300,In_2871,In_3550);
xor U3301 (N_3301,In_2047,In_607);
and U3302 (N_3302,In_4059,In_4364);
xor U3303 (N_3303,In_724,In_1463);
and U3304 (N_3304,In_1026,In_1519);
nand U3305 (N_3305,In_2101,In_3112);
nand U3306 (N_3306,In_3261,In_4864);
xnor U3307 (N_3307,In_3658,In_3703);
nor U3308 (N_3308,In_3123,In_1882);
nor U3309 (N_3309,In_3068,In_4173);
and U3310 (N_3310,In_2719,In_2316);
nand U3311 (N_3311,In_2002,In_2407);
xor U3312 (N_3312,In_639,In_4240);
xnor U3313 (N_3313,In_4497,In_3482);
xor U3314 (N_3314,In_3639,In_63);
or U3315 (N_3315,In_1885,In_3176);
or U3316 (N_3316,In_3665,In_3414);
or U3317 (N_3317,In_2562,In_4232);
nand U3318 (N_3318,In_4072,In_2137);
xnor U3319 (N_3319,In_3636,In_1170);
xnor U3320 (N_3320,In_4888,In_4724);
nand U3321 (N_3321,In_1239,In_3457);
and U3322 (N_3322,In_2508,In_2028);
nor U3323 (N_3323,In_3376,In_4616);
and U3324 (N_3324,In_717,In_142);
or U3325 (N_3325,In_4584,In_4242);
and U3326 (N_3326,In_4005,In_4266);
or U3327 (N_3327,In_3649,In_4134);
nand U3328 (N_3328,In_1018,In_3374);
nand U3329 (N_3329,In_3216,In_3676);
xnor U3330 (N_3330,In_2732,In_3175);
or U3331 (N_3331,In_1800,In_4918);
xor U3332 (N_3332,In_704,In_3589);
nand U3333 (N_3333,In_1310,In_4191);
nor U3334 (N_3334,In_347,In_2608);
and U3335 (N_3335,In_3579,In_704);
nor U3336 (N_3336,In_4875,In_1303);
nor U3337 (N_3337,In_1098,In_1502);
and U3338 (N_3338,In_1512,In_1989);
xor U3339 (N_3339,In_360,In_482);
and U3340 (N_3340,In_193,In_1015);
nand U3341 (N_3341,In_456,In_2135);
xnor U3342 (N_3342,In_3378,In_2020);
nor U3343 (N_3343,In_2086,In_4247);
nor U3344 (N_3344,In_0,In_712);
or U3345 (N_3345,In_762,In_3183);
or U3346 (N_3346,In_4036,In_1873);
and U3347 (N_3347,In_2454,In_913);
xor U3348 (N_3348,In_1264,In_1969);
and U3349 (N_3349,In_4595,In_1153);
or U3350 (N_3350,In_667,In_2052);
and U3351 (N_3351,In_2692,In_4030);
nor U3352 (N_3352,In_2709,In_903);
xnor U3353 (N_3353,In_4107,In_2281);
nand U3354 (N_3354,In_1804,In_4726);
xor U3355 (N_3355,In_1939,In_1174);
nand U3356 (N_3356,In_329,In_3899);
or U3357 (N_3357,In_1220,In_3919);
xor U3358 (N_3358,In_275,In_1384);
nor U3359 (N_3359,In_3849,In_1284);
nand U3360 (N_3360,In_2752,In_4433);
and U3361 (N_3361,In_1144,In_1724);
nor U3362 (N_3362,In_2617,In_2557);
nand U3363 (N_3363,In_347,In_2175);
nand U3364 (N_3364,In_343,In_4922);
nor U3365 (N_3365,In_550,In_456);
nand U3366 (N_3366,In_3678,In_3654);
nand U3367 (N_3367,In_3439,In_3460);
xor U3368 (N_3368,In_3927,In_1919);
xnor U3369 (N_3369,In_4239,In_1658);
xnor U3370 (N_3370,In_1228,In_2195);
xor U3371 (N_3371,In_655,In_3568);
xnor U3372 (N_3372,In_2477,In_2326);
nand U3373 (N_3373,In_1160,In_3887);
xor U3374 (N_3374,In_2741,In_2259);
or U3375 (N_3375,In_4029,In_1940);
or U3376 (N_3376,In_156,In_1215);
xnor U3377 (N_3377,In_3834,In_1471);
and U3378 (N_3378,In_4997,In_2239);
xor U3379 (N_3379,In_4919,In_4004);
and U3380 (N_3380,In_4582,In_976);
nor U3381 (N_3381,In_1807,In_1179);
or U3382 (N_3382,In_1840,In_3242);
or U3383 (N_3383,In_683,In_2369);
nor U3384 (N_3384,In_4904,In_2466);
nand U3385 (N_3385,In_2484,In_1171);
nand U3386 (N_3386,In_4271,In_3816);
nor U3387 (N_3387,In_1783,In_2079);
xnor U3388 (N_3388,In_3931,In_2052);
nand U3389 (N_3389,In_574,In_3743);
and U3390 (N_3390,In_1646,In_1137);
nand U3391 (N_3391,In_4789,In_4326);
or U3392 (N_3392,In_2755,In_185);
nand U3393 (N_3393,In_1253,In_3219);
and U3394 (N_3394,In_2763,In_1414);
xor U3395 (N_3395,In_3386,In_2692);
nor U3396 (N_3396,In_2495,In_3260);
nor U3397 (N_3397,In_2253,In_3565);
and U3398 (N_3398,In_331,In_101);
and U3399 (N_3399,In_3569,In_3793);
nor U3400 (N_3400,In_4032,In_3803);
nand U3401 (N_3401,In_3146,In_296);
nor U3402 (N_3402,In_3848,In_3145);
and U3403 (N_3403,In_1529,In_4444);
or U3404 (N_3404,In_4829,In_3528);
or U3405 (N_3405,In_1262,In_3365);
nor U3406 (N_3406,In_1815,In_925);
and U3407 (N_3407,In_448,In_4961);
and U3408 (N_3408,In_4807,In_131);
nand U3409 (N_3409,In_113,In_591);
xor U3410 (N_3410,In_3241,In_1351);
or U3411 (N_3411,In_2284,In_3402);
nor U3412 (N_3412,In_4337,In_722);
or U3413 (N_3413,In_4296,In_2109);
xnor U3414 (N_3414,In_2676,In_4242);
nor U3415 (N_3415,In_2387,In_3509);
xnor U3416 (N_3416,In_4874,In_3643);
nor U3417 (N_3417,In_396,In_2177);
and U3418 (N_3418,In_1912,In_23);
nand U3419 (N_3419,In_51,In_1699);
nor U3420 (N_3420,In_1654,In_589);
nand U3421 (N_3421,In_1567,In_4743);
or U3422 (N_3422,In_3301,In_94);
or U3423 (N_3423,In_4144,In_3741);
nor U3424 (N_3424,In_1856,In_3863);
or U3425 (N_3425,In_1500,In_2609);
or U3426 (N_3426,In_2675,In_1466);
or U3427 (N_3427,In_1371,In_2521);
and U3428 (N_3428,In_312,In_1385);
xor U3429 (N_3429,In_3723,In_3332);
or U3430 (N_3430,In_2000,In_4390);
xnor U3431 (N_3431,In_2263,In_4776);
nand U3432 (N_3432,In_2179,In_2399);
or U3433 (N_3433,In_4801,In_1713);
and U3434 (N_3434,In_3984,In_1675);
and U3435 (N_3435,In_1328,In_2264);
or U3436 (N_3436,In_3390,In_2247);
nand U3437 (N_3437,In_2080,In_1101);
xor U3438 (N_3438,In_4205,In_2508);
nor U3439 (N_3439,In_100,In_1266);
and U3440 (N_3440,In_683,In_916);
xnor U3441 (N_3441,In_1391,In_1090);
or U3442 (N_3442,In_2213,In_4916);
or U3443 (N_3443,In_797,In_3876);
xor U3444 (N_3444,In_4849,In_2179);
or U3445 (N_3445,In_2929,In_3913);
or U3446 (N_3446,In_724,In_1280);
or U3447 (N_3447,In_306,In_926);
nor U3448 (N_3448,In_1892,In_3212);
nor U3449 (N_3449,In_1145,In_2716);
and U3450 (N_3450,In_843,In_115);
and U3451 (N_3451,In_3811,In_395);
and U3452 (N_3452,In_2667,In_3078);
nor U3453 (N_3453,In_1669,In_469);
xor U3454 (N_3454,In_888,In_228);
or U3455 (N_3455,In_4833,In_1222);
nor U3456 (N_3456,In_3266,In_4903);
xnor U3457 (N_3457,In_4716,In_1272);
nor U3458 (N_3458,In_1182,In_127);
nor U3459 (N_3459,In_3219,In_1267);
nand U3460 (N_3460,In_4361,In_4104);
nand U3461 (N_3461,In_3210,In_2440);
and U3462 (N_3462,In_795,In_722);
nor U3463 (N_3463,In_3311,In_1200);
and U3464 (N_3464,In_2705,In_4504);
nand U3465 (N_3465,In_4708,In_4935);
nor U3466 (N_3466,In_3266,In_863);
and U3467 (N_3467,In_2839,In_4688);
nand U3468 (N_3468,In_3751,In_3681);
nand U3469 (N_3469,In_4968,In_4262);
xnor U3470 (N_3470,In_3118,In_4362);
and U3471 (N_3471,In_3885,In_1540);
nand U3472 (N_3472,In_4151,In_3483);
and U3473 (N_3473,In_220,In_2398);
xor U3474 (N_3474,In_3664,In_2331);
nand U3475 (N_3475,In_2317,In_3823);
or U3476 (N_3476,In_4476,In_4969);
xnor U3477 (N_3477,In_2072,In_1604);
and U3478 (N_3478,In_2570,In_2614);
and U3479 (N_3479,In_1654,In_1071);
nor U3480 (N_3480,In_1172,In_3194);
and U3481 (N_3481,In_4192,In_342);
nand U3482 (N_3482,In_3717,In_3660);
and U3483 (N_3483,In_2173,In_4195);
nand U3484 (N_3484,In_2898,In_1026);
nand U3485 (N_3485,In_2018,In_2846);
nand U3486 (N_3486,In_4767,In_2387);
nand U3487 (N_3487,In_896,In_586);
nand U3488 (N_3488,In_3260,In_1979);
and U3489 (N_3489,In_3539,In_2462);
nand U3490 (N_3490,In_3000,In_301);
nand U3491 (N_3491,In_1934,In_721);
nand U3492 (N_3492,In_1131,In_131);
or U3493 (N_3493,In_3683,In_1719);
nand U3494 (N_3494,In_4662,In_4735);
or U3495 (N_3495,In_2217,In_1413);
nor U3496 (N_3496,In_3597,In_682);
and U3497 (N_3497,In_3260,In_2373);
and U3498 (N_3498,In_4325,In_3063);
nor U3499 (N_3499,In_1511,In_1380);
and U3500 (N_3500,In_1552,In_3863);
nor U3501 (N_3501,In_2491,In_575);
nand U3502 (N_3502,In_1385,In_4692);
or U3503 (N_3503,In_2994,In_2060);
nor U3504 (N_3504,In_422,In_759);
nand U3505 (N_3505,In_3620,In_3936);
or U3506 (N_3506,In_2738,In_2889);
nand U3507 (N_3507,In_4963,In_347);
nand U3508 (N_3508,In_1407,In_2771);
and U3509 (N_3509,In_4118,In_1475);
nand U3510 (N_3510,In_3088,In_272);
nor U3511 (N_3511,In_236,In_4018);
or U3512 (N_3512,In_2161,In_3369);
or U3513 (N_3513,In_4793,In_677);
nand U3514 (N_3514,In_4769,In_3383);
nand U3515 (N_3515,In_2047,In_2540);
xor U3516 (N_3516,In_4438,In_1493);
or U3517 (N_3517,In_4183,In_3402);
xnor U3518 (N_3518,In_2461,In_4468);
xnor U3519 (N_3519,In_4120,In_720);
xor U3520 (N_3520,In_593,In_1579);
xor U3521 (N_3521,In_3088,In_4514);
xor U3522 (N_3522,In_1459,In_2750);
or U3523 (N_3523,In_2024,In_3851);
or U3524 (N_3524,In_2794,In_3199);
nand U3525 (N_3525,In_912,In_3532);
xor U3526 (N_3526,In_4643,In_3360);
xor U3527 (N_3527,In_3232,In_1377);
nor U3528 (N_3528,In_143,In_3978);
nand U3529 (N_3529,In_2878,In_2216);
nand U3530 (N_3530,In_3983,In_2842);
and U3531 (N_3531,In_1689,In_1774);
nand U3532 (N_3532,In_2433,In_1712);
nand U3533 (N_3533,In_656,In_587);
nor U3534 (N_3534,In_478,In_1486);
nand U3535 (N_3535,In_4886,In_3151);
and U3536 (N_3536,In_3708,In_734);
or U3537 (N_3537,In_2138,In_3159);
xor U3538 (N_3538,In_11,In_1242);
nand U3539 (N_3539,In_3796,In_210);
nand U3540 (N_3540,In_52,In_1338);
or U3541 (N_3541,In_685,In_4816);
xnor U3542 (N_3542,In_1627,In_652);
or U3543 (N_3543,In_366,In_1338);
nor U3544 (N_3544,In_601,In_4744);
and U3545 (N_3545,In_2888,In_3473);
or U3546 (N_3546,In_1973,In_13);
xnor U3547 (N_3547,In_2610,In_823);
nor U3548 (N_3548,In_3257,In_2538);
nand U3549 (N_3549,In_4500,In_1762);
and U3550 (N_3550,In_4636,In_3303);
or U3551 (N_3551,In_585,In_2946);
or U3552 (N_3552,In_966,In_4954);
xnor U3553 (N_3553,In_213,In_3011);
nor U3554 (N_3554,In_1007,In_921);
or U3555 (N_3555,In_4694,In_3877);
nor U3556 (N_3556,In_3952,In_3933);
xnor U3557 (N_3557,In_3512,In_3783);
or U3558 (N_3558,In_2299,In_2960);
nand U3559 (N_3559,In_2431,In_4017);
xor U3560 (N_3560,In_3460,In_2309);
nand U3561 (N_3561,In_619,In_1775);
or U3562 (N_3562,In_2020,In_2508);
nand U3563 (N_3563,In_1628,In_271);
and U3564 (N_3564,In_2079,In_1705);
nand U3565 (N_3565,In_3178,In_1094);
and U3566 (N_3566,In_2086,In_2179);
xor U3567 (N_3567,In_1762,In_3673);
nand U3568 (N_3568,In_287,In_3589);
or U3569 (N_3569,In_55,In_2938);
or U3570 (N_3570,In_863,In_2065);
or U3571 (N_3571,In_3809,In_1883);
and U3572 (N_3572,In_4198,In_4850);
nand U3573 (N_3573,In_3935,In_3969);
nand U3574 (N_3574,In_787,In_1193);
and U3575 (N_3575,In_2544,In_894);
or U3576 (N_3576,In_1374,In_3028);
xnor U3577 (N_3577,In_2586,In_2566);
or U3578 (N_3578,In_810,In_4532);
and U3579 (N_3579,In_2335,In_3702);
nor U3580 (N_3580,In_1062,In_220);
nor U3581 (N_3581,In_240,In_856);
nor U3582 (N_3582,In_4477,In_1899);
nor U3583 (N_3583,In_1195,In_4424);
xor U3584 (N_3584,In_1092,In_2099);
and U3585 (N_3585,In_1987,In_1571);
nand U3586 (N_3586,In_4547,In_824);
nand U3587 (N_3587,In_3517,In_3619);
nor U3588 (N_3588,In_2523,In_4126);
and U3589 (N_3589,In_266,In_3584);
xnor U3590 (N_3590,In_2479,In_4725);
xor U3591 (N_3591,In_2882,In_1817);
nor U3592 (N_3592,In_1695,In_1273);
and U3593 (N_3593,In_2768,In_3920);
nor U3594 (N_3594,In_2722,In_1544);
xnor U3595 (N_3595,In_4918,In_3046);
nor U3596 (N_3596,In_3881,In_4290);
and U3597 (N_3597,In_2901,In_1710);
and U3598 (N_3598,In_2832,In_1868);
nand U3599 (N_3599,In_233,In_3252);
nor U3600 (N_3600,In_315,In_2680);
nand U3601 (N_3601,In_4575,In_483);
or U3602 (N_3602,In_3930,In_2295);
nor U3603 (N_3603,In_2634,In_3777);
nor U3604 (N_3604,In_3478,In_579);
nor U3605 (N_3605,In_1849,In_1857);
nand U3606 (N_3606,In_3634,In_1051);
nor U3607 (N_3607,In_1378,In_3628);
or U3608 (N_3608,In_4821,In_1634);
xor U3609 (N_3609,In_3332,In_642);
nor U3610 (N_3610,In_1888,In_347);
nand U3611 (N_3611,In_2883,In_1080);
and U3612 (N_3612,In_1863,In_1556);
and U3613 (N_3613,In_3726,In_1316);
or U3614 (N_3614,In_4898,In_2028);
or U3615 (N_3615,In_1500,In_179);
nand U3616 (N_3616,In_1476,In_3901);
and U3617 (N_3617,In_4305,In_2908);
and U3618 (N_3618,In_4029,In_1378);
and U3619 (N_3619,In_702,In_1011);
xnor U3620 (N_3620,In_4674,In_3149);
nand U3621 (N_3621,In_794,In_4828);
nor U3622 (N_3622,In_4561,In_699);
nand U3623 (N_3623,In_3707,In_1704);
xor U3624 (N_3624,In_3262,In_1452);
or U3625 (N_3625,In_4859,In_3937);
and U3626 (N_3626,In_197,In_4778);
nor U3627 (N_3627,In_605,In_3102);
xnor U3628 (N_3628,In_1774,In_4007);
and U3629 (N_3629,In_4279,In_647);
nand U3630 (N_3630,In_4120,In_3145);
nor U3631 (N_3631,In_1569,In_1304);
and U3632 (N_3632,In_2351,In_1062);
nand U3633 (N_3633,In_4175,In_4105);
and U3634 (N_3634,In_2469,In_4194);
xnor U3635 (N_3635,In_169,In_1290);
or U3636 (N_3636,In_2031,In_2705);
nor U3637 (N_3637,In_4456,In_573);
nor U3638 (N_3638,In_1927,In_1536);
nor U3639 (N_3639,In_4734,In_3238);
nor U3640 (N_3640,In_4606,In_1603);
and U3641 (N_3641,In_1406,In_1083);
nor U3642 (N_3642,In_656,In_597);
xor U3643 (N_3643,In_3944,In_4915);
nand U3644 (N_3644,In_1930,In_2810);
nand U3645 (N_3645,In_2581,In_3565);
nor U3646 (N_3646,In_4315,In_558);
xor U3647 (N_3647,In_2674,In_876);
or U3648 (N_3648,In_4046,In_973);
xor U3649 (N_3649,In_2782,In_647);
nand U3650 (N_3650,In_1577,In_2103);
xnor U3651 (N_3651,In_4832,In_4044);
nor U3652 (N_3652,In_2481,In_2283);
nor U3653 (N_3653,In_1217,In_4355);
nor U3654 (N_3654,In_842,In_1205);
and U3655 (N_3655,In_1718,In_3530);
and U3656 (N_3656,In_741,In_3321);
and U3657 (N_3657,In_164,In_1823);
nor U3658 (N_3658,In_3860,In_2663);
or U3659 (N_3659,In_514,In_3853);
nor U3660 (N_3660,In_4860,In_416);
nor U3661 (N_3661,In_2857,In_2354);
nor U3662 (N_3662,In_4087,In_1861);
nand U3663 (N_3663,In_1132,In_2163);
xnor U3664 (N_3664,In_1092,In_4470);
or U3665 (N_3665,In_221,In_1034);
nand U3666 (N_3666,In_2004,In_866);
and U3667 (N_3667,In_904,In_821);
nand U3668 (N_3668,In_4463,In_8);
nand U3669 (N_3669,In_2940,In_3928);
xnor U3670 (N_3670,In_3345,In_1876);
nand U3671 (N_3671,In_3236,In_4577);
nand U3672 (N_3672,In_790,In_1997);
xor U3673 (N_3673,In_2822,In_2495);
xnor U3674 (N_3674,In_2896,In_2300);
nor U3675 (N_3675,In_1108,In_239);
nor U3676 (N_3676,In_289,In_552);
or U3677 (N_3677,In_4937,In_2664);
or U3678 (N_3678,In_2371,In_1943);
nor U3679 (N_3679,In_1766,In_378);
nand U3680 (N_3680,In_877,In_4647);
or U3681 (N_3681,In_693,In_2817);
xor U3682 (N_3682,In_3991,In_1914);
or U3683 (N_3683,In_2606,In_18);
nand U3684 (N_3684,In_2046,In_2211);
xor U3685 (N_3685,In_4866,In_4740);
nor U3686 (N_3686,In_4267,In_2658);
nand U3687 (N_3687,In_1445,In_4395);
nand U3688 (N_3688,In_712,In_3848);
nand U3689 (N_3689,In_2087,In_1203);
nand U3690 (N_3690,In_4763,In_2770);
nand U3691 (N_3691,In_4130,In_2434);
xnor U3692 (N_3692,In_4606,In_1613);
nand U3693 (N_3693,In_2598,In_3204);
nand U3694 (N_3694,In_1109,In_1493);
nor U3695 (N_3695,In_4408,In_1255);
and U3696 (N_3696,In_4924,In_3193);
nor U3697 (N_3697,In_949,In_683);
and U3698 (N_3698,In_4029,In_965);
nand U3699 (N_3699,In_3641,In_3162);
nor U3700 (N_3700,In_3696,In_515);
nor U3701 (N_3701,In_540,In_3095);
and U3702 (N_3702,In_3062,In_555);
xnor U3703 (N_3703,In_3492,In_2939);
or U3704 (N_3704,In_2142,In_2320);
and U3705 (N_3705,In_1823,In_4083);
xor U3706 (N_3706,In_633,In_4658);
or U3707 (N_3707,In_805,In_3645);
or U3708 (N_3708,In_2147,In_2968);
nand U3709 (N_3709,In_138,In_2936);
nand U3710 (N_3710,In_681,In_4093);
nor U3711 (N_3711,In_4251,In_3125);
and U3712 (N_3712,In_1967,In_2085);
and U3713 (N_3713,In_560,In_4532);
nor U3714 (N_3714,In_5,In_1736);
nor U3715 (N_3715,In_4831,In_4523);
nand U3716 (N_3716,In_1254,In_3102);
and U3717 (N_3717,In_2645,In_3701);
xnor U3718 (N_3718,In_3203,In_2925);
xnor U3719 (N_3719,In_1533,In_2974);
nand U3720 (N_3720,In_3064,In_806);
and U3721 (N_3721,In_756,In_2505);
nor U3722 (N_3722,In_2372,In_4743);
and U3723 (N_3723,In_276,In_4414);
nor U3724 (N_3724,In_586,In_4934);
nor U3725 (N_3725,In_2671,In_1068);
nor U3726 (N_3726,In_2521,In_3095);
and U3727 (N_3727,In_1930,In_854);
nand U3728 (N_3728,In_2496,In_573);
xor U3729 (N_3729,In_4715,In_2577);
xnor U3730 (N_3730,In_4502,In_4605);
xnor U3731 (N_3731,In_1008,In_497);
or U3732 (N_3732,In_3662,In_1824);
nor U3733 (N_3733,In_3421,In_2805);
nand U3734 (N_3734,In_2921,In_667);
or U3735 (N_3735,In_2258,In_319);
nand U3736 (N_3736,In_4580,In_3872);
or U3737 (N_3737,In_3429,In_3604);
nor U3738 (N_3738,In_3687,In_3301);
nor U3739 (N_3739,In_1401,In_4494);
xnor U3740 (N_3740,In_2399,In_1759);
nand U3741 (N_3741,In_3204,In_2831);
xnor U3742 (N_3742,In_849,In_468);
or U3743 (N_3743,In_4728,In_4298);
xnor U3744 (N_3744,In_1405,In_4436);
nand U3745 (N_3745,In_4374,In_396);
nor U3746 (N_3746,In_4640,In_4837);
or U3747 (N_3747,In_4019,In_343);
and U3748 (N_3748,In_741,In_4884);
or U3749 (N_3749,In_3789,In_2745);
nor U3750 (N_3750,In_2846,In_3772);
or U3751 (N_3751,In_1032,In_4452);
nor U3752 (N_3752,In_2067,In_3825);
nand U3753 (N_3753,In_4146,In_3428);
nand U3754 (N_3754,In_1577,In_1377);
or U3755 (N_3755,In_302,In_2528);
nand U3756 (N_3756,In_3049,In_3147);
xor U3757 (N_3757,In_1002,In_15);
nand U3758 (N_3758,In_2926,In_936);
nand U3759 (N_3759,In_2826,In_4810);
xor U3760 (N_3760,In_2526,In_3265);
nor U3761 (N_3761,In_1044,In_956);
or U3762 (N_3762,In_2569,In_4771);
nor U3763 (N_3763,In_1842,In_989);
nor U3764 (N_3764,In_3248,In_2164);
and U3765 (N_3765,In_748,In_4390);
and U3766 (N_3766,In_2072,In_3454);
nand U3767 (N_3767,In_841,In_1737);
nor U3768 (N_3768,In_781,In_2108);
nor U3769 (N_3769,In_1593,In_4845);
or U3770 (N_3770,In_4898,In_4941);
nand U3771 (N_3771,In_3258,In_837);
and U3772 (N_3772,In_3232,In_336);
nor U3773 (N_3773,In_2931,In_3054);
nor U3774 (N_3774,In_122,In_3735);
nor U3775 (N_3775,In_664,In_544);
and U3776 (N_3776,In_3256,In_377);
nor U3777 (N_3777,In_9,In_3293);
or U3778 (N_3778,In_2473,In_3990);
nand U3779 (N_3779,In_2172,In_4542);
nand U3780 (N_3780,In_933,In_638);
or U3781 (N_3781,In_3902,In_819);
xor U3782 (N_3782,In_269,In_1980);
and U3783 (N_3783,In_379,In_70);
and U3784 (N_3784,In_2283,In_816);
nor U3785 (N_3785,In_3789,In_314);
nand U3786 (N_3786,In_2996,In_1593);
and U3787 (N_3787,In_1922,In_163);
and U3788 (N_3788,In_4302,In_1920);
nor U3789 (N_3789,In_1802,In_1035);
nor U3790 (N_3790,In_4843,In_3426);
xnor U3791 (N_3791,In_4567,In_965);
nor U3792 (N_3792,In_3333,In_2147);
and U3793 (N_3793,In_3994,In_4225);
and U3794 (N_3794,In_3304,In_4430);
and U3795 (N_3795,In_4113,In_4476);
or U3796 (N_3796,In_2968,In_2639);
and U3797 (N_3797,In_4363,In_742);
nor U3798 (N_3798,In_829,In_1723);
nand U3799 (N_3799,In_825,In_4455);
nor U3800 (N_3800,In_659,In_893);
and U3801 (N_3801,In_3523,In_3362);
nand U3802 (N_3802,In_610,In_1430);
xnor U3803 (N_3803,In_2415,In_4808);
and U3804 (N_3804,In_1784,In_3775);
and U3805 (N_3805,In_2747,In_2272);
or U3806 (N_3806,In_563,In_4709);
nand U3807 (N_3807,In_3548,In_1839);
or U3808 (N_3808,In_3517,In_1628);
or U3809 (N_3809,In_3530,In_1962);
xnor U3810 (N_3810,In_4504,In_379);
and U3811 (N_3811,In_2076,In_2230);
nor U3812 (N_3812,In_3174,In_3074);
or U3813 (N_3813,In_3705,In_4886);
or U3814 (N_3814,In_910,In_1776);
nor U3815 (N_3815,In_4931,In_2331);
nor U3816 (N_3816,In_2058,In_3199);
nor U3817 (N_3817,In_2015,In_3263);
and U3818 (N_3818,In_4321,In_3575);
xor U3819 (N_3819,In_366,In_2576);
nand U3820 (N_3820,In_2698,In_103);
nor U3821 (N_3821,In_4491,In_2806);
nand U3822 (N_3822,In_889,In_990);
nor U3823 (N_3823,In_2088,In_515);
and U3824 (N_3824,In_3417,In_1572);
nand U3825 (N_3825,In_3251,In_3164);
nor U3826 (N_3826,In_2305,In_3460);
and U3827 (N_3827,In_4003,In_4278);
and U3828 (N_3828,In_1921,In_4797);
xnor U3829 (N_3829,In_1540,In_1614);
or U3830 (N_3830,In_2604,In_4381);
or U3831 (N_3831,In_1547,In_2869);
xor U3832 (N_3832,In_1285,In_2335);
and U3833 (N_3833,In_4195,In_4353);
nor U3834 (N_3834,In_3679,In_1754);
nand U3835 (N_3835,In_960,In_742);
or U3836 (N_3836,In_4908,In_1042);
nor U3837 (N_3837,In_4030,In_2952);
xor U3838 (N_3838,In_4896,In_1847);
xor U3839 (N_3839,In_3258,In_2026);
or U3840 (N_3840,In_1206,In_4602);
xnor U3841 (N_3841,In_524,In_891);
xnor U3842 (N_3842,In_4916,In_1057);
or U3843 (N_3843,In_382,In_995);
nand U3844 (N_3844,In_730,In_4581);
nand U3845 (N_3845,In_4630,In_1252);
nor U3846 (N_3846,In_3217,In_979);
nand U3847 (N_3847,In_767,In_3942);
or U3848 (N_3848,In_1977,In_2240);
nand U3849 (N_3849,In_739,In_3923);
or U3850 (N_3850,In_1622,In_4930);
and U3851 (N_3851,In_1340,In_295);
nor U3852 (N_3852,In_1085,In_1177);
and U3853 (N_3853,In_3426,In_2762);
xnor U3854 (N_3854,In_1553,In_2386);
nor U3855 (N_3855,In_3873,In_4474);
and U3856 (N_3856,In_4609,In_4014);
xor U3857 (N_3857,In_2388,In_4924);
and U3858 (N_3858,In_634,In_2215);
nor U3859 (N_3859,In_4465,In_3952);
or U3860 (N_3860,In_2916,In_2037);
nand U3861 (N_3861,In_207,In_388);
nor U3862 (N_3862,In_2695,In_3209);
or U3863 (N_3863,In_119,In_635);
nand U3864 (N_3864,In_1405,In_2239);
xnor U3865 (N_3865,In_2441,In_298);
or U3866 (N_3866,In_3844,In_1652);
nor U3867 (N_3867,In_3485,In_2460);
xor U3868 (N_3868,In_677,In_3826);
and U3869 (N_3869,In_585,In_2827);
or U3870 (N_3870,In_1846,In_1249);
xor U3871 (N_3871,In_4613,In_3085);
or U3872 (N_3872,In_3357,In_3586);
and U3873 (N_3873,In_3493,In_2153);
xor U3874 (N_3874,In_829,In_2370);
nor U3875 (N_3875,In_4255,In_3647);
or U3876 (N_3876,In_3525,In_3042);
xor U3877 (N_3877,In_855,In_103);
xnor U3878 (N_3878,In_1814,In_3655);
or U3879 (N_3879,In_3493,In_2017);
and U3880 (N_3880,In_4074,In_4497);
or U3881 (N_3881,In_624,In_4579);
nor U3882 (N_3882,In_2867,In_1984);
or U3883 (N_3883,In_1076,In_1136);
or U3884 (N_3884,In_1891,In_2872);
nor U3885 (N_3885,In_4394,In_3359);
or U3886 (N_3886,In_4093,In_2965);
xor U3887 (N_3887,In_3892,In_2549);
xor U3888 (N_3888,In_4399,In_4089);
nor U3889 (N_3889,In_3271,In_1754);
nand U3890 (N_3890,In_3662,In_4088);
xor U3891 (N_3891,In_2406,In_1956);
xnor U3892 (N_3892,In_4707,In_456);
or U3893 (N_3893,In_1167,In_4131);
and U3894 (N_3894,In_538,In_204);
nor U3895 (N_3895,In_660,In_129);
xor U3896 (N_3896,In_3350,In_4188);
nor U3897 (N_3897,In_1330,In_47);
nor U3898 (N_3898,In_1212,In_4177);
nand U3899 (N_3899,In_4635,In_2327);
or U3900 (N_3900,In_3275,In_596);
and U3901 (N_3901,In_4694,In_4564);
xnor U3902 (N_3902,In_563,In_2486);
nand U3903 (N_3903,In_907,In_2710);
nand U3904 (N_3904,In_2493,In_1869);
nor U3905 (N_3905,In_1346,In_1688);
nand U3906 (N_3906,In_1655,In_1131);
and U3907 (N_3907,In_1580,In_1329);
nor U3908 (N_3908,In_4246,In_793);
or U3909 (N_3909,In_2424,In_500);
or U3910 (N_3910,In_1811,In_2740);
nand U3911 (N_3911,In_3585,In_4470);
xnor U3912 (N_3912,In_1924,In_1254);
nor U3913 (N_3913,In_1333,In_2375);
nand U3914 (N_3914,In_1543,In_3221);
xnor U3915 (N_3915,In_244,In_116);
nor U3916 (N_3916,In_3765,In_532);
nand U3917 (N_3917,In_321,In_3535);
xnor U3918 (N_3918,In_1360,In_4236);
and U3919 (N_3919,In_2682,In_2988);
or U3920 (N_3920,In_3256,In_2631);
nor U3921 (N_3921,In_3398,In_2037);
nor U3922 (N_3922,In_1875,In_995);
or U3923 (N_3923,In_1573,In_1450);
and U3924 (N_3924,In_392,In_2497);
or U3925 (N_3925,In_4231,In_3129);
and U3926 (N_3926,In_2015,In_2465);
or U3927 (N_3927,In_4991,In_2138);
and U3928 (N_3928,In_275,In_3228);
and U3929 (N_3929,In_4940,In_1947);
nor U3930 (N_3930,In_2285,In_3075);
and U3931 (N_3931,In_2606,In_982);
and U3932 (N_3932,In_2707,In_1417);
and U3933 (N_3933,In_1857,In_3774);
and U3934 (N_3934,In_2885,In_4599);
or U3935 (N_3935,In_4940,In_1147);
and U3936 (N_3936,In_3488,In_4853);
xnor U3937 (N_3937,In_2814,In_2416);
and U3938 (N_3938,In_3182,In_1108);
or U3939 (N_3939,In_457,In_2522);
or U3940 (N_3940,In_4898,In_2505);
xnor U3941 (N_3941,In_1423,In_1268);
or U3942 (N_3942,In_3291,In_2042);
nand U3943 (N_3943,In_4286,In_735);
nand U3944 (N_3944,In_4427,In_993);
xnor U3945 (N_3945,In_1267,In_2880);
and U3946 (N_3946,In_3141,In_261);
or U3947 (N_3947,In_516,In_686);
xor U3948 (N_3948,In_1091,In_1605);
nand U3949 (N_3949,In_2522,In_3593);
nand U3950 (N_3950,In_3925,In_2908);
or U3951 (N_3951,In_3379,In_4329);
or U3952 (N_3952,In_3801,In_3413);
xor U3953 (N_3953,In_4504,In_3782);
xnor U3954 (N_3954,In_768,In_1826);
xor U3955 (N_3955,In_722,In_4122);
xor U3956 (N_3956,In_2260,In_217);
nor U3957 (N_3957,In_1742,In_1552);
xor U3958 (N_3958,In_4466,In_3115);
and U3959 (N_3959,In_2844,In_2929);
or U3960 (N_3960,In_4520,In_3029);
or U3961 (N_3961,In_462,In_469);
and U3962 (N_3962,In_706,In_4677);
or U3963 (N_3963,In_4918,In_529);
nand U3964 (N_3964,In_798,In_3720);
nor U3965 (N_3965,In_3475,In_3543);
xnor U3966 (N_3966,In_3690,In_4992);
nor U3967 (N_3967,In_2393,In_3206);
nand U3968 (N_3968,In_59,In_1017);
xor U3969 (N_3969,In_2304,In_3373);
nand U3970 (N_3970,In_84,In_837);
xor U3971 (N_3971,In_4564,In_1829);
nand U3972 (N_3972,In_2225,In_4165);
and U3973 (N_3973,In_4313,In_1057);
and U3974 (N_3974,In_253,In_1580);
nor U3975 (N_3975,In_805,In_4975);
or U3976 (N_3976,In_3770,In_2424);
or U3977 (N_3977,In_4770,In_4335);
and U3978 (N_3978,In_1633,In_2188);
and U3979 (N_3979,In_369,In_1541);
nor U3980 (N_3980,In_2590,In_3000);
and U3981 (N_3981,In_1772,In_1002);
xnor U3982 (N_3982,In_2821,In_2581);
nor U3983 (N_3983,In_4893,In_1295);
xor U3984 (N_3984,In_2899,In_800);
or U3985 (N_3985,In_4713,In_3597);
xnor U3986 (N_3986,In_4925,In_1697);
and U3987 (N_3987,In_3104,In_1939);
xnor U3988 (N_3988,In_456,In_3584);
or U3989 (N_3989,In_674,In_1094);
or U3990 (N_3990,In_4465,In_506);
xnor U3991 (N_3991,In_3540,In_3918);
nor U3992 (N_3992,In_1173,In_4157);
nor U3993 (N_3993,In_3647,In_3467);
or U3994 (N_3994,In_2004,In_2701);
and U3995 (N_3995,In_4916,In_1309);
nand U3996 (N_3996,In_647,In_4920);
nor U3997 (N_3997,In_3370,In_225);
and U3998 (N_3998,In_4470,In_4717);
and U3999 (N_3999,In_3931,In_156);
and U4000 (N_4000,In_4607,In_2821);
or U4001 (N_4001,In_980,In_4834);
xor U4002 (N_4002,In_3380,In_3533);
or U4003 (N_4003,In_3394,In_2225);
xor U4004 (N_4004,In_3241,In_2009);
nor U4005 (N_4005,In_4498,In_3967);
xor U4006 (N_4006,In_1377,In_2370);
and U4007 (N_4007,In_575,In_2487);
nand U4008 (N_4008,In_2321,In_4968);
or U4009 (N_4009,In_1813,In_1761);
nand U4010 (N_4010,In_1871,In_4807);
xnor U4011 (N_4011,In_3807,In_2646);
and U4012 (N_4012,In_1627,In_4950);
and U4013 (N_4013,In_2550,In_3493);
nor U4014 (N_4014,In_4064,In_2438);
or U4015 (N_4015,In_3949,In_2943);
and U4016 (N_4016,In_940,In_1612);
or U4017 (N_4017,In_4558,In_2127);
or U4018 (N_4018,In_3072,In_2330);
nor U4019 (N_4019,In_3373,In_3903);
xor U4020 (N_4020,In_627,In_1335);
nor U4021 (N_4021,In_2969,In_2562);
or U4022 (N_4022,In_3680,In_4358);
and U4023 (N_4023,In_4921,In_4936);
xnor U4024 (N_4024,In_3096,In_1101);
and U4025 (N_4025,In_1453,In_4514);
nor U4026 (N_4026,In_4807,In_1886);
and U4027 (N_4027,In_1762,In_2092);
or U4028 (N_4028,In_2964,In_3636);
nor U4029 (N_4029,In_2477,In_2173);
nand U4030 (N_4030,In_4110,In_3202);
and U4031 (N_4031,In_3496,In_3695);
nand U4032 (N_4032,In_3767,In_4568);
nor U4033 (N_4033,In_3066,In_2155);
xor U4034 (N_4034,In_1490,In_3934);
nor U4035 (N_4035,In_375,In_3979);
or U4036 (N_4036,In_607,In_1002);
nand U4037 (N_4037,In_4030,In_3054);
nand U4038 (N_4038,In_1119,In_4269);
nor U4039 (N_4039,In_4400,In_4780);
nand U4040 (N_4040,In_2002,In_2377);
nor U4041 (N_4041,In_4535,In_1584);
nand U4042 (N_4042,In_4510,In_3741);
nor U4043 (N_4043,In_453,In_1350);
and U4044 (N_4044,In_488,In_1960);
xnor U4045 (N_4045,In_1761,In_3654);
nor U4046 (N_4046,In_145,In_4154);
xnor U4047 (N_4047,In_4400,In_110);
and U4048 (N_4048,In_4456,In_1448);
or U4049 (N_4049,In_751,In_189);
nand U4050 (N_4050,In_1979,In_506);
nor U4051 (N_4051,In_4802,In_2162);
nand U4052 (N_4052,In_4263,In_944);
xor U4053 (N_4053,In_832,In_4763);
nand U4054 (N_4054,In_1648,In_3040);
and U4055 (N_4055,In_540,In_2284);
and U4056 (N_4056,In_501,In_411);
xnor U4057 (N_4057,In_3794,In_4866);
or U4058 (N_4058,In_1598,In_1722);
xnor U4059 (N_4059,In_1296,In_2935);
xor U4060 (N_4060,In_3999,In_2558);
and U4061 (N_4061,In_844,In_4909);
xnor U4062 (N_4062,In_2771,In_4617);
and U4063 (N_4063,In_2712,In_417);
and U4064 (N_4064,In_1682,In_4922);
nor U4065 (N_4065,In_4376,In_1747);
or U4066 (N_4066,In_106,In_3651);
and U4067 (N_4067,In_1080,In_3309);
nand U4068 (N_4068,In_1705,In_1563);
and U4069 (N_4069,In_2819,In_3611);
xor U4070 (N_4070,In_1210,In_2091);
nor U4071 (N_4071,In_1101,In_1613);
xnor U4072 (N_4072,In_2971,In_586);
or U4073 (N_4073,In_3137,In_983);
nand U4074 (N_4074,In_4410,In_2214);
and U4075 (N_4075,In_1955,In_4348);
nand U4076 (N_4076,In_4302,In_156);
xnor U4077 (N_4077,In_2623,In_4550);
nor U4078 (N_4078,In_2733,In_1239);
nor U4079 (N_4079,In_2851,In_4319);
or U4080 (N_4080,In_83,In_4649);
xor U4081 (N_4081,In_2769,In_2604);
nand U4082 (N_4082,In_2401,In_2244);
nor U4083 (N_4083,In_4505,In_2508);
nand U4084 (N_4084,In_4176,In_2049);
nand U4085 (N_4085,In_1959,In_4594);
and U4086 (N_4086,In_3924,In_392);
and U4087 (N_4087,In_4913,In_4358);
xnor U4088 (N_4088,In_4419,In_643);
and U4089 (N_4089,In_3761,In_2345);
nand U4090 (N_4090,In_2340,In_2893);
xor U4091 (N_4091,In_193,In_1936);
xor U4092 (N_4092,In_2427,In_3259);
xor U4093 (N_4093,In_527,In_4966);
and U4094 (N_4094,In_2588,In_4857);
and U4095 (N_4095,In_1374,In_572);
and U4096 (N_4096,In_1859,In_2459);
or U4097 (N_4097,In_101,In_3187);
xnor U4098 (N_4098,In_1882,In_779);
or U4099 (N_4099,In_2363,In_3355);
and U4100 (N_4100,In_4012,In_1217);
xnor U4101 (N_4101,In_3667,In_1402);
or U4102 (N_4102,In_3625,In_543);
nor U4103 (N_4103,In_3605,In_3946);
nand U4104 (N_4104,In_2135,In_170);
or U4105 (N_4105,In_1192,In_1146);
nand U4106 (N_4106,In_675,In_493);
xnor U4107 (N_4107,In_4583,In_4680);
nand U4108 (N_4108,In_2891,In_2765);
nand U4109 (N_4109,In_1236,In_1723);
or U4110 (N_4110,In_4478,In_1581);
and U4111 (N_4111,In_3351,In_2598);
or U4112 (N_4112,In_746,In_1164);
and U4113 (N_4113,In_2598,In_2550);
and U4114 (N_4114,In_598,In_3869);
nor U4115 (N_4115,In_3980,In_1204);
nor U4116 (N_4116,In_2962,In_1051);
nor U4117 (N_4117,In_2783,In_4782);
xor U4118 (N_4118,In_1465,In_1983);
nor U4119 (N_4119,In_2088,In_3055);
and U4120 (N_4120,In_164,In_1034);
xor U4121 (N_4121,In_2917,In_3228);
nand U4122 (N_4122,In_4872,In_4985);
xor U4123 (N_4123,In_4588,In_3328);
xor U4124 (N_4124,In_2580,In_4469);
nor U4125 (N_4125,In_3314,In_1224);
xor U4126 (N_4126,In_1562,In_1527);
nand U4127 (N_4127,In_3988,In_2433);
xor U4128 (N_4128,In_3497,In_1034);
and U4129 (N_4129,In_3164,In_2503);
nor U4130 (N_4130,In_1366,In_24);
and U4131 (N_4131,In_3894,In_695);
or U4132 (N_4132,In_4944,In_4624);
nand U4133 (N_4133,In_970,In_34);
nor U4134 (N_4134,In_3023,In_25);
nand U4135 (N_4135,In_2336,In_2819);
nor U4136 (N_4136,In_789,In_9);
xor U4137 (N_4137,In_1556,In_486);
or U4138 (N_4138,In_1197,In_3185);
or U4139 (N_4139,In_3196,In_2650);
and U4140 (N_4140,In_217,In_4306);
nand U4141 (N_4141,In_1431,In_1862);
nand U4142 (N_4142,In_607,In_4743);
or U4143 (N_4143,In_3178,In_1821);
nor U4144 (N_4144,In_3284,In_3604);
nand U4145 (N_4145,In_211,In_2841);
or U4146 (N_4146,In_1366,In_1534);
or U4147 (N_4147,In_280,In_3535);
nand U4148 (N_4148,In_2321,In_1281);
or U4149 (N_4149,In_1568,In_2318);
nor U4150 (N_4150,In_4963,In_1196);
or U4151 (N_4151,In_3469,In_3903);
and U4152 (N_4152,In_55,In_373);
and U4153 (N_4153,In_1122,In_4546);
nor U4154 (N_4154,In_4568,In_2729);
nand U4155 (N_4155,In_1898,In_4109);
nand U4156 (N_4156,In_2823,In_1432);
and U4157 (N_4157,In_3550,In_2902);
nand U4158 (N_4158,In_3533,In_795);
and U4159 (N_4159,In_3935,In_885);
xnor U4160 (N_4160,In_4753,In_183);
nand U4161 (N_4161,In_2406,In_495);
and U4162 (N_4162,In_934,In_352);
and U4163 (N_4163,In_502,In_4183);
nor U4164 (N_4164,In_3087,In_3199);
nor U4165 (N_4165,In_4790,In_1041);
xnor U4166 (N_4166,In_1286,In_2664);
nand U4167 (N_4167,In_4892,In_883);
nor U4168 (N_4168,In_486,In_1258);
and U4169 (N_4169,In_3250,In_1958);
and U4170 (N_4170,In_2560,In_3035);
and U4171 (N_4171,In_4213,In_217);
or U4172 (N_4172,In_1952,In_4864);
xor U4173 (N_4173,In_3358,In_2121);
nand U4174 (N_4174,In_1635,In_2362);
nor U4175 (N_4175,In_3576,In_2210);
nor U4176 (N_4176,In_4362,In_2316);
xor U4177 (N_4177,In_1044,In_4670);
or U4178 (N_4178,In_1130,In_2166);
or U4179 (N_4179,In_2998,In_3787);
nor U4180 (N_4180,In_4817,In_948);
nor U4181 (N_4181,In_2509,In_658);
xnor U4182 (N_4182,In_2173,In_3720);
nor U4183 (N_4183,In_2659,In_2427);
or U4184 (N_4184,In_4336,In_3436);
xor U4185 (N_4185,In_505,In_940);
nand U4186 (N_4186,In_3083,In_361);
nand U4187 (N_4187,In_3673,In_1774);
nand U4188 (N_4188,In_707,In_581);
or U4189 (N_4189,In_2375,In_4440);
and U4190 (N_4190,In_2200,In_3021);
nand U4191 (N_4191,In_825,In_3574);
and U4192 (N_4192,In_1362,In_1850);
nand U4193 (N_4193,In_47,In_3306);
and U4194 (N_4194,In_2846,In_766);
nor U4195 (N_4195,In_708,In_436);
nor U4196 (N_4196,In_3378,In_800);
and U4197 (N_4197,In_4966,In_1296);
xor U4198 (N_4198,In_2925,In_4539);
nand U4199 (N_4199,In_3455,In_2777);
or U4200 (N_4200,In_169,In_3672);
nor U4201 (N_4201,In_3525,In_2216);
xor U4202 (N_4202,In_2600,In_1222);
nand U4203 (N_4203,In_632,In_4131);
xor U4204 (N_4204,In_765,In_251);
nor U4205 (N_4205,In_972,In_2204);
nand U4206 (N_4206,In_1115,In_1473);
nand U4207 (N_4207,In_2488,In_484);
and U4208 (N_4208,In_2035,In_2817);
nor U4209 (N_4209,In_4308,In_377);
xor U4210 (N_4210,In_2880,In_4249);
and U4211 (N_4211,In_2350,In_4418);
or U4212 (N_4212,In_4933,In_965);
or U4213 (N_4213,In_3650,In_3593);
or U4214 (N_4214,In_3875,In_563);
nand U4215 (N_4215,In_2372,In_2556);
xnor U4216 (N_4216,In_2369,In_1519);
or U4217 (N_4217,In_1770,In_1641);
nor U4218 (N_4218,In_431,In_4965);
or U4219 (N_4219,In_2226,In_1390);
nor U4220 (N_4220,In_181,In_157);
and U4221 (N_4221,In_3311,In_4887);
nand U4222 (N_4222,In_1813,In_2435);
or U4223 (N_4223,In_2984,In_3132);
nand U4224 (N_4224,In_815,In_4499);
or U4225 (N_4225,In_3817,In_616);
or U4226 (N_4226,In_3675,In_4497);
nor U4227 (N_4227,In_2945,In_4142);
nand U4228 (N_4228,In_1617,In_2565);
nand U4229 (N_4229,In_835,In_3506);
nor U4230 (N_4230,In_2227,In_2765);
and U4231 (N_4231,In_879,In_3049);
xor U4232 (N_4232,In_633,In_4277);
nor U4233 (N_4233,In_4909,In_1083);
or U4234 (N_4234,In_1345,In_1917);
or U4235 (N_4235,In_568,In_3440);
and U4236 (N_4236,In_1428,In_681);
or U4237 (N_4237,In_2975,In_3040);
nor U4238 (N_4238,In_986,In_1479);
nor U4239 (N_4239,In_3249,In_3046);
nor U4240 (N_4240,In_2077,In_2318);
xnor U4241 (N_4241,In_3891,In_2935);
nor U4242 (N_4242,In_2772,In_982);
nand U4243 (N_4243,In_1560,In_3652);
and U4244 (N_4244,In_926,In_177);
nand U4245 (N_4245,In_4491,In_476);
nor U4246 (N_4246,In_743,In_3431);
or U4247 (N_4247,In_4555,In_4152);
nor U4248 (N_4248,In_3328,In_3580);
nand U4249 (N_4249,In_1828,In_1097);
xnor U4250 (N_4250,In_4037,In_1440);
nor U4251 (N_4251,In_4442,In_4051);
xnor U4252 (N_4252,In_4305,In_1168);
nor U4253 (N_4253,In_4464,In_4685);
xnor U4254 (N_4254,In_4798,In_1015);
xnor U4255 (N_4255,In_2998,In_4703);
and U4256 (N_4256,In_3568,In_2041);
nand U4257 (N_4257,In_1667,In_4144);
or U4258 (N_4258,In_4401,In_3899);
nand U4259 (N_4259,In_594,In_2881);
nand U4260 (N_4260,In_2430,In_3524);
nand U4261 (N_4261,In_965,In_3411);
and U4262 (N_4262,In_3811,In_1603);
or U4263 (N_4263,In_3081,In_2519);
and U4264 (N_4264,In_4684,In_2204);
and U4265 (N_4265,In_3598,In_1242);
and U4266 (N_4266,In_4329,In_2030);
xnor U4267 (N_4267,In_898,In_328);
or U4268 (N_4268,In_1139,In_3723);
or U4269 (N_4269,In_1700,In_2517);
or U4270 (N_4270,In_1740,In_4906);
nor U4271 (N_4271,In_1071,In_3101);
and U4272 (N_4272,In_1600,In_229);
or U4273 (N_4273,In_3188,In_3842);
nand U4274 (N_4274,In_2867,In_1402);
nand U4275 (N_4275,In_3904,In_4188);
nand U4276 (N_4276,In_2457,In_2619);
xnor U4277 (N_4277,In_1831,In_1322);
and U4278 (N_4278,In_4509,In_2025);
nor U4279 (N_4279,In_3225,In_3195);
nor U4280 (N_4280,In_3674,In_1817);
nor U4281 (N_4281,In_4909,In_3711);
xor U4282 (N_4282,In_1185,In_4460);
and U4283 (N_4283,In_1215,In_3148);
and U4284 (N_4284,In_2056,In_3136);
or U4285 (N_4285,In_1720,In_2134);
or U4286 (N_4286,In_1066,In_387);
nor U4287 (N_4287,In_4439,In_2820);
and U4288 (N_4288,In_2747,In_4926);
or U4289 (N_4289,In_3708,In_856);
nand U4290 (N_4290,In_1683,In_1383);
nor U4291 (N_4291,In_4121,In_431);
xor U4292 (N_4292,In_4316,In_4363);
and U4293 (N_4293,In_4723,In_3567);
or U4294 (N_4294,In_3130,In_3574);
xor U4295 (N_4295,In_3868,In_1290);
and U4296 (N_4296,In_171,In_216);
or U4297 (N_4297,In_2834,In_7);
or U4298 (N_4298,In_2251,In_4739);
or U4299 (N_4299,In_2956,In_1778);
nand U4300 (N_4300,In_2822,In_1088);
nor U4301 (N_4301,In_999,In_362);
or U4302 (N_4302,In_4260,In_1781);
nand U4303 (N_4303,In_3825,In_2548);
or U4304 (N_4304,In_3647,In_2396);
and U4305 (N_4305,In_1059,In_3279);
and U4306 (N_4306,In_329,In_82);
nor U4307 (N_4307,In_4543,In_2676);
or U4308 (N_4308,In_271,In_1024);
nand U4309 (N_4309,In_2541,In_308);
xnor U4310 (N_4310,In_1096,In_1593);
or U4311 (N_4311,In_3477,In_2717);
nor U4312 (N_4312,In_1790,In_3255);
and U4313 (N_4313,In_230,In_2496);
and U4314 (N_4314,In_4372,In_1190);
and U4315 (N_4315,In_3767,In_163);
xor U4316 (N_4316,In_2311,In_666);
nand U4317 (N_4317,In_3838,In_2455);
nor U4318 (N_4318,In_3694,In_3004);
nor U4319 (N_4319,In_2595,In_528);
and U4320 (N_4320,In_360,In_1490);
nor U4321 (N_4321,In_4121,In_4249);
and U4322 (N_4322,In_3380,In_4439);
nand U4323 (N_4323,In_1253,In_547);
xor U4324 (N_4324,In_4491,In_3292);
nand U4325 (N_4325,In_1297,In_4744);
or U4326 (N_4326,In_2540,In_4752);
nor U4327 (N_4327,In_1762,In_3380);
or U4328 (N_4328,In_260,In_3350);
and U4329 (N_4329,In_726,In_4095);
nand U4330 (N_4330,In_2570,In_1245);
nor U4331 (N_4331,In_3518,In_1072);
and U4332 (N_4332,In_1021,In_2860);
nor U4333 (N_4333,In_1332,In_4545);
nand U4334 (N_4334,In_1745,In_3765);
nor U4335 (N_4335,In_2311,In_4328);
and U4336 (N_4336,In_2437,In_132);
or U4337 (N_4337,In_846,In_2603);
xor U4338 (N_4338,In_4223,In_4210);
or U4339 (N_4339,In_2416,In_259);
nor U4340 (N_4340,In_2471,In_1294);
nand U4341 (N_4341,In_1009,In_1041);
xor U4342 (N_4342,In_3709,In_270);
nor U4343 (N_4343,In_578,In_3507);
or U4344 (N_4344,In_1673,In_3218);
or U4345 (N_4345,In_2733,In_967);
nor U4346 (N_4346,In_2888,In_1757);
nor U4347 (N_4347,In_171,In_1636);
and U4348 (N_4348,In_3935,In_524);
nand U4349 (N_4349,In_2934,In_3294);
nand U4350 (N_4350,In_2067,In_3764);
xnor U4351 (N_4351,In_691,In_462);
nor U4352 (N_4352,In_1207,In_3358);
nand U4353 (N_4353,In_3683,In_4369);
and U4354 (N_4354,In_2925,In_373);
or U4355 (N_4355,In_4126,In_493);
or U4356 (N_4356,In_4120,In_1138);
or U4357 (N_4357,In_1559,In_4870);
nor U4358 (N_4358,In_3184,In_1977);
nor U4359 (N_4359,In_2850,In_2282);
and U4360 (N_4360,In_3608,In_829);
xor U4361 (N_4361,In_1399,In_670);
nor U4362 (N_4362,In_743,In_1011);
and U4363 (N_4363,In_1639,In_3392);
nor U4364 (N_4364,In_663,In_4514);
nor U4365 (N_4365,In_3862,In_1965);
nand U4366 (N_4366,In_2632,In_1627);
nand U4367 (N_4367,In_649,In_2042);
or U4368 (N_4368,In_2324,In_234);
nor U4369 (N_4369,In_1483,In_47);
nor U4370 (N_4370,In_1909,In_1846);
nand U4371 (N_4371,In_1012,In_2636);
nand U4372 (N_4372,In_2390,In_3413);
nand U4373 (N_4373,In_2836,In_3794);
nand U4374 (N_4374,In_2464,In_3430);
xnor U4375 (N_4375,In_4103,In_394);
or U4376 (N_4376,In_4545,In_4220);
nand U4377 (N_4377,In_929,In_998);
or U4378 (N_4378,In_2099,In_452);
and U4379 (N_4379,In_3670,In_3343);
xor U4380 (N_4380,In_4169,In_2619);
and U4381 (N_4381,In_520,In_2073);
or U4382 (N_4382,In_505,In_1081);
nand U4383 (N_4383,In_3629,In_3087);
and U4384 (N_4384,In_108,In_1198);
nand U4385 (N_4385,In_1274,In_1508);
nand U4386 (N_4386,In_4898,In_2390);
or U4387 (N_4387,In_121,In_1260);
xor U4388 (N_4388,In_4096,In_4364);
xnor U4389 (N_4389,In_538,In_1604);
nor U4390 (N_4390,In_1053,In_1192);
xnor U4391 (N_4391,In_205,In_971);
nor U4392 (N_4392,In_4131,In_1907);
or U4393 (N_4393,In_3031,In_4610);
nand U4394 (N_4394,In_3827,In_250);
xor U4395 (N_4395,In_2291,In_2390);
or U4396 (N_4396,In_2027,In_3323);
nand U4397 (N_4397,In_1911,In_3219);
nor U4398 (N_4398,In_2338,In_2535);
and U4399 (N_4399,In_815,In_2096);
xnor U4400 (N_4400,In_3135,In_2002);
and U4401 (N_4401,In_4750,In_1224);
and U4402 (N_4402,In_713,In_1749);
nor U4403 (N_4403,In_2958,In_1535);
xor U4404 (N_4404,In_2055,In_4644);
nand U4405 (N_4405,In_1884,In_4767);
or U4406 (N_4406,In_1440,In_1263);
nor U4407 (N_4407,In_4333,In_480);
nor U4408 (N_4408,In_4546,In_2353);
or U4409 (N_4409,In_2908,In_4228);
or U4410 (N_4410,In_3902,In_4455);
and U4411 (N_4411,In_3758,In_2091);
nand U4412 (N_4412,In_3689,In_3935);
xnor U4413 (N_4413,In_3444,In_3309);
and U4414 (N_4414,In_3853,In_517);
and U4415 (N_4415,In_68,In_3438);
or U4416 (N_4416,In_1309,In_4731);
nand U4417 (N_4417,In_3995,In_3941);
nand U4418 (N_4418,In_4996,In_3930);
nor U4419 (N_4419,In_2875,In_885);
nand U4420 (N_4420,In_1689,In_1169);
nor U4421 (N_4421,In_2201,In_1193);
nor U4422 (N_4422,In_1765,In_4257);
or U4423 (N_4423,In_7,In_3119);
nand U4424 (N_4424,In_149,In_3526);
and U4425 (N_4425,In_1349,In_535);
nand U4426 (N_4426,In_796,In_4988);
and U4427 (N_4427,In_1860,In_2689);
xor U4428 (N_4428,In_4740,In_4204);
or U4429 (N_4429,In_3193,In_131);
nand U4430 (N_4430,In_4617,In_1918);
and U4431 (N_4431,In_2340,In_4844);
and U4432 (N_4432,In_2166,In_3693);
nor U4433 (N_4433,In_795,In_1309);
nand U4434 (N_4434,In_2879,In_1410);
nor U4435 (N_4435,In_348,In_398);
xor U4436 (N_4436,In_2852,In_389);
nor U4437 (N_4437,In_1675,In_794);
or U4438 (N_4438,In_2104,In_1803);
and U4439 (N_4439,In_2638,In_1396);
xnor U4440 (N_4440,In_1975,In_1026);
and U4441 (N_4441,In_2429,In_2738);
or U4442 (N_4442,In_4881,In_4564);
or U4443 (N_4443,In_3947,In_2026);
nand U4444 (N_4444,In_1930,In_2688);
and U4445 (N_4445,In_1001,In_880);
nor U4446 (N_4446,In_3908,In_3215);
and U4447 (N_4447,In_2369,In_761);
or U4448 (N_4448,In_1881,In_2987);
and U4449 (N_4449,In_1324,In_3087);
nand U4450 (N_4450,In_4937,In_2671);
nor U4451 (N_4451,In_1958,In_1824);
nand U4452 (N_4452,In_305,In_2942);
xor U4453 (N_4453,In_3323,In_3294);
and U4454 (N_4454,In_344,In_424);
or U4455 (N_4455,In_1270,In_1915);
nand U4456 (N_4456,In_3606,In_3365);
nand U4457 (N_4457,In_1854,In_1398);
or U4458 (N_4458,In_3827,In_3064);
nand U4459 (N_4459,In_3155,In_3549);
and U4460 (N_4460,In_4350,In_894);
nor U4461 (N_4461,In_1585,In_4609);
and U4462 (N_4462,In_2631,In_1143);
or U4463 (N_4463,In_4941,In_408);
nor U4464 (N_4464,In_119,In_2337);
xor U4465 (N_4465,In_4943,In_1535);
xnor U4466 (N_4466,In_258,In_3846);
or U4467 (N_4467,In_29,In_1338);
nor U4468 (N_4468,In_1898,In_958);
nand U4469 (N_4469,In_3234,In_2190);
or U4470 (N_4470,In_4948,In_3620);
and U4471 (N_4471,In_4837,In_2448);
nor U4472 (N_4472,In_4638,In_3656);
nand U4473 (N_4473,In_3028,In_1676);
and U4474 (N_4474,In_4986,In_2539);
xor U4475 (N_4475,In_2360,In_3784);
nand U4476 (N_4476,In_1863,In_4308);
or U4477 (N_4477,In_2823,In_1763);
or U4478 (N_4478,In_1667,In_1494);
or U4479 (N_4479,In_885,In_4109);
xnor U4480 (N_4480,In_3601,In_1243);
or U4481 (N_4481,In_4587,In_3182);
or U4482 (N_4482,In_4975,In_4458);
nor U4483 (N_4483,In_2481,In_3152);
or U4484 (N_4484,In_1697,In_787);
nand U4485 (N_4485,In_3836,In_1694);
nand U4486 (N_4486,In_806,In_952);
xor U4487 (N_4487,In_678,In_415);
nand U4488 (N_4488,In_3777,In_1399);
and U4489 (N_4489,In_108,In_3585);
nand U4490 (N_4490,In_205,In_698);
xor U4491 (N_4491,In_1098,In_990);
nand U4492 (N_4492,In_1109,In_4738);
nand U4493 (N_4493,In_242,In_389);
xnor U4494 (N_4494,In_3909,In_3694);
xnor U4495 (N_4495,In_4802,In_976);
and U4496 (N_4496,In_4075,In_2634);
or U4497 (N_4497,In_4966,In_2642);
and U4498 (N_4498,In_69,In_2955);
nand U4499 (N_4499,In_4587,In_320);
nand U4500 (N_4500,In_197,In_1020);
nand U4501 (N_4501,In_4379,In_3659);
nand U4502 (N_4502,In_3383,In_3090);
and U4503 (N_4503,In_3704,In_3605);
xor U4504 (N_4504,In_1228,In_3989);
or U4505 (N_4505,In_565,In_1072);
nand U4506 (N_4506,In_1982,In_918);
or U4507 (N_4507,In_1239,In_2857);
or U4508 (N_4508,In_2118,In_272);
or U4509 (N_4509,In_436,In_4512);
nand U4510 (N_4510,In_649,In_2910);
or U4511 (N_4511,In_2671,In_3030);
nor U4512 (N_4512,In_4473,In_1287);
nor U4513 (N_4513,In_3697,In_3339);
nand U4514 (N_4514,In_3013,In_1430);
and U4515 (N_4515,In_3302,In_2484);
nand U4516 (N_4516,In_4912,In_4374);
xor U4517 (N_4517,In_371,In_832);
and U4518 (N_4518,In_652,In_3628);
nand U4519 (N_4519,In_2573,In_466);
and U4520 (N_4520,In_4991,In_3695);
or U4521 (N_4521,In_3254,In_3952);
xnor U4522 (N_4522,In_131,In_1093);
and U4523 (N_4523,In_1211,In_2035);
and U4524 (N_4524,In_3535,In_3568);
nand U4525 (N_4525,In_1876,In_2698);
xnor U4526 (N_4526,In_2967,In_3555);
nor U4527 (N_4527,In_4082,In_4994);
nand U4528 (N_4528,In_3917,In_3343);
and U4529 (N_4529,In_342,In_3119);
or U4530 (N_4530,In_249,In_1923);
xor U4531 (N_4531,In_4338,In_758);
nor U4532 (N_4532,In_4790,In_1188);
or U4533 (N_4533,In_4324,In_2299);
and U4534 (N_4534,In_4176,In_3224);
nand U4535 (N_4535,In_4111,In_2101);
and U4536 (N_4536,In_3076,In_254);
nor U4537 (N_4537,In_4485,In_3224);
xnor U4538 (N_4538,In_2884,In_2568);
nand U4539 (N_4539,In_4929,In_518);
or U4540 (N_4540,In_1729,In_3914);
or U4541 (N_4541,In_4,In_4657);
or U4542 (N_4542,In_4695,In_762);
xor U4543 (N_4543,In_951,In_737);
or U4544 (N_4544,In_3745,In_2783);
and U4545 (N_4545,In_3744,In_4593);
xnor U4546 (N_4546,In_1558,In_711);
xnor U4547 (N_4547,In_4423,In_2888);
and U4548 (N_4548,In_1564,In_367);
nor U4549 (N_4549,In_1137,In_3618);
nor U4550 (N_4550,In_4347,In_326);
or U4551 (N_4551,In_3195,In_170);
nand U4552 (N_4552,In_4583,In_4501);
nand U4553 (N_4553,In_1845,In_2928);
xnor U4554 (N_4554,In_4496,In_2673);
nand U4555 (N_4555,In_3478,In_4261);
nor U4556 (N_4556,In_4150,In_1);
and U4557 (N_4557,In_1432,In_2632);
xnor U4558 (N_4558,In_4945,In_816);
nand U4559 (N_4559,In_2447,In_3811);
nand U4560 (N_4560,In_3916,In_912);
or U4561 (N_4561,In_1392,In_2273);
and U4562 (N_4562,In_4629,In_3197);
or U4563 (N_4563,In_580,In_2659);
nand U4564 (N_4564,In_3116,In_306);
or U4565 (N_4565,In_3858,In_1055);
nand U4566 (N_4566,In_847,In_4675);
nor U4567 (N_4567,In_2357,In_739);
and U4568 (N_4568,In_3567,In_678);
nand U4569 (N_4569,In_168,In_149);
nor U4570 (N_4570,In_1814,In_3699);
or U4571 (N_4571,In_1031,In_3835);
or U4572 (N_4572,In_3359,In_4916);
nand U4573 (N_4573,In_4495,In_3467);
or U4574 (N_4574,In_3596,In_3030);
xor U4575 (N_4575,In_4156,In_2784);
nor U4576 (N_4576,In_3394,In_201);
and U4577 (N_4577,In_235,In_3973);
or U4578 (N_4578,In_2096,In_2328);
nand U4579 (N_4579,In_3752,In_74);
nor U4580 (N_4580,In_4669,In_2911);
or U4581 (N_4581,In_4635,In_1535);
and U4582 (N_4582,In_3838,In_565);
or U4583 (N_4583,In_1976,In_1132);
nand U4584 (N_4584,In_2918,In_4007);
nor U4585 (N_4585,In_1169,In_681);
nand U4586 (N_4586,In_4907,In_3539);
nand U4587 (N_4587,In_2219,In_2536);
nor U4588 (N_4588,In_1430,In_590);
nor U4589 (N_4589,In_3792,In_3421);
nor U4590 (N_4590,In_3261,In_2491);
or U4591 (N_4591,In_3421,In_4093);
nor U4592 (N_4592,In_3106,In_2525);
or U4593 (N_4593,In_133,In_521);
and U4594 (N_4594,In_1259,In_3509);
or U4595 (N_4595,In_2336,In_4136);
or U4596 (N_4596,In_535,In_1314);
and U4597 (N_4597,In_1920,In_3521);
nand U4598 (N_4598,In_2035,In_4001);
or U4599 (N_4599,In_4052,In_4920);
and U4600 (N_4600,In_690,In_3491);
nor U4601 (N_4601,In_4488,In_2863);
and U4602 (N_4602,In_4032,In_1595);
or U4603 (N_4603,In_4664,In_1853);
and U4604 (N_4604,In_4916,In_3585);
nor U4605 (N_4605,In_1579,In_1166);
or U4606 (N_4606,In_2258,In_58);
nor U4607 (N_4607,In_3908,In_807);
nand U4608 (N_4608,In_2724,In_4025);
nor U4609 (N_4609,In_679,In_3212);
nor U4610 (N_4610,In_1286,In_4767);
xor U4611 (N_4611,In_327,In_1796);
and U4612 (N_4612,In_3831,In_3520);
xnor U4613 (N_4613,In_4312,In_2117);
nor U4614 (N_4614,In_3044,In_4176);
and U4615 (N_4615,In_3373,In_1061);
xnor U4616 (N_4616,In_635,In_3605);
nor U4617 (N_4617,In_1603,In_1923);
nand U4618 (N_4618,In_3645,In_3967);
or U4619 (N_4619,In_4308,In_407);
nor U4620 (N_4620,In_1781,In_4354);
nor U4621 (N_4621,In_1646,In_3977);
nor U4622 (N_4622,In_2322,In_3159);
and U4623 (N_4623,In_3553,In_1341);
nand U4624 (N_4624,In_1659,In_2604);
and U4625 (N_4625,In_2062,In_4916);
xor U4626 (N_4626,In_4162,In_763);
nand U4627 (N_4627,In_1231,In_854);
xor U4628 (N_4628,In_3143,In_4104);
or U4629 (N_4629,In_100,In_13);
and U4630 (N_4630,In_3443,In_3745);
xnor U4631 (N_4631,In_1569,In_4192);
nor U4632 (N_4632,In_150,In_3403);
xor U4633 (N_4633,In_4243,In_4746);
xnor U4634 (N_4634,In_4389,In_277);
nor U4635 (N_4635,In_1829,In_3105);
and U4636 (N_4636,In_1174,In_2655);
xor U4637 (N_4637,In_995,In_429);
xor U4638 (N_4638,In_1584,In_2351);
and U4639 (N_4639,In_4702,In_4687);
nor U4640 (N_4640,In_2475,In_233);
nor U4641 (N_4641,In_4427,In_2099);
nor U4642 (N_4642,In_798,In_654);
nand U4643 (N_4643,In_2764,In_1832);
nand U4644 (N_4644,In_1858,In_2563);
or U4645 (N_4645,In_4893,In_4662);
and U4646 (N_4646,In_1449,In_2263);
or U4647 (N_4647,In_2206,In_2408);
xnor U4648 (N_4648,In_3340,In_4342);
or U4649 (N_4649,In_416,In_16);
or U4650 (N_4650,In_3284,In_3930);
nand U4651 (N_4651,In_3246,In_3738);
or U4652 (N_4652,In_694,In_4271);
nor U4653 (N_4653,In_4333,In_364);
or U4654 (N_4654,In_4112,In_2075);
or U4655 (N_4655,In_3726,In_29);
and U4656 (N_4656,In_2705,In_539);
nor U4657 (N_4657,In_4639,In_3745);
nand U4658 (N_4658,In_1101,In_3603);
nor U4659 (N_4659,In_2645,In_1571);
xnor U4660 (N_4660,In_912,In_1955);
or U4661 (N_4661,In_1088,In_3287);
or U4662 (N_4662,In_1411,In_4319);
and U4663 (N_4663,In_1924,In_3665);
xor U4664 (N_4664,In_1707,In_917);
and U4665 (N_4665,In_4696,In_45);
nand U4666 (N_4666,In_4767,In_3276);
nand U4667 (N_4667,In_1752,In_4294);
nor U4668 (N_4668,In_3682,In_220);
nand U4669 (N_4669,In_3364,In_2913);
nor U4670 (N_4670,In_4623,In_2571);
nor U4671 (N_4671,In_3441,In_4643);
nand U4672 (N_4672,In_4209,In_3123);
xor U4673 (N_4673,In_1629,In_4235);
or U4674 (N_4674,In_3103,In_4761);
or U4675 (N_4675,In_2879,In_4044);
nor U4676 (N_4676,In_342,In_4754);
or U4677 (N_4677,In_4662,In_922);
and U4678 (N_4678,In_3357,In_4788);
nand U4679 (N_4679,In_1836,In_2500);
or U4680 (N_4680,In_2826,In_3758);
nor U4681 (N_4681,In_599,In_1701);
or U4682 (N_4682,In_2920,In_3479);
xnor U4683 (N_4683,In_1156,In_1803);
or U4684 (N_4684,In_674,In_1271);
nor U4685 (N_4685,In_3934,In_1155);
and U4686 (N_4686,In_196,In_366);
xnor U4687 (N_4687,In_3790,In_115);
nor U4688 (N_4688,In_2648,In_1439);
nor U4689 (N_4689,In_4523,In_1208);
nand U4690 (N_4690,In_4288,In_1668);
nand U4691 (N_4691,In_66,In_812);
and U4692 (N_4692,In_4239,In_1657);
and U4693 (N_4693,In_2187,In_1980);
xor U4694 (N_4694,In_1839,In_3143);
nor U4695 (N_4695,In_4336,In_3598);
or U4696 (N_4696,In_1066,In_2891);
xnor U4697 (N_4697,In_253,In_409);
and U4698 (N_4698,In_4704,In_2635);
nor U4699 (N_4699,In_1904,In_3274);
nand U4700 (N_4700,In_857,In_4893);
and U4701 (N_4701,In_4580,In_3517);
nand U4702 (N_4702,In_754,In_740);
nand U4703 (N_4703,In_4755,In_3441);
or U4704 (N_4704,In_4532,In_4817);
or U4705 (N_4705,In_1786,In_4254);
nand U4706 (N_4706,In_859,In_2525);
and U4707 (N_4707,In_1111,In_4081);
nor U4708 (N_4708,In_3514,In_2635);
nand U4709 (N_4709,In_3158,In_1705);
nor U4710 (N_4710,In_990,In_524);
nand U4711 (N_4711,In_1924,In_4607);
or U4712 (N_4712,In_19,In_3529);
and U4713 (N_4713,In_3793,In_4792);
and U4714 (N_4714,In_2886,In_4685);
or U4715 (N_4715,In_1302,In_4830);
nor U4716 (N_4716,In_1879,In_654);
nand U4717 (N_4717,In_2677,In_280);
and U4718 (N_4718,In_4,In_3631);
nand U4719 (N_4719,In_4832,In_1695);
or U4720 (N_4720,In_2481,In_4841);
and U4721 (N_4721,In_2573,In_2597);
or U4722 (N_4722,In_3935,In_4079);
or U4723 (N_4723,In_174,In_4967);
or U4724 (N_4724,In_494,In_2732);
and U4725 (N_4725,In_4376,In_1972);
and U4726 (N_4726,In_2971,In_2187);
and U4727 (N_4727,In_2806,In_4817);
nor U4728 (N_4728,In_4323,In_1897);
nand U4729 (N_4729,In_67,In_2400);
nand U4730 (N_4730,In_868,In_3232);
or U4731 (N_4731,In_1461,In_4544);
and U4732 (N_4732,In_1169,In_2783);
nor U4733 (N_4733,In_2193,In_1365);
nor U4734 (N_4734,In_4576,In_2339);
or U4735 (N_4735,In_62,In_170);
nand U4736 (N_4736,In_3809,In_4962);
nor U4737 (N_4737,In_4350,In_3750);
or U4738 (N_4738,In_4158,In_115);
nand U4739 (N_4739,In_2455,In_1953);
or U4740 (N_4740,In_1147,In_923);
nand U4741 (N_4741,In_4802,In_1203);
and U4742 (N_4742,In_1809,In_288);
and U4743 (N_4743,In_3176,In_2943);
or U4744 (N_4744,In_3083,In_543);
or U4745 (N_4745,In_4877,In_201);
and U4746 (N_4746,In_3886,In_89);
or U4747 (N_4747,In_3959,In_3902);
nor U4748 (N_4748,In_117,In_1738);
and U4749 (N_4749,In_2453,In_3234);
or U4750 (N_4750,In_2727,In_231);
or U4751 (N_4751,In_3355,In_270);
xnor U4752 (N_4752,In_2450,In_2201);
xor U4753 (N_4753,In_2813,In_1933);
and U4754 (N_4754,In_3171,In_4719);
xnor U4755 (N_4755,In_816,In_1532);
and U4756 (N_4756,In_1546,In_3558);
or U4757 (N_4757,In_965,In_1433);
nand U4758 (N_4758,In_3823,In_1999);
or U4759 (N_4759,In_1543,In_2417);
or U4760 (N_4760,In_3213,In_3296);
nor U4761 (N_4761,In_2854,In_3034);
nand U4762 (N_4762,In_3912,In_3234);
nor U4763 (N_4763,In_2727,In_511);
xor U4764 (N_4764,In_4089,In_289);
or U4765 (N_4765,In_3438,In_4472);
nor U4766 (N_4766,In_619,In_1757);
nor U4767 (N_4767,In_1147,In_4937);
nor U4768 (N_4768,In_4894,In_2284);
xnor U4769 (N_4769,In_2423,In_4422);
nand U4770 (N_4770,In_4215,In_885);
xor U4771 (N_4771,In_2160,In_1829);
and U4772 (N_4772,In_1416,In_353);
or U4773 (N_4773,In_1917,In_1087);
xnor U4774 (N_4774,In_4493,In_4720);
nor U4775 (N_4775,In_1289,In_1354);
and U4776 (N_4776,In_1640,In_4238);
nor U4777 (N_4777,In_1693,In_4116);
or U4778 (N_4778,In_1467,In_3280);
and U4779 (N_4779,In_3283,In_1752);
and U4780 (N_4780,In_1061,In_2941);
and U4781 (N_4781,In_1655,In_2497);
nand U4782 (N_4782,In_1457,In_1716);
nand U4783 (N_4783,In_4176,In_1012);
nand U4784 (N_4784,In_3618,In_699);
nor U4785 (N_4785,In_3264,In_3852);
xor U4786 (N_4786,In_3252,In_873);
or U4787 (N_4787,In_2059,In_4076);
xor U4788 (N_4788,In_445,In_1351);
xnor U4789 (N_4789,In_3054,In_4080);
nor U4790 (N_4790,In_3530,In_539);
or U4791 (N_4791,In_832,In_3142);
nand U4792 (N_4792,In_4252,In_3891);
nor U4793 (N_4793,In_1209,In_2585);
nor U4794 (N_4794,In_426,In_3456);
nor U4795 (N_4795,In_972,In_1730);
and U4796 (N_4796,In_2774,In_4744);
and U4797 (N_4797,In_2133,In_916);
nor U4798 (N_4798,In_3753,In_568);
and U4799 (N_4799,In_4332,In_4406);
or U4800 (N_4800,In_204,In_408);
xor U4801 (N_4801,In_1705,In_1121);
and U4802 (N_4802,In_2267,In_4494);
and U4803 (N_4803,In_4775,In_424);
xnor U4804 (N_4804,In_130,In_4189);
and U4805 (N_4805,In_834,In_4306);
xor U4806 (N_4806,In_2406,In_4236);
and U4807 (N_4807,In_3643,In_3394);
xnor U4808 (N_4808,In_4174,In_3499);
nor U4809 (N_4809,In_826,In_2134);
and U4810 (N_4810,In_4509,In_1322);
and U4811 (N_4811,In_894,In_4652);
nand U4812 (N_4812,In_2258,In_794);
or U4813 (N_4813,In_102,In_1389);
and U4814 (N_4814,In_3042,In_144);
or U4815 (N_4815,In_4529,In_1287);
nor U4816 (N_4816,In_2266,In_4378);
and U4817 (N_4817,In_61,In_4672);
or U4818 (N_4818,In_564,In_2855);
nand U4819 (N_4819,In_4937,In_3380);
or U4820 (N_4820,In_2217,In_3052);
or U4821 (N_4821,In_1262,In_2308);
nor U4822 (N_4822,In_1358,In_3980);
and U4823 (N_4823,In_4670,In_832);
xor U4824 (N_4824,In_2154,In_2183);
or U4825 (N_4825,In_1759,In_1092);
nand U4826 (N_4826,In_4194,In_4074);
nand U4827 (N_4827,In_3137,In_510);
or U4828 (N_4828,In_2524,In_3746);
nor U4829 (N_4829,In_2955,In_4771);
xnor U4830 (N_4830,In_4319,In_2341);
nand U4831 (N_4831,In_1333,In_2452);
nand U4832 (N_4832,In_60,In_4634);
nor U4833 (N_4833,In_2059,In_3647);
nor U4834 (N_4834,In_2729,In_1553);
nor U4835 (N_4835,In_846,In_4409);
and U4836 (N_4836,In_3674,In_3957);
or U4837 (N_4837,In_68,In_3800);
nor U4838 (N_4838,In_1001,In_3364);
xor U4839 (N_4839,In_3001,In_2351);
and U4840 (N_4840,In_1238,In_4890);
nor U4841 (N_4841,In_263,In_3752);
xnor U4842 (N_4842,In_4004,In_2297);
xnor U4843 (N_4843,In_4281,In_4752);
or U4844 (N_4844,In_3135,In_4453);
nand U4845 (N_4845,In_3945,In_2990);
or U4846 (N_4846,In_2387,In_2019);
and U4847 (N_4847,In_4198,In_2602);
or U4848 (N_4848,In_4042,In_4660);
nand U4849 (N_4849,In_786,In_2328);
nand U4850 (N_4850,In_4259,In_213);
or U4851 (N_4851,In_1633,In_1437);
nor U4852 (N_4852,In_3980,In_2718);
and U4853 (N_4853,In_4622,In_4340);
or U4854 (N_4854,In_4005,In_4393);
nor U4855 (N_4855,In_1319,In_4439);
nor U4856 (N_4856,In_933,In_2874);
nor U4857 (N_4857,In_1861,In_281);
or U4858 (N_4858,In_1128,In_4472);
xnor U4859 (N_4859,In_4449,In_572);
nand U4860 (N_4860,In_2309,In_2098);
nand U4861 (N_4861,In_4190,In_2172);
and U4862 (N_4862,In_4883,In_1921);
or U4863 (N_4863,In_4329,In_2525);
and U4864 (N_4864,In_3668,In_4522);
xor U4865 (N_4865,In_1958,In_4048);
nand U4866 (N_4866,In_3987,In_4058);
or U4867 (N_4867,In_2548,In_3983);
or U4868 (N_4868,In_2384,In_4176);
nor U4869 (N_4869,In_1614,In_691);
xor U4870 (N_4870,In_1046,In_769);
xor U4871 (N_4871,In_2237,In_454);
xor U4872 (N_4872,In_2297,In_1923);
or U4873 (N_4873,In_442,In_3788);
or U4874 (N_4874,In_595,In_2098);
nor U4875 (N_4875,In_1880,In_561);
xor U4876 (N_4876,In_2013,In_3101);
nand U4877 (N_4877,In_1559,In_3713);
nor U4878 (N_4878,In_4673,In_562);
nor U4879 (N_4879,In_2551,In_1739);
nor U4880 (N_4880,In_1659,In_2774);
nor U4881 (N_4881,In_561,In_2057);
or U4882 (N_4882,In_844,In_2678);
or U4883 (N_4883,In_3709,In_3172);
and U4884 (N_4884,In_3076,In_2053);
nand U4885 (N_4885,In_2157,In_1767);
xor U4886 (N_4886,In_1147,In_3348);
nor U4887 (N_4887,In_2701,In_1789);
xnor U4888 (N_4888,In_140,In_327);
and U4889 (N_4889,In_2271,In_552);
and U4890 (N_4890,In_2801,In_2223);
xor U4891 (N_4891,In_2150,In_799);
or U4892 (N_4892,In_4406,In_846);
nand U4893 (N_4893,In_1799,In_2493);
xnor U4894 (N_4894,In_4966,In_4713);
nor U4895 (N_4895,In_2784,In_100);
xor U4896 (N_4896,In_4793,In_1274);
nand U4897 (N_4897,In_3533,In_4877);
nand U4898 (N_4898,In_2792,In_187);
or U4899 (N_4899,In_4199,In_903);
nand U4900 (N_4900,In_311,In_120);
or U4901 (N_4901,In_843,In_1569);
or U4902 (N_4902,In_3437,In_3134);
and U4903 (N_4903,In_1924,In_477);
or U4904 (N_4904,In_2075,In_1864);
xnor U4905 (N_4905,In_2234,In_3010);
or U4906 (N_4906,In_4680,In_3487);
and U4907 (N_4907,In_1566,In_1906);
nor U4908 (N_4908,In_3081,In_4006);
nor U4909 (N_4909,In_258,In_3152);
nand U4910 (N_4910,In_548,In_2920);
nor U4911 (N_4911,In_262,In_3190);
xor U4912 (N_4912,In_855,In_1237);
or U4913 (N_4913,In_396,In_3112);
and U4914 (N_4914,In_3644,In_2660);
and U4915 (N_4915,In_2990,In_3620);
xnor U4916 (N_4916,In_4988,In_192);
or U4917 (N_4917,In_861,In_727);
xnor U4918 (N_4918,In_2999,In_418);
or U4919 (N_4919,In_2673,In_521);
and U4920 (N_4920,In_4715,In_2155);
nand U4921 (N_4921,In_3189,In_4791);
nor U4922 (N_4922,In_360,In_2290);
or U4923 (N_4923,In_2427,In_1117);
nand U4924 (N_4924,In_2925,In_4711);
nor U4925 (N_4925,In_3674,In_4390);
or U4926 (N_4926,In_2814,In_1655);
and U4927 (N_4927,In_237,In_2433);
nand U4928 (N_4928,In_535,In_4425);
nor U4929 (N_4929,In_3963,In_25);
or U4930 (N_4930,In_1419,In_3048);
or U4931 (N_4931,In_2249,In_567);
or U4932 (N_4932,In_67,In_2897);
nor U4933 (N_4933,In_832,In_2985);
nand U4934 (N_4934,In_3402,In_2986);
nand U4935 (N_4935,In_3129,In_3630);
xnor U4936 (N_4936,In_1872,In_4071);
nand U4937 (N_4937,In_29,In_2377);
xor U4938 (N_4938,In_3591,In_121);
nor U4939 (N_4939,In_908,In_4104);
nor U4940 (N_4940,In_165,In_4723);
xor U4941 (N_4941,In_4922,In_2687);
nor U4942 (N_4942,In_4558,In_585);
nor U4943 (N_4943,In_800,In_4978);
or U4944 (N_4944,In_1854,In_4882);
or U4945 (N_4945,In_2641,In_1646);
or U4946 (N_4946,In_773,In_1545);
xnor U4947 (N_4947,In_3811,In_4313);
xor U4948 (N_4948,In_1684,In_3911);
and U4949 (N_4949,In_4804,In_336);
nand U4950 (N_4950,In_3620,In_2912);
nor U4951 (N_4951,In_384,In_1344);
xnor U4952 (N_4952,In_3667,In_4704);
and U4953 (N_4953,In_4062,In_202);
nor U4954 (N_4954,In_904,In_3307);
nand U4955 (N_4955,In_19,In_1865);
xnor U4956 (N_4956,In_965,In_3261);
nand U4957 (N_4957,In_3302,In_1171);
nor U4958 (N_4958,In_3171,In_925);
nand U4959 (N_4959,In_4081,In_4318);
nand U4960 (N_4960,In_4596,In_758);
nand U4961 (N_4961,In_3670,In_981);
nand U4962 (N_4962,In_2716,In_1813);
nor U4963 (N_4963,In_1417,In_3668);
nand U4964 (N_4964,In_4176,In_723);
and U4965 (N_4965,In_1680,In_2057);
and U4966 (N_4966,In_117,In_1386);
nor U4967 (N_4967,In_2537,In_4647);
xnor U4968 (N_4968,In_3308,In_842);
or U4969 (N_4969,In_1600,In_2136);
and U4970 (N_4970,In_50,In_3416);
xnor U4971 (N_4971,In_3733,In_1062);
and U4972 (N_4972,In_4899,In_4700);
nand U4973 (N_4973,In_996,In_3548);
nand U4974 (N_4974,In_3370,In_2890);
or U4975 (N_4975,In_3082,In_1556);
nor U4976 (N_4976,In_4321,In_2047);
and U4977 (N_4977,In_4437,In_2043);
xnor U4978 (N_4978,In_559,In_1695);
or U4979 (N_4979,In_489,In_4397);
and U4980 (N_4980,In_3408,In_197);
xnor U4981 (N_4981,In_2165,In_3922);
and U4982 (N_4982,In_631,In_3394);
nor U4983 (N_4983,In_179,In_350);
xnor U4984 (N_4984,In_3419,In_3370);
xnor U4985 (N_4985,In_3267,In_872);
nand U4986 (N_4986,In_2037,In_3231);
and U4987 (N_4987,In_3916,In_4416);
and U4988 (N_4988,In_390,In_966);
or U4989 (N_4989,In_223,In_4611);
or U4990 (N_4990,In_526,In_1874);
nor U4991 (N_4991,In_235,In_3287);
and U4992 (N_4992,In_3253,In_2527);
nor U4993 (N_4993,In_716,In_527);
and U4994 (N_4994,In_2387,In_474);
and U4995 (N_4995,In_2182,In_1334);
xor U4996 (N_4996,In_1693,In_1224);
and U4997 (N_4997,In_3333,In_1671);
nand U4998 (N_4998,In_269,In_3397);
nor U4999 (N_4999,In_132,In_151);
or U5000 (N_5000,N_2879,N_98);
and U5001 (N_5001,N_4079,N_1598);
and U5002 (N_5002,N_4153,N_2006);
and U5003 (N_5003,N_2873,N_3539);
nor U5004 (N_5004,N_1344,N_4854);
xor U5005 (N_5005,N_4692,N_2143);
nor U5006 (N_5006,N_4935,N_1083);
and U5007 (N_5007,N_4511,N_3380);
nor U5008 (N_5008,N_2785,N_4028);
xor U5009 (N_5009,N_347,N_3593);
and U5010 (N_5010,N_1823,N_3468);
nand U5011 (N_5011,N_3661,N_2965);
nand U5012 (N_5012,N_237,N_4505);
nor U5013 (N_5013,N_3592,N_755);
xnor U5014 (N_5014,N_1479,N_4922);
and U5015 (N_5015,N_4482,N_1700);
and U5016 (N_5016,N_1876,N_4494);
nand U5017 (N_5017,N_498,N_2048);
and U5018 (N_5018,N_3718,N_4977);
xnor U5019 (N_5019,N_1570,N_1683);
nor U5020 (N_5020,N_3395,N_3148);
and U5021 (N_5021,N_1157,N_3596);
or U5022 (N_5022,N_834,N_2061);
nor U5023 (N_5023,N_2763,N_1052);
and U5024 (N_5024,N_2177,N_4197);
nor U5025 (N_5025,N_3102,N_1381);
nand U5026 (N_5026,N_3473,N_4286);
nand U5027 (N_5027,N_1580,N_2255);
and U5028 (N_5028,N_4044,N_1502);
nand U5029 (N_5029,N_1872,N_2779);
or U5030 (N_5030,N_262,N_3039);
or U5031 (N_5031,N_635,N_2246);
xnor U5032 (N_5032,N_1739,N_272);
and U5033 (N_5033,N_1684,N_2810);
nand U5034 (N_5034,N_1702,N_2844);
or U5035 (N_5035,N_550,N_3553);
and U5036 (N_5036,N_249,N_2482);
and U5037 (N_5037,N_4576,N_1875);
or U5038 (N_5038,N_912,N_2588);
or U5039 (N_5039,N_2921,N_3507);
and U5040 (N_5040,N_4885,N_1676);
or U5041 (N_5041,N_306,N_4292);
or U5042 (N_5042,N_4160,N_2804);
nand U5043 (N_5043,N_4604,N_3470);
nor U5044 (N_5044,N_343,N_4451);
nand U5045 (N_5045,N_4696,N_3526);
and U5046 (N_5046,N_3945,N_2562);
and U5047 (N_5047,N_3589,N_1153);
nor U5048 (N_5048,N_4655,N_3022);
nand U5049 (N_5049,N_4860,N_1449);
or U5050 (N_5050,N_2712,N_749);
nand U5051 (N_5051,N_663,N_1483);
nor U5052 (N_5052,N_3780,N_2869);
and U5053 (N_5053,N_3610,N_4296);
or U5054 (N_5054,N_108,N_1377);
nand U5055 (N_5055,N_977,N_1627);
and U5056 (N_5056,N_3578,N_3571);
nor U5057 (N_5057,N_131,N_1250);
or U5058 (N_5058,N_3678,N_3434);
nand U5059 (N_5059,N_1279,N_4512);
xnor U5060 (N_5060,N_4502,N_985);
nor U5061 (N_5061,N_4087,N_3546);
nand U5062 (N_5062,N_1681,N_596);
and U5063 (N_5063,N_1977,N_3160);
or U5064 (N_5064,N_4058,N_4617);
and U5065 (N_5065,N_81,N_3574);
nand U5066 (N_5066,N_4788,N_3189);
and U5067 (N_5067,N_4312,N_565);
xnor U5068 (N_5068,N_1431,N_610);
and U5069 (N_5069,N_3585,N_567);
xor U5070 (N_5070,N_3796,N_3831);
nand U5071 (N_5071,N_3629,N_2248);
and U5072 (N_5072,N_1557,N_3449);
xnor U5073 (N_5073,N_1675,N_4546);
nor U5074 (N_5074,N_1240,N_1630);
nand U5075 (N_5075,N_2990,N_4104);
nand U5076 (N_5076,N_1649,N_2529);
nand U5077 (N_5077,N_3698,N_4179);
nor U5078 (N_5078,N_3535,N_4510);
nand U5079 (N_5079,N_3794,N_1738);
or U5080 (N_5080,N_1399,N_4279);
nand U5081 (N_5081,N_3351,N_4839);
nor U5082 (N_5082,N_119,N_2372);
xor U5083 (N_5083,N_1108,N_3634);
or U5084 (N_5084,N_2633,N_430);
and U5085 (N_5085,N_745,N_2442);
or U5086 (N_5086,N_2789,N_1162);
xnor U5087 (N_5087,N_2877,N_43);
xnor U5088 (N_5088,N_2101,N_701);
nor U5089 (N_5089,N_4049,N_4402);
nor U5090 (N_5090,N_4262,N_691);
xor U5091 (N_5091,N_250,N_3943);
nor U5092 (N_5092,N_1165,N_2882);
and U5093 (N_5093,N_1476,N_1861);
xor U5094 (N_5094,N_2000,N_1520);
or U5095 (N_5095,N_3472,N_1424);
nand U5096 (N_5096,N_3566,N_3904);
xnor U5097 (N_5097,N_1025,N_1439);
nand U5098 (N_5098,N_978,N_4660);
nor U5099 (N_5099,N_4877,N_4543);
nand U5100 (N_5100,N_1597,N_1716);
xor U5101 (N_5101,N_930,N_1981);
and U5102 (N_5102,N_4073,N_3327);
nor U5103 (N_5103,N_3726,N_2262);
nand U5104 (N_5104,N_3662,N_1632);
nand U5105 (N_5105,N_3813,N_355);
and U5106 (N_5106,N_463,N_1940);
nor U5107 (N_5107,N_4361,N_4478);
or U5108 (N_5108,N_3016,N_412);
or U5109 (N_5109,N_943,N_4973);
or U5110 (N_5110,N_458,N_1111);
or U5111 (N_5111,N_3443,N_79);
xor U5112 (N_5112,N_1934,N_3847);
nand U5113 (N_5113,N_3930,N_535);
or U5114 (N_5114,N_3776,N_2135);
and U5115 (N_5115,N_4649,N_3488);
nand U5116 (N_5116,N_2540,N_11);
and U5117 (N_5117,N_4100,N_257);
nand U5118 (N_5118,N_1420,N_4497);
xor U5119 (N_5119,N_3205,N_4957);
nand U5120 (N_5120,N_4389,N_3533);
nor U5121 (N_5121,N_4932,N_2075);
or U5122 (N_5122,N_1709,N_4955);
and U5123 (N_5123,N_86,N_1236);
nor U5124 (N_5124,N_1554,N_988);
or U5125 (N_5125,N_4679,N_3287);
nor U5126 (N_5126,N_4670,N_951);
xor U5127 (N_5127,N_804,N_3693);
or U5128 (N_5128,N_2799,N_3707);
and U5129 (N_5129,N_2522,N_4567);
nand U5130 (N_5130,N_4875,N_3834);
and U5131 (N_5131,N_3751,N_4607);
nand U5132 (N_5132,N_2014,N_3128);
xor U5133 (N_5133,N_1835,N_248);
nor U5134 (N_5134,N_2934,N_4491);
xnor U5135 (N_5135,N_766,N_160);
and U5136 (N_5136,N_780,N_1774);
or U5137 (N_5137,N_1751,N_651);
or U5138 (N_5138,N_3106,N_823);
and U5139 (N_5139,N_1574,N_709);
and U5140 (N_5140,N_4254,N_2485);
xnor U5141 (N_5141,N_4564,N_1072);
or U5142 (N_5142,N_3021,N_2387);
or U5143 (N_5143,N_1271,N_4643);
nor U5144 (N_5144,N_3263,N_494);
nor U5145 (N_5145,N_2251,N_335);
or U5146 (N_5146,N_4676,N_2123);
or U5147 (N_5147,N_2284,N_278);
nor U5148 (N_5148,N_4059,N_35);
and U5149 (N_5149,N_4407,N_1543);
and U5150 (N_5150,N_3802,N_2777);
xnor U5151 (N_5151,N_935,N_609);
nand U5152 (N_5152,N_3795,N_2527);
nor U5153 (N_5153,N_1039,N_3699);
or U5154 (N_5154,N_2150,N_3451);
or U5155 (N_5155,N_4615,N_3142);
nor U5156 (N_5156,N_3940,N_3753);
nand U5157 (N_5157,N_1813,N_4014);
nor U5158 (N_5158,N_3427,N_3992);
or U5159 (N_5159,N_33,N_3994);
nand U5160 (N_5160,N_3147,N_4919);
or U5161 (N_5161,N_3027,N_3757);
nand U5162 (N_5162,N_1053,N_4560);
nor U5163 (N_5163,N_2734,N_2096);
nand U5164 (N_5164,N_2681,N_4193);
xor U5165 (N_5165,N_416,N_4062);
nand U5166 (N_5166,N_1801,N_689);
xor U5167 (N_5167,N_1281,N_717);
nand U5168 (N_5168,N_4295,N_1219);
nor U5169 (N_5169,N_2408,N_4359);
xor U5170 (N_5170,N_538,N_3230);
or U5171 (N_5171,N_3176,N_354);
and U5172 (N_5172,N_2563,N_2698);
nand U5173 (N_5173,N_1752,N_2126);
nor U5174 (N_5174,N_2122,N_3630);
and U5175 (N_5175,N_1247,N_1747);
and U5176 (N_5176,N_3722,N_3956);
or U5177 (N_5177,N_3090,N_744);
or U5178 (N_5178,N_1191,N_2535);
and U5179 (N_5179,N_1892,N_846);
and U5180 (N_5180,N_2596,N_4818);
and U5181 (N_5181,N_1354,N_4826);
xnor U5182 (N_5182,N_1489,N_2600);
nor U5183 (N_5183,N_2250,N_1990);
xor U5184 (N_5184,N_1440,N_3264);
and U5185 (N_5185,N_4256,N_2967);
nand U5186 (N_5186,N_2922,N_4527);
and U5187 (N_5187,N_140,N_3942);
and U5188 (N_5188,N_1,N_59);
and U5189 (N_5189,N_2275,N_3639);
nand U5190 (N_5190,N_4164,N_4988);
and U5191 (N_5191,N_1831,N_2863);
xor U5192 (N_5192,N_1372,N_1558);
nand U5193 (N_5193,N_4594,N_1211);
xnor U5194 (N_5194,N_1565,N_3014);
nor U5195 (N_5195,N_4620,N_4903);
and U5196 (N_5196,N_2895,N_1532);
nand U5197 (N_5197,N_1624,N_4908);
or U5198 (N_5198,N_4481,N_3156);
nor U5199 (N_5199,N_3980,N_2927);
xnor U5200 (N_5200,N_168,N_4410);
xor U5201 (N_5201,N_2003,N_161);
or U5202 (N_5202,N_2860,N_1104);
xnor U5203 (N_5203,N_1722,N_4091);
nor U5204 (N_5204,N_1169,N_388);
nand U5205 (N_5205,N_1051,N_1056);
nand U5206 (N_5206,N_619,N_1559);
nor U5207 (N_5207,N_4470,N_4005);
xor U5208 (N_5208,N_92,N_503);
or U5209 (N_5209,N_1343,N_3950);
and U5210 (N_5210,N_3807,N_2621);
nand U5211 (N_5211,N_3150,N_3354);
and U5212 (N_5212,N_1155,N_3116);
xor U5213 (N_5213,N_1304,N_4325);
and U5214 (N_5214,N_2825,N_1694);
nor U5215 (N_5215,N_4868,N_1481);
or U5216 (N_5216,N_3217,N_3213);
nand U5217 (N_5217,N_3317,N_4559);
xor U5218 (N_5218,N_4269,N_3987);
nor U5219 (N_5219,N_4037,N_1326);
nand U5220 (N_5220,N_1112,N_2243);
and U5221 (N_5221,N_3764,N_2585);
nor U5222 (N_5222,N_3700,N_1814);
nor U5223 (N_5223,N_1190,N_4626);
xor U5224 (N_5224,N_615,N_1297);
or U5225 (N_5225,N_3181,N_305);
xor U5226 (N_5226,N_4392,N_4215);
or U5227 (N_5227,N_1468,N_478);
and U5228 (N_5228,N_1874,N_747);
or U5229 (N_5229,N_3816,N_114);
or U5230 (N_5230,N_4943,N_4414);
and U5231 (N_5231,N_147,N_2911);
and U5232 (N_5232,N_3259,N_841);
nand U5233 (N_5233,N_1750,N_4724);
xnor U5234 (N_5234,N_4320,N_3607);
and U5235 (N_5235,N_2127,N_1827);
or U5236 (N_5236,N_3360,N_4961);
nor U5237 (N_5237,N_3626,N_1631);
or U5238 (N_5238,N_1446,N_267);
nor U5239 (N_5239,N_4427,N_4600);
or U5240 (N_5240,N_4161,N_3513);
xor U5241 (N_5241,N_4827,N_2261);
xor U5242 (N_5242,N_2302,N_2132);
and U5243 (N_5243,N_1786,N_3328);
xor U5244 (N_5244,N_4319,N_4820);
nor U5245 (N_5245,N_3918,N_4157);
nor U5246 (N_5246,N_880,N_815);
or U5247 (N_5247,N_1095,N_725);
and U5248 (N_5248,N_496,N_3570);
nor U5249 (N_5249,N_3517,N_135);
and U5250 (N_5250,N_206,N_2446);
xnor U5251 (N_5251,N_684,N_1059);
or U5252 (N_5252,N_4814,N_1176);
or U5253 (N_5253,N_2136,N_4612);
nand U5254 (N_5254,N_3081,N_4586);
nor U5255 (N_5255,N_792,N_653);
nor U5256 (N_5256,N_3050,N_4631);
and U5257 (N_5257,N_3408,N_932);
nor U5258 (N_5258,N_1859,N_126);
nand U5259 (N_5259,N_3197,N_1715);
and U5260 (N_5260,N_403,N_239);
or U5261 (N_5261,N_3364,N_1229);
and U5262 (N_5262,N_1454,N_1746);
nand U5263 (N_5263,N_1885,N_2245);
nand U5264 (N_5264,N_2183,N_2549);
nor U5265 (N_5265,N_4916,N_1825);
nand U5266 (N_5266,N_2793,N_2340);
and U5267 (N_5267,N_616,N_2313);
and U5268 (N_5268,N_4998,N_2656);
xor U5269 (N_5269,N_199,N_294);
and U5270 (N_5270,N_3872,N_428);
nand U5271 (N_5271,N_4298,N_95);
or U5272 (N_5272,N_353,N_4314);
and U5273 (N_5273,N_2159,N_1719);
or U5274 (N_5274,N_1736,N_60);
nand U5275 (N_5275,N_2818,N_2885);
xor U5276 (N_5276,N_2521,N_2500);
nand U5277 (N_5277,N_898,N_4270);
nor U5278 (N_5278,N_2272,N_1414);
nor U5279 (N_5279,N_222,N_1070);
nand U5280 (N_5280,N_4458,N_3387);
and U5281 (N_5281,N_1006,N_4796);
xnor U5282 (N_5282,N_15,N_3411);
or U5283 (N_5283,N_2182,N_2821);
or U5284 (N_5284,N_4188,N_2117);
and U5285 (N_5285,N_2497,N_2983);
nor U5286 (N_5286,N_1980,N_3322);
or U5287 (N_5287,N_1171,N_2084);
or U5288 (N_5288,N_1878,N_2627);
xor U5289 (N_5289,N_825,N_1090);
nor U5290 (N_5290,N_500,N_752);
xnor U5291 (N_5291,N_1259,N_986);
and U5292 (N_5292,N_3685,N_417);
nand U5293 (N_5293,N_3618,N_205);
xor U5294 (N_5294,N_2568,N_4504);
xnor U5295 (N_5295,N_2209,N_2597);
and U5296 (N_5296,N_3867,N_2756);
and U5297 (N_5297,N_2267,N_4452);
and U5298 (N_5298,N_4486,N_3854);
nor U5299 (N_5299,N_1926,N_133);
nand U5300 (N_5300,N_3686,N_3031);
nor U5301 (N_5301,N_3278,N_4343);
and U5302 (N_5302,N_763,N_3551);
nand U5303 (N_5303,N_3073,N_185);
nand U5304 (N_5304,N_38,N_854);
and U5305 (N_5305,N_4758,N_4630);
and U5306 (N_5306,N_1121,N_3540);
xnor U5307 (N_5307,N_800,N_1436);
xnor U5308 (N_5308,N_1886,N_1034);
xnor U5309 (N_5309,N_4332,N_3399);
xor U5310 (N_5310,N_1351,N_323);
and U5311 (N_5311,N_97,N_3774);
or U5312 (N_5312,N_3727,N_3199);
xnor U5313 (N_5313,N_4236,N_4180);
nor U5314 (N_5314,N_4734,N_631);
nand U5315 (N_5315,N_2839,N_2450);
and U5316 (N_5316,N_2155,N_4151);
or U5317 (N_5317,N_1928,N_1817);
or U5318 (N_5318,N_3061,N_279);
and U5319 (N_5319,N_3193,N_3300);
nand U5320 (N_5320,N_2192,N_2021);
and U5321 (N_5321,N_1525,N_1612);
and U5322 (N_5322,N_1541,N_3382);
xor U5323 (N_5323,N_3746,N_4201);
xor U5324 (N_5324,N_1088,N_2888);
nand U5325 (N_5325,N_564,N_961);
xor U5326 (N_5326,N_220,N_4233);
nand U5327 (N_5327,N_3967,N_1415);
and U5328 (N_5328,N_2494,N_3799);
or U5329 (N_5329,N_3186,N_1332);
and U5330 (N_5330,N_1201,N_4387);
or U5331 (N_5331,N_2374,N_2291);
or U5332 (N_5332,N_579,N_4728);
nor U5333 (N_5333,N_3255,N_4130);
nand U5334 (N_5334,N_1772,N_2750);
xnor U5335 (N_5335,N_2541,N_711);
and U5336 (N_5336,N_4095,N_1042);
nand U5337 (N_5337,N_1316,N_177);
nand U5338 (N_5338,N_4646,N_1067);
and U5339 (N_5339,N_2841,N_4872);
nor U5340 (N_5340,N_3695,N_2931);
nand U5341 (N_5341,N_3497,N_4408);
nand U5342 (N_5342,N_327,N_838);
xnor U5343 (N_5343,N_3243,N_1726);
nor U5344 (N_5344,N_2448,N_1895);
nor U5345 (N_5345,N_64,N_3273);
and U5346 (N_5346,N_724,N_3909);
or U5347 (N_5347,N_3801,N_284);
nand U5348 (N_5348,N_3284,N_967);
or U5349 (N_5349,N_4847,N_2655);
nor U5350 (N_5350,N_3544,N_4134);
and U5351 (N_5351,N_1196,N_4240);
nand U5352 (N_5352,N_4082,N_3232);
or U5353 (N_5353,N_990,N_2773);
nor U5354 (N_5354,N_3966,N_2214);
nor U5355 (N_5355,N_674,N_2795);
or U5356 (N_5356,N_4303,N_1788);
or U5357 (N_5357,N_2912,N_2378);
xor U5358 (N_5358,N_1089,N_2998);
nor U5359 (N_5359,N_4810,N_4550);
or U5360 (N_5360,N_76,N_1593);
nand U5361 (N_5361,N_2315,N_3237);
and U5362 (N_5362,N_3792,N_4918);
xor U5363 (N_5363,N_3149,N_2066);
nand U5364 (N_5364,N_3173,N_137);
xnor U5365 (N_5365,N_2131,N_3682);
xnor U5366 (N_5366,N_3803,N_2964);
nand U5367 (N_5367,N_1704,N_3219);
nor U5368 (N_5368,N_2537,N_605);
or U5369 (N_5369,N_620,N_4386);
xnor U5370 (N_5370,N_4742,N_4686);
or U5371 (N_5371,N_1288,N_1617);
nand U5372 (N_5372,N_4553,N_1376);
nand U5373 (N_5373,N_2137,N_3366);
xnor U5374 (N_5374,N_1935,N_2817);
and U5375 (N_5375,N_2306,N_4107);
xnor U5376 (N_5376,N_807,N_3941);
nor U5377 (N_5377,N_1139,N_4232);
and U5378 (N_5378,N_2016,N_2216);
xnor U5379 (N_5379,N_4819,N_240);
nand U5380 (N_5380,N_3358,N_983);
or U5381 (N_5381,N_2830,N_3439);
xor U5382 (N_5382,N_3934,N_4135);
nand U5383 (N_5383,N_3295,N_820);
and U5384 (N_5384,N_4640,N_2511);
nor U5385 (N_5385,N_3673,N_389);
xnor U5386 (N_5386,N_2564,N_3270);
or U5387 (N_5387,N_2984,N_36);
nand U5388 (N_5388,N_626,N_361);
nor U5389 (N_5389,N_2560,N_668);
and U5390 (N_5390,N_4710,N_942);
or U5391 (N_5391,N_828,N_4490);
and U5392 (N_5392,N_1445,N_2980);
and U5393 (N_5393,N_3800,N_4341);
nand U5394 (N_5394,N_1670,N_1303);
nor U5395 (N_5395,N_115,N_681);
and U5396 (N_5396,N_336,N_2711);
and U5397 (N_5397,N_3818,N_976);
nor U5398 (N_5398,N_793,N_3778);
xnor U5399 (N_5399,N_944,N_3155);
nand U5400 (N_5400,N_2373,N_1319);
and U5401 (N_5401,N_2082,N_4124);
nor U5402 (N_5402,N_4396,N_3077);
or U5403 (N_5403,N_2832,N_4335);
xnor U5404 (N_5404,N_863,N_4950);
or U5405 (N_5405,N_4508,N_1368);
xor U5406 (N_5406,N_2491,N_3336);
and U5407 (N_5407,N_2188,N_688);
xor U5408 (N_5408,N_2812,N_4162);
or U5409 (N_5409,N_2996,N_3025);
nand U5410 (N_5410,N_2667,N_2115);
or U5411 (N_5411,N_1129,N_4609);
nor U5412 (N_5412,N_399,N_3002);
nand U5413 (N_5413,N_2056,N_3158);
and U5414 (N_5414,N_2571,N_845);
and U5415 (N_5415,N_4148,N_3836);
nor U5416 (N_5416,N_905,N_4024);
or U5417 (N_5417,N_1869,N_218);
xnor U5418 (N_5418,N_4390,N_3787);
nor U5419 (N_5419,N_2089,N_3388);
and U5420 (N_5420,N_2002,N_2827);
or U5421 (N_5421,N_4739,N_4380);
nand U5422 (N_5422,N_3309,N_3761);
nor U5423 (N_5423,N_2544,N_4196);
nor U5424 (N_5424,N_3644,N_1272);
xnor U5425 (N_5425,N_1447,N_639);
xnor U5426 (N_5426,N_1273,N_200);
nor U5427 (N_5427,N_4579,N_1962);
and U5428 (N_5428,N_34,N_1579);
or U5429 (N_5429,N_4176,N_1918);
and U5430 (N_5430,N_1727,N_3483);
or U5431 (N_5431,N_4789,N_933);
or U5432 (N_5432,N_2359,N_4150);
nor U5433 (N_5433,N_2686,N_2189);
xnor U5434 (N_5434,N_1115,N_4467);
or U5435 (N_5435,N_634,N_3144);
nor U5436 (N_5436,N_4801,N_4338);
xnor U5437 (N_5437,N_4763,N_134);
nor U5438 (N_5438,N_4717,N_286);
nor U5439 (N_5439,N_3337,N_3582);
nand U5440 (N_5440,N_4699,N_4178);
xor U5441 (N_5441,N_1920,N_992);
or U5442 (N_5442,N_1514,N_3107);
nand U5443 (N_5443,N_2580,N_3845);
nand U5444 (N_5444,N_4962,N_2133);
nor U5445 (N_5445,N_4367,N_4433);
nor U5446 (N_5446,N_4561,N_734);
nor U5447 (N_5447,N_773,N_2977);
nand U5448 (N_5448,N_1173,N_3015);
and U5449 (N_5449,N_2874,N_413);
or U5450 (N_5450,N_1884,N_3837);
nor U5451 (N_5451,N_4566,N_4666);
and U5452 (N_5452,N_2816,N_1030);
or U5453 (N_5453,N_4281,N_2153);
and U5454 (N_5454,N_3064,N_2266);
nand U5455 (N_5455,N_3040,N_1324);
nor U5456 (N_5456,N_799,N_743);
xor U5457 (N_5457,N_2249,N_4991);
xor U5458 (N_5458,N_2556,N_3588);
and U5459 (N_5459,N_170,N_2467);
nor U5460 (N_5460,N_4799,N_774);
xor U5461 (N_5461,N_1055,N_1922);
nand U5462 (N_5462,N_2758,N_2871);
nand U5463 (N_5463,N_4887,N_991);
or U5464 (N_5464,N_904,N_2629);
nor U5465 (N_5465,N_2447,N_1976);
or U5466 (N_5466,N_4811,N_301);
or U5467 (N_5467,N_2501,N_3172);
and U5468 (N_5468,N_39,N_1560);
nand U5469 (N_5469,N_3032,N_3897);
nor U5470 (N_5470,N_3239,N_4925);
nor U5471 (N_5471,N_3342,N_1542);
and U5472 (N_5472,N_3314,N_1228);
nand U5473 (N_5473,N_3622,N_1494);
and U5474 (N_5474,N_425,N_3353);
xor U5475 (N_5475,N_441,N_1050);
and U5476 (N_5476,N_897,N_148);
nand U5477 (N_5477,N_172,N_467);
or U5478 (N_5478,N_2053,N_2583);
xor U5479 (N_5479,N_1652,N_3215);
nor U5480 (N_5480,N_2952,N_3931);
xnor U5481 (N_5481,N_1673,N_19);
xnor U5482 (N_5482,N_926,N_4867);
nor U5483 (N_5483,N_1703,N_2649);
nor U5484 (N_5484,N_3963,N_3690);
nand U5485 (N_5485,N_592,N_3480);
nand U5486 (N_5486,N_312,N_2038);
or U5487 (N_5487,N_958,N_4778);
or U5488 (N_5488,N_4019,N_3789);
nand U5489 (N_5489,N_1671,N_1309);
or U5490 (N_5490,N_4397,N_613);
or U5491 (N_5491,N_3231,N_4085);
nand U5492 (N_5492,N_3367,N_3549);
xnor U5493 (N_5493,N_3720,N_4723);
nor U5494 (N_5494,N_292,N_3249);
and U5495 (N_5495,N_1122,N_31);
nor U5496 (N_5496,N_543,N_3694);
nor U5497 (N_5497,N_2805,N_3572);
and U5498 (N_5498,N_732,N_2105);
and U5499 (N_5499,N_1331,N_1983);
or U5500 (N_5500,N_3974,N_121);
nor U5501 (N_5501,N_2187,N_1946);
xor U5502 (N_5502,N_1465,N_304);
or U5503 (N_5503,N_3119,N_4103);
or U5504 (N_5504,N_524,N_1352);
or U5505 (N_5505,N_3806,N_2751);
and U5506 (N_5506,N_2069,N_2226);
xnor U5507 (N_5507,N_1566,N_2577);
or U5508 (N_5508,N_3777,N_2203);
and U5509 (N_5509,N_4886,N_2303);
xnor U5510 (N_5510,N_4967,N_4117);
and U5511 (N_5511,N_3613,N_703);
and U5512 (N_5512,N_2211,N_3140);
and U5513 (N_5513,N_2684,N_3579);
and U5514 (N_5514,N_1100,N_1383);
and U5515 (N_5515,N_554,N_591);
xor U5516 (N_5516,N_4580,N_4558);
xnor U5517 (N_5517,N_2916,N_865);
nand U5518 (N_5518,N_1855,N_683);
nor U5519 (N_5519,N_1216,N_4572);
nor U5520 (N_5520,N_1537,N_438);
xnor U5521 (N_5521,N_372,N_2487);
or U5522 (N_5522,N_4726,N_4437);
or U5523 (N_5523,N_1320,N_3381);
nor U5524 (N_5524,N_2443,N_314);
or U5525 (N_5525,N_652,N_2088);
or U5526 (N_5526,N_195,N_664);
xor U5527 (N_5527,N_2968,N_810);
nor U5528 (N_5528,N_2472,N_4732);
nor U5529 (N_5529,N_3089,N_3597);
nor U5530 (N_5530,N_2988,N_998);
nand U5531 (N_5531,N_4479,N_4638);
xnor U5532 (N_5532,N_1893,N_520);
xor U5533 (N_5533,N_4250,N_886);
xor U5534 (N_5534,N_2095,N_4434);
and U5535 (N_5535,N_4419,N_3453);
nand U5536 (N_5536,N_3069,N_4483);
nor U5537 (N_5537,N_1371,N_3609);
and U5538 (N_5538,N_4695,N_1531);
xor U5539 (N_5539,N_3870,N_1997);
and U5540 (N_5540,N_2887,N_2747);
or U5541 (N_5541,N_4782,N_563);
or U5542 (N_5542,N_3001,N_885);
nand U5543 (N_5543,N_3502,N_1947);
and U5544 (N_5544,N_785,N_1578);
and U5545 (N_5545,N_2508,N_1852);
nand U5546 (N_5546,N_4182,N_4283);
or U5547 (N_5547,N_3413,N_995);
nor U5548 (N_5548,N_736,N_1732);
and U5549 (N_5549,N_1170,N_2702);
and U5550 (N_5550,N_1607,N_589);
or U5551 (N_5551,N_3188,N_3088);
nand U5552 (N_5552,N_2923,N_655);
nor U5553 (N_5553,N_3898,N_2550);
xnor U5554 (N_5554,N_1661,N_505);
nand U5555 (N_5555,N_2552,N_6);
and U5556 (N_5556,N_1016,N_2671);
xor U5557 (N_5557,N_223,N_3936);
and U5558 (N_5558,N_2426,N_4424);
nor U5559 (N_5559,N_1906,N_1184);
and U5560 (N_5560,N_1158,N_315);
or U5561 (N_5561,N_385,N_4542);
nor U5562 (N_5562,N_945,N_999);
and U5563 (N_5563,N_3482,N_4128);
and U5564 (N_5564,N_2584,N_812);
and U5565 (N_5565,N_4074,N_275);
nor U5566 (N_5566,N_2835,N_1283);
xor U5567 (N_5567,N_3233,N_1120);
nor U5568 (N_5568,N_4009,N_2323);
nand U5569 (N_5569,N_1057,N_3524);
or U5570 (N_5570,N_3520,N_993);
and U5571 (N_5571,N_2754,N_3130);
nand U5572 (N_5572,N_2463,N_4942);
nor U5573 (N_5573,N_1896,N_3729);
and U5574 (N_5574,N_3078,N_3616);
xor U5575 (N_5575,N_1699,N_4484);
nand U5576 (N_5576,N_2416,N_4842);
xnor U5577 (N_5577,N_2409,N_4704);
and U5578 (N_5578,N_2200,N_264);
nor U5579 (N_5579,N_1390,N_2397);
and U5580 (N_5580,N_4227,N_556);
nor U5581 (N_5581,N_1576,N_2548);
nand U5582 (N_5582,N_2402,N_2784);
nand U5583 (N_5583,N_1382,N_1099);
xor U5584 (N_5584,N_4994,N_4779);
or U5585 (N_5585,N_4588,N_3591);
nand U5586 (N_5586,N_1858,N_4964);
or U5587 (N_5587,N_3320,N_490);
nand U5588 (N_5588,N_4606,N_4013);
nor U5589 (N_5589,N_829,N_4767);
or U5590 (N_5590,N_3606,N_2739);
nand U5591 (N_5591,N_3528,N_1660);
and U5592 (N_5592,N_273,N_2140);
nor U5593 (N_5593,N_4665,N_4873);
and U5594 (N_5594,N_1779,N_881);
nand U5595 (N_5595,N_4366,N_3341);
and U5596 (N_5596,N_4625,N_3891);
nand U5597 (N_5597,N_3620,N_802);
and U5598 (N_5598,N_1101,N_2166);
or U5599 (N_5599,N_2910,N_1214);
nor U5600 (N_5600,N_255,N_3771);
nand U5601 (N_5601,N_3759,N_2380);
xor U5602 (N_5602,N_3146,N_4904);
xor U5603 (N_5603,N_851,N_1080);
or U5604 (N_5604,N_227,N_3619);
nor U5605 (N_5605,N_499,N_2030);
nor U5606 (N_5606,N_2699,N_4783);
nand U5607 (N_5607,N_910,N_714);
or U5608 (N_5608,N_266,N_501);
nor U5609 (N_5609,N_2247,N_4708);
nor U5610 (N_5610,N_866,N_4574);
nor U5611 (N_5611,N_3719,N_1460);
nand U5612 (N_5612,N_3044,N_4822);
nor U5613 (N_5613,N_260,N_2714);
nor U5614 (N_5614,N_4584,N_3652);
nor U5615 (N_5615,N_1182,N_3325);
nand U5616 (N_5616,N_679,N_3074);
and U5617 (N_5617,N_2351,N_594);
and U5618 (N_5618,N_3245,N_179);
or U5619 (N_5619,N_4378,N_2349);
nor U5620 (N_5620,N_3663,N_4092);
and U5621 (N_5621,N_2429,N_832);
or U5622 (N_5622,N_2111,N_1984);
nand U5623 (N_5623,N_4099,N_3548);
or U5624 (N_5624,N_1711,N_4555);
and U5625 (N_5625,N_947,N_4828);
and U5626 (N_5626,N_1148,N_1871);
or U5627 (N_5627,N_972,N_1282);
xnor U5628 (N_5628,N_4220,N_1096);
or U5629 (N_5629,N_1975,N_1138);
or U5630 (N_5630,N_4,N_4290);
nand U5631 (N_5631,N_3334,N_2528);
or U5632 (N_5632,N_3083,N_1754);
or U5633 (N_5633,N_1767,N_1863);
or U5634 (N_5634,N_4455,N_3175);
nand U5635 (N_5635,N_1118,N_1640);
or U5636 (N_5636,N_3305,N_2607);
nand U5637 (N_5637,N_2886,N_4264);
or U5638 (N_5638,N_830,N_767);
xor U5639 (N_5639,N_4803,N_4537);
and U5640 (N_5640,N_4773,N_2217);
or U5641 (N_5641,N_1164,N_186);
nor U5642 (N_5642,N_3852,N_4064);
nand U5643 (N_5643,N_1815,N_495);
xnor U5644 (N_5644,N_345,N_540);
and U5645 (N_5645,N_3860,N_3244);
nor U5646 (N_5646,N_3989,N_3151);
or U5647 (N_5647,N_3752,N_1359);
xor U5648 (N_5648,N_2026,N_3724);
nor U5649 (N_5649,N_2776,N_1669);
and U5650 (N_5650,N_572,N_340);
or U5651 (N_5651,N_4745,N_349);
xnor U5652 (N_5652,N_4192,N_4171);
nor U5653 (N_5653,N_3604,N_2142);
xor U5654 (N_5654,N_2461,N_2434);
nand U5655 (N_5655,N_2308,N_1695);
and U5656 (N_5656,N_4812,N_3056);
nor U5657 (N_5657,N_735,N_690);
or U5658 (N_5658,N_777,N_2915);
and U5659 (N_5659,N_398,N_3948);
nor U5660 (N_5660,N_4525,N_4945);
and U5661 (N_5661,N_770,N_3889);
nand U5662 (N_5662,N_4246,N_42);
nand U5663 (N_5663,N_779,N_803);
or U5664 (N_5664,N_2256,N_3766);
and U5665 (N_5665,N_2958,N_2043);
and U5666 (N_5666,N_118,N_4540);
and U5667 (N_5667,N_1294,N_4509);
nor U5668 (N_5668,N_1741,N_2542);
nor U5669 (N_5669,N_3331,N_721);
nand U5670 (N_5670,N_4506,N_3208);
xor U5671 (N_5671,N_2280,N_422);
nand U5672 (N_5672,N_587,N_3508);
nor U5673 (N_5673,N_2044,N_1925);
or U5674 (N_5674,N_1085,N_2525);
or U5675 (N_5675,N_2098,N_2352);
or U5676 (N_5676,N_1713,N_2496);
nand U5677 (N_5677,N_641,N_1701);
nand U5678 (N_5678,N_1160,N_1475);
and U5679 (N_5679,N_242,N_504);
nor U5680 (N_5680,N_4003,N_4947);
and U5681 (N_5681,N_4816,N_298);
xor U5682 (N_5682,N_3895,N_1724);
nor U5683 (N_5683,N_2715,N_1234);
nor U5684 (N_5684,N_4531,N_3184);
or U5685 (N_5685,N_2897,N_69);
nand U5686 (N_5686,N_2460,N_2360);
and U5687 (N_5687,N_4422,N_754);
or U5688 (N_5688,N_4677,N_4897);
nand U5689 (N_5689,N_2415,N_4460);
or U5690 (N_5690,N_2543,N_2492);
nor U5691 (N_5691,N_1828,N_4989);
and U5692 (N_5692,N_2748,N_2225);
or U5693 (N_5693,N_693,N_414);
nand U5694 (N_5694,N_4173,N_2059);
xor U5695 (N_5695,N_3552,N_617);
or U5696 (N_5696,N_874,N_1195);
and U5697 (N_5697,N_400,N_4893);
or U5698 (N_5698,N_1255,N_2190);
xor U5699 (N_5699,N_4321,N_1492);
or U5700 (N_5700,N_1426,N_4443);
or U5701 (N_5701,N_1403,N_4235);
nand U5702 (N_5702,N_3736,N_3436);
or U5703 (N_5703,N_3750,N_1049);
or U5704 (N_5704,N_2108,N_771);
or U5705 (N_5705,N_4899,N_4858);
or U5706 (N_5706,N_686,N_1462);
and U5707 (N_5707,N_654,N_1765);
nor U5708 (N_5708,N_2565,N_4159);
nand U5709 (N_5709,N_1936,N_4619);
or U5710 (N_5710,N_2640,N_1608);
nor U5711 (N_5711,N_3712,N_1318);
and U5712 (N_5712,N_2456,N_1964);
and U5713 (N_5713,N_583,N_2695);
or U5714 (N_5714,N_868,N_545);
or U5715 (N_5715,N_3007,N_4775);
or U5716 (N_5716,N_847,N_4924);
nor U5717 (N_5717,N_87,N_3674);
nor U5718 (N_5718,N_2424,N_887);
nor U5719 (N_5719,N_670,N_1974);
nand U5720 (N_5720,N_1186,N_2304);
nand U5721 (N_5721,N_3534,N_3683);
nand U5722 (N_5722,N_2829,N_1960);
nand U5723 (N_5723,N_902,N_1346);
nand U5724 (N_5724,N_1028,N_4517);
xnor U5725 (N_5725,N_1071,N_751);
and U5726 (N_5726,N_2036,N_4068);
xnor U5727 (N_5727,N_2760,N_2093);
and U5728 (N_5728,N_3060,N_3444);
xor U5729 (N_5729,N_1092,N_4992);
and U5730 (N_5730,N_4154,N_2168);
and U5731 (N_5731,N_2361,N_173);
nor U5732 (N_5732,N_4365,N_4888);
or U5733 (N_5733,N_2431,N_608);
nand U5734 (N_5734,N_3046,N_2840);
nand U5735 (N_5735,N_2994,N_4821);
nor U5736 (N_5736,N_4047,N_3815);
or U5737 (N_5737,N_644,N_1452);
xnor U5738 (N_5738,N_1045,N_3880);
nor U5739 (N_5739,N_1843,N_4413);
nand U5740 (N_5740,N_1613,N_1197);
nor U5741 (N_5741,N_3456,N_1522);
and U5742 (N_5742,N_2417,N_575);
nand U5743 (N_5743,N_4857,N_3441);
nand U5744 (N_5744,N_3326,N_3995);
xor U5745 (N_5745,N_2792,N_4012);
nor U5746 (N_5746,N_1499,N_1839);
nand U5747 (N_5747,N_88,N_1411);
and U5748 (N_5748,N_3976,N_3790);
xnor U5749 (N_5749,N_3969,N_420);
or U5750 (N_5750,N_2932,N_2233);
and U5751 (N_5751,N_4342,N_3059);
xnor U5752 (N_5752,N_2332,N_4769);
nor U5753 (N_5753,N_2039,N_1509);
nand U5754 (N_5754,N_2338,N_2878);
and U5755 (N_5755,N_3696,N_1404);
and U5756 (N_5756,N_3023,N_862);
and U5757 (N_5757,N_4063,N_4194);
nand U5758 (N_5758,N_16,N_460);
nand U5759 (N_5759,N_2680,N_1757);
nor U5760 (N_5760,N_955,N_2422);
nand U5761 (N_5761,N_3153,N_4444);
and U5762 (N_5762,N_837,N_879);
xor U5763 (N_5763,N_4911,N_3018);
or U5764 (N_5764,N_1198,N_357);
nand U5765 (N_5765,N_3228,N_2198);
and U5766 (N_5766,N_4850,N_3122);
nor U5767 (N_5767,N_2713,N_2974);
nand U5768 (N_5768,N_1958,N_3899);
xor U5769 (N_5769,N_2669,N_3740);
and U5770 (N_5770,N_511,N_3345);
nand U5771 (N_5771,N_1620,N_4895);
and U5772 (N_5772,N_366,N_1450);
xnor U5773 (N_5773,N_2908,N_3214);
and U5774 (N_5774,N_1275,N_1939);
nor U5775 (N_5775,N_2295,N_2489);
xnor U5776 (N_5776,N_392,N_3840);
nor U5777 (N_5777,N_598,N_4403);
or U5778 (N_5778,N_899,N_1312);
nand U5779 (N_5779,N_4231,N_1742);
nor U5780 (N_5780,N_1023,N_21);
or U5781 (N_5781,N_2570,N_3768);
xor U5782 (N_5782,N_2334,N_4718);
nor U5783 (N_5783,N_25,N_1014);
nor U5784 (N_5784,N_1510,N_4187);
or U5785 (N_5785,N_1277,N_547);
and U5786 (N_5786,N_3971,N_1914);
and U5787 (N_5787,N_3062,N_395);
nor U5788 (N_5788,N_4979,N_4733);
xnor U5789 (N_5789,N_1202,N_3730);
nand U5790 (N_5790,N_1396,N_1851);
nor U5791 (N_5791,N_4363,N_4571);
or U5792 (N_5792,N_2421,N_1880);
xnor U5793 (N_5793,N_4224,N_164);
nand U5794 (N_5794,N_3094,N_4084);
nor U5795 (N_5795,N_559,N_103);
nand U5796 (N_5796,N_1032,N_1956);
xor U5797 (N_5797,N_3583,N_1749);
and U5798 (N_5798,N_2946,N_2925);
nor U5799 (N_5799,N_2985,N_3428);
nor U5800 (N_5800,N_3211,N_1725);
nor U5801 (N_5801,N_3418,N_4690);
nand U5802 (N_5802,N_4815,N_824);
nor U5803 (N_5803,N_1310,N_1137);
nor U5804 (N_5804,N_4689,N_4532);
nand U5805 (N_5805,N_1970,N_2112);
nor U5806 (N_5806,N_3398,N_1013);
or U5807 (N_5807,N_2722,N_1800);
xor U5808 (N_5808,N_1325,N_4524);
or U5809 (N_5809,N_74,N_2731);
nand U5810 (N_5810,N_3762,N_3135);
and U5811 (N_5811,N_2757,N_2644);
nor U5812 (N_5812,N_2305,N_2040);
nand U5813 (N_5813,N_786,N_4184);
xnor U5814 (N_5814,N_2367,N_4302);
nor U5815 (N_5815,N_728,N_4682);
xnor U5816 (N_5816,N_4268,N_3392);
nand U5817 (N_5817,N_2594,N_3143);
and U5818 (N_5818,N_4057,N_720);
or U5819 (N_5819,N_4891,N_2738);
and U5820 (N_5820,N_2310,N_3907);
or U5821 (N_5821,N_4447,N_3157);
nor U5822 (N_5822,N_2516,N_4285);
nand U5823 (N_5823,N_1866,N_4045);
or U5824 (N_5824,N_2276,N_1221);
xor U5825 (N_5825,N_602,N_162);
nor U5826 (N_5826,N_2979,N_4759);
nand U5827 (N_5827,N_1175,N_581);
and U5828 (N_5828,N_3560,N_2301);
xnor U5829 (N_5829,N_4177,N_183);
xor U5830 (N_5830,N_974,N_1533);
xnor U5831 (N_5831,N_356,N_380);
nor U5832 (N_5832,N_1305,N_787);
and U5833 (N_5833,N_150,N_4432);
nor U5834 (N_5834,N_3177,N_1552);
nor U5835 (N_5835,N_508,N_358);
and U5836 (N_5836,N_2471,N_1894);
xor U5837 (N_5837,N_2328,N_1066);
xor U5838 (N_5838,N_219,N_4306);
or U5839 (N_5839,N_4097,N_276);
nor U5840 (N_5840,N_1902,N_3033);
nand U5841 (N_5841,N_3671,N_4834);
nand U5842 (N_5842,N_3717,N_1513);
and U5843 (N_5843,N_57,N_3821);
and U5844 (N_5844,N_4720,N_2437);
nor U5845 (N_5845,N_1291,N_4382);
and U5846 (N_5846,N_2451,N_194);
or U5847 (N_5847,N_1524,N_677);
or U5848 (N_5848,N_1209,N_128);
nor U5849 (N_5849,N_4790,N_4959);
and U5850 (N_5850,N_332,N_2076);
nand U5851 (N_5851,N_840,N_4464);
and U5852 (N_5852,N_542,N_449);
nor U5853 (N_5853,N_231,N_1549);
or U5854 (N_5854,N_4694,N_225);
and U5855 (N_5855,N_2458,N_860);
nor U5856 (N_5856,N_2220,N_3169);
xor U5857 (N_5857,N_4056,N_2330);
and U5858 (N_5858,N_2843,N_1490);
or U5859 (N_5859,N_3123,N_3055);
nand U5860 (N_5860,N_4282,N_4190);
and U5861 (N_5861,N_1834,N_3704);
nor U5862 (N_5862,N_3152,N_4678);
nor U5863 (N_5863,N_3393,N_3210);
nor U5864 (N_5864,N_2412,N_3464);
xor U5865 (N_5865,N_4070,N_1708);
nand U5866 (N_5866,N_2484,N_241);
or U5867 (N_5867,N_1215,N_169);
or U5868 (N_5868,N_2094,N_4841);
nor U5869 (N_5869,N_4420,N_1022);
and U5870 (N_5870,N_368,N_890);
nand U5871 (N_5871,N_4518,N_2726);
nor U5872 (N_5872,N_3183,N_3246);
nand U5873 (N_5873,N_196,N_3573);
nand U5874 (N_5874,N_2682,N_2466);
xnor U5875 (N_5875,N_4487,N_3734);
nand U5876 (N_5876,N_4002,N_3356);
nor U5877 (N_5877,N_1086,N_232);
nor U5878 (N_5878,N_850,N_3594);
xnor U5879 (N_5879,N_919,N_117);
xnor U5880 (N_5880,N_658,N_3126);
or U5881 (N_5881,N_3567,N_562);
nand U5882 (N_5882,N_1758,N_2819);
and U5883 (N_5883,N_4987,N_618);
nand U5884 (N_5884,N_145,N_265);
nor U5885 (N_5885,N_2202,N_809);
xnor U5886 (N_5886,N_1585,N_1375);
and U5887 (N_5887,N_4914,N_277);
and U5888 (N_5888,N_4851,N_3095);
nand U5889 (N_5889,N_3558,N_2517);
or U5890 (N_5890,N_479,N_4495);
nand U5891 (N_5891,N_2928,N_1140);
nand U5892 (N_5892,N_719,N_339);
and U5893 (N_5893,N_4119,N_917);
xor U5894 (N_5894,N_2278,N_4656);
nor U5895 (N_5895,N_4348,N_1781);
xor U5896 (N_5896,N_1226,N_1289);
or U5897 (N_5897,N_2240,N_1595);
nor U5898 (N_5898,N_3713,N_4352);
nor U5899 (N_5899,N_3580,N_3271);
or U5900 (N_5900,N_2023,N_2164);
xnor U5901 (N_5901,N_1339,N_3332);
and U5902 (N_5902,N_625,N_2012);
or U5903 (N_5903,N_470,N_1504);
xor U5904 (N_5904,N_4421,N_3405);
nor U5905 (N_5905,N_4463,N_2474);
or U5906 (N_5906,N_1194,N_2611);
xor U5907 (N_5907,N_1891,N_4501);
and U5908 (N_5908,N_2371,N_903);
xor U5909 (N_5909,N_1795,N_2703);
xnor U5910 (N_5910,N_3675,N_3052);
nand U5911 (N_5911,N_4806,N_3310);
nand U5912 (N_5912,N_4798,N_3797);
and U5913 (N_5913,N_1647,N_3471);
nand U5914 (N_5914,N_1245,N_2464);
and U5915 (N_5915,N_3306,N_2641);
nor U5916 (N_5916,N_4145,N_1905);
and U5917 (N_5917,N_3823,N_2382);
xnor U5918 (N_5918,N_805,N_2480);
nor U5919 (N_5919,N_308,N_3159);
nor U5920 (N_5920,N_3396,N_4889);
xor U5921 (N_5921,N_3145,N_2636);
xor U5922 (N_5922,N_1979,N_2951);
nor U5923 (N_5923,N_4534,N_4657);
xor U5924 (N_5924,N_2956,N_4549);
or U5925 (N_5925,N_1555,N_1929);
nor U5926 (N_5926,N_775,N_1730);
or U5927 (N_5927,N_1653,N_3611);
xor U5928 (N_5928,N_3601,N_2582);
nor U5929 (N_5929,N_4258,N_2943);
and U5930 (N_5930,N_4211,N_3672);
nor U5931 (N_5931,N_1753,N_1840);
nand U5932 (N_5932,N_2231,N_1686);
and U5933 (N_5933,N_4853,N_3955);
xnor U5934 (N_5934,N_78,N_1605);
nor U5935 (N_5935,N_814,N_2706);
nor U5936 (N_5936,N_75,N_1087);
nand U5937 (N_5937,N_1646,N_2872);
or U5938 (N_5938,N_2708,N_4687);
nand U5939 (N_5939,N_3105,N_570);
nor U5940 (N_5940,N_1790,N_3238);
or U5941 (N_5941,N_3042,N_408);
nand U5942 (N_5942,N_3689,N_2152);
or U5943 (N_5943,N_1544,N_3518);
xnor U5944 (N_5944,N_2677,N_4216);
nand U5945 (N_5945,N_2212,N_3391);
xor U5946 (N_5946,N_3058,N_3912);
nor U5947 (N_5947,N_4175,N_3112);
and U5948 (N_5948,N_1307,N_216);
nor U5949 (N_5949,N_1223,N_4780);
nand U5950 (N_5950,N_2842,N_480);
or U5951 (N_5951,N_1285,N_3543);
nor U5952 (N_5952,N_397,N_3125);
nor U5953 (N_5953,N_3262,N_4713);
nor U5954 (N_5954,N_4228,N_4714);
xnor U5955 (N_5955,N_3484,N_704);
and U5956 (N_5956,N_4133,N_4393);
xnor U5957 (N_5957,N_62,N_1625);
xor U5958 (N_5958,N_661,N_3203);
or U5959 (N_5959,N_3763,N_1931);
nand U5960 (N_5960,N_1882,N_3440);
and U5961 (N_5961,N_1188,N_37);
or U5962 (N_5962,N_1105,N_4844);
nor U5963 (N_5963,N_2366,N_4802);
or U5964 (N_5964,N_3770,N_96);
nor U5965 (N_5965,N_3798,N_4592);
xor U5966 (N_5966,N_1952,N_4652);
nand U5967 (N_5967,N_1930,N_1917);
nor U5968 (N_5968,N_3226,N_2989);
nand U5969 (N_5969,N_2746,N_1688);
nor U5970 (N_5970,N_3915,N_229);
and U5971 (N_5971,N_2595,N_3086);
nand U5972 (N_5972,N_697,N_4754);
nand U5973 (N_5973,N_2796,N_2553);
nand U5974 (N_5974,N_1648,N_2883);
or U5975 (N_5975,N_2343,N_1623);
xnor U5976 (N_5976,N_3833,N_1908);
or U5977 (N_5977,N_1218,N_3000);
nand U5978 (N_5978,N_521,N_953);
and U5979 (N_5979,N_896,N_4461);
or U5980 (N_5980,N_4140,N_2486);
nor U5981 (N_5981,N_1799,N_2536);
nor U5982 (N_5982,N_1463,N_3091);
nor U5983 (N_5983,N_3137,N_827);
nor U5984 (N_5984,N_1212,N_4036);
and U5985 (N_5985,N_383,N_1058);
or U5986 (N_5986,N_1618,N_2926);
and U5987 (N_5987,N_4831,N_4774);
nand U5988 (N_5988,N_2647,N_665);
nand U5989 (N_5989,N_4896,N_2128);
or U5990 (N_5990,N_4337,N_151);
or U5991 (N_5991,N_2176,N_1938);
or U5992 (N_5992,N_1060,N_1847);
and U5993 (N_5993,N_2608,N_937);
xor U5994 (N_5994,N_2862,N_296);
or U5995 (N_5995,N_638,N_155);
xnor U5996 (N_5996,N_274,N_726);
and U5997 (N_5997,N_853,N_1803);
nand U5998 (N_5998,N_4462,N_4547);
nor U5999 (N_5999,N_1760,N_1639);
or U6000 (N_6000,N_4311,N_1338);
nor U6001 (N_6001,N_1172,N_485);
xor U6002 (N_6002,N_3825,N_2368);
nand U6003 (N_6003,N_710,N_1123);
nor U6004 (N_6004,N_2283,N_2743);
nor U6005 (N_6005,N_4777,N_245);
and U6006 (N_6006,N_869,N_4010);
nor U6007 (N_6007,N_2678,N_2025);
and U6008 (N_6008,N_3224,N_3034);
xor U6009 (N_6009,N_2558,N_963);
nand U6010 (N_6010,N_5,N_3009);
or U6011 (N_6011,N_3600,N_1659);
nor U6012 (N_6012,N_3340,N_1841);
xnor U6013 (N_6013,N_1480,N_2613);
nand U6014 (N_6014,N_2507,N_3038);
xor U6015 (N_6015,N_3114,N_694);
or U6016 (N_6016,N_3856,N_3035);
nand U6017 (N_6017,N_3598,N_1340);
and U6018 (N_6018,N_4751,N_3758);
nor U6019 (N_6019,N_1256,N_811);
or U6020 (N_6020,N_379,N_1110);
nand U6021 (N_6021,N_2638,N_806);
and U6022 (N_6022,N_3330,N_2478);
nor U6023 (N_6023,N_3503,N_26);
nand U6024 (N_6024,N_3749,N_4174);
nand U6025 (N_6025,N_3161,N_202);
and U6026 (N_6026,N_675,N_636);
or U6027 (N_6027,N_190,N_364);
nand U6028 (N_6028,N_1199,N_1538);
nand U6029 (N_6029,N_3476,N_3883);
nor U6030 (N_6030,N_4906,N_377);
xor U6031 (N_6031,N_1642,N_1584);
nor U6032 (N_6032,N_3474,N_4766);
and U6033 (N_6033,N_175,N_4881);
xor U6034 (N_6034,N_127,N_4500);
nand U6035 (N_6035,N_1082,N_1192);
xnor U6036 (N_6036,N_1567,N_3769);
xnor U6037 (N_6037,N_3557,N_497);
xor U6038 (N_6038,N_2742,N_4650);
nand U6039 (N_6039,N_4876,N_4204);
xor U6040 (N_6040,N_1193,N_4533);
nand U6041 (N_6041,N_952,N_2064);
nand U6042 (N_6042,N_901,N_1526);
xnor U6043 (N_6043,N_878,N_580);
xor U6044 (N_6044,N_3925,N_3422);
xnor U6045 (N_6045,N_1398,N_2683);
xor U6046 (N_6046,N_922,N_158);
xor U6047 (N_6047,N_893,N_1369);
nand U6048 (N_6048,N_4053,N_2870);
or U6049 (N_6049,N_3485,N_1563);
nor U6050 (N_6050,N_2125,N_224);
or U6051 (N_6051,N_2418,N_530);
nor U6052 (N_6052,N_997,N_4156);
and U6053 (N_6053,N_2399,N_2975);
nand U6054 (N_6054,N_629,N_4354);
xnor U6055 (N_6055,N_4046,N_1363);
nand U6056 (N_6056,N_921,N_3532);
nor U6057 (N_6057,N_1141,N_2772);
xnor U6058 (N_6058,N_1069,N_3442);
nor U6059 (N_6059,N_1008,N_334);
nand U6060 (N_6060,N_3462,N_423);
or U6061 (N_6061,N_848,N_3527);
nor U6062 (N_6062,N_1116,N_1515);
nand U6063 (N_6063,N_2254,N_1737);
nor U6064 (N_6064,N_936,N_3827);
or U6065 (N_6065,N_198,N_1911);
nand U6066 (N_6066,N_2725,N_4257);
and U6067 (N_6067,N_2612,N_125);
nor U6068 (N_6068,N_1263,N_2893);
or U6069 (N_6069,N_2369,N_2224);
or U6070 (N_6070,N_1395,N_3333);
nand U6071 (N_6071,N_4629,N_3201);
xor U6072 (N_6072,N_3373,N_4539);
or U6073 (N_6073,N_971,N_394);
or U6074 (N_6074,N_2252,N_1644);
xnor U6075 (N_6075,N_2578,N_45);
xnor U6076 (N_6076,N_2139,N_4123);
nor U6077 (N_6077,N_4288,N_3093);
and U6078 (N_6078,N_201,N_1775);
or U6079 (N_6079,N_1955,N_4636);
nor U6080 (N_6080,N_2384,N_3313);
nor U6081 (N_6081,N_1179,N_419);
or U6082 (N_6082,N_2258,N_3377);
or U6083 (N_6083,N_3922,N_4223);
or U6084 (N_6084,N_2318,N_1007);
or U6085 (N_6085,N_360,N_1500);
nand U6086 (N_6086,N_3665,N_1987);
and U6087 (N_6087,N_2953,N_1668);
nand U6088 (N_6088,N_790,N_4929);
and U6089 (N_6089,N_4118,N_3865);
or U6090 (N_6090,N_4394,N_4226);
nand U6091 (N_6091,N_4557,N_3920);
and U6092 (N_6092,N_1601,N_342);
nand U6093 (N_6093,N_1818,N_2995);
nor U6094 (N_6094,N_875,N_831);
nand U6095 (N_6095,N_2697,N_4086);
and U6096 (N_6096,N_4622,N_915);
xor U6097 (N_6097,N_2533,N_4144);
xor U6098 (N_6098,N_742,N_4535);
and U6099 (N_6099,N_2960,N_3368);
and U6100 (N_6100,N_70,N_1350);
or U6101 (N_6101,N_2894,N_4040);
or U6102 (N_6102,N_359,N_3493);
xnor U6103 (N_6103,N_4331,N_2087);
xor U6104 (N_6104,N_1473,N_1832);
nand U6105 (N_6105,N_3065,N_4737);
nor U6106 (N_6106,N_889,N_3076);
nand U6107 (N_6107,N_4096,N_3460);
nand U6108 (N_6108,N_1328,N_3383);
and U6109 (N_6109,N_4234,N_585);
nand U6110 (N_6110,N_3653,N_916);
or U6111 (N_6111,N_3202,N_1276);
or U6112 (N_6112,N_2438,N_293);
nor U6113 (N_6113,N_1591,N_1322);
nor U6114 (N_6114,N_1854,N_3012);
nor U6115 (N_6115,N_624,N_4623);
nor U6116 (N_6116,N_489,N_373);
nor U6117 (N_6117,N_4603,N_3293);
nor U6118 (N_6118,N_2518,N_2820);
nand U6119 (N_6119,N_920,N_3655);
xnor U6120 (N_6120,N_577,N_303);
nand U6121 (N_6121,N_1540,N_4102);
or U6122 (N_6122,N_2205,N_941);
nand U6123 (N_6123,N_4293,N_2178);
and U6124 (N_6124,N_4516,N_4949);
or U6125 (N_6125,N_2147,N_3808);
xor U6126 (N_6126,N_3084,N_4214);
or U6127 (N_6127,N_409,N_4890);
and U6128 (N_6128,N_1031,N_4377);
nor U6129 (N_6129,N_1487,N_3841);
and U6130 (N_6130,N_1836,N_442);
xnor U6131 (N_6131,N_3857,N_1043);
xnor U6132 (N_6132,N_4078,N_2196);
and U6133 (N_6133,N_4041,N_3242);
nand U6134 (N_6134,N_1658,N_3603);
or U6135 (N_6135,N_329,N_2701);
or U6136 (N_6136,N_2737,N_4195);
nor U6137 (N_6137,N_2118,N_1516);
nor U6138 (N_6138,N_685,N_3466);
nand U6139 (N_6139,N_3347,N_4212);
and U6140 (N_6140,N_557,N_2892);
and U6141 (N_6141,N_1614,N_1425);
and U6142 (N_6142,N_3410,N_3097);
and U6143 (N_6143,N_560,N_2358);
and U6144 (N_6144,N_1370,N_4642);
or U6145 (N_6145,N_4514,N_3647);
xor U6146 (N_6146,N_2767,N_642);
or U6147 (N_6147,N_2232,N_4445);
or U6148 (N_6148,N_2824,N_1507);
and U6149 (N_6149,N_4705,N_1262);
xor U6150 (N_6150,N_3481,N_1456);
or U6151 (N_6151,N_3839,N_4308);
and U6152 (N_6152,N_3786,N_17);
nand U6153 (N_6153,N_2475,N_2902);
and U6154 (N_6154,N_1707,N_4304);
or U6155 (N_6155,N_3394,N_3426);
xor U6156 (N_6156,N_649,N_680);
nand U6157 (N_6157,N_2337,N_3869);
nand U6158 (N_6158,N_3688,N_2615);
nor U6159 (N_6159,N_2477,N_4653);
nor U6160 (N_6160,N_2065,N_3812);
nand U6161 (N_6161,N_980,N_4391);
nand U6162 (N_6162,N_4275,N_1040);
and U6163 (N_6163,N_1804,N_656);
nor U6164 (N_6164,N_3783,N_4883);
nor U6165 (N_6165,N_3636,N_4229);
xnor U6166 (N_6166,N_1587,N_124);
and U6167 (N_6167,N_4971,N_1257);
xnor U6168 (N_6168,N_2569,N_3645);
xor U6169 (N_6169,N_2022,N_4855);
and U6170 (N_6170,N_4083,N_4746);
and U6171 (N_6171,N_192,N_2439);
nand U6172 (N_6172,N_3926,N_491);
and U6173 (N_6173,N_1178,N_1602);
nor U6174 (N_6174,N_2156,N_2253);
xnor U6175 (N_6175,N_2499,N_4244);
xnor U6176 (N_6176,N_4031,N_4344);
nor U6177 (N_6177,N_44,N_2586);
and U6178 (N_6178,N_2389,N_3677);
and U6179 (N_6179,N_3953,N_764);
nor U6180 (N_6180,N_2700,N_4598);
and U6181 (N_6181,N_2538,N_1027);
nand U6182 (N_6182,N_2290,N_1146);
nand U6183 (N_6183,N_696,N_960);
nand U6184 (N_6184,N_8,N_4385);
nor U6185 (N_6185,N_1996,N_4997);
xnor U6186 (N_6186,N_4672,N_645);
xor U6187 (N_6187,N_3861,N_3063);
or U6188 (N_6188,N_4248,N_3096);
xnor U6189 (N_6189,N_90,N_2289);
nor U6190 (N_6190,N_3277,N_2070);
xnor U6191 (N_6191,N_4669,N_234);
or U6192 (N_6192,N_4611,N_2037);
nand U6193 (N_6193,N_4926,N_894);
nor U6194 (N_6194,N_1313,N_4591);
nand U6195 (N_6195,N_3397,N_1771);
nor U6196 (N_6196,N_2554,N_4218);
and U6197 (N_6197,N_52,N_2959);
xnor U6198 (N_6198,N_895,N_3505);
or U6199 (N_6199,N_3495,N_1941);
nor U6200 (N_6200,N_3164,N_1606);
or U6201 (N_6201,N_1054,N_10);
nor U6202 (N_6202,N_309,N_1017);
xnor U6203 (N_6203,N_4700,N_2031);
or U6204 (N_6204,N_4706,N_99);
nand U6205 (N_6205,N_3913,N_3465);
and U6206 (N_6206,N_2392,N_4750);
xor U6207 (N_6207,N_3701,N_3804);
nand U6208 (N_6208,N_595,N_1599);
or U6209 (N_6209,N_3416,N_2279);
xor U6210 (N_6210,N_2719,N_1654);
nand U6211 (N_6211,N_2274,N_2599);
or U6212 (N_6212,N_3939,N_4015);
nor U6213 (N_6213,N_3221,N_122);
and U6214 (N_6214,N_1994,N_4995);
nor U6215 (N_6215,N_0,N_4569);
or U6216 (N_6216,N_1315,N_393);
nand U6217 (N_6217,N_1366,N_4785);
nand U6218 (N_6218,N_4760,N_4305);
nor U6219 (N_6219,N_1434,N_2898);
or U6220 (N_6220,N_2400,N_434);
and U6221 (N_6221,N_2317,N_4442);
and U6222 (N_6222,N_4126,N_2425);
nand U6223 (N_6223,N_2555,N_84);
nor U6224 (N_6224,N_3110,N_436);
xnor U6225 (N_6225,N_2194,N_4974);
and U6226 (N_6226,N_80,N_1405);
nand U6227 (N_6227,N_1879,N_2299);
nor U6228 (N_6228,N_1971,N_1081);
and U6229 (N_6229,N_3236,N_3129);
and U6230 (N_6230,N_1254,N_20);
or U6231 (N_6231,N_852,N_507);
or U6232 (N_6232,N_2331,N_2045);
or U6233 (N_6233,N_2889,N_288);
nor U6234 (N_6234,N_873,N_1392);
xnor U6235 (N_6235,N_1244,N_970);
nand U6236 (N_6236,N_4744,N_968);
nor U6237 (N_6237,N_835,N_2311);
nand U6238 (N_6238,N_3584,N_2435);
nand U6239 (N_6239,N_2602,N_1418);
xor U6240 (N_6240,N_3744,N_2173);
nor U6241 (N_6241,N_1621,N_1530);
and U6242 (N_6242,N_3384,N_363);
or U6243 (N_6243,N_3457,N_1144);
or U6244 (N_6244,N_2801,N_3972);
and U6245 (N_6245,N_1989,N_1367);
nand U6246 (N_6246,N_513,N_4120);
or U6247 (N_6247,N_2504,N_3072);
nor U6248 (N_6248,N_269,N_3011);
and U6249 (N_6249,N_475,N_3602);
nand U6250 (N_6250,N_1225,N_632);
and U6251 (N_6251,N_1455,N_1098);
nor U6252 (N_6252,N_4329,N_2962);
nand U6253 (N_6253,N_855,N_3478);
nor U6254 (N_6254,N_3307,N_4781);
or U6255 (N_6255,N_3849,N_1933);
or U6256 (N_6256,N_1714,N_4139);
or U6257 (N_6257,N_666,N_4132);
nor U6258 (N_6258,N_4878,N_53);
or U6259 (N_6259,N_882,N_964);
and U6260 (N_6260,N_1796,N_253);
xnor U6261 (N_6261,N_1260,N_3561);
nor U6262 (N_6262,N_3386,N_4265);
xor U6263 (N_6263,N_698,N_4289);
nor U6264 (N_6264,N_2079,N_2420);
nand U6265 (N_6265,N_551,N_877);
nand U6266 (N_6266,N_3937,N_1564);
xor U6267 (N_6267,N_300,N_2904);
xor U6268 (N_6268,N_2324,N_2074);
nand U6269 (N_6269,N_1407,N_4836);
nor U6270 (N_6270,N_3303,N_528);
nor U6271 (N_6271,N_282,N_1762);
and U6272 (N_6272,N_1478,N_3010);
and U6273 (N_6273,N_3053,N_3928);
xor U6274 (N_6274,N_4595,N_973);
xnor U6275 (N_6275,N_3414,N_531);
nor U6276 (N_6276,N_4050,N_3168);
xor U6277 (N_6277,N_3984,N_4105);
and U6278 (N_6278,N_4207,N_1068);
or U6279 (N_6279,N_1266,N_116);
and U6280 (N_6280,N_4953,N_1109);
or U6281 (N_6281,N_506,N_2042);
or U6282 (N_6282,N_1084,N_702);
or U6283 (N_6283,N_1529,N_2356);
or U6284 (N_6284,N_867,N_2099);
and U6285 (N_6285,N_4405,N_1972);
and U6286 (N_6286,N_1845,N_418);
nand U6287 (N_6287,N_322,N_4469);
nand U6288 (N_6288,N_3670,N_3876);
nand U6289 (N_6289,N_4829,N_3469);
or U6290 (N_6290,N_4259,N_3559);
or U6291 (N_6291,N_4225,N_3706);
nand U6292 (N_6292,N_1000,N_4384);
xnor U6293 (N_6293,N_1238,N_1784);
xor U6294 (N_6294,N_3445,N_3917);
or U6295 (N_6295,N_1029,N_2648);
nor U6296 (N_6296,N_872,N_4712);
xnor U6297 (N_6297,N_965,N_4975);
xor U6298 (N_6298,N_4731,N_4538);
nand U6299 (N_6299,N_4381,N_700);
nor U6300 (N_6300,N_1662,N_3492);
nor U6301 (N_6301,N_2286,N_4871);
nor U6302 (N_6302,N_3890,N_1389);
and U6303 (N_6303,N_4610,N_2639);
xor U6304 (N_6304,N_1718,N_307);
xnor U6305 (N_6305,N_4753,N_4349);
xor U6306 (N_6306,N_648,N_102);
or U6307 (N_6307,N_4169,N_3265);
nor U6308 (N_6308,N_4772,N_3660);
nor U6309 (N_6309,N_3182,N_4017);
nor U6310 (N_6310,N_481,N_302);
xor U6311 (N_6311,N_2411,N_4954);
xor U6312 (N_6312,N_211,N_29);
or U6313 (N_6313,N_4770,N_1705);
or U6314 (N_6314,N_316,N_4277);
and U6315 (N_6315,N_4920,N_1734);
and U6316 (N_6316,N_1985,N_1927);
nor U6317 (N_6317,N_367,N_2452);
nand U6318 (N_6318,N_4939,N_2185);
nand U6319 (N_6319,N_1848,N_723);
and U6320 (N_6320,N_483,N_553);
and U6321 (N_6321,N_1650,N_892);
xnor U6322 (N_6322,N_23,N_2092);
nor U6323 (N_6323,N_1573,N_3666);
nor U6324 (N_6324,N_454,N_2797);
and U6325 (N_6325,N_130,N_68);
nand U6326 (N_6326,N_2459,N_3043);
nand U6327 (N_6327,N_344,N_931);
and U6328 (N_6328,N_457,N_4928);
and U6329 (N_6329,N_4898,N_4685);
xnor U6330 (N_6330,N_4601,N_784);
or U6331 (N_6331,N_3075,N_2495);
and U6332 (N_6332,N_4416,N_1290);
nor U6333 (N_6333,N_1978,N_2341);
and U6334 (N_6334,N_2530,N_3372);
or U6335 (N_6335,N_1959,N_1002);
or U6336 (N_6336,N_159,N_1556);
nand U6337 (N_6337,N_883,N_1517);
xor U6338 (N_6338,N_3132,N_2336);
and U6339 (N_6339,N_3299,N_4373);
nand U6340 (N_6340,N_1870,N_3248);
and U6341 (N_6341,N_3864,N_2462);
nor U6342 (N_6342,N_2561,N_4969);
or U6343 (N_6343,N_2891,N_1957);
nand U6344 (N_6344,N_1664,N_3741);
and U6345 (N_6345,N_1690,N_1829);
nand U6346 (N_6346,N_861,N_2567);
and U6347 (N_6347,N_381,N_2204);
or U6348 (N_6348,N_1076,N_221);
nand U6349 (N_6349,N_4200,N_593);
nand U6350 (N_6350,N_2445,N_4738);
nor U6351 (N_6351,N_788,N_1001);
or U6352 (N_6352,N_529,N_3859);
nor U6353 (N_6353,N_2179,N_2657);
nand U6354 (N_6354,N_3509,N_3791);
or U6355 (N_6355,N_4599,N_166);
nor U6356 (N_6356,N_4597,N_3862);
or U6357 (N_6357,N_4912,N_1471);
nor U6358 (N_6358,N_1867,N_4202);
nand U6359 (N_6359,N_1019,N_822);
or U6360 (N_6360,N_337,N_2106);
nand U6361 (N_6361,N_2309,N_4562);
or U6362 (N_6362,N_4261,N_3887);
xnor U6363 (N_6363,N_2919,N_3115);
nand U6364 (N_6364,N_1921,N_3900);
and U6365 (N_6365,N_1422,N_913);
nor U6366 (N_6366,N_3538,N_1583);
nand U6367 (N_6367,N_3586,N_2740);
xor U6368 (N_6368,N_3198,N_2782);
nor U6369 (N_6369,N_836,N_3196);
and U6370 (N_6370,N_2213,N_3978);
xnor U6371 (N_6371,N_1437,N_4129);
or U6372 (N_6372,N_54,N_3234);
nand U6373 (N_6373,N_3192,N_4741);
xnor U6374 (N_6374,N_2783,N_669);
nand U6375 (N_6375,N_2781,N_844);
nand U6376 (N_6376,N_4541,N_614);
nor U6377 (N_6377,N_4252,N_1174);
or U6378 (N_6378,N_3047,N_4976);
or U6379 (N_6379,N_2981,N_2945);
xor U6380 (N_6380,N_2362,N_1503);
nor U6381 (N_6381,N_2078,N_3279);
and U6382 (N_6382,N_1954,N_258);
xnor U6383 (N_6383,N_3851,N_2019);
nand U6384 (N_6384,N_487,N_3850);
or U6385 (N_6385,N_2573,N_2288);
or U6386 (N_6386,N_1020,N_586);
nand U6387 (N_6387,N_1268,N_71);
nand U6388 (N_6388,N_4651,N_129);
and U6389 (N_6389,N_996,N_4866);
or U6390 (N_6390,N_3631,N_351);
or U6391 (N_6391,N_4488,N_156);
nand U6392 (N_6392,N_2509,N_3648);
or U6393 (N_6393,N_2195,N_3679);
xor U6394 (N_6394,N_2162,N_1429);
xor U6395 (N_6395,N_517,N_3374);
nor U6396 (N_6396,N_510,N_2661);
nor U6397 (N_6397,N_311,N_2157);
nand U6398 (N_6398,N_7,N_4570);
and U6399 (N_6399,N_2481,N_778);
xor U6400 (N_6400,N_3500,N_3350);
and U6401 (N_6401,N_4923,N_4297);
nor U6402 (N_6402,N_3363,N_2610);
and U6403 (N_6403,N_1397,N_3048);
or U6404 (N_6404,N_4869,N_512);
and U6405 (N_6405,N_4884,N_4892);
and U6406 (N_6406,N_1306,N_1356);
xnor U6407 (N_6407,N_1444,N_4055);
or U6408 (N_6408,N_4034,N_1527);
and U6409 (N_6409,N_4251,N_4917);
nand U6410 (N_6410,N_526,N_2724);
xnor U6411 (N_6411,N_4011,N_261);
or U6412 (N_6412,N_660,N_1127);
nor U6413 (N_6413,N_1242,N_2692);
and U6414 (N_6414,N_2293,N_4360);
xnor U6415 (N_6415,N_370,N_4616);
xnor U6416 (N_6416,N_391,N_3614);
or U6417 (N_6417,N_4480,N_4838);
nand U6418 (N_6418,N_4996,N_2282);
or U6419 (N_6419,N_2938,N_533);
nor U6420 (N_6420,N_48,N_4353);
xnor U6421 (N_6421,N_230,N_461);
nor U6422 (N_6422,N_4242,N_4115);
nor U6423 (N_6423,N_348,N_2972);
or U6424 (N_6424,N_3501,N_3283);
nor U6425 (N_6425,N_3747,N_3390);
nor U6426 (N_6426,N_2077,N_4417);
and U6427 (N_6427,N_1384,N_3525);
xor U6428 (N_6428,N_2032,N_4007);
and U6429 (N_6429,N_2163,N_3868);
xor U6430 (N_6430,N_1258,N_1820);
or U6431 (N_6431,N_3635,N_621);
or U6432 (N_6432,N_2591,N_331);
xor U6433 (N_6433,N_4401,N_1547);
nand U6434 (N_6434,N_1677,N_163);
nor U6435 (N_6435,N_285,N_1988);
nor U6436 (N_6436,N_759,N_2836);
or U6437 (N_6437,N_3068,N_2653);
or U6438 (N_6438,N_750,N_2314);
nand U6439 (N_6439,N_4749,N_1808);
or U6440 (N_6440,N_3024,N_3136);
and U6441 (N_6441,N_676,N_2524);
or U6442 (N_6442,N_2502,N_67);
or U6443 (N_6443,N_369,N_2449);
nand U6444 (N_6444,N_2193,N_4715);
nor U6445 (N_6445,N_839,N_515);
nor U6446 (N_6446,N_4848,N_2320);
nand U6447 (N_6447,N_3355,N_3748);
xnor U6448 (N_6448,N_3921,N_374);
or U6449 (N_6449,N_1562,N_2710);
xnor U6450 (N_6450,N_746,N_2780);
xnor U6451 (N_6451,N_3595,N_2181);
and U6452 (N_6452,N_3329,N_3565);
and U6453 (N_6453,N_2559,N_2800);
xnor U6454 (N_6454,N_1949,N_2009);
and U6455 (N_6455,N_1044,N_3649);
or U6456 (N_6456,N_3866,N_297);
or U6457 (N_6457,N_1857,N_3251);
nand U6458 (N_6458,N_2809,N_929);
nor U6459 (N_6459,N_783,N_1093);
nand U6460 (N_6460,N_4436,N_706);
or U6461 (N_6461,N_1177,N_2503);
nor U6462 (N_6462,N_3873,N_601);
nor U6463 (N_6463,N_3990,N_3389);
or U6464 (N_6464,N_2875,N_2924);
xnor U6465 (N_6465,N_4071,N_2120);
or U6466 (N_6466,N_3343,N_2665);
and U6467 (N_6467,N_2469,N_1777);
and U6468 (N_6468,N_2976,N_30);
xor U6469 (N_6469,N_2010,N_208);
nand U6470 (N_6470,N_4634,N_1301);
and U6471 (N_6471,N_4978,N_4627);
nand U6472 (N_6472,N_3433,N_2786);
and U6473 (N_6473,N_4439,N_1518);
and U6474 (N_6474,N_2342,N_2950);
nor U6475 (N_6475,N_729,N_4339);
nand U6476 (N_6476,N_3743,N_3087);
or U6477 (N_6477,N_3319,N_900);
and U6478 (N_6478,N_3285,N_523);
nor U6479 (N_6479,N_476,N_1508);
xnor U6480 (N_6480,N_2730,N_939);
xor U6481 (N_6481,N_1901,N_946);
or U6482 (N_6482,N_482,N_3338);
xnor U6483 (N_6483,N_3454,N_519);
and U6484 (N_6484,N_1041,N_1887);
and U6485 (N_6485,N_3216,N_3691);
and U6486 (N_6486,N_4824,N_4476);
nor U6487 (N_6487,N_2814,N_2206);
xnor U6488 (N_6488,N_4809,N_643);
xnor U6489 (N_6489,N_4901,N_2978);
nand U6490 (N_6490,N_352,N_2693);
or U6491 (N_6491,N_433,N_2490);
or U6492 (N_6492,N_191,N_3832);
nor U6493 (N_6493,N_2929,N_2557);
xor U6494 (N_6494,N_1995,N_2526);
or U6495 (N_6495,N_1015,N_2881);
nand U6496 (N_6496,N_4088,N_3755);
nand U6497 (N_6497,N_2357,N_4519);
xor U6498 (N_6498,N_4804,N_2219);
and U6499 (N_6499,N_1787,N_4249);
xnor U6500 (N_6500,N_2834,N_165);
nand U6501 (N_6501,N_2865,N_2775);
or U6502 (N_6502,N_1416,N_2028);
nand U6503 (N_6503,N_440,N_4035);
nor U6504 (N_6504,N_4023,N_2268);
xnor U6505 (N_6505,N_657,N_3844);
or U6506 (N_6506,N_4364,N_2468);
xnor U6507 (N_6507,N_1442,N_1249);
and U6508 (N_6508,N_4430,N_1417);
and U6509 (N_6509,N_2498,N_2327);
nand U6510 (N_6510,N_1577,N_455);
nor U6511 (N_6511,N_2210,N_2630);
or U6512 (N_6512,N_4907,N_3605);
xnor U6513 (N_6513,N_104,N_1150);
nand U6514 (N_6514,N_3805,N_1785);
xor U6515 (N_6515,N_2271,N_2646);
xor U6516 (N_6516,N_671,N_1833);
xnor U6517 (N_6517,N_3510,N_682);
nand U6518 (N_6518,N_2345,N_3842);
or U6519 (N_6519,N_959,N_180);
nor U6520 (N_6520,N_4429,N_217);
and U6521 (N_6521,N_1937,N_2470);
nand U6522 (N_6522,N_2020,N_4552);
nand U6523 (N_6523,N_722,N_4794);
or U6524 (N_6524,N_4213,N_41);
nor U6525 (N_6525,N_3171,N_576);
and U6526 (N_6526,N_2770,N_2547);
nor U6527 (N_6527,N_3404,N_1047);
xor U6528 (N_6528,N_105,N_2344);
nor U6529 (N_6529,N_1333,N_3431);
and U6530 (N_6530,N_4941,N_4940);
nor U6531 (N_6531,N_1142,N_647);
nand U6532 (N_6532,N_2806,N_4880);
xor U6533 (N_6533,N_4155,N_2913);
and U6534 (N_6534,N_4340,N_4702);
xnor U6535 (N_6535,N_243,N_2666);
nand U6536 (N_6536,N_782,N_4415);
nand U6537 (N_6537,N_91,N_3830);
nand U6538 (N_6538,N_2707,N_1311);
nor U6539 (N_6539,N_4273,N_299);
or U6540 (N_6540,N_1837,N_144);
xnor U6541 (N_6541,N_2263,N_1026);
or U6542 (N_6542,N_4496,N_207);
or U6543 (N_6543,N_3999,N_4181);
and U6544 (N_6544,N_2228,N_2068);
nand U6545 (N_6545,N_4921,N_2407);
and U6546 (N_6546,N_3323,N_3256);
or U6547 (N_6547,N_1519,N_842);
and U6548 (N_6548,N_4111,N_760);
or U6549 (N_6549,N_4805,N_2047);
nor U6550 (N_6550,N_4663,N_2376);
and U6551 (N_6551,N_4412,N_2102);
or U6552 (N_6552,N_2124,N_2171);
nor U6553 (N_6553,N_189,N_2852);
nor U6554 (N_6554,N_1293,N_2222);
nand U6555 (N_6555,N_2060,N_4032);
nand U6556 (N_6556,N_753,N_4948);
and U6557 (N_6557,N_3489,N_3207);
nand U6558 (N_6558,N_4983,N_544);
or U6559 (N_6559,N_4667,N_1347);
or U6560 (N_6560,N_1594,N_2574);
and U6561 (N_6561,N_1075,N_110);
xnor U6562 (N_6562,N_3335,N_4448);
or U6563 (N_6563,N_1284,N_3365);
and U6564 (N_6564,N_1308,N_3166);
or U6565 (N_6565,N_2546,N_2257);
and U6566 (N_6566,N_4832,N_4127);
and U6567 (N_6567,N_1035,N_1535);
nor U6568 (N_6568,N_1393,N_404);
and U6569 (N_6569,N_4933,N_1021);
nor U6570 (N_6570,N_3117,N_3250);
nor U6571 (N_6571,N_659,N_4934);
nand U6572 (N_6572,N_3511,N_2523);
nor U6573 (N_6573,N_4985,N_2052);
nor U6574 (N_6574,N_1913,N_3029);
and U6575 (N_6575,N_2119,N_3923);
nand U6576 (N_6576,N_3438,N_3983);
and U6577 (N_6577,N_1024,N_3282);
nand U6578 (N_6578,N_2062,N_1780);
nor U6579 (N_6579,N_4243,N_2774);
nor U6580 (N_6580,N_2428,N_1973);
and U6581 (N_6581,N_3131,N_2510);
nor U6582 (N_6582,N_32,N_2129);
nor U6583 (N_6583,N_2234,N_2920);
and U6584 (N_6584,N_3888,N_4747);
nand U6585 (N_6585,N_1830,N_536);
xnor U6586 (N_6586,N_2970,N_4637);
xor U6587 (N_6587,N_3723,N_3993);
nor U6588 (N_6588,N_2033,N_1469);
nor U6589 (N_6589,N_2476,N_2822);
and U6590 (N_6590,N_3853,N_3985);
xnor U6591 (N_6591,N_705,N_1635);
and U6592 (N_6592,N_4568,N_2221);
or U6593 (N_6593,N_3906,N_1149);
xor U6594 (N_6594,N_1505,N_2762);
and U6595 (N_6595,N_3809,N_3893);
and U6596 (N_6596,N_1074,N_3667);
nor U6597 (N_6597,N_2572,N_4526);
or U6598 (N_6598,N_3979,N_210);
xnor U6599 (N_6599,N_2717,N_1134);
or U6600 (N_6600,N_4647,N_3139);
nand U6601 (N_6601,N_3829,N_1220);
nand U6602 (N_6602,N_2864,N_969);
nand U6603 (N_6603,N_415,N_3858);
nor U6604 (N_6604,N_1496,N_2479);
nand U6605 (N_6605,N_762,N_4324);
or U6606 (N_6606,N_3947,N_2335);
or U6607 (N_6607,N_2807,N_1168);
nand U6608 (N_6608,N_3111,N_2744);
and U6609 (N_6609,N_3946,N_3266);
nor U6610 (N_6610,N_715,N_3933);
nor U6611 (N_6611,N_4830,N_3435);
or U6612 (N_6612,N_3627,N_4077);
or U6613 (N_6613,N_1187,N_3092);
xor U6614 (N_6614,N_3521,N_3272);
nor U6615 (N_6615,N_4477,N_3773);
or U6616 (N_6616,N_2905,N_1846);
and U6617 (N_6617,N_3281,N_3965);
xnor U6618 (N_6618,N_350,N_3716);
nor U6619 (N_6619,N_3054,N_1136);
and U6620 (N_6620,N_2576,N_558);
nor U6621 (N_6621,N_4418,N_673);
nor U6622 (N_6622,N_4345,N_188);
xor U6623 (N_6623,N_1412,N_1467);
or U6624 (N_6624,N_1672,N_2161);
nand U6625 (N_6625,N_3057,N_3779);
nor U6626 (N_6626,N_2353,N_1181);
or U6627 (N_6627,N_2388,N_3467);
and U6628 (N_6628,N_2846,N_975);
xor U6629 (N_6629,N_4051,N_3019);
and U6630 (N_6630,N_468,N_4428);
or U6631 (N_6631,N_2687,N_3218);
xnor U6632 (N_6632,N_3529,N_3514);
and U6633 (N_6633,N_3975,N_4219);
xnor U6634 (N_6634,N_1330,N_2326);
or U6635 (N_6635,N_2034,N_4379);
nand U6636 (N_6636,N_1423,N_3669);
xor U6637 (N_6637,N_93,N_1342);
nand U6638 (N_6638,N_4170,N_1641);
and U6639 (N_6639,N_4237,N_1125);
nand U6640 (N_6640,N_4370,N_2237);
nor U6641 (N_6641,N_2721,N_4186);
nor U6642 (N_6642,N_4165,N_421);
nand U6643 (N_6643,N_4328,N_1720);
and U6644 (N_6644,N_4054,N_4563);
nor U6645 (N_6645,N_3296,N_1912);
and U6646 (N_6646,N_4661,N_3811);
nor U6647 (N_6647,N_3138,N_4138);
nand U6648 (N_6648,N_2890,N_2999);
or U6649 (N_6649,N_4322,N_2532);
nand U6650 (N_6650,N_1501,N_1167);
or U6651 (N_6651,N_4984,N_1791);
nor U6652 (N_6652,N_4183,N_2319);
nor U6653 (N_6653,N_4369,N_3448);
xor U6654 (N_6654,N_3623,N_864);
or U6655 (N_6655,N_2154,N_1361);
or U6656 (N_6656,N_1298,N_2623);
nand U6657 (N_6657,N_2265,N_3986);
and U6658 (N_6658,N_2,N_2993);
nand U6659 (N_6659,N_1287,N_387);
and U6660 (N_6660,N_3970,N_514);
or U6661 (N_6661,N_4004,N_4596);
or U6662 (N_6662,N_3599,N_1916);
nor U6663 (N_6663,N_2618,N_3714);
nand U6664 (N_6664,N_197,N_1235);
nor U6665 (N_6665,N_1470,N_1102);
or U6666 (N_6666,N_1435,N_2575);
nand U6667 (N_6667,N_966,N_4825);
or U6668 (N_6668,N_290,N_1299);
or U6669 (N_6669,N_452,N_1682);
nor U6670 (N_6670,N_3680,N_2160);
nand U6671 (N_6671,N_2855,N_4109);
nand U6672 (N_6672,N_1161,N_1865);
nor U6673 (N_6673,N_3697,N_3463);
xnor U6674 (N_6674,N_3163,N_3257);
nand U6675 (N_6675,N_139,N_4203);
and U6676 (N_6676,N_2940,N_2645);
and U6677 (N_6677,N_451,N_427);
and U6678 (N_6678,N_1743,N_522);
or U6679 (N_6679,N_1778,N_3362);
xnor U6680 (N_6680,N_3446,N_3297);
xor U6681 (N_6681,N_4668,N_3657);
or U6682 (N_6682,N_4301,N_136);
xor U6683 (N_6683,N_3108,N_24);
nand U6684 (N_6684,N_4530,N_3709);
nor U6685 (N_6685,N_789,N_1413);
xor U6686 (N_6686,N_3569,N_612);
nand U6687 (N_6687,N_2083,N_4768);
or U6688 (N_6688,N_181,N_4284);
and U6689 (N_6689,N_2808,N_2732);
nor U6690 (N_6690,N_4960,N_2901);
nand U6691 (N_6691,N_818,N_539);
and U6692 (N_6692,N_1457,N_699);
nand U6693 (N_6693,N_1610,N_2514);
or U6694 (N_6694,N_1862,N_4466);
xnor U6695 (N_6695,N_1798,N_3908);
and U6696 (N_6696,N_1408,N_4241);
and U6697 (N_6697,N_1378,N_3407);
and U6698 (N_6698,N_4315,N_3274);
nor U6699 (N_6699,N_2454,N_2823);
nand U6700 (N_6700,N_142,N_769);
or U6701 (N_6701,N_3437,N_1548);
nand U6702 (N_6702,N_4276,N_4946);
and U6703 (N_6703,N_2676,N_3916);
nor U6704 (N_6704,N_909,N_4608);
xnor U6705 (N_6705,N_4618,N_4172);
nor U6706 (N_6706,N_2593,N_113);
nand U6707 (N_6707,N_801,N_4937);
nor U6708 (N_6708,N_1636,N_4454);
xnor U6709 (N_6709,N_4554,N_3109);
xor U6710 (N_6710,N_4435,N_3348);
xnor U6711 (N_6711,N_291,N_4067);
or U6712 (N_6712,N_1461,N_1609);
nor U6713 (N_6713,N_4052,N_101);
or U6714 (N_6714,N_2628,N_1678);
nand U6715 (N_6715,N_4544,N_2027);
xnor U6716 (N_6716,N_566,N_324);
nor U6717 (N_6717,N_2624,N_908);
xnor U6718 (N_6718,N_1793,N_923);
and U6719 (N_6719,N_2696,N_4870);
or U6720 (N_6720,N_1923,N_607);
xor U6721 (N_6721,N_678,N_2370);
xnor U6722 (N_6722,N_375,N_1323);
nor U6723 (N_6723,N_4238,N_1764);
or U6724 (N_6724,N_3855,N_1296);
and U6725 (N_6725,N_1651,N_2277);
nand U6726 (N_6726,N_1251,N_3871);
nand U6727 (N_6727,N_1217,N_424);
or U6728 (N_6728,N_317,N_2850);
or U6729 (N_6729,N_1864,N_3369);
and U6730 (N_6730,N_2513,N_2637);
and U6731 (N_6731,N_471,N_2900);
nand U6732 (N_6732,N_2614,N_2377);
nand U6733 (N_6733,N_4879,N_4915);
or U6734 (N_6734,N_3998,N_2281);
and U6735 (N_6735,N_4468,N_708);
nand U6736 (N_6736,N_3814,N_2294);
nand U6737 (N_6737,N_2632,N_2379);
nor U6738 (N_6738,N_4291,N_2691);
and U6739 (N_6739,N_1731,N_2207);
xor U6740 (N_6740,N_4807,N_365);
nand U6741 (N_6741,N_1373,N_1355);
and U6742 (N_6742,N_1770,N_3370);
or U6743 (N_6743,N_772,N_4837);
and U6744 (N_6744,N_49,N_1337);
nor U6745 (N_6745,N_2395,N_2845);
xnor U6746 (N_6746,N_2081,N_4465);
nor U6747 (N_6747,N_4472,N_2169);
xor U6748 (N_6748,N_646,N_9);
or U6749 (N_6749,N_3400,N_3731);
or U6750 (N_6750,N_2622,N_1477);
and U6751 (N_6751,N_4859,N_870);
nand U6752 (N_6752,N_3530,N_3760);
or U6753 (N_6753,N_3103,N_254);
and U6754 (N_6754,N_623,N_791);
or U6755 (N_6755,N_4936,N_3458);
and U6756 (N_6756,N_2741,N_1345);
and U6757 (N_6757,N_2049,N_268);
nor U6758 (N_6758,N_1982,N_3051);
xor U6759 (N_6759,N_2404,N_1521);
nor U6760 (N_6760,N_443,N_3581);
xor U6761 (N_6761,N_819,N_3550);
nand U6762 (N_6762,N_2802,N_3537);
or U6763 (N_6763,N_382,N_2385);
and U6764 (N_6764,N_259,N_4383);
nand U6765 (N_6765,N_2296,N_1274);
or U6766 (N_6766,N_439,N_4861);
xnor U6767 (N_6767,N_1364,N_4362);
nor U6768 (N_6768,N_2297,N_3910);
xnor U6769 (N_6769,N_2457,N_2018);
xor U6770 (N_6770,N_1710,N_4585);
or U6771 (N_6771,N_2058,N_281);
and U6772 (N_6772,N_1877,N_94);
and U6773 (N_6773,N_3952,N_3782);
nor U6774 (N_6774,N_2007,N_106);
and U6775 (N_6775,N_3824,N_3376);
and U6776 (N_6776,N_3882,N_3419);
xnor U6777 (N_6777,N_4166,N_2790);
and U6778 (N_6778,N_3499,N_611);
and U6779 (N_6779,N_4800,N_3450);
nor U6780 (N_6780,N_2679,N_3542);
nor U6781 (N_6781,N_2720,N_2488);
nor U6782 (N_6782,N_2241,N_3357);
or U6783 (N_6783,N_4374,N_3846);
nand U6784 (N_6784,N_2046,N_407);
and U6785 (N_6785,N_2348,N_4310);
and U6786 (N_6786,N_2430,N_2322);
nor U6787 (N_6787,N_1062,N_3461);
and U6788 (N_6788,N_4578,N_4239);
and U6789 (N_6789,N_4475,N_667);
nor U6790 (N_6790,N_4823,N_3254);
nor U6791 (N_6791,N_1126,N_1227);
xor U6792 (N_6792,N_1512,N_1655);
xnor U6793 (N_6793,N_1464,N_2230);
or U6794 (N_6794,N_3927,N_4757);
nor U6795 (N_6795,N_1881,N_4318);
and U6796 (N_6796,N_1292,N_263);
and U6797 (N_6797,N_1802,N_4965);
xor U6798 (N_6798,N_1948,N_1810);
and U6799 (N_6799,N_14,N_858);
nor U6800 (N_6800,N_4247,N_4735);
nor U6801 (N_6801,N_2803,N_4528);
and U6802 (N_6802,N_4411,N_1239);
xnor U6803 (N_6803,N_4108,N_1756);
nand U6804 (N_6804,N_3003,N_1117);
xor U6805 (N_6805,N_3101,N_1207);
or U6806 (N_6806,N_12,N_2986);
or U6807 (N_6807,N_3767,N_3049);
nand U6808 (N_6808,N_111,N_4459);
nand U6809 (N_6809,N_1592,N_2778);
nand U6810 (N_6810,N_3371,N_1868);
xnor U6811 (N_6811,N_4198,N_326);
nand U6812 (N_6812,N_4536,N_3810);
nand U6813 (N_6813,N_174,N_4664);
and U6814 (N_6814,N_2339,N_2545);
nand U6815 (N_6815,N_2158,N_4375);
xor U6816 (N_6816,N_2598,N_962);
nand U6817 (N_6817,N_2041,N_1094);
or U6818 (N_6818,N_2833,N_154);
nand U6819 (N_6819,N_2321,N_1965);
nand U6820 (N_6820,N_4253,N_4209);
or U6821 (N_6821,N_3378,N_2091);
nand U6822 (N_6822,N_4756,N_18);
xor U6823 (N_6823,N_2401,N_4909);
or U6824 (N_6824,N_2144,N_3252);
nor U6825 (N_6825,N_1061,N_1097);
nand U6826 (N_6826,N_3312,N_4409);
or U6827 (N_6827,N_2427,N_3957);
xor U6828 (N_6828,N_4033,N_2664);
xnor U6829 (N_6829,N_3017,N_3554);
and U6830 (N_6830,N_1821,N_1850);
and U6831 (N_6831,N_3637,N_204);
nand U6832 (N_6832,N_4515,N_712);
and U6833 (N_6833,N_138,N_2876);
xnor U6834 (N_6834,N_2072,N_1269);
or U6835 (N_6835,N_1132,N_1907);
nand U6836 (N_6836,N_3541,N_3612);
nand U6837 (N_6837,N_2441,N_280);
and U6838 (N_6838,N_1064,N_2654);
xor U6839 (N_6839,N_3134,N_1474);
or U6840 (N_6840,N_4688,N_3028);
nand U6841 (N_6841,N_3070,N_3608);
nand U6842 (N_6842,N_740,N_4951);
or U6843 (N_6843,N_4026,N_630);
or U6844 (N_6844,N_4523,N_1204);
nor U6845 (N_6845,N_4093,N_1409);
and U6846 (N_6846,N_1679,N_4307);
nor U6847 (N_6847,N_796,N_1561);
or U6848 (N_6848,N_2838,N_4065);
or U6849 (N_6849,N_1341,N_2997);
nor U6850 (N_6850,N_2086,N_4817);
xor U6851 (N_6851,N_1616,N_3996);
and U6852 (N_6852,N_3321,N_2287);
or U6853 (N_6853,N_1486,N_2410);
nand U6854 (N_6854,N_3737,N_4372);
and U6855 (N_6855,N_748,N_2473);
xor U6856 (N_6856,N_1130,N_3951);
or U6857 (N_6857,N_798,N_4147);
xor U6858 (N_6858,N_429,N_3536);
or U6859 (N_6859,N_2604,N_50);
xnor U6860 (N_6860,N_2723,N_1386);
and U6861 (N_6861,N_58,N_3884);
and U6862 (N_6862,N_47,N_4399);
nand U6863 (N_6863,N_2914,N_2055);
nand U6864 (N_6864,N_1586,N_4648);
and U6865 (N_6865,N_3066,N_1374);
or U6866 (N_6866,N_3935,N_2506);
nor U6867 (N_6867,N_2579,N_1603);
nor U6868 (N_6868,N_1432,N_1844);
nor U6869 (N_6869,N_2201,N_2148);
and U6870 (N_6870,N_61,N_1485);
xnor U6871 (N_6871,N_3006,N_2292);
or U6872 (N_6872,N_149,N_1231);
nand U6873 (N_6873,N_3632,N_233);
xnor U6874 (N_6874,N_2436,N_3258);
nor U6875 (N_6875,N_1809,N_4846);
nor U6876 (N_6876,N_3621,N_146);
nand U6877 (N_6877,N_1077,N_3886);
nand U6878 (N_6878,N_1805,N_1119);
and U6879 (N_6879,N_100,N_1628);
or U6880 (N_6880,N_2650,N_4094);
nor U6881 (N_6881,N_3642,N_1159);
nor U6882 (N_6882,N_4577,N_1590);
and U6883 (N_6883,N_2512,N_152);
and U6884 (N_6884,N_4784,N_2109);
xnor U6885 (N_6885,N_450,N_4621);
and U6886 (N_6886,N_4614,N_1782);
or U6887 (N_6887,N_1991,N_4956);
xnor U6888 (N_6888,N_120,N_1717);
nor U6889 (N_6889,N_3733,N_1484);
nand U6890 (N_6890,N_2668,N_2259);
nor U6891 (N_6891,N_2987,N_3929);
xor U6892 (N_6892,N_1797,N_2116);
or U6893 (N_6893,N_469,N_4189);
nor U6894 (N_6894,N_1998,N_2620);
and U6895 (N_6895,N_843,N_3784);
xnor U6896 (N_6896,N_4691,N_1491);
nor U6897 (N_6897,N_4163,N_3291);
or U6898 (N_6898,N_1924,N_2013);
or U6899 (N_6899,N_1572,N_1849);
nor U6900 (N_6900,N_474,N_1999);
nor U6901 (N_6901,N_2505,N_2346);
nand U6902 (N_6902,N_3728,N_1459);
nand U6903 (N_6903,N_1932,N_1888);
nor U6904 (N_6904,N_2051,N_1993);
xnor U6905 (N_6905,N_386,N_4080);
and U6906 (N_6906,N_289,N_1691);
xnor U6907 (N_6907,N_4431,N_738);
nor U6908 (N_6908,N_1819,N_1759);
xor U6909 (N_6909,N_2609,N_3531);
or U6910 (N_6910,N_2761,N_2390);
nand U6911 (N_6911,N_3286,N_3406);
nand U6912 (N_6912,N_2617,N_1443);
and U6913 (N_6913,N_2300,N_2944);
nor U6914 (N_6914,N_3968,N_1166);
nand U6915 (N_6915,N_3961,N_525);
nor U6916 (N_6916,N_4503,N_1963);
or U6917 (N_6917,N_954,N_1046);
xnor U6918 (N_6918,N_927,N_2165);
nor U6919 (N_6919,N_3225,N_252);
xnor U6920 (N_6920,N_2906,N_4593);
nor U6921 (N_6921,N_1036,N_184);
nor U6922 (N_6922,N_633,N_313);
xnor U6923 (N_6923,N_3475,N_4098);
and U6924 (N_6924,N_3124,N_956);
and U6925 (N_6925,N_56,N_4874);
or U6926 (N_6926,N_3902,N_2191);
or U6927 (N_6927,N_3772,N_1622);
nand U6928 (N_6928,N_4639,N_4635);
xnor U6929 (N_6929,N_3903,N_4963);
nand U6930 (N_6930,N_1611,N_1261);
or U6931 (N_6931,N_1546,N_4149);
or U6932 (N_6932,N_4185,N_2008);
nand U6933 (N_6933,N_672,N_3555);
or U6934 (N_6934,N_2673,N_1657);
or U6935 (N_6935,N_1794,N_2218);
and U6936 (N_6936,N_3681,N_1553);
and U6937 (N_6937,N_4426,N_3651);
nor U6938 (N_6938,N_546,N_1685);
nand U6939 (N_6939,N_4582,N_2935);
xor U6940 (N_6940,N_924,N_2768);
and U6941 (N_6941,N_3008,N_4716);
nor U6942 (N_6942,N_4022,N_1550);
nor U6943 (N_6943,N_2917,N_4210);
xnor U6944 (N_6944,N_3324,N_4245);
or U6945 (N_6945,N_3079,N_4334);
and U6946 (N_6946,N_4313,N_994);
xor U6947 (N_6947,N_3315,N_2727);
or U6948 (N_6948,N_4520,N_2141);
or U6949 (N_6949,N_4573,N_1807);
nor U6950 (N_6950,N_4222,N_1674);
or U6951 (N_6951,N_3276,N_2798);
or U6952 (N_6952,N_1003,N_2483);
nor U6953 (N_6953,N_3429,N_3977);
and U6954 (N_6954,N_3835,N_3165);
or U6955 (N_6955,N_1723,N_3268);
and U6956 (N_6956,N_4060,N_957);
nor U6957 (N_6957,N_1349,N_4008);
xor U6958 (N_6958,N_1493,N_4797);
xor U6959 (N_6959,N_157,N_4628);
xor U6960 (N_6960,N_1321,N_2238);
or U6961 (N_6961,N_733,N_3292);
and U6962 (N_6962,N_143,N_516);
and U6963 (N_6963,N_4982,N_3924);
nand U6964 (N_6964,N_3568,N_4395);
nor U6965 (N_6965,N_2394,N_1387);
xor U6966 (N_6966,N_1816,N_3352);
nand U6967 (N_6967,N_3896,N_1073);
or U6968 (N_6968,N_2138,N_3421);
and U6969 (N_6969,N_2398,N_2433);
or U6970 (N_6970,N_4125,N_3711);
xnor U6971 (N_6971,N_492,N_4167);
nor U6972 (N_6972,N_330,N_532);
xor U6973 (N_6973,N_4260,N_502);
or U6974 (N_6974,N_3459,N_85);
nor U6975 (N_6975,N_3954,N_1944);
or U6976 (N_6976,N_2626,N_4485);
or U6977 (N_6977,N_4755,N_2634);
nand U6978 (N_6978,N_1909,N_1400);
and U6979 (N_6979,N_4136,N_4707);
nor U6980 (N_6980,N_4675,N_3894);
nor U6981 (N_6981,N_4351,N_3756);
or U6982 (N_6982,N_3981,N_3487);
and U6983 (N_6983,N_1943,N_4350);
nor U6984 (N_6984,N_1353,N_2866);
xor U6985 (N_6985,N_4076,N_410);
nand U6986 (N_6986,N_2199,N_2347);
or U6987 (N_6987,N_2625,N_2355);
or U6988 (N_6988,N_1156,N_4371);
nand U6989 (N_6989,N_4752,N_4116);
and U6990 (N_6990,N_2991,N_3417);
xor U6991 (N_6991,N_3643,N_2759);
nand U6992 (N_6992,N_1773,N_2957);
or U6993 (N_6993,N_2235,N_1143);
nor U6994 (N_6994,N_3,N_3412);
xor U6995 (N_6995,N_1968,N_1634);
xor U6996 (N_6996,N_1402,N_1915);
nor U6997 (N_6997,N_2090,N_1812);
or U6998 (N_6998,N_4787,N_193);
xor U6999 (N_6999,N_1037,N_776);
xnor U7000 (N_7000,N_2813,N_1689);
and U7001 (N_7001,N_2071,N_109);
or U7002 (N_7002,N_3179,N_1860);
nor U7003 (N_7003,N_1889,N_590);
nand U7004 (N_7004,N_716,N_1472);
nand U7005 (N_7005,N_695,N_1899);
or U7006 (N_7006,N_1210,N_2606);
or U7007 (N_7007,N_2771,N_3735);
and U7008 (N_7008,N_107,N_849);
xor U7009 (N_7009,N_1766,N_1388);
xor U7010 (N_7010,N_3878,N_1545);
or U7011 (N_7011,N_3687,N_1744);
nor U7012 (N_7012,N_2581,N_2391);
or U7013 (N_7013,N_2969,N_2130);
nand U7014 (N_7014,N_1329,N_3240);
nand U7015 (N_7015,N_1645,N_2145);
nand U7016 (N_7016,N_3624,N_4450);
nor U7017 (N_7017,N_4590,N_582);
and U7018 (N_7018,N_597,N_2854);
and U7019 (N_7019,N_2050,N_2973);
nor U7020 (N_7020,N_600,N_3174);
nand U7021 (N_7021,N_4624,N_456);
and U7022 (N_7022,N_3781,N_13);
or U7023 (N_7023,N_3220,N_4090);
and U7024 (N_7024,N_4548,N_246);
nor U7025 (N_7025,N_599,N_3490);
xnor U7026 (N_7026,N_4565,N_2264);
and U7027 (N_7027,N_1633,N_3838);
nand U7028 (N_7028,N_1536,N_3280);
and U7029 (N_7029,N_3067,N_3013);
or U7030 (N_7030,N_4346,N_3575);
nand U7031 (N_7031,N_3515,N_4762);
nand U7032 (N_7032,N_4990,N_914);
nand U7033 (N_7033,N_4894,N_214);
nand U7034 (N_7034,N_4066,N_4355);
and U7035 (N_7035,N_2239,N_1264);
nand U7036 (N_7036,N_1453,N_4280);
xnor U7037 (N_7037,N_3964,N_1466);
nor U7038 (N_7038,N_4793,N_3223);
nand U7039 (N_7039,N_473,N_4018);
nor U7040 (N_7040,N_3819,N_817);
or U7041 (N_7041,N_3361,N_4199);
and U7042 (N_7042,N_3877,N_1581);
or U7043 (N_7043,N_3099,N_1776);
or U7044 (N_7044,N_3447,N_4602);
and U7045 (N_7045,N_1314,N_3739);
or U7046 (N_7046,N_1379,N_1488);
nor U7047 (N_7047,N_1033,N_741);
and U7048 (N_7048,N_2603,N_3732);
xor U7049 (N_7049,N_1604,N_2764);
nor U7050 (N_7050,N_63,N_3113);
xor U7051 (N_7051,N_4446,N_2592);
xor U7052 (N_7052,N_3879,N_4027);
and U7053 (N_7053,N_3045,N_3991);
nor U7054 (N_7054,N_1822,N_4581);
nor U7055 (N_7055,N_1203,N_4333);
or U7056 (N_7056,N_1890,N_4736);
nor U7057 (N_7057,N_27,N_4039);
nor U7058 (N_7058,N_1335,N_3562);
or U7059 (N_7059,N_1792,N_727);
nor U7060 (N_7060,N_4061,N_3874);
and U7061 (N_7061,N_4589,N_4727);
xor U7062 (N_7062,N_569,N_2942);
or U7063 (N_7063,N_2690,N_765);
nand U7064 (N_7064,N_77,N_465);
or U7065 (N_7065,N_295,N_1523);
and U7066 (N_7066,N_4016,N_606);
and U7067 (N_7067,N_2444,N_3187);
nor U7068 (N_7068,N_1385,N_3496);
xor U7069 (N_7069,N_4278,N_432);
nor U7070 (N_7070,N_4938,N_2728);
or U7071 (N_7071,N_4440,N_2643);
and U7072 (N_7072,N_4697,N_406);
and U7073 (N_7073,N_1232,N_4230);
and U7074 (N_7074,N_1992,N_938);
nand U7075 (N_7075,N_2107,N_4684);
or U7076 (N_7076,N_3646,N_1224);
or U7077 (N_7077,N_2688,N_2939);
xnor U7078 (N_7078,N_4358,N_2899);
or U7079 (N_7079,N_568,N_2174);
and U7080 (N_7080,N_4765,N_2856);
nor U7081 (N_7081,N_4703,N_325);
and U7082 (N_7082,N_2005,N_911);
nand U7083 (N_7083,N_4081,N_1133);
xor U7084 (N_7084,N_2227,N_1665);
or U7085 (N_7085,N_1213,N_3576);
or U7086 (N_7086,N_574,N_650);
xnor U7087 (N_7087,N_1151,N_3959);
nand U7088 (N_7088,N_739,N_4217);
or U7089 (N_7089,N_2229,N_3036);
nand U7090 (N_7090,N_3167,N_4191);
or U7091 (N_7091,N_3311,N_628);
nor U7092 (N_7092,N_2631,N_2652);
nor U7093 (N_7093,N_2672,N_2364);
nor U7094 (N_7094,N_1693,N_1643);
and U7095 (N_7095,N_3190,N_4972);
xnor U7096 (N_7096,N_1280,N_1421);
nor U7097 (N_7097,N_484,N_1588);
or U7098 (N_7098,N_2393,N_2175);
nand U7099 (N_7099,N_4221,N_3615);
nand U7100 (N_7100,N_3304,N_4711);
xnor U7101 (N_7101,N_3185,N_65);
nand U7102 (N_7102,N_83,N_627);
xnor U7103 (N_7103,N_1838,N_4698);
nand U7104 (N_7104,N_1233,N_4168);
nand U7105 (N_7105,N_3742,N_1497);
xnor U7106 (N_7106,N_2551,N_1721);
xor U7107 (N_7107,N_1495,N_2403);
nor U7108 (N_7108,N_2432,N_1113);
and U7109 (N_7109,N_4709,N_2861);
and U7110 (N_7110,N_1327,N_4644);
and U7111 (N_7111,N_3863,N_1919);
nor U7112 (N_7112,N_3997,N_346);
or U7113 (N_7113,N_4336,N_2186);
xnor U7114 (N_7114,N_153,N_2375);
xor U7115 (N_7115,N_1667,N_1551);
xor U7116 (N_7116,N_73,N_4471);
nand U7117 (N_7117,N_3692,N_1163);
xnor U7118 (N_7118,N_3919,N_411);
nor U7119 (N_7119,N_1183,N_2642);
nand U7120 (N_7120,N_1011,N_4101);
and U7121 (N_7121,N_1103,N_3650);
or U7122 (N_7122,N_2197,N_1428);
xor U7123 (N_7123,N_1656,N_2675);
or U7124 (N_7124,N_987,N_3030);
xor U7125 (N_7125,N_244,N_4900);
and U7126 (N_7126,N_271,N_4862);
xor U7127 (N_7127,N_2534,N_2519);
xor U7128 (N_7128,N_2419,N_1692);
or U7129 (N_7129,N_548,N_4020);
or U7130 (N_7130,N_2930,N_4507);
nor U7131 (N_7131,N_1728,N_4813);
and U7132 (N_7132,N_1265,N_934);
or U7133 (N_7133,N_2884,N_1114);
or U7134 (N_7134,N_2493,N_1568);
nand U7135 (N_7135,N_4952,N_251);
nand U7136 (N_7136,N_4910,N_2662);
nor U7137 (N_7137,N_2029,N_2151);
and U7138 (N_7138,N_3346,N_622);
and U7139 (N_7139,N_1124,N_2704);
or U7140 (N_7140,N_3715,N_1433);
or U7141 (N_7141,N_2333,N_781);
nor U7142 (N_7142,N_123,N_426);
or U7143 (N_7143,N_3658,N_4000);
nor U7144 (N_7144,N_4856,N_4404);
and U7145 (N_7145,N_4743,N_4843);
nor U7146 (N_7146,N_2531,N_4958);
and U7147 (N_7147,N_1278,N_3275);
and U7148 (N_7148,N_2729,N_1706);
nor U7149 (N_7149,N_3379,N_3654);
and U7150 (N_7150,N_2017,N_4294);
nor U7151 (N_7151,N_891,N_1806);
nor U7152 (N_7152,N_2455,N_4966);
and U7153 (N_7153,N_1967,N_2001);
nor U7154 (N_7154,N_2236,N_4141);
nand U7155 (N_7155,N_4263,N_4043);
nand U7156 (N_7156,N_3204,N_4357);
xor U7157 (N_7157,N_3037,N_2947);
or U7158 (N_7158,N_2982,N_4993);
nor U7159 (N_7159,N_3261,N_55);
nand U7160 (N_7160,N_761,N_2587);
xnor U7161 (N_7161,N_328,N_3004);
nand U7162 (N_7162,N_3793,N_4721);
or U7163 (N_7163,N_4740,N_4764);
and U7164 (N_7164,N_3641,N_1063);
nand U7165 (N_7165,N_3294,N_1883);
xnor U7166 (N_7166,N_1697,N_256);
or U7167 (N_7167,N_1128,N_1241);
xor U7168 (N_7168,N_1200,N_3820);
nand U7169 (N_7169,N_4272,N_3725);
xor U7170 (N_7170,N_1910,N_3409);
nor U7171 (N_7171,N_1430,N_2223);
and U7172 (N_7172,N_2907,N_2414);
or U7173 (N_7173,N_477,N_4722);
and U7174 (N_7174,N_4529,N_3154);
and U7175 (N_7175,N_4545,N_2651);
nor U7176 (N_7176,N_2100,N_2685);
nor U7177 (N_7177,N_3944,N_1904);
xor U7178 (N_7178,N_3973,N_3479);
nand U7179 (N_7179,N_453,N_4449);
nand U7180 (N_7180,N_1038,N_182);
and U7181 (N_7181,N_1575,N_3267);
and U7182 (N_7182,N_4299,N_731);
or U7183 (N_7183,N_1131,N_2080);
and U7184 (N_7184,N_1945,N_2011);
nand U7185 (N_7185,N_2766,N_4492);
or U7186 (N_7186,N_2539,N_40);
nand U7187 (N_7187,N_2811,N_578);
or U7188 (N_7188,N_2909,N_176);
nor U7189 (N_7189,N_4089,N_3349);
nand U7190 (N_7190,N_1295,N_1853);
nand U7191 (N_7191,N_2396,N_3721);
and U7192 (N_7192,N_2405,N_212);
and U7193 (N_7193,N_287,N_112);
nand U7194 (N_7194,N_3881,N_1482);
xnor U7195 (N_7195,N_2114,N_2386);
nor U7196 (N_7196,N_2170,N_1528);
nor U7197 (N_7197,N_808,N_541);
nand U7198 (N_7198,N_4833,N_3843);
nor U7199 (N_7199,N_1511,N_3705);
and U7200 (N_7200,N_2755,N_3425);
nand U7201 (N_7201,N_4456,N_1663);
or U7202 (N_7202,N_226,N_1735);
xnor U7203 (N_7203,N_2113,N_1761);
xor U7204 (N_7204,N_310,N_1401);
or U7205 (N_7205,N_4029,N_1745);
or U7206 (N_7206,N_2566,N_2363);
nor U7207 (N_7207,N_4255,N_4680);
nor U7208 (N_7208,N_4970,N_3587);
nand U7209 (N_7209,N_3423,N_3754);
or U7210 (N_7210,N_1012,N_4683);
xor U7211 (N_7211,N_2857,N_3026);
xor U7212 (N_7212,N_1009,N_4388);
xnor U7213 (N_7213,N_235,N_1079);
or U7214 (N_7214,N_22,N_1391);
xor U7215 (N_7215,N_1362,N_2918);
nand U7216 (N_7216,N_4863,N_1589);
or U7217 (N_7217,N_209,N_1961);
or U7218 (N_7218,N_4980,N_3247);
nor U7219 (N_7219,N_3127,N_1438);
nand U7220 (N_7220,N_187,N_444);
xor U7221 (N_7221,N_1004,N_3498);
xnor U7222 (N_7222,N_362,N_2660);
nand U7223 (N_7223,N_2961,N_4323);
nand U7224 (N_7224,N_2381,N_4441);
and U7225 (N_7225,N_4398,N_2848);
or U7226 (N_7226,N_4356,N_4267);
or U7227 (N_7227,N_3905,N_2966);
or U7228 (N_7228,N_4999,N_3617);
and U7229 (N_7229,N_3703,N_4632);
xor U7230 (N_7230,N_3005,N_1419);
xor U7231 (N_7231,N_1451,N_378);
nand U7232 (N_7232,N_3938,N_3775);
xnor U7233 (N_7233,N_1267,N_2880);
and U7234 (N_7234,N_4048,N_1302);
nor U7235 (N_7235,N_2242,N_1448);
nand U7236 (N_7236,N_4208,N_1206);
nor U7237 (N_7237,N_3875,N_1638);
nor U7238 (N_7238,N_1856,N_4152);
or U7239 (N_7239,N_3402,N_3638);
xor U7240 (N_7240,N_238,N_1842);
and U7241 (N_7241,N_2383,N_3625);
and U7242 (N_7242,N_2868,N_4453);
nor U7243 (N_7243,N_396,N_4001);
xor U7244 (N_7244,N_1768,N_3628);
xor U7245 (N_7245,N_4521,N_1615);
xor U7246 (N_7246,N_462,N_4021);
xor U7247 (N_7247,N_1410,N_2589);
nor U7248 (N_7248,N_493,N_3512);
or U7249 (N_7249,N_3301,N_2167);
or U7250 (N_7250,N_89,N_4274);
xor U7251 (N_7251,N_3100,N_1789);
or U7252 (N_7252,N_549,N_3235);
or U7253 (N_7253,N_3180,N_884);
nor U7254 (N_7254,N_730,N_2413);
or U7255 (N_7255,N_2590,N_51);
and U7256 (N_7256,N_3227,N_2270);
nor U7257 (N_7257,N_4927,N_3133);
and U7258 (N_7258,N_3206,N_1358);
nand U7259 (N_7259,N_215,N_2948);
xor U7260 (N_7260,N_687,N_2709);
xor U7261 (N_7261,N_435,N_1336);
xor U7262 (N_7262,N_989,N_2971);
and U7263 (N_7263,N_447,N_2015);
or U7264 (N_7264,N_3229,N_3269);
and U7265 (N_7265,N_3141,N_3401);
xor U7266 (N_7266,N_3085,N_1755);
or U7267 (N_7267,N_4438,N_3911);
nor U7268 (N_7268,N_2067,N_4376);
and U7269 (N_7269,N_1152,N_1394);
nand U7270 (N_7270,N_718,N_2736);
or U7271 (N_7271,N_4158,N_3982);
xor U7272 (N_7272,N_3403,N_4038);
nand U7273 (N_7273,N_2954,N_757);
xor U7274 (N_7274,N_3222,N_2705);
nor U7275 (N_7275,N_4206,N_3308);
and U7276 (N_7276,N_3178,N_437);
xor U7277 (N_7277,N_588,N_459);
xnor U7278 (N_7278,N_1903,N_821);
xnor U7279 (N_7279,N_1205,N_3316);
nand U7280 (N_7280,N_1317,N_236);
or U7281 (N_7281,N_228,N_2073);
nand U7282 (N_7282,N_445,N_1107);
xnor U7283 (N_7283,N_2735,N_4587);
or U7284 (N_7284,N_2605,N_1145);
or U7285 (N_7285,N_3590,N_3200);
xor U7286 (N_7286,N_979,N_509);
nand U7287 (N_7287,N_3080,N_2749);
and U7288 (N_7288,N_4498,N_2244);
nor U7289 (N_7289,N_552,N_2896);
nor U7290 (N_7290,N_4845,N_4330);
and U7291 (N_7291,N_2941,N_3344);
or U7292 (N_7292,N_1252,N_1712);
nor U7293 (N_7293,N_3577,N_4368);
nor U7294 (N_7294,N_2787,N_2791);
nor U7295 (N_7295,N_1458,N_981);
xnor U7296 (N_7296,N_4849,N_4522);
and U7297 (N_7297,N_2670,N_2849);
or U7298 (N_7298,N_466,N_3633);
xnor U7299 (N_7299,N_573,N_871);
nand U7300 (N_7300,N_940,N_3302);
xor U7301 (N_7301,N_2269,N_4513);
or U7302 (N_7302,N_4006,N_1498);
or U7303 (N_7303,N_3041,N_2674);
nand U7304 (N_7304,N_2110,N_1969);
or U7305 (N_7305,N_4730,N_4326);
nand U7306 (N_7306,N_3988,N_4654);
xor U7307 (N_7307,N_3848,N_4131);
and U7308 (N_7308,N_1078,N_813);
xor U7309 (N_7309,N_2035,N_3785);
xnor U7310 (N_7310,N_3545,N_4406);
nor U7311 (N_7311,N_3385,N_1571);
nand U7312 (N_7312,N_3901,N_3708);
nand U7313 (N_7313,N_4551,N_3949);
and U7314 (N_7314,N_4121,N_1237);
or U7315 (N_7315,N_662,N_1010);
or U7316 (N_7316,N_4613,N_3194);
or U7317 (N_7317,N_1406,N_3098);
nor U7318 (N_7318,N_132,N_2440);
or U7319 (N_7319,N_3486,N_1582);
xnor U7320 (N_7320,N_2663,N_1897);
xnor U7321 (N_7321,N_3118,N_1569);
nand U7322 (N_7322,N_4931,N_320);
and U7323 (N_7323,N_2867,N_1733);
nand U7324 (N_7324,N_472,N_856);
xor U7325 (N_7325,N_1696,N_1154);
xor U7326 (N_7326,N_3958,N_2515);
nor U7327 (N_7327,N_1986,N_4719);
nor U7328 (N_7328,N_3522,N_1380);
nor U7329 (N_7329,N_4072,N_1596);
or U7330 (N_7330,N_2465,N_758);
or U7331 (N_7331,N_2659,N_4633);
or U7332 (N_7332,N_4792,N_3885);
and U7333 (N_7333,N_2406,N_203);
and U7334 (N_7334,N_4662,N_2828);
or U7335 (N_7335,N_1065,N_4905);
nand U7336 (N_7336,N_4659,N_4423);
nor U7337 (N_7337,N_4317,N_3494);
nand U7338 (N_7338,N_4681,N_1953);
and U7339 (N_7339,N_1180,N_2054);
and U7340 (N_7340,N_795,N_3640);
and U7341 (N_7341,N_3071,N_1189);
or U7342 (N_7342,N_402,N_341);
nor U7343 (N_7343,N_2859,N_2769);
and U7344 (N_7344,N_4122,N_555);
or U7345 (N_7345,N_2329,N_3477);
nand U7346 (N_7346,N_213,N_3170);
and U7347 (N_7347,N_1951,N_4110);
nand U7348 (N_7348,N_4106,N_4902);
nor U7349 (N_7349,N_3676,N_141);
xnor U7350 (N_7350,N_906,N_3289);
nor U7351 (N_7351,N_857,N_1666);
and U7352 (N_7352,N_2149,N_3506);
nand U7353 (N_7353,N_1360,N_4693);
or U7354 (N_7354,N_2063,N_2963);
or U7355 (N_7355,N_4981,N_794);
and U7356 (N_7356,N_2718,N_1005);
nand U7357 (N_7357,N_1048,N_1427);
nand U7358 (N_7358,N_384,N_1230);
nand U7359 (N_7359,N_1942,N_318);
nand U7360 (N_7360,N_534,N_603);
or U7361 (N_7361,N_4701,N_333);
or U7362 (N_7362,N_2619,N_3359);
or U7363 (N_7363,N_1763,N_2733);
xnor U7364 (N_7364,N_4583,N_4112);
nor U7365 (N_7365,N_4671,N_4489);
xnor U7366 (N_7366,N_2752,N_3253);
and U7367 (N_7367,N_3519,N_4776);
nor U7368 (N_7368,N_2788,N_949);
xnor U7369 (N_7369,N_3817,N_2933);
and U7370 (N_7370,N_2365,N_4143);
and U7371 (N_7371,N_4316,N_3288);
or U7372 (N_7372,N_1729,N_72);
nand U7373 (N_7373,N_888,N_1898);
nor U7374 (N_7374,N_1243,N_2316);
nor U7375 (N_7375,N_3415,N_1680);
and U7376 (N_7376,N_3491,N_371);
or U7377 (N_7377,N_4771,N_4674);
or U7378 (N_7378,N_3668,N_2955);
nor U7379 (N_7379,N_3162,N_2903);
or U7380 (N_7380,N_756,N_3020);
or U7381 (N_7381,N_321,N_640);
nor U7382 (N_7382,N_907,N_4075);
nand U7383 (N_7383,N_405,N_3702);
and U7384 (N_7384,N_3564,N_66);
or U7385 (N_7385,N_1208,N_3298);
xnor U7386 (N_7386,N_2831,N_3828);
or U7387 (N_7387,N_4645,N_28);
nor U7388 (N_7388,N_1253,N_4556);
nor U7389 (N_7389,N_4113,N_3914);
xnor U7390 (N_7390,N_1698,N_2146);
and U7391 (N_7391,N_3339,N_4347);
xor U7392 (N_7392,N_4748,N_2815);
nor U7393 (N_7393,N_3420,N_3318);
xor U7394 (N_7394,N_3209,N_3504);
or U7395 (N_7395,N_3120,N_876);
nor U7396 (N_7396,N_3191,N_2851);
and U7397 (N_7397,N_319,N_4795);
or U7398 (N_7398,N_486,N_3547);
or U7399 (N_7399,N_401,N_2745);
xor U7400 (N_7400,N_3738,N_1769);
and U7401 (N_7401,N_4425,N_4575);
nand U7402 (N_7402,N_4266,N_3765);
or U7403 (N_7403,N_4473,N_3452);
or U7404 (N_7404,N_2658,N_4986);
nor U7405 (N_7405,N_2103,N_4913);
and U7406 (N_7406,N_2635,N_2104);
nand U7407 (N_7407,N_925,N_1950);
nor U7408 (N_7408,N_3104,N_2837);
nor U7409 (N_7409,N_2694,N_4865);
nand U7410 (N_7410,N_3659,N_604);
xnor U7411 (N_7411,N_2024,N_1619);
nand U7412 (N_7412,N_4271,N_2273);
nand U7413 (N_7413,N_1626,N_2423);
xnor U7414 (N_7414,N_376,N_2753);
and U7415 (N_7415,N_4761,N_4791);
nor U7416 (N_7416,N_2853,N_3516);
nor U7417 (N_7417,N_1248,N_768);
xor U7418 (N_7418,N_3822,N_826);
xnor U7419 (N_7419,N_4808,N_431);
xnor U7420 (N_7420,N_2097,N_737);
and U7421 (N_7421,N_1246,N_4400);
or U7422 (N_7422,N_2858,N_2312);
nor U7423 (N_7423,N_178,N_4030);
nand U7424 (N_7424,N_637,N_918);
or U7425 (N_7425,N_1348,N_4137);
nand U7426 (N_7426,N_1600,N_537);
xor U7427 (N_7427,N_4641,N_3684);
and U7428 (N_7428,N_446,N_4673);
xnor U7429 (N_7429,N_464,N_859);
nor U7430 (N_7430,N_4300,N_713);
nor U7431 (N_7431,N_2325,N_692);
and U7432 (N_7432,N_1300,N_338);
or U7433 (N_7433,N_1135,N_4864);
nand U7434 (N_7434,N_2057,N_3710);
nor U7435 (N_7435,N_2184,N_3960);
nor U7436 (N_7436,N_3892,N_1185);
or U7437 (N_7437,N_4493,N_4882);
or U7438 (N_7438,N_1222,N_4852);
xnor U7439 (N_7439,N_1286,N_561);
nand U7440 (N_7440,N_1966,N_4309);
or U7441 (N_7441,N_2616,N_4944);
nor U7442 (N_7442,N_1637,N_1873);
xor U7443 (N_7443,N_2949,N_3082);
xor U7444 (N_7444,N_488,N_2260);
nand U7445 (N_7445,N_2936,N_1687);
or U7446 (N_7446,N_2937,N_4142);
nor U7447 (N_7447,N_2992,N_3424);
and U7448 (N_7448,N_3556,N_3260);
nand U7449 (N_7449,N_2172,N_4786);
nor U7450 (N_7450,N_948,N_82);
nor U7451 (N_7451,N_2134,N_4725);
or U7452 (N_7452,N_2215,N_3962);
nor U7453 (N_7453,N_2601,N_950);
nand U7454 (N_7454,N_390,N_2354);
nand U7455 (N_7455,N_1365,N_928);
and U7456 (N_7456,N_518,N_1740);
nor U7457 (N_7457,N_2121,N_584);
and U7458 (N_7458,N_4146,N_2453);
nor U7459 (N_7459,N_4729,N_2285);
xor U7460 (N_7460,N_1441,N_2689);
nor U7461 (N_7461,N_816,N_1629);
and U7462 (N_7462,N_984,N_3826);
nand U7463 (N_7463,N_1106,N_4835);
nor U7464 (N_7464,N_171,N_2765);
xor U7465 (N_7465,N_2180,N_1506);
xnor U7466 (N_7466,N_4025,N_1811);
nor U7467 (N_7467,N_4457,N_3430);
or U7468 (N_7468,N_2847,N_4474);
or U7469 (N_7469,N_3121,N_2004);
or U7470 (N_7470,N_2716,N_2350);
xnor U7471 (N_7471,N_283,N_1748);
nand U7472 (N_7472,N_3212,N_2520);
and U7473 (N_7473,N_1900,N_4658);
xor U7474 (N_7474,N_982,N_1539);
nor U7475 (N_7475,N_2208,N_1534);
or U7476 (N_7476,N_2298,N_167);
nor U7477 (N_7477,N_2826,N_4968);
or U7478 (N_7478,N_2307,N_3745);
and U7479 (N_7479,N_1091,N_1334);
xor U7480 (N_7480,N_3195,N_3932);
xnor U7481 (N_7481,N_3563,N_4605);
nand U7482 (N_7482,N_3432,N_3241);
and U7483 (N_7483,N_3664,N_1018);
and U7484 (N_7484,N_3290,N_247);
and U7485 (N_7485,N_1270,N_448);
nor U7486 (N_7486,N_1826,N_3375);
and U7487 (N_7487,N_270,N_1357);
nand U7488 (N_7488,N_4042,N_4114);
nand U7489 (N_7489,N_833,N_2085);
nor U7490 (N_7490,N_4840,N_527);
xnor U7491 (N_7491,N_3788,N_571);
xnor U7492 (N_7492,N_797,N_4499);
xor U7493 (N_7493,N_4069,N_707);
nor U7494 (N_7494,N_46,N_4327);
or U7495 (N_7495,N_4930,N_2794);
xor U7496 (N_7496,N_1147,N_3523);
or U7497 (N_7497,N_3656,N_4205);
xnor U7498 (N_7498,N_3455,N_1783);
and U7499 (N_7499,N_1824,N_4287);
xor U7500 (N_7500,N_951,N_2296);
nand U7501 (N_7501,N_1528,N_727);
and U7502 (N_7502,N_1126,N_2019);
or U7503 (N_7503,N_3603,N_4839);
nor U7504 (N_7504,N_3403,N_2250);
and U7505 (N_7505,N_3202,N_3011);
xnor U7506 (N_7506,N_951,N_2378);
or U7507 (N_7507,N_491,N_4805);
nor U7508 (N_7508,N_4550,N_4835);
and U7509 (N_7509,N_2856,N_4144);
nor U7510 (N_7510,N_3776,N_2187);
xnor U7511 (N_7511,N_2501,N_211);
and U7512 (N_7512,N_3096,N_4951);
or U7513 (N_7513,N_472,N_2769);
or U7514 (N_7514,N_3052,N_616);
nand U7515 (N_7515,N_4837,N_2944);
and U7516 (N_7516,N_2974,N_1884);
xnor U7517 (N_7517,N_1295,N_2574);
nor U7518 (N_7518,N_848,N_3928);
xor U7519 (N_7519,N_1199,N_526);
and U7520 (N_7520,N_4978,N_1091);
or U7521 (N_7521,N_356,N_2721);
xnor U7522 (N_7522,N_2952,N_73);
nand U7523 (N_7523,N_4855,N_4843);
or U7524 (N_7524,N_204,N_3912);
or U7525 (N_7525,N_3570,N_2015);
or U7526 (N_7526,N_3118,N_2769);
nor U7527 (N_7527,N_3725,N_501);
or U7528 (N_7528,N_3407,N_4589);
and U7529 (N_7529,N_3758,N_440);
nor U7530 (N_7530,N_4324,N_54);
nand U7531 (N_7531,N_936,N_3254);
xnor U7532 (N_7532,N_685,N_2576);
xnor U7533 (N_7533,N_3479,N_4172);
nor U7534 (N_7534,N_606,N_4164);
nor U7535 (N_7535,N_980,N_2049);
xnor U7536 (N_7536,N_2041,N_2524);
xor U7537 (N_7537,N_2039,N_2019);
or U7538 (N_7538,N_4895,N_704);
nor U7539 (N_7539,N_4205,N_36);
nand U7540 (N_7540,N_2830,N_3710);
nor U7541 (N_7541,N_525,N_3217);
xnor U7542 (N_7542,N_513,N_2708);
nor U7543 (N_7543,N_2677,N_768);
and U7544 (N_7544,N_4542,N_2936);
or U7545 (N_7545,N_237,N_1654);
and U7546 (N_7546,N_2333,N_2006);
nand U7547 (N_7547,N_4163,N_920);
xor U7548 (N_7548,N_3978,N_2164);
xnor U7549 (N_7549,N_1481,N_4972);
nand U7550 (N_7550,N_2024,N_1687);
or U7551 (N_7551,N_677,N_1951);
and U7552 (N_7552,N_2988,N_2329);
xnor U7553 (N_7553,N_445,N_3267);
and U7554 (N_7554,N_1807,N_3612);
or U7555 (N_7555,N_767,N_2194);
or U7556 (N_7556,N_4979,N_919);
nand U7557 (N_7557,N_4751,N_1689);
nand U7558 (N_7558,N_594,N_2193);
or U7559 (N_7559,N_2899,N_1899);
nand U7560 (N_7560,N_3256,N_4197);
and U7561 (N_7561,N_3308,N_2486);
nor U7562 (N_7562,N_3214,N_1284);
nor U7563 (N_7563,N_1397,N_1678);
and U7564 (N_7564,N_2510,N_2697);
or U7565 (N_7565,N_2173,N_872);
or U7566 (N_7566,N_1822,N_4800);
or U7567 (N_7567,N_3477,N_4464);
or U7568 (N_7568,N_1539,N_1498);
nand U7569 (N_7569,N_4341,N_134);
and U7570 (N_7570,N_1639,N_1814);
and U7571 (N_7571,N_3593,N_4922);
and U7572 (N_7572,N_4456,N_2865);
nor U7573 (N_7573,N_3904,N_2805);
xnor U7574 (N_7574,N_1094,N_191);
or U7575 (N_7575,N_2633,N_1372);
xor U7576 (N_7576,N_4539,N_876);
nand U7577 (N_7577,N_525,N_2593);
nand U7578 (N_7578,N_1378,N_39);
xor U7579 (N_7579,N_1808,N_3709);
nand U7580 (N_7580,N_3025,N_2092);
and U7581 (N_7581,N_3943,N_3103);
nor U7582 (N_7582,N_4395,N_53);
and U7583 (N_7583,N_947,N_2521);
and U7584 (N_7584,N_3056,N_3448);
or U7585 (N_7585,N_1009,N_2023);
xnor U7586 (N_7586,N_4501,N_2091);
and U7587 (N_7587,N_1354,N_4925);
xnor U7588 (N_7588,N_3113,N_3636);
or U7589 (N_7589,N_595,N_4979);
nand U7590 (N_7590,N_762,N_2561);
nor U7591 (N_7591,N_1258,N_2939);
xnor U7592 (N_7592,N_3239,N_4465);
or U7593 (N_7593,N_1544,N_2600);
nand U7594 (N_7594,N_2096,N_647);
and U7595 (N_7595,N_2855,N_3961);
or U7596 (N_7596,N_4062,N_366);
nor U7597 (N_7597,N_4106,N_354);
and U7598 (N_7598,N_453,N_912);
xor U7599 (N_7599,N_3560,N_3594);
nand U7600 (N_7600,N_2776,N_3515);
and U7601 (N_7601,N_693,N_3415);
xnor U7602 (N_7602,N_390,N_4430);
and U7603 (N_7603,N_2349,N_4266);
and U7604 (N_7604,N_2723,N_4283);
xnor U7605 (N_7605,N_662,N_73);
nor U7606 (N_7606,N_2339,N_2399);
xnor U7607 (N_7607,N_2580,N_1605);
and U7608 (N_7608,N_3820,N_2406);
and U7609 (N_7609,N_1912,N_4705);
and U7610 (N_7610,N_4587,N_2986);
nor U7611 (N_7611,N_2616,N_3917);
nor U7612 (N_7612,N_94,N_1685);
or U7613 (N_7613,N_2645,N_1686);
or U7614 (N_7614,N_2676,N_347);
nand U7615 (N_7615,N_400,N_3960);
xnor U7616 (N_7616,N_4816,N_817);
and U7617 (N_7617,N_2241,N_1481);
nand U7618 (N_7618,N_1945,N_2639);
and U7619 (N_7619,N_1351,N_4610);
or U7620 (N_7620,N_2929,N_1948);
or U7621 (N_7621,N_4009,N_4653);
and U7622 (N_7622,N_1463,N_2669);
nor U7623 (N_7623,N_3564,N_319);
xor U7624 (N_7624,N_954,N_484);
nor U7625 (N_7625,N_2501,N_901);
and U7626 (N_7626,N_1671,N_3387);
xor U7627 (N_7627,N_3436,N_2769);
nand U7628 (N_7628,N_3707,N_2967);
nor U7629 (N_7629,N_1428,N_237);
nor U7630 (N_7630,N_448,N_2411);
xor U7631 (N_7631,N_4837,N_1540);
nand U7632 (N_7632,N_1217,N_4715);
or U7633 (N_7633,N_3716,N_3610);
and U7634 (N_7634,N_3871,N_3394);
xor U7635 (N_7635,N_1329,N_4768);
or U7636 (N_7636,N_3418,N_4733);
nor U7637 (N_7637,N_175,N_133);
nand U7638 (N_7638,N_1602,N_3614);
nor U7639 (N_7639,N_4186,N_1605);
nand U7640 (N_7640,N_2251,N_4665);
and U7641 (N_7641,N_2174,N_2861);
and U7642 (N_7642,N_946,N_351);
or U7643 (N_7643,N_4504,N_987);
nor U7644 (N_7644,N_4172,N_3074);
nor U7645 (N_7645,N_1613,N_467);
or U7646 (N_7646,N_2673,N_249);
xor U7647 (N_7647,N_772,N_1423);
nand U7648 (N_7648,N_1687,N_631);
or U7649 (N_7649,N_1601,N_2204);
and U7650 (N_7650,N_4951,N_828);
nand U7651 (N_7651,N_2986,N_3435);
or U7652 (N_7652,N_4396,N_1126);
xor U7653 (N_7653,N_2015,N_3534);
nand U7654 (N_7654,N_2902,N_3265);
xor U7655 (N_7655,N_1248,N_424);
nand U7656 (N_7656,N_3532,N_574);
nor U7657 (N_7657,N_2543,N_2477);
nand U7658 (N_7658,N_2959,N_3853);
and U7659 (N_7659,N_54,N_4335);
xor U7660 (N_7660,N_4115,N_3933);
or U7661 (N_7661,N_2616,N_2790);
nand U7662 (N_7662,N_1135,N_3341);
and U7663 (N_7663,N_471,N_4999);
nor U7664 (N_7664,N_296,N_2545);
nand U7665 (N_7665,N_4295,N_3679);
nand U7666 (N_7666,N_920,N_2288);
nand U7667 (N_7667,N_4658,N_4668);
and U7668 (N_7668,N_2860,N_118);
nor U7669 (N_7669,N_4427,N_4165);
xnor U7670 (N_7670,N_2462,N_617);
nand U7671 (N_7671,N_848,N_900);
or U7672 (N_7672,N_2232,N_3208);
nand U7673 (N_7673,N_1101,N_2697);
nor U7674 (N_7674,N_1727,N_3765);
xor U7675 (N_7675,N_1355,N_3141);
and U7676 (N_7676,N_3807,N_3423);
or U7677 (N_7677,N_1808,N_1316);
and U7678 (N_7678,N_4435,N_382);
or U7679 (N_7679,N_4355,N_2825);
and U7680 (N_7680,N_1935,N_1381);
and U7681 (N_7681,N_3372,N_4516);
nand U7682 (N_7682,N_2972,N_3863);
and U7683 (N_7683,N_1552,N_234);
and U7684 (N_7684,N_3523,N_3824);
xnor U7685 (N_7685,N_1891,N_3929);
or U7686 (N_7686,N_4893,N_3887);
xnor U7687 (N_7687,N_4836,N_2621);
and U7688 (N_7688,N_4027,N_1008);
and U7689 (N_7689,N_1158,N_1734);
nor U7690 (N_7690,N_3731,N_2030);
nand U7691 (N_7691,N_2868,N_1534);
xor U7692 (N_7692,N_3706,N_1131);
and U7693 (N_7693,N_3025,N_2322);
xor U7694 (N_7694,N_523,N_477);
xnor U7695 (N_7695,N_3442,N_2194);
or U7696 (N_7696,N_4779,N_1250);
or U7697 (N_7697,N_568,N_4479);
xor U7698 (N_7698,N_3459,N_2660);
xor U7699 (N_7699,N_1217,N_50);
nor U7700 (N_7700,N_4355,N_4904);
nand U7701 (N_7701,N_4040,N_3343);
nor U7702 (N_7702,N_493,N_2674);
nand U7703 (N_7703,N_2331,N_2574);
nor U7704 (N_7704,N_1800,N_2537);
xor U7705 (N_7705,N_4593,N_1752);
and U7706 (N_7706,N_4307,N_3468);
or U7707 (N_7707,N_2034,N_323);
or U7708 (N_7708,N_3585,N_1362);
nand U7709 (N_7709,N_494,N_641);
or U7710 (N_7710,N_2493,N_499);
or U7711 (N_7711,N_1140,N_2165);
and U7712 (N_7712,N_2415,N_1009);
nand U7713 (N_7713,N_1397,N_1273);
or U7714 (N_7714,N_2394,N_2531);
nor U7715 (N_7715,N_679,N_548);
xor U7716 (N_7716,N_2056,N_3452);
xor U7717 (N_7717,N_2107,N_4929);
xor U7718 (N_7718,N_2227,N_1423);
xnor U7719 (N_7719,N_171,N_4687);
or U7720 (N_7720,N_211,N_3809);
xnor U7721 (N_7721,N_817,N_2349);
nand U7722 (N_7722,N_4281,N_956);
nand U7723 (N_7723,N_4998,N_3795);
nand U7724 (N_7724,N_4535,N_1692);
or U7725 (N_7725,N_3684,N_3072);
nor U7726 (N_7726,N_4573,N_3104);
nor U7727 (N_7727,N_3596,N_4833);
nand U7728 (N_7728,N_3539,N_2394);
nand U7729 (N_7729,N_4989,N_3825);
nor U7730 (N_7730,N_3327,N_3214);
or U7731 (N_7731,N_3202,N_495);
nor U7732 (N_7732,N_489,N_3972);
xnor U7733 (N_7733,N_3535,N_2054);
xnor U7734 (N_7734,N_2208,N_4031);
and U7735 (N_7735,N_989,N_3282);
or U7736 (N_7736,N_2086,N_1332);
nor U7737 (N_7737,N_4959,N_1363);
xnor U7738 (N_7738,N_1124,N_3947);
or U7739 (N_7739,N_2095,N_2590);
xor U7740 (N_7740,N_479,N_2954);
or U7741 (N_7741,N_4621,N_110);
xor U7742 (N_7742,N_2544,N_1040);
nand U7743 (N_7743,N_1026,N_4046);
xor U7744 (N_7744,N_4667,N_228);
and U7745 (N_7745,N_956,N_3047);
and U7746 (N_7746,N_1890,N_4329);
nand U7747 (N_7747,N_2617,N_655);
or U7748 (N_7748,N_4943,N_1028);
or U7749 (N_7749,N_2737,N_4681);
or U7750 (N_7750,N_4949,N_4654);
xor U7751 (N_7751,N_490,N_2953);
nand U7752 (N_7752,N_1568,N_871);
nor U7753 (N_7753,N_4993,N_1837);
or U7754 (N_7754,N_4161,N_3381);
nand U7755 (N_7755,N_781,N_1181);
xnor U7756 (N_7756,N_1504,N_4835);
nand U7757 (N_7757,N_293,N_4505);
nor U7758 (N_7758,N_4788,N_4627);
nor U7759 (N_7759,N_1387,N_2245);
and U7760 (N_7760,N_4319,N_2247);
xnor U7761 (N_7761,N_4042,N_2124);
nor U7762 (N_7762,N_327,N_3289);
nand U7763 (N_7763,N_761,N_1468);
or U7764 (N_7764,N_2365,N_859);
nand U7765 (N_7765,N_1141,N_1307);
or U7766 (N_7766,N_3856,N_1507);
or U7767 (N_7767,N_3054,N_897);
nor U7768 (N_7768,N_767,N_614);
nand U7769 (N_7769,N_4557,N_2217);
nor U7770 (N_7770,N_1677,N_3394);
xor U7771 (N_7771,N_1874,N_4107);
nor U7772 (N_7772,N_4427,N_2818);
xnor U7773 (N_7773,N_1333,N_2480);
nor U7774 (N_7774,N_4772,N_2894);
nand U7775 (N_7775,N_2097,N_3221);
nand U7776 (N_7776,N_4910,N_4978);
or U7777 (N_7777,N_997,N_2855);
xor U7778 (N_7778,N_143,N_4987);
and U7779 (N_7779,N_4896,N_4911);
nor U7780 (N_7780,N_4643,N_1634);
xor U7781 (N_7781,N_4193,N_3047);
xor U7782 (N_7782,N_4683,N_1304);
nor U7783 (N_7783,N_2362,N_1728);
and U7784 (N_7784,N_1003,N_2156);
or U7785 (N_7785,N_783,N_2465);
nor U7786 (N_7786,N_2375,N_4517);
and U7787 (N_7787,N_1957,N_1545);
and U7788 (N_7788,N_1902,N_1091);
nor U7789 (N_7789,N_3662,N_717);
nor U7790 (N_7790,N_3861,N_2067);
nor U7791 (N_7791,N_3453,N_90);
nor U7792 (N_7792,N_157,N_2500);
xnor U7793 (N_7793,N_4690,N_2345);
nor U7794 (N_7794,N_3891,N_3067);
nor U7795 (N_7795,N_4256,N_1019);
nand U7796 (N_7796,N_4599,N_3940);
nor U7797 (N_7797,N_1053,N_3520);
nor U7798 (N_7798,N_3125,N_3248);
nor U7799 (N_7799,N_1321,N_2398);
nor U7800 (N_7800,N_4072,N_3611);
or U7801 (N_7801,N_4996,N_3624);
and U7802 (N_7802,N_4111,N_2869);
or U7803 (N_7803,N_1366,N_2062);
and U7804 (N_7804,N_2219,N_2773);
nand U7805 (N_7805,N_4134,N_191);
and U7806 (N_7806,N_972,N_457);
or U7807 (N_7807,N_1666,N_2684);
nor U7808 (N_7808,N_849,N_4087);
xnor U7809 (N_7809,N_3295,N_590);
and U7810 (N_7810,N_3991,N_2955);
or U7811 (N_7811,N_82,N_633);
xor U7812 (N_7812,N_904,N_4031);
and U7813 (N_7813,N_3389,N_2290);
nand U7814 (N_7814,N_1738,N_4211);
nand U7815 (N_7815,N_2315,N_165);
nor U7816 (N_7816,N_3491,N_2228);
nor U7817 (N_7817,N_3871,N_3857);
nand U7818 (N_7818,N_2280,N_538);
nand U7819 (N_7819,N_103,N_218);
nor U7820 (N_7820,N_2545,N_4585);
nand U7821 (N_7821,N_1470,N_4840);
nor U7822 (N_7822,N_1654,N_4326);
or U7823 (N_7823,N_1023,N_446);
nor U7824 (N_7824,N_2208,N_2054);
nand U7825 (N_7825,N_3972,N_3172);
and U7826 (N_7826,N_1898,N_784);
or U7827 (N_7827,N_3464,N_3056);
nor U7828 (N_7828,N_4183,N_3839);
or U7829 (N_7829,N_1027,N_3516);
or U7830 (N_7830,N_4830,N_997);
xor U7831 (N_7831,N_3119,N_3616);
nand U7832 (N_7832,N_1822,N_4771);
and U7833 (N_7833,N_2625,N_3948);
xnor U7834 (N_7834,N_2910,N_2706);
and U7835 (N_7835,N_4723,N_3539);
xor U7836 (N_7836,N_2134,N_1139);
and U7837 (N_7837,N_2047,N_3860);
nor U7838 (N_7838,N_496,N_4087);
nor U7839 (N_7839,N_4681,N_4352);
nand U7840 (N_7840,N_1568,N_4678);
or U7841 (N_7841,N_411,N_4201);
or U7842 (N_7842,N_2926,N_4611);
nor U7843 (N_7843,N_301,N_4625);
and U7844 (N_7844,N_2777,N_3184);
and U7845 (N_7845,N_1167,N_2873);
xor U7846 (N_7846,N_1920,N_4284);
or U7847 (N_7847,N_2585,N_1763);
nor U7848 (N_7848,N_2641,N_2723);
nand U7849 (N_7849,N_2172,N_1775);
nor U7850 (N_7850,N_733,N_1173);
and U7851 (N_7851,N_3416,N_4685);
or U7852 (N_7852,N_3463,N_4029);
xor U7853 (N_7853,N_3954,N_4239);
and U7854 (N_7854,N_3120,N_3228);
xnor U7855 (N_7855,N_1262,N_1465);
nand U7856 (N_7856,N_906,N_2581);
nor U7857 (N_7857,N_3311,N_2899);
nand U7858 (N_7858,N_4803,N_364);
nor U7859 (N_7859,N_275,N_479);
nor U7860 (N_7860,N_4807,N_3305);
nand U7861 (N_7861,N_1784,N_3098);
nand U7862 (N_7862,N_4391,N_23);
nor U7863 (N_7863,N_364,N_573);
or U7864 (N_7864,N_1797,N_1233);
nor U7865 (N_7865,N_3410,N_4491);
nand U7866 (N_7866,N_4617,N_459);
xnor U7867 (N_7867,N_4563,N_961);
nor U7868 (N_7868,N_2638,N_811);
xor U7869 (N_7869,N_666,N_4673);
nor U7870 (N_7870,N_2081,N_142);
nand U7871 (N_7871,N_3125,N_1557);
xor U7872 (N_7872,N_3767,N_1722);
or U7873 (N_7873,N_944,N_4483);
and U7874 (N_7874,N_3179,N_2862);
xnor U7875 (N_7875,N_3905,N_1698);
and U7876 (N_7876,N_3376,N_3650);
nand U7877 (N_7877,N_807,N_3951);
nand U7878 (N_7878,N_1901,N_1057);
or U7879 (N_7879,N_1419,N_220);
nor U7880 (N_7880,N_1596,N_666);
and U7881 (N_7881,N_691,N_1136);
xor U7882 (N_7882,N_143,N_4394);
xnor U7883 (N_7883,N_4388,N_1319);
and U7884 (N_7884,N_4413,N_3271);
xnor U7885 (N_7885,N_690,N_2484);
or U7886 (N_7886,N_788,N_3030);
nand U7887 (N_7887,N_3267,N_1385);
and U7888 (N_7888,N_506,N_1494);
and U7889 (N_7889,N_637,N_3606);
nand U7890 (N_7890,N_4429,N_2359);
or U7891 (N_7891,N_4858,N_1745);
and U7892 (N_7892,N_2251,N_3556);
and U7893 (N_7893,N_1054,N_4805);
nor U7894 (N_7894,N_293,N_3246);
or U7895 (N_7895,N_4667,N_1011);
nor U7896 (N_7896,N_3161,N_176);
xor U7897 (N_7897,N_1961,N_3679);
nor U7898 (N_7898,N_1742,N_3904);
and U7899 (N_7899,N_2171,N_2007);
or U7900 (N_7900,N_230,N_3455);
and U7901 (N_7901,N_4803,N_4051);
or U7902 (N_7902,N_2533,N_1658);
and U7903 (N_7903,N_4615,N_2148);
nor U7904 (N_7904,N_245,N_904);
or U7905 (N_7905,N_4327,N_3617);
nand U7906 (N_7906,N_4863,N_1624);
and U7907 (N_7907,N_1757,N_798);
and U7908 (N_7908,N_1227,N_699);
xnor U7909 (N_7909,N_4628,N_1207);
nand U7910 (N_7910,N_4462,N_1290);
or U7911 (N_7911,N_2423,N_288);
xor U7912 (N_7912,N_971,N_2684);
and U7913 (N_7913,N_878,N_843);
nand U7914 (N_7914,N_1179,N_4066);
xnor U7915 (N_7915,N_3503,N_4030);
nor U7916 (N_7916,N_3058,N_2789);
xor U7917 (N_7917,N_3999,N_1862);
nor U7918 (N_7918,N_4526,N_2108);
and U7919 (N_7919,N_1321,N_3788);
or U7920 (N_7920,N_1858,N_2993);
and U7921 (N_7921,N_892,N_2816);
and U7922 (N_7922,N_4703,N_2573);
xor U7923 (N_7923,N_696,N_2915);
nor U7924 (N_7924,N_203,N_2490);
or U7925 (N_7925,N_4488,N_366);
nand U7926 (N_7926,N_2066,N_456);
or U7927 (N_7927,N_355,N_3841);
nor U7928 (N_7928,N_2558,N_295);
and U7929 (N_7929,N_1590,N_890);
and U7930 (N_7930,N_2177,N_2612);
xnor U7931 (N_7931,N_4450,N_1598);
nand U7932 (N_7932,N_3233,N_452);
nand U7933 (N_7933,N_2766,N_3039);
nor U7934 (N_7934,N_913,N_4471);
and U7935 (N_7935,N_4909,N_1396);
nor U7936 (N_7936,N_3368,N_299);
or U7937 (N_7937,N_417,N_1321);
and U7938 (N_7938,N_2551,N_1043);
xnor U7939 (N_7939,N_2757,N_542);
xor U7940 (N_7940,N_73,N_652);
and U7941 (N_7941,N_2208,N_2349);
and U7942 (N_7942,N_2255,N_3946);
and U7943 (N_7943,N_465,N_1405);
xnor U7944 (N_7944,N_2026,N_4782);
xor U7945 (N_7945,N_3792,N_4015);
nand U7946 (N_7946,N_4226,N_2810);
and U7947 (N_7947,N_855,N_4495);
nand U7948 (N_7948,N_1929,N_4048);
or U7949 (N_7949,N_934,N_1921);
nand U7950 (N_7950,N_4148,N_3037);
or U7951 (N_7951,N_4983,N_4686);
nor U7952 (N_7952,N_236,N_53);
nor U7953 (N_7953,N_256,N_1720);
xnor U7954 (N_7954,N_3264,N_3863);
nand U7955 (N_7955,N_4626,N_2235);
or U7956 (N_7956,N_1821,N_2387);
and U7957 (N_7957,N_4741,N_190);
xnor U7958 (N_7958,N_3577,N_1932);
nor U7959 (N_7959,N_1045,N_3171);
nor U7960 (N_7960,N_1560,N_647);
xor U7961 (N_7961,N_560,N_606);
xor U7962 (N_7962,N_1483,N_4603);
and U7963 (N_7963,N_172,N_4981);
nand U7964 (N_7964,N_433,N_4147);
nand U7965 (N_7965,N_2729,N_3082);
or U7966 (N_7966,N_569,N_1393);
or U7967 (N_7967,N_53,N_2599);
nor U7968 (N_7968,N_890,N_2342);
and U7969 (N_7969,N_1556,N_476);
xor U7970 (N_7970,N_4058,N_4442);
nand U7971 (N_7971,N_2592,N_1127);
nand U7972 (N_7972,N_1534,N_1787);
nand U7973 (N_7973,N_3771,N_2912);
and U7974 (N_7974,N_589,N_526);
nand U7975 (N_7975,N_3000,N_2587);
nor U7976 (N_7976,N_185,N_4248);
nor U7977 (N_7977,N_4834,N_1488);
nor U7978 (N_7978,N_843,N_1432);
xor U7979 (N_7979,N_4849,N_2451);
nor U7980 (N_7980,N_977,N_1675);
nand U7981 (N_7981,N_2192,N_3804);
xnor U7982 (N_7982,N_1084,N_4635);
nor U7983 (N_7983,N_2008,N_1541);
and U7984 (N_7984,N_3996,N_3216);
xor U7985 (N_7985,N_2594,N_4970);
nor U7986 (N_7986,N_4933,N_4038);
xor U7987 (N_7987,N_718,N_352);
xor U7988 (N_7988,N_3780,N_1995);
xnor U7989 (N_7989,N_3406,N_4647);
nor U7990 (N_7990,N_4151,N_101);
or U7991 (N_7991,N_4280,N_2531);
xnor U7992 (N_7992,N_1286,N_4852);
xor U7993 (N_7993,N_159,N_703);
and U7994 (N_7994,N_2264,N_4624);
and U7995 (N_7995,N_3956,N_2620);
and U7996 (N_7996,N_4115,N_4523);
nor U7997 (N_7997,N_3954,N_2325);
or U7998 (N_7998,N_1502,N_300);
xnor U7999 (N_7999,N_3561,N_4028);
nor U8000 (N_8000,N_2294,N_3731);
or U8001 (N_8001,N_2212,N_1794);
or U8002 (N_8002,N_3692,N_653);
or U8003 (N_8003,N_2159,N_245);
xnor U8004 (N_8004,N_4531,N_657);
and U8005 (N_8005,N_4106,N_1221);
xnor U8006 (N_8006,N_4278,N_1034);
xnor U8007 (N_8007,N_2345,N_913);
and U8008 (N_8008,N_4320,N_496);
or U8009 (N_8009,N_2837,N_54);
or U8010 (N_8010,N_1048,N_660);
and U8011 (N_8011,N_4218,N_3821);
or U8012 (N_8012,N_3914,N_4154);
or U8013 (N_8013,N_95,N_4289);
and U8014 (N_8014,N_4485,N_4063);
xnor U8015 (N_8015,N_449,N_1316);
nor U8016 (N_8016,N_489,N_4872);
xnor U8017 (N_8017,N_3966,N_1959);
and U8018 (N_8018,N_1683,N_267);
nand U8019 (N_8019,N_4242,N_2704);
nor U8020 (N_8020,N_229,N_2776);
nor U8021 (N_8021,N_2344,N_2991);
and U8022 (N_8022,N_2931,N_2204);
and U8023 (N_8023,N_1808,N_1344);
or U8024 (N_8024,N_2769,N_1375);
or U8025 (N_8025,N_4685,N_1902);
nand U8026 (N_8026,N_2091,N_840);
and U8027 (N_8027,N_1953,N_3981);
and U8028 (N_8028,N_1430,N_4513);
xnor U8029 (N_8029,N_2692,N_3666);
nand U8030 (N_8030,N_2976,N_1748);
nand U8031 (N_8031,N_339,N_832);
nor U8032 (N_8032,N_707,N_398);
nor U8033 (N_8033,N_1161,N_4923);
nor U8034 (N_8034,N_2647,N_2717);
xnor U8035 (N_8035,N_1443,N_4022);
nor U8036 (N_8036,N_4540,N_1494);
and U8037 (N_8037,N_10,N_3216);
xnor U8038 (N_8038,N_2762,N_1889);
xor U8039 (N_8039,N_744,N_4984);
or U8040 (N_8040,N_573,N_706);
or U8041 (N_8041,N_153,N_178);
and U8042 (N_8042,N_1598,N_217);
nor U8043 (N_8043,N_2505,N_1093);
nor U8044 (N_8044,N_3015,N_3014);
nor U8045 (N_8045,N_1133,N_3904);
xor U8046 (N_8046,N_3042,N_233);
nor U8047 (N_8047,N_3685,N_3460);
xnor U8048 (N_8048,N_2015,N_1723);
and U8049 (N_8049,N_4715,N_3960);
nor U8050 (N_8050,N_1205,N_1882);
nand U8051 (N_8051,N_4209,N_4964);
or U8052 (N_8052,N_4027,N_4895);
and U8053 (N_8053,N_2977,N_959);
and U8054 (N_8054,N_4107,N_2127);
xnor U8055 (N_8055,N_1772,N_609);
xor U8056 (N_8056,N_2420,N_2103);
or U8057 (N_8057,N_1655,N_1469);
nor U8058 (N_8058,N_3956,N_1889);
nor U8059 (N_8059,N_2572,N_1255);
xnor U8060 (N_8060,N_1750,N_507);
xor U8061 (N_8061,N_3073,N_813);
or U8062 (N_8062,N_400,N_1884);
nor U8063 (N_8063,N_1445,N_2824);
xor U8064 (N_8064,N_2677,N_1982);
and U8065 (N_8065,N_1770,N_3622);
or U8066 (N_8066,N_136,N_4779);
nand U8067 (N_8067,N_758,N_3838);
nor U8068 (N_8068,N_4696,N_1094);
nand U8069 (N_8069,N_470,N_474);
xnor U8070 (N_8070,N_2486,N_4581);
nor U8071 (N_8071,N_1306,N_1980);
nor U8072 (N_8072,N_2248,N_1761);
nand U8073 (N_8073,N_3326,N_4710);
or U8074 (N_8074,N_2710,N_4607);
and U8075 (N_8075,N_2565,N_2397);
or U8076 (N_8076,N_2581,N_2056);
or U8077 (N_8077,N_1399,N_3234);
and U8078 (N_8078,N_1465,N_4261);
or U8079 (N_8079,N_3418,N_1454);
nor U8080 (N_8080,N_474,N_842);
or U8081 (N_8081,N_4155,N_580);
nor U8082 (N_8082,N_266,N_1462);
nand U8083 (N_8083,N_4514,N_2485);
and U8084 (N_8084,N_2228,N_2439);
nand U8085 (N_8085,N_2563,N_1506);
nor U8086 (N_8086,N_2855,N_3797);
nor U8087 (N_8087,N_3713,N_3840);
nand U8088 (N_8088,N_4146,N_3112);
or U8089 (N_8089,N_4886,N_1646);
and U8090 (N_8090,N_459,N_1423);
xor U8091 (N_8091,N_3146,N_1385);
and U8092 (N_8092,N_1435,N_4898);
nor U8093 (N_8093,N_1471,N_2846);
and U8094 (N_8094,N_4374,N_2307);
nor U8095 (N_8095,N_2429,N_6);
or U8096 (N_8096,N_3461,N_4176);
or U8097 (N_8097,N_487,N_441);
xnor U8098 (N_8098,N_2845,N_3966);
nand U8099 (N_8099,N_4516,N_2558);
xor U8100 (N_8100,N_3050,N_385);
nor U8101 (N_8101,N_2425,N_3870);
and U8102 (N_8102,N_4619,N_4133);
or U8103 (N_8103,N_3405,N_4122);
and U8104 (N_8104,N_4213,N_3560);
xor U8105 (N_8105,N_2917,N_4370);
nor U8106 (N_8106,N_1128,N_2400);
nand U8107 (N_8107,N_3158,N_4450);
nor U8108 (N_8108,N_1078,N_2074);
nor U8109 (N_8109,N_1514,N_1081);
or U8110 (N_8110,N_664,N_4933);
or U8111 (N_8111,N_1494,N_4859);
nand U8112 (N_8112,N_4779,N_1914);
nor U8113 (N_8113,N_2079,N_4050);
nand U8114 (N_8114,N_3453,N_3395);
or U8115 (N_8115,N_2859,N_3087);
or U8116 (N_8116,N_102,N_1360);
nand U8117 (N_8117,N_2229,N_529);
nand U8118 (N_8118,N_3722,N_1256);
or U8119 (N_8119,N_3377,N_1588);
nand U8120 (N_8120,N_3863,N_113);
and U8121 (N_8121,N_1967,N_2084);
xnor U8122 (N_8122,N_1573,N_4727);
xor U8123 (N_8123,N_2422,N_4232);
or U8124 (N_8124,N_35,N_4431);
nand U8125 (N_8125,N_3680,N_3731);
or U8126 (N_8126,N_4571,N_2127);
nand U8127 (N_8127,N_2605,N_227);
nand U8128 (N_8128,N_2362,N_3419);
xnor U8129 (N_8129,N_4692,N_4477);
and U8130 (N_8130,N_2133,N_950);
nand U8131 (N_8131,N_1792,N_4244);
nand U8132 (N_8132,N_1083,N_1220);
nand U8133 (N_8133,N_2697,N_1934);
and U8134 (N_8134,N_2911,N_2679);
nand U8135 (N_8135,N_1770,N_2526);
nand U8136 (N_8136,N_4638,N_1147);
and U8137 (N_8137,N_1670,N_4652);
or U8138 (N_8138,N_1010,N_4020);
or U8139 (N_8139,N_1144,N_3302);
xnor U8140 (N_8140,N_23,N_2759);
xnor U8141 (N_8141,N_2803,N_669);
and U8142 (N_8142,N_539,N_2561);
nor U8143 (N_8143,N_3883,N_3576);
or U8144 (N_8144,N_334,N_3002);
nand U8145 (N_8145,N_4790,N_983);
or U8146 (N_8146,N_4209,N_1374);
xnor U8147 (N_8147,N_1908,N_4648);
or U8148 (N_8148,N_2947,N_4837);
nor U8149 (N_8149,N_3982,N_1161);
xor U8150 (N_8150,N_3596,N_1700);
xnor U8151 (N_8151,N_4870,N_1006);
xnor U8152 (N_8152,N_4572,N_3847);
or U8153 (N_8153,N_3331,N_4020);
nor U8154 (N_8154,N_279,N_4768);
xnor U8155 (N_8155,N_4704,N_3077);
or U8156 (N_8156,N_4376,N_3153);
nand U8157 (N_8157,N_2134,N_4927);
xnor U8158 (N_8158,N_4194,N_4937);
xnor U8159 (N_8159,N_2738,N_4539);
xor U8160 (N_8160,N_85,N_799);
and U8161 (N_8161,N_815,N_4253);
xor U8162 (N_8162,N_2388,N_3770);
xor U8163 (N_8163,N_3477,N_3691);
nor U8164 (N_8164,N_2873,N_1014);
nand U8165 (N_8165,N_2337,N_4887);
or U8166 (N_8166,N_2433,N_550);
nand U8167 (N_8167,N_3509,N_3818);
xor U8168 (N_8168,N_579,N_4037);
nor U8169 (N_8169,N_1619,N_1878);
and U8170 (N_8170,N_950,N_4848);
nand U8171 (N_8171,N_1513,N_4071);
or U8172 (N_8172,N_2887,N_3515);
nand U8173 (N_8173,N_517,N_145);
xor U8174 (N_8174,N_3142,N_1903);
or U8175 (N_8175,N_487,N_2492);
or U8176 (N_8176,N_181,N_1742);
or U8177 (N_8177,N_803,N_1378);
xor U8178 (N_8178,N_1707,N_602);
nand U8179 (N_8179,N_4492,N_2069);
and U8180 (N_8180,N_2747,N_4269);
and U8181 (N_8181,N_4404,N_4049);
nand U8182 (N_8182,N_3938,N_3316);
nor U8183 (N_8183,N_4289,N_4187);
or U8184 (N_8184,N_4085,N_724);
or U8185 (N_8185,N_2648,N_3571);
or U8186 (N_8186,N_945,N_1850);
nor U8187 (N_8187,N_3168,N_2055);
and U8188 (N_8188,N_4593,N_4749);
or U8189 (N_8189,N_3371,N_714);
xor U8190 (N_8190,N_1962,N_4994);
and U8191 (N_8191,N_4471,N_1157);
nand U8192 (N_8192,N_3564,N_4999);
nand U8193 (N_8193,N_4926,N_2323);
nand U8194 (N_8194,N_3365,N_1126);
or U8195 (N_8195,N_1013,N_553);
xnor U8196 (N_8196,N_1655,N_4884);
nand U8197 (N_8197,N_1601,N_1612);
nor U8198 (N_8198,N_556,N_4775);
nand U8199 (N_8199,N_2681,N_4646);
xor U8200 (N_8200,N_3279,N_4924);
xor U8201 (N_8201,N_2280,N_408);
xor U8202 (N_8202,N_4731,N_3123);
or U8203 (N_8203,N_405,N_1721);
nand U8204 (N_8204,N_2019,N_1401);
or U8205 (N_8205,N_3813,N_3186);
or U8206 (N_8206,N_2801,N_3076);
nand U8207 (N_8207,N_4795,N_3280);
nand U8208 (N_8208,N_1427,N_598);
and U8209 (N_8209,N_3837,N_1798);
or U8210 (N_8210,N_2658,N_3563);
nand U8211 (N_8211,N_4642,N_4233);
or U8212 (N_8212,N_1681,N_1758);
xnor U8213 (N_8213,N_279,N_3445);
nor U8214 (N_8214,N_3032,N_2701);
xnor U8215 (N_8215,N_468,N_1979);
xor U8216 (N_8216,N_2308,N_3048);
or U8217 (N_8217,N_2876,N_4104);
and U8218 (N_8218,N_3804,N_2215);
xnor U8219 (N_8219,N_3307,N_2660);
or U8220 (N_8220,N_1754,N_371);
nor U8221 (N_8221,N_4393,N_4059);
nor U8222 (N_8222,N_265,N_553);
and U8223 (N_8223,N_1580,N_666);
nor U8224 (N_8224,N_642,N_415);
xnor U8225 (N_8225,N_1911,N_4426);
nor U8226 (N_8226,N_4375,N_2373);
nand U8227 (N_8227,N_3345,N_4849);
nor U8228 (N_8228,N_2999,N_1127);
nand U8229 (N_8229,N_726,N_563);
or U8230 (N_8230,N_4122,N_2202);
nand U8231 (N_8231,N_320,N_4521);
nand U8232 (N_8232,N_2668,N_2426);
or U8233 (N_8233,N_4856,N_3924);
nor U8234 (N_8234,N_3601,N_2499);
nand U8235 (N_8235,N_3713,N_4142);
xor U8236 (N_8236,N_4340,N_600);
nand U8237 (N_8237,N_2464,N_747);
nand U8238 (N_8238,N_4175,N_799);
and U8239 (N_8239,N_436,N_2061);
nor U8240 (N_8240,N_3874,N_4030);
nand U8241 (N_8241,N_3250,N_4871);
and U8242 (N_8242,N_2198,N_2240);
xnor U8243 (N_8243,N_1603,N_1967);
or U8244 (N_8244,N_1203,N_4833);
nor U8245 (N_8245,N_4679,N_1006);
or U8246 (N_8246,N_2199,N_406);
xor U8247 (N_8247,N_264,N_4775);
or U8248 (N_8248,N_3927,N_1662);
nor U8249 (N_8249,N_2804,N_633);
xor U8250 (N_8250,N_877,N_4729);
nand U8251 (N_8251,N_1912,N_4951);
xor U8252 (N_8252,N_2506,N_3640);
and U8253 (N_8253,N_1269,N_4375);
or U8254 (N_8254,N_4669,N_1539);
and U8255 (N_8255,N_3259,N_893);
or U8256 (N_8256,N_3608,N_892);
or U8257 (N_8257,N_3823,N_2236);
xor U8258 (N_8258,N_1961,N_4339);
and U8259 (N_8259,N_1586,N_1340);
nand U8260 (N_8260,N_4149,N_4161);
nor U8261 (N_8261,N_143,N_4456);
nand U8262 (N_8262,N_2642,N_910);
and U8263 (N_8263,N_1642,N_2796);
xnor U8264 (N_8264,N_741,N_4529);
and U8265 (N_8265,N_1985,N_1465);
or U8266 (N_8266,N_2747,N_3551);
xor U8267 (N_8267,N_4301,N_261);
and U8268 (N_8268,N_2744,N_1753);
and U8269 (N_8269,N_1821,N_4995);
or U8270 (N_8270,N_3765,N_384);
nor U8271 (N_8271,N_3494,N_2402);
xor U8272 (N_8272,N_1818,N_3819);
and U8273 (N_8273,N_1744,N_2195);
nor U8274 (N_8274,N_2096,N_2520);
nor U8275 (N_8275,N_3934,N_1574);
and U8276 (N_8276,N_3157,N_1392);
or U8277 (N_8277,N_3598,N_3739);
and U8278 (N_8278,N_2305,N_2064);
nor U8279 (N_8279,N_4405,N_3828);
xor U8280 (N_8280,N_3738,N_1201);
nand U8281 (N_8281,N_183,N_4813);
xnor U8282 (N_8282,N_4633,N_1205);
nor U8283 (N_8283,N_905,N_2784);
xnor U8284 (N_8284,N_4748,N_3396);
nand U8285 (N_8285,N_490,N_1192);
and U8286 (N_8286,N_4004,N_71);
or U8287 (N_8287,N_808,N_2247);
nand U8288 (N_8288,N_4186,N_4281);
xnor U8289 (N_8289,N_4402,N_1577);
nor U8290 (N_8290,N_1951,N_1878);
xnor U8291 (N_8291,N_3376,N_1327);
nand U8292 (N_8292,N_4989,N_2581);
nand U8293 (N_8293,N_4160,N_2650);
and U8294 (N_8294,N_4481,N_1070);
nor U8295 (N_8295,N_34,N_2768);
and U8296 (N_8296,N_3872,N_3469);
xnor U8297 (N_8297,N_3694,N_3536);
xnor U8298 (N_8298,N_715,N_3139);
and U8299 (N_8299,N_2599,N_4204);
or U8300 (N_8300,N_4317,N_3267);
or U8301 (N_8301,N_445,N_1570);
and U8302 (N_8302,N_2331,N_3158);
or U8303 (N_8303,N_4964,N_3155);
xnor U8304 (N_8304,N_1300,N_4410);
or U8305 (N_8305,N_2184,N_4698);
nor U8306 (N_8306,N_4036,N_2524);
nand U8307 (N_8307,N_4572,N_2251);
nand U8308 (N_8308,N_1815,N_3779);
nand U8309 (N_8309,N_3416,N_3879);
xor U8310 (N_8310,N_1633,N_3223);
nor U8311 (N_8311,N_4946,N_2212);
or U8312 (N_8312,N_3428,N_1977);
and U8313 (N_8313,N_4580,N_4566);
nand U8314 (N_8314,N_3938,N_2594);
xor U8315 (N_8315,N_855,N_2699);
or U8316 (N_8316,N_4568,N_534);
nand U8317 (N_8317,N_4252,N_4305);
xnor U8318 (N_8318,N_4750,N_3162);
nor U8319 (N_8319,N_4861,N_1294);
or U8320 (N_8320,N_4843,N_1737);
nand U8321 (N_8321,N_3955,N_1800);
and U8322 (N_8322,N_4860,N_2809);
nor U8323 (N_8323,N_2180,N_1073);
nor U8324 (N_8324,N_198,N_2409);
nand U8325 (N_8325,N_2683,N_677);
and U8326 (N_8326,N_4103,N_634);
or U8327 (N_8327,N_543,N_213);
nor U8328 (N_8328,N_2749,N_2584);
and U8329 (N_8329,N_2947,N_4060);
nand U8330 (N_8330,N_1523,N_708);
or U8331 (N_8331,N_3597,N_4982);
or U8332 (N_8332,N_2192,N_1841);
and U8333 (N_8333,N_1871,N_4918);
nand U8334 (N_8334,N_4471,N_675);
or U8335 (N_8335,N_1285,N_1687);
nand U8336 (N_8336,N_3174,N_2875);
xor U8337 (N_8337,N_4489,N_200);
xor U8338 (N_8338,N_2899,N_3593);
nor U8339 (N_8339,N_15,N_4084);
nand U8340 (N_8340,N_2804,N_1163);
or U8341 (N_8341,N_3703,N_2061);
nor U8342 (N_8342,N_2487,N_1300);
nor U8343 (N_8343,N_4314,N_620);
or U8344 (N_8344,N_3009,N_2735);
nor U8345 (N_8345,N_365,N_2349);
xnor U8346 (N_8346,N_1511,N_4832);
xor U8347 (N_8347,N_2734,N_218);
xnor U8348 (N_8348,N_4560,N_2224);
and U8349 (N_8349,N_1392,N_1500);
nor U8350 (N_8350,N_4544,N_3175);
nor U8351 (N_8351,N_2915,N_4600);
xnor U8352 (N_8352,N_459,N_3953);
and U8353 (N_8353,N_4089,N_4983);
xnor U8354 (N_8354,N_1517,N_858);
nor U8355 (N_8355,N_3339,N_4315);
nor U8356 (N_8356,N_4990,N_3838);
nor U8357 (N_8357,N_1605,N_3792);
and U8358 (N_8358,N_3621,N_2425);
or U8359 (N_8359,N_4787,N_1587);
xor U8360 (N_8360,N_1346,N_531);
and U8361 (N_8361,N_4494,N_305);
or U8362 (N_8362,N_172,N_953);
xnor U8363 (N_8363,N_4885,N_1480);
xor U8364 (N_8364,N_588,N_4155);
and U8365 (N_8365,N_2161,N_3594);
nand U8366 (N_8366,N_4997,N_3123);
nand U8367 (N_8367,N_162,N_774);
nand U8368 (N_8368,N_4695,N_1832);
nor U8369 (N_8369,N_3613,N_3420);
nor U8370 (N_8370,N_4741,N_1019);
and U8371 (N_8371,N_3154,N_3322);
nand U8372 (N_8372,N_4912,N_2190);
or U8373 (N_8373,N_32,N_2493);
xor U8374 (N_8374,N_532,N_4157);
and U8375 (N_8375,N_3467,N_2502);
xor U8376 (N_8376,N_3593,N_1526);
xor U8377 (N_8377,N_1519,N_126);
nor U8378 (N_8378,N_2984,N_2018);
and U8379 (N_8379,N_2786,N_1456);
and U8380 (N_8380,N_4165,N_3560);
xnor U8381 (N_8381,N_2652,N_3452);
nand U8382 (N_8382,N_4454,N_2536);
xor U8383 (N_8383,N_1633,N_748);
and U8384 (N_8384,N_2365,N_3740);
nor U8385 (N_8385,N_4139,N_1466);
or U8386 (N_8386,N_4373,N_2511);
nand U8387 (N_8387,N_2315,N_1219);
or U8388 (N_8388,N_1524,N_1446);
and U8389 (N_8389,N_2100,N_1084);
xor U8390 (N_8390,N_2585,N_4249);
nor U8391 (N_8391,N_3825,N_4845);
xnor U8392 (N_8392,N_4023,N_1522);
nand U8393 (N_8393,N_4277,N_1843);
nand U8394 (N_8394,N_1841,N_149);
nand U8395 (N_8395,N_909,N_4471);
and U8396 (N_8396,N_2555,N_4549);
and U8397 (N_8397,N_1309,N_362);
nor U8398 (N_8398,N_2880,N_3363);
nor U8399 (N_8399,N_1645,N_1043);
xor U8400 (N_8400,N_2668,N_2473);
xor U8401 (N_8401,N_4202,N_4833);
and U8402 (N_8402,N_4497,N_4797);
xnor U8403 (N_8403,N_3184,N_1530);
nor U8404 (N_8404,N_2603,N_1272);
nand U8405 (N_8405,N_3057,N_4269);
nand U8406 (N_8406,N_4377,N_3197);
or U8407 (N_8407,N_2740,N_1016);
nand U8408 (N_8408,N_851,N_3240);
or U8409 (N_8409,N_4904,N_3765);
xor U8410 (N_8410,N_4900,N_4928);
nor U8411 (N_8411,N_2981,N_3161);
xnor U8412 (N_8412,N_1750,N_1825);
xor U8413 (N_8413,N_3142,N_4180);
or U8414 (N_8414,N_1466,N_1660);
nor U8415 (N_8415,N_1577,N_4448);
or U8416 (N_8416,N_1614,N_279);
nand U8417 (N_8417,N_1294,N_1585);
or U8418 (N_8418,N_4143,N_1804);
or U8419 (N_8419,N_641,N_897);
nand U8420 (N_8420,N_3285,N_3064);
or U8421 (N_8421,N_4974,N_623);
nand U8422 (N_8422,N_4907,N_636);
xor U8423 (N_8423,N_2843,N_4801);
and U8424 (N_8424,N_1096,N_68);
nor U8425 (N_8425,N_3123,N_1248);
nor U8426 (N_8426,N_2528,N_3136);
or U8427 (N_8427,N_3471,N_1981);
nor U8428 (N_8428,N_2461,N_2542);
or U8429 (N_8429,N_309,N_4202);
nor U8430 (N_8430,N_3941,N_1640);
and U8431 (N_8431,N_1803,N_2680);
nand U8432 (N_8432,N_2602,N_907);
xor U8433 (N_8433,N_4762,N_1654);
and U8434 (N_8434,N_1558,N_4499);
nor U8435 (N_8435,N_321,N_3897);
xnor U8436 (N_8436,N_3153,N_52);
and U8437 (N_8437,N_1878,N_3920);
nor U8438 (N_8438,N_3170,N_4144);
nor U8439 (N_8439,N_3353,N_1839);
xnor U8440 (N_8440,N_2864,N_3931);
nor U8441 (N_8441,N_2464,N_4555);
xor U8442 (N_8442,N_4742,N_3310);
nor U8443 (N_8443,N_2934,N_1731);
xnor U8444 (N_8444,N_871,N_2964);
and U8445 (N_8445,N_14,N_3142);
xor U8446 (N_8446,N_3318,N_51);
xor U8447 (N_8447,N_280,N_1607);
xnor U8448 (N_8448,N_4982,N_1803);
nor U8449 (N_8449,N_1012,N_1876);
nand U8450 (N_8450,N_4617,N_4515);
and U8451 (N_8451,N_4524,N_1523);
nand U8452 (N_8452,N_3226,N_3666);
nor U8453 (N_8453,N_3455,N_2733);
and U8454 (N_8454,N_1235,N_3208);
nand U8455 (N_8455,N_3410,N_2047);
nor U8456 (N_8456,N_1541,N_47);
nand U8457 (N_8457,N_2497,N_4027);
and U8458 (N_8458,N_294,N_3009);
nor U8459 (N_8459,N_3499,N_2246);
nor U8460 (N_8460,N_2881,N_1486);
or U8461 (N_8461,N_2735,N_2189);
and U8462 (N_8462,N_774,N_2817);
nand U8463 (N_8463,N_1865,N_792);
and U8464 (N_8464,N_1895,N_1801);
nor U8465 (N_8465,N_1399,N_2083);
and U8466 (N_8466,N_1241,N_2000);
nor U8467 (N_8467,N_4835,N_2652);
and U8468 (N_8468,N_1242,N_3079);
nor U8469 (N_8469,N_21,N_2882);
nor U8470 (N_8470,N_246,N_4863);
nor U8471 (N_8471,N_3891,N_2926);
nand U8472 (N_8472,N_1994,N_2115);
nor U8473 (N_8473,N_3872,N_4406);
nand U8474 (N_8474,N_4340,N_454);
and U8475 (N_8475,N_149,N_642);
or U8476 (N_8476,N_1405,N_4682);
xnor U8477 (N_8477,N_4460,N_4146);
nand U8478 (N_8478,N_2957,N_900);
nor U8479 (N_8479,N_1921,N_2800);
nor U8480 (N_8480,N_3958,N_4254);
and U8481 (N_8481,N_1772,N_2151);
nor U8482 (N_8482,N_3059,N_4796);
xor U8483 (N_8483,N_3565,N_4664);
nand U8484 (N_8484,N_950,N_3784);
or U8485 (N_8485,N_4841,N_3685);
xor U8486 (N_8486,N_3871,N_1066);
nor U8487 (N_8487,N_2215,N_1187);
nor U8488 (N_8488,N_3436,N_1059);
and U8489 (N_8489,N_439,N_1661);
or U8490 (N_8490,N_2889,N_1472);
and U8491 (N_8491,N_988,N_1758);
and U8492 (N_8492,N_3916,N_2312);
or U8493 (N_8493,N_3331,N_2385);
xnor U8494 (N_8494,N_2609,N_2196);
nand U8495 (N_8495,N_890,N_3949);
xnor U8496 (N_8496,N_4773,N_4137);
and U8497 (N_8497,N_1183,N_2194);
or U8498 (N_8498,N_4064,N_4262);
nand U8499 (N_8499,N_451,N_4891);
nand U8500 (N_8500,N_1234,N_1897);
nor U8501 (N_8501,N_1589,N_2312);
nand U8502 (N_8502,N_4683,N_4958);
nand U8503 (N_8503,N_239,N_2968);
nor U8504 (N_8504,N_1303,N_4610);
and U8505 (N_8505,N_151,N_3844);
xnor U8506 (N_8506,N_775,N_258);
and U8507 (N_8507,N_3805,N_956);
xnor U8508 (N_8508,N_1209,N_1527);
nand U8509 (N_8509,N_2883,N_1664);
xnor U8510 (N_8510,N_4715,N_1299);
and U8511 (N_8511,N_4641,N_2866);
and U8512 (N_8512,N_4208,N_4721);
nand U8513 (N_8513,N_3338,N_2661);
and U8514 (N_8514,N_4097,N_3043);
and U8515 (N_8515,N_2826,N_4028);
nand U8516 (N_8516,N_3934,N_954);
nor U8517 (N_8517,N_4145,N_1216);
and U8518 (N_8518,N_1975,N_2757);
nor U8519 (N_8519,N_4284,N_1375);
nor U8520 (N_8520,N_581,N_2674);
nand U8521 (N_8521,N_3140,N_934);
nor U8522 (N_8522,N_4946,N_4795);
nor U8523 (N_8523,N_1749,N_2264);
and U8524 (N_8524,N_3148,N_3711);
xor U8525 (N_8525,N_2823,N_501);
nor U8526 (N_8526,N_3681,N_1914);
xnor U8527 (N_8527,N_3150,N_849);
nor U8528 (N_8528,N_4126,N_3882);
xnor U8529 (N_8529,N_2239,N_4808);
or U8530 (N_8530,N_4987,N_2291);
nor U8531 (N_8531,N_1212,N_144);
and U8532 (N_8532,N_4869,N_838);
xor U8533 (N_8533,N_135,N_3904);
or U8534 (N_8534,N_670,N_1814);
or U8535 (N_8535,N_248,N_2763);
xnor U8536 (N_8536,N_3735,N_3653);
or U8537 (N_8537,N_2689,N_454);
or U8538 (N_8538,N_1271,N_4509);
nand U8539 (N_8539,N_2791,N_2376);
xnor U8540 (N_8540,N_1468,N_1971);
xnor U8541 (N_8541,N_879,N_385);
or U8542 (N_8542,N_4793,N_4268);
nor U8543 (N_8543,N_1879,N_3725);
nor U8544 (N_8544,N_280,N_4737);
and U8545 (N_8545,N_455,N_864);
xnor U8546 (N_8546,N_1637,N_4832);
xnor U8547 (N_8547,N_438,N_1982);
and U8548 (N_8548,N_83,N_1062);
and U8549 (N_8549,N_4920,N_2346);
nand U8550 (N_8550,N_4735,N_4715);
xnor U8551 (N_8551,N_4142,N_390);
and U8552 (N_8552,N_2351,N_593);
nor U8553 (N_8553,N_2692,N_963);
or U8554 (N_8554,N_2319,N_1683);
nand U8555 (N_8555,N_4656,N_668);
or U8556 (N_8556,N_3953,N_4134);
nand U8557 (N_8557,N_2197,N_3779);
and U8558 (N_8558,N_1181,N_4975);
or U8559 (N_8559,N_3152,N_2514);
and U8560 (N_8560,N_497,N_637);
xor U8561 (N_8561,N_2640,N_3049);
and U8562 (N_8562,N_3751,N_3772);
nand U8563 (N_8563,N_1473,N_576);
nand U8564 (N_8564,N_134,N_2789);
or U8565 (N_8565,N_278,N_3547);
and U8566 (N_8566,N_1372,N_2330);
nand U8567 (N_8567,N_4486,N_4975);
and U8568 (N_8568,N_145,N_4825);
xor U8569 (N_8569,N_2771,N_331);
xnor U8570 (N_8570,N_3491,N_4007);
and U8571 (N_8571,N_2338,N_2028);
or U8572 (N_8572,N_1506,N_3757);
xor U8573 (N_8573,N_2922,N_2748);
or U8574 (N_8574,N_2008,N_67);
nor U8575 (N_8575,N_1657,N_2817);
nor U8576 (N_8576,N_2677,N_4990);
nand U8577 (N_8577,N_4724,N_4886);
nor U8578 (N_8578,N_3417,N_2416);
nor U8579 (N_8579,N_1572,N_1185);
and U8580 (N_8580,N_4987,N_2112);
and U8581 (N_8581,N_3649,N_4486);
or U8582 (N_8582,N_472,N_3698);
and U8583 (N_8583,N_2513,N_1691);
nand U8584 (N_8584,N_392,N_1312);
nor U8585 (N_8585,N_2169,N_1711);
nor U8586 (N_8586,N_3140,N_2615);
xnor U8587 (N_8587,N_4806,N_53);
and U8588 (N_8588,N_1972,N_714);
nor U8589 (N_8589,N_3716,N_4906);
or U8590 (N_8590,N_133,N_338);
nand U8591 (N_8591,N_1267,N_1511);
and U8592 (N_8592,N_1811,N_466);
or U8593 (N_8593,N_4467,N_998);
nand U8594 (N_8594,N_2786,N_1275);
nand U8595 (N_8595,N_1267,N_1535);
nor U8596 (N_8596,N_826,N_1721);
nand U8597 (N_8597,N_2061,N_1864);
nand U8598 (N_8598,N_934,N_3428);
xor U8599 (N_8599,N_4931,N_3288);
nor U8600 (N_8600,N_4158,N_3950);
and U8601 (N_8601,N_4183,N_1762);
nand U8602 (N_8602,N_170,N_646);
nand U8603 (N_8603,N_4064,N_2818);
nor U8604 (N_8604,N_2436,N_4460);
nand U8605 (N_8605,N_2936,N_245);
or U8606 (N_8606,N_224,N_2896);
xnor U8607 (N_8607,N_3227,N_650);
or U8608 (N_8608,N_3899,N_753);
xor U8609 (N_8609,N_3185,N_4123);
xnor U8610 (N_8610,N_2190,N_3119);
nor U8611 (N_8611,N_1349,N_4464);
nor U8612 (N_8612,N_780,N_4843);
nand U8613 (N_8613,N_2539,N_3793);
nor U8614 (N_8614,N_908,N_2610);
xor U8615 (N_8615,N_2839,N_759);
or U8616 (N_8616,N_1410,N_650);
nand U8617 (N_8617,N_546,N_1066);
and U8618 (N_8618,N_396,N_2487);
nand U8619 (N_8619,N_1331,N_3015);
xnor U8620 (N_8620,N_3901,N_4082);
and U8621 (N_8621,N_1099,N_3078);
nor U8622 (N_8622,N_4312,N_2771);
and U8623 (N_8623,N_4190,N_185);
xor U8624 (N_8624,N_3788,N_3276);
and U8625 (N_8625,N_932,N_2803);
nor U8626 (N_8626,N_1252,N_3397);
and U8627 (N_8627,N_3038,N_2910);
nand U8628 (N_8628,N_1601,N_4116);
xnor U8629 (N_8629,N_2877,N_4982);
nor U8630 (N_8630,N_4196,N_2795);
and U8631 (N_8631,N_3394,N_1238);
nor U8632 (N_8632,N_3796,N_4304);
or U8633 (N_8633,N_2336,N_2973);
or U8634 (N_8634,N_210,N_4523);
xor U8635 (N_8635,N_1295,N_2769);
xnor U8636 (N_8636,N_4668,N_1670);
and U8637 (N_8637,N_4405,N_3575);
nor U8638 (N_8638,N_4126,N_3784);
or U8639 (N_8639,N_2192,N_2050);
or U8640 (N_8640,N_4259,N_4120);
and U8641 (N_8641,N_1986,N_993);
or U8642 (N_8642,N_600,N_2823);
and U8643 (N_8643,N_2299,N_2927);
nor U8644 (N_8644,N_1685,N_1546);
and U8645 (N_8645,N_3116,N_3552);
or U8646 (N_8646,N_3456,N_3974);
nor U8647 (N_8647,N_2726,N_1404);
or U8648 (N_8648,N_3401,N_2693);
xnor U8649 (N_8649,N_696,N_1700);
xnor U8650 (N_8650,N_3210,N_2350);
or U8651 (N_8651,N_4643,N_3211);
or U8652 (N_8652,N_243,N_776);
nand U8653 (N_8653,N_3285,N_4513);
nor U8654 (N_8654,N_4257,N_2946);
or U8655 (N_8655,N_1797,N_4114);
and U8656 (N_8656,N_4325,N_2430);
nor U8657 (N_8657,N_1962,N_3462);
nor U8658 (N_8658,N_2883,N_1584);
nand U8659 (N_8659,N_4061,N_2952);
nand U8660 (N_8660,N_3183,N_453);
nor U8661 (N_8661,N_4351,N_3735);
xor U8662 (N_8662,N_1128,N_2808);
xor U8663 (N_8663,N_3715,N_3318);
nor U8664 (N_8664,N_3324,N_1974);
xor U8665 (N_8665,N_220,N_3879);
xnor U8666 (N_8666,N_4913,N_132);
and U8667 (N_8667,N_4929,N_4937);
and U8668 (N_8668,N_4542,N_1920);
nand U8669 (N_8669,N_4078,N_4529);
nand U8670 (N_8670,N_3101,N_4530);
xor U8671 (N_8671,N_4940,N_4229);
xnor U8672 (N_8672,N_2904,N_3393);
or U8673 (N_8673,N_4776,N_1653);
xor U8674 (N_8674,N_1069,N_4955);
nor U8675 (N_8675,N_2981,N_4129);
nor U8676 (N_8676,N_3804,N_3654);
nor U8677 (N_8677,N_2636,N_4675);
and U8678 (N_8678,N_3365,N_4744);
nor U8679 (N_8679,N_610,N_1596);
and U8680 (N_8680,N_1685,N_3961);
nand U8681 (N_8681,N_3616,N_2057);
nand U8682 (N_8682,N_1750,N_2007);
nor U8683 (N_8683,N_4886,N_2803);
nand U8684 (N_8684,N_457,N_4805);
nand U8685 (N_8685,N_839,N_163);
nor U8686 (N_8686,N_1459,N_1025);
xnor U8687 (N_8687,N_2259,N_2823);
and U8688 (N_8688,N_3015,N_4382);
nor U8689 (N_8689,N_640,N_1549);
nor U8690 (N_8690,N_1047,N_1444);
or U8691 (N_8691,N_623,N_171);
nand U8692 (N_8692,N_3531,N_3523);
nor U8693 (N_8693,N_4011,N_2257);
xor U8694 (N_8694,N_4663,N_3088);
nor U8695 (N_8695,N_173,N_2047);
or U8696 (N_8696,N_1455,N_4720);
nor U8697 (N_8697,N_4890,N_4201);
or U8698 (N_8698,N_2072,N_796);
nor U8699 (N_8699,N_1585,N_1077);
and U8700 (N_8700,N_1248,N_4746);
xor U8701 (N_8701,N_1444,N_3832);
nor U8702 (N_8702,N_3259,N_1391);
xor U8703 (N_8703,N_2597,N_3652);
and U8704 (N_8704,N_4764,N_3816);
nor U8705 (N_8705,N_11,N_2960);
xnor U8706 (N_8706,N_4411,N_351);
or U8707 (N_8707,N_3943,N_3626);
and U8708 (N_8708,N_695,N_1881);
nor U8709 (N_8709,N_4204,N_1764);
xnor U8710 (N_8710,N_754,N_551);
or U8711 (N_8711,N_3478,N_2014);
nor U8712 (N_8712,N_3272,N_2814);
or U8713 (N_8713,N_4977,N_4219);
and U8714 (N_8714,N_4697,N_4965);
nand U8715 (N_8715,N_3506,N_410);
nand U8716 (N_8716,N_1797,N_1364);
xor U8717 (N_8717,N_2682,N_2150);
and U8718 (N_8718,N_3052,N_267);
nor U8719 (N_8719,N_4774,N_4165);
or U8720 (N_8720,N_269,N_2230);
nand U8721 (N_8721,N_3083,N_458);
nand U8722 (N_8722,N_1503,N_1039);
nand U8723 (N_8723,N_1864,N_706);
nor U8724 (N_8724,N_1759,N_4875);
nand U8725 (N_8725,N_2917,N_4900);
xnor U8726 (N_8726,N_2189,N_1745);
nand U8727 (N_8727,N_2741,N_2688);
xnor U8728 (N_8728,N_3755,N_2793);
and U8729 (N_8729,N_4895,N_883);
and U8730 (N_8730,N_989,N_4580);
xnor U8731 (N_8731,N_742,N_4707);
xnor U8732 (N_8732,N_3990,N_675);
xor U8733 (N_8733,N_3335,N_50);
nand U8734 (N_8734,N_1457,N_2865);
and U8735 (N_8735,N_1432,N_1917);
and U8736 (N_8736,N_3776,N_3644);
nor U8737 (N_8737,N_2826,N_3510);
nor U8738 (N_8738,N_3284,N_3191);
nand U8739 (N_8739,N_3515,N_862);
or U8740 (N_8740,N_1084,N_2201);
or U8741 (N_8741,N_540,N_3359);
nor U8742 (N_8742,N_43,N_4511);
nor U8743 (N_8743,N_2850,N_4217);
and U8744 (N_8744,N_1834,N_2111);
nand U8745 (N_8745,N_1169,N_4286);
and U8746 (N_8746,N_4124,N_268);
nor U8747 (N_8747,N_369,N_4645);
nor U8748 (N_8748,N_3415,N_3729);
or U8749 (N_8749,N_3861,N_4826);
xnor U8750 (N_8750,N_2573,N_791);
xor U8751 (N_8751,N_4807,N_703);
and U8752 (N_8752,N_1905,N_441);
or U8753 (N_8753,N_153,N_2175);
nand U8754 (N_8754,N_2972,N_3603);
and U8755 (N_8755,N_132,N_2118);
or U8756 (N_8756,N_996,N_266);
or U8757 (N_8757,N_1640,N_1043);
and U8758 (N_8758,N_2925,N_2555);
xor U8759 (N_8759,N_287,N_694);
xnor U8760 (N_8760,N_2654,N_988);
or U8761 (N_8761,N_2333,N_4719);
xor U8762 (N_8762,N_553,N_3301);
xor U8763 (N_8763,N_491,N_1820);
nand U8764 (N_8764,N_3238,N_3381);
and U8765 (N_8765,N_1375,N_1290);
nand U8766 (N_8766,N_2750,N_1194);
nor U8767 (N_8767,N_2174,N_3068);
xnor U8768 (N_8768,N_537,N_4542);
or U8769 (N_8769,N_1065,N_49);
nand U8770 (N_8770,N_1371,N_1165);
xnor U8771 (N_8771,N_2783,N_1655);
xnor U8772 (N_8772,N_3129,N_3487);
and U8773 (N_8773,N_4408,N_3995);
nand U8774 (N_8774,N_4924,N_716);
or U8775 (N_8775,N_2035,N_4829);
or U8776 (N_8776,N_1962,N_2398);
nor U8777 (N_8777,N_660,N_1470);
xnor U8778 (N_8778,N_3329,N_2112);
and U8779 (N_8779,N_4804,N_3740);
nand U8780 (N_8780,N_2150,N_3796);
nor U8781 (N_8781,N_3001,N_4574);
and U8782 (N_8782,N_2019,N_1703);
xor U8783 (N_8783,N_2702,N_2891);
xor U8784 (N_8784,N_2513,N_1599);
and U8785 (N_8785,N_1822,N_613);
and U8786 (N_8786,N_2686,N_4105);
or U8787 (N_8787,N_4338,N_751);
nor U8788 (N_8788,N_4438,N_1407);
xor U8789 (N_8789,N_2663,N_3092);
and U8790 (N_8790,N_2337,N_2236);
xor U8791 (N_8791,N_3308,N_3567);
and U8792 (N_8792,N_4916,N_1015);
xnor U8793 (N_8793,N_2818,N_1343);
and U8794 (N_8794,N_1723,N_154);
xor U8795 (N_8795,N_613,N_811);
xnor U8796 (N_8796,N_1769,N_1390);
nand U8797 (N_8797,N_3360,N_3661);
nand U8798 (N_8798,N_3430,N_2791);
or U8799 (N_8799,N_99,N_2388);
or U8800 (N_8800,N_719,N_4308);
xnor U8801 (N_8801,N_1754,N_1575);
and U8802 (N_8802,N_2425,N_1486);
or U8803 (N_8803,N_4845,N_871);
and U8804 (N_8804,N_2858,N_4084);
xnor U8805 (N_8805,N_113,N_3766);
xor U8806 (N_8806,N_658,N_4760);
and U8807 (N_8807,N_1872,N_797);
nor U8808 (N_8808,N_3579,N_4317);
and U8809 (N_8809,N_1828,N_1208);
or U8810 (N_8810,N_294,N_3701);
nor U8811 (N_8811,N_1043,N_4953);
and U8812 (N_8812,N_4337,N_3932);
and U8813 (N_8813,N_2653,N_2158);
nand U8814 (N_8814,N_4836,N_2054);
nand U8815 (N_8815,N_4302,N_273);
or U8816 (N_8816,N_4746,N_3033);
nor U8817 (N_8817,N_316,N_44);
or U8818 (N_8818,N_3748,N_1187);
and U8819 (N_8819,N_44,N_2606);
xnor U8820 (N_8820,N_2288,N_4046);
and U8821 (N_8821,N_206,N_595);
nand U8822 (N_8822,N_1940,N_2867);
nor U8823 (N_8823,N_3267,N_1104);
or U8824 (N_8824,N_769,N_4597);
and U8825 (N_8825,N_362,N_2704);
or U8826 (N_8826,N_1586,N_1277);
nand U8827 (N_8827,N_3286,N_2747);
and U8828 (N_8828,N_2533,N_2817);
or U8829 (N_8829,N_678,N_4652);
or U8830 (N_8830,N_1870,N_4114);
nand U8831 (N_8831,N_4383,N_4953);
nor U8832 (N_8832,N_1279,N_932);
and U8833 (N_8833,N_3726,N_2288);
nand U8834 (N_8834,N_2012,N_1959);
and U8835 (N_8835,N_2491,N_2375);
xor U8836 (N_8836,N_2212,N_4506);
or U8837 (N_8837,N_4832,N_3170);
xor U8838 (N_8838,N_2356,N_4059);
and U8839 (N_8839,N_4800,N_4201);
xor U8840 (N_8840,N_599,N_1728);
nand U8841 (N_8841,N_1694,N_3810);
nand U8842 (N_8842,N_2411,N_1023);
or U8843 (N_8843,N_2748,N_4699);
and U8844 (N_8844,N_960,N_4332);
xor U8845 (N_8845,N_3232,N_1329);
nand U8846 (N_8846,N_2585,N_2132);
nand U8847 (N_8847,N_4401,N_192);
nand U8848 (N_8848,N_3012,N_1412);
nor U8849 (N_8849,N_1461,N_658);
xor U8850 (N_8850,N_3984,N_4412);
nand U8851 (N_8851,N_2460,N_3914);
or U8852 (N_8852,N_232,N_3735);
nor U8853 (N_8853,N_4201,N_4631);
nand U8854 (N_8854,N_3618,N_3799);
xor U8855 (N_8855,N_3628,N_4530);
xor U8856 (N_8856,N_1665,N_3565);
or U8857 (N_8857,N_1823,N_2046);
nand U8858 (N_8858,N_1438,N_3631);
and U8859 (N_8859,N_1868,N_905);
or U8860 (N_8860,N_1711,N_3810);
or U8861 (N_8861,N_2879,N_167);
nand U8862 (N_8862,N_4113,N_4474);
and U8863 (N_8863,N_432,N_4391);
nor U8864 (N_8864,N_3064,N_157);
xnor U8865 (N_8865,N_3586,N_2425);
nor U8866 (N_8866,N_3296,N_1568);
or U8867 (N_8867,N_1181,N_3581);
or U8868 (N_8868,N_593,N_1264);
and U8869 (N_8869,N_357,N_2729);
nand U8870 (N_8870,N_4831,N_598);
nand U8871 (N_8871,N_251,N_1195);
nand U8872 (N_8872,N_1214,N_3177);
or U8873 (N_8873,N_1912,N_4753);
and U8874 (N_8874,N_2756,N_2216);
or U8875 (N_8875,N_655,N_4477);
or U8876 (N_8876,N_227,N_2976);
nor U8877 (N_8877,N_1625,N_3916);
nand U8878 (N_8878,N_3349,N_4995);
nand U8879 (N_8879,N_44,N_911);
nor U8880 (N_8880,N_3164,N_2256);
nand U8881 (N_8881,N_2991,N_85);
or U8882 (N_8882,N_1621,N_3810);
nor U8883 (N_8883,N_2814,N_2545);
nor U8884 (N_8884,N_2837,N_3483);
xor U8885 (N_8885,N_3300,N_274);
nand U8886 (N_8886,N_4283,N_542);
nor U8887 (N_8887,N_1754,N_2894);
nand U8888 (N_8888,N_280,N_2752);
xnor U8889 (N_8889,N_640,N_911);
or U8890 (N_8890,N_2400,N_4698);
nor U8891 (N_8891,N_915,N_2575);
or U8892 (N_8892,N_2985,N_3203);
and U8893 (N_8893,N_4698,N_587);
nor U8894 (N_8894,N_4517,N_1600);
or U8895 (N_8895,N_2239,N_1375);
nand U8896 (N_8896,N_522,N_4139);
nand U8897 (N_8897,N_1929,N_2817);
and U8898 (N_8898,N_4694,N_1909);
or U8899 (N_8899,N_2681,N_4736);
or U8900 (N_8900,N_621,N_248);
and U8901 (N_8901,N_837,N_2643);
xnor U8902 (N_8902,N_2770,N_2358);
nand U8903 (N_8903,N_4605,N_4097);
nor U8904 (N_8904,N_1870,N_3012);
nand U8905 (N_8905,N_4865,N_639);
nor U8906 (N_8906,N_1310,N_2579);
xnor U8907 (N_8907,N_2484,N_3107);
or U8908 (N_8908,N_3018,N_4870);
nor U8909 (N_8909,N_761,N_1059);
and U8910 (N_8910,N_1874,N_1138);
xor U8911 (N_8911,N_617,N_25);
and U8912 (N_8912,N_2318,N_259);
xnor U8913 (N_8913,N_2107,N_2468);
xnor U8914 (N_8914,N_1431,N_4921);
xor U8915 (N_8915,N_608,N_2566);
and U8916 (N_8916,N_1799,N_2212);
and U8917 (N_8917,N_1330,N_2880);
xor U8918 (N_8918,N_1934,N_1884);
nand U8919 (N_8919,N_3351,N_275);
or U8920 (N_8920,N_1426,N_814);
and U8921 (N_8921,N_824,N_1738);
nand U8922 (N_8922,N_3681,N_46);
nand U8923 (N_8923,N_987,N_1467);
nor U8924 (N_8924,N_1599,N_2106);
nor U8925 (N_8925,N_3547,N_4423);
xor U8926 (N_8926,N_1015,N_3921);
xor U8927 (N_8927,N_1129,N_3428);
xor U8928 (N_8928,N_3985,N_1481);
nand U8929 (N_8929,N_4829,N_3090);
and U8930 (N_8930,N_3664,N_38);
or U8931 (N_8931,N_3070,N_3564);
nor U8932 (N_8932,N_3881,N_2715);
or U8933 (N_8933,N_4891,N_3172);
xor U8934 (N_8934,N_918,N_4847);
and U8935 (N_8935,N_2947,N_2063);
xnor U8936 (N_8936,N_885,N_3803);
nor U8937 (N_8937,N_3725,N_4808);
and U8938 (N_8938,N_4664,N_255);
or U8939 (N_8939,N_4574,N_581);
nor U8940 (N_8940,N_1587,N_4509);
and U8941 (N_8941,N_3950,N_1613);
xnor U8942 (N_8942,N_2751,N_4034);
nand U8943 (N_8943,N_3204,N_2046);
xor U8944 (N_8944,N_4310,N_2821);
or U8945 (N_8945,N_2031,N_1910);
nand U8946 (N_8946,N_3151,N_82);
nor U8947 (N_8947,N_3637,N_2511);
and U8948 (N_8948,N_630,N_4760);
xor U8949 (N_8949,N_211,N_4366);
or U8950 (N_8950,N_1854,N_4389);
or U8951 (N_8951,N_3492,N_3556);
or U8952 (N_8952,N_4618,N_1400);
and U8953 (N_8953,N_287,N_4677);
xnor U8954 (N_8954,N_2446,N_3250);
nand U8955 (N_8955,N_629,N_3855);
nor U8956 (N_8956,N_2503,N_3230);
nor U8957 (N_8957,N_4296,N_775);
xnor U8958 (N_8958,N_4509,N_1109);
or U8959 (N_8959,N_8,N_15);
nor U8960 (N_8960,N_3219,N_1745);
nor U8961 (N_8961,N_4989,N_3510);
xnor U8962 (N_8962,N_2166,N_1745);
nor U8963 (N_8963,N_415,N_1610);
nor U8964 (N_8964,N_3063,N_4021);
nand U8965 (N_8965,N_3349,N_281);
xnor U8966 (N_8966,N_583,N_1403);
nor U8967 (N_8967,N_850,N_1728);
nor U8968 (N_8968,N_4808,N_3088);
and U8969 (N_8969,N_1408,N_243);
or U8970 (N_8970,N_2279,N_1895);
and U8971 (N_8971,N_4694,N_3819);
xnor U8972 (N_8972,N_496,N_781);
and U8973 (N_8973,N_2928,N_2056);
nand U8974 (N_8974,N_1364,N_2123);
or U8975 (N_8975,N_92,N_1108);
and U8976 (N_8976,N_4392,N_2226);
or U8977 (N_8977,N_3048,N_4872);
nand U8978 (N_8978,N_790,N_4131);
and U8979 (N_8979,N_1292,N_4372);
xnor U8980 (N_8980,N_1909,N_3631);
nor U8981 (N_8981,N_4934,N_2931);
or U8982 (N_8982,N_770,N_3800);
nand U8983 (N_8983,N_4182,N_1328);
nand U8984 (N_8984,N_3176,N_4215);
or U8985 (N_8985,N_1977,N_1824);
nor U8986 (N_8986,N_1584,N_2387);
and U8987 (N_8987,N_824,N_200);
xor U8988 (N_8988,N_4547,N_3666);
xor U8989 (N_8989,N_1005,N_1732);
and U8990 (N_8990,N_3315,N_2073);
nand U8991 (N_8991,N_3276,N_1621);
nand U8992 (N_8992,N_4921,N_133);
xnor U8993 (N_8993,N_2989,N_3164);
xnor U8994 (N_8994,N_1518,N_1425);
or U8995 (N_8995,N_885,N_25);
and U8996 (N_8996,N_4850,N_898);
nand U8997 (N_8997,N_2774,N_1985);
xor U8998 (N_8998,N_4613,N_3286);
nor U8999 (N_8999,N_4562,N_361);
xor U9000 (N_9000,N_873,N_3384);
nand U9001 (N_9001,N_794,N_200);
or U9002 (N_9002,N_3911,N_3994);
xnor U9003 (N_9003,N_4549,N_1415);
xnor U9004 (N_9004,N_4356,N_3079);
or U9005 (N_9005,N_357,N_3330);
nor U9006 (N_9006,N_2249,N_4355);
nand U9007 (N_9007,N_372,N_418);
nor U9008 (N_9008,N_275,N_1218);
or U9009 (N_9009,N_4657,N_4690);
nor U9010 (N_9010,N_4884,N_4510);
nor U9011 (N_9011,N_3973,N_4658);
xor U9012 (N_9012,N_4141,N_1419);
nand U9013 (N_9013,N_3292,N_4290);
xnor U9014 (N_9014,N_3082,N_2913);
xnor U9015 (N_9015,N_3491,N_1571);
xor U9016 (N_9016,N_3764,N_2689);
and U9017 (N_9017,N_1025,N_1552);
xor U9018 (N_9018,N_4067,N_2025);
nand U9019 (N_9019,N_3047,N_3894);
and U9020 (N_9020,N_1804,N_4340);
xor U9021 (N_9021,N_2576,N_4825);
and U9022 (N_9022,N_3559,N_3119);
nand U9023 (N_9023,N_4155,N_4016);
or U9024 (N_9024,N_2526,N_4660);
or U9025 (N_9025,N_1618,N_1934);
and U9026 (N_9026,N_929,N_4903);
nand U9027 (N_9027,N_2640,N_3601);
and U9028 (N_9028,N_4773,N_1967);
nor U9029 (N_9029,N_949,N_3931);
xnor U9030 (N_9030,N_701,N_4466);
nand U9031 (N_9031,N_4578,N_670);
and U9032 (N_9032,N_1118,N_4160);
and U9033 (N_9033,N_1169,N_2459);
xor U9034 (N_9034,N_47,N_3520);
nor U9035 (N_9035,N_3692,N_3387);
or U9036 (N_9036,N_4790,N_68);
and U9037 (N_9037,N_2962,N_2742);
nor U9038 (N_9038,N_2291,N_3404);
nor U9039 (N_9039,N_3541,N_1345);
and U9040 (N_9040,N_3928,N_3891);
or U9041 (N_9041,N_4059,N_4222);
nor U9042 (N_9042,N_4352,N_1792);
nand U9043 (N_9043,N_2337,N_2424);
and U9044 (N_9044,N_3015,N_1701);
nor U9045 (N_9045,N_59,N_1271);
nor U9046 (N_9046,N_1571,N_3250);
nor U9047 (N_9047,N_4206,N_4144);
and U9048 (N_9048,N_388,N_4914);
nand U9049 (N_9049,N_2069,N_2814);
and U9050 (N_9050,N_1680,N_4835);
nand U9051 (N_9051,N_4823,N_1265);
nor U9052 (N_9052,N_4174,N_2525);
and U9053 (N_9053,N_1609,N_619);
and U9054 (N_9054,N_1655,N_920);
nor U9055 (N_9055,N_4654,N_4247);
nand U9056 (N_9056,N_2015,N_304);
and U9057 (N_9057,N_3313,N_2285);
xnor U9058 (N_9058,N_847,N_2695);
xor U9059 (N_9059,N_4461,N_3691);
or U9060 (N_9060,N_3112,N_3855);
nand U9061 (N_9061,N_457,N_2731);
nand U9062 (N_9062,N_1067,N_4843);
xnor U9063 (N_9063,N_3559,N_784);
nand U9064 (N_9064,N_4708,N_919);
and U9065 (N_9065,N_526,N_1014);
xnor U9066 (N_9066,N_2545,N_368);
and U9067 (N_9067,N_4343,N_1087);
and U9068 (N_9068,N_3581,N_2125);
or U9069 (N_9069,N_2761,N_3553);
nor U9070 (N_9070,N_3541,N_3319);
nor U9071 (N_9071,N_440,N_1222);
nand U9072 (N_9072,N_707,N_4754);
nand U9073 (N_9073,N_2393,N_593);
nand U9074 (N_9074,N_949,N_249);
nand U9075 (N_9075,N_3655,N_4555);
or U9076 (N_9076,N_449,N_4644);
and U9077 (N_9077,N_4088,N_4511);
and U9078 (N_9078,N_2777,N_2209);
and U9079 (N_9079,N_217,N_4430);
and U9080 (N_9080,N_1267,N_4746);
nor U9081 (N_9081,N_4171,N_3418);
xnor U9082 (N_9082,N_3784,N_4741);
and U9083 (N_9083,N_2067,N_2900);
or U9084 (N_9084,N_2606,N_2011);
and U9085 (N_9085,N_500,N_1848);
nand U9086 (N_9086,N_723,N_919);
and U9087 (N_9087,N_4303,N_360);
xor U9088 (N_9088,N_28,N_1725);
xor U9089 (N_9089,N_194,N_3111);
nor U9090 (N_9090,N_2267,N_1043);
nand U9091 (N_9091,N_1713,N_135);
xnor U9092 (N_9092,N_4072,N_1592);
nand U9093 (N_9093,N_4159,N_4780);
nor U9094 (N_9094,N_2084,N_1608);
nand U9095 (N_9095,N_1642,N_1424);
nand U9096 (N_9096,N_2867,N_907);
and U9097 (N_9097,N_3022,N_561);
or U9098 (N_9098,N_2514,N_3654);
nand U9099 (N_9099,N_401,N_2880);
nand U9100 (N_9100,N_1355,N_4754);
nand U9101 (N_9101,N_244,N_3890);
and U9102 (N_9102,N_1440,N_1752);
xor U9103 (N_9103,N_4876,N_1538);
or U9104 (N_9104,N_1471,N_3977);
xnor U9105 (N_9105,N_2632,N_467);
xor U9106 (N_9106,N_2976,N_3447);
nor U9107 (N_9107,N_600,N_1829);
nor U9108 (N_9108,N_1896,N_3524);
or U9109 (N_9109,N_2240,N_367);
nand U9110 (N_9110,N_3101,N_2548);
nor U9111 (N_9111,N_1858,N_3306);
nor U9112 (N_9112,N_3364,N_2866);
or U9113 (N_9113,N_3696,N_3313);
nor U9114 (N_9114,N_1551,N_3927);
nand U9115 (N_9115,N_3941,N_2730);
xor U9116 (N_9116,N_1430,N_2551);
nand U9117 (N_9117,N_1515,N_3191);
nor U9118 (N_9118,N_1403,N_109);
xor U9119 (N_9119,N_3927,N_380);
or U9120 (N_9120,N_4187,N_2744);
nand U9121 (N_9121,N_2400,N_3019);
nor U9122 (N_9122,N_342,N_2880);
nor U9123 (N_9123,N_2871,N_4034);
or U9124 (N_9124,N_4148,N_622);
nand U9125 (N_9125,N_4122,N_2042);
nand U9126 (N_9126,N_698,N_424);
nor U9127 (N_9127,N_218,N_2650);
xor U9128 (N_9128,N_4505,N_2975);
nor U9129 (N_9129,N_3810,N_1237);
nor U9130 (N_9130,N_4881,N_376);
nand U9131 (N_9131,N_46,N_2354);
nor U9132 (N_9132,N_1185,N_2633);
nor U9133 (N_9133,N_4958,N_31);
nand U9134 (N_9134,N_36,N_2178);
or U9135 (N_9135,N_2409,N_1334);
xor U9136 (N_9136,N_1708,N_1967);
nand U9137 (N_9137,N_2507,N_4408);
and U9138 (N_9138,N_1568,N_2864);
and U9139 (N_9139,N_3811,N_2601);
xnor U9140 (N_9140,N_279,N_4836);
and U9141 (N_9141,N_3944,N_4101);
nor U9142 (N_9142,N_2313,N_550);
nand U9143 (N_9143,N_4526,N_4824);
xor U9144 (N_9144,N_1745,N_4632);
or U9145 (N_9145,N_2093,N_4622);
and U9146 (N_9146,N_75,N_4963);
xor U9147 (N_9147,N_989,N_182);
and U9148 (N_9148,N_3249,N_947);
or U9149 (N_9149,N_2694,N_3144);
or U9150 (N_9150,N_4847,N_4965);
and U9151 (N_9151,N_4243,N_583);
xnor U9152 (N_9152,N_2136,N_828);
nor U9153 (N_9153,N_4659,N_3874);
and U9154 (N_9154,N_295,N_4313);
or U9155 (N_9155,N_266,N_2633);
xnor U9156 (N_9156,N_2386,N_1334);
nand U9157 (N_9157,N_2595,N_3407);
nor U9158 (N_9158,N_3630,N_2398);
nand U9159 (N_9159,N_358,N_4388);
nor U9160 (N_9160,N_681,N_947);
or U9161 (N_9161,N_4517,N_4364);
xnor U9162 (N_9162,N_780,N_4660);
nand U9163 (N_9163,N_611,N_2217);
nand U9164 (N_9164,N_1697,N_3885);
xor U9165 (N_9165,N_4956,N_2305);
or U9166 (N_9166,N_103,N_766);
or U9167 (N_9167,N_3783,N_2642);
or U9168 (N_9168,N_3542,N_1866);
nor U9169 (N_9169,N_1243,N_4981);
or U9170 (N_9170,N_1129,N_3215);
nand U9171 (N_9171,N_3512,N_755);
nor U9172 (N_9172,N_2171,N_3695);
xor U9173 (N_9173,N_3808,N_4694);
or U9174 (N_9174,N_736,N_3725);
or U9175 (N_9175,N_123,N_2839);
xor U9176 (N_9176,N_650,N_118);
nand U9177 (N_9177,N_2706,N_1897);
or U9178 (N_9178,N_1552,N_411);
and U9179 (N_9179,N_734,N_4517);
nand U9180 (N_9180,N_2399,N_2223);
nand U9181 (N_9181,N_4153,N_4746);
and U9182 (N_9182,N_3227,N_4046);
and U9183 (N_9183,N_4676,N_1925);
xor U9184 (N_9184,N_451,N_2058);
nand U9185 (N_9185,N_1403,N_3113);
and U9186 (N_9186,N_3207,N_4657);
nor U9187 (N_9187,N_2014,N_1726);
and U9188 (N_9188,N_4712,N_3277);
xnor U9189 (N_9189,N_4084,N_2676);
and U9190 (N_9190,N_2664,N_4309);
nand U9191 (N_9191,N_840,N_1322);
or U9192 (N_9192,N_2428,N_3969);
xnor U9193 (N_9193,N_897,N_1990);
nand U9194 (N_9194,N_2997,N_3045);
xor U9195 (N_9195,N_3761,N_3529);
or U9196 (N_9196,N_4523,N_3485);
nand U9197 (N_9197,N_3263,N_2400);
nor U9198 (N_9198,N_4930,N_1723);
xor U9199 (N_9199,N_1860,N_3);
and U9200 (N_9200,N_1486,N_3883);
nor U9201 (N_9201,N_3947,N_1046);
or U9202 (N_9202,N_1007,N_1256);
and U9203 (N_9203,N_1484,N_2894);
nor U9204 (N_9204,N_1881,N_1089);
and U9205 (N_9205,N_1046,N_1390);
and U9206 (N_9206,N_4317,N_134);
nor U9207 (N_9207,N_3017,N_3543);
xnor U9208 (N_9208,N_1280,N_2787);
xor U9209 (N_9209,N_4869,N_81);
and U9210 (N_9210,N_3123,N_3499);
xnor U9211 (N_9211,N_25,N_1858);
xor U9212 (N_9212,N_2394,N_2144);
xor U9213 (N_9213,N_1084,N_2082);
and U9214 (N_9214,N_4665,N_2598);
or U9215 (N_9215,N_3441,N_2376);
xor U9216 (N_9216,N_3343,N_3365);
nor U9217 (N_9217,N_1137,N_4321);
nor U9218 (N_9218,N_1241,N_1056);
and U9219 (N_9219,N_956,N_1672);
nand U9220 (N_9220,N_1305,N_3342);
nand U9221 (N_9221,N_3990,N_3168);
and U9222 (N_9222,N_1502,N_479);
and U9223 (N_9223,N_4730,N_119);
xnor U9224 (N_9224,N_1664,N_4293);
or U9225 (N_9225,N_1260,N_801);
and U9226 (N_9226,N_3960,N_4633);
or U9227 (N_9227,N_3798,N_1281);
and U9228 (N_9228,N_297,N_1934);
xor U9229 (N_9229,N_4051,N_14);
xnor U9230 (N_9230,N_4312,N_3056);
or U9231 (N_9231,N_826,N_1056);
xnor U9232 (N_9232,N_1637,N_1284);
nor U9233 (N_9233,N_1305,N_4959);
and U9234 (N_9234,N_3027,N_4586);
and U9235 (N_9235,N_1314,N_2832);
nand U9236 (N_9236,N_1905,N_2532);
and U9237 (N_9237,N_2553,N_3057);
or U9238 (N_9238,N_3054,N_1953);
xnor U9239 (N_9239,N_3672,N_4387);
nor U9240 (N_9240,N_1324,N_2792);
or U9241 (N_9241,N_2090,N_2003);
or U9242 (N_9242,N_3080,N_3470);
and U9243 (N_9243,N_4983,N_1509);
xnor U9244 (N_9244,N_856,N_4896);
xor U9245 (N_9245,N_2300,N_2987);
or U9246 (N_9246,N_1491,N_1960);
and U9247 (N_9247,N_874,N_2001);
or U9248 (N_9248,N_453,N_3137);
nand U9249 (N_9249,N_3419,N_819);
nand U9250 (N_9250,N_357,N_3792);
nor U9251 (N_9251,N_1940,N_4766);
xnor U9252 (N_9252,N_4578,N_3420);
nand U9253 (N_9253,N_4102,N_3390);
nor U9254 (N_9254,N_17,N_1977);
or U9255 (N_9255,N_1719,N_915);
nor U9256 (N_9256,N_2818,N_1319);
nand U9257 (N_9257,N_775,N_3979);
or U9258 (N_9258,N_937,N_3479);
xnor U9259 (N_9259,N_273,N_2116);
nor U9260 (N_9260,N_978,N_563);
nor U9261 (N_9261,N_565,N_1551);
and U9262 (N_9262,N_3501,N_870);
or U9263 (N_9263,N_2524,N_4723);
and U9264 (N_9264,N_1867,N_1996);
xnor U9265 (N_9265,N_1450,N_3133);
nor U9266 (N_9266,N_1995,N_3011);
nor U9267 (N_9267,N_1498,N_3031);
and U9268 (N_9268,N_505,N_3920);
nand U9269 (N_9269,N_1445,N_3782);
nand U9270 (N_9270,N_1443,N_4180);
nand U9271 (N_9271,N_103,N_1114);
nand U9272 (N_9272,N_4422,N_1227);
or U9273 (N_9273,N_285,N_99);
xor U9274 (N_9274,N_2613,N_1299);
nor U9275 (N_9275,N_720,N_4484);
xnor U9276 (N_9276,N_4022,N_4226);
nand U9277 (N_9277,N_386,N_2130);
and U9278 (N_9278,N_3286,N_4520);
or U9279 (N_9279,N_3405,N_4064);
nand U9280 (N_9280,N_416,N_4282);
xor U9281 (N_9281,N_2925,N_109);
and U9282 (N_9282,N_4284,N_1340);
nand U9283 (N_9283,N_1703,N_3408);
nand U9284 (N_9284,N_3797,N_19);
nand U9285 (N_9285,N_147,N_3473);
nand U9286 (N_9286,N_643,N_2123);
nand U9287 (N_9287,N_4605,N_175);
or U9288 (N_9288,N_850,N_4489);
or U9289 (N_9289,N_1121,N_2128);
or U9290 (N_9290,N_3627,N_2299);
and U9291 (N_9291,N_4394,N_1703);
nor U9292 (N_9292,N_4814,N_4134);
and U9293 (N_9293,N_3111,N_549);
or U9294 (N_9294,N_1153,N_2849);
or U9295 (N_9295,N_2467,N_4510);
and U9296 (N_9296,N_4985,N_1730);
or U9297 (N_9297,N_429,N_300);
xnor U9298 (N_9298,N_3147,N_1549);
and U9299 (N_9299,N_2664,N_3343);
nand U9300 (N_9300,N_643,N_2991);
and U9301 (N_9301,N_3360,N_4265);
xnor U9302 (N_9302,N_3336,N_3694);
or U9303 (N_9303,N_3006,N_2184);
or U9304 (N_9304,N_4832,N_496);
and U9305 (N_9305,N_1523,N_4424);
nand U9306 (N_9306,N_2320,N_4965);
and U9307 (N_9307,N_1318,N_2206);
nand U9308 (N_9308,N_1202,N_1102);
nand U9309 (N_9309,N_3502,N_3489);
and U9310 (N_9310,N_2017,N_4632);
and U9311 (N_9311,N_4056,N_523);
and U9312 (N_9312,N_4673,N_1650);
and U9313 (N_9313,N_2453,N_3850);
nand U9314 (N_9314,N_4416,N_2150);
xor U9315 (N_9315,N_3944,N_4058);
xnor U9316 (N_9316,N_3780,N_1930);
and U9317 (N_9317,N_1060,N_907);
xnor U9318 (N_9318,N_1225,N_185);
xor U9319 (N_9319,N_4536,N_4901);
nor U9320 (N_9320,N_3204,N_1436);
xor U9321 (N_9321,N_4307,N_2174);
xor U9322 (N_9322,N_2761,N_4054);
xor U9323 (N_9323,N_1533,N_1858);
nor U9324 (N_9324,N_4436,N_280);
or U9325 (N_9325,N_4978,N_4519);
or U9326 (N_9326,N_4511,N_195);
xor U9327 (N_9327,N_2719,N_801);
nor U9328 (N_9328,N_880,N_2835);
or U9329 (N_9329,N_4314,N_632);
xnor U9330 (N_9330,N_3435,N_2982);
nand U9331 (N_9331,N_4431,N_3165);
nor U9332 (N_9332,N_4578,N_1194);
xnor U9333 (N_9333,N_3927,N_932);
xor U9334 (N_9334,N_3942,N_1251);
and U9335 (N_9335,N_784,N_1623);
xnor U9336 (N_9336,N_1363,N_1741);
nor U9337 (N_9337,N_309,N_1791);
and U9338 (N_9338,N_1419,N_3264);
xor U9339 (N_9339,N_1702,N_4377);
nand U9340 (N_9340,N_4235,N_105);
nand U9341 (N_9341,N_3236,N_270);
nor U9342 (N_9342,N_2680,N_4669);
nor U9343 (N_9343,N_2926,N_3183);
xor U9344 (N_9344,N_338,N_4840);
xnor U9345 (N_9345,N_1665,N_2642);
xnor U9346 (N_9346,N_3002,N_1875);
or U9347 (N_9347,N_4970,N_4374);
nor U9348 (N_9348,N_2097,N_54);
nor U9349 (N_9349,N_3412,N_4804);
xor U9350 (N_9350,N_8,N_4832);
nor U9351 (N_9351,N_3510,N_4136);
and U9352 (N_9352,N_1332,N_2021);
and U9353 (N_9353,N_2531,N_3157);
or U9354 (N_9354,N_2612,N_3919);
or U9355 (N_9355,N_637,N_3686);
or U9356 (N_9356,N_985,N_3886);
and U9357 (N_9357,N_257,N_2123);
xnor U9358 (N_9358,N_4810,N_3080);
nand U9359 (N_9359,N_3803,N_3993);
or U9360 (N_9360,N_2407,N_2209);
nand U9361 (N_9361,N_4405,N_489);
or U9362 (N_9362,N_4630,N_3227);
nor U9363 (N_9363,N_3535,N_3029);
or U9364 (N_9364,N_1709,N_1706);
nand U9365 (N_9365,N_579,N_3059);
and U9366 (N_9366,N_2742,N_4420);
xor U9367 (N_9367,N_994,N_3282);
nor U9368 (N_9368,N_77,N_585);
or U9369 (N_9369,N_1483,N_2351);
and U9370 (N_9370,N_4386,N_4438);
and U9371 (N_9371,N_109,N_4092);
nor U9372 (N_9372,N_1217,N_746);
and U9373 (N_9373,N_4606,N_4010);
or U9374 (N_9374,N_2248,N_4481);
or U9375 (N_9375,N_301,N_3180);
nand U9376 (N_9376,N_3034,N_2379);
nor U9377 (N_9377,N_3412,N_1147);
nand U9378 (N_9378,N_1106,N_1915);
nand U9379 (N_9379,N_1277,N_3702);
or U9380 (N_9380,N_4994,N_3487);
and U9381 (N_9381,N_2400,N_4776);
xnor U9382 (N_9382,N_425,N_1934);
nand U9383 (N_9383,N_763,N_1859);
or U9384 (N_9384,N_2888,N_3304);
and U9385 (N_9385,N_4600,N_4640);
or U9386 (N_9386,N_1695,N_2286);
and U9387 (N_9387,N_794,N_3874);
and U9388 (N_9388,N_4806,N_3804);
or U9389 (N_9389,N_1089,N_801);
xnor U9390 (N_9390,N_3183,N_110);
nor U9391 (N_9391,N_4612,N_1760);
nand U9392 (N_9392,N_4689,N_2772);
xor U9393 (N_9393,N_1333,N_4937);
xnor U9394 (N_9394,N_54,N_3003);
and U9395 (N_9395,N_4088,N_2523);
and U9396 (N_9396,N_4908,N_2533);
xnor U9397 (N_9397,N_1504,N_2785);
nor U9398 (N_9398,N_4729,N_3621);
xnor U9399 (N_9399,N_2897,N_3460);
xor U9400 (N_9400,N_2632,N_2771);
and U9401 (N_9401,N_2266,N_2458);
and U9402 (N_9402,N_4817,N_603);
nor U9403 (N_9403,N_3147,N_3040);
or U9404 (N_9404,N_391,N_4682);
nor U9405 (N_9405,N_1784,N_2628);
and U9406 (N_9406,N_1095,N_509);
and U9407 (N_9407,N_4568,N_3648);
nand U9408 (N_9408,N_2058,N_340);
and U9409 (N_9409,N_4889,N_2240);
or U9410 (N_9410,N_1036,N_600);
nor U9411 (N_9411,N_1865,N_1417);
nand U9412 (N_9412,N_3177,N_594);
nand U9413 (N_9413,N_3302,N_1659);
nand U9414 (N_9414,N_4479,N_1122);
or U9415 (N_9415,N_1080,N_3894);
nand U9416 (N_9416,N_3778,N_3672);
xor U9417 (N_9417,N_2716,N_3243);
and U9418 (N_9418,N_3422,N_1767);
xnor U9419 (N_9419,N_4033,N_3759);
xnor U9420 (N_9420,N_4036,N_2749);
or U9421 (N_9421,N_1034,N_388);
xor U9422 (N_9422,N_3856,N_3708);
and U9423 (N_9423,N_3778,N_1174);
or U9424 (N_9424,N_3504,N_802);
and U9425 (N_9425,N_1255,N_3604);
and U9426 (N_9426,N_4680,N_2994);
xor U9427 (N_9427,N_4354,N_1324);
nor U9428 (N_9428,N_115,N_1789);
nor U9429 (N_9429,N_3630,N_4518);
or U9430 (N_9430,N_3096,N_4284);
xor U9431 (N_9431,N_2869,N_3331);
xor U9432 (N_9432,N_3633,N_3041);
nor U9433 (N_9433,N_1749,N_4012);
or U9434 (N_9434,N_3086,N_202);
or U9435 (N_9435,N_1612,N_3410);
nand U9436 (N_9436,N_2602,N_2742);
nand U9437 (N_9437,N_4250,N_2403);
nor U9438 (N_9438,N_4422,N_262);
nor U9439 (N_9439,N_1030,N_757);
nor U9440 (N_9440,N_786,N_3765);
or U9441 (N_9441,N_1173,N_3950);
and U9442 (N_9442,N_51,N_3091);
nor U9443 (N_9443,N_2496,N_192);
or U9444 (N_9444,N_4879,N_811);
or U9445 (N_9445,N_1967,N_2863);
nor U9446 (N_9446,N_1195,N_1431);
and U9447 (N_9447,N_1038,N_3730);
nor U9448 (N_9448,N_1123,N_954);
xor U9449 (N_9449,N_1337,N_1668);
or U9450 (N_9450,N_2851,N_4361);
nor U9451 (N_9451,N_4657,N_283);
nand U9452 (N_9452,N_3280,N_2172);
nand U9453 (N_9453,N_2126,N_563);
nand U9454 (N_9454,N_2827,N_1294);
nor U9455 (N_9455,N_3864,N_2633);
or U9456 (N_9456,N_4995,N_1909);
nand U9457 (N_9457,N_1186,N_2466);
nor U9458 (N_9458,N_4803,N_1853);
xor U9459 (N_9459,N_4997,N_4526);
or U9460 (N_9460,N_3439,N_1452);
nand U9461 (N_9461,N_3897,N_1595);
nor U9462 (N_9462,N_1441,N_2665);
or U9463 (N_9463,N_4942,N_144);
or U9464 (N_9464,N_2166,N_3530);
nor U9465 (N_9465,N_4960,N_3093);
and U9466 (N_9466,N_3248,N_3848);
and U9467 (N_9467,N_4703,N_111);
and U9468 (N_9468,N_3671,N_4348);
nor U9469 (N_9469,N_4060,N_3550);
and U9470 (N_9470,N_3553,N_4936);
nand U9471 (N_9471,N_3699,N_1821);
nand U9472 (N_9472,N_1009,N_3593);
nand U9473 (N_9473,N_3557,N_4943);
or U9474 (N_9474,N_205,N_1894);
nand U9475 (N_9475,N_2256,N_1849);
and U9476 (N_9476,N_4290,N_2934);
xnor U9477 (N_9477,N_2577,N_989);
xnor U9478 (N_9478,N_2278,N_2256);
xnor U9479 (N_9479,N_362,N_4209);
nand U9480 (N_9480,N_2119,N_1966);
nand U9481 (N_9481,N_2832,N_4940);
or U9482 (N_9482,N_762,N_3444);
and U9483 (N_9483,N_4771,N_3603);
xor U9484 (N_9484,N_646,N_1156);
or U9485 (N_9485,N_3426,N_2474);
nand U9486 (N_9486,N_185,N_2079);
xor U9487 (N_9487,N_248,N_3769);
and U9488 (N_9488,N_2831,N_4432);
xor U9489 (N_9489,N_1596,N_3150);
xor U9490 (N_9490,N_3713,N_3093);
or U9491 (N_9491,N_4996,N_478);
or U9492 (N_9492,N_2613,N_778);
or U9493 (N_9493,N_2976,N_1841);
nor U9494 (N_9494,N_3730,N_2844);
or U9495 (N_9495,N_4272,N_235);
nor U9496 (N_9496,N_1835,N_1915);
and U9497 (N_9497,N_1702,N_1019);
xnor U9498 (N_9498,N_1079,N_3329);
nor U9499 (N_9499,N_1348,N_1616);
xnor U9500 (N_9500,N_4013,N_3339);
nor U9501 (N_9501,N_365,N_2504);
nand U9502 (N_9502,N_4225,N_3497);
nor U9503 (N_9503,N_4669,N_465);
xor U9504 (N_9504,N_559,N_2690);
and U9505 (N_9505,N_273,N_765);
nor U9506 (N_9506,N_1992,N_911);
or U9507 (N_9507,N_144,N_289);
or U9508 (N_9508,N_750,N_66);
or U9509 (N_9509,N_4386,N_727);
nor U9510 (N_9510,N_2086,N_1685);
xor U9511 (N_9511,N_973,N_4628);
xor U9512 (N_9512,N_1488,N_626);
nand U9513 (N_9513,N_1102,N_3229);
and U9514 (N_9514,N_2429,N_1873);
and U9515 (N_9515,N_2287,N_3344);
or U9516 (N_9516,N_150,N_1088);
nand U9517 (N_9517,N_3274,N_1970);
and U9518 (N_9518,N_3515,N_1268);
nand U9519 (N_9519,N_571,N_4082);
xnor U9520 (N_9520,N_667,N_2519);
and U9521 (N_9521,N_4898,N_118);
or U9522 (N_9522,N_4528,N_3957);
and U9523 (N_9523,N_3580,N_991);
nand U9524 (N_9524,N_2280,N_3558);
and U9525 (N_9525,N_1182,N_3523);
xor U9526 (N_9526,N_2289,N_4287);
nor U9527 (N_9527,N_1611,N_1582);
and U9528 (N_9528,N_4905,N_2064);
nor U9529 (N_9529,N_1776,N_706);
nor U9530 (N_9530,N_3836,N_3561);
and U9531 (N_9531,N_4420,N_44);
nand U9532 (N_9532,N_3127,N_743);
or U9533 (N_9533,N_4546,N_3283);
or U9534 (N_9534,N_2336,N_3894);
nor U9535 (N_9535,N_2231,N_4248);
or U9536 (N_9536,N_4674,N_4064);
nand U9537 (N_9537,N_2322,N_4458);
and U9538 (N_9538,N_402,N_2985);
xor U9539 (N_9539,N_2319,N_2139);
or U9540 (N_9540,N_1542,N_824);
or U9541 (N_9541,N_523,N_1904);
nor U9542 (N_9542,N_1137,N_3625);
nand U9543 (N_9543,N_812,N_4326);
or U9544 (N_9544,N_4560,N_2682);
nor U9545 (N_9545,N_2354,N_295);
xnor U9546 (N_9546,N_2608,N_383);
or U9547 (N_9547,N_4105,N_774);
nand U9548 (N_9548,N_188,N_4237);
and U9549 (N_9549,N_4094,N_1990);
nor U9550 (N_9550,N_4793,N_2363);
nor U9551 (N_9551,N_1771,N_4482);
nor U9552 (N_9552,N_1167,N_2493);
nor U9553 (N_9553,N_4566,N_4881);
or U9554 (N_9554,N_3444,N_4226);
nor U9555 (N_9555,N_3161,N_2572);
xnor U9556 (N_9556,N_3482,N_4725);
nand U9557 (N_9557,N_391,N_2503);
or U9558 (N_9558,N_3111,N_22);
nor U9559 (N_9559,N_4613,N_1235);
and U9560 (N_9560,N_4609,N_4892);
or U9561 (N_9561,N_3914,N_4373);
and U9562 (N_9562,N_3261,N_4715);
or U9563 (N_9563,N_3127,N_109);
nand U9564 (N_9564,N_2710,N_1480);
and U9565 (N_9565,N_3765,N_4218);
or U9566 (N_9566,N_2436,N_1456);
nand U9567 (N_9567,N_438,N_1978);
or U9568 (N_9568,N_1166,N_1227);
and U9569 (N_9569,N_2303,N_3767);
and U9570 (N_9570,N_3345,N_3478);
nor U9571 (N_9571,N_573,N_3359);
nor U9572 (N_9572,N_201,N_3874);
nor U9573 (N_9573,N_3377,N_4700);
nor U9574 (N_9574,N_2764,N_2568);
and U9575 (N_9575,N_562,N_4570);
xnor U9576 (N_9576,N_793,N_3829);
or U9577 (N_9577,N_2011,N_61);
and U9578 (N_9578,N_3695,N_2783);
nand U9579 (N_9579,N_2764,N_3786);
xnor U9580 (N_9580,N_3455,N_4116);
xor U9581 (N_9581,N_4796,N_2679);
or U9582 (N_9582,N_2382,N_3146);
nor U9583 (N_9583,N_1816,N_2722);
xnor U9584 (N_9584,N_492,N_65);
or U9585 (N_9585,N_4600,N_3273);
and U9586 (N_9586,N_3153,N_1833);
xnor U9587 (N_9587,N_4093,N_2209);
or U9588 (N_9588,N_3990,N_2435);
and U9589 (N_9589,N_4710,N_1297);
or U9590 (N_9590,N_2258,N_4909);
nor U9591 (N_9591,N_2140,N_3017);
nor U9592 (N_9592,N_2082,N_247);
nor U9593 (N_9593,N_1557,N_3247);
xnor U9594 (N_9594,N_1409,N_312);
and U9595 (N_9595,N_4287,N_1908);
or U9596 (N_9596,N_1460,N_1929);
xor U9597 (N_9597,N_827,N_2891);
and U9598 (N_9598,N_3258,N_1604);
and U9599 (N_9599,N_2233,N_1231);
and U9600 (N_9600,N_1120,N_1977);
nand U9601 (N_9601,N_4986,N_2970);
or U9602 (N_9602,N_1840,N_2483);
and U9603 (N_9603,N_895,N_3428);
nor U9604 (N_9604,N_4963,N_4119);
nand U9605 (N_9605,N_3789,N_1376);
nand U9606 (N_9606,N_3360,N_4503);
and U9607 (N_9607,N_2397,N_1908);
and U9608 (N_9608,N_4392,N_1868);
nor U9609 (N_9609,N_1549,N_273);
xor U9610 (N_9610,N_3294,N_364);
xnor U9611 (N_9611,N_1475,N_3355);
or U9612 (N_9612,N_2871,N_4430);
nand U9613 (N_9613,N_2749,N_2);
xnor U9614 (N_9614,N_3478,N_355);
nand U9615 (N_9615,N_3431,N_3166);
or U9616 (N_9616,N_1844,N_570);
xnor U9617 (N_9617,N_476,N_871);
and U9618 (N_9618,N_753,N_2697);
and U9619 (N_9619,N_3899,N_2631);
or U9620 (N_9620,N_352,N_4824);
nor U9621 (N_9621,N_2125,N_2480);
nor U9622 (N_9622,N_3631,N_1584);
nor U9623 (N_9623,N_1559,N_1024);
and U9624 (N_9624,N_4804,N_1050);
xor U9625 (N_9625,N_779,N_3278);
or U9626 (N_9626,N_2997,N_4515);
nand U9627 (N_9627,N_2031,N_319);
or U9628 (N_9628,N_1943,N_2159);
nand U9629 (N_9629,N_4969,N_1707);
nand U9630 (N_9630,N_1593,N_980);
nor U9631 (N_9631,N_266,N_1787);
and U9632 (N_9632,N_3377,N_4824);
xor U9633 (N_9633,N_2742,N_1401);
nor U9634 (N_9634,N_4591,N_1748);
and U9635 (N_9635,N_3300,N_3358);
and U9636 (N_9636,N_982,N_4529);
nand U9637 (N_9637,N_3781,N_4351);
xor U9638 (N_9638,N_3792,N_3881);
and U9639 (N_9639,N_1727,N_1804);
and U9640 (N_9640,N_1356,N_590);
nand U9641 (N_9641,N_1893,N_1152);
xor U9642 (N_9642,N_73,N_1125);
nand U9643 (N_9643,N_3372,N_2444);
and U9644 (N_9644,N_4180,N_4870);
nand U9645 (N_9645,N_2192,N_2870);
and U9646 (N_9646,N_2059,N_645);
or U9647 (N_9647,N_2951,N_3733);
xor U9648 (N_9648,N_4173,N_3806);
and U9649 (N_9649,N_1623,N_4162);
or U9650 (N_9650,N_330,N_4191);
and U9651 (N_9651,N_3767,N_719);
nor U9652 (N_9652,N_950,N_2155);
xor U9653 (N_9653,N_1327,N_3706);
or U9654 (N_9654,N_1236,N_3187);
and U9655 (N_9655,N_2645,N_1784);
or U9656 (N_9656,N_1464,N_1287);
or U9657 (N_9657,N_3181,N_4952);
and U9658 (N_9658,N_2180,N_517);
or U9659 (N_9659,N_2628,N_2672);
and U9660 (N_9660,N_1862,N_4797);
xnor U9661 (N_9661,N_1367,N_3633);
nor U9662 (N_9662,N_1251,N_4751);
or U9663 (N_9663,N_1902,N_332);
and U9664 (N_9664,N_691,N_2820);
nand U9665 (N_9665,N_4611,N_3735);
nand U9666 (N_9666,N_1889,N_730);
nand U9667 (N_9667,N_1394,N_703);
xor U9668 (N_9668,N_3745,N_4207);
nand U9669 (N_9669,N_3862,N_268);
nand U9670 (N_9670,N_3976,N_4192);
nand U9671 (N_9671,N_1486,N_4898);
nor U9672 (N_9672,N_2141,N_4622);
nor U9673 (N_9673,N_3584,N_3922);
nand U9674 (N_9674,N_1941,N_556);
nor U9675 (N_9675,N_4093,N_4976);
and U9676 (N_9676,N_2384,N_906);
and U9677 (N_9677,N_1466,N_4074);
xnor U9678 (N_9678,N_2645,N_1193);
and U9679 (N_9679,N_2605,N_176);
or U9680 (N_9680,N_3614,N_4554);
nand U9681 (N_9681,N_2795,N_3834);
and U9682 (N_9682,N_2877,N_488);
xor U9683 (N_9683,N_1554,N_3696);
nor U9684 (N_9684,N_4720,N_610);
nor U9685 (N_9685,N_62,N_3925);
and U9686 (N_9686,N_4608,N_1693);
xnor U9687 (N_9687,N_1414,N_1630);
nor U9688 (N_9688,N_3443,N_3588);
nand U9689 (N_9689,N_1682,N_573);
nand U9690 (N_9690,N_255,N_3035);
xor U9691 (N_9691,N_4346,N_720);
nor U9692 (N_9692,N_1029,N_1225);
xor U9693 (N_9693,N_4340,N_1513);
and U9694 (N_9694,N_4484,N_1374);
or U9695 (N_9695,N_3398,N_1716);
nand U9696 (N_9696,N_2697,N_3936);
and U9697 (N_9697,N_1401,N_2584);
and U9698 (N_9698,N_4170,N_4707);
xor U9699 (N_9699,N_2344,N_277);
nor U9700 (N_9700,N_3044,N_2524);
or U9701 (N_9701,N_4220,N_2300);
xnor U9702 (N_9702,N_4560,N_284);
nand U9703 (N_9703,N_1105,N_143);
or U9704 (N_9704,N_2220,N_3282);
or U9705 (N_9705,N_1652,N_3574);
or U9706 (N_9706,N_1971,N_2070);
xor U9707 (N_9707,N_1499,N_1444);
xnor U9708 (N_9708,N_4522,N_2889);
and U9709 (N_9709,N_2291,N_4126);
xnor U9710 (N_9710,N_1090,N_920);
nor U9711 (N_9711,N_2614,N_1507);
or U9712 (N_9712,N_2074,N_607);
and U9713 (N_9713,N_470,N_1047);
or U9714 (N_9714,N_3672,N_4643);
nor U9715 (N_9715,N_3489,N_4479);
or U9716 (N_9716,N_737,N_548);
nor U9717 (N_9717,N_2958,N_3169);
xnor U9718 (N_9718,N_2083,N_3847);
xnor U9719 (N_9719,N_2219,N_1177);
nor U9720 (N_9720,N_3967,N_2363);
and U9721 (N_9721,N_4560,N_1735);
nand U9722 (N_9722,N_2764,N_558);
and U9723 (N_9723,N_1307,N_1897);
xor U9724 (N_9724,N_1280,N_974);
nand U9725 (N_9725,N_1833,N_4283);
nor U9726 (N_9726,N_1559,N_4352);
nor U9727 (N_9727,N_2316,N_3643);
or U9728 (N_9728,N_3826,N_3937);
xor U9729 (N_9729,N_1186,N_4930);
nor U9730 (N_9730,N_4412,N_4071);
or U9731 (N_9731,N_3942,N_3374);
xnor U9732 (N_9732,N_393,N_3136);
nand U9733 (N_9733,N_387,N_3745);
or U9734 (N_9734,N_487,N_2169);
and U9735 (N_9735,N_2828,N_1734);
or U9736 (N_9736,N_1626,N_3789);
and U9737 (N_9737,N_3143,N_2818);
and U9738 (N_9738,N_642,N_762);
nand U9739 (N_9739,N_3728,N_2794);
or U9740 (N_9740,N_1410,N_1580);
xor U9741 (N_9741,N_738,N_4661);
nor U9742 (N_9742,N_2436,N_4242);
nand U9743 (N_9743,N_937,N_12);
and U9744 (N_9744,N_882,N_3384);
and U9745 (N_9745,N_4239,N_3070);
or U9746 (N_9746,N_1301,N_1528);
and U9747 (N_9747,N_4179,N_3259);
nand U9748 (N_9748,N_2976,N_3773);
nand U9749 (N_9749,N_278,N_99);
and U9750 (N_9750,N_1118,N_4311);
nor U9751 (N_9751,N_2390,N_4110);
xnor U9752 (N_9752,N_3616,N_4295);
and U9753 (N_9753,N_199,N_1168);
and U9754 (N_9754,N_1842,N_3099);
or U9755 (N_9755,N_1897,N_1782);
and U9756 (N_9756,N_3528,N_3462);
xnor U9757 (N_9757,N_995,N_4270);
and U9758 (N_9758,N_1622,N_2210);
and U9759 (N_9759,N_3629,N_1096);
nor U9760 (N_9760,N_1731,N_4193);
or U9761 (N_9761,N_827,N_3040);
nand U9762 (N_9762,N_3484,N_1324);
nor U9763 (N_9763,N_1412,N_1746);
or U9764 (N_9764,N_4275,N_3437);
or U9765 (N_9765,N_1960,N_3211);
and U9766 (N_9766,N_2447,N_2333);
or U9767 (N_9767,N_1526,N_4394);
and U9768 (N_9768,N_217,N_2261);
xor U9769 (N_9769,N_1982,N_4616);
xor U9770 (N_9770,N_4572,N_623);
nor U9771 (N_9771,N_229,N_2867);
or U9772 (N_9772,N_1404,N_3129);
and U9773 (N_9773,N_3114,N_2446);
or U9774 (N_9774,N_2106,N_2130);
and U9775 (N_9775,N_1824,N_881);
or U9776 (N_9776,N_4282,N_4740);
nand U9777 (N_9777,N_1282,N_2439);
xor U9778 (N_9778,N_4819,N_4325);
xnor U9779 (N_9779,N_4328,N_4618);
xnor U9780 (N_9780,N_328,N_3186);
xnor U9781 (N_9781,N_3786,N_2728);
nor U9782 (N_9782,N_597,N_3527);
nand U9783 (N_9783,N_4818,N_1678);
or U9784 (N_9784,N_2498,N_4442);
nor U9785 (N_9785,N_4131,N_3306);
xor U9786 (N_9786,N_1375,N_1196);
or U9787 (N_9787,N_455,N_3392);
and U9788 (N_9788,N_4754,N_2313);
nand U9789 (N_9789,N_3179,N_2044);
nor U9790 (N_9790,N_1707,N_32);
and U9791 (N_9791,N_4769,N_3912);
xnor U9792 (N_9792,N_2970,N_955);
nand U9793 (N_9793,N_3862,N_2560);
nor U9794 (N_9794,N_4984,N_537);
and U9795 (N_9795,N_1055,N_2441);
and U9796 (N_9796,N_4702,N_2311);
xnor U9797 (N_9797,N_4957,N_3704);
or U9798 (N_9798,N_3417,N_1342);
or U9799 (N_9799,N_2470,N_135);
and U9800 (N_9800,N_3393,N_2666);
xnor U9801 (N_9801,N_1457,N_2461);
nand U9802 (N_9802,N_2225,N_2085);
nor U9803 (N_9803,N_4544,N_4065);
or U9804 (N_9804,N_410,N_1315);
and U9805 (N_9805,N_898,N_4288);
and U9806 (N_9806,N_1902,N_3243);
nor U9807 (N_9807,N_1628,N_2274);
nand U9808 (N_9808,N_2734,N_4524);
nor U9809 (N_9809,N_4396,N_1858);
xnor U9810 (N_9810,N_2284,N_2224);
nand U9811 (N_9811,N_745,N_3525);
and U9812 (N_9812,N_3428,N_4164);
nand U9813 (N_9813,N_3019,N_2574);
nor U9814 (N_9814,N_2678,N_831);
or U9815 (N_9815,N_1788,N_4705);
xnor U9816 (N_9816,N_4534,N_4315);
nand U9817 (N_9817,N_4631,N_4074);
and U9818 (N_9818,N_4985,N_4996);
or U9819 (N_9819,N_78,N_2910);
nand U9820 (N_9820,N_3877,N_4920);
or U9821 (N_9821,N_4163,N_2333);
or U9822 (N_9822,N_2353,N_2777);
and U9823 (N_9823,N_286,N_2087);
nand U9824 (N_9824,N_1966,N_4505);
xor U9825 (N_9825,N_3432,N_2407);
or U9826 (N_9826,N_4690,N_4040);
xor U9827 (N_9827,N_3839,N_1643);
and U9828 (N_9828,N_4483,N_4973);
nor U9829 (N_9829,N_4209,N_882);
and U9830 (N_9830,N_609,N_1206);
xnor U9831 (N_9831,N_3393,N_1972);
nor U9832 (N_9832,N_1504,N_4686);
and U9833 (N_9833,N_1795,N_2603);
nand U9834 (N_9834,N_3807,N_1160);
and U9835 (N_9835,N_1489,N_2394);
xnor U9836 (N_9836,N_4580,N_1669);
xnor U9837 (N_9837,N_1937,N_3849);
xor U9838 (N_9838,N_3589,N_4567);
xnor U9839 (N_9839,N_3231,N_498);
nand U9840 (N_9840,N_361,N_1645);
and U9841 (N_9841,N_3034,N_666);
or U9842 (N_9842,N_694,N_2725);
nand U9843 (N_9843,N_1087,N_1348);
and U9844 (N_9844,N_2837,N_3472);
xor U9845 (N_9845,N_1385,N_1019);
nor U9846 (N_9846,N_3384,N_2639);
and U9847 (N_9847,N_4487,N_3715);
nor U9848 (N_9848,N_1704,N_1524);
or U9849 (N_9849,N_906,N_4643);
or U9850 (N_9850,N_3348,N_2625);
xor U9851 (N_9851,N_4128,N_4647);
and U9852 (N_9852,N_545,N_1007);
or U9853 (N_9853,N_792,N_1596);
nand U9854 (N_9854,N_4471,N_1843);
nor U9855 (N_9855,N_1276,N_3821);
xnor U9856 (N_9856,N_2334,N_2653);
nor U9857 (N_9857,N_657,N_3205);
and U9858 (N_9858,N_1608,N_2664);
xor U9859 (N_9859,N_1933,N_4938);
nand U9860 (N_9860,N_3042,N_104);
nor U9861 (N_9861,N_2393,N_967);
and U9862 (N_9862,N_4872,N_3308);
and U9863 (N_9863,N_66,N_4859);
and U9864 (N_9864,N_2284,N_3590);
nor U9865 (N_9865,N_3872,N_2757);
xor U9866 (N_9866,N_3548,N_2215);
nand U9867 (N_9867,N_565,N_1351);
nor U9868 (N_9868,N_3409,N_1757);
nor U9869 (N_9869,N_2257,N_2458);
nand U9870 (N_9870,N_1427,N_1239);
xnor U9871 (N_9871,N_2532,N_3966);
or U9872 (N_9872,N_3547,N_2600);
and U9873 (N_9873,N_3638,N_3255);
and U9874 (N_9874,N_3968,N_1401);
xor U9875 (N_9875,N_1606,N_1865);
or U9876 (N_9876,N_3409,N_1768);
xnor U9877 (N_9877,N_1264,N_4273);
nand U9878 (N_9878,N_1707,N_4033);
or U9879 (N_9879,N_1020,N_1019);
or U9880 (N_9880,N_1844,N_1053);
nand U9881 (N_9881,N_2527,N_4536);
nor U9882 (N_9882,N_3965,N_1228);
nor U9883 (N_9883,N_2438,N_213);
xor U9884 (N_9884,N_1221,N_4075);
or U9885 (N_9885,N_3476,N_500);
or U9886 (N_9886,N_2139,N_1958);
nand U9887 (N_9887,N_1904,N_3032);
nand U9888 (N_9888,N_3774,N_1234);
or U9889 (N_9889,N_1193,N_1368);
and U9890 (N_9890,N_3771,N_2795);
or U9891 (N_9891,N_133,N_2340);
and U9892 (N_9892,N_3880,N_268);
or U9893 (N_9893,N_1225,N_2391);
and U9894 (N_9894,N_3654,N_431);
nor U9895 (N_9895,N_1095,N_4593);
or U9896 (N_9896,N_3807,N_0);
nand U9897 (N_9897,N_3057,N_1844);
xor U9898 (N_9898,N_4622,N_1997);
nor U9899 (N_9899,N_2320,N_1965);
xnor U9900 (N_9900,N_4702,N_2094);
or U9901 (N_9901,N_2823,N_1002);
nand U9902 (N_9902,N_24,N_3701);
nor U9903 (N_9903,N_4685,N_1426);
nand U9904 (N_9904,N_438,N_659);
or U9905 (N_9905,N_407,N_4881);
and U9906 (N_9906,N_4694,N_255);
nor U9907 (N_9907,N_4576,N_182);
or U9908 (N_9908,N_2972,N_667);
xnor U9909 (N_9909,N_3642,N_279);
or U9910 (N_9910,N_1841,N_1837);
nor U9911 (N_9911,N_3138,N_2090);
or U9912 (N_9912,N_4763,N_916);
or U9913 (N_9913,N_57,N_3339);
or U9914 (N_9914,N_4512,N_3241);
xor U9915 (N_9915,N_307,N_1444);
or U9916 (N_9916,N_2531,N_4867);
or U9917 (N_9917,N_3686,N_1356);
and U9918 (N_9918,N_4205,N_2184);
and U9919 (N_9919,N_4560,N_3258);
nor U9920 (N_9920,N_4693,N_2152);
and U9921 (N_9921,N_832,N_2888);
nand U9922 (N_9922,N_2479,N_2055);
nor U9923 (N_9923,N_4515,N_4585);
xor U9924 (N_9924,N_2633,N_2172);
nor U9925 (N_9925,N_3671,N_677);
xor U9926 (N_9926,N_889,N_4476);
xnor U9927 (N_9927,N_767,N_3590);
xnor U9928 (N_9928,N_2795,N_2214);
and U9929 (N_9929,N_4886,N_4183);
nor U9930 (N_9930,N_4601,N_2733);
or U9931 (N_9931,N_1413,N_4413);
and U9932 (N_9932,N_4820,N_367);
and U9933 (N_9933,N_697,N_3278);
and U9934 (N_9934,N_4380,N_1057);
nand U9935 (N_9935,N_4948,N_1168);
nor U9936 (N_9936,N_593,N_4935);
and U9937 (N_9937,N_2154,N_2910);
or U9938 (N_9938,N_3392,N_3372);
and U9939 (N_9939,N_1836,N_1094);
and U9940 (N_9940,N_1215,N_885);
xor U9941 (N_9941,N_2250,N_3776);
nor U9942 (N_9942,N_4879,N_4570);
nor U9943 (N_9943,N_4541,N_2420);
or U9944 (N_9944,N_3860,N_3919);
nand U9945 (N_9945,N_4548,N_2291);
or U9946 (N_9946,N_2740,N_4625);
nand U9947 (N_9947,N_38,N_2756);
nand U9948 (N_9948,N_919,N_172);
or U9949 (N_9949,N_3157,N_1998);
or U9950 (N_9950,N_3912,N_1763);
xor U9951 (N_9951,N_2349,N_3343);
or U9952 (N_9952,N_327,N_4279);
nor U9953 (N_9953,N_4121,N_3802);
xor U9954 (N_9954,N_2670,N_1905);
nor U9955 (N_9955,N_695,N_3891);
and U9956 (N_9956,N_411,N_1514);
xor U9957 (N_9957,N_907,N_4263);
and U9958 (N_9958,N_1792,N_1135);
or U9959 (N_9959,N_4242,N_1003);
and U9960 (N_9960,N_485,N_1787);
or U9961 (N_9961,N_3866,N_1871);
nor U9962 (N_9962,N_2034,N_4363);
nand U9963 (N_9963,N_4971,N_4139);
xnor U9964 (N_9964,N_4641,N_4849);
xnor U9965 (N_9965,N_3701,N_4220);
nand U9966 (N_9966,N_2005,N_1336);
xnor U9967 (N_9967,N_1996,N_3564);
and U9968 (N_9968,N_3238,N_2399);
nor U9969 (N_9969,N_1526,N_4481);
or U9970 (N_9970,N_4031,N_4235);
nor U9971 (N_9971,N_37,N_146);
nand U9972 (N_9972,N_4814,N_1027);
xor U9973 (N_9973,N_3352,N_3261);
nand U9974 (N_9974,N_4424,N_4303);
and U9975 (N_9975,N_1734,N_2693);
nor U9976 (N_9976,N_4491,N_1013);
nand U9977 (N_9977,N_4998,N_907);
or U9978 (N_9978,N_3855,N_587);
and U9979 (N_9979,N_3731,N_1361);
and U9980 (N_9980,N_3352,N_1090);
or U9981 (N_9981,N_1647,N_2968);
and U9982 (N_9982,N_1525,N_3846);
xnor U9983 (N_9983,N_4236,N_2946);
nor U9984 (N_9984,N_2041,N_509);
and U9985 (N_9985,N_4594,N_2925);
nor U9986 (N_9986,N_4089,N_3652);
or U9987 (N_9987,N_4125,N_1915);
nor U9988 (N_9988,N_2109,N_3090);
nor U9989 (N_9989,N_477,N_557);
nor U9990 (N_9990,N_3209,N_1088);
nand U9991 (N_9991,N_4061,N_3028);
and U9992 (N_9992,N_189,N_4902);
nor U9993 (N_9993,N_1863,N_3749);
nor U9994 (N_9994,N_3986,N_2418);
nand U9995 (N_9995,N_3629,N_495);
and U9996 (N_9996,N_4922,N_2876);
or U9997 (N_9997,N_1343,N_621);
nor U9998 (N_9998,N_755,N_542);
xnor U9999 (N_9999,N_798,N_3947);
and U10000 (N_10000,N_6212,N_6007);
nand U10001 (N_10001,N_5285,N_9667);
xor U10002 (N_10002,N_8334,N_5404);
xor U10003 (N_10003,N_9291,N_7657);
nor U10004 (N_10004,N_8836,N_5445);
and U10005 (N_10005,N_9278,N_7781);
nand U10006 (N_10006,N_5969,N_5028);
and U10007 (N_10007,N_9181,N_9151);
nor U10008 (N_10008,N_5549,N_8830);
and U10009 (N_10009,N_9671,N_8828);
or U10010 (N_10010,N_7530,N_8464);
nor U10011 (N_10011,N_5794,N_6320);
or U10012 (N_10012,N_5482,N_5496);
or U10013 (N_10013,N_5121,N_6996);
or U10014 (N_10014,N_5552,N_7143);
and U10015 (N_10015,N_7582,N_7770);
nand U10016 (N_10016,N_8640,N_9322);
and U10017 (N_10017,N_8617,N_7252);
or U10018 (N_10018,N_7383,N_8506);
xnor U10019 (N_10019,N_8267,N_7815);
or U10020 (N_10020,N_8575,N_6621);
xor U10021 (N_10021,N_7200,N_6453);
and U10022 (N_10022,N_6850,N_6956);
xnor U10023 (N_10023,N_6823,N_7532);
and U10024 (N_10024,N_7328,N_5506);
nand U10025 (N_10025,N_9900,N_7754);
or U10026 (N_10026,N_8119,N_6716);
xnor U10027 (N_10027,N_7984,N_7416);
or U10028 (N_10028,N_9432,N_6395);
and U10029 (N_10029,N_9785,N_8672);
and U10030 (N_10030,N_7730,N_7878);
xnor U10031 (N_10031,N_8991,N_7660);
nor U10032 (N_10032,N_9566,N_8317);
nor U10033 (N_10033,N_5034,N_6458);
xor U10034 (N_10034,N_5278,N_8168);
or U10035 (N_10035,N_9150,N_5633);
nand U10036 (N_10036,N_7405,N_5171);
nor U10037 (N_10037,N_7159,N_7685);
or U10038 (N_10038,N_7947,N_6069);
and U10039 (N_10039,N_6442,N_9142);
nand U10040 (N_10040,N_5555,N_8905);
nor U10041 (N_10041,N_8588,N_6822);
nor U10042 (N_10042,N_7182,N_6142);
or U10043 (N_10043,N_5775,N_8998);
xnor U10044 (N_10044,N_5889,N_6265);
nor U10045 (N_10045,N_8893,N_7459);
or U10046 (N_10046,N_7933,N_5917);
nor U10047 (N_10047,N_7264,N_8897);
xnor U10048 (N_10048,N_6665,N_8148);
nand U10049 (N_10049,N_9551,N_8476);
xor U10050 (N_10050,N_8356,N_7964);
nor U10051 (N_10051,N_7958,N_6372);
and U10052 (N_10052,N_5959,N_7742);
and U10053 (N_10053,N_6494,N_6163);
or U10054 (N_10054,N_5948,N_8070);
and U10055 (N_10055,N_9219,N_8077);
or U10056 (N_10056,N_7084,N_9032);
xnor U10057 (N_10057,N_6539,N_5411);
nand U10058 (N_10058,N_5668,N_9310);
and U10059 (N_10059,N_6405,N_5999);
nand U10060 (N_10060,N_8207,N_9362);
and U10061 (N_10061,N_7192,N_5085);
nand U10062 (N_10062,N_8773,N_9969);
and U10063 (N_10063,N_9029,N_8565);
or U10064 (N_10064,N_6726,N_6485);
xnor U10065 (N_10065,N_7825,N_5058);
or U10066 (N_10066,N_9554,N_5540);
or U10067 (N_10067,N_8795,N_5813);
or U10068 (N_10068,N_9617,N_7032);
xnor U10069 (N_10069,N_7807,N_5421);
nand U10070 (N_10070,N_7583,N_7544);
xnor U10071 (N_10071,N_6607,N_5080);
or U10072 (N_10072,N_6098,N_6826);
nand U10073 (N_10073,N_7491,N_9556);
nand U10074 (N_10074,N_9696,N_7028);
nand U10075 (N_10075,N_8099,N_9862);
nor U10076 (N_10076,N_8601,N_9709);
nor U10077 (N_10077,N_8697,N_7727);
and U10078 (N_10078,N_5911,N_7251);
or U10079 (N_10079,N_8004,N_9393);
and U10080 (N_10080,N_6290,N_9620);
nand U10081 (N_10081,N_5339,N_6410);
and U10082 (N_10082,N_7374,N_7434);
nor U10083 (N_10083,N_5871,N_7848);
or U10084 (N_10084,N_8243,N_5606);
nor U10085 (N_10085,N_6421,N_6868);
xnor U10086 (N_10086,N_9914,N_6100);
or U10087 (N_10087,N_7981,N_8212);
xnor U10088 (N_10088,N_8360,N_7750);
nor U10089 (N_10089,N_5806,N_6640);
nor U10090 (N_10090,N_8739,N_8282);
or U10091 (N_10091,N_8481,N_5050);
nand U10092 (N_10092,N_9192,N_6579);
and U10093 (N_10093,N_8999,N_5043);
and U10094 (N_10094,N_5897,N_9640);
nand U10095 (N_10095,N_9416,N_6363);
nor U10096 (N_10096,N_6993,N_6364);
xor U10097 (N_10097,N_6240,N_8125);
or U10098 (N_10098,N_7323,N_7978);
or U10099 (N_10099,N_7077,N_6351);
nand U10100 (N_10100,N_8072,N_9853);
and U10101 (N_10101,N_6157,N_9560);
xnor U10102 (N_10102,N_8911,N_9692);
xor U10103 (N_10103,N_9272,N_5756);
nand U10104 (N_10104,N_6710,N_6377);
nand U10105 (N_10105,N_7334,N_8771);
xor U10106 (N_10106,N_9741,N_6629);
xor U10107 (N_10107,N_8044,N_8545);
and U10108 (N_10108,N_9833,N_9835);
nor U10109 (N_10109,N_5112,N_6548);
nand U10110 (N_10110,N_7123,N_7139);
xnor U10111 (N_10111,N_7505,N_9501);
or U10112 (N_10112,N_6269,N_7589);
xnor U10113 (N_10113,N_8711,N_7749);
xor U10114 (N_10114,N_7438,N_9541);
nor U10115 (N_10115,N_7164,N_9378);
or U10116 (N_10116,N_5861,N_9120);
nor U10117 (N_10117,N_8966,N_7795);
nand U10118 (N_10118,N_5183,N_8386);
xnor U10119 (N_10119,N_5648,N_6368);
nor U10120 (N_10120,N_5545,N_8139);
and U10121 (N_10121,N_5637,N_5597);
and U10122 (N_10122,N_7454,N_9894);
and U10123 (N_10123,N_6662,N_6695);
and U10124 (N_10124,N_9852,N_7635);
and U10125 (N_10125,N_7518,N_8537);
or U10126 (N_10126,N_8986,N_9847);
nand U10127 (N_10127,N_8400,N_6319);
and U10128 (N_10128,N_5995,N_8604);
or U10129 (N_10129,N_8889,N_6119);
and U10130 (N_10130,N_5521,N_9703);
and U10131 (N_10131,N_7724,N_5136);
or U10132 (N_10132,N_9413,N_6281);
nand U10133 (N_10133,N_8655,N_6615);
xnor U10134 (N_10134,N_5898,N_7350);
and U10135 (N_10135,N_7510,N_8758);
nand U10136 (N_10136,N_9866,N_6706);
and U10137 (N_10137,N_6602,N_7876);
and U10138 (N_10138,N_8598,N_5440);
and U10139 (N_10139,N_9173,N_5566);
xor U10140 (N_10140,N_7128,N_5417);
or U10141 (N_10141,N_8131,N_5685);
nand U10142 (N_10142,N_6914,N_6236);
and U10143 (N_10143,N_9713,N_6849);
nand U10144 (N_10144,N_7983,N_8814);
nand U10145 (N_10145,N_9925,N_9724);
nor U10146 (N_10146,N_9731,N_9759);
xnor U10147 (N_10147,N_9238,N_8549);
or U10148 (N_10148,N_9545,N_5732);
nor U10149 (N_10149,N_9936,N_9086);
nor U10150 (N_10150,N_8877,N_8230);
nand U10151 (N_10151,N_9816,N_8257);
xnor U10152 (N_10152,N_8067,N_8762);
xor U10153 (N_10153,N_6392,N_8487);
nor U10154 (N_10154,N_9654,N_6278);
nand U10155 (N_10155,N_6501,N_8741);
and U10156 (N_10156,N_8263,N_5922);
and U10157 (N_10157,N_5193,N_7569);
or U10158 (N_10158,N_7254,N_7609);
and U10159 (N_10159,N_8766,N_7331);
or U10160 (N_10160,N_7073,N_9448);
or U10161 (N_10161,N_7675,N_5746);
xnor U10162 (N_10162,N_5124,N_9186);
xor U10163 (N_10163,N_9243,N_6759);
and U10164 (N_10164,N_8443,N_7606);
nand U10165 (N_10165,N_5645,N_9528);
or U10166 (N_10166,N_9353,N_5832);
and U10167 (N_10167,N_6530,N_7414);
and U10168 (N_10168,N_8406,N_7037);
and U10169 (N_10169,N_8985,N_9022);
nor U10170 (N_10170,N_6027,N_7783);
or U10171 (N_10171,N_8523,N_6166);
xor U10172 (N_10172,N_6730,N_5131);
and U10173 (N_10173,N_5736,N_6468);
or U10174 (N_10174,N_5067,N_7697);
or U10175 (N_10175,N_9806,N_8394);
nand U10176 (N_10176,N_7101,N_8756);
xor U10177 (N_10177,N_5579,N_8731);
or U10178 (N_10178,N_6896,N_6630);
nand U10179 (N_10179,N_5011,N_9758);
nor U10180 (N_10180,N_9846,N_5338);
or U10181 (N_10181,N_9779,N_5992);
xnor U10182 (N_10182,N_9776,N_6591);
nor U10183 (N_10183,N_9331,N_9233);
nand U10184 (N_10184,N_9817,N_8325);
nor U10185 (N_10185,N_9146,N_9348);
xnor U10186 (N_10186,N_5610,N_5647);
and U10187 (N_10187,N_6198,N_5369);
nor U10188 (N_10188,N_6937,N_6891);
nor U10189 (N_10189,N_7113,N_9295);
nor U10190 (N_10190,N_8436,N_6248);
nand U10191 (N_10191,N_6291,N_5457);
and U10192 (N_10192,N_8793,N_8621);
nor U10193 (N_10193,N_5570,N_8913);
nand U10194 (N_10194,N_9625,N_7721);
or U10195 (N_10195,N_6857,N_9477);
and U10196 (N_10196,N_6418,N_8231);
xor U10197 (N_10197,N_8922,N_8181);
and U10198 (N_10198,N_8433,N_8339);
xnor U10199 (N_10199,N_7492,N_8603);
or U10200 (N_10200,N_5517,N_5209);
and U10201 (N_10201,N_5912,N_6385);
nor U10202 (N_10202,N_5475,N_7812);
xor U10203 (N_10203,N_5270,N_7311);
xnor U10204 (N_10204,N_7064,N_8554);
nor U10205 (N_10205,N_7584,N_9898);
or U10206 (N_10206,N_9190,N_6981);
xor U10207 (N_10207,N_7805,N_8473);
or U10208 (N_10208,N_5965,N_7295);
nor U10209 (N_10209,N_9434,N_5079);
and U10210 (N_10210,N_6231,N_6671);
or U10211 (N_10211,N_7508,N_5086);
nand U10212 (N_10212,N_9287,N_8422);
and U10213 (N_10213,N_5151,N_5788);
or U10214 (N_10214,N_7000,N_5013);
and U10215 (N_10215,N_7130,N_7687);
xnor U10216 (N_10216,N_6177,N_8191);
or U10217 (N_10217,N_8728,N_7118);
nor U10218 (N_10218,N_6354,N_8313);
xor U10219 (N_10219,N_5681,N_6712);
xor U10220 (N_10220,N_8201,N_9168);
and U10221 (N_10221,N_7081,N_9574);
or U10222 (N_10222,N_7935,N_5114);
nand U10223 (N_10223,N_5925,N_8918);
and U10224 (N_10224,N_9543,N_6005);
xor U10225 (N_10225,N_8624,N_9182);
nor U10226 (N_10226,N_9156,N_8724);
nand U10227 (N_10227,N_5162,N_5296);
nor U10228 (N_10228,N_9910,N_6229);
and U10229 (N_10229,N_7752,N_9125);
nor U10230 (N_10230,N_6070,N_9447);
and U10231 (N_10231,N_8306,N_8264);
and U10232 (N_10232,N_5614,N_5840);
xor U10233 (N_10233,N_9368,N_8428);
nor U10234 (N_10234,N_8145,N_5102);
and U10235 (N_10235,N_9949,N_9922);
nand U10236 (N_10236,N_8687,N_6725);
nor U10237 (N_10237,N_7571,N_8032);
or U10238 (N_10238,N_6031,N_5370);
nor U10239 (N_10239,N_9937,N_7355);
xnor U10240 (N_10240,N_5918,N_5282);
or U10241 (N_10241,N_8546,N_9444);
xor U10242 (N_10242,N_5656,N_5327);
nand U10243 (N_10243,N_6599,N_7605);
xnor U10244 (N_10244,N_5913,N_7865);
xor U10245 (N_10245,N_6958,N_9811);
or U10246 (N_10246,N_7940,N_6645);
or U10247 (N_10247,N_6397,N_6301);
nor U10248 (N_10248,N_5315,N_9431);
or U10249 (N_10249,N_9356,N_5763);
nand U10250 (N_10250,N_9657,N_7133);
nand U10251 (N_10251,N_9335,N_5800);
or U10252 (N_10252,N_6089,N_5373);
xnor U10253 (N_10253,N_8752,N_5699);
or U10254 (N_10254,N_6417,N_7757);
xnor U10255 (N_10255,N_8853,N_7973);
xnor U10256 (N_10256,N_6106,N_9481);
and U10257 (N_10257,N_9347,N_7124);
or U10258 (N_10258,N_9460,N_6636);
xnor U10259 (N_10259,N_8717,N_7803);
nor U10260 (N_10260,N_5405,N_9651);
and U10261 (N_10261,N_9145,N_6347);
nor U10262 (N_10262,N_5444,N_5748);
or U10263 (N_10263,N_6499,N_8579);
nor U10264 (N_10264,N_5608,N_8097);
nor U10265 (N_10265,N_5236,N_6147);
or U10266 (N_10266,N_8708,N_7900);
nand U10267 (N_10267,N_9496,N_8248);
xor U10268 (N_10268,N_9225,N_8699);
xor U10269 (N_10269,N_7796,N_7937);
xor U10270 (N_10270,N_7855,N_9301);
and U10271 (N_10271,N_7404,N_7849);
or U10272 (N_10272,N_8103,N_8748);
nand U10273 (N_10273,N_7247,N_5352);
nor U10274 (N_10274,N_7718,N_6552);
and U10275 (N_10275,N_9942,N_8530);
nor U10276 (N_10276,N_6964,N_5300);
nand U10277 (N_10277,N_6804,N_7633);
xor U10278 (N_10278,N_9637,N_7282);
xor U10279 (N_10279,N_9318,N_6832);
xnor U10280 (N_10280,N_8484,N_9209);
or U10281 (N_10281,N_9716,N_8471);
and U10282 (N_10282,N_7108,N_9215);
nand U10283 (N_10283,N_8517,N_7991);
or U10284 (N_10284,N_5558,N_5189);
or U10285 (N_10285,N_6718,N_9178);
xor U10286 (N_10286,N_7104,N_9672);
and U10287 (N_10287,N_7686,N_8767);
xnor U10288 (N_10288,N_7408,N_6673);
nand U10289 (N_10289,N_9237,N_7538);
and U10290 (N_10290,N_6855,N_8178);
and U10291 (N_10291,N_9730,N_5509);
nand U10292 (N_10292,N_8492,N_5795);
xnor U10293 (N_10293,N_6529,N_6437);
or U10294 (N_10294,N_6039,N_9061);
xor U10295 (N_10295,N_9329,N_7594);
and U10296 (N_10296,N_5764,N_5895);
nor U10297 (N_10297,N_8040,N_6181);
and U10298 (N_10298,N_8206,N_6952);
nand U10299 (N_10299,N_6776,N_9189);
or U10300 (N_10300,N_6332,N_6409);
xnor U10301 (N_10301,N_8623,N_7612);
nand U10302 (N_10302,N_6924,N_6035);
nand U10303 (N_10303,N_6722,N_6191);
xnor U10304 (N_10304,N_6666,N_6566);
nor U10305 (N_10305,N_6061,N_7776);
nand U10306 (N_10306,N_6935,N_8886);
xnor U10307 (N_10307,N_9154,N_5152);
and U10308 (N_10308,N_6481,N_7548);
and U10309 (N_10309,N_8126,N_6909);
or U10310 (N_10310,N_9712,N_9558);
nor U10311 (N_10311,N_8210,N_6279);
or U10312 (N_10312,N_5516,N_6321);
xor U10313 (N_10313,N_8254,N_9748);
xor U10314 (N_10314,N_9803,N_7047);
or U10315 (N_10315,N_6114,N_8496);
xnor U10316 (N_10316,N_8234,N_9899);
nand U10317 (N_10317,N_5265,N_5063);
or U10318 (N_10318,N_5602,N_9139);
and U10319 (N_10319,N_9786,N_5505);
xnor U10320 (N_10320,N_6985,N_9208);
nor U10321 (N_10321,N_9793,N_6155);
xor U10322 (N_10322,N_9170,N_7533);
nand U10323 (N_10323,N_9955,N_6327);
or U10324 (N_10324,N_8096,N_9406);
or U10325 (N_10325,N_7216,N_9913);
nor U10326 (N_10326,N_8246,N_9661);
xnor U10327 (N_10327,N_7648,N_8029);
or U10328 (N_10328,N_5293,N_5256);
nand U10329 (N_10329,N_9921,N_9599);
nand U10330 (N_10330,N_8668,N_5858);
nand U10331 (N_10331,N_8714,N_6498);
and U10332 (N_10332,N_9924,N_8020);
nand U10333 (N_10333,N_7570,N_7075);
and U10334 (N_10334,N_7246,N_7483);
nand U10335 (N_10335,N_6145,N_9603);
nor U10336 (N_10336,N_7762,N_5447);
and U10337 (N_10337,N_8883,N_9658);
and U10338 (N_10338,N_5829,N_6919);
nor U10339 (N_10339,N_9777,N_9941);
nor U10340 (N_10340,N_5423,N_7674);
nand U10341 (N_10341,N_6553,N_6340);
nor U10342 (N_10342,N_7440,N_6307);
nor U10343 (N_10343,N_8352,N_8896);
xor U10344 (N_10344,N_5228,N_7470);
or U10345 (N_10345,N_8785,N_7860);
nand U10346 (N_10346,N_9166,N_9263);
nor U10347 (N_10347,N_7289,N_5587);
or U10348 (N_10348,N_6842,N_7156);
or U10349 (N_10349,N_7550,N_7751);
or U10350 (N_10350,N_8713,N_6173);
and U10351 (N_10351,N_6831,N_9693);
or U10352 (N_10352,N_5479,N_5468);
xor U10353 (N_10353,N_5975,N_7877);
xnor U10354 (N_10354,N_5119,N_5808);
and U10355 (N_10355,N_9380,N_5810);
nand U10356 (N_10356,N_5461,N_6918);
or U10357 (N_10357,N_8875,N_9026);
and U10358 (N_10358,N_7952,N_6475);
nand U10359 (N_10359,N_5288,N_9122);
or U10360 (N_10360,N_6911,N_8784);
nor U10361 (N_10361,N_9733,N_5357);
and U10362 (N_10362,N_5707,N_7337);
and U10363 (N_10363,N_7103,N_8887);
nor U10364 (N_10364,N_5534,N_9371);
or U10365 (N_10365,N_5585,N_8845);
xor U10366 (N_10366,N_6976,N_6339);
nor U10367 (N_10367,N_9751,N_7050);
or U10368 (N_10368,N_6510,N_5919);
or U10369 (N_10369,N_6219,N_8482);
nor U10370 (N_10370,N_6803,N_9152);
or U10371 (N_10371,N_5693,N_5100);
and U10372 (N_10372,N_9979,N_9388);
nor U10373 (N_10373,N_6003,N_8380);
xor U10374 (N_10374,N_7627,N_8150);
xor U10375 (N_10375,N_8102,N_6205);
and U10376 (N_10376,N_5432,N_6051);
and U10377 (N_10377,N_7689,N_8894);
and U10378 (N_10378,N_7562,N_6491);
nand U10379 (N_10379,N_8904,N_9052);
nor U10380 (N_10380,N_9149,N_6777);
nand U10381 (N_10381,N_5845,N_9333);
xnor U10382 (N_10382,N_5298,N_5531);
nor U10383 (N_10383,N_6611,N_8121);
xor U10384 (N_10384,N_9714,N_9246);
xor U10385 (N_10385,N_9115,N_9462);
nor U10386 (N_10386,N_6528,N_6495);
nor U10387 (N_10387,N_5786,N_6605);
nand U10388 (N_10388,N_8123,N_6006);
nand U10389 (N_10389,N_5695,N_7632);
or U10390 (N_10390,N_5787,N_6882);
nor U10391 (N_10391,N_7154,N_9196);
nand U10392 (N_10392,N_6478,N_5044);
xor U10393 (N_10393,N_9267,N_9988);
nor U10394 (N_10394,N_7843,N_7198);
nand U10395 (N_10395,N_7052,N_5957);
or U10396 (N_10396,N_9705,N_6268);
or U10397 (N_10397,N_6818,N_9389);
and U10398 (N_10398,N_8445,N_5053);
nand U10399 (N_10399,N_8650,N_5723);
nor U10400 (N_10400,N_6677,N_8223);
xnor U10401 (N_10401,N_7960,N_7391);
and U10402 (N_10402,N_7402,N_5933);
nor U10403 (N_10403,N_6598,N_7946);
nor U10404 (N_10404,N_7189,N_6391);
nor U10405 (N_10405,N_8089,N_6572);
and U10406 (N_10406,N_8388,N_8671);
xnor U10407 (N_10407,N_7939,N_7305);
nand U10408 (N_10408,N_7953,N_6900);
nand U10409 (N_10409,N_5462,N_6427);
and U10410 (N_10410,N_6564,N_6751);
xnor U10411 (N_10411,N_6692,N_6245);
nand U10412 (N_10412,N_5138,N_6997);
or U10413 (N_10413,N_6056,N_5223);
nand U10414 (N_10414,N_6073,N_9334);
and U10415 (N_10415,N_8943,N_5660);
and U10416 (N_10416,N_8541,N_9831);
xor U10417 (N_10417,N_8982,N_8417);
and U10418 (N_10418,N_9297,N_5014);
xor U10419 (N_10419,N_8002,N_7021);
nor U10420 (N_10420,N_6595,N_9597);
nor U10421 (N_10421,N_6578,N_5567);
nand U10422 (N_10422,N_8910,N_6953);
nand U10423 (N_10423,N_7679,N_9126);
or U10424 (N_10424,N_5499,N_9083);
nand U10425 (N_10425,N_7814,N_7654);
nand U10426 (N_10426,N_5409,N_9236);
nand U10427 (N_10427,N_7925,N_9670);
or U10428 (N_10428,N_6330,N_7703);
nor U10429 (N_10429,N_9782,N_5269);
and U10430 (N_10430,N_6134,N_6833);
and U10431 (N_10431,N_5002,N_8408);
and U10432 (N_10432,N_9283,N_5560);
and U10433 (N_10433,N_7363,N_6542);
nand U10434 (N_10434,N_9858,N_6667);
nand U10435 (N_10435,N_8618,N_5064);
and U10436 (N_10436,N_8000,N_9884);
or U10437 (N_10437,N_6715,N_5205);
xnor U10438 (N_10438,N_9679,N_8049);
or U10439 (N_10439,N_5562,N_5007);
nor U10440 (N_10440,N_6717,N_5759);
nand U10441 (N_10441,N_9517,N_8439);
nand U10442 (N_10442,N_5953,N_6102);
nand U10443 (N_10443,N_5493,N_5535);
or U10444 (N_10444,N_9983,N_5692);
nor U10445 (N_10445,N_7857,N_9935);
nor U10446 (N_10446,N_7065,N_6511);
and U10447 (N_10447,N_8151,N_6011);
or U10448 (N_10448,N_6954,N_8790);
nand U10449 (N_10449,N_9970,N_8494);
and U10450 (N_10450,N_6258,N_6854);
or U10451 (N_10451,N_7788,N_5816);
nor U10452 (N_10452,N_7928,N_8751);
nand U10453 (N_10453,N_6786,N_7996);
xor U10454 (N_10454,N_9342,N_5978);
nor U10455 (N_10455,N_5783,N_8147);
and U10456 (N_10456,N_5422,N_7437);
xnor U10457 (N_10457,N_7327,N_9435);
nor U10458 (N_10458,N_8085,N_9093);
nor U10459 (N_10459,N_9338,N_7560);
or U10460 (N_10460,N_6772,N_8686);
xnor U10461 (N_10461,N_7922,N_8971);
and U10462 (N_10462,N_5330,N_5197);
xnor U10463 (N_10463,N_5230,N_9953);
xor U10464 (N_10464,N_9877,N_8050);
xor U10465 (N_10465,N_9259,N_9856);
nand U10466 (N_10466,N_5239,N_8120);
nor U10467 (N_10467,N_9091,N_8843);
and U10468 (N_10468,N_7817,N_9619);
nor U10469 (N_10469,N_7333,N_7856);
xnor U10470 (N_10470,N_9140,N_6685);
nand U10471 (N_10471,N_6209,N_5908);
nor U10472 (N_10472,N_5546,N_6654);
xnor U10473 (N_10473,N_7708,N_6783);
nand U10474 (N_10474,N_9804,N_7593);
or U10475 (N_10475,N_5945,N_6676);
nor U10476 (N_10476,N_5356,N_6570);
or U10477 (N_10477,N_6461,N_7135);
nor U10478 (N_10478,N_8721,N_5024);
nand U10479 (N_10479,N_8582,N_7672);
and U10480 (N_10480,N_9212,N_6086);
nand U10481 (N_10481,N_7668,N_5711);
or U10482 (N_10482,N_8193,N_7810);
nand U10483 (N_10483,N_5891,N_9162);
nand U10484 (N_10484,N_8727,N_8434);
xnor U10485 (N_10485,N_6479,N_9036);
nor U10486 (N_10486,N_9621,N_5888);
or U10487 (N_10487,N_7565,N_9017);
and U10488 (N_10488,N_8303,N_9198);
nand U10489 (N_10489,N_9454,N_8399);
nor U10490 (N_10490,N_8340,N_7442);
or U10491 (N_10491,N_9085,N_8684);
xnor U10492 (N_10492,N_5122,N_6420);
and U10493 (N_10493,N_9644,N_6210);
or U10494 (N_10494,N_6423,N_7448);
nand U10495 (N_10495,N_7986,N_6447);
nand U10496 (N_10496,N_6293,N_5433);
or U10497 (N_10497,N_8689,N_7869);
and U10498 (N_10498,N_8202,N_5618);
nor U10499 (N_10499,N_7870,N_6022);
and U10500 (N_10500,N_9702,N_8683);
or U10501 (N_10501,N_7255,N_9773);
xnor U10502 (N_10502,N_8415,N_8309);
nand U10503 (N_10503,N_7944,N_5182);
and U10504 (N_10504,N_6913,N_6451);
nor U10505 (N_10505,N_8286,N_5176);
xor U10506 (N_10506,N_9881,N_5156);
nor U10507 (N_10507,N_6249,N_9616);
or U10508 (N_10508,N_5773,N_9129);
and U10509 (N_10509,N_7656,N_9601);
xor U10510 (N_10510,N_7203,N_7961);
or U10511 (N_10511,N_9655,N_9766);
or U10512 (N_10512,N_6619,N_9019);
nor U10513 (N_10513,N_9094,N_8364);
nand U10514 (N_10514,N_9893,N_6805);
or U10515 (N_10515,N_7759,N_9700);
xor U10516 (N_10516,N_9211,N_5986);
or U10517 (N_10517,N_7932,N_9131);
and U10518 (N_10518,N_8874,N_7617);
and U10519 (N_10519,N_8581,N_9442);
or U10520 (N_10520,N_6257,N_6160);
xnor U10521 (N_10521,N_5510,N_8074);
nor U10522 (N_10522,N_9926,N_6734);
nand U10523 (N_10523,N_7060,N_6659);
nand U10524 (N_10524,N_8110,N_8700);
or U10525 (N_10525,N_6674,N_9028);
nand U10526 (N_10526,N_8284,N_7144);
or U10527 (N_10527,N_9401,N_6502);
xnor U10528 (N_10528,N_6225,N_9155);
and U10529 (N_10529,N_7951,N_8957);
and U10530 (N_10530,N_8869,N_9227);
xor U10531 (N_10531,N_8323,N_6262);
or U10532 (N_10532,N_5353,N_5295);
and U10533 (N_10533,N_8937,N_7998);
or U10534 (N_10534,N_6273,N_7469);
nand U10535 (N_10535,N_5881,N_8602);
xnor U10536 (N_10536,N_8587,N_7340);
xor U10537 (N_10537,N_6661,N_7300);
nor U10538 (N_10538,N_8108,N_5803);
or U10539 (N_10539,N_6897,N_5848);
and U10540 (N_10540,N_7704,N_9947);
nand U10541 (N_10541,N_6524,N_8631);
nand U10542 (N_10542,N_6756,N_7006);
and U10543 (N_10543,N_9127,N_5514);
or U10544 (N_10544,N_8091,N_6193);
and U10545 (N_10545,N_8827,N_6038);
nor U10546 (N_10546,N_5244,N_9684);
xor U10547 (N_10547,N_5082,N_5669);
nand U10548 (N_10548,N_6400,N_8558);
nor U10549 (N_10549,N_6250,N_7163);
nor U10550 (N_10550,N_5492,N_7005);
nand U10551 (N_10551,N_8539,N_9873);
xnor U10552 (N_10552,N_9066,N_8167);
nor U10553 (N_10553,N_8307,N_6691);
or U10554 (N_10554,N_5657,N_8591);
xor U10555 (N_10555,N_8393,N_8805);
or U10556 (N_10556,N_7030,N_8955);
nor U10557 (N_10557,N_9531,N_7468);
nand U10558 (N_10558,N_9521,N_9213);
and U10559 (N_10559,N_8373,N_7755);
and U10560 (N_10560,N_9499,N_8759);
nor U10561 (N_10561,N_5283,N_8124);
nand U10562 (N_10562,N_6713,N_7314);
and U10563 (N_10563,N_5859,N_5989);
xor U10564 (N_10564,N_7445,N_7186);
or U10565 (N_10565,N_5905,N_8787);
and U10566 (N_10566,N_6892,N_9830);
nand U10567 (N_10567,N_8462,N_8101);
nand U10568 (N_10568,N_5988,N_9891);
or U10569 (N_10569,N_9157,N_7572);
and U10570 (N_10570,N_6525,N_6276);
or U10571 (N_10571,N_7224,N_9252);
and U10572 (N_10572,N_5456,N_6184);
nand U10573 (N_10573,N_6312,N_8118);
and U10574 (N_10574,N_7033,N_5257);
nand U10575 (N_10575,N_5181,N_5104);
and U10576 (N_10576,N_8941,N_8540);
nor U10577 (N_10577,N_9195,N_5682);
or U10578 (N_10578,N_5751,N_9916);
and U10579 (N_10579,N_8132,N_9544);
xor U10580 (N_10580,N_8543,N_9859);
and U10581 (N_10581,N_7578,N_5233);
nand U10582 (N_10582,N_6176,N_7839);
or U10583 (N_10583,N_9999,N_7899);
nor U10584 (N_10584,N_8857,N_9842);
or U10585 (N_10585,N_8807,N_7158);
or U10586 (N_10586,N_8651,N_8600);
and U10587 (N_10587,N_5718,N_9070);
and U10588 (N_10588,N_8038,N_6370);
and U10589 (N_10589,N_9372,N_8486);
and U10590 (N_10590,N_9418,N_9271);
nor U10591 (N_10591,N_8336,N_5304);
nand U10592 (N_10592,N_7769,N_5714);
or U10593 (N_10593,N_5247,N_7592);
xor U10594 (N_10594,N_7142,N_5850);
nor U10595 (N_10595,N_5446,N_9270);
and U10596 (N_10596,N_7741,N_9948);
or U10597 (N_10597,N_8653,N_8674);
and U10598 (N_10598,N_9719,N_9582);
nor U10599 (N_10599,N_7979,N_8753);
and U10600 (N_10600,N_8521,N_9732);
xor U10601 (N_10601,N_5110,N_8789);
nand U10602 (N_10602,N_8738,N_8022);
nand U10603 (N_10603,N_7464,N_7458);
nand U10604 (N_10604,N_7017,N_5092);
or U10605 (N_10605,N_6845,N_5224);
xnor U10606 (N_10606,N_5191,N_7357);
nor U10607 (N_10607,N_6887,N_7036);
nor U10608 (N_10608,N_6190,N_9137);
or U10609 (N_10609,N_6969,N_7371);
and U10610 (N_10610,N_7054,N_5069);
nor U10611 (N_10611,N_8607,N_6681);
nor U10612 (N_10612,N_9929,N_7456);
or U10613 (N_10613,N_8750,N_7919);
nand U10614 (N_10614,N_8823,N_6575);
nor U10615 (N_10615,N_7479,N_5812);
xnor U10616 (N_10616,N_5164,N_6592);
nand U10617 (N_10617,N_8391,N_5862);
or U10618 (N_10618,N_7955,N_6890);
xor U10619 (N_10619,N_8329,N_7670);
nor U10620 (N_10620,N_8791,N_8289);
or U10621 (N_10621,N_7649,N_7179);
nor U10622 (N_10622,N_7829,N_7520);
nand U10623 (N_10623,N_5821,N_8536);
and U10624 (N_10624,N_6207,N_8172);
xnor U10625 (N_10625,N_7819,N_5441);
and U10626 (N_10626,N_7267,N_6237);
and U10627 (N_10627,N_7014,N_6886);
xnor U10628 (N_10628,N_5267,N_7738);
xnor U10629 (N_10629,N_6698,N_5753);
or U10630 (N_10630,N_6424,N_9459);
and U10631 (N_10631,N_9174,N_7471);
xnor U10632 (N_10632,N_6213,N_5039);
and U10633 (N_10633,N_7909,N_9647);
and U10634 (N_10634,N_8184,N_9863);
and U10635 (N_10635,N_7547,N_5167);
nor U10636 (N_10636,N_8405,N_5512);
nand U10637 (N_10637,N_8271,N_8662);
and U10638 (N_10638,N_9191,N_6241);
nor U10639 (N_10639,N_5569,N_8940);
nor U10640 (N_10640,N_8259,N_9218);
and U10641 (N_10641,N_6084,N_9183);
xnor U10642 (N_10642,N_5939,N_7926);
or U10643 (N_10643,N_5683,N_8799);
xor U10644 (N_10644,N_6927,N_5573);
and U10645 (N_10645,N_9102,N_6302);
nand U10646 (N_10646,N_6457,N_6353);
and U10647 (N_10647,N_8116,N_7949);
nand U10648 (N_10648,N_6083,N_5297);
nand U10649 (N_10649,N_9886,N_7862);
xnor U10650 (N_10650,N_5469,N_5649);
and U10651 (N_10651,N_7324,N_6104);
nand U10652 (N_10652,N_9476,N_7098);
nor U10653 (N_10653,N_5674,N_6840);
or U10654 (N_10654,N_9665,N_8235);
and U10655 (N_10655,N_8547,N_7826);
xnor U10656 (N_10656,N_5650,N_8967);
nand U10657 (N_10657,N_8636,N_7356);
xnor U10658 (N_10658,N_7901,N_7574);
nand U10659 (N_10659,N_8308,N_8765);
or U10660 (N_10660,N_5609,N_8083);
xnor U10661 (N_10661,N_5463,N_5201);
or U10662 (N_10662,N_7339,N_6693);
xnor U10663 (N_10663,N_6381,N_8693);
or U10664 (N_10664,N_7141,N_9728);
nand U10665 (N_10665,N_7431,N_5883);
nand U10666 (N_10666,N_7699,N_6757);
xor U10667 (N_10667,N_5839,N_6224);
nand U10668 (N_10668,N_9557,N_8338);
nor U10669 (N_10669,N_9855,N_9510);
nand U10670 (N_10670,N_9682,N_6150);
nand U10671 (N_10671,N_6226,N_6095);
or U10672 (N_10672,N_6851,N_9905);
nor U10673 (N_10673,N_7588,N_9355);
or U10674 (N_10674,N_8048,N_5684);
and U10675 (N_10675,N_7873,N_9888);
and U10676 (N_10676,N_5291,N_6382);
nand U10677 (N_10677,N_7284,N_9014);
nand U10678 (N_10678,N_5670,N_6120);
and U10679 (N_10679,N_9967,N_9286);
xnor U10680 (N_10680,N_5500,N_7969);
and U10681 (N_10681,N_8115,N_9033);
and U10682 (N_10682,N_9653,N_5252);
xnor U10683 (N_10683,N_6148,N_6483);
xor U10684 (N_10684,N_9740,N_9135);
and U10685 (N_10685,N_6168,N_6508);
and U10686 (N_10686,N_9928,N_5589);
or U10687 (N_10687,N_8045,N_7982);
or U10688 (N_10688,N_7793,N_9345);
nor U10689 (N_10689,N_7972,N_9051);
or U10690 (N_10690,N_8114,N_6135);
and U10691 (N_10691,N_6577,N_9711);
and U10692 (N_10692,N_7426,N_7507);
xor U10693 (N_10693,N_5385,N_6632);
xnor U10694 (N_10694,N_6813,N_6652);
nor U10695 (N_10695,N_6182,N_6308);
and U10696 (N_10696,N_7669,N_6439);
nor U10697 (N_10697,N_6346,N_5076);
nor U10698 (N_10698,N_9718,N_5188);
nand U10699 (N_10699,N_5084,N_7066);
xor U10700 (N_10700,N_8834,N_5915);
xnor U10701 (N_10701,N_9755,N_7097);
nor U10702 (N_10702,N_8295,N_9176);
xor U10703 (N_10703,N_7667,N_8312);
nand U10704 (N_10704,N_6318,N_8780);
and U10705 (N_10705,N_5466,N_8198);
and U10706 (N_10706,N_7038,N_6446);
and U10707 (N_10707,N_9379,N_5792);
or U10708 (N_10708,N_9715,N_5936);
nand U10709 (N_10709,N_7702,N_7515);
nand U10710 (N_10710,N_8559,N_5120);
or U10711 (N_10711,N_8171,N_9633);
nor U10712 (N_10712,N_9055,N_7119);
nor U10713 (N_10713,N_7923,N_6796);
xor U10714 (N_10714,N_7837,N_9317);
nor U10715 (N_10715,N_5153,N_7076);
or U10716 (N_10716,N_8855,N_6774);
and U10717 (N_10717,N_7830,N_6864);
nand U10718 (N_10718,N_8626,N_5113);
and U10719 (N_10719,N_5276,N_6093);
nand U10720 (N_10720,N_7147,N_5166);
xor U10721 (N_10721,N_9717,N_8898);
and U10722 (N_10722,N_8163,N_7595);
nor U10723 (N_10723,N_9902,N_5460);
and U10724 (N_10724,N_8993,N_7536);
xnor U10725 (N_10725,N_7622,N_6675);
nor U10726 (N_10726,N_8228,N_6580);
or U10727 (N_10727,N_8095,N_6137);
and U10728 (N_10728,N_9750,N_9753);
and U10729 (N_10729,N_6023,N_5822);
nand U10730 (N_10730,N_9160,N_8001);
or U10731 (N_10731,N_9324,N_5501);
xor U10732 (N_10732,N_5074,N_5761);
nor U10733 (N_10733,N_9296,N_9819);
and U10734 (N_10734,N_9944,N_7338);
xor U10735 (N_10735,N_6739,N_9165);
xor U10736 (N_10736,N_9080,N_5524);
nor U10737 (N_10737,N_5018,N_7963);
and U10738 (N_10738,N_6438,N_8880);
xnor U10739 (N_10739,N_8696,N_8705);
nor U10740 (N_10740,N_8774,N_5379);
xor U10741 (N_10741,N_8324,N_5782);
nor U10742 (N_10742,N_5318,N_8299);
xnor U10743 (N_10743,N_7231,N_6999);
nor U10744 (N_10744,N_9484,N_9456);
xor U10745 (N_10745,N_8681,N_7872);
nor U10746 (N_10746,N_5068,N_6477);
xor U10747 (N_10747,N_9527,N_5680);
xor U10748 (N_10748,N_5778,N_8007);
and U10749 (N_10749,N_7466,N_8735);
xor U10750 (N_10750,N_6720,N_7364);
xor U10751 (N_10751,N_9792,N_6723);
nor U10752 (N_10752,N_6081,N_8361);
nor U10753 (N_10753,N_5326,N_9791);
nand U10754 (N_10754,N_7765,N_5321);
nand U10755 (N_10755,N_8963,N_7265);
nand U10756 (N_10756,N_8796,N_9638);
xnor U10757 (N_10757,N_5582,N_7740);
nand U10758 (N_10758,N_7106,N_5192);
and U10759 (N_10759,N_5486,N_7858);
xnor U10760 (N_10760,N_6445,N_9870);
nor U10761 (N_10761,N_7304,N_7245);
or U10762 (N_10762,N_5745,N_7537);
nand U10763 (N_10763,N_9232,N_5442);
nor U10764 (N_10764,N_8497,N_8291);
nor U10765 (N_10765,N_9171,N_7748);
nand U10766 (N_10766,N_7171,N_5200);
or U10767 (N_10767,N_5434,N_9167);
and U10768 (N_10768,N_8768,N_7867);
or U10769 (N_10769,N_8818,N_9265);
and U10770 (N_10770,N_9666,N_6802);
and U10771 (N_10771,N_8638,N_7117);
nor U10772 (N_10772,N_7087,N_7244);
and U10773 (N_10773,N_8844,N_7987);
nor U10774 (N_10774,N_5094,N_5655);
xnor U10775 (N_10775,N_5578,N_6972);
or U10776 (N_10776,N_5144,N_5346);
nor U10777 (N_10777,N_7904,N_7274);
or U10778 (N_10778,N_7618,N_7063);
or U10779 (N_10779,N_8915,N_9562);
or U10780 (N_10780,N_9974,N_5343);
nand U10781 (N_10781,N_6747,N_5117);
xor U10782 (N_10782,N_9593,N_5632);
and U10783 (N_10783,N_5332,N_7840);
xor U10784 (N_10784,N_6811,N_7678);
or U10785 (N_10785,N_9344,N_5355);
and U10786 (N_10786,N_6300,N_5667);
nor U10787 (N_10787,N_9503,N_9995);
nor U10788 (N_10788,N_5474,N_7013);
nor U10789 (N_10789,N_6781,N_8865);
xnor U10790 (N_10790,N_6108,N_8528);
xor U10791 (N_10791,N_5366,N_9683);
nand U10792 (N_10792,N_5942,N_8890);
and U10793 (N_10793,N_5708,N_7966);
xnor U10794 (N_10794,N_6537,N_9095);
or U10795 (N_10795,N_7372,N_8572);
or U10796 (N_10796,N_5967,N_8188);
or U10797 (N_10797,N_9626,N_9253);
nand U10798 (N_10798,N_7166,N_7027);
or U10799 (N_10799,N_6429,N_7423);
and U10800 (N_10800,N_9896,N_5926);
or U10801 (N_10801,N_5586,N_6222);
nand U10802 (N_10802,N_5738,N_8973);
nand U10803 (N_10803,N_9341,N_6709);
and U10804 (N_10804,N_8734,N_5254);
xnor U10805 (N_10805,N_9402,N_6779);
nand U10806 (N_10806,N_8195,N_9725);
nor U10807 (N_10807,N_6889,N_8846);
xor U10808 (N_10808,N_5438,N_5303);
xor U10809 (N_10809,N_7975,N_9563);
and U10810 (N_10810,N_9883,N_9478);
or U10811 (N_10811,N_9770,N_9537);
nor U10812 (N_10812,N_6103,N_9734);
or U10813 (N_10813,N_5335,N_7576);
nand U10814 (N_10814,N_9300,N_9980);
or U10815 (N_10815,N_7908,N_9203);
nor U10816 (N_10816,N_6275,N_6711);
and U10817 (N_10817,N_6144,N_7619);
nand U10818 (N_10818,N_5863,N_8838);
and U10819 (N_10819,N_8117,N_5981);
nand U10820 (N_10820,N_7237,N_5354);
and U10821 (N_10821,N_8518,N_5616);
or U10822 (N_10822,N_7779,N_9204);
nor U10823 (N_10823,N_9294,N_9072);
or U10824 (N_10824,N_5319,N_5729);
nand U10825 (N_10825,N_9071,N_7348);
or U10826 (N_10826,N_6770,N_6655);
nand U10827 (N_10827,N_8276,N_9871);
or U10828 (N_10828,N_6430,N_9039);
nor U10829 (N_10829,N_7816,N_6928);
and U10830 (N_10830,N_6597,N_6639);
xor U10831 (N_10831,N_5001,N_6390);
or U10832 (N_10832,N_5984,N_6380);
xnor U10833 (N_10833,N_5481,N_5825);
and U10834 (N_10834,N_6202,N_6841);
nand U10835 (N_10835,N_9704,N_8888);
and U10836 (N_10836,N_7173,N_9450);
and U10837 (N_10837,N_5838,N_7362);
xor U10838 (N_10838,N_9112,N_6428);
nand U10839 (N_10839,N_7497,N_8891);
xnor U10840 (N_10840,N_6917,N_9312);
and U10841 (N_10841,N_7145,N_9321);
nor U10842 (N_10842,N_7771,N_6844);
nand U10843 (N_10843,N_5245,N_9078);
xnor U10844 (N_10844,N_7380,N_8354);
xor U10845 (N_10845,N_9801,N_9445);
or U10846 (N_10846,N_9643,N_8457);
and U10847 (N_10847,N_8129,N_8692);
and U10848 (N_10848,N_9954,N_7732);
and U10849 (N_10849,N_6132,N_9482);
and U10850 (N_10850,N_7346,N_9124);
or U10851 (N_10851,N_7652,N_8157);
nand U10852 (N_10852,N_6355,N_7152);
nand U10853 (N_10853,N_6771,N_9604);
or U10854 (N_10854,N_6067,N_8863);
nand U10855 (N_10855,N_7519,N_8611);
and U10856 (N_10856,N_7428,N_5664);
or U10857 (N_10857,N_7555,N_7099);
xor U10858 (N_10858,N_8297,N_5940);
nand U10859 (N_10859,N_9463,N_9461);
and U10860 (N_10860,N_5471,N_6738);
and U10861 (N_10861,N_5542,N_6609);
or U10862 (N_10862,N_8413,N_9367);
xnor U10863 (N_10863,N_7489,N_6124);
nor U10864 (N_10864,N_9396,N_7382);
xnor U10865 (N_10865,N_7131,N_9119);
or U10866 (N_10866,N_6366,N_6812);
nor U10867 (N_10867,N_5884,N_5931);
and U10868 (N_10868,N_5857,N_6130);
nand U10869 (N_10869,N_9529,N_8777);
nor U10870 (N_10870,N_7475,N_8763);
xor U10871 (N_10871,N_8994,N_6326);
nor U10872 (N_10872,N_8311,N_5211);
nand U10873 (N_10873,N_6036,N_5742);
and U10874 (N_10874,N_5676,N_9539);
or U10875 (N_10875,N_5075,N_5396);
nand U10876 (N_10876,N_9710,N_7398);
xor U10877 (N_10877,N_5459,N_7653);
nand U10878 (N_10878,N_8669,N_6538);
nor U10879 (N_10879,N_7903,N_9760);
nor U10880 (N_10880,N_5870,N_8667);
nor U10881 (N_10881,N_7009,N_6383);
nand U10882 (N_10882,N_6670,N_5021);
xor U10883 (N_10883,N_9132,N_8255);
nor U10884 (N_10884,N_5219,N_8226);
nor U10885 (N_10885,N_9809,N_6215);
nand U10886 (N_10886,N_9285,N_7883);
and U10887 (N_10887,N_6565,N_9098);
nand U10888 (N_10888,N_8702,N_7746);
nand U10889 (N_10889,N_6071,N_6338);
xor U10890 (N_10890,N_9964,N_8016);
xnor U10891 (N_10891,N_7174,N_8811);
or U10892 (N_10892,N_7293,N_8238);
nor U10893 (N_10893,N_9951,N_5993);
xor U10894 (N_10894,N_7546,N_9920);
nor U10895 (N_10895,N_9069,N_6413);
and U10896 (N_10896,N_8566,N_7210);
or U10897 (N_10897,N_6568,N_8314);
xor U10898 (N_10898,N_8961,N_9262);
nand U10899 (N_10899,N_7474,N_6456);
xnor U10900 (N_10900,N_5946,N_9689);
nor U10901 (N_10901,N_6118,N_5090);
or U10902 (N_10902,N_8794,N_7859);
xor U10903 (N_10903,N_9581,N_7226);
xor U10904 (N_10904,N_8164,N_6522);
nor U10905 (N_10905,N_6087,N_7310);
nand U10906 (N_10906,N_5581,N_9507);
xor U10907 (N_10907,N_5900,N_6863);
nand U10908 (N_10908,N_7874,N_9595);
nor U10909 (N_10909,N_7494,N_5056);
nand U10910 (N_10910,N_5246,N_6955);
and U10911 (N_10911,N_9838,N_9184);
or U10912 (N_10912,N_8958,N_8701);
nand U10913 (N_10913,N_7439,N_8087);
xnor U10914 (N_10914,N_6365,N_5344);
and U10915 (N_10915,N_5161,N_5391);
xnor U10916 (N_10916,N_5488,N_5323);
nor U10917 (N_10917,N_5322,N_7002);
nor U10918 (N_10918,N_9850,N_6728);
or U10919 (N_10919,N_8064,N_6204);
nand U10920 (N_10920,N_9749,N_9547);
nor U10921 (N_10921,N_8414,N_7787);
xor U10922 (N_10922,N_9480,N_6107);
xnor U10923 (N_10923,N_8011,N_8449);
nor U10924 (N_10924,N_6583,N_8519);
or U10925 (N_10925,N_7435,N_7785);
nor U10926 (N_10926,N_7160,N_5450);
and U10927 (N_10927,N_9015,N_7239);
nand U10928 (N_10928,N_5613,N_5174);
and U10929 (N_10929,N_9269,N_6853);
xor U10930 (N_10930,N_5134,N_8635);
nor U10931 (N_10931,N_7389,N_5386);
xor U10932 (N_10932,N_9984,N_8786);
nor U10933 (N_10933,N_9251,N_9832);
nor U10934 (N_10934,N_8984,N_6412);
and U10935 (N_10935,N_5735,N_7934);
or U10936 (N_10936,N_9049,N_7756);
xnor U10937 (N_10937,N_8008,N_9370);
and U10938 (N_10938,N_7281,N_7229);
or U10939 (N_10939,N_8813,N_5636);
and U10940 (N_10940,N_5097,N_9177);
xnor U10941 (N_10941,N_7834,N_6612);
nand U10942 (N_10942,N_6860,N_5458);
or U10943 (N_10943,N_5491,N_8948);
nand U10944 (N_10944,N_6721,N_5378);
nor U10945 (N_10945,N_6987,N_7650);
or U10946 (N_10946,N_9245,N_6870);
nor U10947 (N_10947,N_7664,N_6778);
nand U10948 (N_10948,N_8500,N_7285);
xor U10949 (N_10949,N_7418,N_5132);
xor U10950 (N_10950,N_6852,N_7259);
and U10951 (N_10951,N_6876,N_6943);
and U10952 (N_10952,N_6359,N_8710);
and U10953 (N_10953,N_8932,N_5158);
and U10954 (N_10954,N_6925,N_5921);
or U10955 (N_10955,N_5962,N_9101);
xor U10956 (N_10956,N_7954,N_7378);
nor U10957 (N_10957,N_9062,N_9385);
or U10958 (N_10958,N_7450,N_6443);
nand U10959 (N_10959,N_8835,N_6014);
xor U10960 (N_10960,N_8570,N_9316);
xnor U10961 (N_10961,N_9076,N_9440);
nor U10962 (N_10962,N_6936,N_9876);
or U10963 (N_10963,N_6862,N_9538);
nand U10964 (N_10964,N_7121,N_7778);
nor U10965 (N_10965,N_8858,N_7493);
nor U10966 (N_10966,N_6828,N_8232);
nor U10967 (N_10967,N_8899,N_7370);
nor U10968 (N_10968,N_5604,N_8300);
xor U10969 (N_10969,N_6506,N_8010);
nor U10970 (N_10970,N_9996,N_9968);
nor U10971 (N_10971,N_6057,N_8320);
nand U10972 (N_10972,N_7710,N_5728);
nor U10973 (N_10973,N_7988,N_8782);
nor U10974 (N_10974,N_9239,N_7488);
nand U10975 (N_10975,N_6650,N_9532);
or U10976 (N_10976,N_8366,N_9231);
and U10977 (N_10977,N_7831,N_5772);
xnor U10978 (N_10978,N_7449,N_5554);
and U10979 (N_10979,N_8798,N_7938);
nor U10980 (N_10980,N_6096,N_5412);
and U10981 (N_10981,N_8371,N_9598);
nand U10982 (N_10982,N_8479,N_8936);
and U10983 (N_10983,N_9874,N_8832);
or U10984 (N_10984,N_9089,N_6131);
nand U10985 (N_10985,N_8358,N_8363);
nor U10986 (N_10986,N_8627,N_5073);
nand U10987 (N_10987,N_5563,N_5876);
nor U10988 (N_10988,N_9360,N_9464);
nand U10989 (N_10989,N_6903,N_8808);
and U10990 (N_10990,N_8395,N_8504);
or U10991 (N_10991,N_7197,N_7109);
nand U10992 (N_10992,N_7780,N_5210);
or U10993 (N_10993,N_7061,N_7607);
xnor U10994 (N_10994,N_5363,N_5416);
xnor U10995 (N_10995,N_5599,N_6901);
nor U10996 (N_10996,N_7563,N_5490);
nor U10997 (N_10997,N_6604,N_5072);
xor U10998 (N_10998,N_5739,N_7178);
and U10999 (N_10999,N_8273,N_9488);
or U11000 (N_11000,N_8350,N_6866);
nand U11001 (N_11001,N_7945,N_7671);
nand U11002 (N_11002,N_5846,N_6459);
and U11003 (N_11003,N_7581,N_9207);
nand U11004 (N_11004,N_5081,N_8847);
nand U11005 (N_11005,N_5414,N_7291);
xnor U11006 (N_11006,N_8030,N_6623);
nor U11007 (N_11007,N_6244,N_8508);
nand U11008 (N_11008,N_7789,N_7602);
nand U11009 (N_11009,N_9848,N_5368);
and U11010 (N_11010,N_7529,N_8344);
nand U11011 (N_11011,N_9153,N_7316);
nor U11012 (N_11012,N_8704,N_9727);
or U11013 (N_11013,N_5077,N_6221);
xnor U11014 (N_11014,N_9646,N_5495);
xor U11015 (N_11015,N_8376,N_7524);
and U11016 (N_11016,N_5802,N_7344);
nand U11017 (N_11017,N_6492,N_6705);
and U11018 (N_11018,N_5199,N_6545);
nor U11019 (N_11019,N_8006,N_8718);
nor U11020 (N_11020,N_9624,N_5515);
or U11021 (N_11021,N_7095,N_7421);
or U11022 (N_11022,N_6957,N_7092);
and U11023 (N_11023,N_7149,N_9918);
nor U11024 (N_11024,N_5779,N_8047);
nor U11025 (N_11025,N_7278,N_8628);
or U11026 (N_11026,N_5638,N_7481);
and U11027 (N_11027,N_5204,N_6610);
and U11028 (N_11028,N_8105,N_9820);
nor U11029 (N_11029,N_7041,N_8909);
nand U11030 (N_11030,N_8241,N_7248);
xor U11031 (N_11031,N_8058,N_8256);
or U11032 (N_11032,N_7797,N_8285);
xor U11033 (N_11033,N_8469,N_5406);
and U11034 (N_11034,N_6052,N_8448);
or U11035 (N_11035,N_5123,N_5830);
xnor U11036 (N_11036,N_9971,N_7709);
xnor U11037 (N_11037,N_9214,N_9796);
nand U11038 (N_11038,N_6745,N_6884);
nand U11039 (N_11039,N_6898,N_5098);
and U11040 (N_11040,N_7885,N_9869);
or U11041 (N_11041,N_5827,N_7238);
and U11042 (N_11042,N_8186,N_6063);
nor U11043 (N_11043,N_8778,N_5932);
nand U11044 (N_11044,N_8560,N_9991);
xor U11045 (N_11045,N_8031,N_8341);
nor U11046 (N_11046,N_8456,N_8330);
nor U11047 (N_11047,N_7503,N_5347);
nand U11048 (N_11048,N_7794,N_9771);
or U11049 (N_11049,N_7441,N_6700);
or U11050 (N_11050,N_9768,N_6940);
nand U11051 (N_11051,N_6349,N_6358);
and U11052 (N_11052,N_7567,N_9060);
nor U11053 (N_11053,N_7965,N_8493);
nor U11054 (N_11054,N_6872,N_8665);
nand U11055 (N_11055,N_6348,N_6753);
or U11056 (N_11056,N_6333,N_6782);
xnor U11057 (N_11057,N_5964,N_6990);
xnor U11058 (N_11058,N_5583,N_6970);
xnor U11059 (N_11059,N_9409,N_9774);
nor U11060 (N_11060,N_9425,N_7941);
xnor U11061 (N_11061,N_7682,N_5099);
and U11062 (N_11062,N_9860,N_5093);
nor U11063 (N_11063,N_8061,N_9933);
nand U11064 (N_11064,N_7614,N_9810);
or U11065 (N_11065,N_6388,N_5580);
xnor U11066 (N_11066,N_9258,N_5994);
nor U11067 (N_11067,N_8140,N_8698);
nor U11068 (N_11068,N_8068,N_5971);
and U11069 (N_11069,N_7535,N_5642);
xor U11070 (N_11070,N_7396,N_5596);
nand U11071 (N_11071,N_8090,N_7722);
nand U11072 (N_11072,N_9934,N_5436);
and U11073 (N_11073,N_9424,N_9141);
nand U11074 (N_11074,N_8460,N_5678);
nand U11075 (N_11075,N_5880,N_9056);
nand U11076 (N_11076,N_9892,N_8615);
nor U11077 (N_11077,N_5837,N_7658);
and U11078 (N_11078,N_9880,N_6488);
xnor U11079 (N_11079,N_8645,N_8037);
nand U11080 (N_11080,N_7462,N_5853);
nor U11081 (N_11081,N_5671,N_8599);
nor U11082 (N_11082,N_5847,N_6719);
xnor U11083 (N_11083,N_9365,N_9872);
or U11084 (N_11084,N_7821,N_8564);
xnor U11085 (N_11085,N_9708,N_9764);
nor U11086 (N_11086,N_5377,N_8141);
xnor U11087 (N_11087,N_5047,N_9530);
nand U11088 (N_11088,N_7049,N_9542);
nand U11089 (N_11089,N_7071,N_6791);
and U11090 (N_11090,N_5275,N_6907);
or U11091 (N_11091,N_9997,N_7598);
nand U11092 (N_11092,N_8176,N_7062);
xor U11093 (N_11093,N_7551,N_7838);
xor U11094 (N_11094,N_6414,N_6614);
xnor U11095 (N_11095,N_5284,N_5968);
or U11096 (N_11096,N_8441,N_8298);
xor U11097 (N_11097,N_8076,N_5584);
or U11098 (N_11098,N_6550,N_9946);
and U11099 (N_11099,N_8179,N_9325);
nand U11100 (N_11100,N_6214,N_6571);
nor U11101 (N_11101,N_8661,N_9468);
nor U11102 (N_11102,N_9457,N_8633);
and U11103 (N_11103,N_8729,N_6780);
nor U11104 (N_11104,N_8249,N_9485);
nand U11105 (N_11105,N_8515,N_9011);
or U11106 (N_11106,N_9492,N_6931);
and U11107 (N_11107,N_5004,N_8712);
nand U11108 (N_11108,N_6010,N_7368);
and U11109 (N_11109,N_9584,N_6920);
xnor U11110 (N_11110,N_9821,N_8079);
nand U11111 (N_11111,N_6277,N_9426);
xor U11112 (N_11112,N_5154,N_5195);
nand U11113 (N_11113,N_8929,N_5532);
xor U11114 (N_11114,N_5710,N_6724);
and U11115 (N_11115,N_9660,N_8639);
nor U11116 (N_11116,N_7206,N_9423);
or U11117 (N_11117,N_5998,N_6895);
or U11118 (N_11118,N_9264,N_7115);
and U11119 (N_11119,N_5494,N_7916);
xnor U11120 (N_11120,N_9549,N_6255);
and U11121 (N_11121,N_5991,N_7974);
xnor U11122 (N_11122,N_7343,N_8194);
and U11123 (N_11123,N_9572,N_7484);
or U11124 (N_11124,N_5186,N_9144);
or U11125 (N_11125,N_7035,N_7628);
nor U11126 (N_11126,N_6651,N_8820);
or U11127 (N_11127,N_7552,N_5487);
nor U11128 (N_11128,N_6966,N_5615);
xnor U11129 (N_11129,N_6256,N_7580);
nand U11130 (N_11130,N_8419,N_5452);
or U11131 (N_11131,N_5342,N_9087);
nor U11132 (N_11132,N_5805,N_6317);
and U11133 (N_11133,N_6068,N_9673);
nand U11134 (N_11134,N_9221,N_6247);
and U11135 (N_11135,N_6861,N_6873);
xor U11136 (N_11136,N_8073,N_9386);
xnor U11137 (N_11137,N_5622,N_9407);
xor U11138 (N_11138,N_6151,N_6527);
xnor U11139 (N_11139,N_7545,N_5274);
and U11140 (N_11140,N_8850,N_9082);
nand U11141 (N_11141,N_6696,N_6252);
and U11142 (N_11142,N_9739,N_5801);
nand U11143 (N_11143,N_5611,N_7879);
nor U11144 (N_11144,N_6294,N_5892);
xnor U11145 (N_11145,N_7644,N_9698);
xnor U11146 (N_11146,N_5949,N_5910);
nor U11147 (N_11147,N_5798,N_7392);
and U11148 (N_11148,N_6159,N_7927);
and U11149 (N_11149,N_9756,N_5425);
and U11150 (N_11150,N_8018,N_9723);
or U11151 (N_11151,N_8740,N_5654);
nand U11152 (N_11152,N_6616,N_6110);
nand U11153 (N_11153,N_7126,N_5038);
nor U11154 (N_11154,N_8885,N_7272);
or U11155 (N_11155,N_7335,N_6658);
or U11156 (N_11156,N_5277,N_5525);
nand U11157 (N_11157,N_8960,N_5249);
nand U11158 (N_11158,N_7712,N_9650);
nor U11159 (N_11159,N_6304,N_5215);
and U11160 (N_11160,N_9890,N_9021);
or U11161 (N_11161,N_7055,N_5896);
nand U11162 (N_11162,N_6998,N_7707);
and U11163 (N_11163,N_7694,N_9622);
and U11164 (N_11164,N_5790,N_7615);
xnor U11165 (N_11165,N_8556,N_6376);
and U11166 (N_11166,N_7824,N_6543);
xnor U11167 (N_11167,N_7125,N_9315);
nand U11168 (N_11168,N_6075,N_5336);
nand U11169 (N_11169,N_5006,N_6807);
and U11170 (N_11170,N_8368,N_6201);
nor U11171 (N_11171,N_9609,N_5328);
nor U11172 (N_11172,N_7773,N_5894);
nand U11173 (N_11173,N_5485,N_8612);
or U11174 (N_11174,N_6633,N_6644);
nand U11175 (N_11175,N_8279,N_8781);
xnor U11176 (N_11176,N_7390,N_6425);
and U11177 (N_11177,N_9762,N_9938);
xor U11178 (N_11178,N_7365,N_5313);
nor U11179 (N_11179,N_8111,N_5071);
nor U11180 (N_11180,N_9930,N_5697);
or U11181 (N_11181,N_9398,N_8901);
nor U11182 (N_11182,N_7111,N_5408);
and U11183 (N_11183,N_8474,N_6839);
and U11184 (N_11184,N_5221,N_7184);
xnor U11185 (N_11185,N_8542,N_6641);
or U11186 (N_11186,N_8833,N_8654);
and U11187 (N_11187,N_9199,N_9512);
nand U11188 (N_11188,N_6624,N_7811);
xnor U11189 (N_11189,N_8574,N_7786);
and U11190 (N_11190,N_9958,N_9068);
nand U11191 (N_11191,N_7561,N_7260);
nand U11192 (N_11192,N_9885,N_9610);
and U11193 (N_11193,N_8378,N_8137);
nor U11194 (N_11194,N_5163,N_8480);
and U11195 (N_11195,N_6647,N_8754);
nor U11196 (N_11196,N_9746,N_6589);
and U11197 (N_11197,N_6206,N_8217);
xor U11198 (N_11198,N_5527,N_9511);
and U11199 (N_11199,N_6323,N_9299);
nor U11200 (N_11200,N_5914,N_5523);
and U11201 (N_11201,N_8453,N_6267);
nand U11202 (N_11202,N_6360,N_9466);
nand U11203 (N_11203,N_6473,N_5133);
nor U11204 (N_11204,N_5796,N_7057);
and U11205 (N_11205,N_5954,N_9433);
or U11206 (N_11206,N_7880,N_6978);
and U11207 (N_11207,N_6744,N_5592);
or U11208 (N_11208,N_5937,N_8321);
and U11209 (N_11209,N_7100,N_6441);
nand U11210 (N_11210,N_6556,N_8156);
and U11211 (N_11211,N_6544,N_9417);
xor U11212 (N_11212,N_9109,N_5799);
nand U11213 (N_11213,N_6497,N_7813);
or U11214 (N_11214,N_6684,N_9111);
xor U11215 (N_11215,N_6289,N_9909);
or U11216 (N_11216,N_5537,N_9179);
nor U11217 (N_11217,N_5078,N_7715);
and U11218 (N_11218,N_7463,N_5793);
xor U11219 (N_11219,N_8138,N_7659);
or U11220 (N_11220,N_9669,N_9897);
or U11221 (N_11221,N_7429,N_8328);
nand U11222 (N_11222,N_6555,N_6362);
or U11223 (N_11223,N_8342,N_5508);
nand U11224 (N_11224,N_9040,N_7436);
nor U11225 (N_11225,N_9747,N_5747);
xnor U11226 (N_11226,N_8930,N_5744);
xor U11227 (N_11227,N_5145,N_7743);
and U11228 (N_11228,N_9241,N_7587);
nand U11229 (N_11229,N_9031,N_5612);
xnor U11230 (N_11230,N_9524,N_5776);
or U11231 (N_11231,N_5717,N_7526);
and U11232 (N_11232,N_7320,N_6161);
nand U11233 (N_11233,N_6112,N_9992);
nor U11234 (N_11234,N_8976,N_7263);
and U11235 (N_11235,N_7384,N_9006);
or U11236 (N_11236,N_7299,N_9737);
nand U11237 (N_11237,N_9629,N_9769);
xnor U11238 (N_11238,N_9694,N_7072);
nor U11239 (N_11239,N_9540,N_5143);
and U11240 (N_11240,N_6755,N_6171);
xor U11241 (N_11241,N_5901,N_5553);
nand U11242 (N_11242,N_7539,N_8252);
nand U11243 (N_11243,N_8594,N_5854);
nor U11244 (N_11244,N_7161,N_5757);
nor U11245 (N_11245,N_8027,N_6493);
nor U11246 (N_11246,N_6587,N_5400);
nand U11247 (N_11247,N_7956,N_8082);
or U11248 (N_11248,N_5208,N_7074);
xor U11249 (N_11249,N_6769,N_6708);
nor U11250 (N_11250,N_7381,N_7325);
and U11251 (N_11251,N_7782,N_9397);
or U11252 (N_11252,N_5216,N_8876);
and U11253 (N_11253,N_7303,N_9815);
nor U11254 (N_11254,N_5904,N_9663);
nand U11255 (N_11255,N_7808,N_7764);
or U11256 (N_11256,N_8801,N_5541);
nand U11257 (N_11257,N_6795,N_5393);
xnor U11258 (N_11258,N_6762,N_5448);
nand U11259 (N_11259,N_6378,N_7801);
nand U11260 (N_11260,N_8647,N_6266);
nor U11261 (N_11261,N_5951,N_8397);
or U11262 (N_11262,N_9118,N_5083);
and U11263 (N_11263,N_5561,N_6569);
nor U11264 (N_11264,N_5690,N_5175);
and U11265 (N_11265,N_8071,N_8347);
nor U11266 (N_11266,N_8987,N_5952);
or U11267 (N_11267,N_7427,N_8902);
or U11268 (N_11268,N_5886,N_7213);
nor U11269 (N_11269,N_7287,N_6020);
or U11270 (N_11270,N_9840,N_6341);
nand U11271 (N_11271,N_5052,N_9889);
nor U11272 (N_11272,N_8287,N_5916);
nor U11273 (N_11273,N_7465,N_7992);
and U11274 (N_11274,N_7089,N_8296);
nor U11275 (N_11275,N_5168,N_9350);
and U11276 (N_11276,N_8383,N_6581);
and U11277 (N_11277,N_8824,N_5818);
and U11278 (N_11278,N_8092,N_9548);
and U11279 (N_11279,N_5415,N_7134);
and U11280 (N_11280,N_6227,N_6357);
or U11281 (N_11281,N_6179,N_6573);
or U11282 (N_11282,N_9430,N_9568);
and U11283 (N_11283,N_5384,N_8900);
nand U11284 (N_11284,N_7138,N_9138);
nor U11285 (N_11285,N_8335,N_7353);
or U11286 (N_11286,N_5877,N_9826);
or U11287 (N_11287,N_8872,N_7007);
or U11288 (N_11288,N_8586,N_9513);
nand U11289 (N_11289,N_7444,N_8351);
and U11290 (N_11290,N_6054,N_7070);
or U11291 (N_11291,N_7112,N_5712);
or U11292 (N_11292,N_7720,N_9053);
nand U11293 (N_11293,N_6748,N_7034);
or U11294 (N_11294,N_8968,N_9577);
xnor U11295 (N_11295,N_6398,N_9084);
and U11296 (N_11296,N_9180,N_6123);
nand U11297 (N_11297,N_7107,N_7590);
and U11298 (N_11298,N_7646,N_5941);
and U11299 (N_11299,N_5997,N_6037);
and U11300 (N_11300,N_9281,N_9659);
nand U11301 (N_11301,N_6620,N_5828);
nand U11302 (N_11302,N_5351,N_6763);
or U11303 (N_11303,N_6959,N_9354);
nand U11304 (N_11304,N_5180,N_8390);
or U11305 (N_11305,N_5557,N_8213);
xor U11306 (N_11306,N_5944,N_8365);
and U11307 (N_11307,N_6386,N_5268);
or U11308 (N_11308,N_9010,N_9590);
or U11309 (N_11309,N_8589,N_7150);
or U11310 (N_11310,N_8737,N_7351);
or U11311 (N_11311,N_6264,N_8881);
nor U11312 (N_11312,N_5139,N_6242);
and U11313 (N_11313,N_5030,N_6028);
xnor U11314 (N_11314,N_5334,N_9534);
nor U11315 (N_11315,N_5522,N_5961);
nand U11316 (N_11316,N_7719,N_6663);
nor U11317 (N_11317,N_5727,N_8196);
xor U11318 (N_11318,N_8158,N_9303);
nor U11319 (N_11319,N_8430,N_7102);
nand U11320 (N_11320,N_9453,N_9228);
and U11321 (N_11321,N_7393,N_9065);
xnor U11322 (N_11322,N_8679,N_7997);
nand U11323 (N_11323,N_5627,N_7640);
and U11324 (N_11324,N_9526,N_7504);
nand U11325 (N_11325,N_6013,N_7585);
xnor U11326 (N_11326,N_8418,N_9438);
nor U11327 (N_11327,N_8440,N_7257);
nand U11328 (N_11328,N_9636,N_8225);
nor U11329 (N_11329,N_8005,N_9172);
and U11330 (N_11330,N_7457,N_5791);
or U11331 (N_11331,N_6019,N_6758);
nor U11332 (N_11332,N_7898,N_8903);
nor U11333 (N_11333,N_8499,N_5724);
or U11334 (N_11334,N_9304,N_8507);
xor U11335 (N_11335,N_7673,N_5263);
or U11336 (N_11336,N_9037,N_7736);
nand U11337 (N_11337,N_7082,N_7168);
nor U11338 (N_11338,N_8275,N_8995);
or U11339 (N_11339,N_9400,N_7717);
xnor U11340 (N_11340,N_5551,N_5766);
or U11341 (N_11341,N_6183,N_7046);
or U11342 (N_11342,N_7688,N_8245);
or U11343 (N_11343,N_5588,N_9305);
nor U11344 (N_11344,N_9514,N_6631);
and U11345 (N_11345,N_9075,N_8265);
xor U11346 (N_11346,N_9775,N_8203);
or U11347 (N_11347,N_7326,N_9346);
nand U11348 (N_11348,N_5826,N_7053);
nand U11349 (N_11349,N_7419,N_6760);
nand U11350 (N_11350,N_8513,N_7286);
or U11351 (N_11351,N_8907,N_5042);
and U11352 (N_11352,N_5634,N_6156);
and U11353 (N_11353,N_9244,N_5519);
xor U11354 (N_11354,N_6283,N_9875);
nand U11355 (N_11355,N_8802,N_8086);
and U11356 (N_11356,N_7011,N_8216);
and U11357 (N_11357,N_8656,N_9108);
xnor U11358 (N_11358,N_8402,N_7322);
and U11359 (N_11359,N_9814,N_8389);
nor U11360 (N_11360,N_6299,N_9117);
xnor U11361 (N_11361,N_6149,N_5141);
or U11362 (N_11362,N_6315,N_9578);
xor U11363 (N_11363,N_6974,N_5635);
nand U11364 (N_11364,N_6334,N_9013);
nor U11365 (N_11365,N_6680,N_5142);
nor U11366 (N_11366,N_7369,N_6313);
nor U11367 (N_11367,N_8316,N_7411);
and U11368 (N_11368,N_8879,N_7629);
nand U11369 (N_11369,N_5626,N_8377);
xnor U11370 (N_11370,N_7792,N_7199);
and U11371 (N_11371,N_9977,N_9163);
or U11372 (N_11372,N_8109,N_5577);
nand U11373 (N_11373,N_6002,N_7999);
xor U11374 (N_11374,N_9161,N_8028);
and U11375 (N_11375,N_5835,N_6152);
nand U11376 (N_11376,N_6526,N_8036);
or U11377 (N_11377,N_9735,N_9743);
nor U11378 (N_11378,N_9754,N_5111);
xor U11379 (N_11379,N_9726,N_5234);
or U11380 (N_11380,N_9364,N_9474);
and U11381 (N_11381,N_8526,N_8841);
and U11382 (N_11382,N_5392,N_9783);
nand U11383 (N_11383,N_7185,N_8975);
or U11384 (N_11384,N_7473,N_7375);
and U11385 (N_11385,N_7406,N_8166);
nor U11386 (N_11386,N_9608,N_7798);
nor U11387 (N_11387,N_8817,N_5741);
nand U11388 (N_11388,N_6766,N_6373);
nand U11389 (N_11389,N_9077,N_7443);
nor U11390 (N_11390,N_6480,N_9678);
or U11391 (N_11391,N_6465,N_9185);
and U11392 (N_11392,N_5048,N_6858);
xor U11393 (N_11393,N_6503,N_7003);
xnor U11394 (N_11394,N_8258,N_6174);
or U11395 (N_11395,N_6452,N_7698);
or U11396 (N_11396,N_9340,N_8538);
or U11397 (N_11397,N_6690,N_9497);
nand U11398 (N_11398,N_7201,N_9867);
or U11399 (N_11399,N_8792,N_7850);
or U11400 (N_11400,N_9002,N_8242);
nand U11401 (N_11401,N_7165,N_8510);
or U11402 (N_11402,N_5371,N_6074);
nand U11403 (N_11403,N_8459,N_8084);
xnor U11404 (N_11404,N_8153,N_8260);
nand U11405 (N_11405,N_9351,N_7895);
xor U11406 (N_11406,N_5630,N_8003);
xor U11407 (N_11407,N_7890,N_5401);
nand U11408 (N_11408,N_8381,N_7385);
nand U11409 (N_11409,N_8175,N_9390);
and U11410 (N_11410,N_8677,N_5700);
nor U11411 (N_11411,N_9339,N_7514);
nand U11412 (N_11412,N_7564,N_7553);
and U11413 (N_11413,N_7487,N_6239);
and U11414 (N_11414,N_5593,N_7774);
or U11415 (N_11415,N_7332,N_7288);
nor U11416 (N_11416,N_5253,N_8927);
nor U11417 (N_11417,N_8042,N_8732);
or U11418 (N_11418,N_8100,N_9044);
nand U11419 (N_11419,N_7085,N_7296);
nor U11420 (N_11420,N_9047,N_5885);
xnor U11421 (N_11421,N_8214,N_5719);
nand U11422 (N_11422,N_8568,N_9580);
nor U11423 (N_11423,N_7846,N_5899);
nor U11424 (N_11424,N_7379,N_8039);
nand U11425 (N_11425,N_5427,N_9631);
and U11426 (N_11426,N_9048,N_6435);
and U11427 (N_11427,N_6843,N_9784);
xor U11428 (N_11428,N_7059,N_8590);
or U11429 (N_11429,N_5231,N_9288);
or U11430 (N_11430,N_9395,N_7499);
or U11431 (N_11431,N_8197,N_9436);
or U11432 (N_11432,N_7977,N_5873);
xnor U11433 (N_11433,N_8154,N_7994);
xnor U11434 (N_11434,N_8990,N_9965);
xor U11435 (N_11435,N_9159,N_8608);
xor U11436 (N_11436,N_6646,N_9956);
nand U11437 (N_11437,N_9634,N_7242);
and U11438 (N_11438,N_6761,N_5600);
xnor U11439 (N_11439,N_8788,N_6816);
xnor U11440 (N_11440,N_9465,N_9323);
nor U11441 (N_11441,N_9676,N_6618);
and U11442 (N_11442,N_6371,N_7665);
and U11443 (N_11443,N_7892,N_6588);
nand U11444 (N_11444,N_5947,N_8035);
nand U11445 (N_11445,N_5280,N_6995);
nor U11446 (N_11446,N_9987,N_6560);
nor U11447 (N_11447,N_6211,N_5015);
nand U11448 (N_11448,N_7894,N_9043);
or U11449 (N_11449,N_5314,N_6170);
nor U11450 (N_11450,N_9943,N_6158);
nand U11451 (N_11451,N_6448,N_5372);
or U11452 (N_11452,N_9128,N_8641);
and U11453 (N_11453,N_7601,N_8595);
or U11454 (N_11454,N_5768,N_5923);
xor U11455 (N_11455,N_6402,N_5666);
xnor U11456 (N_11456,N_8660,N_6474);
and U11457 (N_11457,N_8988,N_6938);
nor U11458 (N_11458,N_5403,N_8596);
nor U11459 (N_11459,N_5359,N_9522);
xnor U11460 (N_11460,N_7214,N_8747);
or U11461 (N_11461,N_5420,N_6128);
or U11462 (N_11462,N_7302,N_7096);
or U11463 (N_11463,N_8892,N_5159);
nand U11464 (N_11464,N_8529,N_5777);
nand U11465 (N_11465,N_5927,N_7495);
nand U11466 (N_11466,N_8412,N_7884);
xor U11467 (N_11467,N_7235,N_8024);
nor U11468 (N_11468,N_6322,N_5785);
nand U11469 (N_11469,N_9357,N_7845);
or U11470 (N_11470,N_9825,N_9571);
or U11471 (N_11471,N_8842,N_8065);
nand U11472 (N_11472,N_7680,N_6933);
nand U11473 (N_11473,N_9561,N_5536);
nor U11474 (N_11474,N_6921,N_8691);
xnor U11475 (N_11475,N_8466,N_7048);
nor U11476 (N_11476,N_6136,N_9494);
and U11477 (N_11477,N_9523,N_7319);
nor U11478 (N_11478,N_6848,N_9116);
nor U11479 (N_11479,N_8928,N_8577);
or U11480 (N_11480,N_5867,N_7525);
nand U11481 (N_11481,N_5758,N_9961);
nor U11482 (N_11482,N_5294,N_5040);
nand U11483 (N_11483,N_5864,N_9088);
or U11484 (N_11484,N_9405,N_8619);
nor U11485 (N_11485,N_8112,N_8182);
and U11486 (N_11486,N_9491,N_6416);
and U11487 (N_11487,N_9419,N_7114);
or U11488 (N_11488,N_5709,N_5169);
xnor U11489 (N_11489,N_7624,N_6746);
nor U11490 (N_11490,N_7403,N_7620);
nor U11491 (N_11491,N_9256,N_9202);
and U11492 (N_11492,N_5672,N_9046);
xor U11493 (N_11493,N_9836,N_9613);
or U11494 (N_11494,N_9518,N_9612);
or U11495 (N_11495,N_5943,N_6584);
and U11496 (N_11496,N_6883,N_8730);
nand U11497 (N_11497,N_8416,N_8359);
and U11498 (N_11498,N_7266,N_6101);
or U11499 (N_11499,N_7625,N_5155);
nand U11500 (N_11500,N_7029,N_7623);
xnor U11501 (N_11501,N_5619,N_5118);
nor U11502 (N_11502,N_8673,N_8442);
or U11503 (N_11503,N_9767,N_7957);
and U11504 (N_11504,N_5856,N_7243);
xnor U11505 (N_11505,N_6837,N_9428);
or U11506 (N_11506,N_7268,N_6507);
or U11507 (N_11507,N_7410,N_7527);
or U11508 (N_11508,N_5271,N_6046);
nand U11509 (N_11509,N_8859,N_5691);
and U11510 (N_11510,N_8849,N_7039);
nor U11511 (N_11511,N_8444,N_9248);
or U11512 (N_11512,N_8017,N_5218);
nand U11513 (N_11513,N_8578,N_6874);
xnor U11514 (N_11514,N_6449,N_6531);
xor U11515 (N_11515,N_5128,N_6523);
or U11516 (N_11516,N_9280,N_6657);
xor U11517 (N_11517,N_7424,N_6467);
or U11518 (N_11518,N_8634,N_5974);
xor U11519 (N_11519,N_6856,N_8063);
and U11520 (N_11520,N_6835,N_7407);
nand U11521 (N_11521,N_8675,N_5824);
xor U11522 (N_11522,N_9579,N_8133);
and U11523 (N_11523,N_9978,N_5305);
xnor U11524 (N_11524,N_7067,N_6687);
xor U11525 (N_11525,N_8614,N_5804);
xnor U11526 (N_11526,N_9266,N_6806);
and U11527 (N_11527,N_9475,N_8247);
and U11528 (N_11528,N_9515,N_7621);
xnor U11529 (N_11529,N_6984,N_8348);
and U11530 (N_11530,N_7451,N_7476);
xnor U11531 (N_11531,N_5762,N_7768);
or U11532 (N_11532,N_6932,N_7212);
and U11533 (N_11533,N_6590,N_9045);
and U11534 (N_11534,N_6015,N_7528);
nor U11535 (N_11535,N_8404,N_9535);
or U11536 (N_11536,N_6603,N_6309);
or U11537 (N_11537,N_9982,N_7307);
nor U11538 (N_11538,N_5116,N_5929);
xor U11539 (N_11539,N_8387,N_7486);
or U11540 (N_11540,N_5887,N_6941);
nand U11541 (N_11541,N_6079,N_5027);
xor U11542 (N_11542,N_7016,N_6484);
and U11543 (N_11543,N_8657,N_9945);
nor U11544 (N_11544,N_9408,N_9470);
nor U11545 (N_11545,N_5679,N_8951);
or U11546 (N_11546,N_7502,N_8557);
xor U11547 (N_11547,N_8573,N_8609);
nand U11548 (N_11548,N_7980,N_9824);
or U11549 (N_11549,N_6001,N_9675);
or U11550 (N_11550,N_6973,N_9973);
nor U11551 (N_11551,N_8310,N_7318);
nand U11552 (N_11552,N_7897,N_5470);
nand U11553 (N_11553,N_8562,N_5722);
xnor U11554 (N_11554,N_8809,N_9134);
or U11555 (N_11555,N_7701,N_5307);
or U11556 (N_11556,N_5771,N_7120);
nor U11557 (N_11557,N_7616,N_5849);
nor U11558 (N_11558,N_9802,N_7270);
or U11559 (N_11559,N_5769,N_8972);
and U11560 (N_11560,N_6518,N_5449);
and U11561 (N_11561,N_9908,N_7557);
or U11562 (N_11562,N_7763,N_6469);
or U11563 (N_11563,N_8812,N_6520);
nor U11564 (N_11564,N_9596,N_8127);
and U11565 (N_11565,N_6916,N_8165);
nand U11566 (N_11566,N_8362,N_5140);
xor U11567 (N_11567,N_6407,N_5726);
nor U11568 (N_11568,N_8826,N_7995);
and U11569 (N_11569,N_8821,N_9343);
or U11570 (N_11570,N_8200,N_8041);
and U11571 (N_11571,N_8804,N_9550);
nand U11572 (N_11572,N_8426,N_5130);
nand U11573 (N_11573,N_6271,N_8427);
and U11574 (N_11574,N_6464,N_6923);
nand U11575 (N_11575,N_6880,N_6613);
or U11576 (N_11576,N_8561,N_6847);
and U11577 (N_11577,N_8423,N_7162);
nor U11578 (N_11578,N_5286,N_8262);
xnor U11579 (N_11579,N_9446,N_7275);
and U11580 (N_11580,N_6305,N_6626);
or U11581 (N_11581,N_8219,N_5976);
and U11582 (N_11582,N_5629,N_8592);
nor U11583 (N_11583,N_8629,N_5465);
and U11584 (N_11584,N_7010,N_6741);
and U11585 (N_11585,N_7359,N_8746);
nor U11586 (N_11586,N_6902,N_7875);
or U11587 (N_11587,N_8866,N_8189);
nand U11588 (N_11588,N_7045,N_5287);
nand U11589 (N_11589,N_9882,N_6547);
nand U11590 (N_11590,N_9114,N_6133);
or U11591 (N_11591,N_9635,N_9169);
xor U11592 (N_11592,N_7256,N_8349);
nor U11593 (N_11593,N_9649,N_9276);
or U11594 (N_11594,N_8622,N_9567);
nor U11595 (N_11595,N_6608,N_5157);
xnor U11596 (N_11596,N_9143,N_9210);
nor U11597 (N_11597,N_5507,N_5150);
and U11598 (N_11598,N_9024,N_9387);
nor U11599 (N_11599,N_5108,N_5310);
xor U11600 (N_11600,N_8916,N_5572);
nand U11601 (N_11601,N_9648,N_9255);
nor U11602 (N_11602,N_7187,N_5760);
and U11603 (N_11603,N_9133,N_5767);
or U11604 (N_11604,N_8204,N_7700);
and U11605 (N_11605,N_9067,N_8379);
nor U11606 (N_11606,N_7726,N_6554);
xnor U11607 (N_11607,N_9903,N_8337);
and U11608 (N_11608,N_6337,N_9690);
and U11609 (N_11609,N_8919,N_7516);
xor U11610 (N_11610,N_5095,N_6532);
or U11611 (N_11611,N_9645,N_7153);
xnor U11612 (N_11612,N_9193,N_7559);
xor U11613 (N_11613,N_9605,N_9962);
and U11614 (N_11614,N_7637,N_6797);
or U11615 (N_11615,N_7044,N_8772);
and U11616 (N_11616,N_7541,N_6091);
xnor U11617 (N_11617,N_5057,N_6350);
nor U11618 (N_11618,N_6208,N_8658);
nor U11619 (N_11619,N_8800,N_8725);
nor U11620 (N_11620,N_9090,N_7447);
xor U11621 (N_11621,N_5834,N_7148);
nor U11622 (N_11622,N_5852,N_5950);
xor U11623 (N_11623,N_9242,N_8488);
xor U11624 (N_11624,N_8989,N_6470);
nand U11625 (N_11625,N_7818,N_9788);
xor U11626 (N_11626,N_8749,N_6296);
xnor U11627 (N_11627,N_5533,N_9377);
nand U11628 (N_11628,N_5055,N_6324);
or U11629 (N_11629,N_7088,N_9059);
nor U11630 (N_11630,N_7600,N_6930);
nor U11631 (N_11631,N_8938,N_5009);
and U11632 (N_11632,N_9957,N_6165);
nand U11633 (N_11633,N_6945,N_7744);
or U11634 (N_11634,N_7180,N_7086);
and U11635 (N_11635,N_6217,N_8924);
xor U11636 (N_11636,N_9851,N_6126);
nand U11637 (N_11637,N_7227,N_7155);
nor U11638 (N_11638,N_5350,N_8643);
or U11639 (N_11639,N_7784,N_5088);
xor U11640 (N_11640,N_8884,N_8438);
or U11641 (N_11641,N_5105,N_7677);
and U11642 (N_11642,N_9222,N_6092);
xnor U11643 (N_11643,N_8062,N_7611);
and U11644 (N_11644,N_7271,N_8921);
nor U11645 (N_11645,N_7193,N_6533);
nor U11646 (N_11646,N_6444,N_6707);
and U11647 (N_11647,N_6336,N_6638);
nand U11648 (N_11648,N_8637,N_5774);
or U11649 (N_11649,N_6234,N_8914);
nand U11650 (N_11650,N_8113,N_7836);
nand U11651 (N_11651,N_8353,N_8501);
and U11652 (N_11652,N_5362,N_5844);
xor U11653 (N_11653,N_7040,N_7734);
xnor U11654 (N_11654,N_9843,N_5528);
nor U11655 (N_11655,N_6146,N_5317);
nor U11656 (N_11656,N_9293,N_6419);
nand U11657 (N_11657,N_5127,N_6045);
or U11658 (N_11658,N_6463,N_9373);
xor U11659 (N_11659,N_8161,N_5031);
nand U11660 (N_11660,N_8779,N_7250);
nor U11661 (N_11661,N_8694,N_9765);
or U11662 (N_11662,N_6090,N_5429);
or U11663 (N_11663,N_9284,N_6965);
nor U11664 (N_11664,N_5539,N_7127);
and U11665 (N_11665,N_5930,N_6328);
nand U11666 (N_11666,N_6910,N_8424);
or U11667 (N_11667,N_5309,N_9467);
or U11668 (N_11668,N_7232,N_5365);
and U11669 (N_11669,N_6021,N_8146);
nor U11670 (N_11670,N_8224,N_9486);
nor U11671 (N_11671,N_6218,N_8177);
nand U11672 (N_11672,N_7228,N_5424);
nand U11673 (N_11673,N_6961,N_9757);
and U11674 (N_11674,N_7993,N_9668);
xnor U11675 (N_11675,N_7262,N_9904);
and U11676 (N_11676,N_9394,N_9487);
nand U11677 (N_11677,N_8104,N_6669);
nand U11678 (N_11678,N_7042,N_5511);
nor U11679 (N_11679,N_7341,N_8490);
xnor U11680 (N_11680,N_5734,N_5241);
nor U11681 (N_11681,N_7747,N_8535);
nor U11682 (N_11682,N_6367,N_7948);
and U11683 (N_11683,N_6316,N_5410);
nor U11684 (N_11684,N_8569,N_6113);
and U11685 (N_11685,N_9414,N_9455);
nor U11686 (N_11686,N_8060,N_6042);
xor U11687 (N_11687,N_9781,N_5662);
or U11688 (N_11688,N_6331,N_6825);
xnor U11689 (N_11689,N_8056,N_8553);
or U11690 (N_11690,N_6809,N_6697);
nand U11691 (N_11691,N_8769,N_6117);
nor U11692 (N_11692,N_7276,N_9100);
and U11693 (N_11693,N_8770,N_7477);
nor U11694 (N_11694,N_8080,N_9807);
nor U11695 (N_11695,N_5478,N_9504);
xnor U11696 (N_11696,N_5387,N_8716);
or U11697 (N_11697,N_8409,N_6838);
or U11698 (N_11698,N_7176,N_5595);
or U11699 (N_11699,N_8190,N_7833);
nand U11700 (N_11700,N_8567,N_5996);
nor U11701 (N_11701,N_6635,N_6836);
nand U11702 (N_11702,N_5065,N_8078);
xnor U11703 (N_11703,N_8912,N_7761);
xnor U11704 (N_11704,N_5419,N_8776);
nand U11705 (N_11705,N_7208,N_5399);
xor U11706 (N_11706,N_8435,N_6732);
xnor U11707 (N_11707,N_8864,N_5376);
nand U11708 (N_11708,N_9583,N_8454);
xnor U11709 (N_11709,N_5019,N_5646);
nand U11710 (N_11710,N_8327,N_7976);
or U11711 (N_11711,N_9564,N_6950);
and U11712 (N_11712,N_9662,N_8726);
and U11713 (N_11713,N_9591,N_9383);
xnor U11714 (N_11714,N_6668,N_5817);
and U11715 (N_11715,N_7018,N_9939);
xnor U11716 (N_11716,N_8946,N_5046);
xnor U11717 (N_11717,N_6789,N_8550);
nor U11718 (N_11718,N_9041,N_7852);
or U11719 (N_11719,N_5833,N_6129);
or U11720 (N_11720,N_5272,N_7279);
or U11721 (N_11721,N_5367,N_8514);
nand U11722 (N_11722,N_9546,N_7568);
and U11723 (N_11723,N_5025,N_5576);
or U11724 (N_11724,N_8280,N_6154);
or U11725 (N_11725,N_7500,N_9516);
nor U11726 (N_11726,N_9923,N_7358);
nand U11727 (N_11727,N_8851,N_8860);
nand U11728 (N_11728,N_5324,N_6403);
or U11729 (N_11729,N_7223,N_8997);
xnor U11730 (N_11730,N_8945,N_9573);
or U11731 (N_11731,N_6164,N_5173);
and U11732 (N_11732,N_8625,N_5160);
and U11733 (N_11733,N_6977,N_7655);
xnor U11734 (N_11734,N_6815,N_5990);
or U11735 (N_11735,N_9273,N_8917);
or U11736 (N_11736,N_7758,N_7420);
or U11737 (N_11737,N_9422,N_9812);
or U11738 (N_11738,N_7822,N_7638);
xor U11739 (N_11739,N_8331,N_8326);
xnor U11740 (N_11740,N_6773,N_5418);
nor U11741 (N_11741,N_6238,N_9575);
nand U11742 (N_11742,N_6032,N_7681);
or U11743 (N_11743,N_5235,N_7019);
and U11744 (N_11744,N_5435,N_7094);
and U11745 (N_11745,N_8261,N_9194);
or U11746 (N_11746,N_8848,N_7985);
or U11747 (N_11747,N_5497,N_7706);
or U11748 (N_11748,N_6765,N_7566);
or U11749 (N_11749,N_5526,N_5698);
nor U11750 (N_11750,N_8229,N_9778);
xor U11751 (N_11751,N_6197,N_6082);
nand U11752 (N_11752,N_6097,N_7373);
xor U11753 (N_11753,N_9292,N_7222);
and U11754 (N_11754,N_8533,N_7731);
or U11755 (N_11755,N_6875,N_8659);
or U11756 (N_11756,N_7573,N_7556);
nand U11757 (N_11757,N_8054,N_7853);
xor U11758 (N_11758,N_5225,N_7841);
nand U11759 (N_11759,N_8355,N_9656);
nor U11760 (N_11760,N_6384,N_7760);
xnor U11761 (N_11761,N_9701,N_6440);
xnor U11762 (N_11762,N_9106,N_5675);
xnor U11763 (N_11763,N_6790,N_6934);
nor U11764 (N_11764,N_6387,N_5260);
nand U11765 (N_11765,N_6846,N_9412);
and U11766 (N_11766,N_8066,N_6535);
or U11767 (N_11767,N_9012,N_8944);
or U11768 (N_11768,N_6737,N_7871);
nand U11769 (N_11769,N_5380,N_7886);
or U11770 (N_11770,N_5202,N_8411);
and U11771 (N_11771,N_5935,N_8503);
xor U11772 (N_11772,N_6455,N_7219);
nand U11773 (N_11773,N_6065,N_6139);
or U11774 (N_11774,N_9823,N_7645);
nand U11775 (N_11775,N_7129,N_7766);
nand U11776 (N_11776,N_5631,N_5242);
xor U11777 (N_11777,N_6162,N_5431);
nand U11778 (N_11778,N_5982,N_5187);
xor U11779 (N_11779,N_5005,N_6024);
xor U11780 (N_11780,N_5395,N_6169);
nor U11781 (N_11781,N_9761,N_5564);
and U11782 (N_11782,N_9411,N_5966);
and U11783 (N_11783,N_8505,N_5374);
nor U11784 (N_11784,N_6704,N_7820);
or U11785 (N_11785,N_7330,N_7827);
and U11786 (N_11786,N_7599,N_7604);
nand U11787 (N_11787,N_9410,N_6625);
and U11788 (N_11788,N_9473,N_8491);
xnor U11789 (N_11789,N_8437,N_5963);
xor U11790 (N_11790,N_5658,N_6504);
xor U11791 (N_11791,N_8463,N_6399);
nand U11792 (N_11792,N_5036,N_5902);
nor U11793 (N_11793,N_8978,N_8452);
nor U11794 (N_11794,N_6975,N_7294);
nor U11795 (N_11795,N_8690,N_6515);
and U11796 (N_11796,N_7360,N_9308);
nor U11797 (N_11797,N_7799,N_9404);
nand U11798 (N_11798,N_6072,N_7642);
and U11799 (N_11799,N_9738,N_7395);
or U11800 (N_11800,N_7920,N_5623);
xnor U11801 (N_11801,N_9495,N_5428);
nor U11802 (N_11802,N_5008,N_9427);
nor U11803 (N_11803,N_5621,N_8318);
nand U11804 (N_11804,N_6314,N_5289);
and U11805 (N_11805,N_9763,N_9274);
nor U11806 (N_11806,N_6968,N_9506);
and U11807 (N_11807,N_6066,N_9861);
xor U11808 (N_11808,N_5797,N_5641);
nand U11809 (N_11809,N_7989,N_7802);
nor U11810 (N_11810,N_7024,N_8954);
or U11811 (N_11811,N_8644,N_6798);
xor U11812 (N_11812,N_7367,N_5190);
nand U11813 (N_11813,N_5565,N_5390);
nor U11814 (N_11814,N_7432,N_6274);
or U11815 (N_11815,N_5251,N_9057);
nand U11816 (N_11816,N_7586,N_7651);
nor U11817 (N_11817,N_5972,N_6767);
xor U11818 (N_11818,N_7015,N_5843);
nand U11819 (N_11819,N_7177,N_8906);
nor U11820 (N_11820,N_5227,N_7723);
nor U11821 (N_11821,N_7485,N_9123);
and U11822 (N_11822,N_7313,N_8451);
and U11823 (N_11823,N_9614,N_6824);
nand U11824 (N_11824,N_7577,N_5643);
nand U11825 (N_11825,N_8288,N_7397);
nor U11826 (N_11826,N_9627,N_5146);
nand U11827 (N_11827,N_8375,N_5617);
nor U11828 (N_11828,N_6298,N_7790);
nand U11829 (N_11829,N_9600,N_6223);
nand U11830 (N_11830,N_5574,N_6792);
nor U11831 (N_11831,N_6285,N_8666);
nor U11832 (N_11832,N_5311,N_6048);
nand U11833 (N_11833,N_8332,N_7221);
and U11834 (N_11834,N_6344,N_7215);
or U11835 (N_11835,N_7691,N_7241);
or U11836 (N_11836,N_5149,N_6487);
nand U11837 (N_11837,N_7083,N_5665);
and U11838 (N_11838,N_9797,N_9677);
and U11839 (N_11839,N_7220,N_6345);
xnor U11840 (N_11840,N_9254,N_8021);
nand U11841 (N_11841,N_5217,N_7888);
and U11842 (N_11842,N_6018,N_8760);
or U11843 (N_11843,N_5413,N_8680);
xor U11844 (N_11844,N_5607,N_9986);
and U11845 (N_11845,N_9330,N_6942);
nor U11846 (N_11846,N_9003,N_7942);
nand U11847 (N_11847,N_6513,N_5041);
nor U11848 (N_11848,N_8870,N_5185);
nand U11849 (N_11849,N_8301,N_7696);
nand U11850 (N_11850,N_9391,N_8270);
or U11851 (N_11851,N_9309,N_9691);
nand U11852 (N_11852,N_9569,N_5439);
and U11853 (N_11853,N_8450,N_8107);
nand U11854 (N_11854,N_8253,N_8816);
nor U11855 (N_11855,N_6394,N_6648);
or U11856 (N_11856,N_8563,N_8571);
nor U11857 (N_11857,N_5550,N_6379);
or U11858 (N_11858,N_6122,N_7591);
and U11859 (N_11859,N_6342,N_6029);
xor U11860 (N_11860,N_7705,N_7234);
nand U11861 (N_11861,N_7399,N_8128);
xor U11862 (N_11862,N_7713,N_7079);
xor U11863 (N_11863,N_5820,N_8281);
xor U11864 (N_11864,N_7800,N_9994);
nand U11865 (N_11865,N_5455,N_6817);
nand U11866 (N_11866,N_6682,N_5381);
xnor U11867 (N_11867,N_7968,N_7342);
xor U11868 (N_11868,N_5333,N_9200);
and U11869 (N_11869,N_9536,N_6310);
or U11870 (N_11870,N_8455,N_8333);
nor U11871 (N_11871,N_7692,N_5220);
and U11872 (N_11872,N_9813,N_8761);
and U11873 (N_11873,N_7354,N_5087);
or U11874 (N_11874,N_8733,N_9615);
or U11875 (N_11875,N_5814,N_7205);
xor U11876 (N_11876,N_5530,N_5261);
and U11877 (N_11877,N_9827,N_5696);
xor U11878 (N_11878,N_9319,N_7230);
or U11879 (N_11879,N_8840,N_5713);
and U11880 (N_11880,N_5059,N_5851);
nor U11881 (N_11881,N_8192,N_5591);
and U11882 (N_11882,N_9865,N_8135);
xor U11883 (N_11883,N_8173,N_8719);
xor U11884 (N_11884,N_9868,N_6233);
and U11885 (N_11885,N_7315,N_9298);
or U11886 (N_11886,N_5970,N_7366);
nor U11887 (N_11887,N_9652,N_9981);
nor U11888 (N_11888,N_7641,N_7967);
nor U11889 (N_11889,N_9729,N_7151);
nand U11890 (N_11890,N_6125,N_6141);
xnor U11891 (N_11891,N_6489,N_9025);
or U11892 (N_11892,N_6601,N_6251);
or U11893 (N_11893,N_6865,N_8169);
xor U11894 (N_11894,N_8837,N_5430);
xor U11895 (N_11895,N_6596,N_6742);
or U11896 (N_11896,N_8678,N_7191);
nor U11897 (N_11897,N_6594,N_5866);
and U11898 (N_11898,N_8294,N_7861);
xor U11899 (N_11899,N_6944,N_5872);
xnor U11900 (N_11900,N_8522,N_9828);
and U11901 (N_11901,N_5842,N_9443);
xnor U11902 (N_11902,N_5716,N_7881);
nand U11903 (N_11903,N_9917,N_5109);
or U11904 (N_11904,N_9375,N_6546);
nor U11905 (N_11905,N_6664,N_5890);
and U11906 (N_11906,N_6030,N_5869);
xor U11907 (N_11907,N_5135,N_8420);
nor U11908 (N_11908,N_5628,N_8369);
xnor U11909 (N_11909,N_9697,N_5598);
nor U11910 (N_11910,N_6971,N_6516);
nand U11911 (N_11911,N_8663,N_7915);
nor U11912 (N_11912,N_6192,N_5243);
nand U11913 (N_11913,N_8149,N_9906);
nand U11914 (N_11914,N_9932,N_9332);
or U11915 (N_11915,N_5721,N_7490);
or U11916 (N_11916,N_8446,N_5754);
xnor U11917 (N_11917,N_9588,N_7211);
nor U11918 (N_11918,N_9960,N_5906);
and U11919 (N_11919,N_9587,N_7943);
xor U11920 (N_11920,N_5443,N_5394);
and U11921 (N_11921,N_5103,N_7558);
xnor U11922 (N_11922,N_7676,N_6094);
and U11923 (N_11923,N_6871,N_5704);
and U11924 (N_11924,N_5979,N_5222);
nor U11925 (N_11925,N_6178,N_6167);
nand U11926 (N_11926,N_8278,N_8034);
nand U11927 (N_11927,N_5836,N_9260);
nand U11928 (N_11928,N_8878,N_7513);
xor U11929 (N_11929,N_5934,N_7931);
nand U11930 (N_11930,N_6536,N_5060);
and U11931 (N_11931,N_8969,N_8051);
or U11932 (N_11932,N_9226,N_6235);
or U11933 (N_11933,N_8755,N_6743);
xnor U11934 (N_11934,N_9618,N_6422);
or U11935 (N_11935,N_6228,N_8873);
nor U11936 (N_11936,N_7001,N_8583);
or U11937 (N_11937,N_6980,N_9632);
nor U11938 (N_11938,N_8970,N_9306);
xnor U11939 (N_11939,N_8142,N_6509);
nand U11940 (N_11940,N_5725,N_9403);
nand U11941 (N_11941,N_9686,N_8852);
xnor U11942 (N_11942,N_7217,N_7031);
or U11943 (N_11943,N_6586,N_7912);
xor U11944 (N_11944,N_9034,N_5137);
xnor U11945 (N_11945,N_7896,N_9381);
xor U11946 (N_11946,N_8274,N_9907);
nand U11947 (N_11947,N_7422,N_6270);
nand U11948 (N_11948,N_9500,N_8720);
xnor U11949 (N_11949,N_5229,N_5720);
nand U11950 (N_11950,N_7297,N_7767);
nand U11951 (N_11951,N_8868,N_5250);
nor U11952 (N_11952,N_9437,N_6908);
nor U11953 (N_11953,N_8015,N_6044);
or U11954 (N_11954,N_7695,N_5781);
nand U11955 (N_11955,N_9079,N_9376);
xor U11956 (N_11956,N_8829,N_8136);
xor U11957 (N_11957,N_6490,N_6820);
or U11958 (N_11958,N_9234,N_8979);
xor U11959 (N_11959,N_6175,N_8964);
xor U11960 (N_11960,N_8396,N_6814);
nand U11961 (N_11961,N_6801,N_6979);
and U11962 (N_11962,N_8292,N_5706);
and U11963 (N_11963,N_6784,N_9493);
or U11964 (N_11964,N_9229,N_7349);
nand U11965 (N_11965,N_8839,N_6894);
nand U11966 (N_11966,N_5473,N_5644);
or U11967 (N_11967,N_7218,N_5980);
or U11968 (N_11968,N_7690,N_7804);
nor U11969 (N_11969,N_7401,N_8215);
nand U11970 (N_11970,N_5489,N_5232);
or U11971 (N_11971,N_9038,N_5348);
and U11972 (N_11972,N_8831,N_9469);
nor U11973 (N_11973,N_6551,N_6375);
or U11974 (N_11974,N_8211,N_8057);
and U11975 (N_11975,N_9744,N_9103);
and U11976 (N_11976,N_9439,N_6172);
xor U11977 (N_11977,N_5375,N_7661);
nor U11978 (N_11978,N_6810,N_5513);
or U11979 (N_11979,N_9555,N_7480);
nand U11980 (N_11980,N_7921,N_8470);
nand U11981 (N_11981,N_9752,N_9050);
xnor U11982 (N_11982,N_9798,N_7172);
nand U11983 (N_11983,N_8199,N_6076);
nor U11984 (N_11984,N_5498,N_5504);
or U11985 (N_11985,N_6983,N_5179);
and U11986 (N_11986,N_9058,N_5559);
nor U11987 (N_11987,N_7613,N_5312);
and U11988 (N_11988,N_7844,N_8033);
nor U11989 (N_11989,N_6922,N_9399);
xor U11990 (N_11990,N_8512,N_9854);
nand U11991 (N_11991,N_7647,N_7534);
and U11992 (N_11992,N_9027,N_6562);
or U11993 (N_11993,N_8685,N_8606);
xnor U11994 (N_11994,N_7430,N_6482);
or U11995 (N_11995,N_8736,N_9736);
and U11996 (N_11996,N_7352,N_5207);
nor U11997 (N_11997,N_6220,N_5568);
or U11998 (N_11998,N_6951,N_9326);
or U11999 (N_11999,N_5823,N_7258);
nor U12000 (N_12000,N_7929,N_6195);
or U12001 (N_12001,N_6396,N_6541);
nand U12002 (N_12002,N_5026,N_7280);
nor U12003 (N_12003,N_8458,N_9479);
or U12004 (N_12004,N_8272,N_6750);
and U12005 (N_12005,N_7851,N_7400);
or U12006 (N_12006,N_7188,N_8950);
xor U12007 (N_12007,N_9745,N_5397);
nor U12008 (N_12008,N_9664,N_5687);
nor U12009 (N_12009,N_6187,N_7336);
and U12010 (N_12010,N_6617,N_6727);
nand U12011 (N_12011,N_7729,N_5544);
or U12012 (N_12012,N_9187,N_8597);
xnor U12013 (N_12013,N_9097,N_9525);
xnor U12014 (N_12014,N_7361,N_8992);
nand U12015 (N_12015,N_8953,N_5529);
and U12016 (N_12016,N_9985,N_6050);
nor U12017 (N_12017,N_8227,N_5882);
nand U12018 (N_12018,N_6111,N_7167);
or U12019 (N_12019,N_7554,N_5341);
and U12020 (N_12020,N_8019,N_8088);
or U12021 (N_12021,N_8534,N_5686);
xor U12022 (N_12022,N_5860,N_8980);
xor U12023 (N_12023,N_6060,N_9121);
nand U12024 (N_12024,N_5089,N_7828);
or U12025 (N_12025,N_8304,N_7971);
nor U12026 (N_12026,N_5784,N_5170);
xor U12027 (N_12027,N_5985,N_5477);
nor U12028 (N_12028,N_5907,N_7345);
xnor U12029 (N_12029,N_8797,N_5702);
nand U12030 (N_12030,N_7196,N_8965);
nor U12031 (N_12031,N_6426,N_5106);
or U12032 (N_12032,N_9887,N_7596);
and U12033 (N_12033,N_9327,N_8485);
or U12034 (N_12034,N_6701,N_8707);
nand U12035 (N_12035,N_6272,N_8208);
or U12036 (N_12036,N_6561,N_6634);
nand U12037 (N_12037,N_7733,N_6678);
and U12038 (N_12038,N_6043,N_5194);
nand U12039 (N_12039,N_7522,N_7579);
nand U12040 (N_12040,N_8996,N_6454);
nor U12041 (N_12041,N_8695,N_6053);
or U12042 (N_12042,N_7460,N_7043);
or U12043 (N_12043,N_9113,N_5819);
xor U12044 (N_12044,N_5196,N_7023);
or U12045 (N_12045,N_9594,N_5360);
xor U12046 (N_12046,N_5281,N_8706);
or U12047 (N_12047,N_8552,N_9592);
xnor U12048 (N_12048,N_9966,N_5035);
nand U12049 (N_12049,N_5299,N_9290);
or U12050 (N_12050,N_9105,N_6140);
or U12051 (N_12051,N_7864,N_7321);
or U12052 (N_12052,N_9081,N_8283);
xor U12053 (N_12053,N_5502,N_7482);
xnor U12054 (N_12054,N_9441,N_6476);
and U12055 (N_12055,N_8745,N_6827);
and U12056 (N_12056,N_8425,N_6878);
xor U12057 (N_12057,N_9520,N_7329);
nand U12058 (N_12058,N_8585,N_9829);
and U12059 (N_12059,N_5032,N_9834);
xnor U12060 (N_12060,N_6058,N_5868);
nor U12061 (N_12061,N_9498,N_6025);
or U12062 (N_12062,N_6188,N_9837);
and U12063 (N_12063,N_8555,N_9268);
nor U12064 (N_12064,N_5402,N_8502);
xnor U12065 (N_12065,N_9864,N_6521);
nand U12066 (N_12066,N_6768,N_6243);
or U12067 (N_12067,N_8392,N_5809);
nand U12068 (N_12068,N_9164,N_8410);
or U12069 (N_12069,N_6261,N_5673);
nand U12070 (N_12070,N_8185,N_6361);
nor U12071 (N_12071,N_6199,N_8315);
and U12072 (N_12072,N_6292,N_9320);
nand U12073 (N_12073,N_5749,N_6295);
and U12074 (N_12074,N_8947,N_8981);
nor U12075 (N_12075,N_7913,N_8664);
nand U12076 (N_12076,N_7542,N_5070);
or U12077 (N_12077,N_6694,N_8676);
nor U12078 (N_12078,N_7194,N_6962);
xnor U12079 (N_12079,N_5603,N_8421);
and U12080 (N_12080,N_8682,N_9586);
nand U12081 (N_12081,N_7290,N_9197);
nor U12082 (N_12082,N_6593,N_6189);
xnor U12083 (N_12083,N_9302,N_7080);
or U12084 (N_12084,N_9589,N_5292);
or U12085 (N_12085,N_8023,N_9004);
xnor U12086 (N_12086,N_8250,N_9384);
or U12087 (N_12087,N_9249,N_9483);
or U12088 (N_12088,N_5061,N_8527);
nor U12089 (N_12089,N_8218,N_8134);
xor U12090 (N_12090,N_7907,N_8616);
xor U12091 (N_12091,N_6628,N_5955);
xor U12092 (N_12092,N_6683,N_9449);
or U12093 (N_12093,N_6799,N_9509);
nand U12094 (N_12094,N_7549,N_6200);
xnor U12095 (N_12095,N_8483,N_6062);
xnor U12096 (N_12096,N_8939,N_9699);
nor U12097 (N_12097,N_6749,N_6534);
nor U12098 (N_12098,N_8155,N_9064);
nand U12099 (N_12099,N_6563,N_6606);
nand U12100 (N_12100,N_6600,N_6033);
or U12101 (N_12101,N_8046,N_6472);
or U12102 (N_12102,N_5752,N_8081);
nand U12103 (N_12103,N_5977,N_7478);
nor U12104 (N_12104,N_5480,N_7714);
xnor U12105 (N_12105,N_9505,N_5651);
xor U12106 (N_12106,N_5029,N_5238);
xnor U12107 (N_12107,N_6585,N_7540);
and U12108 (N_12108,N_6500,N_7868);
or U12109 (N_12109,N_5184,N_7936);
or U12110 (N_12110,N_5663,N_9508);
nor U12111 (N_12111,N_7990,N_9787);
nand U12112 (N_12112,N_5878,N_6415);
nand U12113 (N_12113,N_7225,N_8180);
nand U12114 (N_12114,N_8584,N_8382);
and U12115 (N_12115,N_9630,N_9680);
or U12116 (N_12116,N_8983,N_6016);
or U12117 (N_12117,N_5301,N_5543);
and U12118 (N_12118,N_8170,N_8610);
and U12119 (N_12119,N_6949,N_6703);
or U12120 (N_12120,N_6881,N_6369);
nor U12121 (N_12121,N_5620,N_8925);
nand U12122 (N_12122,N_9009,N_7970);
nor U12123 (N_12123,N_5476,N_8861);
nand U12124 (N_12124,N_8703,N_5320);
nor U12125 (N_12125,N_6808,N_5206);
xnor U12126 (N_12126,N_6519,N_8959);
and U12127 (N_12127,N_6967,N_5453);
nor U12128 (N_12128,N_8544,N_8069);
nand U12129 (N_12129,N_9235,N_8075);
nand U12130 (N_12130,N_8268,N_8498);
nand U12131 (N_12131,N_6754,N_9136);
nand U12132 (N_12132,N_9845,N_8367);
and U12133 (N_12133,N_6906,N_5841);
and U12134 (N_12134,N_6656,N_9818);
and U12135 (N_12135,N_7269,N_6411);
xor U12136 (N_12136,N_6138,N_9585);
or U12137 (N_12137,N_5049,N_8221);
and U12138 (N_12138,N_5625,N_8931);
xnor U12139 (N_12139,N_6127,N_9607);
nor U12140 (N_12140,N_5973,N_6306);
nand U12141 (N_12141,N_7914,N_5503);
xor U12142 (N_12142,N_8305,N_5705);
xnor U12143 (N_12143,N_6702,N_5147);
nor U12144 (N_12144,N_9261,N_5388);
or U12145 (N_12145,N_7377,N_6899);
and U12146 (N_12146,N_8162,N_7387);
and U12147 (N_12147,N_7608,N_7725);
nor U12148 (N_12148,N_9130,N_9950);
or U12149 (N_12149,N_6401,N_9311);
or U12150 (N_12150,N_7091,N_9707);
nor U12151 (N_12151,N_8013,N_5624);
or U12152 (N_12152,N_6988,N_5743);
or U12153 (N_12153,N_5398,N_7893);
xnor U12154 (N_12154,N_5000,N_7745);
xnor U12155 (N_12155,N_8895,N_8977);
or U12156 (N_12156,N_7051,N_5451);
or U12157 (N_12157,N_5337,N_7735);
nand U12158 (N_12158,N_6819,N_6672);
nand U12159 (N_12159,N_6888,N_6558);
nor U12160 (N_12160,N_5472,N_5126);
nor U12161 (N_12161,N_5601,N_7634);
nand U12162 (N_12162,N_9250,N_6335);
nand U12163 (N_12163,N_5258,N_7630);
nor U12164 (N_12164,N_9959,N_7277);
xor U12165 (N_12165,N_7190,N_9559);
nand U12166 (N_12166,N_5815,N_6230);
or U12167 (N_12167,N_6834,N_5361);
and U12168 (N_12168,N_7347,N_6540);
nor U12169 (N_12169,N_8398,N_8620);
and U12170 (N_12170,N_9458,N_6688);
or U12171 (N_12171,N_5701,N_7412);
and U12172 (N_12172,N_6196,N_8026);
and U12173 (N_12173,N_8882,N_5983);
nor U12174 (N_12174,N_5575,N_9993);
nand U12175 (N_12175,N_8239,N_6280);
and U12176 (N_12176,N_9224,N_9361);
nand U12177 (N_12177,N_9429,N_8593);
nand U12178 (N_12178,N_7891,N_8357);
and U12179 (N_12179,N_6877,N_6432);
and U12180 (N_12180,N_6466,N_5920);
nor U12181 (N_12181,N_7835,N_7918);
and U12182 (N_12182,N_9220,N_9952);
xnor U12183 (N_12183,N_8806,N_9639);
nor U12184 (N_12184,N_5037,N_5677);
nor U12185 (N_12185,N_8343,N_7684);
xor U12186 (N_12186,N_8220,N_6735);
nor U12187 (N_12187,N_6764,N_6460);
or U12188 (N_12188,N_6505,N_7004);
xor U12189 (N_12189,N_6622,N_5325);
nand U12190 (N_12190,N_6642,N_6406);
and U12191 (N_12191,N_5924,N_8949);
or U12192 (N_12192,N_7472,N_9674);
and U12193 (N_12193,N_8942,N_7020);
or U12194 (N_12194,N_7906,N_8952);
or U12195 (N_12195,N_8871,N_6041);
xnor U12196 (N_12196,N_8236,N_6040);
nand U12197 (N_12197,N_7863,N_8302);
and U12198 (N_12198,N_5661,N_6740);
xnor U12199 (N_12199,N_7388,N_6343);
nand U12200 (N_12200,N_7146,N_9074);
or U12201 (N_12201,N_7298,N_5426);
nand U12202 (N_12202,N_7753,N_7950);
or U12203 (N_12203,N_6263,N_5054);
nor U12204 (N_12204,N_9313,N_5571);
nor U12205 (N_12205,N_5266,N_5737);
xnor U12206 (N_12206,N_5062,N_8183);
xor U12207 (N_12207,N_6088,N_8477);
xnor U12208 (N_12208,N_5688,N_5956);
nor U12209 (N_12209,N_5022,N_6085);
nand U12210 (N_12210,N_9606,N_7455);
nor U12211 (N_12211,N_9989,N_9628);
nor U12212 (N_12212,N_5770,N_8551);
nor U12213 (N_12213,N_6582,N_8548);
nor U12214 (N_12214,N_9008,N_9552);
xor U12215 (N_12215,N_8478,N_6049);
and U12216 (N_12216,N_5765,N_5340);
nand U12217 (N_12217,N_7959,N_5066);
xor U12218 (N_12218,N_5958,N_9205);
nand U12219 (N_12219,N_7905,N_9092);
nor U12220 (N_12220,N_6408,N_6325);
nand U12221 (N_12221,N_9158,N_7711);
nand U12222 (N_12222,N_5879,N_7433);
xnor U12223 (N_12223,N_6714,N_8251);
nor U12224 (N_12224,N_8744,N_5329);
or U12225 (N_12225,N_6660,N_8447);
nor U12226 (N_12226,N_5107,N_6574);
nand U12227 (N_12227,N_7626,N_8319);
and U12228 (N_12228,N_7008,N_9148);
nor U12229 (N_12229,N_6729,N_6356);
nor U12230 (N_12230,N_8346,N_5987);
nor U12231 (N_12231,N_7204,N_7170);
nor U12232 (N_12232,N_8385,N_8757);
and U12233 (N_12233,N_7012,N_5331);
xor U12234 (N_12234,N_6989,N_8630);
xor U12235 (N_12235,N_7292,N_5855);
xnor U12236 (N_12236,N_6963,N_8642);
xnor U12237 (N_12237,N_7663,N_9533);
nand U12238 (N_12238,N_7962,N_9790);
xor U12239 (N_12239,N_9314,N_6047);
and U12240 (N_12240,N_5255,N_9451);
and U12241 (N_12241,N_9794,N_7308);
nand U12242 (N_12242,N_7772,N_6143);
xor U12243 (N_12243,N_6679,N_5316);
and U12244 (N_12244,N_8059,N_7847);
nand U12245 (N_12245,N_9016,N_6303);
nor U12246 (N_12246,N_5659,N_7376);
xor U12247 (N_12247,N_6433,N_9808);
nand U12248 (N_12248,N_5590,N_8511);
nand U12249 (N_12249,N_8465,N_8923);
and U12250 (N_12250,N_9392,N_7597);
or U12251 (N_12251,N_8775,N_6282);
and U12252 (N_12252,N_8290,N_8576);
or U12253 (N_12253,N_7512,N_7110);
xnor U12254 (N_12254,N_8648,N_9247);
nor U12255 (N_12255,N_9844,N_5115);
or U12256 (N_12256,N_6431,N_9611);
or U12257 (N_12257,N_8432,N_5520);
nand U12258 (N_12258,N_9849,N_8209);
or U12259 (N_12259,N_6752,N_6653);
nand U12260 (N_12260,N_7639,N_6787);
and U12261 (N_12261,N_6867,N_5538);
or U12262 (N_12262,N_6078,N_6288);
and U12263 (N_12263,N_7415,N_6991);
or U12264 (N_12264,N_8495,N_5703);
nor U12265 (N_12265,N_6254,N_5017);
nor U12266 (N_12266,N_9073,N_7136);
xor U12267 (N_12267,N_5454,N_6947);
or U12268 (N_12268,N_6960,N_8822);
nand U12269 (N_12269,N_5051,N_9289);
and U12270 (N_12270,N_8742,N_5547);
or U12271 (N_12271,N_9415,N_5938);
or U12272 (N_12272,N_6017,N_5407);
or U12273 (N_12273,N_9201,N_5020);
or U12274 (N_12274,N_6627,N_9104);
or U12275 (N_12275,N_5484,N_6637);
nor U12276 (N_12276,N_8856,N_6004);
xor U12277 (N_12277,N_7823,N_6450);
and U12278 (N_12278,N_6436,N_9805);
or U12279 (N_12279,N_9998,N_9147);
nor U12280 (N_12280,N_6829,N_5290);
and U12281 (N_12281,N_9502,N_7777);
or U12282 (N_12282,N_8431,N_8130);
nor U12283 (N_12283,N_5045,N_8429);
nor U12284 (N_12284,N_5129,N_7093);
and U12285 (N_12285,N_6994,N_7501);
xnor U12286 (N_12286,N_7025,N_5715);
and U12287 (N_12287,N_8009,N_8233);
and U12288 (N_12288,N_9282,N_6008);
nand U12289 (N_12289,N_8815,N_7511);
nor U12290 (N_12290,N_9570,N_5789);
and U12291 (N_12291,N_9001,N_9839);
nor U12292 (N_12292,N_8244,N_6253);
xnor U12293 (N_12293,N_5556,N_9721);
and U12294 (N_12294,N_6462,N_9349);
nor U12295 (N_12295,N_7889,N_9230);
xor U12296 (N_12296,N_6121,N_9927);
nand U12297 (N_12297,N_7791,N_5279);
nand U12298 (N_12298,N_9000,N_6287);
xnor U12299 (N_12299,N_6260,N_5259);
nand U12300 (N_12300,N_5731,N_9489);
nor U12301 (N_12301,N_6194,N_9911);
xor U12302 (N_12302,N_5177,N_9688);
or U12303 (N_12303,N_6986,N_8269);
and U12304 (N_12304,N_9277,N_6009);
or U12305 (N_12305,N_7775,N_5101);
nor U12306 (N_12306,N_9063,N_8803);
nor U12307 (N_12307,N_8403,N_8926);
nor U12308 (N_12308,N_7317,N_5364);
or U12309 (N_12309,N_9901,N_7506);
xor U12310 (N_12310,N_7461,N_5306);
nand U12311 (N_12311,N_5213,N_9175);
and U12312 (N_12312,N_5023,N_9020);
xnor U12313 (N_12313,N_5091,N_6389);
nand U12314 (N_12314,N_7137,N_8908);
nand U12315 (N_12315,N_6180,N_8670);
and U12316 (N_12316,N_9685,N_7056);
nor U12317 (N_12317,N_8580,N_8467);
nand U12318 (N_12318,N_8532,N_9275);
xor U12319 (N_12319,N_9706,N_7240);
or U12320 (N_12320,N_5755,N_5389);
nor U12321 (N_12321,N_6912,N_9328);
and U12322 (N_12322,N_7236,N_5148);
or U12323 (N_12323,N_8920,N_7882);
or U12324 (N_12324,N_7413,N_9054);
and U12325 (N_12325,N_8345,N_7058);
xnor U12326 (N_12326,N_6246,N_8867);
nor U12327 (N_12327,N_5010,N_7523);
and U12328 (N_12328,N_7169,N_6404);
nand U12329 (N_12329,N_6775,N_9841);
xnor U12330 (N_12330,N_9366,N_7924);
or U12331 (N_12331,N_7887,N_7910);
nor U12332 (N_12332,N_8509,N_6232);
nand U12333 (N_12333,N_8525,N_9772);
xor U12334 (N_12334,N_7666,N_8174);
nand U12335 (N_12335,N_9352,N_8934);
and U12336 (N_12336,N_5750,N_6286);
or U12337 (N_12337,N_9337,N_5464);
nor U12338 (N_12338,N_7175,N_7643);
xnor U12339 (N_12339,N_8722,N_9915);
nand U12340 (N_12340,N_6699,N_6821);
and U12341 (N_12341,N_7069,N_7209);
nand U12342 (N_12342,N_6297,N_9099);
and U12343 (N_12343,N_6059,N_9789);
nor U12344 (N_12344,N_5909,N_7728);
or U12345 (N_12345,N_8974,N_5345);
and U12346 (N_12346,N_5893,N_5012);
nor U12347 (N_12347,N_6915,N_8646);
xor U12348 (N_12348,N_6788,N_8370);
nor U12349 (N_12349,N_8055,N_7603);
and U12350 (N_12350,N_5212,N_5652);
xnor U12351 (N_12351,N_9452,N_7283);
or U12352 (N_12352,N_7543,N_6064);
nor U12353 (N_12353,N_9553,N_7806);
and U12354 (N_12354,N_7842,N_5653);
xnor U12355 (N_12355,N_9007,N_8613);
nor U12356 (N_12356,N_7132,N_8962);
and U12357 (N_12357,N_7233,N_5226);
nor U12358 (N_12358,N_9369,N_6686);
nand U12359 (N_12359,N_8862,N_5096);
or U12360 (N_12360,N_6557,N_9822);
nor U12361 (N_12361,N_8293,N_5302);
xor U12362 (N_12362,N_8144,N_9576);
nand U12363 (N_12363,N_5467,N_9681);
nor U12364 (N_12364,N_7693,N_5198);
or U12365 (N_12365,N_7683,N_9421);
xor U12366 (N_12366,N_6736,N_8854);
nand U12367 (N_12367,N_6080,N_9018);
nor U12368 (N_12368,N_9471,N_5874);
xnor U12369 (N_12369,N_7452,N_6486);
and U12370 (N_12370,N_6284,N_6929);
and U12371 (N_12371,N_8374,N_9359);
nor U12372 (N_12372,N_8159,N_7911);
and U12373 (N_12373,N_8472,N_9931);
or U12374 (N_12374,N_9382,N_6649);
xnor U12375 (N_12375,N_6946,N_7453);
nor U12376 (N_12376,N_6352,N_6948);
and U12377 (N_12377,N_8407,N_7417);
xnor U12378 (N_12378,N_6939,N_5730);
nor U12379 (N_12379,N_7917,N_5264);
nand U12380 (N_12380,N_6185,N_9279);
xor U12381 (N_12381,N_9307,N_5349);
and U12382 (N_12382,N_5165,N_9895);
nor U12383 (N_12383,N_5358,N_7517);
and U12384 (N_12384,N_8652,N_5605);
nand U12385 (N_12385,N_7068,N_9799);
nand U12386 (N_12386,N_6000,N_7181);
xnor U12387 (N_12387,N_9720,N_6576);
nor U12388 (N_12388,N_9963,N_6859);
nor U12389 (N_12389,N_9358,N_5382);
nand U12390 (N_12390,N_6026,N_8277);
and U12391 (N_12391,N_7832,N_9742);
and U12392 (N_12392,N_7716,N_6434);
nand U12393 (N_12393,N_6115,N_8322);
nand U12394 (N_12394,N_8520,N_6800);
or U12395 (N_12395,N_7809,N_7273);
or U12396 (N_12396,N_8819,N_6153);
nand U12397 (N_12397,N_9800,N_8384);
nand U12398 (N_12398,N_7930,N_7105);
nand U12399 (N_12399,N_5865,N_6869);
nand U12400 (N_12400,N_7078,N_8649);
nand U12401 (N_12401,N_5807,N_7394);
xor U12402 (N_12402,N_9976,N_8524);
or U12403 (N_12403,N_5875,N_9420);
and U12404 (N_12404,N_8461,N_9641);
nand U12405 (N_12405,N_5811,N_7509);
nor U12406 (N_12406,N_9990,N_7531);
or U12407 (N_12407,N_9005,N_9110);
or U12408 (N_12408,N_6793,N_7610);
nor U12409 (N_12409,N_7662,N_7631);
and U12410 (N_12410,N_5960,N_8531);
nand U12411 (N_12411,N_9623,N_7386);
or U12412 (N_12412,N_6311,N_9879);
xor U12413 (N_12413,N_5237,N_7496);
nor U12414 (N_12414,N_8266,N_5548);
nand U12415 (N_12415,N_9919,N_6904);
xor U12416 (N_12416,N_6982,N_7140);
nand U12417 (N_12417,N_6517,N_8043);
and U12418 (N_12418,N_8715,N_7207);
or U12419 (N_12419,N_9336,N_7521);
or U12420 (N_12420,N_5594,N_6496);
xor U12421 (N_12421,N_7312,N_7022);
nor U12422 (N_12422,N_7195,N_9257);
xnor U12423 (N_12423,N_8143,N_6905);
nand U12424 (N_12424,N_7202,N_7026);
or U12425 (N_12425,N_6785,N_9687);
nand U12426 (N_12426,N_6216,N_6116);
nor U12427 (N_12427,N_9363,N_8052);
and U12428 (N_12428,N_8160,N_6393);
nor U12429 (N_12429,N_8098,N_8053);
or U12430 (N_12430,N_5733,N_7498);
and U12431 (N_12431,N_7446,N_9035);
and U12432 (N_12432,N_8401,N_9795);
or U12433 (N_12433,N_8372,N_9642);
or U12434 (N_12434,N_7739,N_8605);
and U12435 (N_12435,N_9780,N_6055);
nor U12436 (N_12436,N_5016,N_6689);
and U12437 (N_12437,N_8106,N_6567);
nand U12438 (N_12438,N_9878,N_7183);
and U12439 (N_12439,N_5248,N_7866);
or U12440 (N_12440,N_9217,N_7157);
and U12441 (N_12441,N_5033,N_6549);
and U12442 (N_12442,N_5125,N_6830);
or U12443 (N_12443,N_9972,N_9519);
or U12444 (N_12444,N_8014,N_5240);
nand U12445 (N_12445,N_8152,N_8688);
nor U12446 (N_12446,N_6559,N_8632);
nor U12447 (N_12447,N_7253,N_6109);
or U12448 (N_12448,N_7636,N_9472);
nand U12449 (N_12449,N_6259,N_6512);
and U12450 (N_12450,N_6077,N_6374);
nor U12451 (N_12451,N_9096,N_9030);
nand U12452 (N_12452,N_8012,N_8237);
xor U12453 (N_12453,N_6186,N_9565);
xnor U12454 (N_12454,N_8743,N_8475);
or U12455 (N_12455,N_9216,N_9602);
nor U12456 (N_12456,N_5308,N_5831);
or U12457 (N_12457,N_5483,N_7309);
nand U12458 (N_12458,N_5689,N_9490);
and U12459 (N_12459,N_7116,N_7249);
and U12460 (N_12460,N_9722,N_8468);
nand U12461 (N_12461,N_8094,N_6105);
or U12462 (N_12462,N_8516,N_7467);
xor U12463 (N_12463,N_9374,N_8489);
nor U12464 (N_12464,N_8205,N_8723);
xnor U12465 (N_12465,N_7409,N_9223);
and U12466 (N_12466,N_6514,N_5203);
xor U12467 (N_12467,N_8093,N_7854);
and U12468 (N_12468,N_9975,N_5262);
or U12469 (N_12469,N_6471,N_5694);
xnor U12470 (N_12470,N_7122,N_6879);
nand U12471 (N_12471,N_5780,N_5383);
nand U12472 (N_12472,N_5172,N_9940);
or U12473 (N_12473,N_5178,N_5740);
xor U12474 (N_12474,N_8187,N_8935);
nand U12475 (N_12475,N_5273,N_6733);
nor U12476 (N_12476,N_7902,N_5640);
xor U12477 (N_12477,N_8709,N_7425);
nand U12478 (N_12478,N_9107,N_6893);
xor U12479 (N_12479,N_5518,N_8810);
nand U12480 (N_12480,N_6885,N_5903);
and U12481 (N_12481,N_6731,N_7261);
xnor U12482 (N_12482,N_8240,N_8933);
xnor U12483 (N_12483,N_6329,N_5003);
nand U12484 (N_12484,N_5437,N_8956);
nand U12485 (N_12485,N_7575,N_6099);
or U12486 (N_12486,N_5639,N_6926);
or U12487 (N_12487,N_8122,N_9857);
or U12488 (N_12488,N_8222,N_8764);
xnor U12489 (N_12489,N_6203,N_9042);
and U12490 (N_12490,N_7737,N_8025);
and U12491 (N_12491,N_9695,N_9206);
and U12492 (N_12492,N_8783,N_9188);
or U12493 (N_12493,N_6034,N_7301);
nor U12494 (N_12494,N_9240,N_6012);
nand U12495 (N_12495,N_6992,N_5928);
nand U12496 (N_12496,N_8825,N_6643);
nor U12497 (N_12497,N_7306,N_9912);
and U12498 (N_12498,N_7090,N_6794);
and U12499 (N_12499,N_9023,N_5214);
xor U12500 (N_12500,N_7961,N_7250);
or U12501 (N_12501,N_6821,N_7227);
or U12502 (N_12502,N_6535,N_6170);
or U12503 (N_12503,N_5782,N_5146);
or U12504 (N_12504,N_6504,N_5038);
nand U12505 (N_12505,N_7746,N_9054);
nor U12506 (N_12506,N_8623,N_9661);
nor U12507 (N_12507,N_6305,N_6767);
and U12508 (N_12508,N_8144,N_8684);
or U12509 (N_12509,N_8965,N_9077);
xnor U12510 (N_12510,N_8018,N_9817);
and U12511 (N_12511,N_9346,N_5639);
and U12512 (N_12512,N_5891,N_7646);
and U12513 (N_12513,N_7013,N_7477);
or U12514 (N_12514,N_8558,N_6733);
or U12515 (N_12515,N_8572,N_5398);
and U12516 (N_12516,N_7972,N_5227);
or U12517 (N_12517,N_7464,N_7802);
nor U12518 (N_12518,N_7999,N_8985);
nor U12519 (N_12519,N_9014,N_6103);
and U12520 (N_12520,N_5171,N_8590);
nand U12521 (N_12521,N_9307,N_9319);
nand U12522 (N_12522,N_8315,N_7157);
nand U12523 (N_12523,N_7577,N_8916);
nor U12524 (N_12524,N_8026,N_5216);
or U12525 (N_12525,N_6858,N_9348);
or U12526 (N_12526,N_7521,N_9289);
nor U12527 (N_12527,N_5778,N_6028);
nand U12528 (N_12528,N_7113,N_7746);
or U12529 (N_12529,N_8927,N_5843);
xor U12530 (N_12530,N_9569,N_5545);
xnor U12531 (N_12531,N_7419,N_6188);
nor U12532 (N_12532,N_9751,N_7852);
xnor U12533 (N_12533,N_6025,N_8056);
nor U12534 (N_12534,N_5967,N_6658);
nor U12535 (N_12535,N_6335,N_6462);
nand U12536 (N_12536,N_5476,N_5054);
or U12537 (N_12537,N_6465,N_6811);
xor U12538 (N_12538,N_5673,N_8544);
nor U12539 (N_12539,N_5314,N_7759);
or U12540 (N_12540,N_5275,N_9725);
xor U12541 (N_12541,N_8824,N_9767);
or U12542 (N_12542,N_9996,N_6625);
or U12543 (N_12543,N_8609,N_9350);
and U12544 (N_12544,N_6328,N_7047);
and U12545 (N_12545,N_8855,N_9135);
nor U12546 (N_12546,N_6736,N_9061);
nand U12547 (N_12547,N_9576,N_5197);
nand U12548 (N_12548,N_9020,N_7350);
xnor U12549 (N_12549,N_6228,N_8387);
and U12550 (N_12550,N_9726,N_6612);
and U12551 (N_12551,N_8199,N_8468);
nor U12552 (N_12552,N_9607,N_7802);
nand U12553 (N_12553,N_6404,N_5922);
nand U12554 (N_12554,N_9034,N_9142);
or U12555 (N_12555,N_9301,N_6948);
nand U12556 (N_12556,N_8601,N_5486);
or U12557 (N_12557,N_6053,N_5560);
nor U12558 (N_12558,N_5109,N_8829);
nor U12559 (N_12559,N_8118,N_7514);
and U12560 (N_12560,N_8572,N_8457);
xor U12561 (N_12561,N_6378,N_5736);
and U12562 (N_12562,N_9189,N_6890);
xor U12563 (N_12563,N_7392,N_7437);
and U12564 (N_12564,N_6799,N_9668);
nor U12565 (N_12565,N_5575,N_8348);
nor U12566 (N_12566,N_6252,N_5357);
nand U12567 (N_12567,N_8277,N_6181);
xnor U12568 (N_12568,N_6595,N_6494);
nor U12569 (N_12569,N_8585,N_8314);
nor U12570 (N_12570,N_8537,N_5737);
nor U12571 (N_12571,N_8419,N_8479);
and U12572 (N_12572,N_5678,N_7555);
nor U12573 (N_12573,N_7031,N_6048);
xnor U12574 (N_12574,N_9252,N_9514);
nand U12575 (N_12575,N_7441,N_7809);
xor U12576 (N_12576,N_5181,N_9665);
xnor U12577 (N_12577,N_6765,N_7932);
nor U12578 (N_12578,N_7748,N_5059);
or U12579 (N_12579,N_8445,N_5400);
nor U12580 (N_12580,N_7293,N_8916);
or U12581 (N_12581,N_8685,N_5394);
xnor U12582 (N_12582,N_9791,N_8076);
nor U12583 (N_12583,N_8324,N_6704);
and U12584 (N_12584,N_7111,N_7341);
or U12585 (N_12585,N_7809,N_9681);
and U12586 (N_12586,N_5782,N_5347);
xnor U12587 (N_12587,N_5699,N_8451);
or U12588 (N_12588,N_7345,N_5773);
xnor U12589 (N_12589,N_6463,N_6922);
xnor U12590 (N_12590,N_6736,N_9650);
and U12591 (N_12591,N_9064,N_7621);
or U12592 (N_12592,N_7188,N_5506);
or U12593 (N_12593,N_5285,N_9924);
or U12594 (N_12594,N_7430,N_6980);
or U12595 (N_12595,N_8125,N_7380);
xor U12596 (N_12596,N_9185,N_5112);
nor U12597 (N_12597,N_5256,N_8954);
nor U12598 (N_12598,N_7005,N_7044);
xor U12599 (N_12599,N_5971,N_6827);
nand U12600 (N_12600,N_8191,N_7259);
and U12601 (N_12601,N_8504,N_8813);
and U12602 (N_12602,N_7034,N_5196);
xor U12603 (N_12603,N_8752,N_5676);
and U12604 (N_12604,N_9907,N_7829);
or U12605 (N_12605,N_5948,N_5513);
nand U12606 (N_12606,N_5643,N_8681);
nor U12607 (N_12607,N_5424,N_9874);
and U12608 (N_12608,N_8051,N_8600);
or U12609 (N_12609,N_6007,N_7107);
nand U12610 (N_12610,N_8686,N_6334);
xnor U12611 (N_12611,N_8930,N_6833);
nor U12612 (N_12612,N_7016,N_5097);
nand U12613 (N_12613,N_5667,N_6977);
xnor U12614 (N_12614,N_5427,N_7868);
or U12615 (N_12615,N_7002,N_8889);
nand U12616 (N_12616,N_7000,N_6695);
nor U12617 (N_12617,N_8027,N_6613);
xor U12618 (N_12618,N_6215,N_5604);
nand U12619 (N_12619,N_8445,N_8389);
or U12620 (N_12620,N_8841,N_5770);
nor U12621 (N_12621,N_7509,N_7074);
nand U12622 (N_12622,N_9254,N_5397);
xnor U12623 (N_12623,N_6909,N_7897);
and U12624 (N_12624,N_5076,N_6164);
nand U12625 (N_12625,N_8782,N_5620);
or U12626 (N_12626,N_9910,N_7266);
or U12627 (N_12627,N_5033,N_6881);
or U12628 (N_12628,N_8725,N_6698);
nor U12629 (N_12629,N_5769,N_5037);
or U12630 (N_12630,N_5658,N_8807);
xnor U12631 (N_12631,N_7230,N_8843);
nor U12632 (N_12632,N_9297,N_6504);
nand U12633 (N_12633,N_6158,N_7550);
nor U12634 (N_12634,N_9505,N_8368);
nor U12635 (N_12635,N_6764,N_6795);
and U12636 (N_12636,N_8608,N_6419);
xnor U12637 (N_12637,N_8280,N_8641);
nand U12638 (N_12638,N_7691,N_8213);
nand U12639 (N_12639,N_6023,N_9209);
nand U12640 (N_12640,N_5147,N_6174);
or U12641 (N_12641,N_7464,N_5149);
nor U12642 (N_12642,N_6144,N_6641);
or U12643 (N_12643,N_6156,N_8952);
or U12644 (N_12644,N_8240,N_8910);
or U12645 (N_12645,N_7159,N_9634);
xor U12646 (N_12646,N_9536,N_8261);
nor U12647 (N_12647,N_9871,N_6462);
xor U12648 (N_12648,N_9170,N_7933);
and U12649 (N_12649,N_7113,N_8584);
nand U12650 (N_12650,N_6860,N_9695);
nand U12651 (N_12651,N_5083,N_6394);
nand U12652 (N_12652,N_7552,N_7625);
nor U12653 (N_12653,N_7255,N_7747);
nor U12654 (N_12654,N_6068,N_5083);
or U12655 (N_12655,N_5858,N_7628);
and U12656 (N_12656,N_8255,N_5350);
xnor U12657 (N_12657,N_7927,N_7914);
xor U12658 (N_12658,N_7177,N_8852);
nand U12659 (N_12659,N_8680,N_9298);
nand U12660 (N_12660,N_7758,N_5931);
nor U12661 (N_12661,N_5488,N_5933);
and U12662 (N_12662,N_7919,N_9472);
xnor U12663 (N_12663,N_5712,N_5954);
and U12664 (N_12664,N_8336,N_9832);
nor U12665 (N_12665,N_6100,N_5284);
or U12666 (N_12666,N_5477,N_6620);
nand U12667 (N_12667,N_8019,N_9939);
or U12668 (N_12668,N_9921,N_7086);
or U12669 (N_12669,N_7594,N_9844);
and U12670 (N_12670,N_8050,N_5304);
nor U12671 (N_12671,N_8610,N_8138);
nor U12672 (N_12672,N_5372,N_6669);
or U12673 (N_12673,N_8611,N_5173);
nand U12674 (N_12674,N_5157,N_5499);
or U12675 (N_12675,N_8382,N_6383);
and U12676 (N_12676,N_7384,N_8241);
or U12677 (N_12677,N_6681,N_9117);
and U12678 (N_12678,N_5649,N_5544);
or U12679 (N_12679,N_5620,N_9706);
xor U12680 (N_12680,N_6707,N_5219);
nor U12681 (N_12681,N_7881,N_5168);
nand U12682 (N_12682,N_9603,N_9080);
xnor U12683 (N_12683,N_6748,N_8835);
and U12684 (N_12684,N_5824,N_7975);
nand U12685 (N_12685,N_5315,N_9530);
nand U12686 (N_12686,N_9683,N_8671);
xnor U12687 (N_12687,N_6006,N_9466);
nand U12688 (N_12688,N_9908,N_7955);
nand U12689 (N_12689,N_5475,N_9446);
nand U12690 (N_12690,N_6077,N_5308);
nor U12691 (N_12691,N_6482,N_7815);
nor U12692 (N_12692,N_6876,N_7810);
or U12693 (N_12693,N_9629,N_7277);
nand U12694 (N_12694,N_8273,N_8905);
or U12695 (N_12695,N_9373,N_9824);
xor U12696 (N_12696,N_7096,N_8488);
or U12697 (N_12697,N_9366,N_7899);
nand U12698 (N_12698,N_8667,N_6449);
xnor U12699 (N_12699,N_5764,N_9209);
nand U12700 (N_12700,N_5807,N_6466);
nand U12701 (N_12701,N_7677,N_7760);
nor U12702 (N_12702,N_9976,N_8446);
nor U12703 (N_12703,N_7385,N_7523);
xnor U12704 (N_12704,N_5320,N_7112);
xor U12705 (N_12705,N_7299,N_5353);
nor U12706 (N_12706,N_7105,N_5870);
xnor U12707 (N_12707,N_9395,N_6929);
xor U12708 (N_12708,N_8252,N_9119);
nand U12709 (N_12709,N_6870,N_9681);
or U12710 (N_12710,N_7785,N_6261);
nor U12711 (N_12711,N_5813,N_7135);
or U12712 (N_12712,N_5853,N_7104);
nor U12713 (N_12713,N_6453,N_7606);
and U12714 (N_12714,N_9669,N_9590);
nand U12715 (N_12715,N_8689,N_6676);
or U12716 (N_12716,N_5018,N_8817);
xnor U12717 (N_12717,N_7522,N_6689);
nand U12718 (N_12718,N_8335,N_6993);
and U12719 (N_12719,N_7360,N_6030);
and U12720 (N_12720,N_9488,N_6727);
nor U12721 (N_12721,N_6116,N_9973);
or U12722 (N_12722,N_8703,N_9030);
or U12723 (N_12723,N_5530,N_5693);
xor U12724 (N_12724,N_6852,N_7659);
and U12725 (N_12725,N_5825,N_9572);
and U12726 (N_12726,N_5107,N_6337);
or U12727 (N_12727,N_9950,N_5789);
nand U12728 (N_12728,N_6639,N_7616);
and U12729 (N_12729,N_9898,N_5297);
xor U12730 (N_12730,N_7224,N_8607);
nor U12731 (N_12731,N_5726,N_8674);
and U12732 (N_12732,N_9852,N_7382);
nand U12733 (N_12733,N_7457,N_7640);
nand U12734 (N_12734,N_9664,N_6893);
and U12735 (N_12735,N_5664,N_6417);
nor U12736 (N_12736,N_6736,N_6334);
xnor U12737 (N_12737,N_5041,N_8173);
or U12738 (N_12738,N_5023,N_6654);
or U12739 (N_12739,N_8600,N_7766);
nand U12740 (N_12740,N_8721,N_9988);
nand U12741 (N_12741,N_8492,N_7338);
nand U12742 (N_12742,N_5015,N_6447);
or U12743 (N_12743,N_9118,N_6385);
nand U12744 (N_12744,N_9877,N_7352);
and U12745 (N_12745,N_6894,N_7799);
nor U12746 (N_12746,N_6768,N_7024);
and U12747 (N_12747,N_5123,N_6984);
xnor U12748 (N_12748,N_7817,N_8263);
and U12749 (N_12749,N_9237,N_9929);
nand U12750 (N_12750,N_5540,N_7423);
nand U12751 (N_12751,N_7456,N_8899);
and U12752 (N_12752,N_9086,N_6722);
and U12753 (N_12753,N_6135,N_8269);
nor U12754 (N_12754,N_8348,N_5030);
and U12755 (N_12755,N_6173,N_7619);
and U12756 (N_12756,N_8322,N_5763);
nand U12757 (N_12757,N_5821,N_9481);
nand U12758 (N_12758,N_5178,N_8568);
and U12759 (N_12759,N_6567,N_8311);
nand U12760 (N_12760,N_9403,N_6137);
xor U12761 (N_12761,N_6987,N_8120);
and U12762 (N_12762,N_6045,N_6649);
and U12763 (N_12763,N_7082,N_6302);
and U12764 (N_12764,N_6242,N_7914);
xnor U12765 (N_12765,N_7749,N_5602);
xor U12766 (N_12766,N_6635,N_6625);
and U12767 (N_12767,N_7115,N_9079);
or U12768 (N_12768,N_7156,N_8133);
nand U12769 (N_12769,N_7617,N_6463);
and U12770 (N_12770,N_6422,N_5109);
nor U12771 (N_12771,N_5704,N_6371);
nand U12772 (N_12772,N_7066,N_9859);
and U12773 (N_12773,N_9631,N_6832);
nor U12774 (N_12774,N_8517,N_8076);
and U12775 (N_12775,N_5255,N_5155);
xnor U12776 (N_12776,N_7234,N_5749);
nand U12777 (N_12777,N_9536,N_7330);
or U12778 (N_12778,N_7875,N_6138);
nand U12779 (N_12779,N_9821,N_5253);
and U12780 (N_12780,N_5934,N_5805);
or U12781 (N_12781,N_8306,N_9819);
nand U12782 (N_12782,N_6549,N_9770);
nand U12783 (N_12783,N_9254,N_5204);
nand U12784 (N_12784,N_6488,N_8800);
or U12785 (N_12785,N_6327,N_6487);
nand U12786 (N_12786,N_5019,N_9100);
or U12787 (N_12787,N_9551,N_6888);
xnor U12788 (N_12788,N_9828,N_7190);
nor U12789 (N_12789,N_5965,N_9115);
and U12790 (N_12790,N_8919,N_9295);
and U12791 (N_12791,N_8837,N_6848);
nor U12792 (N_12792,N_5260,N_6934);
xnor U12793 (N_12793,N_9620,N_7645);
xor U12794 (N_12794,N_6911,N_9530);
and U12795 (N_12795,N_6922,N_9172);
nand U12796 (N_12796,N_9492,N_7136);
nor U12797 (N_12797,N_7619,N_8411);
xor U12798 (N_12798,N_7717,N_7243);
and U12799 (N_12799,N_8975,N_8648);
and U12800 (N_12800,N_9909,N_7453);
nor U12801 (N_12801,N_5813,N_7247);
and U12802 (N_12802,N_9181,N_8691);
xnor U12803 (N_12803,N_5102,N_8093);
nor U12804 (N_12804,N_7271,N_7167);
xor U12805 (N_12805,N_9299,N_8074);
nor U12806 (N_12806,N_7397,N_8199);
or U12807 (N_12807,N_5171,N_7850);
nor U12808 (N_12808,N_9742,N_8515);
and U12809 (N_12809,N_9922,N_8204);
and U12810 (N_12810,N_5421,N_8064);
nand U12811 (N_12811,N_7037,N_6303);
or U12812 (N_12812,N_5571,N_7529);
nor U12813 (N_12813,N_5608,N_7954);
nand U12814 (N_12814,N_5421,N_5618);
nor U12815 (N_12815,N_6658,N_5963);
or U12816 (N_12816,N_7702,N_6901);
xnor U12817 (N_12817,N_8949,N_8906);
or U12818 (N_12818,N_5494,N_8749);
xor U12819 (N_12819,N_8200,N_7438);
and U12820 (N_12820,N_7026,N_6282);
nand U12821 (N_12821,N_7770,N_5965);
or U12822 (N_12822,N_6635,N_6426);
nor U12823 (N_12823,N_8357,N_9959);
nor U12824 (N_12824,N_9937,N_6154);
or U12825 (N_12825,N_7536,N_6331);
nand U12826 (N_12826,N_5251,N_7532);
nand U12827 (N_12827,N_6416,N_7448);
xor U12828 (N_12828,N_8568,N_8974);
or U12829 (N_12829,N_5338,N_9765);
nand U12830 (N_12830,N_6868,N_7309);
nand U12831 (N_12831,N_8754,N_7008);
nand U12832 (N_12832,N_9254,N_6801);
or U12833 (N_12833,N_9569,N_7488);
xor U12834 (N_12834,N_5729,N_8548);
or U12835 (N_12835,N_8392,N_5160);
or U12836 (N_12836,N_9536,N_5877);
nand U12837 (N_12837,N_5132,N_9676);
and U12838 (N_12838,N_9580,N_7276);
or U12839 (N_12839,N_7577,N_8629);
or U12840 (N_12840,N_5787,N_6640);
or U12841 (N_12841,N_9716,N_5101);
nor U12842 (N_12842,N_8021,N_9921);
and U12843 (N_12843,N_7173,N_8664);
xor U12844 (N_12844,N_6880,N_7697);
or U12845 (N_12845,N_6322,N_9091);
nor U12846 (N_12846,N_8526,N_5352);
nand U12847 (N_12847,N_9284,N_8970);
and U12848 (N_12848,N_9651,N_8500);
nor U12849 (N_12849,N_7989,N_9824);
nand U12850 (N_12850,N_9642,N_9865);
xor U12851 (N_12851,N_7973,N_7998);
nor U12852 (N_12852,N_5814,N_9707);
nand U12853 (N_12853,N_5597,N_5430);
xor U12854 (N_12854,N_9282,N_9482);
nand U12855 (N_12855,N_8726,N_9463);
nand U12856 (N_12856,N_5650,N_9290);
and U12857 (N_12857,N_8758,N_9189);
nand U12858 (N_12858,N_9650,N_8103);
or U12859 (N_12859,N_6437,N_5569);
nor U12860 (N_12860,N_5638,N_7103);
xnor U12861 (N_12861,N_5821,N_6279);
nand U12862 (N_12862,N_5286,N_7304);
nand U12863 (N_12863,N_7300,N_5912);
nand U12864 (N_12864,N_8095,N_6264);
or U12865 (N_12865,N_5340,N_5590);
xor U12866 (N_12866,N_5934,N_5394);
or U12867 (N_12867,N_5249,N_8769);
nand U12868 (N_12868,N_9262,N_6795);
and U12869 (N_12869,N_6583,N_5233);
and U12870 (N_12870,N_5263,N_6267);
and U12871 (N_12871,N_6243,N_9971);
nand U12872 (N_12872,N_5788,N_6455);
or U12873 (N_12873,N_9299,N_5469);
or U12874 (N_12874,N_5867,N_9289);
or U12875 (N_12875,N_8608,N_5007);
or U12876 (N_12876,N_5849,N_5413);
nor U12877 (N_12877,N_5406,N_5024);
nor U12878 (N_12878,N_7628,N_6184);
nor U12879 (N_12879,N_6547,N_9208);
or U12880 (N_12880,N_8574,N_7031);
nor U12881 (N_12881,N_9005,N_6522);
nand U12882 (N_12882,N_7074,N_7577);
nand U12883 (N_12883,N_7625,N_9567);
or U12884 (N_12884,N_6167,N_6428);
nand U12885 (N_12885,N_5108,N_5220);
or U12886 (N_12886,N_7320,N_7885);
nand U12887 (N_12887,N_8233,N_7604);
nor U12888 (N_12888,N_8254,N_7115);
xnor U12889 (N_12889,N_6182,N_6707);
or U12890 (N_12890,N_8034,N_8899);
or U12891 (N_12891,N_9858,N_6552);
and U12892 (N_12892,N_5712,N_8473);
and U12893 (N_12893,N_9635,N_5321);
nand U12894 (N_12894,N_7477,N_6325);
or U12895 (N_12895,N_8127,N_6468);
nand U12896 (N_12896,N_9651,N_7308);
nand U12897 (N_12897,N_9215,N_8497);
nor U12898 (N_12898,N_8716,N_9446);
or U12899 (N_12899,N_7470,N_8639);
and U12900 (N_12900,N_5374,N_7560);
nor U12901 (N_12901,N_9808,N_8243);
or U12902 (N_12902,N_7230,N_6225);
or U12903 (N_12903,N_8408,N_7135);
nand U12904 (N_12904,N_5364,N_8428);
nor U12905 (N_12905,N_6880,N_8243);
and U12906 (N_12906,N_9187,N_5637);
nand U12907 (N_12907,N_9094,N_7730);
and U12908 (N_12908,N_5910,N_8917);
nor U12909 (N_12909,N_8503,N_7653);
nor U12910 (N_12910,N_7675,N_9505);
xor U12911 (N_12911,N_7125,N_9170);
nand U12912 (N_12912,N_6399,N_8868);
nor U12913 (N_12913,N_5789,N_6612);
xnor U12914 (N_12914,N_7062,N_7401);
xor U12915 (N_12915,N_9080,N_5771);
nand U12916 (N_12916,N_5817,N_7601);
or U12917 (N_12917,N_6561,N_5581);
nand U12918 (N_12918,N_8287,N_5848);
nor U12919 (N_12919,N_5599,N_7925);
and U12920 (N_12920,N_6144,N_6855);
nor U12921 (N_12921,N_6942,N_7954);
nand U12922 (N_12922,N_9041,N_6182);
or U12923 (N_12923,N_6056,N_5927);
or U12924 (N_12924,N_9365,N_8249);
nor U12925 (N_12925,N_5829,N_8410);
and U12926 (N_12926,N_5676,N_9576);
nor U12927 (N_12927,N_5309,N_8652);
nor U12928 (N_12928,N_7331,N_8729);
xor U12929 (N_12929,N_6487,N_9554);
and U12930 (N_12930,N_6354,N_5775);
or U12931 (N_12931,N_7768,N_7280);
nor U12932 (N_12932,N_6465,N_9411);
nor U12933 (N_12933,N_7414,N_8469);
nand U12934 (N_12934,N_6509,N_7208);
nor U12935 (N_12935,N_9131,N_8778);
or U12936 (N_12936,N_7364,N_5978);
and U12937 (N_12937,N_6598,N_6103);
nand U12938 (N_12938,N_8898,N_5293);
nor U12939 (N_12939,N_8473,N_7216);
nand U12940 (N_12940,N_8230,N_5287);
nor U12941 (N_12941,N_6012,N_6950);
nor U12942 (N_12942,N_6606,N_7420);
xnor U12943 (N_12943,N_6798,N_6930);
nand U12944 (N_12944,N_6759,N_5871);
nor U12945 (N_12945,N_5426,N_7109);
xor U12946 (N_12946,N_6876,N_7640);
or U12947 (N_12947,N_9064,N_8735);
nand U12948 (N_12948,N_9289,N_7464);
xnor U12949 (N_12949,N_7984,N_7059);
and U12950 (N_12950,N_8991,N_6753);
nor U12951 (N_12951,N_9311,N_8202);
nor U12952 (N_12952,N_6965,N_6119);
and U12953 (N_12953,N_7111,N_9208);
xor U12954 (N_12954,N_9315,N_9189);
xnor U12955 (N_12955,N_8775,N_5583);
and U12956 (N_12956,N_6382,N_6732);
and U12957 (N_12957,N_9222,N_8667);
nor U12958 (N_12958,N_9757,N_5957);
and U12959 (N_12959,N_6512,N_9537);
xor U12960 (N_12960,N_9409,N_8666);
and U12961 (N_12961,N_6657,N_5746);
or U12962 (N_12962,N_7711,N_8558);
nor U12963 (N_12963,N_6318,N_6723);
and U12964 (N_12964,N_8118,N_8196);
xnor U12965 (N_12965,N_8303,N_8001);
nor U12966 (N_12966,N_5500,N_8330);
xnor U12967 (N_12967,N_8891,N_7818);
and U12968 (N_12968,N_5783,N_5093);
xor U12969 (N_12969,N_7937,N_6683);
nand U12970 (N_12970,N_8281,N_8802);
and U12971 (N_12971,N_9813,N_5221);
nand U12972 (N_12972,N_9921,N_5444);
xnor U12973 (N_12973,N_8094,N_5743);
nand U12974 (N_12974,N_9387,N_8194);
nor U12975 (N_12975,N_8401,N_7282);
nand U12976 (N_12976,N_9623,N_7594);
xor U12977 (N_12977,N_7221,N_6250);
nor U12978 (N_12978,N_5593,N_9629);
and U12979 (N_12979,N_5371,N_7543);
or U12980 (N_12980,N_7679,N_5365);
nand U12981 (N_12981,N_9090,N_8277);
nor U12982 (N_12982,N_5058,N_5012);
nor U12983 (N_12983,N_5737,N_5291);
or U12984 (N_12984,N_6946,N_9154);
nor U12985 (N_12985,N_8534,N_6469);
and U12986 (N_12986,N_9636,N_8571);
xnor U12987 (N_12987,N_9816,N_6983);
and U12988 (N_12988,N_6115,N_6012);
nand U12989 (N_12989,N_5999,N_5235);
or U12990 (N_12990,N_5898,N_5378);
and U12991 (N_12991,N_9547,N_6412);
xor U12992 (N_12992,N_8058,N_6989);
and U12993 (N_12993,N_8868,N_5083);
xor U12994 (N_12994,N_8359,N_9822);
nor U12995 (N_12995,N_8812,N_5399);
and U12996 (N_12996,N_6649,N_6127);
nor U12997 (N_12997,N_8765,N_9376);
and U12998 (N_12998,N_5625,N_7358);
and U12999 (N_12999,N_8755,N_8263);
or U13000 (N_13000,N_7005,N_5799);
nand U13001 (N_13001,N_5752,N_7836);
or U13002 (N_13002,N_7940,N_9590);
nor U13003 (N_13003,N_5185,N_6567);
or U13004 (N_13004,N_7549,N_7478);
and U13005 (N_13005,N_7737,N_6352);
nor U13006 (N_13006,N_8483,N_6592);
xor U13007 (N_13007,N_8172,N_5082);
nand U13008 (N_13008,N_5117,N_5444);
xor U13009 (N_13009,N_8869,N_6727);
or U13010 (N_13010,N_7820,N_8877);
xnor U13011 (N_13011,N_7287,N_9378);
xor U13012 (N_13012,N_7551,N_8690);
or U13013 (N_13013,N_9128,N_8131);
or U13014 (N_13014,N_6869,N_9931);
nor U13015 (N_13015,N_8537,N_9944);
and U13016 (N_13016,N_7808,N_5289);
xor U13017 (N_13017,N_8605,N_7318);
nor U13018 (N_13018,N_7465,N_6312);
and U13019 (N_13019,N_6950,N_9753);
and U13020 (N_13020,N_8109,N_6773);
nand U13021 (N_13021,N_5568,N_9893);
nor U13022 (N_13022,N_7607,N_7992);
nor U13023 (N_13023,N_5420,N_5203);
or U13024 (N_13024,N_9575,N_5140);
nor U13025 (N_13025,N_8503,N_7669);
nand U13026 (N_13026,N_9372,N_9867);
xor U13027 (N_13027,N_7280,N_8065);
or U13028 (N_13028,N_8357,N_6127);
or U13029 (N_13029,N_9874,N_9420);
nor U13030 (N_13030,N_7646,N_8060);
nand U13031 (N_13031,N_6574,N_6515);
xnor U13032 (N_13032,N_7780,N_7136);
and U13033 (N_13033,N_7371,N_6189);
nor U13034 (N_13034,N_5832,N_9430);
or U13035 (N_13035,N_5965,N_5286);
and U13036 (N_13036,N_9981,N_6839);
nand U13037 (N_13037,N_6703,N_6049);
nor U13038 (N_13038,N_9103,N_6398);
nand U13039 (N_13039,N_5834,N_7133);
nand U13040 (N_13040,N_6852,N_9413);
nand U13041 (N_13041,N_7684,N_8818);
nor U13042 (N_13042,N_9408,N_8392);
and U13043 (N_13043,N_5014,N_9749);
or U13044 (N_13044,N_7259,N_5011);
xor U13045 (N_13045,N_7559,N_6156);
or U13046 (N_13046,N_8663,N_8977);
nand U13047 (N_13047,N_7130,N_9503);
or U13048 (N_13048,N_5871,N_5083);
xnor U13049 (N_13049,N_9717,N_5444);
xnor U13050 (N_13050,N_6567,N_5829);
xnor U13051 (N_13051,N_7992,N_5132);
nand U13052 (N_13052,N_9492,N_6236);
and U13053 (N_13053,N_5686,N_7019);
or U13054 (N_13054,N_6407,N_8827);
and U13055 (N_13055,N_5533,N_8740);
nor U13056 (N_13056,N_6206,N_7022);
or U13057 (N_13057,N_5009,N_9896);
xor U13058 (N_13058,N_7710,N_6412);
xnor U13059 (N_13059,N_9049,N_7093);
nor U13060 (N_13060,N_7570,N_9443);
xnor U13061 (N_13061,N_8933,N_8027);
and U13062 (N_13062,N_5635,N_7037);
and U13063 (N_13063,N_6652,N_8282);
and U13064 (N_13064,N_5727,N_5618);
xor U13065 (N_13065,N_9317,N_9417);
or U13066 (N_13066,N_9315,N_7161);
or U13067 (N_13067,N_7215,N_7504);
nor U13068 (N_13068,N_8377,N_6698);
or U13069 (N_13069,N_9445,N_9206);
nor U13070 (N_13070,N_8563,N_9158);
and U13071 (N_13071,N_8637,N_8444);
or U13072 (N_13072,N_8336,N_5652);
xnor U13073 (N_13073,N_5711,N_7020);
and U13074 (N_13074,N_8170,N_8368);
or U13075 (N_13075,N_7991,N_9051);
nor U13076 (N_13076,N_9371,N_8105);
nand U13077 (N_13077,N_8440,N_9806);
nand U13078 (N_13078,N_9969,N_5160);
nand U13079 (N_13079,N_6496,N_5055);
nand U13080 (N_13080,N_9102,N_5974);
nand U13081 (N_13081,N_5480,N_8642);
and U13082 (N_13082,N_6156,N_8635);
or U13083 (N_13083,N_7565,N_8427);
and U13084 (N_13084,N_6838,N_6660);
nor U13085 (N_13085,N_7448,N_7568);
or U13086 (N_13086,N_6636,N_6503);
and U13087 (N_13087,N_7061,N_7684);
and U13088 (N_13088,N_6837,N_6112);
or U13089 (N_13089,N_8251,N_7180);
xor U13090 (N_13090,N_9719,N_6945);
nand U13091 (N_13091,N_8695,N_7812);
nor U13092 (N_13092,N_9100,N_7957);
nand U13093 (N_13093,N_8137,N_7554);
xor U13094 (N_13094,N_5516,N_7275);
or U13095 (N_13095,N_7672,N_6336);
nand U13096 (N_13096,N_6239,N_8842);
or U13097 (N_13097,N_7444,N_9889);
nor U13098 (N_13098,N_9945,N_5151);
nor U13099 (N_13099,N_7085,N_5655);
xnor U13100 (N_13100,N_5253,N_6673);
nand U13101 (N_13101,N_6215,N_5704);
and U13102 (N_13102,N_5606,N_5957);
nor U13103 (N_13103,N_6794,N_8489);
or U13104 (N_13104,N_6838,N_6318);
nand U13105 (N_13105,N_7280,N_5775);
nand U13106 (N_13106,N_6312,N_5158);
nor U13107 (N_13107,N_8821,N_6208);
nand U13108 (N_13108,N_5306,N_8494);
xnor U13109 (N_13109,N_9422,N_5153);
and U13110 (N_13110,N_7334,N_5771);
nand U13111 (N_13111,N_7855,N_8352);
and U13112 (N_13112,N_5058,N_7971);
nor U13113 (N_13113,N_8828,N_8073);
nand U13114 (N_13114,N_7696,N_9889);
or U13115 (N_13115,N_8667,N_9515);
or U13116 (N_13116,N_7486,N_8058);
nor U13117 (N_13117,N_8553,N_9816);
xor U13118 (N_13118,N_9148,N_8202);
nand U13119 (N_13119,N_7010,N_5217);
xnor U13120 (N_13120,N_6428,N_7219);
xnor U13121 (N_13121,N_8925,N_9348);
and U13122 (N_13122,N_5977,N_5649);
nand U13123 (N_13123,N_6919,N_5866);
xnor U13124 (N_13124,N_9744,N_9556);
nor U13125 (N_13125,N_5954,N_9303);
nand U13126 (N_13126,N_9441,N_9872);
xnor U13127 (N_13127,N_7172,N_9395);
xnor U13128 (N_13128,N_5314,N_9680);
xnor U13129 (N_13129,N_5188,N_8049);
nand U13130 (N_13130,N_5280,N_5525);
or U13131 (N_13131,N_8673,N_6438);
and U13132 (N_13132,N_9556,N_7224);
and U13133 (N_13133,N_5396,N_9557);
nor U13134 (N_13134,N_8598,N_9267);
nand U13135 (N_13135,N_6137,N_7895);
nor U13136 (N_13136,N_9531,N_8988);
or U13137 (N_13137,N_5220,N_9706);
nor U13138 (N_13138,N_6992,N_5805);
nor U13139 (N_13139,N_7125,N_9604);
nor U13140 (N_13140,N_7074,N_7146);
nand U13141 (N_13141,N_5418,N_8337);
or U13142 (N_13142,N_8313,N_7345);
nor U13143 (N_13143,N_6495,N_9237);
and U13144 (N_13144,N_5818,N_6061);
nand U13145 (N_13145,N_9444,N_5824);
nor U13146 (N_13146,N_7475,N_8194);
and U13147 (N_13147,N_5050,N_7650);
nor U13148 (N_13148,N_7269,N_8298);
nor U13149 (N_13149,N_7426,N_7029);
nand U13150 (N_13150,N_8561,N_7695);
nor U13151 (N_13151,N_7093,N_6660);
xor U13152 (N_13152,N_8620,N_9738);
nor U13153 (N_13153,N_6939,N_5504);
nand U13154 (N_13154,N_7074,N_5197);
nor U13155 (N_13155,N_7073,N_7684);
nand U13156 (N_13156,N_9504,N_5754);
and U13157 (N_13157,N_9574,N_5755);
and U13158 (N_13158,N_7393,N_5278);
xnor U13159 (N_13159,N_5516,N_9127);
or U13160 (N_13160,N_6189,N_8564);
or U13161 (N_13161,N_9839,N_9744);
or U13162 (N_13162,N_9602,N_9400);
or U13163 (N_13163,N_9989,N_6862);
xnor U13164 (N_13164,N_7347,N_9670);
nand U13165 (N_13165,N_5207,N_5056);
nand U13166 (N_13166,N_8987,N_9876);
nor U13167 (N_13167,N_7185,N_9976);
nor U13168 (N_13168,N_8226,N_6089);
or U13169 (N_13169,N_8393,N_5981);
nor U13170 (N_13170,N_9971,N_9336);
or U13171 (N_13171,N_7920,N_9252);
or U13172 (N_13172,N_9815,N_7504);
and U13173 (N_13173,N_8108,N_9912);
xor U13174 (N_13174,N_5246,N_9135);
nand U13175 (N_13175,N_8083,N_7115);
xor U13176 (N_13176,N_8312,N_8093);
and U13177 (N_13177,N_7249,N_6110);
or U13178 (N_13178,N_6802,N_8290);
xor U13179 (N_13179,N_8986,N_6328);
or U13180 (N_13180,N_8696,N_7255);
and U13181 (N_13181,N_7351,N_9008);
nand U13182 (N_13182,N_9334,N_8029);
or U13183 (N_13183,N_7776,N_6757);
nand U13184 (N_13184,N_5514,N_7888);
or U13185 (N_13185,N_9924,N_5332);
xnor U13186 (N_13186,N_8329,N_7594);
or U13187 (N_13187,N_7364,N_8352);
nand U13188 (N_13188,N_6905,N_9041);
or U13189 (N_13189,N_8704,N_9042);
nand U13190 (N_13190,N_7894,N_6830);
nand U13191 (N_13191,N_7191,N_6487);
nor U13192 (N_13192,N_5513,N_6266);
or U13193 (N_13193,N_7115,N_8258);
xor U13194 (N_13194,N_6542,N_6987);
and U13195 (N_13195,N_6729,N_6910);
nand U13196 (N_13196,N_9782,N_9516);
or U13197 (N_13197,N_6640,N_6061);
nand U13198 (N_13198,N_6415,N_8965);
or U13199 (N_13199,N_7151,N_8842);
xor U13200 (N_13200,N_8392,N_9855);
or U13201 (N_13201,N_9920,N_8279);
xor U13202 (N_13202,N_9783,N_8491);
nor U13203 (N_13203,N_5938,N_7943);
or U13204 (N_13204,N_8411,N_5721);
or U13205 (N_13205,N_6258,N_9012);
or U13206 (N_13206,N_9415,N_8115);
or U13207 (N_13207,N_7375,N_8022);
nand U13208 (N_13208,N_5122,N_5464);
or U13209 (N_13209,N_5797,N_8994);
xor U13210 (N_13210,N_9535,N_7980);
nor U13211 (N_13211,N_5631,N_5938);
xnor U13212 (N_13212,N_7002,N_9521);
and U13213 (N_13213,N_5401,N_9474);
or U13214 (N_13214,N_7417,N_9002);
nand U13215 (N_13215,N_5467,N_8372);
nand U13216 (N_13216,N_8331,N_6802);
nand U13217 (N_13217,N_5072,N_6752);
and U13218 (N_13218,N_7962,N_7095);
xor U13219 (N_13219,N_9420,N_6116);
or U13220 (N_13220,N_7455,N_5983);
or U13221 (N_13221,N_5585,N_7669);
nand U13222 (N_13222,N_5269,N_9103);
nor U13223 (N_13223,N_5444,N_9441);
nand U13224 (N_13224,N_7140,N_9370);
nor U13225 (N_13225,N_5781,N_9171);
xor U13226 (N_13226,N_9330,N_7802);
nand U13227 (N_13227,N_6128,N_5509);
nand U13228 (N_13228,N_7903,N_7037);
or U13229 (N_13229,N_7594,N_5581);
nand U13230 (N_13230,N_5815,N_6004);
nand U13231 (N_13231,N_8187,N_6266);
or U13232 (N_13232,N_7330,N_6458);
nor U13233 (N_13233,N_9429,N_7672);
or U13234 (N_13234,N_5405,N_7235);
or U13235 (N_13235,N_9202,N_5940);
xor U13236 (N_13236,N_9215,N_9931);
or U13237 (N_13237,N_5383,N_9258);
nand U13238 (N_13238,N_9344,N_5000);
or U13239 (N_13239,N_8195,N_5801);
or U13240 (N_13240,N_8630,N_8925);
or U13241 (N_13241,N_8188,N_8962);
nor U13242 (N_13242,N_5411,N_8766);
nor U13243 (N_13243,N_9033,N_7941);
or U13244 (N_13244,N_5061,N_5505);
and U13245 (N_13245,N_5201,N_8515);
nand U13246 (N_13246,N_6029,N_5666);
and U13247 (N_13247,N_9080,N_7643);
or U13248 (N_13248,N_5878,N_7753);
and U13249 (N_13249,N_6621,N_7940);
nand U13250 (N_13250,N_7433,N_5497);
and U13251 (N_13251,N_8039,N_9561);
xor U13252 (N_13252,N_8324,N_6541);
or U13253 (N_13253,N_7707,N_8959);
xor U13254 (N_13254,N_8777,N_5858);
or U13255 (N_13255,N_8750,N_6639);
nand U13256 (N_13256,N_8408,N_5777);
nand U13257 (N_13257,N_5035,N_6340);
xor U13258 (N_13258,N_6516,N_8645);
xnor U13259 (N_13259,N_5590,N_6151);
nor U13260 (N_13260,N_7398,N_9236);
nor U13261 (N_13261,N_8370,N_5282);
and U13262 (N_13262,N_8652,N_9872);
nor U13263 (N_13263,N_6588,N_7319);
or U13264 (N_13264,N_8213,N_6096);
xnor U13265 (N_13265,N_5000,N_5193);
or U13266 (N_13266,N_9198,N_8676);
xnor U13267 (N_13267,N_5407,N_6249);
nor U13268 (N_13268,N_8603,N_7691);
nand U13269 (N_13269,N_8158,N_6654);
xnor U13270 (N_13270,N_8686,N_8836);
nor U13271 (N_13271,N_6006,N_7310);
nor U13272 (N_13272,N_6319,N_8359);
or U13273 (N_13273,N_8245,N_9074);
or U13274 (N_13274,N_5670,N_8661);
and U13275 (N_13275,N_9509,N_7274);
or U13276 (N_13276,N_5791,N_7363);
nor U13277 (N_13277,N_7646,N_8362);
nand U13278 (N_13278,N_6749,N_9911);
or U13279 (N_13279,N_7472,N_6558);
nor U13280 (N_13280,N_9377,N_5111);
nand U13281 (N_13281,N_8781,N_7410);
xnor U13282 (N_13282,N_8917,N_5032);
and U13283 (N_13283,N_6616,N_8584);
and U13284 (N_13284,N_6836,N_8077);
nor U13285 (N_13285,N_8044,N_5572);
xnor U13286 (N_13286,N_6057,N_9250);
or U13287 (N_13287,N_5205,N_6841);
and U13288 (N_13288,N_5505,N_7231);
xnor U13289 (N_13289,N_5478,N_9936);
xnor U13290 (N_13290,N_5610,N_8033);
or U13291 (N_13291,N_7549,N_6119);
nand U13292 (N_13292,N_5231,N_9010);
nand U13293 (N_13293,N_6111,N_7705);
or U13294 (N_13294,N_6499,N_5282);
xnor U13295 (N_13295,N_7954,N_9332);
nor U13296 (N_13296,N_5645,N_7685);
xnor U13297 (N_13297,N_9948,N_7863);
or U13298 (N_13298,N_5008,N_7552);
and U13299 (N_13299,N_5143,N_6101);
or U13300 (N_13300,N_5657,N_5206);
nand U13301 (N_13301,N_8249,N_9590);
nand U13302 (N_13302,N_7784,N_9320);
xor U13303 (N_13303,N_5831,N_7149);
nand U13304 (N_13304,N_5555,N_7230);
xnor U13305 (N_13305,N_6099,N_7957);
nor U13306 (N_13306,N_9911,N_6809);
or U13307 (N_13307,N_7333,N_5434);
and U13308 (N_13308,N_5092,N_9925);
or U13309 (N_13309,N_7856,N_9793);
nand U13310 (N_13310,N_6171,N_7817);
nor U13311 (N_13311,N_6582,N_5826);
nand U13312 (N_13312,N_5170,N_7164);
or U13313 (N_13313,N_7531,N_5249);
nand U13314 (N_13314,N_6443,N_5287);
or U13315 (N_13315,N_6764,N_5396);
or U13316 (N_13316,N_6876,N_5691);
nor U13317 (N_13317,N_7444,N_5610);
nor U13318 (N_13318,N_7148,N_5806);
or U13319 (N_13319,N_7962,N_9577);
or U13320 (N_13320,N_6263,N_6640);
nor U13321 (N_13321,N_7146,N_9817);
or U13322 (N_13322,N_6441,N_6925);
nor U13323 (N_13323,N_9199,N_7216);
nor U13324 (N_13324,N_6987,N_5595);
nor U13325 (N_13325,N_8837,N_8701);
nor U13326 (N_13326,N_9530,N_9858);
nor U13327 (N_13327,N_5774,N_5129);
and U13328 (N_13328,N_9294,N_5907);
nor U13329 (N_13329,N_8421,N_7032);
and U13330 (N_13330,N_6566,N_8523);
or U13331 (N_13331,N_5360,N_9240);
nor U13332 (N_13332,N_6908,N_9683);
or U13333 (N_13333,N_8772,N_8102);
xnor U13334 (N_13334,N_9305,N_5260);
nand U13335 (N_13335,N_6575,N_9710);
nor U13336 (N_13336,N_6848,N_9077);
or U13337 (N_13337,N_9274,N_7812);
xor U13338 (N_13338,N_7213,N_7489);
nor U13339 (N_13339,N_5291,N_8254);
nor U13340 (N_13340,N_7072,N_9374);
nor U13341 (N_13341,N_7196,N_5924);
xnor U13342 (N_13342,N_8364,N_5788);
nor U13343 (N_13343,N_6337,N_5223);
and U13344 (N_13344,N_6004,N_6338);
nor U13345 (N_13345,N_6341,N_7758);
and U13346 (N_13346,N_6263,N_7563);
and U13347 (N_13347,N_9307,N_8037);
nand U13348 (N_13348,N_5562,N_6294);
or U13349 (N_13349,N_6698,N_8487);
and U13350 (N_13350,N_6259,N_5234);
and U13351 (N_13351,N_5335,N_8116);
or U13352 (N_13352,N_5554,N_6984);
nor U13353 (N_13353,N_9038,N_9466);
xor U13354 (N_13354,N_6108,N_9112);
and U13355 (N_13355,N_5429,N_9009);
nand U13356 (N_13356,N_6794,N_9706);
nand U13357 (N_13357,N_7804,N_8277);
and U13358 (N_13358,N_5843,N_6155);
nor U13359 (N_13359,N_8298,N_6091);
nor U13360 (N_13360,N_8678,N_9787);
nand U13361 (N_13361,N_6419,N_9670);
xnor U13362 (N_13362,N_7294,N_5962);
nor U13363 (N_13363,N_8243,N_7444);
xnor U13364 (N_13364,N_6657,N_6999);
nand U13365 (N_13365,N_8794,N_8651);
and U13366 (N_13366,N_7508,N_9252);
and U13367 (N_13367,N_7262,N_8042);
nor U13368 (N_13368,N_6503,N_9126);
and U13369 (N_13369,N_5637,N_7547);
xnor U13370 (N_13370,N_8119,N_7473);
and U13371 (N_13371,N_7158,N_5889);
nor U13372 (N_13372,N_9296,N_7897);
and U13373 (N_13373,N_7719,N_6198);
or U13374 (N_13374,N_6269,N_8290);
xor U13375 (N_13375,N_6157,N_9527);
xor U13376 (N_13376,N_7515,N_9963);
xnor U13377 (N_13377,N_5634,N_5051);
and U13378 (N_13378,N_5583,N_5969);
or U13379 (N_13379,N_8995,N_8981);
or U13380 (N_13380,N_9987,N_5015);
xor U13381 (N_13381,N_8078,N_5529);
xor U13382 (N_13382,N_5751,N_5504);
or U13383 (N_13383,N_9542,N_7684);
nand U13384 (N_13384,N_9828,N_6578);
or U13385 (N_13385,N_6981,N_7600);
nand U13386 (N_13386,N_7934,N_9940);
xor U13387 (N_13387,N_8558,N_8129);
nor U13388 (N_13388,N_5191,N_5006);
nand U13389 (N_13389,N_9984,N_7954);
nand U13390 (N_13390,N_5383,N_8250);
or U13391 (N_13391,N_8153,N_7700);
or U13392 (N_13392,N_7779,N_7409);
nand U13393 (N_13393,N_7328,N_6596);
or U13394 (N_13394,N_5078,N_9193);
nand U13395 (N_13395,N_5640,N_5674);
nor U13396 (N_13396,N_9539,N_9711);
nor U13397 (N_13397,N_9638,N_8637);
and U13398 (N_13398,N_5013,N_6895);
and U13399 (N_13399,N_6703,N_7945);
and U13400 (N_13400,N_5604,N_5176);
nor U13401 (N_13401,N_7951,N_6364);
nand U13402 (N_13402,N_6965,N_6550);
and U13403 (N_13403,N_7679,N_8521);
nor U13404 (N_13404,N_7728,N_6718);
nand U13405 (N_13405,N_6630,N_5304);
and U13406 (N_13406,N_7182,N_6622);
or U13407 (N_13407,N_5992,N_5335);
or U13408 (N_13408,N_8889,N_6978);
nand U13409 (N_13409,N_8643,N_6642);
nand U13410 (N_13410,N_7512,N_7625);
nand U13411 (N_13411,N_9704,N_6429);
and U13412 (N_13412,N_8732,N_5199);
xnor U13413 (N_13413,N_9065,N_5379);
nand U13414 (N_13414,N_5368,N_9103);
nand U13415 (N_13415,N_9749,N_9885);
nand U13416 (N_13416,N_9390,N_8549);
and U13417 (N_13417,N_6270,N_7380);
and U13418 (N_13418,N_9648,N_6588);
nor U13419 (N_13419,N_7153,N_7285);
nand U13420 (N_13420,N_7915,N_9925);
xnor U13421 (N_13421,N_5044,N_9698);
nand U13422 (N_13422,N_9361,N_7484);
or U13423 (N_13423,N_6817,N_6653);
and U13424 (N_13424,N_8765,N_8364);
and U13425 (N_13425,N_8660,N_9145);
and U13426 (N_13426,N_8444,N_7874);
nor U13427 (N_13427,N_5019,N_9412);
xor U13428 (N_13428,N_5829,N_8003);
xor U13429 (N_13429,N_6344,N_5631);
nor U13430 (N_13430,N_6228,N_8619);
xor U13431 (N_13431,N_7887,N_8699);
nand U13432 (N_13432,N_9409,N_5343);
nand U13433 (N_13433,N_7860,N_6747);
nor U13434 (N_13434,N_6016,N_7364);
or U13435 (N_13435,N_5372,N_7071);
nor U13436 (N_13436,N_7487,N_5501);
or U13437 (N_13437,N_5915,N_6229);
xor U13438 (N_13438,N_5129,N_8060);
nor U13439 (N_13439,N_6141,N_5030);
nor U13440 (N_13440,N_7485,N_7707);
nor U13441 (N_13441,N_8559,N_6133);
xor U13442 (N_13442,N_6047,N_9698);
nand U13443 (N_13443,N_6725,N_5900);
nor U13444 (N_13444,N_9149,N_9178);
nor U13445 (N_13445,N_5307,N_7227);
or U13446 (N_13446,N_9973,N_8873);
xnor U13447 (N_13447,N_5139,N_9587);
and U13448 (N_13448,N_8990,N_7373);
nor U13449 (N_13449,N_9654,N_5063);
nor U13450 (N_13450,N_9435,N_9676);
nor U13451 (N_13451,N_9680,N_8388);
nor U13452 (N_13452,N_7109,N_8115);
and U13453 (N_13453,N_6127,N_8881);
or U13454 (N_13454,N_8765,N_5840);
xor U13455 (N_13455,N_8714,N_5478);
or U13456 (N_13456,N_6518,N_8727);
or U13457 (N_13457,N_9339,N_5094);
nand U13458 (N_13458,N_9011,N_5415);
or U13459 (N_13459,N_9829,N_6426);
nand U13460 (N_13460,N_7161,N_8361);
or U13461 (N_13461,N_6186,N_9622);
and U13462 (N_13462,N_5405,N_9606);
nor U13463 (N_13463,N_9806,N_7529);
or U13464 (N_13464,N_9925,N_9427);
nor U13465 (N_13465,N_7682,N_9906);
or U13466 (N_13466,N_7621,N_9862);
and U13467 (N_13467,N_8036,N_9274);
and U13468 (N_13468,N_6712,N_7373);
xor U13469 (N_13469,N_7835,N_7167);
xnor U13470 (N_13470,N_5953,N_7312);
or U13471 (N_13471,N_7845,N_7115);
xnor U13472 (N_13472,N_5873,N_7751);
nor U13473 (N_13473,N_8153,N_9838);
or U13474 (N_13474,N_8198,N_6446);
or U13475 (N_13475,N_8101,N_6459);
or U13476 (N_13476,N_6853,N_8869);
or U13477 (N_13477,N_7921,N_5407);
xor U13478 (N_13478,N_5890,N_9384);
nor U13479 (N_13479,N_6286,N_7980);
nor U13480 (N_13480,N_8734,N_5876);
and U13481 (N_13481,N_7443,N_7274);
and U13482 (N_13482,N_7497,N_5037);
xor U13483 (N_13483,N_9755,N_8129);
or U13484 (N_13484,N_9713,N_5395);
xnor U13485 (N_13485,N_7614,N_5811);
nor U13486 (N_13486,N_7698,N_6714);
and U13487 (N_13487,N_9774,N_9406);
xor U13488 (N_13488,N_5750,N_8243);
and U13489 (N_13489,N_9365,N_8105);
nand U13490 (N_13490,N_6716,N_8527);
nor U13491 (N_13491,N_5691,N_9757);
nand U13492 (N_13492,N_6924,N_9746);
and U13493 (N_13493,N_8128,N_5619);
nor U13494 (N_13494,N_8926,N_8036);
or U13495 (N_13495,N_9817,N_7267);
xnor U13496 (N_13496,N_6890,N_5572);
or U13497 (N_13497,N_6761,N_7447);
and U13498 (N_13498,N_6259,N_7214);
or U13499 (N_13499,N_7112,N_8526);
nand U13500 (N_13500,N_6512,N_6208);
and U13501 (N_13501,N_7153,N_6927);
nor U13502 (N_13502,N_5284,N_8805);
and U13503 (N_13503,N_6075,N_7884);
or U13504 (N_13504,N_6286,N_5597);
xor U13505 (N_13505,N_7704,N_9573);
and U13506 (N_13506,N_9750,N_6564);
or U13507 (N_13507,N_9934,N_9079);
xnor U13508 (N_13508,N_8901,N_5593);
or U13509 (N_13509,N_7778,N_9333);
or U13510 (N_13510,N_8321,N_5588);
nor U13511 (N_13511,N_5249,N_8920);
nand U13512 (N_13512,N_8011,N_5885);
nand U13513 (N_13513,N_8497,N_9799);
and U13514 (N_13514,N_8250,N_9516);
or U13515 (N_13515,N_6223,N_6807);
or U13516 (N_13516,N_6941,N_6684);
nor U13517 (N_13517,N_9880,N_6300);
nand U13518 (N_13518,N_7163,N_7790);
or U13519 (N_13519,N_5492,N_7976);
nand U13520 (N_13520,N_7814,N_7809);
nand U13521 (N_13521,N_7673,N_6721);
or U13522 (N_13522,N_7404,N_6089);
xnor U13523 (N_13523,N_6551,N_8692);
nor U13524 (N_13524,N_7225,N_8678);
and U13525 (N_13525,N_9606,N_6700);
nand U13526 (N_13526,N_8283,N_9340);
or U13527 (N_13527,N_6189,N_7891);
and U13528 (N_13528,N_8638,N_9224);
or U13529 (N_13529,N_8371,N_7952);
nor U13530 (N_13530,N_5410,N_5830);
xor U13531 (N_13531,N_8068,N_6456);
nand U13532 (N_13532,N_9918,N_5048);
nand U13533 (N_13533,N_5691,N_8457);
nand U13534 (N_13534,N_7944,N_9473);
nand U13535 (N_13535,N_5723,N_8008);
xnor U13536 (N_13536,N_9123,N_6580);
and U13537 (N_13537,N_9403,N_7448);
xnor U13538 (N_13538,N_7696,N_5927);
or U13539 (N_13539,N_5209,N_5995);
or U13540 (N_13540,N_6443,N_7136);
nor U13541 (N_13541,N_7179,N_7550);
nand U13542 (N_13542,N_8233,N_6810);
or U13543 (N_13543,N_7249,N_6166);
and U13544 (N_13544,N_9028,N_8819);
xor U13545 (N_13545,N_5174,N_5659);
xnor U13546 (N_13546,N_7677,N_8827);
and U13547 (N_13547,N_8389,N_6706);
nand U13548 (N_13548,N_7388,N_5043);
nor U13549 (N_13549,N_9789,N_5101);
and U13550 (N_13550,N_8575,N_6094);
nand U13551 (N_13551,N_5498,N_8470);
xor U13552 (N_13552,N_5342,N_5253);
xor U13553 (N_13553,N_8405,N_9683);
nor U13554 (N_13554,N_6302,N_8823);
or U13555 (N_13555,N_5097,N_7527);
and U13556 (N_13556,N_7623,N_9615);
xor U13557 (N_13557,N_9200,N_7345);
xnor U13558 (N_13558,N_7195,N_9982);
xnor U13559 (N_13559,N_8609,N_8577);
nand U13560 (N_13560,N_9355,N_6144);
nor U13561 (N_13561,N_7079,N_5335);
nor U13562 (N_13562,N_9089,N_9401);
nor U13563 (N_13563,N_8997,N_6154);
nand U13564 (N_13564,N_6669,N_9570);
nor U13565 (N_13565,N_6115,N_9208);
nor U13566 (N_13566,N_6532,N_5042);
nand U13567 (N_13567,N_9049,N_9567);
xor U13568 (N_13568,N_7691,N_7290);
and U13569 (N_13569,N_6323,N_9958);
xor U13570 (N_13570,N_9184,N_6611);
nand U13571 (N_13571,N_5683,N_8772);
nand U13572 (N_13572,N_5572,N_6276);
nand U13573 (N_13573,N_5148,N_8876);
and U13574 (N_13574,N_9398,N_8502);
or U13575 (N_13575,N_7191,N_7122);
nor U13576 (N_13576,N_7361,N_7887);
xor U13577 (N_13577,N_8169,N_7293);
nor U13578 (N_13578,N_9206,N_9463);
nor U13579 (N_13579,N_6359,N_9170);
xor U13580 (N_13580,N_6323,N_6494);
nor U13581 (N_13581,N_7014,N_9001);
and U13582 (N_13582,N_9011,N_7897);
xnor U13583 (N_13583,N_7236,N_5159);
xor U13584 (N_13584,N_9859,N_8646);
nand U13585 (N_13585,N_5327,N_9568);
nand U13586 (N_13586,N_9001,N_8807);
and U13587 (N_13587,N_7447,N_7271);
xnor U13588 (N_13588,N_6865,N_5108);
nor U13589 (N_13589,N_9265,N_5281);
xor U13590 (N_13590,N_6178,N_5841);
nand U13591 (N_13591,N_5613,N_7303);
nor U13592 (N_13592,N_7838,N_6243);
or U13593 (N_13593,N_7710,N_5517);
or U13594 (N_13594,N_9274,N_9514);
xnor U13595 (N_13595,N_7627,N_8884);
nand U13596 (N_13596,N_8710,N_6772);
nand U13597 (N_13597,N_5618,N_5622);
nor U13598 (N_13598,N_7902,N_7089);
and U13599 (N_13599,N_6057,N_7311);
nand U13600 (N_13600,N_5550,N_9057);
and U13601 (N_13601,N_8293,N_9606);
or U13602 (N_13602,N_5335,N_7885);
nor U13603 (N_13603,N_8675,N_7685);
and U13604 (N_13604,N_8261,N_5591);
and U13605 (N_13605,N_6341,N_5144);
nand U13606 (N_13606,N_5105,N_7576);
nand U13607 (N_13607,N_9862,N_7079);
xor U13608 (N_13608,N_8985,N_6642);
nand U13609 (N_13609,N_9421,N_9492);
nand U13610 (N_13610,N_8449,N_6878);
and U13611 (N_13611,N_9389,N_6624);
xnor U13612 (N_13612,N_5967,N_5049);
or U13613 (N_13613,N_8515,N_9992);
nand U13614 (N_13614,N_6784,N_9489);
nand U13615 (N_13615,N_7099,N_7102);
and U13616 (N_13616,N_9864,N_8050);
or U13617 (N_13617,N_8503,N_9124);
nand U13618 (N_13618,N_5054,N_7442);
nor U13619 (N_13619,N_6896,N_6039);
nor U13620 (N_13620,N_6699,N_6054);
or U13621 (N_13621,N_9005,N_7053);
nand U13622 (N_13622,N_6506,N_8842);
and U13623 (N_13623,N_6281,N_7717);
xnor U13624 (N_13624,N_7674,N_8510);
xnor U13625 (N_13625,N_5092,N_6409);
and U13626 (N_13626,N_7370,N_9139);
nand U13627 (N_13627,N_8186,N_5888);
nand U13628 (N_13628,N_8855,N_5662);
nor U13629 (N_13629,N_8475,N_7431);
or U13630 (N_13630,N_9353,N_5916);
nand U13631 (N_13631,N_9724,N_9081);
nor U13632 (N_13632,N_7101,N_8507);
and U13633 (N_13633,N_7649,N_6465);
or U13634 (N_13634,N_7754,N_7460);
and U13635 (N_13635,N_9579,N_7335);
and U13636 (N_13636,N_9244,N_7842);
and U13637 (N_13637,N_8227,N_9654);
nand U13638 (N_13638,N_7398,N_8890);
nand U13639 (N_13639,N_7378,N_6430);
or U13640 (N_13640,N_7490,N_6626);
and U13641 (N_13641,N_6201,N_6560);
or U13642 (N_13642,N_9133,N_7664);
and U13643 (N_13643,N_9855,N_6535);
or U13644 (N_13644,N_8530,N_9519);
xor U13645 (N_13645,N_8479,N_8320);
nand U13646 (N_13646,N_5638,N_9286);
and U13647 (N_13647,N_5173,N_8088);
xnor U13648 (N_13648,N_8780,N_7259);
xnor U13649 (N_13649,N_5385,N_6147);
nand U13650 (N_13650,N_7703,N_9618);
and U13651 (N_13651,N_8049,N_6083);
nor U13652 (N_13652,N_8338,N_9202);
nor U13653 (N_13653,N_9323,N_5833);
nand U13654 (N_13654,N_8512,N_8019);
and U13655 (N_13655,N_7742,N_6414);
or U13656 (N_13656,N_6798,N_7592);
xor U13657 (N_13657,N_7525,N_6087);
or U13658 (N_13658,N_5731,N_9869);
nand U13659 (N_13659,N_7872,N_6004);
or U13660 (N_13660,N_9228,N_8926);
or U13661 (N_13661,N_5706,N_9920);
nor U13662 (N_13662,N_9418,N_7257);
nand U13663 (N_13663,N_5437,N_6822);
xnor U13664 (N_13664,N_6927,N_5930);
nand U13665 (N_13665,N_9608,N_7311);
nor U13666 (N_13666,N_5405,N_7405);
and U13667 (N_13667,N_8707,N_5179);
nand U13668 (N_13668,N_9667,N_6918);
or U13669 (N_13669,N_9437,N_7423);
and U13670 (N_13670,N_5898,N_5934);
nor U13671 (N_13671,N_8674,N_6945);
nand U13672 (N_13672,N_5736,N_6869);
xor U13673 (N_13673,N_6894,N_9017);
xnor U13674 (N_13674,N_9219,N_9258);
or U13675 (N_13675,N_8631,N_7570);
or U13676 (N_13676,N_7824,N_7678);
nor U13677 (N_13677,N_7941,N_9459);
xnor U13678 (N_13678,N_8953,N_7125);
and U13679 (N_13679,N_6974,N_6264);
nor U13680 (N_13680,N_7952,N_6438);
nand U13681 (N_13681,N_6001,N_8579);
or U13682 (N_13682,N_6462,N_6463);
and U13683 (N_13683,N_9081,N_7769);
nor U13684 (N_13684,N_5355,N_9490);
nand U13685 (N_13685,N_7196,N_7886);
or U13686 (N_13686,N_8744,N_7745);
or U13687 (N_13687,N_8191,N_5460);
nand U13688 (N_13688,N_9343,N_5202);
or U13689 (N_13689,N_5660,N_6632);
xor U13690 (N_13690,N_6253,N_5217);
nor U13691 (N_13691,N_6351,N_6116);
or U13692 (N_13692,N_5869,N_6703);
or U13693 (N_13693,N_7114,N_6659);
nor U13694 (N_13694,N_6669,N_7506);
xnor U13695 (N_13695,N_6935,N_5374);
nor U13696 (N_13696,N_7459,N_9022);
xnor U13697 (N_13697,N_5755,N_5594);
nor U13698 (N_13698,N_5085,N_6068);
nor U13699 (N_13699,N_6260,N_8169);
nor U13700 (N_13700,N_9680,N_5272);
and U13701 (N_13701,N_6189,N_7461);
nand U13702 (N_13702,N_5288,N_5826);
xnor U13703 (N_13703,N_7725,N_6358);
xnor U13704 (N_13704,N_9555,N_5076);
or U13705 (N_13705,N_5835,N_7783);
nand U13706 (N_13706,N_5594,N_7702);
nand U13707 (N_13707,N_7555,N_9563);
or U13708 (N_13708,N_7604,N_8728);
xor U13709 (N_13709,N_5887,N_9938);
nor U13710 (N_13710,N_8430,N_5896);
xor U13711 (N_13711,N_7450,N_9336);
xor U13712 (N_13712,N_9141,N_6040);
nor U13713 (N_13713,N_7490,N_9211);
nor U13714 (N_13714,N_7228,N_6842);
nand U13715 (N_13715,N_8618,N_9837);
or U13716 (N_13716,N_5040,N_9651);
xnor U13717 (N_13717,N_8727,N_6783);
xnor U13718 (N_13718,N_5479,N_7735);
nor U13719 (N_13719,N_6547,N_7949);
xnor U13720 (N_13720,N_5271,N_6821);
nor U13721 (N_13721,N_9374,N_9187);
or U13722 (N_13722,N_8362,N_5367);
and U13723 (N_13723,N_7985,N_6362);
and U13724 (N_13724,N_9377,N_8590);
xor U13725 (N_13725,N_8696,N_9926);
nand U13726 (N_13726,N_6217,N_5367);
or U13727 (N_13727,N_6674,N_6923);
xor U13728 (N_13728,N_8704,N_5372);
and U13729 (N_13729,N_7846,N_7009);
nor U13730 (N_13730,N_7289,N_5192);
nand U13731 (N_13731,N_9350,N_8587);
nand U13732 (N_13732,N_7883,N_7291);
xnor U13733 (N_13733,N_6562,N_5472);
or U13734 (N_13734,N_7807,N_5795);
nand U13735 (N_13735,N_8834,N_5414);
or U13736 (N_13736,N_8376,N_9156);
or U13737 (N_13737,N_8203,N_8028);
nand U13738 (N_13738,N_8389,N_9666);
or U13739 (N_13739,N_8846,N_8590);
nand U13740 (N_13740,N_5936,N_5783);
and U13741 (N_13741,N_8609,N_6138);
nor U13742 (N_13742,N_6545,N_9287);
nor U13743 (N_13743,N_8455,N_9096);
nor U13744 (N_13744,N_9830,N_8981);
xnor U13745 (N_13745,N_5864,N_9403);
and U13746 (N_13746,N_9918,N_7292);
nand U13747 (N_13747,N_5226,N_6456);
nand U13748 (N_13748,N_7286,N_7729);
and U13749 (N_13749,N_8845,N_8046);
and U13750 (N_13750,N_5223,N_5239);
or U13751 (N_13751,N_5731,N_6641);
or U13752 (N_13752,N_5809,N_5184);
and U13753 (N_13753,N_8079,N_8133);
and U13754 (N_13754,N_5028,N_8090);
nand U13755 (N_13755,N_9598,N_8366);
nor U13756 (N_13756,N_6928,N_8874);
nor U13757 (N_13757,N_9695,N_6458);
and U13758 (N_13758,N_8589,N_9123);
nor U13759 (N_13759,N_6465,N_6268);
nand U13760 (N_13760,N_5549,N_7829);
and U13761 (N_13761,N_5757,N_8476);
and U13762 (N_13762,N_7523,N_6604);
or U13763 (N_13763,N_8215,N_8220);
nand U13764 (N_13764,N_6152,N_5759);
xnor U13765 (N_13765,N_9413,N_5964);
nor U13766 (N_13766,N_6127,N_8433);
and U13767 (N_13767,N_5621,N_7695);
or U13768 (N_13768,N_5712,N_7269);
nand U13769 (N_13769,N_6460,N_9835);
nor U13770 (N_13770,N_6243,N_6081);
and U13771 (N_13771,N_5759,N_7504);
nor U13772 (N_13772,N_7949,N_7730);
and U13773 (N_13773,N_9206,N_5048);
or U13774 (N_13774,N_5821,N_7703);
or U13775 (N_13775,N_7744,N_8305);
xnor U13776 (N_13776,N_9621,N_9695);
xnor U13777 (N_13777,N_8307,N_7871);
nor U13778 (N_13778,N_9637,N_8331);
nor U13779 (N_13779,N_8233,N_7367);
xor U13780 (N_13780,N_5485,N_6674);
nor U13781 (N_13781,N_8524,N_7813);
or U13782 (N_13782,N_7375,N_5677);
nor U13783 (N_13783,N_8243,N_9984);
nand U13784 (N_13784,N_6540,N_8415);
and U13785 (N_13785,N_7622,N_8121);
nand U13786 (N_13786,N_7505,N_7683);
or U13787 (N_13787,N_6236,N_7423);
xnor U13788 (N_13788,N_6606,N_7605);
nand U13789 (N_13789,N_8556,N_7323);
nor U13790 (N_13790,N_5940,N_5478);
or U13791 (N_13791,N_9183,N_6077);
nand U13792 (N_13792,N_7003,N_5872);
and U13793 (N_13793,N_6613,N_6228);
nand U13794 (N_13794,N_9169,N_5810);
and U13795 (N_13795,N_8401,N_6362);
nand U13796 (N_13796,N_6284,N_8231);
xnor U13797 (N_13797,N_7111,N_5905);
nand U13798 (N_13798,N_9127,N_5733);
or U13799 (N_13799,N_9341,N_6923);
nor U13800 (N_13800,N_8096,N_9805);
nand U13801 (N_13801,N_6167,N_7127);
and U13802 (N_13802,N_7825,N_8802);
nand U13803 (N_13803,N_7862,N_9803);
or U13804 (N_13804,N_6591,N_6596);
nand U13805 (N_13805,N_6179,N_9645);
and U13806 (N_13806,N_6669,N_6868);
xnor U13807 (N_13807,N_8043,N_9953);
xnor U13808 (N_13808,N_6328,N_9501);
xnor U13809 (N_13809,N_7703,N_7066);
or U13810 (N_13810,N_8443,N_9992);
xnor U13811 (N_13811,N_9664,N_6349);
or U13812 (N_13812,N_5788,N_5118);
nor U13813 (N_13813,N_6487,N_7578);
nand U13814 (N_13814,N_7478,N_8117);
nand U13815 (N_13815,N_7626,N_5007);
or U13816 (N_13816,N_7537,N_7461);
xor U13817 (N_13817,N_6036,N_5686);
nand U13818 (N_13818,N_8538,N_6340);
nor U13819 (N_13819,N_8487,N_7173);
nor U13820 (N_13820,N_7341,N_8923);
xor U13821 (N_13821,N_5271,N_7586);
or U13822 (N_13822,N_8404,N_6489);
and U13823 (N_13823,N_5053,N_8422);
or U13824 (N_13824,N_8177,N_7068);
xnor U13825 (N_13825,N_8891,N_9776);
and U13826 (N_13826,N_6841,N_7595);
nand U13827 (N_13827,N_7992,N_7346);
or U13828 (N_13828,N_7520,N_9845);
nor U13829 (N_13829,N_5775,N_9840);
and U13830 (N_13830,N_7631,N_5282);
or U13831 (N_13831,N_9901,N_6041);
nor U13832 (N_13832,N_7564,N_6554);
and U13833 (N_13833,N_8350,N_6333);
nor U13834 (N_13834,N_5449,N_8058);
and U13835 (N_13835,N_8862,N_9864);
xnor U13836 (N_13836,N_8301,N_6340);
nand U13837 (N_13837,N_5418,N_8265);
xor U13838 (N_13838,N_5566,N_9103);
nand U13839 (N_13839,N_6525,N_6800);
nand U13840 (N_13840,N_5342,N_8460);
xor U13841 (N_13841,N_6044,N_9440);
and U13842 (N_13842,N_7489,N_8082);
nand U13843 (N_13843,N_6078,N_7389);
xnor U13844 (N_13844,N_9640,N_9811);
or U13845 (N_13845,N_5220,N_9335);
nor U13846 (N_13846,N_9938,N_6726);
or U13847 (N_13847,N_6587,N_9855);
nor U13848 (N_13848,N_5080,N_6524);
nand U13849 (N_13849,N_8894,N_9649);
nand U13850 (N_13850,N_7924,N_6753);
xnor U13851 (N_13851,N_9600,N_9533);
and U13852 (N_13852,N_9948,N_9036);
nand U13853 (N_13853,N_6075,N_6926);
and U13854 (N_13854,N_9899,N_9595);
nand U13855 (N_13855,N_7341,N_5671);
nand U13856 (N_13856,N_8265,N_6714);
and U13857 (N_13857,N_5472,N_5622);
or U13858 (N_13858,N_9434,N_9572);
or U13859 (N_13859,N_5887,N_8120);
and U13860 (N_13860,N_8453,N_6002);
nor U13861 (N_13861,N_6267,N_8229);
and U13862 (N_13862,N_8337,N_6592);
nand U13863 (N_13863,N_8188,N_9877);
nor U13864 (N_13864,N_8800,N_9483);
xor U13865 (N_13865,N_6099,N_8962);
and U13866 (N_13866,N_9790,N_9437);
nor U13867 (N_13867,N_6715,N_8599);
xnor U13868 (N_13868,N_5570,N_6800);
nand U13869 (N_13869,N_9077,N_6033);
or U13870 (N_13870,N_9437,N_7351);
or U13871 (N_13871,N_5723,N_8100);
nand U13872 (N_13872,N_7901,N_7353);
nand U13873 (N_13873,N_7897,N_8280);
nor U13874 (N_13874,N_6832,N_6413);
nand U13875 (N_13875,N_8321,N_6899);
or U13876 (N_13876,N_9643,N_5350);
and U13877 (N_13877,N_7510,N_7590);
xor U13878 (N_13878,N_9906,N_9614);
nand U13879 (N_13879,N_6955,N_5383);
and U13880 (N_13880,N_5851,N_6742);
nand U13881 (N_13881,N_8668,N_6451);
and U13882 (N_13882,N_8839,N_9316);
xor U13883 (N_13883,N_5962,N_7119);
and U13884 (N_13884,N_9348,N_8560);
and U13885 (N_13885,N_6032,N_8379);
and U13886 (N_13886,N_5267,N_5703);
or U13887 (N_13887,N_5292,N_6896);
nand U13888 (N_13888,N_5562,N_5816);
nor U13889 (N_13889,N_7237,N_9569);
or U13890 (N_13890,N_8738,N_7297);
nor U13891 (N_13891,N_7177,N_5477);
and U13892 (N_13892,N_7310,N_5677);
xnor U13893 (N_13893,N_6517,N_6220);
nor U13894 (N_13894,N_5340,N_7076);
nor U13895 (N_13895,N_7551,N_6853);
or U13896 (N_13896,N_9751,N_6651);
or U13897 (N_13897,N_9961,N_6452);
xor U13898 (N_13898,N_8971,N_6434);
and U13899 (N_13899,N_6317,N_8315);
nor U13900 (N_13900,N_7720,N_7286);
nor U13901 (N_13901,N_9995,N_8097);
or U13902 (N_13902,N_9966,N_5400);
nor U13903 (N_13903,N_7043,N_6082);
and U13904 (N_13904,N_8116,N_9142);
nor U13905 (N_13905,N_7520,N_6525);
nor U13906 (N_13906,N_6533,N_7136);
and U13907 (N_13907,N_8134,N_5024);
or U13908 (N_13908,N_5008,N_7376);
xor U13909 (N_13909,N_5677,N_7306);
and U13910 (N_13910,N_9230,N_9627);
nand U13911 (N_13911,N_7175,N_6537);
nand U13912 (N_13912,N_6076,N_5585);
xor U13913 (N_13913,N_8991,N_5796);
or U13914 (N_13914,N_8708,N_7827);
or U13915 (N_13915,N_6335,N_8651);
or U13916 (N_13916,N_7888,N_6508);
xor U13917 (N_13917,N_9793,N_7671);
or U13918 (N_13918,N_5519,N_9700);
nand U13919 (N_13919,N_6400,N_6216);
nand U13920 (N_13920,N_5250,N_9425);
nand U13921 (N_13921,N_8669,N_5986);
nor U13922 (N_13922,N_7404,N_8552);
nor U13923 (N_13923,N_5598,N_5118);
and U13924 (N_13924,N_5449,N_5155);
nand U13925 (N_13925,N_9660,N_5558);
nand U13926 (N_13926,N_9904,N_5386);
and U13927 (N_13927,N_8410,N_7753);
xnor U13928 (N_13928,N_7224,N_9564);
and U13929 (N_13929,N_9125,N_8274);
and U13930 (N_13930,N_7184,N_7630);
nor U13931 (N_13931,N_9268,N_7669);
or U13932 (N_13932,N_6184,N_7034);
or U13933 (N_13933,N_8105,N_5543);
nor U13934 (N_13934,N_7938,N_7090);
or U13935 (N_13935,N_9330,N_9986);
xnor U13936 (N_13936,N_7404,N_9204);
nand U13937 (N_13937,N_9714,N_6418);
and U13938 (N_13938,N_9738,N_5011);
nor U13939 (N_13939,N_9303,N_6637);
nor U13940 (N_13940,N_6344,N_7994);
nand U13941 (N_13941,N_9788,N_6244);
nor U13942 (N_13942,N_7371,N_9854);
xnor U13943 (N_13943,N_7707,N_6544);
xor U13944 (N_13944,N_5414,N_7748);
and U13945 (N_13945,N_7907,N_6200);
nand U13946 (N_13946,N_8803,N_8613);
and U13947 (N_13947,N_7786,N_6859);
or U13948 (N_13948,N_8642,N_7517);
nor U13949 (N_13949,N_8022,N_8760);
or U13950 (N_13950,N_9568,N_5556);
or U13951 (N_13951,N_9195,N_7184);
nand U13952 (N_13952,N_7889,N_5941);
or U13953 (N_13953,N_5683,N_5294);
and U13954 (N_13954,N_5202,N_6585);
and U13955 (N_13955,N_7633,N_6363);
nand U13956 (N_13956,N_7523,N_9628);
nand U13957 (N_13957,N_8010,N_7439);
and U13958 (N_13958,N_9893,N_6758);
nand U13959 (N_13959,N_7983,N_8026);
and U13960 (N_13960,N_7369,N_6670);
nand U13961 (N_13961,N_5324,N_9991);
or U13962 (N_13962,N_5163,N_8841);
or U13963 (N_13963,N_9294,N_9603);
xor U13964 (N_13964,N_8420,N_6127);
nor U13965 (N_13965,N_6112,N_8001);
and U13966 (N_13966,N_8502,N_5068);
and U13967 (N_13967,N_7101,N_7761);
xor U13968 (N_13968,N_5143,N_9312);
nand U13969 (N_13969,N_5622,N_7227);
or U13970 (N_13970,N_9443,N_5156);
nand U13971 (N_13971,N_6126,N_5084);
xor U13972 (N_13972,N_6340,N_7503);
nor U13973 (N_13973,N_9591,N_5968);
nor U13974 (N_13974,N_9807,N_9320);
and U13975 (N_13975,N_7170,N_7158);
nor U13976 (N_13976,N_9462,N_6003);
nor U13977 (N_13977,N_8454,N_9236);
nand U13978 (N_13978,N_9184,N_5090);
xnor U13979 (N_13979,N_5709,N_5086);
and U13980 (N_13980,N_9877,N_5321);
xnor U13981 (N_13981,N_8049,N_7478);
and U13982 (N_13982,N_9265,N_6599);
or U13983 (N_13983,N_5717,N_7994);
and U13984 (N_13984,N_7199,N_6846);
or U13985 (N_13985,N_8070,N_8086);
nor U13986 (N_13986,N_6439,N_6517);
or U13987 (N_13987,N_9029,N_6809);
nor U13988 (N_13988,N_5344,N_9839);
xor U13989 (N_13989,N_5006,N_5988);
nand U13990 (N_13990,N_6565,N_7330);
or U13991 (N_13991,N_9192,N_9061);
nand U13992 (N_13992,N_8815,N_8124);
and U13993 (N_13993,N_9821,N_5616);
and U13994 (N_13994,N_9887,N_5792);
or U13995 (N_13995,N_9280,N_8362);
and U13996 (N_13996,N_8328,N_6901);
xor U13997 (N_13997,N_8144,N_6336);
nor U13998 (N_13998,N_9608,N_5240);
nand U13999 (N_13999,N_6829,N_5790);
or U14000 (N_14000,N_9714,N_7250);
xor U14001 (N_14001,N_8864,N_5055);
nand U14002 (N_14002,N_8506,N_5966);
and U14003 (N_14003,N_7862,N_5698);
and U14004 (N_14004,N_7663,N_5031);
and U14005 (N_14005,N_5083,N_7881);
nand U14006 (N_14006,N_7050,N_6391);
nor U14007 (N_14007,N_6844,N_9407);
and U14008 (N_14008,N_7170,N_9335);
and U14009 (N_14009,N_5407,N_9306);
and U14010 (N_14010,N_5369,N_8101);
xor U14011 (N_14011,N_5468,N_6942);
nor U14012 (N_14012,N_7574,N_8567);
xor U14013 (N_14013,N_7722,N_8410);
and U14014 (N_14014,N_7698,N_7573);
nand U14015 (N_14015,N_7590,N_8031);
and U14016 (N_14016,N_7005,N_5872);
nor U14017 (N_14017,N_9812,N_6054);
xnor U14018 (N_14018,N_9413,N_8679);
nand U14019 (N_14019,N_5780,N_8557);
or U14020 (N_14020,N_6607,N_7384);
nand U14021 (N_14021,N_7344,N_5073);
nor U14022 (N_14022,N_8448,N_6763);
xor U14023 (N_14023,N_9058,N_6922);
xnor U14024 (N_14024,N_6692,N_9788);
nand U14025 (N_14025,N_9330,N_5468);
and U14026 (N_14026,N_7497,N_6635);
and U14027 (N_14027,N_7278,N_5083);
nand U14028 (N_14028,N_8512,N_5929);
nor U14029 (N_14029,N_6704,N_6833);
nand U14030 (N_14030,N_6018,N_6597);
nor U14031 (N_14031,N_5512,N_9709);
xor U14032 (N_14032,N_7084,N_9634);
xor U14033 (N_14033,N_5363,N_7226);
xnor U14034 (N_14034,N_7206,N_6431);
and U14035 (N_14035,N_8833,N_6059);
nor U14036 (N_14036,N_7269,N_7660);
xor U14037 (N_14037,N_7656,N_5392);
and U14038 (N_14038,N_9864,N_7292);
or U14039 (N_14039,N_9019,N_6131);
or U14040 (N_14040,N_6697,N_8539);
or U14041 (N_14041,N_7730,N_5159);
and U14042 (N_14042,N_9581,N_5564);
and U14043 (N_14043,N_7191,N_5452);
nor U14044 (N_14044,N_5300,N_7412);
or U14045 (N_14045,N_8182,N_7112);
and U14046 (N_14046,N_6847,N_9571);
nor U14047 (N_14047,N_8762,N_9688);
and U14048 (N_14048,N_5620,N_8992);
or U14049 (N_14049,N_9125,N_7595);
and U14050 (N_14050,N_8871,N_9995);
xnor U14051 (N_14051,N_9461,N_6590);
xor U14052 (N_14052,N_6847,N_9530);
or U14053 (N_14053,N_8130,N_6487);
xnor U14054 (N_14054,N_5857,N_7221);
nor U14055 (N_14055,N_5743,N_9362);
xor U14056 (N_14056,N_7138,N_6206);
or U14057 (N_14057,N_7565,N_8654);
nor U14058 (N_14058,N_8564,N_8541);
or U14059 (N_14059,N_8440,N_6257);
xnor U14060 (N_14060,N_5230,N_8357);
and U14061 (N_14061,N_8545,N_6751);
xnor U14062 (N_14062,N_5131,N_7619);
or U14063 (N_14063,N_6737,N_8162);
nand U14064 (N_14064,N_5246,N_5266);
or U14065 (N_14065,N_9430,N_7471);
nand U14066 (N_14066,N_7340,N_9183);
or U14067 (N_14067,N_6162,N_6681);
or U14068 (N_14068,N_6427,N_9444);
xor U14069 (N_14069,N_8881,N_8802);
xnor U14070 (N_14070,N_8518,N_7737);
nand U14071 (N_14071,N_5712,N_7676);
xnor U14072 (N_14072,N_6833,N_8740);
and U14073 (N_14073,N_8803,N_5765);
or U14074 (N_14074,N_6517,N_8121);
or U14075 (N_14075,N_5801,N_7480);
or U14076 (N_14076,N_6839,N_6441);
or U14077 (N_14077,N_6666,N_9751);
or U14078 (N_14078,N_7161,N_7762);
xnor U14079 (N_14079,N_7880,N_7352);
xnor U14080 (N_14080,N_7120,N_9295);
nand U14081 (N_14081,N_7030,N_6529);
and U14082 (N_14082,N_5503,N_9270);
xnor U14083 (N_14083,N_9204,N_6553);
xnor U14084 (N_14084,N_9098,N_9137);
nand U14085 (N_14085,N_7622,N_9188);
or U14086 (N_14086,N_8600,N_7977);
or U14087 (N_14087,N_6257,N_9239);
nor U14088 (N_14088,N_9412,N_7537);
and U14089 (N_14089,N_5453,N_9380);
xor U14090 (N_14090,N_7459,N_6311);
nand U14091 (N_14091,N_9005,N_6071);
or U14092 (N_14092,N_7829,N_6427);
nor U14093 (N_14093,N_8148,N_9568);
or U14094 (N_14094,N_9785,N_7742);
and U14095 (N_14095,N_5258,N_8909);
nor U14096 (N_14096,N_5996,N_9791);
and U14097 (N_14097,N_5996,N_5240);
xnor U14098 (N_14098,N_8116,N_8856);
or U14099 (N_14099,N_8676,N_6280);
and U14100 (N_14100,N_5890,N_9505);
and U14101 (N_14101,N_6975,N_6858);
nand U14102 (N_14102,N_9887,N_9708);
or U14103 (N_14103,N_9999,N_9770);
nor U14104 (N_14104,N_5952,N_7990);
and U14105 (N_14105,N_9173,N_8342);
or U14106 (N_14106,N_8662,N_7135);
or U14107 (N_14107,N_5137,N_8358);
or U14108 (N_14108,N_6015,N_6107);
and U14109 (N_14109,N_9174,N_5016);
or U14110 (N_14110,N_6512,N_7451);
nor U14111 (N_14111,N_8426,N_6840);
nand U14112 (N_14112,N_9474,N_7055);
nor U14113 (N_14113,N_6856,N_6907);
and U14114 (N_14114,N_9636,N_8332);
xnor U14115 (N_14115,N_7959,N_6800);
or U14116 (N_14116,N_7739,N_9540);
nor U14117 (N_14117,N_5709,N_8135);
xor U14118 (N_14118,N_9493,N_6907);
nor U14119 (N_14119,N_7666,N_6173);
and U14120 (N_14120,N_9357,N_8501);
nor U14121 (N_14121,N_8287,N_5687);
xnor U14122 (N_14122,N_7028,N_5172);
and U14123 (N_14123,N_9367,N_8730);
xor U14124 (N_14124,N_6118,N_7095);
xnor U14125 (N_14125,N_5717,N_9170);
nor U14126 (N_14126,N_7502,N_6086);
xnor U14127 (N_14127,N_7360,N_5496);
or U14128 (N_14128,N_5474,N_6099);
and U14129 (N_14129,N_8812,N_8567);
nor U14130 (N_14130,N_6893,N_8082);
nand U14131 (N_14131,N_7481,N_9039);
or U14132 (N_14132,N_6837,N_9537);
or U14133 (N_14133,N_9921,N_6167);
and U14134 (N_14134,N_5226,N_9272);
and U14135 (N_14135,N_7528,N_7703);
or U14136 (N_14136,N_6690,N_8013);
xor U14137 (N_14137,N_5439,N_5880);
and U14138 (N_14138,N_7767,N_7723);
nand U14139 (N_14139,N_9111,N_9022);
and U14140 (N_14140,N_7762,N_6891);
nor U14141 (N_14141,N_8100,N_7116);
nand U14142 (N_14142,N_7232,N_9088);
and U14143 (N_14143,N_7916,N_8656);
or U14144 (N_14144,N_7926,N_7505);
nand U14145 (N_14145,N_8951,N_5385);
and U14146 (N_14146,N_5700,N_7244);
nand U14147 (N_14147,N_5758,N_7251);
and U14148 (N_14148,N_6576,N_8533);
or U14149 (N_14149,N_7261,N_6579);
nand U14150 (N_14150,N_8342,N_9149);
and U14151 (N_14151,N_8207,N_8320);
xnor U14152 (N_14152,N_6386,N_6565);
nor U14153 (N_14153,N_5514,N_7582);
and U14154 (N_14154,N_8117,N_9940);
nor U14155 (N_14155,N_7084,N_8478);
and U14156 (N_14156,N_6869,N_9750);
nand U14157 (N_14157,N_5204,N_8097);
and U14158 (N_14158,N_7180,N_5226);
and U14159 (N_14159,N_9959,N_7763);
nand U14160 (N_14160,N_8094,N_9237);
nand U14161 (N_14161,N_5869,N_8303);
nor U14162 (N_14162,N_6726,N_8341);
nand U14163 (N_14163,N_6852,N_6137);
nand U14164 (N_14164,N_8206,N_6385);
nor U14165 (N_14165,N_8384,N_8616);
or U14166 (N_14166,N_9885,N_5933);
nand U14167 (N_14167,N_7910,N_9680);
and U14168 (N_14168,N_7138,N_5999);
and U14169 (N_14169,N_9969,N_9724);
nand U14170 (N_14170,N_6479,N_7917);
or U14171 (N_14171,N_6570,N_9148);
or U14172 (N_14172,N_5652,N_5851);
nor U14173 (N_14173,N_9084,N_8356);
or U14174 (N_14174,N_5229,N_6124);
or U14175 (N_14175,N_9551,N_7702);
xnor U14176 (N_14176,N_5556,N_9723);
nand U14177 (N_14177,N_6623,N_8602);
nor U14178 (N_14178,N_6913,N_9164);
or U14179 (N_14179,N_7578,N_5392);
nand U14180 (N_14180,N_7348,N_7833);
nand U14181 (N_14181,N_6338,N_9457);
nand U14182 (N_14182,N_5023,N_8195);
or U14183 (N_14183,N_9359,N_8238);
nand U14184 (N_14184,N_8217,N_8079);
nor U14185 (N_14185,N_8577,N_5210);
xnor U14186 (N_14186,N_9842,N_7973);
and U14187 (N_14187,N_5722,N_5913);
or U14188 (N_14188,N_5079,N_6984);
and U14189 (N_14189,N_7384,N_8017);
xnor U14190 (N_14190,N_8745,N_5309);
and U14191 (N_14191,N_8787,N_9211);
nor U14192 (N_14192,N_5349,N_7319);
nand U14193 (N_14193,N_9576,N_9104);
nor U14194 (N_14194,N_8152,N_5825);
xnor U14195 (N_14195,N_8995,N_5821);
xor U14196 (N_14196,N_9318,N_9923);
nor U14197 (N_14197,N_8712,N_9958);
nor U14198 (N_14198,N_8095,N_5274);
nand U14199 (N_14199,N_9202,N_5861);
xnor U14200 (N_14200,N_8694,N_8229);
xnor U14201 (N_14201,N_6744,N_5950);
nor U14202 (N_14202,N_7766,N_7477);
nor U14203 (N_14203,N_6129,N_7021);
and U14204 (N_14204,N_6327,N_6013);
xnor U14205 (N_14205,N_8167,N_9195);
nand U14206 (N_14206,N_7916,N_5939);
or U14207 (N_14207,N_9051,N_5178);
and U14208 (N_14208,N_7647,N_6912);
xor U14209 (N_14209,N_7729,N_5201);
nand U14210 (N_14210,N_9533,N_5345);
nand U14211 (N_14211,N_6431,N_7759);
xor U14212 (N_14212,N_8344,N_9233);
xor U14213 (N_14213,N_7093,N_9905);
or U14214 (N_14214,N_6047,N_5446);
xor U14215 (N_14215,N_9857,N_6103);
xor U14216 (N_14216,N_7816,N_7871);
and U14217 (N_14217,N_7727,N_5915);
xor U14218 (N_14218,N_9843,N_9958);
nand U14219 (N_14219,N_7778,N_6556);
and U14220 (N_14220,N_7609,N_5889);
or U14221 (N_14221,N_6251,N_5213);
xor U14222 (N_14222,N_6082,N_6756);
xnor U14223 (N_14223,N_9002,N_8028);
and U14224 (N_14224,N_5683,N_8461);
nor U14225 (N_14225,N_9413,N_8213);
and U14226 (N_14226,N_9628,N_8420);
xor U14227 (N_14227,N_9079,N_5085);
and U14228 (N_14228,N_6037,N_7169);
nand U14229 (N_14229,N_6941,N_8942);
and U14230 (N_14230,N_8093,N_6989);
nand U14231 (N_14231,N_7651,N_8273);
nor U14232 (N_14232,N_7368,N_6568);
and U14233 (N_14233,N_6193,N_5941);
nor U14234 (N_14234,N_6091,N_5018);
xor U14235 (N_14235,N_9174,N_7935);
nand U14236 (N_14236,N_8314,N_6756);
xor U14237 (N_14237,N_7705,N_7139);
nor U14238 (N_14238,N_5486,N_9407);
nand U14239 (N_14239,N_8027,N_5603);
nand U14240 (N_14240,N_5313,N_7755);
and U14241 (N_14241,N_5510,N_9348);
and U14242 (N_14242,N_7930,N_7862);
nand U14243 (N_14243,N_9662,N_6786);
xor U14244 (N_14244,N_6055,N_5879);
nand U14245 (N_14245,N_5880,N_9836);
nand U14246 (N_14246,N_7418,N_9786);
nor U14247 (N_14247,N_9532,N_7693);
xor U14248 (N_14248,N_8335,N_7748);
nand U14249 (N_14249,N_7941,N_7563);
nor U14250 (N_14250,N_6181,N_7899);
xor U14251 (N_14251,N_8223,N_6268);
or U14252 (N_14252,N_7113,N_8817);
nor U14253 (N_14253,N_7602,N_7545);
nor U14254 (N_14254,N_6675,N_6238);
nor U14255 (N_14255,N_6731,N_6972);
and U14256 (N_14256,N_7705,N_9326);
xnor U14257 (N_14257,N_6598,N_9551);
nor U14258 (N_14258,N_6329,N_5206);
nor U14259 (N_14259,N_5248,N_7114);
nor U14260 (N_14260,N_8822,N_9936);
xnor U14261 (N_14261,N_8669,N_7152);
nor U14262 (N_14262,N_7980,N_8845);
nor U14263 (N_14263,N_5258,N_7859);
nor U14264 (N_14264,N_5216,N_6392);
nor U14265 (N_14265,N_9683,N_7688);
nor U14266 (N_14266,N_5435,N_8680);
nand U14267 (N_14267,N_7296,N_5493);
or U14268 (N_14268,N_8103,N_9448);
or U14269 (N_14269,N_5146,N_6736);
nand U14270 (N_14270,N_8364,N_7481);
nor U14271 (N_14271,N_7627,N_9785);
nor U14272 (N_14272,N_8644,N_8474);
or U14273 (N_14273,N_5513,N_8388);
xor U14274 (N_14274,N_5189,N_9275);
or U14275 (N_14275,N_5841,N_5562);
xnor U14276 (N_14276,N_8583,N_7960);
nor U14277 (N_14277,N_6222,N_7936);
nor U14278 (N_14278,N_8861,N_8482);
nand U14279 (N_14279,N_8151,N_5728);
or U14280 (N_14280,N_5271,N_6621);
or U14281 (N_14281,N_6677,N_7036);
and U14282 (N_14282,N_9200,N_6718);
and U14283 (N_14283,N_8450,N_7352);
or U14284 (N_14284,N_9690,N_9048);
and U14285 (N_14285,N_9240,N_5985);
and U14286 (N_14286,N_5459,N_7295);
and U14287 (N_14287,N_7378,N_9591);
or U14288 (N_14288,N_5524,N_9659);
xor U14289 (N_14289,N_5750,N_7675);
or U14290 (N_14290,N_8118,N_9161);
or U14291 (N_14291,N_7993,N_5267);
xor U14292 (N_14292,N_9319,N_7066);
or U14293 (N_14293,N_9953,N_7525);
or U14294 (N_14294,N_9072,N_7156);
nor U14295 (N_14295,N_6717,N_6198);
and U14296 (N_14296,N_5318,N_5311);
nand U14297 (N_14297,N_6823,N_6363);
nor U14298 (N_14298,N_5539,N_6830);
nand U14299 (N_14299,N_7054,N_5823);
nand U14300 (N_14300,N_8330,N_6632);
nand U14301 (N_14301,N_5691,N_9842);
and U14302 (N_14302,N_5988,N_8459);
xor U14303 (N_14303,N_5108,N_9678);
xor U14304 (N_14304,N_7652,N_6865);
or U14305 (N_14305,N_5837,N_9253);
or U14306 (N_14306,N_5980,N_6709);
xor U14307 (N_14307,N_5584,N_7674);
or U14308 (N_14308,N_5126,N_8949);
or U14309 (N_14309,N_9629,N_9304);
or U14310 (N_14310,N_5461,N_7750);
nor U14311 (N_14311,N_9003,N_6991);
nand U14312 (N_14312,N_9365,N_5534);
nor U14313 (N_14313,N_5960,N_6997);
or U14314 (N_14314,N_8799,N_5883);
or U14315 (N_14315,N_9355,N_8902);
xnor U14316 (N_14316,N_8031,N_8349);
nand U14317 (N_14317,N_8608,N_7730);
nand U14318 (N_14318,N_6662,N_5676);
xor U14319 (N_14319,N_6632,N_9089);
or U14320 (N_14320,N_5643,N_7710);
nand U14321 (N_14321,N_6256,N_5239);
nor U14322 (N_14322,N_9447,N_7870);
and U14323 (N_14323,N_7161,N_5927);
nand U14324 (N_14324,N_6374,N_9524);
nand U14325 (N_14325,N_8899,N_9485);
nand U14326 (N_14326,N_5980,N_5135);
nor U14327 (N_14327,N_5784,N_7165);
nor U14328 (N_14328,N_7055,N_5444);
nor U14329 (N_14329,N_9904,N_7374);
xnor U14330 (N_14330,N_7454,N_6108);
nor U14331 (N_14331,N_8854,N_7764);
xor U14332 (N_14332,N_6807,N_9959);
nand U14333 (N_14333,N_5781,N_5769);
nand U14334 (N_14334,N_8438,N_7710);
nand U14335 (N_14335,N_6695,N_7220);
nor U14336 (N_14336,N_7684,N_7676);
or U14337 (N_14337,N_5867,N_7192);
nand U14338 (N_14338,N_7325,N_6609);
nand U14339 (N_14339,N_5920,N_9774);
nor U14340 (N_14340,N_7701,N_7688);
nand U14341 (N_14341,N_8972,N_6855);
and U14342 (N_14342,N_8146,N_7350);
nor U14343 (N_14343,N_9686,N_8210);
xnor U14344 (N_14344,N_5883,N_9500);
and U14345 (N_14345,N_9424,N_6590);
nand U14346 (N_14346,N_8027,N_6873);
nor U14347 (N_14347,N_5090,N_9434);
nor U14348 (N_14348,N_6189,N_8706);
and U14349 (N_14349,N_7240,N_7360);
and U14350 (N_14350,N_9630,N_6448);
or U14351 (N_14351,N_5001,N_7691);
and U14352 (N_14352,N_8280,N_5117);
or U14353 (N_14353,N_8190,N_5227);
nor U14354 (N_14354,N_9256,N_5404);
nor U14355 (N_14355,N_7941,N_5766);
xnor U14356 (N_14356,N_8656,N_5474);
and U14357 (N_14357,N_8222,N_8376);
nand U14358 (N_14358,N_6316,N_8530);
nand U14359 (N_14359,N_7835,N_5957);
nor U14360 (N_14360,N_5070,N_6822);
or U14361 (N_14361,N_8594,N_9699);
and U14362 (N_14362,N_5610,N_5912);
or U14363 (N_14363,N_8454,N_7892);
and U14364 (N_14364,N_8543,N_9731);
nor U14365 (N_14365,N_8562,N_9442);
nor U14366 (N_14366,N_7997,N_9985);
or U14367 (N_14367,N_5516,N_7498);
nor U14368 (N_14368,N_7007,N_9758);
xnor U14369 (N_14369,N_5164,N_5430);
xor U14370 (N_14370,N_8543,N_5514);
nor U14371 (N_14371,N_8647,N_6957);
nor U14372 (N_14372,N_8231,N_7400);
xnor U14373 (N_14373,N_8392,N_6659);
nor U14374 (N_14374,N_9614,N_8005);
xor U14375 (N_14375,N_7308,N_6555);
or U14376 (N_14376,N_5649,N_5004);
and U14377 (N_14377,N_7839,N_8306);
xor U14378 (N_14378,N_8140,N_7010);
and U14379 (N_14379,N_6242,N_9068);
nand U14380 (N_14380,N_5626,N_5660);
nand U14381 (N_14381,N_7824,N_7214);
and U14382 (N_14382,N_7251,N_5784);
xnor U14383 (N_14383,N_7158,N_9851);
nand U14384 (N_14384,N_5208,N_9266);
or U14385 (N_14385,N_6553,N_5132);
or U14386 (N_14386,N_6452,N_6188);
nand U14387 (N_14387,N_5112,N_7935);
nor U14388 (N_14388,N_6388,N_9882);
and U14389 (N_14389,N_9703,N_6665);
nor U14390 (N_14390,N_5428,N_7116);
nand U14391 (N_14391,N_6725,N_7827);
xnor U14392 (N_14392,N_5149,N_8520);
or U14393 (N_14393,N_5649,N_7828);
and U14394 (N_14394,N_5785,N_6775);
nor U14395 (N_14395,N_5382,N_8058);
or U14396 (N_14396,N_5872,N_6862);
nand U14397 (N_14397,N_8424,N_8473);
or U14398 (N_14398,N_5203,N_8266);
xor U14399 (N_14399,N_8293,N_5939);
nand U14400 (N_14400,N_7740,N_7354);
nand U14401 (N_14401,N_5028,N_8079);
nand U14402 (N_14402,N_8300,N_9540);
nor U14403 (N_14403,N_7967,N_9031);
and U14404 (N_14404,N_5810,N_6568);
nor U14405 (N_14405,N_6831,N_9380);
nor U14406 (N_14406,N_8048,N_7778);
nand U14407 (N_14407,N_6297,N_5838);
or U14408 (N_14408,N_8513,N_5937);
nand U14409 (N_14409,N_9925,N_9633);
xor U14410 (N_14410,N_6391,N_8032);
or U14411 (N_14411,N_7978,N_9874);
and U14412 (N_14412,N_9626,N_7866);
or U14413 (N_14413,N_7230,N_5366);
or U14414 (N_14414,N_8670,N_5538);
xnor U14415 (N_14415,N_7589,N_9474);
and U14416 (N_14416,N_7598,N_9431);
or U14417 (N_14417,N_8723,N_6840);
and U14418 (N_14418,N_6813,N_7669);
xnor U14419 (N_14419,N_8949,N_5545);
nand U14420 (N_14420,N_5424,N_8608);
nand U14421 (N_14421,N_6118,N_5970);
and U14422 (N_14422,N_9715,N_8369);
or U14423 (N_14423,N_7363,N_6065);
or U14424 (N_14424,N_5135,N_9306);
nor U14425 (N_14425,N_7691,N_7564);
nor U14426 (N_14426,N_5235,N_5492);
nand U14427 (N_14427,N_6198,N_7009);
nand U14428 (N_14428,N_5402,N_6052);
or U14429 (N_14429,N_7642,N_7480);
xor U14430 (N_14430,N_6816,N_5107);
or U14431 (N_14431,N_9753,N_6481);
or U14432 (N_14432,N_8246,N_7980);
xor U14433 (N_14433,N_6780,N_8474);
nor U14434 (N_14434,N_6606,N_5324);
nor U14435 (N_14435,N_5790,N_8189);
or U14436 (N_14436,N_8739,N_5747);
or U14437 (N_14437,N_5435,N_9905);
or U14438 (N_14438,N_5050,N_9624);
xnor U14439 (N_14439,N_8072,N_6836);
and U14440 (N_14440,N_9843,N_9182);
xnor U14441 (N_14441,N_9063,N_7065);
xor U14442 (N_14442,N_5411,N_5996);
or U14443 (N_14443,N_5865,N_7115);
or U14444 (N_14444,N_6451,N_5950);
or U14445 (N_14445,N_9981,N_5661);
nor U14446 (N_14446,N_5475,N_8779);
nor U14447 (N_14447,N_5597,N_5421);
or U14448 (N_14448,N_5434,N_9780);
nor U14449 (N_14449,N_5288,N_7219);
or U14450 (N_14450,N_6741,N_9275);
and U14451 (N_14451,N_5844,N_7486);
or U14452 (N_14452,N_5872,N_8760);
and U14453 (N_14453,N_5480,N_8291);
nand U14454 (N_14454,N_9134,N_5660);
and U14455 (N_14455,N_5877,N_8558);
and U14456 (N_14456,N_8142,N_8016);
nand U14457 (N_14457,N_9136,N_5744);
nor U14458 (N_14458,N_8305,N_6140);
xnor U14459 (N_14459,N_8948,N_5199);
nand U14460 (N_14460,N_9023,N_9439);
nand U14461 (N_14461,N_8348,N_9788);
nor U14462 (N_14462,N_8969,N_9289);
nand U14463 (N_14463,N_7881,N_5162);
nand U14464 (N_14464,N_7656,N_6214);
nor U14465 (N_14465,N_6275,N_5615);
xnor U14466 (N_14466,N_7998,N_7285);
xnor U14467 (N_14467,N_5863,N_6530);
nand U14468 (N_14468,N_7627,N_5671);
nand U14469 (N_14469,N_7691,N_8788);
nor U14470 (N_14470,N_8601,N_7618);
nand U14471 (N_14471,N_9807,N_8794);
and U14472 (N_14472,N_8342,N_8199);
or U14473 (N_14473,N_6640,N_7481);
xor U14474 (N_14474,N_8791,N_6041);
nand U14475 (N_14475,N_9062,N_9822);
nor U14476 (N_14476,N_9105,N_8587);
or U14477 (N_14477,N_7564,N_5532);
and U14478 (N_14478,N_7886,N_8597);
or U14479 (N_14479,N_8215,N_7664);
xnor U14480 (N_14480,N_8062,N_5374);
or U14481 (N_14481,N_7338,N_6531);
or U14482 (N_14482,N_5359,N_9614);
and U14483 (N_14483,N_8296,N_8733);
nand U14484 (N_14484,N_8632,N_7105);
and U14485 (N_14485,N_9214,N_6999);
nand U14486 (N_14486,N_5033,N_7708);
xnor U14487 (N_14487,N_6407,N_9216);
and U14488 (N_14488,N_6153,N_5313);
or U14489 (N_14489,N_9223,N_8335);
nand U14490 (N_14490,N_7810,N_9796);
xnor U14491 (N_14491,N_6440,N_9211);
nor U14492 (N_14492,N_6478,N_5804);
nor U14493 (N_14493,N_8813,N_9742);
nor U14494 (N_14494,N_9937,N_8061);
or U14495 (N_14495,N_7452,N_8639);
or U14496 (N_14496,N_6504,N_9608);
xor U14497 (N_14497,N_7576,N_9306);
nor U14498 (N_14498,N_6261,N_6704);
nor U14499 (N_14499,N_5121,N_9153);
nor U14500 (N_14500,N_6166,N_5556);
nor U14501 (N_14501,N_5122,N_8425);
nand U14502 (N_14502,N_8380,N_7196);
or U14503 (N_14503,N_5996,N_7880);
nor U14504 (N_14504,N_5905,N_6245);
and U14505 (N_14505,N_5009,N_9352);
or U14506 (N_14506,N_7322,N_7635);
xor U14507 (N_14507,N_8959,N_6350);
and U14508 (N_14508,N_5784,N_9095);
nand U14509 (N_14509,N_9347,N_7627);
nand U14510 (N_14510,N_6035,N_9788);
and U14511 (N_14511,N_9092,N_6715);
xnor U14512 (N_14512,N_9104,N_5243);
xor U14513 (N_14513,N_5025,N_7823);
xnor U14514 (N_14514,N_8845,N_7005);
nand U14515 (N_14515,N_5141,N_9730);
and U14516 (N_14516,N_5503,N_5341);
nor U14517 (N_14517,N_5241,N_7607);
nor U14518 (N_14518,N_7428,N_6602);
nor U14519 (N_14519,N_5849,N_7842);
nand U14520 (N_14520,N_8420,N_7058);
or U14521 (N_14521,N_8127,N_6120);
nand U14522 (N_14522,N_7885,N_7488);
or U14523 (N_14523,N_5643,N_9922);
and U14524 (N_14524,N_9312,N_9356);
nand U14525 (N_14525,N_8513,N_9986);
xor U14526 (N_14526,N_8355,N_8513);
and U14527 (N_14527,N_8723,N_8611);
nor U14528 (N_14528,N_9238,N_9863);
nand U14529 (N_14529,N_9484,N_7259);
and U14530 (N_14530,N_6470,N_9448);
xnor U14531 (N_14531,N_5869,N_8731);
xnor U14532 (N_14532,N_9085,N_6181);
and U14533 (N_14533,N_8684,N_9113);
or U14534 (N_14534,N_9128,N_7288);
xor U14535 (N_14535,N_6756,N_6112);
nor U14536 (N_14536,N_8687,N_6897);
and U14537 (N_14537,N_9323,N_7224);
or U14538 (N_14538,N_6899,N_6842);
nand U14539 (N_14539,N_7848,N_8313);
nor U14540 (N_14540,N_6316,N_9176);
xor U14541 (N_14541,N_7400,N_5071);
and U14542 (N_14542,N_6847,N_7726);
nand U14543 (N_14543,N_5312,N_6961);
nand U14544 (N_14544,N_6046,N_5573);
nor U14545 (N_14545,N_8375,N_9912);
nand U14546 (N_14546,N_7125,N_7574);
and U14547 (N_14547,N_6895,N_7126);
nor U14548 (N_14548,N_6243,N_7465);
or U14549 (N_14549,N_9898,N_6124);
nor U14550 (N_14550,N_9528,N_9211);
nand U14551 (N_14551,N_8805,N_9351);
nor U14552 (N_14552,N_9228,N_5527);
nand U14553 (N_14553,N_5033,N_7808);
and U14554 (N_14554,N_6605,N_7546);
or U14555 (N_14555,N_9477,N_7446);
nor U14556 (N_14556,N_8408,N_5893);
nand U14557 (N_14557,N_6969,N_9893);
xnor U14558 (N_14558,N_6792,N_6691);
xor U14559 (N_14559,N_6940,N_8879);
nor U14560 (N_14560,N_7288,N_8935);
nand U14561 (N_14561,N_8481,N_9842);
nand U14562 (N_14562,N_7342,N_6173);
and U14563 (N_14563,N_9427,N_7179);
or U14564 (N_14564,N_6444,N_6691);
or U14565 (N_14565,N_6567,N_9795);
or U14566 (N_14566,N_8397,N_9661);
nor U14567 (N_14567,N_5650,N_6470);
and U14568 (N_14568,N_9601,N_9345);
and U14569 (N_14569,N_8302,N_5762);
nand U14570 (N_14570,N_6212,N_8879);
nor U14571 (N_14571,N_7025,N_5881);
xor U14572 (N_14572,N_8316,N_7177);
nand U14573 (N_14573,N_6829,N_9732);
xnor U14574 (N_14574,N_9952,N_8759);
and U14575 (N_14575,N_8678,N_5820);
or U14576 (N_14576,N_8501,N_7635);
or U14577 (N_14577,N_5764,N_8824);
xor U14578 (N_14578,N_7885,N_7013);
or U14579 (N_14579,N_7643,N_5885);
and U14580 (N_14580,N_6154,N_8034);
nor U14581 (N_14581,N_5798,N_6381);
and U14582 (N_14582,N_9456,N_9761);
xnor U14583 (N_14583,N_8994,N_9232);
or U14584 (N_14584,N_6009,N_6667);
nand U14585 (N_14585,N_8951,N_8806);
nor U14586 (N_14586,N_5414,N_5065);
nor U14587 (N_14587,N_8219,N_9240);
nand U14588 (N_14588,N_8285,N_6097);
xor U14589 (N_14589,N_8665,N_9661);
nand U14590 (N_14590,N_9872,N_7780);
or U14591 (N_14591,N_9783,N_9688);
nand U14592 (N_14592,N_8145,N_7833);
and U14593 (N_14593,N_5762,N_6971);
xor U14594 (N_14594,N_7943,N_6595);
or U14595 (N_14595,N_8352,N_7116);
and U14596 (N_14596,N_7477,N_8197);
nand U14597 (N_14597,N_9230,N_9701);
nor U14598 (N_14598,N_7505,N_8233);
xnor U14599 (N_14599,N_7106,N_6163);
nand U14600 (N_14600,N_8596,N_7403);
nor U14601 (N_14601,N_8084,N_7623);
or U14602 (N_14602,N_9942,N_5971);
and U14603 (N_14603,N_5177,N_9068);
nor U14604 (N_14604,N_9966,N_8133);
xor U14605 (N_14605,N_8099,N_7451);
nor U14606 (N_14606,N_6395,N_8540);
nor U14607 (N_14607,N_8284,N_9142);
nor U14608 (N_14608,N_9948,N_5683);
nand U14609 (N_14609,N_7789,N_6954);
xor U14610 (N_14610,N_6564,N_7791);
or U14611 (N_14611,N_5578,N_8112);
nor U14612 (N_14612,N_8570,N_5299);
xor U14613 (N_14613,N_8918,N_7812);
nand U14614 (N_14614,N_7746,N_6738);
nand U14615 (N_14615,N_9515,N_5707);
xnor U14616 (N_14616,N_6414,N_6842);
nor U14617 (N_14617,N_6918,N_6183);
and U14618 (N_14618,N_9716,N_8815);
nor U14619 (N_14619,N_5783,N_6206);
nand U14620 (N_14620,N_8393,N_7674);
nand U14621 (N_14621,N_6251,N_6322);
nand U14622 (N_14622,N_7125,N_8998);
xor U14623 (N_14623,N_5863,N_9219);
nand U14624 (N_14624,N_9120,N_7255);
nor U14625 (N_14625,N_7694,N_6418);
nand U14626 (N_14626,N_8160,N_9681);
nor U14627 (N_14627,N_5317,N_5692);
or U14628 (N_14628,N_6911,N_6854);
nor U14629 (N_14629,N_8891,N_6603);
or U14630 (N_14630,N_5722,N_8074);
nor U14631 (N_14631,N_7773,N_9582);
or U14632 (N_14632,N_8051,N_7285);
nor U14633 (N_14633,N_6464,N_6567);
xor U14634 (N_14634,N_6021,N_8204);
nand U14635 (N_14635,N_9833,N_9916);
and U14636 (N_14636,N_5928,N_6166);
nor U14637 (N_14637,N_8628,N_6616);
nor U14638 (N_14638,N_6433,N_6431);
nand U14639 (N_14639,N_5531,N_8248);
nand U14640 (N_14640,N_5804,N_9991);
and U14641 (N_14641,N_8615,N_7193);
xnor U14642 (N_14642,N_9646,N_6433);
and U14643 (N_14643,N_6269,N_7629);
or U14644 (N_14644,N_7457,N_6528);
nor U14645 (N_14645,N_5076,N_9625);
nand U14646 (N_14646,N_6860,N_5286);
nor U14647 (N_14647,N_6911,N_7714);
nor U14648 (N_14648,N_5704,N_5874);
xnor U14649 (N_14649,N_8390,N_7364);
and U14650 (N_14650,N_7117,N_5776);
nand U14651 (N_14651,N_5819,N_7849);
and U14652 (N_14652,N_6515,N_8338);
nand U14653 (N_14653,N_8675,N_7444);
xor U14654 (N_14654,N_6820,N_5464);
and U14655 (N_14655,N_8878,N_7703);
and U14656 (N_14656,N_6600,N_8464);
nor U14657 (N_14657,N_8831,N_5604);
xnor U14658 (N_14658,N_9060,N_5571);
nand U14659 (N_14659,N_9337,N_8590);
or U14660 (N_14660,N_9597,N_6097);
nor U14661 (N_14661,N_6535,N_5662);
xor U14662 (N_14662,N_6842,N_8612);
or U14663 (N_14663,N_9846,N_9845);
or U14664 (N_14664,N_7092,N_7335);
nand U14665 (N_14665,N_9143,N_7456);
or U14666 (N_14666,N_5999,N_9903);
nand U14667 (N_14667,N_5875,N_9545);
or U14668 (N_14668,N_7958,N_8933);
and U14669 (N_14669,N_5610,N_8092);
nor U14670 (N_14670,N_9174,N_9135);
and U14671 (N_14671,N_8382,N_6410);
nor U14672 (N_14672,N_9705,N_9843);
xnor U14673 (N_14673,N_8544,N_9677);
nand U14674 (N_14674,N_6385,N_5891);
xnor U14675 (N_14675,N_5942,N_5780);
nand U14676 (N_14676,N_6625,N_7924);
nand U14677 (N_14677,N_8797,N_5983);
nand U14678 (N_14678,N_7925,N_9342);
nand U14679 (N_14679,N_8157,N_5897);
xor U14680 (N_14680,N_7767,N_5706);
xnor U14681 (N_14681,N_5608,N_9358);
nand U14682 (N_14682,N_6368,N_6762);
or U14683 (N_14683,N_8524,N_6152);
or U14684 (N_14684,N_6244,N_7545);
nor U14685 (N_14685,N_5130,N_6314);
nand U14686 (N_14686,N_8899,N_5976);
or U14687 (N_14687,N_9584,N_5022);
and U14688 (N_14688,N_8445,N_5021);
or U14689 (N_14689,N_7748,N_9201);
nand U14690 (N_14690,N_8474,N_6957);
and U14691 (N_14691,N_5379,N_8525);
or U14692 (N_14692,N_8654,N_9044);
or U14693 (N_14693,N_9361,N_8429);
or U14694 (N_14694,N_7644,N_7539);
nand U14695 (N_14695,N_5633,N_6687);
or U14696 (N_14696,N_7367,N_9895);
or U14697 (N_14697,N_7667,N_9927);
xnor U14698 (N_14698,N_7615,N_8245);
nand U14699 (N_14699,N_5646,N_6148);
xnor U14700 (N_14700,N_9601,N_6296);
xnor U14701 (N_14701,N_9618,N_9309);
or U14702 (N_14702,N_7789,N_8623);
and U14703 (N_14703,N_7217,N_5441);
or U14704 (N_14704,N_8279,N_7798);
nand U14705 (N_14705,N_5095,N_8068);
and U14706 (N_14706,N_7696,N_8217);
and U14707 (N_14707,N_5913,N_6983);
nand U14708 (N_14708,N_9513,N_5942);
or U14709 (N_14709,N_6864,N_7473);
xnor U14710 (N_14710,N_5238,N_9502);
nand U14711 (N_14711,N_8865,N_6097);
nor U14712 (N_14712,N_8886,N_5092);
xor U14713 (N_14713,N_7956,N_8691);
nor U14714 (N_14714,N_8561,N_8052);
xnor U14715 (N_14715,N_8437,N_8347);
or U14716 (N_14716,N_9040,N_9794);
xnor U14717 (N_14717,N_8517,N_5995);
nor U14718 (N_14718,N_7704,N_6903);
or U14719 (N_14719,N_8660,N_5244);
and U14720 (N_14720,N_6865,N_8527);
xnor U14721 (N_14721,N_5061,N_8586);
nor U14722 (N_14722,N_6818,N_5893);
nand U14723 (N_14723,N_9937,N_9697);
xor U14724 (N_14724,N_5081,N_9106);
xnor U14725 (N_14725,N_7287,N_5793);
nand U14726 (N_14726,N_7586,N_8750);
and U14727 (N_14727,N_9812,N_7635);
and U14728 (N_14728,N_8321,N_6915);
nand U14729 (N_14729,N_7973,N_6749);
and U14730 (N_14730,N_9278,N_7243);
or U14731 (N_14731,N_7780,N_5646);
or U14732 (N_14732,N_8166,N_9573);
nand U14733 (N_14733,N_8190,N_6737);
or U14734 (N_14734,N_9808,N_9377);
and U14735 (N_14735,N_5381,N_6922);
nor U14736 (N_14736,N_7391,N_7445);
or U14737 (N_14737,N_6099,N_7077);
and U14738 (N_14738,N_9986,N_9682);
or U14739 (N_14739,N_8623,N_9324);
or U14740 (N_14740,N_7933,N_5707);
and U14741 (N_14741,N_5023,N_5026);
xor U14742 (N_14742,N_9365,N_7504);
nand U14743 (N_14743,N_7894,N_5375);
xnor U14744 (N_14744,N_8550,N_8289);
nand U14745 (N_14745,N_8060,N_5521);
and U14746 (N_14746,N_9625,N_8548);
xor U14747 (N_14747,N_6770,N_8618);
or U14748 (N_14748,N_5951,N_7489);
or U14749 (N_14749,N_5130,N_5782);
or U14750 (N_14750,N_7970,N_9122);
or U14751 (N_14751,N_5265,N_9185);
and U14752 (N_14752,N_6039,N_6739);
xor U14753 (N_14753,N_5409,N_6082);
nand U14754 (N_14754,N_5399,N_9212);
xor U14755 (N_14755,N_5479,N_5090);
nand U14756 (N_14756,N_5573,N_5113);
nor U14757 (N_14757,N_5054,N_5912);
nand U14758 (N_14758,N_8226,N_5620);
nand U14759 (N_14759,N_6500,N_8032);
xnor U14760 (N_14760,N_9073,N_6661);
xnor U14761 (N_14761,N_8975,N_5637);
nor U14762 (N_14762,N_6294,N_5058);
and U14763 (N_14763,N_6833,N_9359);
nand U14764 (N_14764,N_7732,N_9142);
nor U14765 (N_14765,N_6634,N_8757);
nor U14766 (N_14766,N_6938,N_6183);
nand U14767 (N_14767,N_8788,N_5008);
or U14768 (N_14768,N_6805,N_9072);
nor U14769 (N_14769,N_9700,N_8763);
nor U14770 (N_14770,N_9039,N_6528);
xnor U14771 (N_14771,N_6847,N_7753);
xor U14772 (N_14772,N_8824,N_6393);
or U14773 (N_14773,N_7922,N_9717);
xnor U14774 (N_14774,N_8710,N_8351);
or U14775 (N_14775,N_9308,N_6458);
or U14776 (N_14776,N_8576,N_7145);
nand U14777 (N_14777,N_5693,N_6885);
xor U14778 (N_14778,N_5570,N_5428);
and U14779 (N_14779,N_6650,N_7799);
nor U14780 (N_14780,N_5560,N_5720);
and U14781 (N_14781,N_8524,N_6443);
or U14782 (N_14782,N_5060,N_7228);
nand U14783 (N_14783,N_6340,N_8754);
xor U14784 (N_14784,N_8109,N_7394);
and U14785 (N_14785,N_8135,N_5298);
nand U14786 (N_14786,N_5453,N_8491);
or U14787 (N_14787,N_6102,N_8416);
and U14788 (N_14788,N_7121,N_5886);
nor U14789 (N_14789,N_8973,N_9134);
nand U14790 (N_14790,N_7447,N_5225);
nand U14791 (N_14791,N_8842,N_5718);
and U14792 (N_14792,N_6592,N_6342);
nand U14793 (N_14793,N_9656,N_7908);
and U14794 (N_14794,N_8615,N_7014);
xor U14795 (N_14795,N_5942,N_8546);
nor U14796 (N_14796,N_5440,N_7263);
nor U14797 (N_14797,N_6271,N_5960);
xor U14798 (N_14798,N_6663,N_9112);
nand U14799 (N_14799,N_8589,N_6404);
or U14800 (N_14800,N_9866,N_9296);
nor U14801 (N_14801,N_8201,N_5243);
or U14802 (N_14802,N_8769,N_6969);
xor U14803 (N_14803,N_6134,N_9188);
nor U14804 (N_14804,N_6587,N_7378);
xnor U14805 (N_14805,N_7280,N_7849);
or U14806 (N_14806,N_8916,N_9559);
or U14807 (N_14807,N_9100,N_7232);
and U14808 (N_14808,N_7757,N_8390);
and U14809 (N_14809,N_9119,N_9454);
nand U14810 (N_14810,N_5694,N_6581);
nor U14811 (N_14811,N_5866,N_6489);
nand U14812 (N_14812,N_6796,N_7819);
xnor U14813 (N_14813,N_8757,N_6641);
and U14814 (N_14814,N_9160,N_9934);
or U14815 (N_14815,N_8329,N_7648);
or U14816 (N_14816,N_8299,N_7351);
nor U14817 (N_14817,N_9227,N_5587);
and U14818 (N_14818,N_8884,N_7997);
nor U14819 (N_14819,N_5629,N_8996);
xor U14820 (N_14820,N_9937,N_7353);
xor U14821 (N_14821,N_8137,N_9368);
nand U14822 (N_14822,N_9156,N_7350);
and U14823 (N_14823,N_8154,N_7510);
xor U14824 (N_14824,N_5485,N_7741);
xnor U14825 (N_14825,N_8392,N_8246);
and U14826 (N_14826,N_7014,N_6311);
or U14827 (N_14827,N_9660,N_8047);
nor U14828 (N_14828,N_5052,N_7056);
and U14829 (N_14829,N_9958,N_5310);
nand U14830 (N_14830,N_9445,N_7975);
or U14831 (N_14831,N_7202,N_8702);
nand U14832 (N_14832,N_6059,N_8973);
or U14833 (N_14833,N_6624,N_6188);
and U14834 (N_14834,N_6595,N_7907);
nand U14835 (N_14835,N_5043,N_9876);
or U14836 (N_14836,N_7349,N_6938);
xor U14837 (N_14837,N_8819,N_5777);
and U14838 (N_14838,N_5538,N_5350);
and U14839 (N_14839,N_9085,N_8009);
and U14840 (N_14840,N_8388,N_6399);
nor U14841 (N_14841,N_8124,N_6299);
nand U14842 (N_14842,N_9586,N_5214);
xnor U14843 (N_14843,N_8327,N_7007);
and U14844 (N_14844,N_5130,N_8028);
xor U14845 (N_14845,N_5301,N_9339);
or U14846 (N_14846,N_8412,N_8892);
or U14847 (N_14847,N_9831,N_7633);
and U14848 (N_14848,N_5586,N_9162);
xnor U14849 (N_14849,N_9232,N_7885);
xor U14850 (N_14850,N_7846,N_7421);
nor U14851 (N_14851,N_9182,N_5219);
and U14852 (N_14852,N_9914,N_6465);
nor U14853 (N_14853,N_9617,N_5126);
nor U14854 (N_14854,N_7410,N_9870);
or U14855 (N_14855,N_8535,N_5856);
and U14856 (N_14856,N_7740,N_5923);
or U14857 (N_14857,N_8866,N_7611);
nor U14858 (N_14858,N_8712,N_9834);
or U14859 (N_14859,N_5270,N_6564);
xor U14860 (N_14860,N_5969,N_7212);
nand U14861 (N_14861,N_7119,N_7873);
and U14862 (N_14862,N_6328,N_7889);
xnor U14863 (N_14863,N_8892,N_9049);
and U14864 (N_14864,N_8825,N_7069);
xor U14865 (N_14865,N_6486,N_8427);
or U14866 (N_14866,N_6982,N_6071);
and U14867 (N_14867,N_5876,N_6089);
xnor U14868 (N_14868,N_8735,N_8964);
nand U14869 (N_14869,N_9658,N_8220);
nor U14870 (N_14870,N_6041,N_9918);
and U14871 (N_14871,N_8695,N_7549);
nor U14872 (N_14872,N_7207,N_9338);
nand U14873 (N_14873,N_8073,N_8108);
xor U14874 (N_14874,N_9147,N_9348);
and U14875 (N_14875,N_8793,N_5404);
or U14876 (N_14876,N_9454,N_7075);
or U14877 (N_14877,N_9088,N_5519);
nor U14878 (N_14878,N_5896,N_5742);
nor U14879 (N_14879,N_9890,N_6573);
or U14880 (N_14880,N_5581,N_7864);
nand U14881 (N_14881,N_6249,N_9290);
nor U14882 (N_14882,N_6115,N_9409);
nand U14883 (N_14883,N_7783,N_6697);
xnor U14884 (N_14884,N_9290,N_6197);
nor U14885 (N_14885,N_9712,N_5351);
or U14886 (N_14886,N_9657,N_9534);
or U14887 (N_14887,N_5700,N_9949);
nand U14888 (N_14888,N_7890,N_8998);
xnor U14889 (N_14889,N_9089,N_8236);
nor U14890 (N_14890,N_9914,N_5084);
nor U14891 (N_14891,N_8624,N_6761);
or U14892 (N_14892,N_7236,N_6121);
nand U14893 (N_14893,N_8156,N_5135);
nor U14894 (N_14894,N_6547,N_6232);
nand U14895 (N_14895,N_7094,N_9696);
xor U14896 (N_14896,N_7151,N_5858);
or U14897 (N_14897,N_9090,N_5777);
nor U14898 (N_14898,N_8240,N_9885);
xnor U14899 (N_14899,N_7794,N_8865);
or U14900 (N_14900,N_7323,N_9720);
and U14901 (N_14901,N_6350,N_9445);
and U14902 (N_14902,N_8728,N_9535);
xor U14903 (N_14903,N_6473,N_6837);
nand U14904 (N_14904,N_5650,N_9532);
xnor U14905 (N_14905,N_5964,N_6792);
or U14906 (N_14906,N_5669,N_8545);
or U14907 (N_14907,N_9642,N_7347);
nor U14908 (N_14908,N_8580,N_9138);
xor U14909 (N_14909,N_9396,N_8633);
xor U14910 (N_14910,N_9801,N_8860);
or U14911 (N_14911,N_8950,N_7360);
nand U14912 (N_14912,N_5605,N_5644);
or U14913 (N_14913,N_5496,N_7063);
or U14914 (N_14914,N_7370,N_6470);
xnor U14915 (N_14915,N_8994,N_5181);
and U14916 (N_14916,N_5897,N_6963);
or U14917 (N_14917,N_9608,N_7090);
nor U14918 (N_14918,N_8573,N_6187);
or U14919 (N_14919,N_6598,N_9723);
xnor U14920 (N_14920,N_7545,N_7855);
nor U14921 (N_14921,N_9454,N_6547);
and U14922 (N_14922,N_7104,N_6043);
and U14923 (N_14923,N_9477,N_8389);
nand U14924 (N_14924,N_7749,N_9977);
nor U14925 (N_14925,N_9048,N_6408);
or U14926 (N_14926,N_6311,N_6021);
nor U14927 (N_14927,N_9394,N_7999);
or U14928 (N_14928,N_9468,N_6649);
and U14929 (N_14929,N_5809,N_5005);
and U14930 (N_14930,N_9402,N_7169);
nand U14931 (N_14931,N_6422,N_5831);
nand U14932 (N_14932,N_8695,N_8562);
and U14933 (N_14933,N_9231,N_9539);
or U14934 (N_14934,N_5617,N_5521);
or U14935 (N_14935,N_5255,N_6518);
xor U14936 (N_14936,N_8806,N_5629);
or U14937 (N_14937,N_8781,N_7229);
or U14938 (N_14938,N_5220,N_5828);
xor U14939 (N_14939,N_9290,N_7265);
nand U14940 (N_14940,N_6906,N_8238);
and U14941 (N_14941,N_8573,N_8025);
xnor U14942 (N_14942,N_7009,N_9631);
and U14943 (N_14943,N_8550,N_9621);
and U14944 (N_14944,N_8908,N_6785);
nand U14945 (N_14945,N_7416,N_7928);
xnor U14946 (N_14946,N_7578,N_5528);
nor U14947 (N_14947,N_7262,N_7729);
or U14948 (N_14948,N_5093,N_9634);
xnor U14949 (N_14949,N_8277,N_7570);
nand U14950 (N_14950,N_7862,N_8161);
xor U14951 (N_14951,N_9640,N_8825);
and U14952 (N_14952,N_8845,N_9609);
nor U14953 (N_14953,N_8489,N_6620);
or U14954 (N_14954,N_6256,N_6192);
xor U14955 (N_14955,N_7312,N_7172);
or U14956 (N_14956,N_8591,N_6968);
xor U14957 (N_14957,N_8244,N_5419);
nor U14958 (N_14958,N_8862,N_6994);
nand U14959 (N_14959,N_7904,N_6291);
xor U14960 (N_14960,N_7582,N_6849);
or U14961 (N_14961,N_8317,N_7486);
or U14962 (N_14962,N_8856,N_7219);
nand U14963 (N_14963,N_5115,N_9690);
nand U14964 (N_14964,N_5384,N_9684);
xnor U14965 (N_14965,N_6028,N_9736);
nand U14966 (N_14966,N_6908,N_6445);
and U14967 (N_14967,N_6127,N_7320);
xnor U14968 (N_14968,N_9475,N_9113);
or U14969 (N_14969,N_7496,N_8233);
xor U14970 (N_14970,N_8381,N_6028);
nand U14971 (N_14971,N_6471,N_5359);
nand U14972 (N_14972,N_5018,N_8862);
and U14973 (N_14973,N_7852,N_7411);
nor U14974 (N_14974,N_8778,N_9359);
nor U14975 (N_14975,N_8243,N_9059);
xnor U14976 (N_14976,N_9909,N_6113);
nand U14977 (N_14977,N_8100,N_7473);
and U14978 (N_14978,N_6390,N_7997);
or U14979 (N_14979,N_7305,N_6659);
or U14980 (N_14980,N_8147,N_9725);
and U14981 (N_14981,N_8661,N_8715);
nand U14982 (N_14982,N_7731,N_9613);
and U14983 (N_14983,N_5587,N_7002);
or U14984 (N_14984,N_6685,N_6776);
or U14985 (N_14985,N_9597,N_7968);
nand U14986 (N_14986,N_8874,N_9185);
and U14987 (N_14987,N_6911,N_9466);
and U14988 (N_14988,N_9963,N_6853);
xor U14989 (N_14989,N_9468,N_6366);
or U14990 (N_14990,N_7879,N_7764);
nand U14991 (N_14991,N_5366,N_9116);
and U14992 (N_14992,N_6653,N_7185);
and U14993 (N_14993,N_7970,N_6813);
and U14994 (N_14994,N_6915,N_9964);
nor U14995 (N_14995,N_7369,N_6711);
or U14996 (N_14996,N_9563,N_8613);
nor U14997 (N_14997,N_8217,N_6348);
or U14998 (N_14998,N_8529,N_5153);
nor U14999 (N_14999,N_6105,N_7677);
nand U15000 (N_15000,N_11376,N_12554);
nand U15001 (N_15001,N_12310,N_11224);
xnor U15002 (N_15002,N_10898,N_14633);
xor U15003 (N_15003,N_10343,N_13974);
and U15004 (N_15004,N_12701,N_12475);
nor U15005 (N_15005,N_10695,N_13028);
nor U15006 (N_15006,N_13708,N_13246);
or U15007 (N_15007,N_11317,N_11504);
xor U15008 (N_15008,N_12488,N_14165);
and U15009 (N_15009,N_10203,N_14013);
nor U15010 (N_15010,N_10029,N_11795);
nor U15011 (N_15011,N_11764,N_14915);
and U15012 (N_15012,N_11236,N_13543);
xnor U15013 (N_15013,N_11731,N_14523);
and U15014 (N_15014,N_12532,N_12582);
xnor U15015 (N_15015,N_12404,N_11886);
nand U15016 (N_15016,N_13448,N_12122);
nand U15017 (N_15017,N_14864,N_14166);
nor U15018 (N_15018,N_14702,N_11331);
nor U15019 (N_15019,N_14415,N_12640);
nand U15020 (N_15020,N_14770,N_14392);
xnor U15021 (N_15021,N_10878,N_13113);
and U15022 (N_15022,N_10706,N_12104);
nand U15023 (N_15023,N_14641,N_12023);
nor U15024 (N_15024,N_13923,N_11565);
nor U15025 (N_15025,N_13822,N_10119);
xnor U15026 (N_15026,N_12694,N_13373);
nand U15027 (N_15027,N_13627,N_13789);
nor U15028 (N_15028,N_13542,N_11145);
xor U15029 (N_15029,N_11312,N_13411);
nor U15030 (N_15030,N_14637,N_10676);
xnor U15031 (N_15031,N_14494,N_14146);
or U15032 (N_15032,N_11509,N_14958);
nor U15033 (N_15033,N_10985,N_11086);
nand U15034 (N_15034,N_12092,N_11061);
xnor U15035 (N_15035,N_12621,N_10047);
xor U15036 (N_15036,N_11664,N_12539);
nor U15037 (N_15037,N_12505,N_13804);
or U15038 (N_15038,N_11265,N_11794);
nand U15039 (N_15039,N_10489,N_12825);
nand U15040 (N_15040,N_14480,N_13131);
or U15041 (N_15041,N_13519,N_14881);
xor U15042 (N_15042,N_11448,N_11359);
xnor U15043 (N_15043,N_13532,N_13250);
xor U15044 (N_15044,N_12178,N_12970);
or U15045 (N_15045,N_10429,N_11953);
xnor U15046 (N_15046,N_12879,N_12452);
xnor U15047 (N_15047,N_12735,N_11816);
nor U15048 (N_15048,N_11153,N_10095);
xor U15049 (N_15049,N_10288,N_12135);
xnor U15050 (N_15050,N_11539,N_10351);
nand U15051 (N_15051,N_12343,N_10557);
or U15052 (N_15052,N_14732,N_13092);
nor U15053 (N_15053,N_13317,N_12124);
and U15054 (N_15054,N_14125,N_12171);
or U15055 (N_15055,N_10713,N_12704);
or U15056 (N_15056,N_12821,N_12990);
and U15057 (N_15057,N_10884,N_10425);
nand U15058 (N_15058,N_14466,N_12644);
nor U15059 (N_15059,N_10941,N_12798);
and U15060 (N_15060,N_13468,N_12168);
or U15061 (N_15061,N_12275,N_12056);
nor U15062 (N_15062,N_14357,N_12746);
nor U15063 (N_15063,N_14446,N_14743);
or U15064 (N_15064,N_10322,N_10330);
and U15065 (N_15065,N_14512,N_10460);
or U15066 (N_15066,N_14911,N_14023);
xnor U15067 (N_15067,N_10090,N_12051);
nor U15068 (N_15068,N_11639,N_13563);
or U15069 (N_15069,N_12271,N_14216);
nand U15070 (N_15070,N_11981,N_12829);
and U15071 (N_15071,N_12221,N_10831);
or U15072 (N_15072,N_13692,N_12363);
nor U15073 (N_15073,N_12875,N_12526);
or U15074 (N_15074,N_11056,N_11459);
nor U15075 (N_15075,N_12045,N_14913);
nand U15076 (N_15076,N_14376,N_10862);
or U15077 (N_15077,N_10587,N_12492);
xnor U15078 (N_15078,N_13925,N_11295);
nand U15079 (N_15079,N_11892,N_11353);
nand U15080 (N_15080,N_14812,N_13333);
nand U15081 (N_15081,N_13027,N_13947);
or U15082 (N_15082,N_10163,N_14488);
nor U15083 (N_15083,N_13104,N_11972);
xor U15084 (N_15084,N_11610,N_13331);
nor U15085 (N_15085,N_14140,N_14244);
or U15086 (N_15086,N_12708,N_10164);
nand U15087 (N_15087,N_11782,N_10341);
or U15088 (N_15088,N_10156,N_13485);
nand U15089 (N_15089,N_11567,N_11911);
nor U15090 (N_15090,N_10060,N_10807);
nor U15091 (N_15091,N_11158,N_11860);
nand U15092 (N_15092,N_14282,N_13042);
nor U15093 (N_15093,N_10055,N_14492);
nand U15094 (N_15094,N_13462,N_14416);
xor U15095 (N_15095,N_12066,N_12776);
xor U15096 (N_15096,N_14946,N_12443);
nor U15097 (N_15097,N_10893,N_11307);
xnor U15098 (N_15098,N_13861,N_14631);
xor U15099 (N_15099,N_13157,N_13545);
xnor U15100 (N_15100,N_10499,N_12804);
nand U15101 (N_15101,N_12453,N_12855);
nand U15102 (N_15102,N_10327,N_14226);
nand U15103 (N_15103,N_10923,N_14352);
nor U15104 (N_15104,N_13480,N_14517);
xnor U15105 (N_15105,N_12136,N_10685);
nand U15106 (N_15106,N_10181,N_11470);
and U15107 (N_15107,N_14402,N_14299);
xnor U15108 (N_15108,N_11979,N_14039);
nor U15109 (N_15109,N_14027,N_11793);
nand U15110 (N_15110,N_11568,N_12478);
or U15111 (N_15111,N_11658,N_11582);
nor U15112 (N_15112,N_14481,N_11776);
nor U15113 (N_15113,N_11123,N_12446);
and U15114 (N_15114,N_14590,N_12751);
nand U15115 (N_15115,N_11306,N_13339);
xnor U15116 (N_15116,N_12458,N_11228);
nor U15117 (N_15117,N_12741,N_11573);
or U15118 (N_15118,N_12329,N_13083);
and U15119 (N_15119,N_14869,N_11643);
and U15120 (N_15120,N_12976,N_12146);
or U15121 (N_15121,N_14464,N_10574);
nand U15122 (N_15122,N_13959,N_10751);
or U15123 (N_15123,N_13605,N_12797);
and U15124 (N_15124,N_12083,N_13033);
nor U15125 (N_15125,N_12448,N_11717);
nand U15126 (N_15126,N_11115,N_13016);
nand U15127 (N_15127,N_14180,N_12042);
nor U15128 (N_15128,N_14629,N_10744);
xor U15129 (N_15129,N_14619,N_10073);
nor U15130 (N_15130,N_13522,N_10819);
and U15131 (N_15131,N_12223,N_12713);
xor U15132 (N_15132,N_14826,N_13848);
xor U15133 (N_15133,N_12318,N_13856);
nand U15134 (N_15134,N_11309,N_13548);
nor U15135 (N_15135,N_11695,N_13384);
and U15136 (N_15136,N_13957,N_11308);
and U15137 (N_15137,N_14171,N_10225);
nor U15138 (N_15138,N_12828,N_12913);
or U15139 (N_15139,N_14583,N_14868);
and U15140 (N_15140,N_11476,N_11824);
and U15141 (N_15141,N_12336,N_10357);
or U15142 (N_15142,N_11357,N_10293);
nand U15143 (N_15143,N_13503,N_13224);
nor U15144 (N_15144,N_10767,N_14874);
or U15145 (N_15145,N_10701,N_10222);
nand U15146 (N_15146,N_13364,N_10764);
xor U15147 (N_15147,N_10911,N_14916);
nor U15148 (N_15148,N_10909,N_14181);
and U15149 (N_15149,N_13827,N_10199);
nand U15150 (N_15150,N_14405,N_11447);
nor U15151 (N_15151,N_14752,N_11008);
nand U15152 (N_15152,N_14294,N_13953);
and U15153 (N_15153,N_14432,N_11769);
and U15154 (N_15154,N_10588,N_12173);
and U15155 (N_15155,N_12650,N_10753);
or U15156 (N_15156,N_13460,N_14932);
and U15157 (N_15157,N_10980,N_14143);
xnor U15158 (N_15158,N_10062,N_10715);
nor U15159 (N_15159,N_12624,N_11606);
xor U15160 (N_15160,N_10195,N_13783);
nand U15161 (N_15161,N_10691,N_14960);
xor U15162 (N_15162,N_11190,N_14440);
nand U15163 (N_15163,N_12430,N_13930);
xnor U15164 (N_15164,N_10771,N_13751);
or U15165 (N_15165,N_12962,N_10883);
nor U15166 (N_15166,N_11572,N_11547);
and U15167 (N_15167,N_12327,N_11259);
nor U15168 (N_15168,N_11529,N_13523);
nor U15169 (N_15169,N_14414,N_13035);
nand U15170 (N_15170,N_12082,N_10197);
xnor U15171 (N_15171,N_13866,N_10436);
nor U15172 (N_15172,N_11135,N_13053);
nand U15173 (N_15173,N_13213,N_11413);
xor U15174 (N_15174,N_11460,N_12961);
nor U15175 (N_15175,N_13271,N_14878);
or U15176 (N_15176,N_12369,N_12907);
nand U15177 (N_15177,N_10159,N_14329);
xnor U15178 (N_15178,N_10053,N_10028);
nand U15179 (N_15179,N_11961,N_11918);
or U15180 (N_15180,N_13630,N_10799);
xor U15181 (N_15181,N_12859,N_10537);
and U15182 (N_15182,N_14058,N_11449);
nand U15183 (N_15183,N_14136,N_14311);
and U15184 (N_15184,N_11663,N_11045);
xor U15185 (N_15185,N_12188,N_14444);
xnor U15186 (N_15186,N_10054,N_14876);
xor U15187 (N_15187,N_12884,N_12682);
nand U15188 (N_15188,N_10252,N_12177);
and U15189 (N_15189,N_11399,N_10950);
and U15190 (N_15190,N_13867,N_13119);
nand U15191 (N_15191,N_13290,N_14620);
xor U15192 (N_15192,N_10068,N_14264);
nand U15193 (N_15193,N_11686,N_11724);
nand U15194 (N_15194,N_14062,N_13006);
nand U15195 (N_15195,N_14241,N_12212);
and U15196 (N_15196,N_12528,N_10612);
and U15197 (N_15197,N_11623,N_11131);
xnor U15198 (N_15198,N_10255,N_13628);
or U15199 (N_15199,N_10396,N_11755);
xor U15200 (N_15200,N_10103,N_12189);
xor U15201 (N_15201,N_13977,N_14438);
and U15202 (N_15202,N_10498,N_14575);
nor U15203 (N_15203,N_11942,N_13729);
and U15204 (N_15204,N_12565,N_11429);
nand U15205 (N_15205,N_14778,N_11900);
or U15206 (N_15206,N_11833,N_14727);
and U15207 (N_15207,N_14587,N_13658);
nor U15208 (N_15208,N_12257,N_10920);
nand U15209 (N_15209,N_13836,N_14418);
and U15210 (N_15210,N_10385,N_11347);
xnor U15211 (N_15211,N_13277,N_11469);
xnor U15212 (N_15212,N_14157,N_10270);
and U15213 (N_15213,N_11091,N_13709);
nand U15214 (N_15214,N_11920,N_10345);
and U15215 (N_15215,N_13732,N_10809);
xor U15216 (N_15216,N_14502,N_14212);
nor U15217 (N_15217,N_13539,N_11126);
nor U15218 (N_15218,N_10242,N_12818);
xor U15219 (N_15219,N_13178,N_11600);
nand U15220 (N_15220,N_12549,N_13245);
or U15221 (N_15221,N_12214,N_10021);
xnor U15222 (N_15222,N_14345,N_14367);
or U15223 (N_15223,N_14249,N_10360);
nor U15224 (N_15224,N_11531,N_12808);
nor U15225 (N_15225,N_12249,N_10008);
and U15226 (N_15226,N_10440,N_13349);
nor U15227 (N_15227,N_11859,N_12198);
or U15228 (N_15228,N_10972,N_11074);
nor U15229 (N_15229,N_10863,N_10525);
nor U15230 (N_15230,N_10998,N_14147);
nand U15231 (N_15231,N_13334,N_14597);
and U15232 (N_15232,N_13785,N_10682);
nor U15233 (N_15233,N_10067,N_13014);
nand U15234 (N_15234,N_13886,N_10527);
and U15235 (N_15235,N_14159,N_11311);
and U15236 (N_15236,N_14603,N_12611);
nor U15237 (N_15237,N_14663,N_12282);
nand U15238 (N_15238,N_11798,N_13038);
nand U15239 (N_15239,N_14956,N_10124);
or U15240 (N_15240,N_11327,N_14186);
or U15241 (N_15241,N_10522,N_10412);
nor U15242 (N_15242,N_13499,N_14119);
or U15243 (N_15243,N_11530,N_11473);
xor U15244 (N_15244,N_12344,N_12498);
xnor U15245 (N_15245,N_13447,N_13778);
and U15246 (N_15246,N_14032,N_11551);
and U15247 (N_15247,N_14089,N_12101);
or U15248 (N_15248,N_14493,N_10240);
and U15249 (N_15249,N_12464,N_14269);
xnor U15250 (N_15250,N_10470,N_10613);
and U15251 (N_15251,N_10206,N_10669);
or U15252 (N_15252,N_13336,N_11017);
nor U15253 (N_15253,N_14767,N_12347);
xnor U15254 (N_15254,N_13222,N_12004);
or U15255 (N_15255,N_11758,N_13763);
nand U15256 (N_15256,N_14025,N_13531);
or U15257 (N_15257,N_12634,N_11337);
nor U15258 (N_15258,N_13483,N_10958);
xnor U15259 (N_15259,N_12115,N_14452);
nor U15260 (N_15260,N_12071,N_11648);
nor U15261 (N_15261,N_12424,N_10606);
and U15262 (N_15262,N_11746,N_12956);
nor U15263 (N_15263,N_11070,N_12462);
or U15264 (N_15264,N_14364,N_13425);
and U15265 (N_15265,N_13635,N_14175);
or U15266 (N_15266,N_10916,N_11258);
and U15267 (N_15267,N_11208,N_11174);
and U15268 (N_15268,N_11092,N_10010);
nor U15269 (N_15269,N_14307,N_12312);
nand U15270 (N_15270,N_12372,N_10474);
xor U15271 (N_15271,N_10485,N_11587);
nand U15272 (N_15272,N_10108,N_13444);
nand U15273 (N_15273,N_12264,N_13819);
and U15274 (N_15274,N_10617,N_12158);
xor U15275 (N_15275,N_11986,N_12623);
nand U15276 (N_15276,N_11039,N_13908);
and U15277 (N_15277,N_14694,N_11642);
xnor U15278 (N_15278,N_13674,N_11322);
and U15279 (N_15279,N_12762,N_14983);
xor U15280 (N_15280,N_13897,N_14453);
and U15281 (N_15281,N_13601,N_14592);
xor U15282 (N_15282,N_14951,N_10148);
and U15283 (N_15283,N_13525,N_14534);
xor U15284 (N_15284,N_14542,N_13368);
or U15285 (N_15285,N_10439,N_14532);
nand U15286 (N_15286,N_12721,N_10832);
xor U15287 (N_15287,N_10076,N_10860);
or U15288 (N_15288,N_12631,N_12972);
nor U15289 (N_15289,N_12491,N_12387);
nor U15290 (N_15290,N_14277,N_12468);
nand U15291 (N_15291,N_14483,N_12518);
or U15292 (N_15292,N_10530,N_12924);
nand U15293 (N_15293,N_12848,N_10871);
nor U15294 (N_15294,N_11405,N_11584);
nor U15295 (N_15295,N_10409,N_10660);
or U15296 (N_15296,N_14861,N_10800);
nor U15297 (N_15297,N_12108,N_10447);
nand U15298 (N_15298,N_10504,N_11052);
and U15299 (N_15299,N_13870,N_12227);
nor U15300 (N_15300,N_13585,N_10162);
nor U15301 (N_15301,N_14035,N_10569);
or U15302 (N_15302,N_14191,N_10654);
nand U15303 (N_15303,N_11621,N_10734);
nand U15304 (N_15304,N_11913,N_14061);
nor U15305 (N_15305,N_11006,N_13109);
and U15306 (N_15306,N_10657,N_12166);
nand U15307 (N_15307,N_11738,N_11111);
and U15308 (N_15308,N_12752,N_12703);
and U15309 (N_15309,N_13646,N_11586);
or U15310 (N_15310,N_13849,N_13566);
xor U15311 (N_15311,N_14339,N_11189);
nand U15312 (N_15312,N_12881,N_11958);
or U15313 (N_15313,N_13228,N_10708);
nor U15314 (N_15314,N_12159,N_13593);
and U15315 (N_15315,N_11941,N_11287);
or U15316 (N_15316,N_13798,N_10193);
xor U15317 (N_15317,N_13680,N_14552);
and U15318 (N_15318,N_13576,N_12632);
xnor U15319 (N_15319,N_14717,N_10913);
xnor U15320 (N_15320,N_11614,N_13160);
and U15321 (N_15321,N_12637,N_11791);
nand U15322 (N_15322,N_10297,N_12786);
and U15323 (N_15323,N_11493,N_11015);
and U15324 (N_15324,N_14645,N_12295);
xnor U15325 (N_15325,N_10049,N_11428);
nor U15326 (N_15326,N_11465,N_13636);
nand U15327 (N_15327,N_14780,N_14521);
or U15328 (N_15328,N_13003,N_12936);
xnor U15329 (N_15329,N_13573,N_10126);
and U15330 (N_15330,N_11525,N_14894);
nand U15331 (N_15331,N_13326,N_11212);
and U15332 (N_15332,N_13534,N_11779);
or U15333 (N_15333,N_10895,N_14585);
or U15334 (N_15334,N_14662,N_14949);
nand U15335 (N_15335,N_10141,N_11543);
nand U15336 (N_15336,N_11907,N_13530);
nor U15337 (N_15337,N_12268,N_10122);
and U15338 (N_15338,N_11571,N_10621);
or U15339 (N_15339,N_11381,N_13294);
nor U15340 (N_15340,N_12827,N_13495);
nand U15341 (N_15341,N_12068,N_12375);
or U15342 (N_15342,N_13089,N_14704);
nand U15343 (N_15343,N_10750,N_12814);
xor U15344 (N_15344,N_14297,N_14459);
nor U15345 (N_15345,N_12160,N_11954);
xnor U15346 (N_15346,N_14330,N_14621);
xnor U15347 (N_15347,N_13247,N_10284);
and U15348 (N_15348,N_12809,N_10304);
nor U15349 (N_15349,N_10532,N_14153);
nand U15350 (N_15350,N_13441,N_11687);
nor U15351 (N_15351,N_10512,N_10358);
and U15352 (N_15352,N_10872,N_12061);
or U15353 (N_15353,N_10002,N_14320);
xnor U15354 (N_15354,N_11040,N_11766);
nand U15355 (N_15355,N_14404,N_11897);
nor U15356 (N_15356,N_13390,N_11512);
nand U15357 (N_15357,N_11945,N_10097);
nand U15358 (N_15358,N_14707,N_13196);
nor U15359 (N_15359,N_10575,N_11651);
nor U15360 (N_15360,N_13913,N_12081);
nor U15361 (N_15361,N_12049,N_13017);
nand U15362 (N_15362,N_13845,N_11861);
nand U15363 (N_15363,N_11090,N_12568);
xnor U15364 (N_15364,N_10632,N_10216);
nand U15365 (N_15365,N_11369,N_13350);
nand U15366 (N_15366,N_14562,N_14158);
nor U15367 (N_15367,N_10484,N_11894);
or U15368 (N_15368,N_11303,N_10536);
or U15369 (N_15369,N_13973,N_12945);
nor U15370 (N_15370,N_12197,N_11080);
nand U15371 (N_15371,N_14222,N_12963);
and U15372 (N_15372,N_13116,N_13311);
xnor U15373 (N_15373,N_11083,N_10826);
or U15374 (N_15374,N_10317,N_10600);
nand U15375 (N_15375,N_14126,N_14041);
or U15376 (N_15376,N_13405,N_10093);
nand U15377 (N_15377,N_13182,N_12456);
nand U15378 (N_15378,N_12838,N_11721);
nand U15379 (N_15379,N_14625,N_12931);
nand U15380 (N_15380,N_14824,N_12287);
xor U15381 (N_15381,N_12143,N_14677);
nand U15382 (N_15382,N_10890,N_13514);
nand U15383 (N_15383,N_11455,N_11671);
nand U15384 (N_15384,N_11775,N_13962);
nand U15385 (N_15385,N_12987,N_14178);
nor U15386 (N_15386,N_10325,N_12195);
nor U15387 (N_15387,N_10026,N_11851);
nand U15388 (N_15388,N_11637,N_12683);
xnor U15389 (N_15389,N_11423,N_13359);
nand U15390 (N_15390,N_12733,N_14832);
nor U15391 (N_15391,N_11577,N_12839);
nand U15392 (N_15392,N_10684,N_12933);
nor U15393 (N_15393,N_14624,N_13863);
and U15394 (N_15394,N_13642,N_12350);
and U15395 (N_15395,N_10346,N_13996);
nand U15396 (N_15396,N_14496,N_11225);
nand U15397 (N_15397,N_14786,N_14887);
or U15398 (N_15398,N_13101,N_10280);
xnor U15399 (N_15399,N_14725,N_13800);
and U15400 (N_15400,N_13463,N_12399);
nor U15401 (N_15401,N_13031,N_12661);
nand U15402 (N_15402,N_14337,N_13526);
and U15403 (N_15403,N_11274,N_11827);
nor U15404 (N_15404,N_11757,N_12141);
and U15405 (N_15405,N_13992,N_11919);
nor U15406 (N_15406,N_11800,N_12340);
nand U15407 (N_15407,N_14169,N_11268);
or U15408 (N_15408,N_11703,N_10249);
and U15409 (N_15409,N_10548,N_11646);
and U15410 (N_15410,N_12477,N_10269);
xor U15411 (N_15411,N_10810,N_14421);
and U15412 (N_15412,N_11822,N_11254);
or U15413 (N_15413,N_11235,N_14846);
and U15414 (N_15414,N_14616,N_12604);
or U15415 (N_15415,N_14201,N_13188);
or U15416 (N_15416,N_10031,N_14540);
nand U15417 (N_15417,N_10092,N_14685);
xor U15418 (N_15418,N_13123,N_13637);
nand U15419 (N_15419,N_10271,N_11146);
or U15420 (N_15420,N_14845,N_10417);
or U15421 (N_15421,N_12910,N_12610);
nand U15422 (N_15422,N_10785,N_10843);
and U15423 (N_15423,N_12139,N_10075);
and U15424 (N_15424,N_12130,N_10174);
and U15425 (N_15425,N_13676,N_12888);
nor U15426 (N_15426,N_12847,N_12266);
and U15427 (N_15427,N_12515,N_11773);
nor U15428 (N_15428,N_11089,N_14765);
and U15429 (N_15429,N_12841,N_11397);
xnor U15430 (N_15430,N_14463,N_13043);
nor U15431 (N_15431,N_11088,N_13821);
xor U15432 (N_15432,N_11391,N_11472);
or U15433 (N_15433,N_11046,N_13198);
nor U15434 (N_15434,N_10437,N_14303);
xor U15435 (N_15435,N_13877,N_10789);
xor U15436 (N_15436,N_13618,N_13122);
or U15437 (N_15437,N_12202,N_14766);
nand U15438 (N_15438,N_10449,N_12662);
nor U15439 (N_15439,N_10405,N_14199);
nand U15440 (N_15440,N_14842,N_13980);
nor U15441 (N_15441,N_14000,N_11012);
or U15442 (N_15442,N_10526,N_14172);
and U15443 (N_15443,N_10822,N_12904);
or U15444 (N_15444,N_14315,N_13032);
nand U15445 (N_15445,N_10556,N_13983);
nor U15446 (N_15446,N_13942,N_10518);
or U15447 (N_15447,N_11054,N_14636);
nor U15448 (N_15448,N_13948,N_14608);
and U15449 (N_15449,N_10630,N_14762);
or U15450 (N_15450,N_10703,N_10899);
nand U15451 (N_15451,N_10336,N_13768);
xnor U15452 (N_15452,N_11832,N_13421);
nor U15453 (N_15453,N_12445,N_13341);
nor U15454 (N_15454,N_12359,N_11332);
or U15455 (N_15455,N_12231,N_13533);
nand U15456 (N_15456,N_11768,N_12882);
nand U15457 (N_15457,N_14118,N_12111);
nand U15458 (N_15458,N_11354,N_10529);
nand U15459 (N_15459,N_12357,N_11103);
nor U15460 (N_15460,N_11461,N_10948);
nand U15461 (N_15461,N_13844,N_11380);
xnor U15462 (N_15462,N_12772,N_11415);
and U15463 (N_15463,N_12030,N_12692);
xor U15464 (N_15464,N_14574,N_12314);
and U15465 (N_15465,N_10629,N_12959);
nor U15466 (N_15466,N_11440,N_10411);
nand U15467 (N_15467,N_10992,N_13229);
nor U15468 (N_15468,N_10928,N_11665);
nand U15469 (N_15469,N_14057,N_10263);
nor U15470 (N_15470,N_11513,N_12900);
and U15471 (N_15471,N_14968,N_12503);
or U15472 (N_15472,N_10983,N_14223);
nor U15473 (N_15473,N_13212,N_13385);
and U15474 (N_15474,N_12802,N_11200);
xnor U15475 (N_15475,N_12748,N_13624);
nor U15476 (N_15476,N_14372,N_11930);
and U15477 (N_15477,N_10582,N_12997);
nand U15478 (N_15478,N_13767,N_14467);
nand U15479 (N_15479,N_12754,N_10961);
xor U15480 (N_15480,N_13933,N_13788);
or U15481 (N_15481,N_14412,N_14426);
nor U15482 (N_15482,N_13720,N_13445);
nand U15483 (N_15483,N_11363,N_12932);
and U15484 (N_15484,N_12743,N_10389);
nand U15485 (N_15485,N_14214,N_12309);
and U15486 (N_15486,N_10094,N_13168);
nand U15487 (N_15487,N_12943,N_11857);
or U15488 (N_15488,N_14417,N_13638);
nand U15489 (N_15489,N_14579,N_11427);
or U15490 (N_15490,N_14660,N_13440);
or U15491 (N_15491,N_12636,N_10250);
and U15492 (N_15492,N_11279,N_12406);
and U15493 (N_15493,N_13030,N_10434);
or U15494 (N_15494,N_13126,N_14811);
and U15495 (N_15495,N_10631,N_14942);
xor U15496 (N_15496,N_14858,N_14602);
nor U15497 (N_15497,N_13105,N_14272);
xor U15498 (N_15498,N_11974,N_14782);
nor U15499 (N_15499,N_12673,N_14550);
and U15500 (N_15500,N_11166,N_13107);
or U15501 (N_15501,N_11896,N_10726);
xor U15502 (N_15502,N_11299,N_11917);
or U15503 (N_15503,N_13378,N_14711);
nor U15504 (N_15504,N_12432,N_10342);
and U15505 (N_15505,N_12134,N_14254);
and U15506 (N_15506,N_11444,N_11241);
nand U15507 (N_15507,N_10107,N_12396);
nor U15508 (N_15508,N_12167,N_10312);
nand U15509 (N_15509,N_13860,N_13120);
or U15510 (N_15510,N_12035,N_10403);
nand U15511 (N_15511,N_10072,N_12779);
xor U15512 (N_15512,N_13648,N_12199);
xnor U15513 (N_15513,N_14327,N_10496);
and U15514 (N_15514,N_13494,N_11749);
nand U15515 (N_15515,N_11818,N_13088);
and U15516 (N_15516,N_11626,N_13721);
xnor U15517 (N_15517,N_14112,N_12388);
or U15518 (N_15518,N_11627,N_13437);
xnor U15519 (N_15519,N_14838,N_10724);
xnor U15520 (N_15520,N_13287,N_10004);
xor U15521 (N_15521,N_10374,N_14319);
or U15522 (N_15522,N_13221,N_13050);
and U15523 (N_15523,N_11102,N_14476);
and U15524 (N_15524,N_13832,N_13528);
and U15525 (N_15525,N_11631,N_10605);
or U15526 (N_15526,N_14664,N_10401);
xor U15527 (N_15527,N_14600,N_13871);
and U15528 (N_15528,N_14686,N_12974);
or U15529 (N_15529,N_11227,N_14804);
nor U15530 (N_15530,N_13370,N_14553);
and U15531 (N_15531,N_11005,N_11592);
nand U15532 (N_15532,N_11932,N_13694);
nor U15533 (N_15533,N_12384,N_10756);
and U15534 (N_15534,N_14943,N_14192);
and U15535 (N_15535,N_14643,N_12520);
nor U15536 (N_15536,N_14424,N_11771);
or U15537 (N_15537,N_12415,N_13556);
nand U15538 (N_15538,N_13987,N_11828);
and U15539 (N_15539,N_12089,N_13723);
and U15540 (N_15540,N_10563,N_12088);
nand U15541 (N_15541,N_10817,N_11445);
nand U15542 (N_15542,N_11021,N_11840);
nand U15543 (N_15543,N_13885,N_13399);
nor U15544 (N_15544,N_12527,N_13071);
nand U15545 (N_15545,N_14077,N_14495);
nand U15546 (N_15546,N_10000,N_10473);
nand U15547 (N_15547,N_11772,N_14735);
and U15548 (N_15548,N_10150,N_11993);
xnor U15549 (N_15549,N_10427,N_13295);
and U15550 (N_15550,N_12016,N_13289);
nand U15551 (N_15551,N_10573,N_11097);
or U15552 (N_15552,N_13944,N_14128);
xnor U15553 (N_15553,N_12027,N_13464);
xor U15554 (N_15554,N_11662,N_13203);
or U15555 (N_15555,N_11365,N_13292);
nand U15556 (N_15556,N_14710,N_14996);
xor U15557 (N_15557,N_10435,N_14419);
and U15558 (N_15558,N_12817,N_12484);
nand U15559 (N_15559,N_10558,N_10686);
nand U15560 (N_15560,N_12485,N_14806);
nand U15561 (N_15561,N_10721,N_11220);
nand U15562 (N_15562,N_12429,N_11677);
nor U15563 (N_15563,N_14753,N_13889);
nand U15564 (N_15564,N_12529,N_14817);
and U15565 (N_15565,N_14048,N_11537);
xor U15566 (N_15566,N_11386,N_10069);
and U15567 (N_15567,N_10050,N_14457);
nor U15568 (N_15568,N_11640,N_12991);
nor U15569 (N_15569,N_13675,N_13185);
nor U15570 (N_15570,N_10758,N_14836);
xnor U15571 (N_15571,N_12237,N_10658);
or U15572 (N_15572,N_14069,N_14225);
or U15573 (N_15573,N_12288,N_12587);
and U15574 (N_15574,N_12063,N_13750);
nand U15575 (N_15575,N_14999,N_14683);
xnor U15576 (N_15576,N_12155,N_14567);
and U15577 (N_15577,N_12737,N_10964);
nor U15578 (N_15578,N_10497,N_10295);
xnor U15579 (N_15579,N_11151,N_14322);
or U15580 (N_15580,N_10296,N_11557);
or U15581 (N_15581,N_14866,N_14777);
nor U15582 (N_15582,N_10788,N_10865);
nor U15583 (N_15583,N_11809,N_14377);
nor U15584 (N_15584,N_11510,N_14138);
nor U15585 (N_15585,N_10315,N_14939);
nor U15586 (N_15586,N_14482,N_11977);
or U15587 (N_15587,N_12490,N_13820);
nor U15588 (N_15588,N_12895,N_10262);
or U15589 (N_15589,N_10841,N_14580);
nand U15590 (N_15590,N_12880,N_12966);
nand U15591 (N_15591,N_12711,N_10681);
or U15592 (N_15592,N_13703,N_10578);
and U15593 (N_15593,N_14398,N_13899);
nor U15594 (N_15594,N_10001,N_14623);
xnor U15595 (N_15595,N_11281,N_10083);
and U15596 (N_15596,N_11464,N_10974);
nand U15597 (N_15597,N_14233,N_13135);
xnor U15598 (N_15598,N_12889,N_13409);
nand U15599 (N_15599,N_12908,N_13781);
nor U15600 (N_15600,N_10294,N_10441);
or U15601 (N_15601,N_10639,N_11147);
nor U15602 (N_15602,N_11244,N_12436);
xor U15603 (N_15603,N_14652,N_10386);
nor U15604 (N_15604,N_13291,N_10066);
nor U15605 (N_15605,N_14749,N_14674);
or U15606 (N_15606,N_11028,N_10291);
or U15607 (N_15607,N_12330,N_14468);
or U15608 (N_15608,N_11909,N_14774);
xor U15609 (N_15609,N_10796,N_10641);
or U15610 (N_15610,N_10198,N_12053);
nor U15611 (N_15611,N_11952,N_12393);
and U15612 (N_15612,N_12530,N_12084);
or U15613 (N_15613,N_10272,N_14281);
xor U15614 (N_15614,N_14611,N_11616);
nand U15615 (N_15615,N_10335,N_13148);
and U15616 (N_15616,N_13647,N_12060);
nor U15617 (N_15617,N_13237,N_13610);
and U15618 (N_15618,N_11957,N_14084);
nor U15619 (N_15619,N_10689,N_10638);
nand U15620 (N_15620,N_13875,N_11740);
xor U15621 (N_15621,N_11142,N_10171);
nand U15622 (N_15622,N_11697,N_13649);
and U15623 (N_15623,N_12348,N_10353);
nand U15624 (N_15624,N_14863,N_13645);
nor U15625 (N_15625,N_11216,N_11249);
nand U15626 (N_15626,N_10404,N_13777);
nor U15627 (N_15627,N_13920,N_10671);
nand U15628 (N_15628,N_12165,N_13414);
and U15629 (N_15629,N_14771,N_14271);
xor U15630 (N_15630,N_10384,N_10009);
and U15631 (N_15631,N_13572,N_14588);
or U15632 (N_15632,N_11248,N_12780);
nand U15633 (N_15633,N_12643,N_12472);
nand U15634 (N_15634,N_10808,N_13927);
xnor U15635 (N_15635,N_12710,N_10730);
nand U15636 (N_15636,N_11292,N_12469);
xor U15637 (N_15637,N_12785,N_11785);
or U15638 (N_15638,N_12507,N_13651);
xor U15639 (N_15639,N_12055,N_11393);
nor U15640 (N_15640,N_13738,N_14760);
or U15641 (N_15641,N_10835,N_12355);
and U15642 (N_15642,N_10901,N_13653);
nand U15643 (N_15643,N_13082,N_13201);
nor U15644 (N_15644,N_12728,N_14558);
xnor U15645 (N_15645,N_14291,N_10289);
xnor U15646 (N_15646,N_11990,N_13586);
xnor U15647 (N_15647,N_13209,N_12187);
xor U15648 (N_15648,N_14783,N_13206);
or U15649 (N_15649,N_14794,N_14116);
or U15650 (N_15650,N_13066,N_11434);
and U15651 (N_15651,N_13895,N_13748);
nand U15652 (N_15652,N_10318,N_14831);
xnor U15653 (N_15653,N_13846,N_10041);
nand U15654 (N_15654,N_13354,N_14758);
nor U15655 (N_15655,N_14085,N_11442);
nor U15656 (N_15656,N_10349,N_14024);
and U15657 (N_15657,N_13141,N_12660);
nand U15658 (N_15658,N_14599,N_14802);
and U15659 (N_15659,N_14539,N_12696);
nor U15660 (N_15660,N_13169,N_12020);
or U15661 (N_15661,N_11862,N_12552);
nor U15662 (N_15662,N_13432,N_13714);
and U15663 (N_15663,N_14736,N_13564);
or U15664 (N_15664,N_12979,N_12792);
nand U15665 (N_15665,N_10748,N_12149);
or U15666 (N_15666,N_11546,N_11198);
nand U15667 (N_15667,N_12727,N_14724);
and U15668 (N_15668,N_13069,N_12407);
nand U15669 (N_15669,N_12008,N_11121);
or U15670 (N_15670,N_12607,N_10690);
and U15671 (N_15671,N_10937,N_12534);
and U15672 (N_15672,N_14840,N_14815);
xor U15673 (N_15673,N_13799,N_12397);
nor U15674 (N_15674,N_10743,N_10846);
xnor U15675 (N_15675,N_14998,N_13394);
and U15676 (N_15676,N_13329,N_10472);
and U15677 (N_15677,N_13442,N_11176);
xnor U15678 (N_15678,N_13990,N_13363);
nor U15679 (N_15679,N_11019,N_12927);
nand U15680 (N_15680,N_13652,N_12455);
or U15681 (N_15681,N_14991,N_12985);
nor U15682 (N_15682,N_12277,N_11282);
xnor U15683 (N_15683,N_14381,N_13158);
or U15684 (N_15684,N_10185,N_14789);
and U15685 (N_15685,N_12319,N_12128);
and U15686 (N_15686,N_11723,N_10487);
or U15687 (N_15687,N_12820,N_10024);
nor U15688 (N_15688,N_13391,N_13166);
xor U15689 (N_15689,N_11673,N_10774);
and U15690 (N_15690,N_12698,N_11688);
xor U15691 (N_15691,N_10110,N_12765);
nand U15692 (N_15692,N_14160,N_14856);
nand U15693 (N_15693,N_14746,N_12594);
nor U15694 (N_15694,N_10546,N_13156);
or U15695 (N_15695,N_12164,N_14893);
xor U15696 (N_15696,N_13544,N_14235);
nand U15697 (N_15697,N_11650,N_11812);
nand U15698 (N_15698,N_12342,N_13065);
or U15699 (N_15699,N_11275,N_12890);
nand U15700 (N_15700,N_14564,N_10071);
and U15701 (N_15701,N_11615,N_12509);
or U15702 (N_15702,N_13909,N_12928);
xor U15703 (N_15703,N_12352,N_14504);
nand U15704 (N_15704,N_12590,N_11484);
nand U15705 (N_15705,N_13418,N_14368);
and U15706 (N_15706,N_11521,N_11905);
or U15707 (N_15707,N_11148,N_12510);
xor U15708 (N_15708,N_11997,N_14478);
xnor U15709 (N_15709,N_12331,N_13988);
nor U15710 (N_15710,N_14559,N_14635);
or U15711 (N_15711,N_10656,N_10057);
and U15712 (N_15712,N_14258,N_12395);
nand U15713 (N_15713,N_11973,N_11611);
and U15714 (N_15714,N_14289,N_10452);
nor U15715 (N_15715,N_13840,N_13401);
xnor U15716 (N_15716,N_13745,N_13130);
nand U15717 (N_15717,N_11480,N_10115);
or U15718 (N_15718,N_10303,N_13263);
or U15719 (N_15719,N_13372,N_13803);
or U15720 (N_15720,N_10597,N_13771);
nor U15721 (N_15721,N_13813,N_10868);
nand U15722 (N_15722,N_12648,N_10398);
nand U15723 (N_15723,N_11058,N_13594);
xor U15724 (N_15724,N_12272,N_13453);
xor U15725 (N_15725,N_13281,N_13412);
nand U15726 (N_15726,N_14292,N_12981);
nand U15727 (N_15727,N_13904,N_12885);
or U15728 (N_15728,N_11576,N_13796);
or U15729 (N_15729,N_11802,N_10421);
and U15730 (N_15730,N_13175,N_13426);
nand U15731 (N_15731,N_12580,N_12150);
nand U15732 (N_15732,N_12283,N_10931);
nor U15733 (N_15733,N_13688,N_13711);
and U15734 (N_15734,N_14298,N_11656);
nor U15735 (N_15735,N_10232,N_13562);
and U15736 (N_15736,N_11361,N_13474);
or U15737 (N_15737,N_12794,N_10371);
nand U15738 (N_15738,N_14884,N_13707);
xor U15739 (N_15739,N_12364,N_12433);
nand U15740 (N_15740,N_12465,N_13419);
xnor U15741 (N_15741,N_13226,N_12496);
xnor U15742 (N_15742,N_10453,N_12553);
and U15743 (N_15743,N_14788,N_13625);
xnor U15744 (N_15744,N_10306,N_13002);
xor U15745 (N_15745,N_11847,N_12706);
or U15746 (N_15746,N_11343,N_14224);
and U15747 (N_15747,N_10081,N_12980);
xor U15748 (N_15748,N_11482,N_14678);
and U15749 (N_15749,N_13753,N_12796);
nand U15750 (N_15750,N_12463,N_11871);
nand U15751 (N_15751,N_10048,N_11229);
nor U15752 (N_15752,N_11117,N_13697);
xor U15753 (N_15753,N_12440,N_10542);
or U15754 (N_15754,N_10030,N_10970);
or U15755 (N_15755,N_12756,N_10902);
nor U15756 (N_15756,N_11883,N_14101);
xor U15757 (N_15757,N_10583,N_13055);
nor U15758 (N_15758,N_14309,N_13754);
or U15759 (N_15759,N_10881,N_10814);
xnor U15760 (N_15760,N_12892,N_13874);
nor U15761 (N_15761,N_10572,N_11675);
or U15762 (N_15762,N_12419,N_14986);
xor U15763 (N_15763,N_12599,N_11319);
or U15764 (N_15764,N_10959,N_14284);
and U15765 (N_15765,N_11735,N_14072);
nand U15766 (N_15766,N_14929,N_10534);
or U15767 (N_15767,N_12191,N_12163);
nor U15768 (N_15768,N_12320,N_12075);
or U15769 (N_15769,N_13742,N_13233);
xor U15770 (N_15770,N_11101,N_12586);
nor U15771 (N_15771,N_10422,N_12421);
nor U15772 (N_15772,N_14728,N_12382);
xor U15773 (N_15773,N_13915,N_10194);
nand U15774 (N_15774,N_12201,N_14016);
nand U15775 (N_15775,N_11821,N_11250);
or U15776 (N_15776,N_14507,N_12541);
and U15777 (N_15777,N_12866,N_14052);
nand U15778 (N_15778,N_10191,N_11313);
and U15779 (N_15779,N_11720,N_13579);
nand U15780 (N_15780,N_14650,N_13823);
and U15781 (N_15781,N_13608,N_14930);
nand U15782 (N_15782,N_12098,N_11635);
xor U15783 (N_15783,N_10365,N_12834);
nand U15784 (N_15784,N_11348,N_12439);
or U15785 (N_15785,N_11617,N_10104);
xor U15786 (N_15786,N_10046,N_12921);
xnor U15787 (N_15787,N_12940,N_10754);
xnor U15788 (N_15788,N_13128,N_10577);
xor U15789 (N_15789,N_11106,N_13375);
and U15790 (N_15790,N_10770,N_12575);
xnor U15791 (N_15791,N_10381,N_13174);
nor U15792 (N_15792,N_12058,N_11781);
nand U15793 (N_15793,N_13805,N_12750);
xnor U15794 (N_15794,N_12853,N_10471);
nand U15795 (N_15795,N_14790,N_12069);
nand U15796 (N_15796,N_10922,N_10339);
and U15797 (N_15797,N_12971,N_10173);
and U15798 (N_15798,N_13316,N_12228);
xor U15799 (N_15799,N_12118,N_13376);
xor U15800 (N_15800,N_11588,N_11193);
and U15801 (N_15801,N_10202,N_11412);
and U15802 (N_15802,N_13943,N_12504);
or U15803 (N_15803,N_10917,N_13623);
and U15804 (N_15804,N_13670,N_13802);
or U15805 (N_15805,N_11352,N_13872);
nor U15806 (N_15806,N_13919,N_12274);
nor U15807 (N_15807,N_10151,N_12941);
nand U15808 (N_15808,N_13907,N_13546);
and U15809 (N_15809,N_12595,N_12596);
or U15810 (N_15810,N_13690,N_11409);
xor U15811 (N_15811,N_13137,N_13633);
or U15812 (N_15812,N_11877,N_14433);
xnor U15813 (N_15813,N_12947,N_10866);
xnor U15814 (N_15814,N_10912,N_12719);
nand U15815 (N_15815,N_10729,N_11946);
and U15816 (N_15816,N_11486,N_10746);
xor U15817 (N_15817,N_10372,N_14385);
nand U15818 (N_15818,N_11710,N_13319);
and U15819 (N_15819,N_13550,N_14537);
and U15820 (N_15820,N_12500,N_13780);
nand U15821 (N_15821,N_12234,N_14857);
or U15822 (N_15822,N_10673,N_14251);
nand U15823 (N_15823,N_12285,N_10128);
or U15824 (N_15824,N_14391,N_10815);
nand U15825 (N_15825,N_10239,N_13310);
nor U15826 (N_15826,N_11659,N_10604);
nor U15827 (N_15827,N_14593,N_10904);
or U15828 (N_15828,N_14522,N_10900);
xnor U15829 (N_15829,N_13124,N_11149);
xnor U15830 (N_15830,N_14250,N_10933);
and U15831 (N_15831,N_10585,N_11598);
or U15832 (N_15832,N_10982,N_13583);
and U15833 (N_15833,N_11983,N_10946);
nor U15834 (N_15834,N_12720,N_14713);
nand U15835 (N_15835,N_14355,N_13975);
xnor U15836 (N_15836,N_11839,N_14962);
xor U15837 (N_15837,N_10804,N_12192);
xor U15838 (N_15838,N_14141,N_13217);
or U15839 (N_15839,N_13797,N_11003);
xor U15840 (N_15840,N_11233,N_12258);
and U15841 (N_15841,N_14791,N_14243);
or U15842 (N_15842,N_13467,N_12403);
or U15843 (N_15843,N_12224,N_10618);
nand U15844 (N_15844,N_14239,N_14860);
nand U15845 (N_15845,N_13269,N_14427);
nand U15846 (N_15846,N_12856,N_13286);
nor U15847 (N_15847,N_14926,N_13972);
nor U15848 (N_15848,N_14524,N_14658);
nor U15849 (N_15849,N_13416,N_12919);
nor U15850 (N_15850,N_11715,N_10040);
and U15851 (N_15851,N_10192,N_12039);
or U15852 (N_15852,N_14252,N_11130);
nor U15853 (N_15853,N_14059,N_10149);
xor U15854 (N_15854,N_13616,N_14830);
xor U15855 (N_15855,N_14578,N_11196);
or U15856 (N_15856,N_13132,N_14152);
nor U15857 (N_15857,N_13379,N_11893);
xor U15858 (N_15858,N_12938,N_11456);
xnor U15859 (N_15859,N_13077,N_13381);
xnor U15860 (N_15860,N_13001,N_13746);
and U15861 (N_15861,N_12374,N_10839);
nor U15862 (N_15862,N_12605,N_13606);
nor U15863 (N_15863,N_14665,N_14019);
nor U15864 (N_15864,N_12934,N_13595);
and U15865 (N_15865,N_12615,N_12506);
xnor U15866 (N_15866,N_10244,N_10738);
or U15867 (N_15867,N_14676,N_12975);
nor U15868 (N_15868,N_12531,N_13253);
nor U15869 (N_15869,N_13730,N_13195);
nand U15870 (N_15870,N_10254,N_10633);
nand U15871 (N_15871,N_14397,N_13666);
xor U15872 (N_15872,N_10376,N_10782);
nand U15873 (N_15873,N_11110,N_13728);
and U15874 (N_15874,N_14220,N_10947);
nand U15875 (N_15875,N_14341,N_10739);
nand U15876 (N_15876,N_11554,N_12653);
nor U15877 (N_15877,N_14808,N_10616);
nand U15878 (N_15878,N_11563,N_13695);
or U15879 (N_15879,N_12333,N_13852);
xor U15880 (N_15880,N_14283,N_14867);
and U15881 (N_15881,N_12732,N_12935);
and U15882 (N_15882,N_13917,N_13794);
and U15883 (N_15883,N_11171,N_11387);
nor U15884 (N_15884,N_14921,N_12126);
and U15885 (N_15885,N_14849,N_13835);
and U15886 (N_15886,N_11815,N_12461);
xor U15887 (N_15887,N_13981,N_14185);
nor U15888 (N_15888,N_13747,N_11330);
nand U15889 (N_15889,N_12516,N_14245);
or U15890 (N_15890,N_10943,N_12729);
nor U15891 (N_15891,N_11453,N_11632);
nand U15892 (N_15892,N_10855,N_10380);
xor U15893 (N_15893,N_10571,N_14681);
and U15894 (N_15894,N_13541,N_13307);
or U15895 (N_15895,N_13145,N_10490);
or U15896 (N_15896,N_10319,N_13086);
nor U15897 (N_15897,N_10880,N_14380);
or U15898 (N_15898,N_13099,N_14670);
or U15899 (N_15899,N_13504,N_13516);
xnor U15900 (N_15900,N_10951,N_14852);
or U15901 (N_15901,N_13869,N_11071);
and U15902 (N_15902,N_10454,N_12473);
xnor U15903 (N_15903,N_13152,N_11133);
or U15904 (N_15904,N_11107,N_11706);
nor U15905 (N_15905,N_12874,N_10873);
nor U15906 (N_15906,N_10442,N_13734);
and U15907 (N_15907,N_12912,N_10020);
and U15908 (N_15908,N_14449,N_11305);
or U15909 (N_15909,N_13374,N_13926);
or U15910 (N_15910,N_11712,N_11967);
or U15911 (N_15911,N_14606,N_14503);
nor U15912 (N_15912,N_12086,N_10752);
xor U15913 (N_15913,N_13939,N_12865);
xnor U15914 (N_15914,N_14471,N_13716);
xor U15915 (N_15915,N_11257,N_14012);
nor U15916 (N_15916,N_11439,N_14657);
or U15917 (N_15917,N_14374,N_13165);
xor U15918 (N_15918,N_11013,N_11033);
nor U15919 (N_15919,N_13760,N_11503);
and U15920 (N_15920,N_13664,N_12219);
nand U15921 (N_15921,N_10736,N_14228);
and U15922 (N_15922,N_11559,N_11589);
nand U15923 (N_15923,N_11085,N_14304);
or U15924 (N_15924,N_13187,N_10395);
xnor U15925 (N_15925,N_13142,N_11105);
nand U15926 (N_15926,N_14518,N_10292);
nor U15927 (N_15927,N_13815,N_12172);
or U15928 (N_15928,N_11261,N_10074);
xor U15929 (N_15929,N_13219,N_11813);
and U15930 (N_15930,N_14055,N_12054);
nand U15931 (N_15931,N_11183,N_12062);
and U15932 (N_15932,N_10942,N_12153);
and U15933 (N_15933,N_14182,N_13810);
nand U15934 (N_15934,N_14556,N_10233);
and U15935 (N_15935,N_14064,N_10200);
xnor U15936 (N_15936,N_13323,N_13214);
nor U15937 (N_15937,N_10519,N_10735);
and U15938 (N_15938,N_13884,N_12993);
nor U15939 (N_15939,N_11654,N_14231);
nor U15940 (N_15940,N_11137,N_10230);
and U15941 (N_15941,N_12181,N_14088);
and U15942 (N_15942,N_10853,N_12216);
and U15943 (N_15943,N_10390,N_12511);
and U15944 (N_15944,N_13510,N_10476);
xor U15945 (N_15945,N_12428,N_13784);
or U15946 (N_15946,N_12113,N_12398);
nor U15947 (N_15947,N_14900,N_14561);
or U15948 (N_15948,N_13265,N_13656);
nand U15949 (N_15949,N_11205,N_13041);
xor U15950 (N_15950,N_11751,N_13581);
and U15951 (N_15951,N_10611,N_12992);
xnor U15952 (N_15952,N_10777,N_10973);
xnor U15953 (N_15953,N_14536,N_13338);
xnor U15954 (N_15954,N_14953,N_11256);
or U15955 (N_15955,N_12401,N_10803);
and U15956 (N_15956,N_13328,N_13170);
nor U15957 (N_15957,N_10521,N_13428);
or U15958 (N_15958,N_12246,N_11485);
nor U15959 (N_15959,N_12583,N_10366);
or U15960 (N_15960,N_12523,N_13344);
nor U15961 (N_15961,N_13911,N_13979);
xnor U15962 (N_15962,N_10759,N_13561);
nor U15963 (N_15963,N_12481,N_10361);
and U15964 (N_15964,N_10844,N_12044);
nand U15965 (N_15965,N_10326,N_13950);
or U15966 (N_15966,N_13893,N_14668);
nor U15967 (N_15967,N_13582,N_10477);
nand U15968 (N_15968,N_11081,N_10266);
or U15969 (N_15969,N_11944,N_14622);
nor U15970 (N_15970,N_11417,N_11786);
and U15971 (N_15971,N_10121,N_13842);
xor U15972 (N_15972,N_13814,N_12722);
and U15973 (N_15973,N_12801,N_10231);
nor U15974 (N_15974,N_10889,N_13045);
or U15975 (N_15975,N_14068,N_10801);
and U15976 (N_15976,N_11566,N_14948);
and U15977 (N_15977,N_13779,N_14697);
xor U15978 (N_15978,N_14193,N_14306);
nor U15979 (N_15979,N_10338,N_14441);
or U15980 (N_15980,N_13918,N_12863);
nor U15981 (N_15981,N_10968,N_11167);
nand U15982 (N_15982,N_14198,N_12712);
xor U15983 (N_15983,N_11320,N_11518);
nor U15984 (N_15984,N_12040,N_14074);
and U15985 (N_15985,N_13239,N_11392);
and U15986 (N_15986,N_12536,N_12296);
or U15987 (N_15987,N_12031,N_11032);
or U15988 (N_15988,N_11155,N_12899);
nand U15989 (N_15989,N_12253,N_11674);
and U15990 (N_15990,N_12758,N_13200);
nand U15991 (N_15991,N_12542,N_14940);
nor U15992 (N_15992,N_11996,N_10061);
xor U15993 (N_15993,N_14454,N_14257);
nor U15994 (N_15994,N_14111,N_11187);
xnor U15995 (N_15995,N_11394,N_11416);
nand U15996 (N_15996,N_13793,N_14335);
or U15997 (N_15997,N_12744,N_13584);
nand U15998 (N_15998,N_13896,N_12116);
nor U15999 (N_15999,N_10379,N_10209);
nand U16000 (N_16000,N_13811,N_11964);
and U16001 (N_16001,N_14267,N_14596);
or U16002 (N_16002,N_12132,N_10382);
nand U16003 (N_16003,N_13759,N_13816);
and U16004 (N_16004,N_13537,N_14646);
xor U16005 (N_16005,N_14626,N_12090);
xor U16006 (N_16006,N_10154,N_12579);
nand U16007 (N_16007,N_12731,N_13061);
xnor U16008 (N_16008,N_14378,N_11878);
nor U16009 (N_16009,N_13770,N_12259);
and U16010 (N_16010,N_13698,N_10364);
xnor U16011 (N_16011,N_11505,N_12891);
nor U16012 (N_16012,N_13912,N_10514);
xor U16013 (N_16013,N_14325,N_10457);
xor U16014 (N_16014,N_12613,N_11018);
or U16015 (N_16015,N_13257,N_10570);
nand U16016 (N_16016,N_14403,N_12078);
and U16017 (N_16017,N_11360,N_10082);
nor U16018 (N_16018,N_10934,N_11010);
nand U16019 (N_16019,N_10927,N_11134);
and U16020 (N_16020,N_14486,N_12842);
or U16021 (N_16021,N_11599,N_12194);
xnor U16022 (N_16022,N_11432,N_10623);
xnor U16023 (N_16023,N_11988,N_12738);
xnor U16024 (N_16024,N_11884,N_12423);
or U16025 (N_16025,N_10806,N_10495);
and U16026 (N_16026,N_14535,N_13410);
nor U16027 (N_16027,N_14918,N_11628);
nor U16028 (N_16028,N_12289,N_10503);
or U16029 (N_16029,N_13070,N_14897);
or U16030 (N_16030,N_14966,N_13881);
or U16031 (N_16031,N_14033,N_11315);
or U16032 (N_16032,N_12784,N_10464);
nor U16033 (N_16033,N_11514,N_10993);
nand U16034 (N_16034,N_12358,N_10400);
and U16035 (N_16035,N_13540,N_11825);
nor U16036 (N_16036,N_10888,N_12734);
nand U16037 (N_16037,N_14952,N_14912);
or U16038 (N_16038,N_14268,N_10876);
xor U16039 (N_16039,N_13735,N_10956);
nor U16040 (N_16040,N_10089,N_13431);
or U16041 (N_16041,N_11708,N_11752);
xnor U16042 (N_16042,N_10674,N_11914);
nor U16043 (N_16043,N_12386,N_13111);
nand U16044 (N_16044,N_13699,N_14754);
nor U16045 (N_16045,N_14151,N_13505);
or U16046 (N_16046,N_11441,N_14183);
nor U16047 (N_16047,N_11084,N_14028);
xnor U16048 (N_16048,N_13769,N_14078);
and U16049 (N_16049,N_12592,N_14569);
and U16050 (N_16050,N_11291,N_11001);
or U16051 (N_16051,N_11406,N_10599);
and U16052 (N_16052,N_11601,N_10553);
xnor U16053 (N_16053,N_14666,N_11845);
nand U16054 (N_16054,N_11120,N_11169);
nand U16055 (N_16055,N_12392,N_11578);
xnor U16056 (N_16056,N_14370,N_13617);
or U16057 (N_16057,N_10700,N_13262);
nor U16058 (N_16058,N_11494,N_10125);
and U16059 (N_16059,N_14508,N_11209);
xor U16060 (N_16060,N_12517,N_14684);
and U16061 (N_16061,N_11022,N_11808);
nor U16062 (N_16062,N_11246,N_14627);
nor U16063 (N_16063,N_13529,N_14576);
and U16064 (N_16064,N_14350,N_11678);
and U16065 (N_16065,N_14359,N_12742);
nor U16066 (N_16066,N_14447,N_14821);
and U16067 (N_16067,N_13136,N_11744);
nand U16068 (N_16068,N_13691,N_12242);
xor U16069 (N_16069,N_12148,N_14994);
nor U16070 (N_16070,N_10710,N_10042);
nand U16071 (N_16071,N_12543,N_12988);
nand U16072 (N_16072,N_10659,N_14469);
nor U16073 (N_16073,N_14642,N_11756);
nor U16074 (N_16074,N_13817,N_13549);
xnor U16075 (N_16075,N_10481,N_13756);
or U16076 (N_16076,N_14708,N_14527);
and U16077 (N_16077,N_14287,N_11185);
or U16078 (N_16078,N_14109,N_13577);
nor U16079 (N_16079,N_11575,N_12292);
or U16080 (N_16080,N_12810,N_10038);
xor U16081 (N_16081,N_14689,N_10885);
xnor U16082 (N_16082,N_11076,N_11962);
xnor U16083 (N_16083,N_10967,N_13971);
and U16084 (N_16084,N_13833,N_13600);
nand U16085 (N_16085,N_11247,N_13012);
and U16086 (N_16086,N_11263,N_13591);
or U16087 (N_16087,N_14835,N_12304);
or U16088 (N_16088,N_14259,N_11774);
and U16089 (N_16089,N_13782,N_13599);
nand U16090 (N_16090,N_12840,N_13484);
xor U16091 (N_16091,N_14551,N_11328);
nand U16092 (N_16092,N_12457,N_10562);
xnor U16093 (N_16093,N_11879,N_13236);
or U16094 (N_16094,N_14133,N_14818);
nor U16095 (N_16095,N_12002,N_11214);
xor U16096 (N_16096,N_11466,N_12026);
nand U16097 (N_16097,N_13283,N_14699);
or U16098 (N_16098,N_12028,N_10234);
or U16099 (N_16099,N_12180,N_14979);
or U16100 (N_16100,N_10509,N_13868);
or U16101 (N_16101,N_14737,N_10652);
and U16102 (N_16102,N_14389,N_10430);
or U16103 (N_16103,N_11410,N_13057);
and U16104 (N_16104,N_10424,N_14354);
nand U16105 (N_16105,N_12117,N_10994);
xor U16106 (N_16106,N_13427,N_12341);
or U16107 (N_16107,N_11239,N_14066);
or U16108 (N_16108,N_13138,N_10367);
nor U16109 (N_16109,N_13244,N_10698);
nor U16110 (N_16110,N_12955,N_13194);
nand U16111 (N_16111,N_14582,N_14560);
nor U16112 (N_16112,N_11283,N_13080);
nand U16113 (N_16113,N_12495,N_10035);
nand U16114 (N_16114,N_14734,N_10954);
nand U16115 (N_16115,N_13679,N_10494);
nor U16116 (N_16116,N_12210,N_14029);
or U16117 (N_16117,N_13151,N_11939);
nor U16118 (N_16118,N_12593,N_10636);
or U16119 (N_16119,N_10733,N_11419);
and U16120 (N_16120,N_12778,N_12824);
or U16121 (N_16121,N_14555,N_12373);
or U16122 (N_16122,N_11834,N_10725);
nor U16123 (N_16123,N_12826,N_12564);
and U16124 (N_16124,N_11730,N_11910);
nor U16125 (N_16125,N_11316,N_10377);
nor U16126 (N_16126,N_10143,N_10276);
or U16127 (N_16127,N_14134,N_13007);
nor U16128 (N_16128,N_14963,N_10845);
and U16129 (N_16129,N_14529,N_13190);
nand U16130 (N_16130,N_14757,N_13040);
and U16131 (N_16131,N_12871,N_10776);
and U16132 (N_16132,N_10106,N_12730);
nor U16133 (N_16133,N_10135,N_14989);
xor U16134 (N_16134,N_12620,N_12830);
or U16135 (N_16135,N_13524,N_10969);
nor U16136 (N_16136,N_13108,N_11273);
nand U16137 (N_16137,N_12379,N_12659);
nor U16138 (N_16138,N_14362,N_11660);
nand U16139 (N_16139,N_12647,N_13517);
nor U16140 (N_16140,N_10875,N_11865);
xnor U16141 (N_16141,N_13318,N_14744);
or U16142 (N_16142,N_10953,N_14351);
and U16143 (N_16143,N_12100,N_12482);
and U16144 (N_16144,N_12793,N_13408);
nand U16145 (N_16145,N_10773,N_11202);
nor U16146 (N_16146,N_12764,N_13074);
nor U16147 (N_16147,N_12193,N_11890);
or U16148 (N_16148,N_11345,N_10086);
nand U16149 (N_16149,N_12876,N_12639);
nand U16150 (N_16150,N_12581,N_12273);
nand U16151 (N_16151,N_12589,N_13435);
or U16152 (N_16152,N_12845,N_10480);
nor U16153 (N_16153,N_12602,N_13851);
and U16154 (N_16154,N_12822,N_12046);
xnor U16155 (N_16155,N_13332,N_13365);
or U16156 (N_16156,N_10590,N_14423);
xnor U16157 (N_16157,N_12145,N_13826);
or U16158 (N_16158,N_11079,N_10704);
and U16159 (N_16159,N_14144,N_11542);
or U16160 (N_16160,N_10099,N_14781);
nand U16161 (N_16161,N_11206,N_10840);
nor U16162 (N_16162,N_13087,N_14190);
or U16163 (N_16163,N_12263,N_10428);
or U16164 (N_16164,N_11995,N_10580);
xnor U16165 (N_16165,N_13924,N_10626);
or U16166 (N_16166,N_13668,N_14021);
xnor U16167 (N_16167,N_11297,N_14675);
and U16168 (N_16168,N_11655,N_14290);
and U16169 (N_16169,N_13383,N_14018);
or U16170 (N_16170,N_10134,N_10705);
nor U16171 (N_16171,N_12766,N_14647);
or U16172 (N_16172,N_12725,N_11255);
nor U16173 (N_16173,N_11344,N_13960);
or U16174 (N_16174,N_11063,N_12977);
or U16175 (N_16175,N_10120,N_11852);
nand U16176 (N_16176,N_13932,N_14104);
and U16177 (N_16177,N_12665,N_11817);
xnor U16178 (N_16178,N_14669,N_10105);
or U16179 (N_16179,N_10737,N_12232);
nor U16180 (N_16180,N_11116,N_14721);
or U16181 (N_16181,N_12501,N_13184);
nor U16182 (N_16182,N_10445,N_13211);
and U16183 (N_16183,N_10896,N_12011);
nor U16184 (N_16184,N_11716,N_10663);
xor U16185 (N_16185,N_10907,N_12811);
or U16186 (N_16186,N_11750,N_11414);
nor U16187 (N_16187,N_11679,N_14967);
and U16188 (N_16188,N_12603,N_12771);
or U16189 (N_16189,N_10544,N_12402);
nor U16190 (N_16190,N_11044,N_12072);
and U16191 (N_16191,N_13267,N_10145);
xor U16192 (N_16192,N_12843,N_14848);
nor U16193 (N_16193,N_10467,N_13891);
or U16194 (N_16194,N_11237,N_11629);
xnor U16195 (N_16195,N_10305,N_13325);
nor U16196 (N_16196,N_12850,N_10755);
xor U16197 (N_16197,N_12585,N_12411);
or U16198 (N_16198,N_12186,N_11057);
or U16199 (N_16199,N_14396,N_11866);
and U16200 (N_16200,N_11524,N_10745);
nor U16201 (N_16201,N_12617,N_13093);
or U16202 (N_16202,N_10170,N_14437);
nor U16203 (N_16203,N_12470,N_11156);
or U16204 (N_16204,N_13554,N_11581);
or U16205 (N_16205,N_11855,N_12179);
nor U16206 (N_16206,N_10559,N_10827);
nor U16207 (N_16207,N_11732,N_14236);
and U16208 (N_16208,N_10283,N_10634);
and U16209 (N_16209,N_14081,N_10279);
xor U16210 (N_16210,N_11797,N_13471);
or U16211 (N_16211,N_13496,N_10227);
nor U16212 (N_16212,N_13970,N_13812);
and U16213 (N_16213,N_12849,N_11558);
xor U16214 (N_16214,N_10019,N_12024);
or U16215 (N_16215,N_10127,N_11869);
and U16216 (N_16216,N_13740,N_10935);
xnor U16217 (N_16217,N_11014,N_13013);
nor U16218 (N_16218,N_13058,N_14045);
and U16219 (N_16219,N_14870,N_14516);
xnor U16220 (N_16220,N_13386,N_12431);
and U16221 (N_16221,N_13662,N_13521);
or U16222 (N_16222,N_10211,N_14407);
and U16223 (N_16223,N_13931,N_13005);
or U16224 (N_16224,N_12705,N_12915);
nor U16225 (N_16225,N_11048,N_13486);
nand U16226 (N_16226,N_14408,N_11355);
nand U16227 (N_16227,N_11916,N_13882);
nor U16228 (N_16228,N_12356,N_11684);
nor U16229 (N_16229,N_12265,N_13607);
nor U16230 (N_16230,N_10795,N_11560);
or U16231 (N_16231,N_11574,N_13901);
nor U16232 (N_16232,N_10201,N_12366);
or U16233 (N_16233,N_10650,N_14751);
or U16234 (N_16234,N_12573,N_12260);
nand U16235 (N_16235,N_12887,N_11763);
nand U16236 (N_16236,N_14187,N_13705);
and U16237 (N_16237,N_13527,N_10456);
nor U16238 (N_16238,N_10334,N_11082);
nand U16239 (N_16239,N_13587,N_10615);
and U16240 (N_16240,N_12654,N_11976);
nor U16241 (N_16241,N_12942,N_14461);
nand U16242 (N_16242,N_12036,N_14107);
and U16243 (N_16243,N_14591,N_11727);
nor U16244 (N_16244,N_11994,N_10651);
xnor U16245 (N_16245,N_13459,N_10627);
and U16246 (N_16246,N_10757,N_10984);
nor U16247 (N_16247,N_11759,N_10241);
and U16248 (N_16248,N_12322,N_10607);
nand U16249 (N_16249,N_11339,N_12416);
nand U16250 (N_16250,N_13403,N_12598);
nor U16251 (N_16251,N_14248,N_12519);
and U16252 (N_16252,N_13596,N_11334);
xor U16253 (N_16253,N_12125,N_12013);
and U16254 (N_16254,N_13348,N_12768);
or U16255 (N_16255,N_10543,N_10619);
nand U16256 (N_16256,N_14980,N_10182);
nand U16257 (N_16257,N_12033,N_12467);
and U16258 (N_16258,N_14043,N_10910);
nand U16259 (N_16259,N_13210,N_11424);
and U16260 (N_16260,N_14954,N_13159);
nor U16261 (N_16261,N_11608,N_12290);
nor U16262 (N_16262,N_11221,N_10594);
nand U16263 (N_16263,N_12311,N_13755);
nor U16264 (N_16264,N_11923,N_12057);
or U16265 (N_16265,N_13660,N_14820);
and U16266 (N_16266,N_13661,N_10655);
xnor U16267 (N_16267,N_14044,N_12316);
xor U16268 (N_16268,N_10952,N_14123);
nand U16269 (N_16269,N_11215,N_14273);
xor U16270 (N_16270,N_13273,N_14200);
xor U16271 (N_16271,N_12183,N_12499);
or U16272 (N_16272,N_13475,N_12960);
and U16273 (N_16273,N_13402,N_10179);
and U16274 (N_16274,N_11060,N_14988);
and U16275 (N_16275,N_13989,N_11580);
or U16276 (N_16276,N_11384,N_11168);
nand U16277 (N_16277,N_12034,N_10238);
nand U16278 (N_16278,N_12629,N_14584);
or U16279 (N_16279,N_11544,N_11856);
xor U16280 (N_16280,N_11940,N_13995);
nor U16281 (N_16281,N_12911,N_10561);
nor U16282 (N_16282,N_12211,N_11463);
nor U16283 (N_16283,N_13929,N_10793);
and U16284 (N_16284,N_13180,N_14106);
nor U16285 (N_16285,N_12805,N_11552);
and U16286 (N_16286,N_14993,N_12161);
nand U16287 (N_16287,N_10565,N_14905);
and U16288 (N_16288,N_13091,N_10848);
xnor U16289 (N_16289,N_10207,N_14170);
nor U16290 (N_16290,N_10146,N_12521);
xor U16291 (N_16291,N_11836,N_12513);
nand U16292 (N_16292,N_12739,N_11443);
nand U16293 (N_16293,N_13632,N_10052);
xor U16294 (N_16294,N_10797,N_13191);
nor U16295 (N_16295,N_13458,N_12497);
or U16296 (N_16296,N_13838,N_14361);
nand U16297 (N_16297,N_14654,N_14497);
or U16298 (N_16298,N_13857,N_12480);
nor U16299 (N_16299,N_13146,N_13825);
nand U16300 (N_16300,N_11745,N_10714);
nand U16301 (N_16301,N_13497,N_10741);
xor U16302 (N_16302,N_11481,N_13762);
or U16303 (N_16303,N_11296,N_10158);
or U16304 (N_16304,N_14100,N_12995);
or U16305 (N_16305,N_14923,N_11925);
and U16306 (N_16306,N_12550,N_14937);
and U16307 (N_16307,N_10268,N_10363);
or U16308 (N_16308,N_14071,N_12946);
xor U16309 (N_16309,N_12588,N_10084);
xor U16310 (N_16310,N_12674,N_13176);
xnor U16311 (N_16311,N_12235,N_14972);
nor U16312 (N_16312,N_14379,N_10394);
or U16313 (N_16313,N_12951,N_12858);
xor U16314 (N_16314,N_13461,N_11377);
nand U16315 (N_16315,N_13039,N_12569);
and U16316 (N_16316,N_14110,N_13598);
xnor U16317 (N_16317,N_11284,N_12656);
xnor U16318 (N_16318,N_13204,N_12671);
nand U16319 (N_16319,N_14733,N_11170);
nand U16320 (N_16320,N_11059,N_12868);
or U16321 (N_16321,N_11641,N_13117);
nor U16322 (N_16322,N_10533,N_10102);
xor U16323 (N_16323,N_11943,N_11605);
and U16324 (N_16324,N_13298,N_14568);
nand U16325 (N_16325,N_10720,N_14533);
and U16326 (N_16326,N_13991,N_11038);
nand U16327 (N_16327,N_10301,N_13240);
and U16328 (N_16328,N_13684,N_11490);
nand U16329 (N_16329,N_14121,N_13415);
or U16330 (N_16330,N_11367,N_12964);
nand U16331 (N_16331,N_12618,N_13515);
or U16332 (N_16332,N_10375,N_10811);
and U16333 (N_16333,N_12807,N_12256);
nand U16334 (N_16334,N_12483,N_13047);
or U16335 (N_16335,N_14034,N_14890);
nor U16336 (N_16336,N_14353,N_13243);
or U16337 (N_16337,N_12294,N_10608);
or U16338 (N_16338,N_12251,N_12790);
and U16339 (N_16339,N_11173,N_12442);
nor U16340 (N_16340,N_14997,N_14510);
and U16341 (N_16341,N_13270,N_10792);
nand U16342 (N_16342,N_10647,N_10694);
and U16343 (N_16343,N_10813,N_13199);
nor U16344 (N_16344,N_13859,N_14207);
xnor U16345 (N_16345,N_11496,N_12335);
nand U16346 (N_16346,N_14317,N_13850);
nor U16347 (N_16347,N_13552,N_12140);
nor U16348 (N_16348,N_12570,N_14162);
nor U16349 (N_16349,N_11956,N_10620);
or U16350 (N_16350,N_14079,N_10640);
and U16351 (N_16351,N_13985,N_14598);
nor U16352 (N_16352,N_12270,N_10786);
or U16353 (N_16353,N_13377,N_13388);
and U16354 (N_16354,N_11506,N_13787);
nor U16355 (N_16355,N_14429,N_11109);
and U16356 (N_16356,N_11499,N_10879);
and U16357 (N_16357,N_14435,N_10112);
nor U16358 (N_16358,N_13578,N_12759);
and U16359 (N_16359,N_12441,N_11065);
xor U16360 (N_16360,N_12206,N_14260);
xor U16361 (N_16361,N_14490,N_12957);
or U16362 (N_16362,N_12969,N_10347);
and U16363 (N_16363,N_13862,N_10248);
nor U16364 (N_16364,N_13076,N_11446);
nand U16365 (N_16365,N_11842,N_12323);
xnor U16366 (N_16366,N_14451,N_13171);
nor U16367 (N_16367,N_11922,N_11073);
and U16368 (N_16368,N_13639,N_11743);
xor U16369 (N_16369,N_14885,N_11371);
xnor U16370 (N_16370,N_10517,N_12225);
and U16371 (N_16371,N_11164,N_13024);
nand U16372 (N_16372,N_13352,N_14520);
and U16373 (N_16373,N_14465,N_11680);
nor U16374 (N_16374,N_10564,N_14701);
or U16375 (N_16375,N_11693,N_11887);
and U16376 (N_16376,N_10661,N_13509);
xnor U16377 (N_16377,N_11876,N_12494);
nor U16378 (N_16378,N_11400,N_13011);
and U16379 (N_16379,N_10524,N_11278);
or U16380 (N_16380,N_12948,N_14010);
nand U16381 (N_16381,N_13020,N_10220);
and U16382 (N_16382,N_12354,N_14075);
or U16383 (N_16383,N_11260,N_13371);
nand U16384 (N_16384,N_14745,N_12864);
xnor U16385 (N_16385,N_12435,N_12346);
nor U16386 (N_16386,N_11936,N_12142);
and U16387 (N_16387,N_12209,N_10834);
or U16388 (N_16388,N_10728,N_11304);
xnor U16389 (N_16389,N_14825,N_11179);
nor U16390 (N_16390,N_13133,N_14425);
nor U16391 (N_16391,N_14318,N_13094);
nor U16392 (N_16392,N_14784,N_14139);
xor U16393 (N_16393,N_10281,N_12688);
xnor U16394 (N_16394,N_11780,N_12317);
or U16395 (N_16395,N_11938,N_14047);
and U16396 (N_16396,N_13308,N_12103);
and U16397 (N_16397,N_13490,N_11197);
or U16398 (N_16398,N_11814,N_14557);
xor U16399 (N_16399,N_13547,N_14456);
nor U16400 (N_16400,N_14221,N_14690);
or U16401 (N_16401,N_13162,N_12627);
nor U16402 (N_16402,N_11099,N_12371);
or U16403 (N_16403,N_11880,N_12562);
and U16404 (N_16404,N_14410,N_11034);
nand U16405 (N_16405,N_10667,N_13489);
or U16406 (N_16406,N_12012,N_13276);
nor U16407 (N_16407,N_11398,N_10925);
xor U16408 (N_16408,N_12334,N_13451);
xnor U16409 (N_16409,N_11483,N_12079);
nor U16410 (N_16410,N_12687,N_13036);
xor U16411 (N_16411,N_12920,N_13808);
nor U16412 (N_16412,N_11672,N_14343);
xnor U16413 (N_16413,N_12836,N_13223);
nor U16414 (N_16414,N_13954,N_12308);
xor U16415 (N_16415,N_11201,N_11848);
or U16416 (N_16416,N_12217,N_12451);
nand U16417 (N_16417,N_14712,N_12869);
and U16418 (N_16418,N_13644,N_11041);
or U16419 (N_16419,N_14087,N_12096);
or U16420 (N_16420,N_10707,N_14716);
xor U16421 (N_16421,N_14910,N_14386);
nand U16422 (N_16422,N_14015,N_12684);
nor U16423 (N_16423,N_10406,N_12724);
nor U16424 (N_16424,N_10023,N_12677);
xnor U16425 (N_16425,N_12861,N_10172);
or U16426 (N_16426,N_10554,N_14945);
or U16427 (N_16427,N_14363,N_11982);
nand U16428 (N_16428,N_10256,N_12099);
xor U16429 (N_16429,N_10275,N_14286);
and U16430 (N_16430,N_12286,N_14801);
or U16431 (N_16431,N_12812,N_11585);
nand U16432 (N_16432,N_11603,N_13144);
or U16433 (N_16433,N_14947,N_10538);
and U16434 (N_16434,N_13062,N_14428);
or U16435 (N_16435,N_10137,N_10783);
or U16436 (N_16436,N_11864,N_13025);
nor U16437 (N_16437,N_13682,N_11043);
or U16438 (N_16438,N_12835,N_14229);
and U16439 (N_16439,N_11692,N_11378);
nor U16440 (N_16440,N_12414,N_10309);
xor U16441 (N_16441,N_11326,N_10576);
nand U16442 (N_16442,N_12591,N_12390);
or U16443 (N_16443,N_11612,N_11523);
xor U16444 (N_16444,N_14430,N_10802);
nor U16445 (N_16445,N_10987,N_12293);
and U16446 (N_16446,N_10502,N_11528);
and U16447 (N_16447,N_12806,N_14050);
nor U16448 (N_16448,N_10352,N_10157);
nand U16449 (N_16449,N_13127,N_12169);
nor U16450 (N_16450,N_12156,N_14610);
nor U16451 (N_16451,N_14934,N_12351);
nand U16452 (N_16452,N_10516,N_11823);
nand U16453 (N_16453,N_13790,N_12852);
nand U16454 (N_16454,N_10300,N_14779);
and U16455 (N_16455,N_11407,N_11491);
nand U16456 (N_16456,N_14179,N_10483);
nand U16457 (N_16457,N_13712,N_14276);
nand U16458 (N_16458,N_12297,N_13357);
xnor U16459 (N_16459,N_11534,N_14731);
or U16460 (N_16460,N_11162,N_11960);
or U16461 (N_16461,N_11699,N_10908);
nand U16462 (N_16462,N_11468,N_13634);
and U16463 (N_16463,N_10747,N_14003);
xnor U16464 (N_16464,N_11451,N_10978);
xor U16465 (N_16465,N_14709,N_14399);
and U16466 (N_16466,N_11383,N_11240);
xor U16467 (N_16467,N_14638,N_13230);
and U16468 (N_16468,N_13404,N_11987);
xnor U16469 (N_16469,N_14148,N_14528);
or U16470 (N_16470,N_13830,N_10059);
nor U16471 (N_16471,N_14816,N_13115);
nor U16472 (N_16472,N_13021,N_13064);
nand U16473 (N_16473,N_11532,N_12170);
or U16474 (N_16474,N_11096,N_14730);
or U16475 (N_16475,N_14843,N_13685);
or U16476 (N_16476,N_10333,N_10567);
nor U16477 (N_16477,N_14693,N_14127);
and U16478 (N_16478,N_11553,N_11844);
and U16479 (N_16479,N_13727,N_14519);
nor U16480 (N_16480,N_13103,N_14995);
and U16481 (N_16481,N_14961,N_12572);
xnor U16482 (N_16482,N_10419,N_14460);
nand U16483 (N_16483,N_13887,N_11379);
and U16484 (N_16484,N_10999,N_10070);
or U16485 (N_16485,N_12867,N_10265);
or U16486 (N_16486,N_12967,N_13134);
nor U16487 (N_16487,N_14755,N_14525);
nor U16488 (N_16488,N_10245,N_14748);
and U16489 (N_16489,N_10939,N_14859);
or U16490 (N_16490,N_10399,N_12902);
xnor U16491 (N_16491,N_14813,N_13302);
xor U16492 (N_16492,N_10140,N_11915);
or U16493 (N_16493,N_12717,N_12077);
and U16494 (N_16494,N_10971,N_14442);
nor U16495 (N_16495,N_11288,N_12220);
and U16496 (N_16496,N_12803,N_11066);
and U16497 (N_16497,N_14411,N_10433);
and U16498 (N_16498,N_12524,N_14090);
or U16499 (N_16499,N_10886,N_11796);
xnor U16500 (N_16500,N_11373,N_11437);
nor U16501 (N_16501,N_14395,N_11269);
nand U16502 (N_16502,N_14458,N_11321);
xnor U16503 (N_16503,N_12332,N_14436);
or U16504 (N_16504,N_13312,N_14862);
xor U16505 (N_16505,N_13282,N_13702);
or U16506 (N_16506,N_11487,N_12922);
nor U16507 (N_16507,N_12105,N_11891);
nor U16508 (N_16508,N_10210,N_12616);
or U16509 (N_16509,N_10643,N_12663);
nand U16510 (N_16510,N_13513,N_13015);
and U16511 (N_16511,N_13774,N_14203);
and U16512 (N_16512,N_12204,N_13536);
xnor U16513 (N_16513,N_13655,N_13454);
xnor U16514 (N_16514,N_10138,N_12689);
nor U16515 (N_16515,N_12123,N_14982);
or U16516 (N_16516,N_11569,N_12612);
and U16517 (N_16517,N_12137,N_14382);
or U16518 (N_16518,N_11177,N_13686);
nand U16519 (N_16519,N_11125,N_14499);
or U16520 (N_16520,N_11031,N_12773);
nand U16521 (N_16521,N_12886,N_11998);
and U16522 (N_16522,N_10549,N_11935);
or U16523 (N_16523,N_14445,N_10990);
and U16524 (N_16524,N_11767,N_14406);
nand U16525 (N_16525,N_11020,N_13905);
and U16526 (N_16526,N_13268,N_11157);
nor U16527 (N_16527,N_12196,N_13792);
or U16528 (N_16528,N_13722,N_13997);
nor U16529 (N_16529,N_14773,N_12362);
xnor U16530 (N_16530,N_13683,N_11902);
xor U16531 (N_16531,N_13073,N_10012);
and U16532 (N_16532,N_10903,N_10161);
and U16533 (N_16533,N_12502,N_14120);
nor U16534 (N_16534,N_14763,N_11165);
nand U16535 (N_16535,N_11289,N_13072);
and U16536 (N_16536,N_14810,N_14313);
and U16537 (N_16537,N_11947,N_13994);
nor U16538 (N_16538,N_12851,N_11999);
xnor U16539 (N_16539,N_13749,N_11143);
and U16540 (N_16540,N_14093,N_13834);
nor U16541 (N_16541,N_13879,N_13853);
nand U16542 (N_16542,N_13967,N_10540);
nand U16543 (N_16543,N_14908,N_11364);
nor U16544 (N_16544,N_13669,N_10139);
nand U16545 (N_16545,N_10224,N_14375);
nand U16546 (N_16546,N_13430,N_13389);
or U16547 (N_16547,N_11163,N_14196);
and U16548 (N_16548,N_10116,N_12367);
and U16549 (N_16549,N_12001,N_12361);
xor U16550 (N_16550,N_14970,N_13231);
nor U16551 (N_16551,N_11709,N_12048);
or U16552 (N_16552,N_13518,N_11093);
and U16553 (N_16553,N_13993,N_14484);
xor U16554 (N_16554,N_11969,N_10833);
nor U16555 (N_16555,N_11668,N_13928);
and U16556 (N_16556,N_10290,N_11810);
nand U16557 (N_16557,N_11069,N_12306);
xnor U16558 (N_16558,N_14358,N_12383);
and U16559 (N_16559,N_10257,N_11949);
or U16560 (N_16560,N_12236,N_10218);
xnor U16561 (N_16561,N_13752,N_11211);
and U16562 (N_16562,N_11545,N_14209);
and U16563 (N_16563,N_12474,N_13961);
or U16564 (N_16564,N_10331,N_11975);
nand U16565 (N_16565,N_10027,N_12709);
nor U16566 (N_16566,N_10492,N_11691);
nand U16567 (N_16567,N_11272,N_11570);
nand U16568 (N_16568,N_13075,N_11934);
nor U16569 (N_16569,N_13571,N_12144);
xnor U16570 (N_16570,N_12459,N_14928);
nor U16571 (N_16571,N_10123,N_12015);
nor U16572 (N_16572,N_10535,N_10545);
nand U16573 (N_16573,N_14202,N_10236);
nor U16574 (N_16574,N_11933,N_11517);
or U16575 (N_16575,N_10696,N_11644);
xor U16576 (N_16576,N_12207,N_13149);
or U16577 (N_16577,N_10579,N_14719);
nand U16578 (N_16578,N_13743,N_14360);
nand U16579 (N_16579,N_12245,N_14933);
and U16580 (N_16580,N_10259,N_14601);
and U16581 (N_16581,N_12408,N_14613);
and U16582 (N_16582,N_12038,N_12109);
or U16583 (N_16583,N_13968,N_11454);
nor U16584 (N_16584,N_11222,N_14091);
nor U16585 (N_16585,N_11927,N_13314);
and U16586 (N_16586,N_12832,N_10491);
nand U16587 (N_16587,N_11511,N_10142);
nor U16588 (N_16588,N_11501,N_12761);
nor U16589 (N_16589,N_10510,N_14570);
nor U16590 (N_16590,N_13609,N_11805);
xnor U16591 (N_16591,N_14595,N_13487);
and U16592 (N_16592,N_10877,N_11068);
or U16593 (N_16593,N_13916,N_11652);
nor U16594 (N_16594,N_14698,N_14274);
or U16595 (N_16595,N_12315,N_12901);
or U16596 (N_16596,N_12622,N_12321);
and U16597 (N_16597,N_11912,N_10838);
xnor U16598 (N_16598,N_14238,N_13465);
xor U16599 (N_16599,N_13614,N_13078);
nand U16600 (N_16600,N_12787,N_11872);
xor U16601 (N_16601,N_11906,N_10478);
xor U16602 (N_16602,N_13955,N_14031);
and U16603 (N_16603,N_10957,N_11590);
xnor U16604 (N_16604,N_11108,N_10592);
xnor U16605 (N_16605,N_14577,N_13551);
nor U16606 (N_16606,N_14394,N_13986);
and U16607 (N_16607,N_13186,N_11356);
or U16608 (N_16608,N_11850,N_10273);
xnor U16609 (N_16609,N_14927,N_12360);
and U16610 (N_16610,N_10393,N_13249);
nand U16611 (N_16611,N_13673,N_12338);
nor U16612 (N_16612,N_10551,N_10812);
and U16613 (N_16613,N_14124,N_10531);
nor U16614 (N_16614,N_10794,N_14300);
and U16615 (N_16615,N_11624,N_10356);
nand U16616 (N_16616,N_10932,N_14017);
or U16617 (N_16617,N_13396,N_10167);
nor U16618 (N_16618,N_13112,N_12449);
nor U16619 (N_16619,N_13324,N_13876);
or U16620 (N_16620,N_11742,N_11000);
or U16621 (N_16621,N_11488,N_12093);
nor U16622 (N_16622,N_14827,N_13343);
xnor U16623 (N_16623,N_12625,N_11498);
or U16624 (N_16624,N_12777,N_11024);
or U16625 (N_16625,N_14401,N_11803);
and U16626 (N_16626,N_12200,N_14131);
nand U16627 (N_16627,N_10625,N_12065);
nor U16628 (N_16628,N_14917,N_10818);
xnor U16629 (N_16629,N_10861,N_11667);
or U16630 (N_16630,N_11704,N_11985);
or U16631 (N_16631,N_12353,N_10340);
or U16632 (N_16632,N_12691,N_10949);
or U16633 (N_16633,N_13567,N_12645);
and U16634 (N_16634,N_14409,N_10426);
nor U16635 (N_16635,N_11374,N_12305);
nor U16636 (N_16636,N_14280,N_11049);
nand U16637 (N_16637,N_10085,N_11219);
xor U16638 (N_16638,N_10719,N_11489);
nand U16639 (N_16639,N_10450,N_12567);
nor U16640 (N_16640,N_10508,N_10155);
nand U16641 (N_16641,N_12047,N_13741);
and U16642 (N_16642,N_10486,N_12418);
nand U16643 (N_16643,N_13758,N_10215);
nand U16644 (N_16644,N_11889,N_14526);
or U16645 (N_16645,N_11556,N_14393);
xnor U16646 (N_16646,N_10287,N_10513);
nor U16647 (N_16647,N_14987,N_13824);
and U16648 (N_16648,N_11404,N_13717);
or U16649 (N_16649,N_11868,N_14255);
nor U16650 (N_16650,N_13890,N_13018);
xor U16651 (N_16651,N_12190,N_11495);
nand U16652 (N_16652,N_10017,N_14772);
nand U16653 (N_16653,N_13397,N_14614);
xor U16654 (N_16654,N_14137,N_13677);
or U16655 (N_16655,N_14919,N_14546);
or U16656 (N_16656,N_14544,N_10603);
or U16657 (N_16657,N_13102,N_10805);
xor U16658 (N_16658,N_13641,N_13183);
or U16659 (N_16659,N_12984,N_12059);
or U16660 (N_16660,N_10402,N_12635);
and U16661 (N_16661,N_12278,N_14227);
nand U16662 (N_16662,N_11141,N_14609);
or U16663 (N_16663,N_10882,N_13938);
or U16664 (N_16664,N_13864,N_11991);
and U16665 (N_16665,N_14803,N_10847);
and U16666 (N_16666,N_14924,N_11430);
or U16667 (N_16667,N_13613,N_12999);
nand U16668 (N_16668,N_12437,N_11375);
and U16669 (N_16669,N_12512,N_11403);
xor U16670 (N_16670,N_14950,N_11199);
xnor U16671 (N_16671,N_10852,N_13272);
and U16672 (N_16672,N_11854,N_14922);
and U16673 (N_16673,N_13010,N_14981);
nand U16674 (N_16674,N_13177,N_10664);
nand U16675 (N_16675,N_13161,N_12560);
and U16676 (N_16676,N_10261,N_10891);
nor U16677 (N_16677,N_13417,N_14971);
nor U16678 (N_16678,N_12666,N_11271);
and U16679 (N_16679,N_14880,N_12655);
nand U16680 (N_16680,N_11218,N_13023);
nor U16681 (N_16681,N_13678,N_10989);
xor U16682 (N_16682,N_12767,N_13258);
xor U16683 (N_16683,N_10034,N_14197);
and U16684 (N_16684,N_13865,N_13079);
nor U16685 (N_16685,N_11516,N_11118);
and U16686 (N_16686,N_11950,N_12690);
and U16687 (N_16687,N_12345,N_13737);
and U16688 (N_16688,N_11114,N_13477);
xor U16689 (N_16689,N_12091,N_11077);
or U16690 (N_16690,N_14833,N_13037);
and U16691 (N_16691,N_14883,N_11055);
and U16692 (N_16692,N_14008,N_10205);
and U16693 (N_16693,N_13153,N_11396);
nand U16694 (N_16694,N_12675,N_12789);
nand U16695 (N_16695,N_12646,N_13284);
or U16696 (N_16696,N_13260,N_12937);
xnor U16697 (N_16697,N_11100,N_10763);
and U16698 (N_16698,N_11607,N_10966);
or U16699 (N_16699,N_10063,N_13726);
nand U16700 (N_16700,N_12576,N_12548);
or U16701 (N_16701,N_12559,N_12010);
or U16702 (N_16702,N_10644,N_14305);
nand U16703 (N_16703,N_14891,N_12667);
nand U16704 (N_16704,N_12325,N_10391);
xor U16705 (N_16705,N_11182,N_14547);
and U16706 (N_16706,N_12037,N_10416);
or U16707 (N_16707,N_10388,N_14369);
xnor U16708 (N_16708,N_11042,N_14500);
xnor U16709 (N_16709,N_10918,N_12162);
and U16710 (N_16710,N_13369,N_13951);
nor U16711 (N_16711,N_10830,N_11178);
or U16712 (N_16712,N_12916,N_14215);
nor U16713 (N_16713,N_11098,N_14741);
nor U16714 (N_16714,N_11002,N_13252);
nor U16715 (N_16715,N_14607,N_13275);
nor U16716 (N_16716,N_14554,N_11806);
and U16717 (N_16717,N_14720,N_14333);
and U16718 (N_16718,N_14964,N_14899);
xor U16719 (N_16719,N_12007,N_13557);
nor U16720 (N_16720,N_13831,N_10392);
and U16721 (N_16721,N_13347,N_12400);
and U16722 (N_16722,N_12508,N_12872);
nor U16723 (N_16723,N_12715,N_10302);
or U16724 (N_16724,N_13090,N_14195);
xor U16725 (N_16725,N_14822,N_12854);
or U16726 (N_16726,N_10328,N_14056);
and U16727 (N_16727,N_10821,N_14054);
nor U16728 (N_16728,N_12823,N_12996);
xor U16729 (N_16729,N_12479,N_10032);
xnor U16730 (N_16730,N_12276,N_14634);
or U16731 (N_16731,N_12247,N_13619);
nand U16732 (N_16732,N_10829,N_10598);
or U16733 (N_16733,N_14740,N_10337);
or U16734 (N_16734,N_11801,N_14718);
or U16735 (N_16735,N_10602,N_10560);
and U16736 (N_16736,N_13801,N_13657);
and U16737 (N_16737,N_14722,N_14312);
nor U16738 (N_16738,N_12313,N_11408);
and U16739 (N_16739,N_10836,N_14388);
xor U16740 (N_16740,N_11661,N_12370);
and U16741 (N_16741,N_10168,N_11733);
or U16742 (N_16742,N_12944,N_13921);
nor U16743 (N_16743,N_14756,N_14020);
nor U16744 (N_16744,N_13098,N_14256);
nor U16745 (N_16745,N_13570,N_10462);
and U16746 (N_16746,N_12112,N_12695);
and U16747 (N_16747,N_13858,N_12781);
nand U16748 (N_16748,N_10614,N_12668);
or U16749 (N_16749,N_11718,N_12608);
and U16750 (N_16750,N_13309,N_10282);
nor U16751 (N_16751,N_12837,N_13631);
nand U16752 (N_16752,N_14892,N_11633);
nand U16753 (N_16753,N_14854,N_11719);
and U16754 (N_16754,N_14566,N_13940);
nor U16755 (N_16755,N_12676,N_14814);
xnor U16756 (N_16756,N_14513,N_11290);
nand U16757 (N_16757,N_12412,N_14142);
or U16758 (N_16758,N_13969,N_10362);
nor U16759 (N_16759,N_13367,N_10344);
nand U16760 (N_16760,N_11966,N_10387);
and U16761 (N_16761,N_12630,N_11707);
and U16762 (N_16762,N_10423,N_11242);
nor U16763 (N_16763,N_11037,N_12679);
xnor U16764 (N_16764,N_13555,N_14612);
and U16765 (N_16765,N_10332,N_11095);
or U16766 (N_16766,N_12269,N_14844);
xnor U16767 (N_16767,N_13667,N_10894);
nand U16768 (N_16768,N_14334,N_11789);
xor U16769 (N_16769,N_12422,N_12898);
or U16770 (N_16770,N_12107,N_12417);
nand U16771 (N_16771,N_12563,N_10680);
xnor U16772 (N_16772,N_10114,N_13097);
nor U16773 (N_16773,N_11112,N_11368);
and U16774 (N_16774,N_11984,N_13296);
xnor U16775 (N_16775,N_14775,N_12250);
or U16776 (N_16776,N_10446,N_10936);
or U16777 (N_16777,N_14237,N_11252);
nor U16778 (N_16778,N_11700,N_11450);
xor U16779 (N_16779,N_12240,N_14648);
or U16780 (N_16780,N_14649,N_11533);
and U16781 (N_16781,N_13393,N_11188);
or U16782 (N_16782,N_11203,N_12685);
nand U16783 (N_16783,N_14042,N_12244);
nand U16784 (N_16784,N_10769,N_13663);
nand U16785 (N_16785,N_11026,N_13492);
and U16786 (N_16786,N_10555,N_12337);
and U16787 (N_16787,N_11426,N_13046);
and U16788 (N_16788,N_10668,N_11285);
xnor U16789 (N_16789,N_10919,N_14103);
and U16790 (N_16790,N_13216,N_14729);
nand U16791 (N_16791,N_10410,N_12385);
and U16792 (N_16792,N_10056,N_14004);
or U16793 (N_16793,N_12298,N_11186);
and U16794 (N_16794,N_13847,N_12074);
nand U16795 (N_16795,N_13629,N_13903);
or U16796 (N_16796,N_13322,N_12986);
or U16797 (N_16797,N_12699,N_12525);
xnor U16798 (N_16798,N_14931,N_10646);
and U16799 (N_16799,N_13400,N_11747);
or U16800 (N_16800,N_10383,N_12229);
or U16801 (N_16801,N_11159,N_14130);
or U16802 (N_16802,N_14161,N_10550);
nand U16803 (N_16803,N_14135,N_13818);
and U16804 (N_16804,N_11402,N_10854);
nand U16805 (N_16805,N_12413,N_11471);
nor U16806 (N_16806,N_10960,N_11181);
xnor U16807 (N_16807,N_13976,N_14242);
or U16808 (N_16808,N_14797,N_13665);
nor U16809 (N_16809,N_11690,N_13914);
nor U16810 (N_16810,N_11310,N_11669);
and U16811 (N_16811,N_14189,N_13208);
and U16812 (N_16812,N_11094,N_11604);
or U16813 (N_16813,N_13202,N_12522);
xnor U16814 (N_16814,N_13068,N_12138);
nor U16815 (N_16815,N_11787,N_12638);
xor U16816 (N_16816,N_11232,N_11152);
and U16817 (N_16817,N_13406,N_13479);
and U16818 (N_16818,N_11194,N_14498);
and U16819 (N_16819,N_11139,N_12670);
or U16820 (N_16820,N_11230,N_14051);
nor U16821 (N_16821,N_11527,N_11507);
xnor U16822 (N_16822,N_10760,N_13878);
and U16823 (N_16823,N_14230,N_13553);
nand U16824 (N_16824,N_12857,N_12450);
nand U16825 (N_16825,N_10176,N_10648);
and U16826 (N_16826,N_14764,N_12816);
nand U16827 (N_16827,N_10475,N_12978);
nand U16828 (N_16828,N_10711,N_12073);
xnor U16829 (N_16829,N_13299,N_14073);
nor U16830 (N_16830,N_10699,N_13342);
or U16831 (N_16831,N_14673,N_13568);
xor U16832 (N_16832,N_14338,N_13251);
or U16833 (N_16833,N_13234,N_11382);
and U16834 (N_16834,N_11522,N_14879);
nand U16835 (N_16835,N_12279,N_11122);
nor U16836 (N_16836,N_14331,N_14889);
and U16837 (N_16837,N_11266,N_13315);
or U16838 (N_16838,N_11765,N_11924);
and U16839 (N_16839,N_12770,N_12681);
or U16840 (N_16840,N_13611,N_11792);
and U16841 (N_16841,N_13337,N_11072);
or U16842 (N_16842,N_10465,N_10451);
and U16843 (N_16843,N_13000,N_10775);
or U16844 (N_16844,N_14413,N_12102);
or U16845 (N_16845,N_14978,N_11175);
nor U16846 (N_16846,N_14349,N_14022);
xor U16847 (N_16847,N_13945,N_10622);
nor U16848 (N_16848,N_13883,N_14819);
nand U16849 (N_16849,N_11597,N_14965);
xnor U16850 (N_16850,N_11401,N_14615);
nand U16851 (N_16851,N_10915,N_10277);
and U16852 (N_16852,N_14070,N_10246);
nand U16853 (N_16853,N_10408,N_14246);
xor U16854 (N_16854,N_12983,N_14366);
xnor U16855 (N_16855,N_14462,N_13687);
nor U16856 (N_16856,N_14747,N_11989);
or U16857 (N_16857,N_14009,N_14545);
nor U16858 (N_16858,N_14829,N_12203);
or U16859 (N_16859,N_11388,N_11820);
nand U16860 (N_16860,N_11064,N_11929);
xnor U16861 (N_16861,N_13382,N_14113);
xor U16862 (N_16862,N_11119,N_14387);
nand U16863 (N_16863,N_13488,N_13026);
and U16864 (N_16864,N_11251,N_10298);
or U16865 (N_16865,N_10523,N_11653);
and U16866 (N_16866,N_14990,N_14875);
nand U16867 (N_16867,N_13558,N_13193);
xnor U16868 (N_16868,N_12218,N_11804);
and U16869 (N_16869,N_12873,N_13303);
and U16870 (N_16870,N_13143,N_11370);
or U16871 (N_16871,N_14959,N_13592);
or U16872 (N_16872,N_14957,N_10018);
xnor U16873 (N_16873,N_10712,N_13500);
and U16874 (N_16874,N_10468,N_14188);
and U16875 (N_16875,N_14247,N_12929);
xor U16876 (N_16876,N_11921,N_12121);
nor U16877 (N_16877,N_13129,N_14723);
and U16878 (N_16878,N_14096,N_13672);
nor U16879 (N_16879,N_11184,N_11425);
xor U16880 (N_16880,N_11029,N_10635);
nor U16881 (N_16881,N_13164,N_14473);
xor U16882 (N_16882,N_10870,N_11267);
nor U16883 (N_16883,N_11325,N_11366);
nor U16884 (N_16884,N_11849,N_12795);
nor U16885 (N_16885,N_12571,N_12716);
xnor U16886 (N_16886,N_12255,N_12949);
and U16887 (N_16887,N_14515,N_13671);
nand U16888 (N_16888,N_13084,N_13110);
and U16889 (N_16889,N_12774,N_10311);
nor U16890 (N_16890,N_11422,N_11595);
xnor U16891 (N_16891,N_14049,N_11009);
nor U16892 (N_16892,N_14914,N_10975);
and U16893 (N_16893,N_11670,N_11475);
xnor U16894 (N_16894,N_13476,N_13724);
nor U16895 (N_16895,N_13227,N_11734);
and U16896 (N_16896,N_14667,N_12686);
xnor U16897 (N_16897,N_11418,N_13446);
nand U16898 (N_16898,N_10432,N_13235);
and U16899 (N_16899,N_13650,N_14543);
nand U16900 (N_16900,N_13559,N_10466);
nor U16901 (N_16901,N_13327,N_14293);
nor U16902 (N_16902,N_11385,N_10058);
xnor U16903 (N_16903,N_10469,N_12998);
or U16904 (N_16904,N_12749,N_14108);
nand U16905 (N_16905,N_13081,N_12005);
xnor U16906 (N_16906,N_14316,N_10180);
nand U16907 (N_16907,N_14935,N_10213);
or U16908 (N_16908,N_12846,N_14253);
nand U16909 (N_16909,N_14275,N_10595);
and U16910 (N_16910,N_10022,N_10938);
or U16911 (N_16911,N_12003,N_12860);
or U16912 (N_16912,N_13854,N_13096);
nand U16913 (N_16913,N_13044,N_14985);
xor U16914 (N_16914,N_11705,N_10850);
nand U16915 (N_16915,N_14092,N_11739);
or U16916 (N_16916,N_11207,N_14594);
and U16917 (N_16917,N_14439,N_12328);
nor U16918 (N_16918,N_13978,N_14925);
xnor U16919 (N_16919,N_13575,N_11682);
xnor U16920 (N_16920,N_10716,N_13956);
and U16921 (N_16921,N_11980,N_11618);
or U16922 (N_16922,N_14302,N_13118);
xor U16923 (N_16923,N_10169,N_11195);
or U16924 (N_16924,N_11636,N_10274);
xnor U16925 (N_16925,N_14177,N_12394);
nand U16926 (N_16926,N_12299,N_14509);
xnor U16927 (N_16927,N_12434,N_11508);
nand U16928 (N_16928,N_12087,N_10314);
xnor U16929 (N_16929,N_12076,N_14390);
nand U16930 (N_16930,N_12471,N_11349);
nor U16931 (N_16931,N_13498,N_13713);
and U16932 (N_16932,N_13689,N_10766);
or U16933 (N_16933,N_12968,N_11234);
nor U16934 (N_16934,N_11602,N_10986);
and U16935 (N_16935,N_11853,N_10662);
nor U16936 (N_16936,N_13356,N_11799);
xor U16937 (N_16937,N_13085,N_14589);
and U16938 (N_16938,N_12018,N_10991);
nand U16939 (N_16939,N_10589,N_11276);
or U16940 (N_16940,N_11837,N_11591);
xnor U16941 (N_16941,N_10697,N_10368);
nand U16942 (N_16942,N_12953,N_13280);
nor U16943 (N_16943,N_10285,N_13574);
xnor U16944 (N_16944,N_11389,N_14902);
or U16945 (N_16945,N_12760,N_10762);
xnor U16946 (N_16946,N_11300,N_14006);
xor U16947 (N_16947,N_12641,N_13640);
nand U16948 (N_16948,N_12176,N_10178);
and U16949 (N_16949,N_13140,N_12844);
or U16950 (N_16950,N_14976,N_11885);
and U16951 (N_16951,N_12918,N_12025);
nand U16952 (N_16952,N_10260,N_10286);
and U16953 (N_16953,N_14038,N_12914);
or U16954 (N_16954,N_10790,N_11075);
xor U16955 (N_16955,N_11324,N_11754);
nor U16956 (N_16956,N_12307,N_13056);
nor U16957 (N_16957,N_14491,N_11124);
and U16958 (N_16958,N_14787,N_11277);
and U16959 (N_16959,N_10183,N_11583);
nand U16960 (N_16960,N_12151,N_14541);
and U16961 (N_16961,N_14265,N_12243);
or U16962 (N_16962,N_10924,N_10226);
xor U16963 (N_16963,N_13242,N_12152);
nor U16964 (N_16964,N_10596,N_13022);
nor U16965 (N_16965,N_11625,N_14630);
xnor U16966 (N_16966,N_14909,N_12578);
nand U16967 (N_16967,N_13218,N_10350);
nor U16968 (N_16968,N_12300,N_10077);
xor U16969 (N_16969,N_12664,N_10237);
xor U16970 (N_16970,N_14278,N_14974);
nor U16971 (N_16971,N_10515,N_12939);
or U16972 (N_16972,N_11753,N_12566);
or U16973 (N_16973,N_12070,N_11245);
nand U16974 (N_16974,N_10323,N_14548);
or U16975 (N_16975,N_13910,N_10036);
nand U16976 (N_16976,N_13321,N_10243);
nand U16977 (N_16977,N_12248,N_12466);
or U16978 (N_16978,N_13320,N_14656);
or U16979 (N_16979,N_12614,N_10479);
nor U16980 (N_16980,N_11819,N_13392);
nand U16981 (N_16981,N_12601,N_11050);
or U16982 (N_16982,N_13330,N_13264);
xor U16983 (N_16983,N_13147,N_13434);
nand U16984 (N_16984,N_14479,N_13207);
or U16985 (N_16985,N_10665,N_10505);
or U16986 (N_16986,N_14487,N_14738);
nand U16987 (N_16987,N_13491,N_14213);
xnor U16988 (N_16988,N_11062,N_12489);
nand U16989 (N_16989,N_14739,N_14443);
or U16990 (N_16990,N_11243,N_11362);
nor U16991 (N_16991,N_12831,N_11888);
nand U16992 (N_16992,N_11536,N_14640);
nand U16993 (N_16993,N_10184,N_11226);
xor U16994 (N_16994,N_13300,N_14855);
and U16995 (N_16995,N_13362,N_10727);
nand U16996 (N_16996,N_12584,N_11596);
and U16997 (N_16997,N_14920,N_14853);
xor U16998 (N_16998,N_11676,N_10065);
nand U16999 (N_16999,N_14098,N_12000);
nand U17000 (N_17000,N_13704,N_11728);
and U17001 (N_17001,N_12545,N_14903);
or U17002 (N_17002,N_11714,N_12909);
and U17003 (N_17003,N_10867,N_10051);
nor U17004 (N_17004,N_11770,N_14348);
nand U17005 (N_17005,N_13189,N_12378);
and U17006 (N_17006,N_11474,N_10568);
and U17007 (N_17007,N_13681,N_12954);
or U17008 (N_17008,N_10175,N_12577);
xnor U17009 (N_17009,N_14455,N_13067);
nor U17010 (N_17010,N_14356,N_13937);
nor U17011 (N_17011,N_11783,N_14572);
xor U17012 (N_17012,N_14563,N_11931);
nor U17013 (N_17013,N_13438,N_13407);
or U17014 (N_17014,N_10324,N_12114);
nor U17015 (N_17015,N_14973,N_13602);
and U17016 (N_17016,N_11035,N_14805);
nor U17017 (N_17017,N_13906,N_13063);
nand U17018 (N_17018,N_13181,N_12702);
nor U17019 (N_17019,N_12324,N_10837);
and U17020 (N_17020,N_14877,N_11467);
xnor U17021 (N_17021,N_13508,N_14422);
xor U17022 (N_17022,N_12427,N_11741);
nor U17023 (N_17023,N_11452,N_13197);
xnor U17024 (N_17024,N_14705,N_11811);
and U17025 (N_17025,N_10945,N_11210);
nand U17026 (N_17026,N_14173,N_10820);
nor U17027 (N_17027,N_12714,N_14617);
xor U17028 (N_17028,N_14944,N_14941);
or U17029 (N_17029,N_12409,N_13100);
xor U17030 (N_17030,N_14263,N_11689);
or U17031 (N_17031,N_10717,N_13452);
xnor U17032 (N_17032,N_10581,N_14167);
xor U17033 (N_17033,N_13952,N_11342);
and U17034 (N_17034,N_10348,N_10709);
nand U17035 (N_17035,N_11790,N_10217);
or U17036 (N_17036,N_10824,N_10117);
nor U17037 (N_17037,N_13121,N_11492);
or U17038 (N_17038,N_13659,N_13710);
nor U17039 (N_17039,N_11338,N_14261);
or U17040 (N_17040,N_10091,N_11683);
nor U17041 (N_17041,N_13693,N_12241);
nand U17042 (N_17042,N_14295,N_11761);
or U17043 (N_17043,N_12157,N_10944);
xnor U17044 (N_17044,N_11701,N_13898);
nor U17045 (N_17045,N_10965,N_12883);
nor U17046 (N_17046,N_14798,N_14715);
xor U17047 (N_17047,N_14204,N_13719);
and U17048 (N_17048,N_12982,N_14285);
nand U17049 (N_17049,N_12377,N_14328);
nor U17050 (N_17050,N_14800,N_11657);
nor U17051 (N_17051,N_14053,N_13470);
nand U17052 (N_17052,N_13220,N_10887);
and U17053 (N_17053,N_11841,N_14659);
xnor U17054 (N_17054,N_10463,N_11696);
xor U17055 (N_17055,N_14969,N_13353);
nand U17056 (N_17056,N_10823,N_11477);
xor U17057 (N_17057,N_13305,N_13278);
or U17058 (N_17058,N_11638,N_13506);
nor U17059 (N_17059,N_12208,N_14761);
and U17060 (N_17060,N_12556,N_10539);
nand U17061 (N_17061,N_11594,N_12281);
nand U17062 (N_17062,N_13241,N_13422);
and U17063 (N_17063,N_12649,N_11314);
and U17064 (N_17064,N_10995,N_11351);
nand U17065 (N_17065,N_11748,N_12693);
xor U17066 (N_17066,N_12697,N_14489);
and U17067 (N_17067,N_14094,N_13285);
nand U17068 (N_17068,N_11784,N_10610);
nand U17069 (N_17069,N_10188,N_10378);
nand U17070 (N_17070,N_14400,N_11535);
nand U17071 (N_17071,N_10679,N_13351);
nand U17072 (N_17072,N_10064,N_12799);
nand U17073 (N_17073,N_10098,N_14115);
or U17074 (N_17074,N_12119,N_10397);
and U17075 (N_17075,N_13482,N_11846);
xor U17076 (N_17076,N_10461,N_10229);
nor U17077 (N_17077,N_10653,N_12019);
or U17078 (N_17078,N_10702,N_10247);
nand U17079 (N_17079,N_13139,N_10187);
and U17080 (N_17080,N_13455,N_14240);
nor U17081 (N_17081,N_12405,N_12094);
or U17082 (N_17082,N_12129,N_13733);
nand U17083 (N_17083,N_13293,N_11901);
nand U17084 (N_17084,N_11270,N_10016);
and U17085 (N_17085,N_14218,N_14644);
nor U17086 (N_17086,N_13481,N_11007);
and U17087 (N_17087,N_14001,N_12994);
or U17088 (N_17088,N_12041,N_12184);
xnor U17089 (N_17089,N_11788,N_12757);
xor U17090 (N_17090,N_13589,N_12574);
and U17091 (N_17091,N_10458,N_14472);
or U17092 (N_17092,N_10541,N_10566);
nor U17093 (N_17093,N_13999,N_10025);
xor U17094 (N_17094,N_14839,N_10828);
or U17095 (N_17095,N_10761,N_12561);
nand U17096 (N_17096,N_10087,N_11217);
and U17097 (N_17097,N_12537,N_12032);
nor U17098 (N_17098,N_10147,N_12672);
nor U17099 (N_17099,N_12339,N_10791);
xor U17100 (N_17100,N_10152,N_10133);
xnor U17101 (N_17101,N_12349,N_10278);
nor U17102 (N_17102,N_12230,N_13855);
nor U17103 (N_17103,N_14618,N_10359);
nand U17104 (N_17104,N_12557,N_11336);
nor U17105 (N_17105,N_13643,N_10851);
and U17106 (N_17106,N_11564,N_11645);
nand U17107 (N_17107,N_13902,N_11548);
nor U17108 (N_17108,N_11965,N_14700);
nor U17109 (N_17109,N_11458,N_14895);
xor U17110 (N_17110,N_14841,N_13706);
xnor U17111 (N_17111,N_13154,N_12633);
xor U17112 (N_17112,N_10420,N_12262);
or U17113 (N_17113,N_14086,N_11843);
nand U17114 (N_17114,N_14651,N_10787);
xor U17115 (N_17115,N_14114,N_13051);
nand U17116 (N_17116,N_13054,N_13259);
xnor U17117 (N_17117,N_12755,N_11681);
xnor U17118 (N_17118,N_14501,N_14691);
and U17119 (N_17119,N_14208,N_11736);
nand U17120 (N_17120,N_14002,N_10160);
xnor U17121 (N_17121,N_14082,N_11762);
xnor U17122 (N_17122,N_13215,N_14332);
nor U17123 (N_17123,N_13949,N_12897);
nand U17124 (N_17124,N_11904,N_13775);
xnor U17125 (N_17125,N_12391,N_11520);
nor U17126 (N_17126,N_12930,N_11634);
nand U17127 (N_17127,N_14549,N_12067);
or U17128 (N_17128,N_13155,N_13736);
nor U17129 (N_17129,N_10642,N_14828);
or U17130 (N_17130,N_14211,N_14682);
xnor U17131 (N_17131,N_10307,N_10088);
nor U17132 (N_17132,N_10929,N_13279);
nor U17133 (N_17133,N_13306,N_12678);
xnor U17134 (N_17134,N_14882,N_13765);
nand U17135 (N_17135,N_12894,N_11959);
or U17136 (N_17136,N_10014,N_14060);
xor U17137 (N_17137,N_14026,N_11760);
or U17138 (N_17138,N_13288,N_14266);
and U17139 (N_17139,N_14262,N_11835);
or U17140 (N_17140,N_10443,N_13095);
and U17141 (N_17141,N_12626,N_14586);
or U17142 (N_17142,N_14888,N_14234);
xnor U17143 (N_17143,N_10628,N_11154);
nor U17144 (N_17144,N_14807,N_14653);
and U17145 (N_17145,N_10190,N_13941);
nor U17146 (N_17146,N_10609,N_13512);
and U17147 (N_17147,N_14448,N_13538);
nor U17148 (N_17148,N_12022,N_12438);
and U17149 (N_17149,N_11562,N_13052);
and U17150 (N_17150,N_14776,N_14680);
nand U17151 (N_17151,N_11036,N_10228);
nor U17152 (N_17152,N_11318,N_14706);
nand U17153 (N_17153,N_11882,N_11538);
xor U17154 (N_17154,N_14795,N_10977);
or U17155 (N_17155,N_10940,N_13615);
and U17156 (N_17156,N_12905,N_14326);
or U17157 (N_17157,N_11436,N_12547);
and U17158 (N_17158,N_13301,N_13622);
nor U17159 (N_17159,N_14505,N_11011);
or U17160 (N_17160,N_11870,N_14324);
nor U17161 (N_17161,N_10444,N_12862);
nand U17162 (N_17162,N_14076,N_10223);
or U17163 (N_17163,N_10415,N_14605);
nor U17164 (N_17164,N_10921,N_11136);
nor U17165 (N_17165,N_14145,N_13700);
nor U17166 (N_17166,N_10677,N_11881);
nand U17167 (N_17167,N_10547,N_13772);
and U17168 (N_17168,N_13807,N_10431);
or U17169 (N_17169,N_13261,N_14154);
and U17170 (N_17170,N_10373,N_14796);
or U17171 (N_17171,N_13423,N_11223);
xor U17172 (N_17172,N_13019,N_14799);
or U17173 (N_17173,N_10369,N_13125);
xnor U17174 (N_17174,N_10100,N_11540);
or U17175 (N_17175,N_12487,N_14450);
xnor U17176 (N_17176,N_13766,N_13880);
and U17177 (N_17177,N_13998,N_10552);
and U17178 (N_17178,N_14164,N_11777);
or U17179 (N_17179,N_10520,N_11004);
and U17180 (N_17180,N_11298,N_13450);
or U17181 (N_17181,N_11067,N_12736);
nor U17182 (N_17182,N_13473,N_12925);
and U17183 (N_17183,N_10493,N_12533);
xnor U17184 (N_17184,N_12131,N_12600);
nand U17185 (N_17185,N_10251,N_12376);
and U17186 (N_17186,N_12652,N_12050);
nor U17187 (N_17187,N_11926,N_10507);
or U17188 (N_17188,N_11264,N_11895);
nor U17189 (N_17189,N_12380,N_14573);
xor U17190 (N_17190,N_13114,N_12267);
and U17191 (N_17191,N_13958,N_10208);
xor U17192 (N_17192,N_10849,N_10109);
or U17193 (N_17193,N_13696,N_14886);
xnor U17194 (N_17194,N_14308,N_14431);
or U17195 (N_17195,N_11593,N_10666);
xnor U17196 (N_17196,N_12213,N_12097);
and U17197 (N_17197,N_13588,N_10731);
nor U17198 (N_17198,N_10996,N_10079);
and U17199 (N_17199,N_11978,N_11713);
and U17200 (N_17200,N_10732,N_13345);
nor U17201 (N_17201,N_13501,N_14117);
or U17202 (N_17202,N_13395,N_13560);
xnor U17203 (N_17203,N_13466,N_14163);
or U17204 (N_17204,N_12326,N_13004);
or U17205 (N_17205,N_12006,N_10780);
nand U17206 (N_17206,N_14703,N_10299);
and U17207 (N_17207,N_10448,N_10649);
or U17208 (N_17208,N_13761,N_14420);
nor U17209 (N_17209,N_13358,N_11140);
nor U17210 (N_17210,N_13059,N_10033);
xnor U17211 (N_17211,N_13478,N_10981);
xnor U17212 (N_17212,N_11903,N_12185);
xnor U17213 (N_17213,N_11702,N_12426);
nand U17214 (N_17214,N_11549,N_14383);
or U17215 (N_17215,N_12368,N_10003);
nor U17216 (N_17216,N_13795,N_12788);
nand U17217 (N_17217,N_11937,N_14896);
and U17218 (N_17218,N_13965,N_13894);
and U17219 (N_17219,N_10784,N_12410);
nand U17220 (N_17220,N_11431,N_10413);
xor U17221 (N_17221,N_14847,N_13380);
and U17222 (N_17222,N_10219,N_14219);
nand U17223 (N_17223,N_14655,N_13626);
nand U17224 (N_17224,N_10857,N_11698);
nand U17225 (N_17225,N_13150,N_13888);
and U17226 (N_17226,N_12301,N_10914);
xor U17227 (N_17227,N_10153,N_14850);
nor U17228 (N_17228,N_10235,N_10687);
and U17229 (N_17229,N_12558,N_10204);
or U17230 (N_17230,N_14984,N_10692);
and U17231 (N_17231,N_13360,N_12239);
and U17232 (N_17232,N_10859,N_12680);
xor U17233 (N_17233,N_14083,N_12813);
nor U17234 (N_17234,N_11948,N_12425);
xor U17235 (N_17235,N_13225,N_13346);
nor U17236 (N_17236,N_12080,N_14336);
or U17237 (N_17237,N_11666,N_14632);
nor U17238 (N_17238,N_11519,N_10688);
nand U17239 (N_17239,N_13773,N_10011);
nor U17240 (N_17240,N_14344,N_11630);
xor U17241 (N_17241,N_10874,N_13304);
nand U17242 (N_17242,N_13565,N_14604);
and U17243 (N_17243,N_12085,N_10988);
and U17244 (N_17244,N_13449,N_14514);
nand U17245 (N_17245,N_10144,N_10329);
or U17246 (N_17246,N_12628,N_12021);
nor U17247 (N_17247,N_12769,N_12514);
xor U17248 (N_17248,N_10869,N_14129);
nand U17249 (N_17249,N_10740,N_10591);
nand U17250 (N_17250,N_13192,N_12877);
nand U17251 (N_17251,N_14661,N_14310);
xor U17252 (N_17252,N_12791,N_10321);
xnor U17253 (N_17253,N_14014,N_14687);
or U17254 (N_17254,N_13612,N_11807);
or U17255 (N_17255,N_12486,N_11204);
nand U17256 (N_17256,N_11346,N_13936);
and U17257 (N_17257,N_14342,N_13535);
and U17258 (N_17258,N_12538,N_14194);
or U17259 (N_17259,N_13049,N_10670);
nor U17260 (N_17260,N_11826,N_10264);
and U17261 (N_17261,N_13167,N_13472);
xnor U17262 (N_17262,N_13313,N_14373);
and U17263 (N_17263,N_12958,N_11579);
nand U17264 (N_17264,N_10511,N_11420);
xnor U17265 (N_17265,N_10825,N_13900);
and U17266 (N_17266,N_14785,N_11725);
xnor U17267 (N_17267,N_14102,N_10459);
and U17268 (N_17268,N_11293,N_14834);
xnor U17269 (N_17269,N_10129,N_12303);
and U17270 (N_17270,N_11722,N_10212);
nand U17271 (N_17271,N_14873,N_10482);
nor U17272 (N_17272,N_13590,N_12906);
and U17273 (N_17273,N_11968,N_12546);
nand U17274 (N_17274,N_14155,N_11253);
and U17275 (N_17275,N_14977,N_10488);
nand U17276 (N_17276,N_10897,N_11372);
or U17277 (N_17277,N_12365,N_11435);
xnor U17278 (N_17278,N_14184,N_12174);
nand U17279 (N_17279,N_13963,N_12460);
nor U17280 (N_17280,N_14105,N_10101);
nand U17281 (N_17281,N_14759,N_10258);
nor U17282 (N_17282,N_10313,N_12535);
and U17283 (N_17283,N_10045,N_14792);
and U17284 (N_17284,N_11144,N_11129);
xnor U17285 (N_17285,N_14030,N_11350);
nor U17286 (N_17286,N_10080,N_12302);
and U17287 (N_17287,N_10267,N_12009);
or U17288 (N_17288,N_13060,N_14232);
and U17289 (N_17289,N_11138,N_12454);
nand U17290 (N_17290,N_11457,N_11899);
xnor U17291 (N_17291,N_11971,N_11550);
nor U17292 (N_17292,N_13456,N_12609);
nor U17293 (N_17293,N_13725,N_14726);
and U17294 (N_17294,N_10693,N_10672);
xnor U17295 (N_17295,N_14321,N_13413);
nand U17296 (N_17296,N_11302,N_11609);
and U17297 (N_17297,N_13828,N_12205);
nor U17298 (N_17298,N_14837,N_12782);
nor U17299 (N_17299,N_13034,N_10407);
nand U17300 (N_17300,N_14475,N_12952);
nor U17301 (N_17301,N_11497,N_14470);
and U17302 (N_17302,N_11778,N_11213);
xnor U17303 (N_17303,N_10044,N_11341);
nand U17304 (N_17304,N_10864,N_12284);
xnor U17305 (N_17305,N_12493,N_13922);
nand U17306 (N_17306,N_14581,N_10118);
nor U17307 (N_17307,N_14936,N_14046);
nand U17308 (N_17308,N_13361,N_12017);
nor U17309 (N_17309,N_12965,N_14279);
and U17310 (N_17310,N_12147,N_12973);
nor U17311 (N_17311,N_14696,N_10130);
nor U17312 (N_17312,N_14992,N_10111);
or U17313 (N_17313,N_10005,N_12127);
nand U17314 (N_17314,N_11047,N_13106);
or U17315 (N_17315,N_11172,N_12540);
nor U17316 (N_17316,N_11928,N_12819);
xnor U17317 (N_17317,N_11478,N_11329);
nor U17318 (N_17318,N_10136,N_13179);
nand U17319 (N_17319,N_12917,N_12669);
nor U17320 (N_17320,N_10308,N_10316);
nor U17321 (N_17321,N_11620,N_10528);
or U17322 (N_17322,N_11908,N_13982);
nor U17323 (N_17323,N_12029,N_11874);
or U17324 (N_17324,N_14906,N_11078);
nand U17325 (N_17325,N_11150,N_10979);
and U17326 (N_17326,N_12014,N_14679);
nand U17327 (N_17327,N_13009,N_13776);
nor U17328 (N_17328,N_14037,N_13433);
and U17329 (N_17329,N_14205,N_13809);
nor U17330 (N_17330,N_10779,N_12052);
or U17331 (N_17331,N_10765,N_12878);
xnor U17332 (N_17332,N_13255,N_11555);
nand U17333 (N_17333,N_14769,N_14346);
and U17334 (N_17334,N_10997,N_10963);
and U17335 (N_17335,N_14768,N_12950);
and U17336 (N_17336,N_14872,N_14149);
and U17337 (N_17337,N_14975,N_12723);
or U17338 (N_17338,N_13266,N_12476);
and U17339 (N_17339,N_10624,N_13837);
or U17340 (N_17340,N_12064,N_11875);
and U17341 (N_17341,N_12657,N_10637);
and U17342 (N_17342,N_13340,N_14714);
and U17343 (N_17343,N_12043,N_13297);
nor U17344 (N_17344,N_12700,N_10500);
nor U17345 (N_17345,N_10858,N_11335);
or U17346 (N_17346,N_10645,N_14371);
and U17347 (N_17347,N_11161,N_12651);
xnor U17348 (N_17348,N_10043,N_10593);
nor U17349 (N_17349,N_13718,N_13238);
or U17350 (N_17350,N_12444,N_11561);
nor U17351 (N_17351,N_13841,N_14511);
xor U17352 (N_17352,N_11970,N_12783);
and U17353 (N_17353,N_14901,N_10186);
and U17354 (N_17354,N_12175,N_12606);
xor U17355 (N_17355,N_11729,N_10798);
nand U17356 (N_17356,N_13839,N_11411);
nor U17357 (N_17357,N_11053,N_14132);
and U17358 (N_17358,N_14955,N_14210);
or U17359 (N_17359,N_14639,N_11863);
and U17360 (N_17360,N_14823,N_14628);
nor U17361 (N_17361,N_12420,N_12726);
and U17362 (N_17362,N_14904,N_14174);
and U17363 (N_17363,N_14695,N_11238);
xnor U17364 (N_17364,N_10506,N_14347);
nand U17365 (N_17365,N_14036,N_10007);
nand U17366 (N_17366,N_13569,N_12389);
nand U17367 (N_17367,N_14672,N_11027);
xnor U17368 (N_17368,N_14217,N_13946);
nor U17369 (N_17369,N_11087,N_14150);
nor U17370 (N_17370,N_12896,N_14099);
and U17371 (N_17371,N_10962,N_14898);
or U17372 (N_17372,N_11113,N_13398);
and U17373 (N_17373,N_10816,N_11160);
xnor U17374 (N_17374,N_14168,N_13387);
nor U17375 (N_17375,N_11838,N_12133);
xor U17376 (N_17376,N_11951,N_10355);
or U17377 (N_17377,N_12989,N_11613);
nor U17378 (N_17378,N_13892,N_14688);
nand U17379 (N_17379,N_12923,N_11301);
xor U17380 (N_17380,N_14365,N_10310);
or U17381 (N_17381,N_13654,N_11829);
nor U17382 (N_17382,N_12642,N_13757);
nand U17383 (N_17383,N_11963,N_11541);
and U17384 (N_17384,N_13469,N_12815);
or U17385 (N_17385,N_13873,N_11831);
and U17386 (N_17386,N_14067,N_12252);
or U17387 (N_17387,N_13274,N_14206);
or U17388 (N_17388,N_10742,N_13984);
and U17389 (N_17389,N_11955,N_14907);
and U17390 (N_17390,N_12775,N_14007);
and U17391 (N_17391,N_14865,N_10683);
or U17392 (N_17392,N_10354,N_14474);
xnor U17393 (N_17393,N_11390,N_10039);
and U17394 (N_17394,N_11526,N_12747);
and U17395 (N_17395,N_13934,N_12226);
xnor U17396 (N_17396,N_14122,N_13172);
nand U17397 (N_17397,N_14384,N_10166);
nand U17398 (N_17398,N_13457,N_13739);
and U17399 (N_17399,N_10778,N_12800);
and U17400 (N_17400,N_13786,N_13420);
xor U17401 (N_17401,N_11500,N_13806);
nand U17402 (N_17402,N_12233,N_13173);
xnor U17403 (N_17403,N_11726,N_13163);
xor U17404 (N_17404,N_11647,N_12551);
and U17405 (N_17405,N_14485,N_14340);
nand U17406 (N_17406,N_13443,N_11191);
or U17407 (N_17407,N_12215,N_10221);
nor U17408 (N_17408,N_14080,N_10905);
nand U17409 (N_17409,N_14005,N_10718);
or U17410 (N_17410,N_14040,N_14477);
or U17411 (N_17411,N_10678,N_10006);
or U17412 (N_17412,N_13048,N_10015);
nand U17413 (N_17413,N_11898,N_10675);
xor U17414 (N_17414,N_12597,N_11231);
xnor U17415 (N_17415,N_12254,N_11438);
and U17416 (N_17416,N_14434,N_11280);
or U17417 (N_17417,N_12718,N_11030);
or U17418 (N_17418,N_11462,N_11294);
nand U17419 (N_17419,N_14809,N_10976);
nand U17420 (N_17420,N_13731,N_11340);
nor U17421 (N_17421,N_12447,N_12261);
nand U17422 (N_17422,N_10177,N_10189);
xor U17423 (N_17423,N_10113,N_10037);
or U17424 (N_17424,N_10955,N_13008);
nor U17425 (N_17425,N_12619,N_10078);
xnor U17426 (N_17426,N_11132,N_10842);
nand U17427 (N_17427,N_12280,N_14742);
nor U17428 (N_17428,N_11127,N_13424);
and U17429 (N_17429,N_10253,N_13493);
xor U17430 (N_17430,N_10601,N_13715);
nand U17431 (N_17431,N_11395,N_14296);
nor U17432 (N_17432,N_11286,N_13256);
and U17433 (N_17433,N_14530,N_12555);
xnor U17434 (N_17434,N_10906,N_12707);
or U17435 (N_17435,N_11694,N_11867);
and U17436 (N_17436,N_13254,N_12544);
nand U17437 (N_17437,N_13366,N_13604);
and U17438 (N_17438,N_14851,N_11023);
and U17439 (N_17439,N_11515,N_13355);
nor U17440 (N_17440,N_12291,N_10013);
nand U17441 (N_17441,N_10438,N_11421);
and U17442 (N_17442,N_10501,N_13597);
or U17443 (N_17443,N_13335,N_12745);
nor U17444 (N_17444,N_13205,N_12120);
xnor U17445 (N_17445,N_14095,N_13764);
nand U17446 (N_17446,N_14270,N_10096);
xor U17447 (N_17447,N_11685,N_10418);
or U17448 (N_17448,N_13621,N_11128);
xnor U17449 (N_17449,N_12658,N_10455);
nor U17450 (N_17450,N_14671,N_13502);
nor U17451 (N_17451,N_11479,N_11358);
or U17452 (N_17452,N_11858,N_13701);
xnor U17453 (N_17453,N_10768,N_14538);
or U17454 (N_17454,N_13248,N_14793);
nand U17455 (N_17455,N_11333,N_10165);
xnor U17456 (N_17456,N_11992,N_11323);
nand U17457 (N_17457,N_10749,N_11873);
nor U17458 (N_17458,N_10781,N_12833);
nor U17459 (N_17459,N_14531,N_12154);
nor U17460 (N_17460,N_13966,N_14692);
xnor U17461 (N_17461,N_10892,N_10722);
xor U17462 (N_17462,N_11737,N_12870);
xnor U17463 (N_17463,N_13580,N_11649);
or U17464 (N_17464,N_14571,N_11830);
xor U17465 (N_17465,N_14288,N_11104);
nor U17466 (N_17466,N_13029,N_13511);
nor U17467 (N_17467,N_12903,N_12222);
nand U17468 (N_17468,N_14063,N_12106);
xor U17469 (N_17469,N_13520,N_10723);
nor U17470 (N_17470,N_10414,N_12110);
xnor U17471 (N_17471,N_10132,N_14156);
xnor U17472 (N_17472,N_12763,N_11502);
or U17473 (N_17473,N_12893,N_13829);
xor U17474 (N_17474,N_10930,N_13964);
nand U17475 (N_17475,N_10856,N_14871);
and U17476 (N_17476,N_12095,N_11622);
xor U17477 (N_17477,N_10370,N_12926);
nand U17478 (N_17478,N_12740,N_11180);
or U17479 (N_17479,N_13507,N_14301);
or U17480 (N_17480,N_13620,N_12381);
or U17481 (N_17481,N_12238,N_14097);
and U17482 (N_17482,N_13791,N_11025);
or U17483 (N_17483,N_10131,N_11433);
and U17484 (N_17484,N_14565,N_14176);
xnor U17485 (N_17485,N_13436,N_10772);
nor U17486 (N_17486,N_10586,N_14506);
or U17487 (N_17487,N_11051,N_12182);
nand U17488 (N_17488,N_10196,N_11711);
nand U17489 (N_17489,N_13744,N_10926);
or U17490 (N_17490,N_14938,N_13843);
and U17491 (N_17491,N_14314,N_10584);
or U17492 (N_17492,N_11016,N_11619);
xor U17493 (N_17493,N_10214,N_13935);
or U17494 (N_17494,N_14065,N_13439);
nor U17495 (N_17495,N_14323,N_14011);
nand U17496 (N_17496,N_11192,N_10320);
nor U17497 (N_17497,N_12753,N_13429);
nor U17498 (N_17498,N_13232,N_14750);
xor U17499 (N_17499,N_13603,N_11262);
nor U17500 (N_17500,N_14755,N_11187);
xnor U17501 (N_17501,N_10192,N_10595);
or U17502 (N_17502,N_11295,N_11138);
xor U17503 (N_17503,N_10844,N_11480);
nand U17504 (N_17504,N_11737,N_14353);
or U17505 (N_17505,N_10598,N_10980);
nor U17506 (N_17506,N_14366,N_14975);
and U17507 (N_17507,N_12219,N_14978);
or U17508 (N_17508,N_13925,N_12535);
and U17509 (N_17509,N_14708,N_11577);
nand U17510 (N_17510,N_14229,N_12107);
nand U17511 (N_17511,N_12451,N_13775);
nor U17512 (N_17512,N_13937,N_12275);
xnor U17513 (N_17513,N_11868,N_10427);
nor U17514 (N_17514,N_11398,N_11111);
and U17515 (N_17515,N_14357,N_10443);
and U17516 (N_17516,N_13851,N_10991);
and U17517 (N_17517,N_10543,N_13960);
nor U17518 (N_17518,N_12072,N_10611);
xnor U17519 (N_17519,N_10350,N_11100);
nor U17520 (N_17520,N_13411,N_10492);
nor U17521 (N_17521,N_10355,N_14840);
and U17522 (N_17522,N_10431,N_11105);
or U17523 (N_17523,N_10634,N_12105);
xnor U17524 (N_17524,N_11009,N_10976);
nand U17525 (N_17525,N_12901,N_10030);
nor U17526 (N_17526,N_10414,N_10700);
nand U17527 (N_17527,N_12758,N_10442);
xnor U17528 (N_17528,N_10468,N_12044);
or U17529 (N_17529,N_11329,N_11202);
or U17530 (N_17530,N_10564,N_12859);
nor U17531 (N_17531,N_10017,N_14814);
and U17532 (N_17532,N_13536,N_13255);
xnor U17533 (N_17533,N_11653,N_14029);
xnor U17534 (N_17534,N_13283,N_11379);
nor U17535 (N_17535,N_12784,N_13319);
or U17536 (N_17536,N_10777,N_14528);
xnor U17537 (N_17537,N_10910,N_12379);
or U17538 (N_17538,N_10105,N_13300);
nor U17539 (N_17539,N_11307,N_10969);
and U17540 (N_17540,N_14831,N_10385);
and U17541 (N_17541,N_11483,N_10610);
nor U17542 (N_17542,N_14096,N_14740);
nand U17543 (N_17543,N_14412,N_10490);
nor U17544 (N_17544,N_14501,N_13459);
nor U17545 (N_17545,N_10824,N_10437);
xnor U17546 (N_17546,N_10473,N_12063);
nor U17547 (N_17547,N_13384,N_14152);
or U17548 (N_17548,N_13550,N_12928);
nor U17549 (N_17549,N_10750,N_13954);
nand U17550 (N_17550,N_12059,N_13252);
nand U17551 (N_17551,N_14778,N_13999);
nor U17552 (N_17552,N_11100,N_13091);
nor U17553 (N_17553,N_10314,N_13148);
nand U17554 (N_17554,N_12080,N_11419);
or U17555 (N_17555,N_13796,N_10749);
nor U17556 (N_17556,N_11684,N_12656);
nand U17557 (N_17557,N_11029,N_13507);
nor U17558 (N_17558,N_14535,N_14347);
and U17559 (N_17559,N_14047,N_14600);
nand U17560 (N_17560,N_11217,N_14201);
nor U17561 (N_17561,N_11505,N_13496);
and U17562 (N_17562,N_12062,N_11149);
nand U17563 (N_17563,N_12101,N_14619);
and U17564 (N_17564,N_12409,N_13503);
and U17565 (N_17565,N_14072,N_12808);
nand U17566 (N_17566,N_12304,N_11617);
or U17567 (N_17567,N_14090,N_10969);
or U17568 (N_17568,N_10289,N_13725);
and U17569 (N_17569,N_13516,N_11413);
or U17570 (N_17570,N_11549,N_14820);
or U17571 (N_17571,N_12958,N_13428);
nand U17572 (N_17572,N_12106,N_13403);
xor U17573 (N_17573,N_10996,N_12235);
xor U17574 (N_17574,N_12849,N_12578);
and U17575 (N_17575,N_14619,N_13840);
nor U17576 (N_17576,N_12193,N_13903);
or U17577 (N_17577,N_11700,N_13062);
xnor U17578 (N_17578,N_14232,N_11028);
nor U17579 (N_17579,N_11586,N_11214);
nor U17580 (N_17580,N_12659,N_13137);
xor U17581 (N_17581,N_12662,N_11331);
nor U17582 (N_17582,N_11178,N_11940);
nor U17583 (N_17583,N_12338,N_12358);
nor U17584 (N_17584,N_13409,N_10304);
and U17585 (N_17585,N_11811,N_12543);
nor U17586 (N_17586,N_14616,N_12394);
or U17587 (N_17587,N_14842,N_12581);
nand U17588 (N_17588,N_14371,N_10153);
xor U17589 (N_17589,N_11603,N_14386);
nand U17590 (N_17590,N_13420,N_14438);
nor U17591 (N_17591,N_10752,N_11828);
or U17592 (N_17592,N_11548,N_13439);
or U17593 (N_17593,N_11884,N_12289);
nor U17594 (N_17594,N_14358,N_12374);
nand U17595 (N_17595,N_10279,N_12167);
or U17596 (N_17596,N_12661,N_11352);
xnor U17597 (N_17597,N_14543,N_12747);
nand U17598 (N_17598,N_12752,N_10830);
or U17599 (N_17599,N_10692,N_11648);
nor U17600 (N_17600,N_12099,N_13496);
nand U17601 (N_17601,N_10729,N_13682);
nand U17602 (N_17602,N_13418,N_14041);
xor U17603 (N_17603,N_14836,N_12179);
nor U17604 (N_17604,N_12538,N_13462);
nand U17605 (N_17605,N_10143,N_10581);
nand U17606 (N_17606,N_11047,N_12427);
nor U17607 (N_17607,N_14118,N_14563);
xor U17608 (N_17608,N_11455,N_10295);
xor U17609 (N_17609,N_11285,N_12988);
xor U17610 (N_17610,N_12379,N_11477);
nor U17611 (N_17611,N_14188,N_12907);
nor U17612 (N_17612,N_10895,N_12236);
nor U17613 (N_17613,N_10903,N_10868);
nand U17614 (N_17614,N_14584,N_12710);
or U17615 (N_17615,N_10187,N_11189);
nor U17616 (N_17616,N_13911,N_13770);
nor U17617 (N_17617,N_12328,N_14632);
nor U17618 (N_17618,N_12954,N_13010);
xor U17619 (N_17619,N_13689,N_14861);
or U17620 (N_17620,N_14791,N_12693);
nor U17621 (N_17621,N_11333,N_14492);
nor U17622 (N_17622,N_12144,N_12540);
nand U17623 (N_17623,N_13926,N_14749);
or U17624 (N_17624,N_11994,N_10571);
nor U17625 (N_17625,N_14762,N_13933);
nand U17626 (N_17626,N_11651,N_12844);
and U17627 (N_17627,N_11274,N_11356);
xnor U17628 (N_17628,N_11703,N_14937);
and U17629 (N_17629,N_14680,N_11944);
xnor U17630 (N_17630,N_12889,N_12307);
or U17631 (N_17631,N_10053,N_13632);
or U17632 (N_17632,N_11737,N_13587);
and U17633 (N_17633,N_13253,N_10439);
and U17634 (N_17634,N_11757,N_14328);
nand U17635 (N_17635,N_10568,N_14902);
xor U17636 (N_17636,N_10344,N_11560);
and U17637 (N_17637,N_14209,N_12710);
xor U17638 (N_17638,N_12248,N_10620);
nand U17639 (N_17639,N_11288,N_14474);
nor U17640 (N_17640,N_13466,N_14209);
nor U17641 (N_17641,N_11499,N_13486);
or U17642 (N_17642,N_10484,N_12854);
or U17643 (N_17643,N_11172,N_12659);
and U17644 (N_17644,N_14828,N_11687);
xor U17645 (N_17645,N_11102,N_14056);
and U17646 (N_17646,N_10035,N_10513);
xor U17647 (N_17647,N_10064,N_10474);
or U17648 (N_17648,N_14018,N_14368);
and U17649 (N_17649,N_11986,N_13205);
xor U17650 (N_17650,N_13101,N_13869);
xnor U17651 (N_17651,N_10103,N_12525);
or U17652 (N_17652,N_13608,N_14734);
and U17653 (N_17653,N_14090,N_12170);
xor U17654 (N_17654,N_12997,N_12446);
and U17655 (N_17655,N_13088,N_13733);
nor U17656 (N_17656,N_12470,N_13292);
nor U17657 (N_17657,N_14493,N_14377);
and U17658 (N_17658,N_12077,N_10854);
nor U17659 (N_17659,N_10445,N_10926);
nand U17660 (N_17660,N_13653,N_10488);
nand U17661 (N_17661,N_13049,N_13472);
nand U17662 (N_17662,N_13650,N_13116);
nor U17663 (N_17663,N_13195,N_13352);
or U17664 (N_17664,N_13363,N_11796);
nand U17665 (N_17665,N_10189,N_14869);
nand U17666 (N_17666,N_13383,N_13747);
nand U17667 (N_17667,N_12520,N_10924);
nor U17668 (N_17668,N_14090,N_11429);
and U17669 (N_17669,N_10758,N_13197);
and U17670 (N_17670,N_11828,N_14096);
or U17671 (N_17671,N_11931,N_11523);
or U17672 (N_17672,N_10984,N_12769);
and U17673 (N_17673,N_13798,N_10320);
or U17674 (N_17674,N_10298,N_10204);
or U17675 (N_17675,N_10984,N_13660);
nor U17676 (N_17676,N_14845,N_11813);
nand U17677 (N_17677,N_11122,N_10217);
or U17678 (N_17678,N_10074,N_13091);
nor U17679 (N_17679,N_13361,N_14178);
xnor U17680 (N_17680,N_14626,N_10927);
or U17681 (N_17681,N_10901,N_14032);
xnor U17682 (N_17682,N_10628,N_10926);
and U17683 (N_17683,N_12588,N_14338);
or U17684 (N_17684,N_10597,N_10298);
or U17685 (N_17685,N_12038,N_14531);
or U17686 (N_17686,N_14967,N_13525);
or U17687 (N_17687,N_12426,N_13225);
nand U17688 (N_17688,N_12158,N_11651);
and U17689 (N_17689,N_12871,N_10792);
xnor U17690 (N_17690,N_12248,N_10006);
nor U17691 (N_17691,N_13225,N_13757);
nand U17692 (N_17692,N_13037,N_11263);
nand U17693 (N_17693,N_13752,N_10600);
and U17694 (N_17694,N_13869,N_12302);
and U17695 (N_17695,N_12509,N_10718);
nand U17696 (N_17696,N_14472,N_10871);
xor U17697 (N_17697,N_10291,N_10356);
and U17698 (N_17698,N_10407,N_10107);
and U17699 (N_17699,N_13029,N_12240);
nand U17700 (N_17700,N_11751,N_12525);
nor U17701 (N_17701,N_14809,N_14286);
xor U17702 (N_17702,N_10912,N_10414);
nand U17703 (N_17703,N_14326,N_11274);
nand U17704 (N_17704,N_14475,N_10487);
nand U17705 (N_17705,N_12257,N_14103);
and U17706 (N_17706,N_11136,N_14169);
xor U17707 (N_17707,N_14078,N_11132);
or U17708 (N_17708,N_11901,N_14921);
nand U17709 (N_17709,N_12166,N_14389);
nor U17710 (N_17710,N_14887,N_13358);
nand U17711 (N_17711,N_10954,N_12079);
nor U17712 (N_17712,N_13666,N_14239);
or U17713 (N_17713,N_14295,N_12313);
nor U17714 (N_17714,N_11584,N_13836);
nor U17715 (N_17715,N_13266,N_13410);
or U17716 (N_17716,N_14572,N_11892);
or U17717 (N_17717,N_10812,N_10912);
nand U17718 (N_17718,N_11292,N_14208);
xnor U17719 (N_17719,N_10622,N_11363);
and U17720 (N_17720,N_11313,N_10233);
nor U17721 (N_17721,N_11946,N_14583);
or U17722 (N_17722,N_14107,N_14653);
nand U17723 (N_17723,N_11016,N_11371);
xnor U17724 (N_17724,N_10761,N_14839);
xnor U17725 (N_17725,N_13348,N_13018);
and U17726 (N_17726,N_10033,N_10978);
nor U17727 (N_17727,N_12090,N_13473);
nor U17728 (N_17728,N_10801,N_13366);
nand U17729 (N_17729,N_11944,N_10003);
and U17730 (N_17730,N_14515,N_11104);
or U17731 (N_17731,N_13226,N_11233);
or U17732 (N_17732,N_13372,N_10622);
nor U17733 (N_17733,N_14271,N_10255);
nand U17734 (N_17734,N_12297,N_13596);
or U17735 (N_17735,N_13996,N_13082);
nand U17736 (N_17736,N_10481,N_13426);
nand U17737 (N_17737,N_14334,N_14890);
nor U17738 (N_17738,N_14077,N_10265);
xnor U17739 (N_17739,N_10778,N_10528);
nand U17740 (N_17740,N_14494,N_12139);
or U17741 (N_17741,N_13684,N_12009);
nand U17742 (N_17742,N_10100,N_10540);
nor U17743 (N_17743,N_12352,N_12055);
and U17744 (N_17744,N_10630,N_12422);
nand U17745 (N_17745,N_12190,N_12333);
nand U17746 (N_17746,N_12465,N_10946);
or U17747 (N_17747,N_14116,N_10993);
nor U17748 (N_17748,N_11892,N_10451);
or U17749 (N_17749,N_13759,N_12310);
xor U17750 (N_17750,N_11645,N_10501);
xnor U17751 (N_17751,N_14760,N_11687);
nor U17752 (N_17752,N_10464,N_10276);
or U17753 (N_17753,N_13973,N_10370);
nor U17754 (N_17754,N_13036,N_13389);
nand U17755 (N_17755,N_10094,N_11295);
xor U17756 (N_17756,N_12194,N_13605);
or U17757 (N_17757,N_14047,N_13913);
nand U17758 (N_17758,N_12824,N_11373);
xnor U17759 (N_17759,N_13816,N_12121);
or U17760 (N_17760,N_12060,N_11568);
nor U17761 (N_17761,N_10111,N_11076);
and U17762 (N_17762,N_13617,N_12239);
nor U17763 (N_17763,N_13704,N_14713);
nor U17764 (N_17764,N_10098,N_12273);
and U17765 (N_17765,N_10307,N_11944);
xor U17766 (N_17766,N_10662,N_12210);
nor U17767 (N_17767,N_14693,N_14732);
nand U17768 (N_17768,N_10892,N_13790);
nand U17769 (N_17769,N_13068,N_14125);
and U17770 (N_17770,N_10490,N_13719);
or U17771 (N_17771,N_11565,N_12677);
and U17772 (N_17772,N_12001,N_10948);
nor U17773 (N_17773,N_10452,N_13820);
nor U17774 (N_17774,N_10313,N_14455);
xor U17775 (N_17775,N_12717,N_12765);
nand U17776 (N_17776,N_13133,N_13119);
nand U17777 (N_17777,N_14065,N_12474);
xor U17778 (N_17778,N_11655,N_12209);
or U17779 (N_17779,N_12516,N_13199);
xor U17780 (N_17780,N_14990,N_11550);
nor U17781 (N_17781,N_14626,N_13011);
nand U17782 (N_17782,N_12055,N_10775);
or U17783 (N_17783,N_12291,N_12957);
and U17784 (N_17784,N_10628,N_13352);
nand U17785 (N_17785,N_12488,N_12074);
xor U17786 (N_17786,N_10953,N_10914);
xor U17787 (N_17787,N_10490,N_13601);
and U17788 (N_17788,N_13851,N_14427);
and U17789 (N_17789,N_13981,N_14494);
or U17790 (N_17790,N_12990,N_10494);
nand U17791 (N_17791,N_13557,N_10375);
xnor U17792 (N_17792,N_11544,N_10148);
xnor U17793 (N_17793,N_14355,N_12626);
and U17794 (N_17794,N_11186,N_10872);
and U17795 (N_17795,N_12535,N_10553);
xnor U17796 (N_17796,N_14642,N_10937);
nand U17797 (N_17797,N_11269,N_14713);
nand U17798 (N_17798,N_13002,N_12718);
nand U17799 (N_17799,N_12656,N_14848);
and U17800 (N_17800,N_14723,N_13079);
or U17801 (N_17801,N_13569,N_11359);
nand U17802 (N_17802,N_10303,N_14365);
xnor U17803 (N_17803,N_13927,N_13985);
nand U17804 (N_17804,N_11891,N_12033);
and U17805 (N_17805,N_10792,N_11007);
nor U17806 (N_17806,N_10656,N_12751);
nand U17807 (N_17807,N_13486,N_13499);
nor U17808 (N_17808,N_11927,N_13683);
nand U17809 (N_17809,N_10346,N_12593);
or U17810 (N_17810,N_11066,N_11016);
nor U17811 (N_17811,N_11356,N_10115);
nor U17812 (N_17812,N_11607,N_10349);
nand U17813 (N_17813,N_12742,N_13386);
or U17814 (N_17814,N_14716,N_12481);
nor U17815 (N_17815,N_10381,N_10831);
nand U17816 (N_17816,N_10150,N_10421);
or U17817 (N_17817,N_12410,N_13908);
and U17818 (N_17818,N_14612,N_10564);
and U17819 (N_17819,N_12561,N_11914);
nand U17820 (N_17820,N_10896,N_11379);
xor U17821 (N_17821,N_14982,N_10541);
or U17822 (N_17822,N_13425,N_14466);
and U17823 (N_17823,N_10600,N_12685);
nand U17824 (N_17824,N_14225,N_13298);
nand U17825 (N_17825,N_13605,N_10077);
nand U17826 (N_17826,N_10163,N_10086);
xor U17827 (N_17827,N_14546,N_12063);
xnor U17828 (N_17828,N_11510,N_12066);
xor U17829 (N_17829,N_10967,N_11462);
nor U17830 (N_17830,N_11659,N_10983);
and U17831 (N_17831,N_10298,N_14289);
or U17832 (N_17832,N_14118,N_11061);
and U17833 (N_17833,N_12107,N_14995);
nor U17834 (N_17834,N_13676,N_12436);
xnor U17835 (N_17835,N_10721,N_14192);
nor U17836 (N_17836,N_12368,N_12608);
xor U17837 (N_17837,N_14855,N_12087);
or U17838 (N_17838,N_14501,N_10678);
xnor U17839 (N_17839,N_11343,N_10781);
xor U17840 (N_17840,N_12733,N_11000);
and U17841 (N_17841,N_11382,N_13521);
nand U17842 (N_17842,N_11300,N_14952);
or U17843 (N_17843,N_12496,N_14922);
xnor U17844 (N_17844,N_10726,N_12200);
or U17845 (N_17845,N_13367,N_14006);
nor U17846 (N_17846,N_11369,N_10336);
xnor U17847 (N_17847,N_13962,N_14350);
xnor U17848 (N_17848,N_12601,N_11116);
nand U17849 (N_17849,N_14692,N_13763);
xnor U17850 (N_17850,N_10417,N_11446);
and U17851 (N_17851,N_10686,N_11727);
or U17852 (N_17852,N_14487,N_12722);
nor U17853 (N_17853,N_11167,N_11191);
xnor U17854 (N_17854,N_11468,N_12176);
and U17855 (N_17855,N_12704,N_11923);
nor U17856 (N_17856,N_10393,N_12083);
or U17857 (N_17857,N_13215,N_12329);
nor U17858 (N_17858,N_13057,N_12474);
nor U17859 (N_17859,N_11054,N_10301);
and U17860 (N_17860,N_14067,N_11618);
nand U17861 (N_17861,N_11440,N_12195);
nand U17862 (N_17862,N_11819,N_10277);
xor U17863 (N_17863,N_14023,N_11342);
or U17864 (N_17864,N_10316,N_11266);
or U17865 (N_17865,N_13093,N_14342);
nand U17866 (N_17866,N_13919,N_12825);
and U17867 (N_17867,N_14459,N_11912);
and U17868 (N_17868,N_13714,N_13112);
xnor U17869 (N_17869,N_13152,N_13446);
xor U17870 (N_17870,N_12027,N_14415);
xnor U17871 (N_17871,N_12100,N_14065);
nand U17872 (N_17872,N_14243,N_14961);
nor U17873 (N_17873,N_10703,N_13158);
and U17874 (N_17874,N_10271,N_13640);
or U17875 (N_17875,N_13350,N_10803);
or U17876 (N_17876,N_13136,N_13271);
and U17877 (N_17877,N_14067,N_12128);
xnor U17878 (N_17878,N_12159,N_11486);
nor U17879 (N_17879,N_10818,N_10950);
nand U17880 (N_17880,N_10462,N_10988);
nand U17881 (N_17881,N_10241,N_11287);
xor U17882 (N_17882,N_12106,N_13040);
or U17883 (N_17883,N_12590,N_14786);
nand U17884 (N_17884,N_13820,N_13914);
or U17885 (N_17885,N_14797,N_13544);
nor U17886 (N_17886,N_11207,N_12107);
nor U17887 (N_17887,N_10360,N_10770);
and U17888 (N_17888,N_12765,N_12804);
nor U17889 (N_17889,N_14122,N_13063);
and U17890 (N_17890,N_12451,N_11615);
nor U17891 (N_17891,N_11906,N_12940);
nand U17892 (N_17892,N_10847,N_10134);
nand U17893 (N_17893,N_14682,N_13354);
and U17894 (N_17894,N_14246,N_10741);
or U17895 (N_17895,N_13490,N_12123);
nor U17896 (N_17896,N_11605,N_10876);
nor U17897 (N_17897,N_12803,N_10449);
xnor U17898 (N_17898,N_14148,N_13629);
or U17899 (N_17899,N_10107,N_14638);
xor U17900 (N_17900,N_10318,N_13274);
nor U17901 (N_17901,N_10012,N_12238);
nand U17902 (N_17902,N_14595,N_11304);
nand U17903 (N_17903,N_13975,N_10111);
or U17904 (N_17904,N_12121,N_13040);
nand U17905 (N_17905,N_14948,N_14294);
and U17906 (N_17906,N_14395,N_10225);
and U17907 (N_17907,N_11076,N_11917);
and U17908 (N_17908,N_10834,N_14208);
xor U17909 (N_17909,N_14356,N_10823);
xor U17910 (N_17910,N_10484,N_10184);
or U17911 (N_17911,N_13619,N_12864);
and U17912 (N_17912,N_13054,N_10727);
nor U17913 (N_17913,N_10604,N_12371);
or U17914 (N_17914,N_13782,N_14287);
nor U17915 (N_17915,N_14342,N_14616);
or U17916 (N_17916,N_13749,N_13786);
nand U17917 (N_17917,N_11441,N_12136);
nand U17918 (N_17918,N_12160,N_11551);
or U17919 (N_17919,N_10148,N_10952);
nor U17920 (N_17920,N_13270,N_11867);
nand U17921 (N_17921,N_11346,N_13608);
nand U17922 (N_17922,N_13427,N_12593);
and U17923 (N_17923,N_12358,N_11003);
nand U17924 (N_17924,N_13559,N_12188);
nand U17925 (N_17925,N_13491,N_11041);
or U17926 (N_17926,N_12564,N_13507);
nor U17927 (N_17927,N_12366,N_11479);
nand U17928 (N_17928,N_11748,N_10047);
nor U17929 (N_17929,N_10986,N_11537);
xor U17930 (N_17930,N_11177,N_14756);
and U17931 (N_17931,N_12526,N_12811);
or U17932 (N_17932,N_12759,N_12460);
nand U17933 (N_17933,N_14877,N_13749);
or U17934 (N_17934,N_13054,N_11806);
and U17935 (N_17935,N_12985,N_11851);
nand U17936 (N_17936,N_13557,N_13623);
nor U17937 (N_17937,N_14987,N_14841);
nand U17938 (N_17938,N_11577,N_14463);
nand U17939 (N_17939,N_12562,N_10304);
and U17940 (N_17940,N_13541,N_11497);
nand U17941 (N_17941,N_12978,N_10979);
nor U17942 (N_17942,N_14367,N_12869);
nor U17943 (N_17943,N_13863,N_13850);
nand U17944 (N_17944,N_11763,N_12371);
or U17945 (N_17945,N_10531,N_12031);
and U17946 (N_17946,N_12436,N_11292);
xor U17947 (N_17947,N_14738,N_11289);
and U17948 (N_17948,N_14731,N_10988);
xnor U17949 (N_17949,N_10442,N_10771);
xnor U17950 (N_17950,N_12723,N_10065);
nand U17951 (N_17951,N_13422,N_10859);
xor U17952 (N_17952,N_14691,N_13270);
nand U17953 (N_17953,N_12858,N_14343);
xnor U17954 (N_17954,N_13810,N_11060);
and U17955 (N_17955,N_13237,N_14451);
and U17956 (N_17956,N_10940,N_11973);
nor U17957 (N_17957,N_10591,N_13086);
and U17958 (N_17958,N_13545,N_11726);
nor U17959 (N_17959,N_14112,N_11961);
nor U17960 (N_17960,N_14626,N_10040);
nor U17961 (N_17961,N_13491,N_10680);
nand U17962 (N_17962,N_10138,N_11288);
nor U17963 (N_17963,N_14930,N_10659);
nor U17964 (N_17964,N_10780,N_11292);
nand U17965 (N_17965,N_13617,N_14433);
and U17966 (N_17966,N_12050,N_12918);
and U17967 (N_17967,N_10319,N_11099);
xnor U17968 (N_17968,N_10101,N_11505);
nor U17969 (N_17969,N_10341,N_14867);
nand U17970 (N_17970,N_11937,N_13476);
or U17971 (N_17971,N_11533,N_13284);
xor U17972 (N_17972,N_12293,N_10103);
and U17973 (N_17973,N_13487,N_14426);
nor U17974 (N_17974,N_10499,N_10968);
or U17975 (N_17975,N_13201,N_12595);
nand U17976 (N_17976,N_10128,N_13332);
nand U17977 (N_17977,N_12472,N_10577);
or U17978 (N_17978,N_12515,N_10728);
or U17979 (N_17979,N_14953,N_13752);
nand U17980 (N_17980,N_13672,N_13487);
nand U17981 (N_17981,N_12496,N_10869);
or U17982 (N_17982,N_12657,N_13980);
or U17983 (N_17983,N_11516,N_10999);
nor U17984 (N_17984,N_10350,N_14386);
xnor U17985 (N_17985,N_13875,N_13410);
nor U17986 (N_17986,N_11883,N_12986);
and U17987 (N_17987,N_12090,N_11533);
or U17988 (N_17988,N_13709,N_12968);
nor U17989 (N_17989,N_14769,N_13715);
and U17990 (N_17990,N_13503,N_10373);
or U17991 (N_17991,N_13446,N_13745);
nand U17992 (N_17992,N_13099,N_10630);
xnor U17993 (N_17993,N_10076,N_12549);
or U17994 (N_17994,N_14121,N_14436);
or U17995 (N_17995,N_14560,N_13271);
nand U17996 (N_17996,N_12874,N_11557);
nor U17997 (N_17997,N_12016,N_10716);
xor U17998 (N_17998,N_13469,N_13118);
and U17999 (N_17999,N_12020,N_11936);
xor U18000 (N_18000,N_14911,N_14079);
nand U18001 (N_18001,N_12027,N_10072);
and U18002 (N_18002,N_14163,N_11327);
nand U18003 (N_18003,N_11892,N_13761);
nor U18004 (N_18004,N_14120,N_13910);
xnor U18005 (N_18005,N_10248,N_13537);
xnor U18006 (N_18006,N_13909,N_12616);
and U18007 (N_18007,N_10332,N_13487);
xor U18008 (N_18008,N_14181,N_13578);
xnor U18009 (N_18009,N_10742,N_13776);
and U18010 (N_18010,N_10346,N_14924);
nor U18011 (N_18011,N_11699,N_13156);
and U18012 (N_18012,N_12819,N_11579);
or U18013 (N_18013,N_12357,N_13088);
or U18014 (N_18014,N_13557,N_14195);
and U18015 (N_18015,N_14508,N_10258);
xor U18016 (N_18016,N_10812,N_12687);
nor U18017 (N_18017,N_11733,N_11914);
nand U18018 (N_18018,N_13108,N_10702);
nand U18019 (N_18019,N_12900,N_14048);
or U18020 (N_18020,N_12964,N_14009);
or U18021 (N_18021,N_13720,N_10179);
or U18022 (N_18022,N_14361,N_11704);
xor U18023 (N_18023,N_12076,N_11998);
xor U18024 (N_18024,N_10292,N_14367);
nand U18025 (N_18025,N_14245,N_14918);
nand U18026 (N_18026,N_13716,N_10824);
and U18027 (N_18027,N_11640,N_14326);
xnor U18028 (N_18028,N_12809,N_13181);
and U18029 (N_18029,N_14923,N_13798);
nand U18030 (N_18030,N_13853,N_13374);
xor U18031 (N_18031,N_11620,N_13914);
or U18032 (N_18032,N_11797,N_10642);
nor U18033 (N_18033,N_13265,N_13388);
xnor U18034 (N_18034,N_10349,N_12560);
nor U18035 (N_18035,N_13550,N_12369);
xor U18036 (N_18036,N_10359,N_10174);
nand U18037 (N_18037,N_11150,N_11058);
nand U18038 (N_18038,N_12132,N_10593);
nor U18039 (N_18039,N_12910,N_13817);
xor U18040 (N_18040,N_11579,N_10381);
and U18041 (N_18041,N_10265,N_12334);
nor U18042 (N_18042,N_13811,N_10367);
xor U18043 (N_18043,N_12652,N_11824);
nand U18044 (N_18044,N_10601,N_13109);
xor U18045 (N_18045,N_10847,N_12609);
or U18046 (N_18046,N_12004,N_12094);
and U18047 (N_18047,N_14462,N_14097);
nor U18048 (N_18048,N_10731,N_11752);
nor U18049 (N_18049,N_11022,N_12936);
nor U18050 (N_18050,N_10042,N_12594);
nor U18051 (N_18051,N_13582,N_11482);
and U18052 (N_18052,N_11302,N_13990);
nand U18053 (N_18053,N_10994,N_10831);
nor U18054 (N_18054,N_10895,N_14895);
nand U18055 (N_18055,N_10400,N_14770);
nand U18056 (N_18056,N_13766,N_11074);
xnor U18057 (N_18057,N_13919,N_11185);
nor U18058 (N_18058,N_14274,N_14048);
nand U18059 (N_18059,N_12905,N_11647);
xnor U18060 (N_18060,N_12365,N_13404);
nand U18061 (N_18061,N_11953,N_12896);
xnor U18062 (N_18062,N_13598,N_13540);
xnor U18063 (N_18063,N_14299,N_10619);
or U18064 (N_18064,N_12979,N_13957);
nor U18065 (N_18065,N_11685,N_10335);
nor U18066 (N_18066,N_14655,N_13525);
nor U18067 (N_18067,N_13343,N_14491);
nor U18068 (N_18068,N_10770,N_10715);
xnor U18069 (N_18069,N_11210,N_10691);
or U18070 (N_18070,N_12749,N_12286);
nor U18071 (N_18071,N_11782,N_10870);
or U18072 (N_18072,N_13410,N_12590);
nor U18073 (N_18073,N_13101,N_10269);
or U18074 (N_18074,N_10170,N_11584);
or U18075 (N_18075,N_13472,N_13217);
nor U18076 (N_18076,N_11038,N_12501);
and U18077 (N_18077,N_14786,N_11151);
nand U18078 (N_18078,N_10513,N_13805);
nor U18079 (N_18079,N_14801,N_10611);
nand U18080 (N_18080,N_10158,N_13776);
and U18081 (N_18081,N_10849,N_11364);
and U18082 (N_18082,N_14794,N_11818);
xor U18083 (N_18083,N_14757,N_13136);
and U18084 (N_18084,N_11961,N_11979);
nor U18085 (N_18085,N_14020,N_14956);
xor U18086 (N_18086,N_11893,N_14449);
and U18087 (N_18087,N_12252,N_14686);
nor U18088 (N_18088,N_11144,N_10950);
xnor U18089 (N_18089,N_10399,N_10493);
or U18090 (N_18090,N_14491,N_12659);
nor U18091 (N_18091,N_11533,N_10818);
and U18092 (N_18092,N_12965,N_13202);
and U18093 (N_18093,N_11423,N_13378);
and U18094 (N_18094,N_12403,N_10904);
nor U18095 (N_18095,N_12032,N_14095);
or U18096 (N_18096,N_13454,N_14336);
and U18097 (N_18097,N_11239,N_14686);
xor U18098 (N_18098,N_14172,N_13984);
nand U18099 (N_18099,N_12186,N_10692);
and U18100 (N_18100,N_10292,N_14047);
nand U18101 (N_18101,N_14658,N_14831);
and U18102 (N_18102,N_12438,N_12034);
xnor U18103 (N_18103,N_14745,N_11440);
nand U18104 (N_18104,N_10376,N_12224);
nor U18105 (N_18105,N_13959,N_12024);
xnor U18106 (N_18106,N_14770,N_14123);
nor U18107 (N_18107,N_12955,N_11316);
or U18108 (N_18108,N_10038,N_14376);
and U18109 (N_18109,N_10818,N_14120);
xor U18110 (N_18110,N_12805,N_12887);
or U18111 (N_18111,N_14213,N_14731);
nor U18112 (N_18112,N_14577,N_11537);
nand U18113 (N_18113,N_10334,N_12705);
xnor U18114 (N_18114,N_12237,N_11421);
nand U18115 (N_18115,N_11552,N_10827);
xnor U18116 (N_18116,N_13977,N_11900);
nor U18117 (N_18117,N_11245,N_14551);
or U18118 (N_18118,N_11045,N_14566);
nand U18119 (N_18119,N_10040,N_11558);
or U18120 (N_18120,N_11916,N_14688);
nor U18121 (N_18121,N_11271,N_10624);
and U18122 (N_18122,N_14467,N_11968);
nand U18123 (N_18123,N_12282,N_11345);
xnor U18124 (N_18124,N_12956,N_11217);
or U18125 (N_18125,N_10750,N_13321);
xor U18126 (N_18126,N_10977,N_12108);
nor U18127 (N_18127,N_14282,N_10790);
and U18128 (N_18128,N_12680,N_11827);
nor U18129 (N_18129,N_12419,N_13290);
or U18130 (N_18130,N_10932,N_13791);
or U18131 (N_18131,N_12260,N_11479);
xor U18132 (N_18132,N_13659,N_10984);
or U18133 (N_18133,N_12141,N_12565);
and U18134 (N_18134,N_13133,N_10424);
and U18135 (N_18135,N_14779,N_11699);
xor U18136 (N_18136,N_11988,N_10563);
nor U18137 (N_18137,N_10487,N_14156);
nand U18138 (N_18138,N_13948,N_13774);
nand U18139 (N_18139,N_10680,N_14086);
or U18140 (N_18140,N_12449,N_14117);
nand U18141 (N_18141,N_14151,N_14594);
or U18142 (N_18142,N_11322,N_11449);
or U18143 (N_18143,N_14660,N_12404);
and U18144 (N_18144,N_13891,N_13910);
and U18145 (N_18145,N_10946,N_12667);
and U18146 (N_18146,N_12476,N_13549);
xnor U18147 (N_18147,N_12659,N_11388);
nand U18148 (N_18148,N_12999,N_13163);
and U18149 (N_18149,N_13197,N_14830);
nor U18150 (N_18150,N_12097,N_10234);
and U18151 (N_18151,N_11289,N_13195);
nand U18152 (N_18152,N_13230,N_14506);
or U18153 (N_18153,N_14014,N_14651);
nor U18154 (N_18154,N_13743,N_10099);
and U18155 (N_18155,N_13134,N_14750);
nand U18156 (N_18156,N_13611,N_11227);
nand U18157 (N_18157,N_11769,N_14743);
or U18158 (N_18158,N_11873,N_13132);
and U18159 (N_18159,N_10448,N_13603);
xnor U18160 (N_18160,N_12967,N_10951);
nor U18161 (N_18161,N_10432,N_12966);
xnor U18162 (N_18162,N_11173,N_12390);
nor U18163 (N_18163,N_12374,N_13510);
or U18164 (N_18164,N_14731,N_13299);
nand U18165 (N_18165,N_11718,N_11227);
or U18166 (N_18166,N_13702,N_10561);
xnor U18167 (N_18167,N_13790,N_11779);
nand U18168 (N_18168,N_11220,N_14997);
nor U18169 (N_18169,N_14023,N_11869);
xnor U18170 (N_18170,N_11414,N_13614);
and U18171 (N_18171,N_10877,N_11251);
and U18172 (N_18172,N_13458,N_13019);
nor U18173 (N_18173,N_12301,N_12627);
and U18174 (N_18174,N_13395,N_11106);
nand U18175 (N_18175,N_11082,N_11660);
nor U18176 (N_18176,N_14416,N_10160);
nor U18177 (N_18177,N_10332,N_13903);
xor U18178 (N_18178,N_11182,N_14823);
xnor U18179 (N_18179,N_10487,N_14985);
nor U18180 (N_18180,N_12467,N_12297);
and U18181 (N_18181,N_11834,N_12926);
xnor U18182 (N_18182,N_12801,N_12233);
or U18183 (N_18183,N_14807,N_10345);
and U18184 (N_18184,N_13394,N_10947);
or U18185 (N_18185,N_12780,N_10777);
xor U18186 (N_18186,N_11956,N_12264);
and U18187 (N_18187,N_12274,N_10195);
nand U18188 (N_18188,N_10185,N_11601);
nand U18189 (N_18189,N_12674,N_11372);
and U18190 (N_18190,N_13694,N_12540);
or U18191 (N_18191,N_14200,N_10448);
or U18192 (N_18192,N_10322,N_14293);
nand U18193 (N_18193,N_14545,N_14136);
nand U18194 (N_18194,N_13777,N_14432);
xor U18195 (N_18195,N_13160,N_11441);
nor U18196 (N_18196,N_14538,N_10349);
xor U18197 (N_18197,N_14250,N_14443);
nand U18198 (N_18198,N_10296,N_11331);
and U18199 (N_18199,N_14443,N_13705);
and U18200 (N_18200,N_12329,N_14783);
and U18201 (N_18201,N_10447,N_13064);
and U18202 (N_18202,N_10198,N_13629);
nand U18203 (N_18203,N_10734,N_10334);
or U18204 (N_18204,N_13056,N_11573);
and U18205 (N_18205,N_13208,N_10772);
and U18206 (N_18206,N_12168,N_14610);
nor U18207 (N_18207,N_13994,N_12584);
xor U18208 (N_18208,N_13844,N_14565);
or U18209 (N_18209,N_14813,N_13709);
or U18210 (N_18210,N_12179,N_12192);
nand U18211 (N_18211,N_12609,N_11259);
nor U18212 (N_18212,N_14157,N_14428);
xnor U18213 (N_18213,N_11698,N_11727);
nand U18214 (N_18214,N_12174,N_13995);
or U18215 (N_18215,N_13342,N_14859);
nand U18216 (N_18216,N_10402,N_14007);
nand U18217 (N_18217,N_10597,N_11298);
nor U18218 (N_18218,N_13136,N_12524);
xor U18219 (N_18219,N_14020,N_10367);
and U18220 (N_18220,N_13017,N_10543);
xor U18221 (N_18221,N_14405,N_10984);
xnor U18222 (N_18222,N_12366,N_14008);
nor U18223 (N_18223,N_14433,N_14579);
nor U18224 (N_18224,N_13760,N_11445);
and U18225 (N_18225,N_12924,N_11456);
and U18226 (N_18226,N_11895,N_12793);
and U18227 (N_18227,N_12661,N_14951);
nand U18228 (N_18228,N_13698,N_11721);
nand U18229 (N_18229,N_12021,N_13050);
xor U18230 (N_18230,N_13614,N_14899);
nand U18231 (N_18231,N_14475,N_12900);
xor U18232 (N_18232,N_14970,N_11862);
nor U18233 (N_18233,N_11132,N_13486);
xnor U18234 (N_18234,N_11002,N_11432);
nand U18235 (N_18235,N_14014,N_12993);
nor U18236 (N_18236,N_10571,N_11180);
and U18237 (N_18237,N_12568,N_10281);
xnor U18238 (N_18238,N_14177,N_11294);
or U18239 (N_18239,N_13257,N_14797);
xnor U18240 (N_18240,N_11435,N_13855);
nor U18241 (N_18241,N_10476,N_11090);
nor U18242 (N_18242,N_12945,N_12198);
and U18243 (N_18243,N_12830,N_11802);
and U18244 (N_18244,N_11000,N_14581);
or U18245 (N_18245,N_14179,N_12312);
or U18246 (N_18246,N_13310,N_12111);
and U18247 (N_18247,N_14606,N_13932);
nand U18248 (N_18248,N_12137,N_10128);
and U18249 (N_18249,N_13655,N_11014);
nand U18250 (N_18250,N_13383,N_14026);
nand U18251 (N_18251,N_12857,N_14060);
nand U18252 (N_18252,N_12559,N_14273);
or U18253 (N_18253,N_12085,N_14836);
nand U18254 (N_18254,N_14533,N_14718);
nand U18255 (N_18255,N_11758,N_14427);
and U18256 (N_18256,N_12226,N_10306);
xnor U18257 (N_18257,N_14394,N_14648);
nand U18258 (N_18258,N_13489,N_13274);
xor U18259 (N_18259,N_14851,N_14475);
xor U18260 (N_18260,N_10822,N_10930);
nand U18261 (N_18261,N_14078,N_12805);
xor U18262 (N_18262,N_10795,N_10834);
nand U18263 (N_18263,N_14090,N_13793);
nand U18264 (N_18264,N_10357,N_13850);
and U18265 (N_18265,N_14570,N_13687);
and U18266 (N_18266,N_14211,N_11584);
or U18267 (N_18267,N_10861,N_14927);
or U18268 (N_18268,N_13370,N_12295);
and U18269 (N_18269,N_10499,N_13333);
and U18270 (N_18270,N_11184,N_12948);
xor U18271 (N_18271,N_13114,N_10229);
and U18272 (N_18272,N_14239,N_12698);
nand U18273 (N_18273,N_10252,N_13580);
nand U18274 (N_18274,N_13496,N_11746);
nand U18275 (N_18275,N_10689,N_11205);
nand U18276 (N_18276,N_13003,N_12074);
nand U18277 (N_18277,N_13075,N_11697);
nor U18278 (N_18278,N_11108,N_10190);
nand U18279 (N_18279,N_12852,N_11732);
and U18280 (N_18280,N_12788,N_13957);
and U18281 (N_18281,N_10063,N_12992);
and U18282 (N_18282,N_14810,N_13669);
and U18283 (N_18283,N_10420,N_14131);
and U18284 (N_18284,N_12340,N_14777);
and U18285 (N_18285,N_12854,N_12219);
nand U18286 (N_18286,N_13260,N_10646);
nor U18287 (N_18287,N_11252,N_11068);
or U18288 (N_18288,N_11942,N_10718);
and U18289 (N_18289,N_13028,N_14016);
or U18290 (N_18290,N_11668,N_13133);
nand U18291 (N_18291,N_14052,N_13575);
nor U18292 (N_18292,N_12174,N_13978);
nand U18293 (N_18293,N_11799,N_11955);
xor U18294 (N_18294,N_12766,N_13541);
nor U18295 (N_18295,N_10649,N_12150);
xor U18296 (N_18296,N_11837,N_11733);
nor U18297 (N_18297,N_12646,N_14485);
and U18298 (N_18298,N_10793,N_10532);
and U18299 (N_18299,N_13279,N_11882);
xor U18300 (N_18300,N_11945,N_13525);
and U18301 (N_18301,N_13886,N_11574);
nand U18302 (N_18302,N_13312,N_12846);
nand U18303 (N_18303,N_11042,N_14327);
nor U18304 (N_18304,N_11756,N_13004);
xnor U18305 (N_18305,N_12539,N_11056);
nand U18306 (N_18306,N_11900,N_14188);
nor U18307 (N_18307,N_12518,N_14548);
and U18308 (N_18308,N_13924,N_10793);
nand U18309 (N_18309,N_11547,N_13297);
or U18310 (N_18310,N_11908,N_11666);
nor U18311 (N_18311,N_12769,N_10799);
nand U18312 (N_18312,N_11678,N_10262);
and U18313 (N_18313,N_13693,N_10530);
or U18314 (N_18314,N_10289,N_11365);
or U18315 (N_18315,N_12548,N_12119);
or U18316 (N_18316,N_13246,N_11137);
xnor U18317 (N_18317,N_13198,N_14165);
nand U18318 (N_18318,N_11866,N_12546);
and U18319 (N_18319,N_12187,N_12244);
or U18320 (N_18320,N_11775,N_10182);
or U18321 (N_18321,N_11274,N_11748);
or U18322 (N_18322,N_14317,N_13517);
or U18323 (N_18323,N_12078,N_14391);
nand U18324 (N_18324,N_10890,N_10566);
nor U18325 (N_18325,N_13774,N_14599);
and U18326 (N_18326,N_13002,N_13722);
and U18327 (N_18327,N_13465,N_14880);
nor U18328 (N_18328,N_10526,N_10749);
xor U18329 (N_18329,N_11890,N_14886);
nand U18330 (N_18330,N_11597,N_12583);
nor U18331 (N_18331,N_13642,N_12460);
and U18332 (N_18332,N_14719,N_13661);
and U18333 (N_18333,N_12604,N_12589);
nand U18334 (N_18334,N_12165,N_12932);
or U18335 (N_18335,N_11859,N_12204);
nor U18336 (N_18336,N_14289,N_10443);
and U18337 (N_18337,N_11761,N_12040);
nand U18338 (N_18338,N_10569,N_12656);
nor U18339 (N_18339,N_13928,N_14364);
xnor U18340 (N_18340,N_12287,N_11199);
or U18341 (N_18341,N_11254,N_13688);
nand U18342 (N_18342,N_14309,N_10816);
or U18343 (N_18343,N_12116,N_11643);
or U18344 (N_18344,N_12432,N_12456);
nor U18345 (N_18345,N_10940,N_14315);
nand U18346 (N_18346,N_13650,N_14576);
nand U18347 (N_18347,N_14680,N_10949);
xnor U18348 (N_18348,N_10852,N_10615);
or U18349 (N_18349,N_11094,N_11145);
nand U18350 (N_18350,N_13101,N_14022);
xor U18351 (N_18351,N_14462,N_12088);
or U18352 (N_18352,N_14908,N_12743);
and U18353 (N_18353,N_11844,N_10809);
nor U18354 (N_18354,N_13959,N_11784);
or U18355 (N_18355,N_12258,N_13446);
and U18356 (N_18356,N_13439,N_14857);
nor U18357 (N_18357,N_11294,N_11744);
or U18358 (N_18358,N_10346,N_10169);
xnor U18359 (N_18359,N_12851,N_13360);
nand U18360 (N_18360,N_11488,N_11449);
xnor U18361 (N_18361,N_11625,N_11909);
and U18362 (N_18362,N_14949,N_12023);
and U18363 (N_18363,N_12032,N_12228);
nor U18364 (N_18364,N_13632,N_10897);
and U18365 (N_18365,N_11452,N_11900);
nor U18366 (N_18366,N_13308,N_14178);
and U18367 (N_18367,N_10694,N_12202);
nand U18368 (N_18368,N_10132,N_12710);
nor U18369 (N_18369,N_14461,N_13827);
xnor U18370 (N_18370,N_13366,N_13173);
xor U18371 (N_18371,N_12380,N_11464);
xor U18372 (N_18372,N_13657,N_11520);
or U18373 (N_18373,N_12946,N_11830);
nor U18374 (N_18374,N_14653,N_11029);
or U18375 (N_18375,N_12274,N_11239);
or U18376 (N_18376,N_10590,N_14691);
or U18377 (N_18377,N_13031,N_13325);
nand U18378 (N_18378,N_13088,N_13186);
or U18379 (N_18379,N_12576,N_13256);
or U18380 (N_18380,N_14445,N_14918);
nand U18381 (N_18381,N_13471,N_10245);
nand U18382 (N_18382,N_10928,N_10345);
nor U18383 (N_18383,N_13391,N_11583);
nor U18384 (N_18384,N_11334,N_13569);
xor U18385 (N_18385,N_14382,N_14709);
xor U18386 (N_18386,N_10980,N_14401);
and U18387 (N_18387,N_12352,N_11103);
and U18388 (N_18388,N_14315,N_11277);
xnor U18389 (N_18389,N_14708,N_13930);
nor U18390 (N_18390,N_12922,N_11542);
xor U18391 (N_18391,N_14397,N_11705);
or U18392 (N_18392,N_11994,N_13483);
nand U18393 (N_18393,N_11398,N_12391);
xnor U18394 (N_18394,N_10325,N_14848);
and U18395 (N_18395,N_13871,N_10056);
or U18396 (N_18396,N_12720,N_14253);
and U18397 (N_18397,N_13541,N_13930);
or U18398 (N_18398,N_10955,N_12495);
nor U18399 (N_18399,N_11836,N_11307);
or U18400 (N_18400,N_10286,N_14245);
xnor U18401 (N_18401,N_12955,N_12976);
or U18402 (N_18402,N_11189,N_10088);
nand U18403 (N_18403,N_13092,N_10732);
or U18404 (N_18404,N_11859,N_14597);
or U18405 (N_18405,N_14440,N_14588);
or U18406 (N_18406,N_13837,N_11323);
nor U18407 (N_18407,N_10039,N_13152);
and U18408 (N_18408,N_14571,N_11393);
xor U18409 (N_18409,N_13537,N_11100);
xor U18410 (N_18410,N_14220,N_11703);
nand U18411 (N_18411,N_13008,N_14741);
xnor U18412 (N_18412,N_11605,N_11661);
xor U18413 (N_18413,N_11783,N_10549);
xor U18414 (N_18414,N_13018,N_12173);
and U18415 (N_18415,N_10511,N_10299);
or U18416 (N_18416,N_13589,N_10050);
nand U18417 (N_18417,N_13181,N_10652);
nand U18418 (N_18418,N_11683,N_14404);
and U18419 (N_18419,N_12277,N_10860);
xnor U18420 (N_18420,N_14354,N_11951);
or U18421 (N_18421,N_14503,N_14502);
nand U18422 (N_18422,N_12452,N_14129);
nor U18423 (N_18423,N_13222,N_10209);
and U18424 (N_18424,N_12565,N_13794);
nor U18425 (N_18425,N_14819,N_11499);
nor U18426 (N_18426,N_10786,N_10234);
xnor U18427 (N_18427,N_12152,N_11421);
or U18428 (N_18428,N_14009,N_11247);
or U18429 (N_18429,N_13538,N_13424);
nor U18430 (N_18430,N_11949,N_13121);
nand U18431 (N_18431,N_14047,N_13977);
nor U18432 (N_18432,N_11118,N_12916);
nand U18433 (N_18433,N_14700,N_14744);
and U18434 (N_18434,N_12513,N_13720);
nand U18435 (N_18435,N_12788,N_11649);
and U18436 (N_18436,N_13924,N_14862);
nor U18437 (N_18437,N_13107,N_10408);
and U18438 (N_18438,N_10491,N_13481);
and U18439 (N_18439,N_14217,N_13871);
xnor U18440 (N_18440,N_13980,N_13679);
nand U18441 (N_18441,N_12361,N_13985);
nand U18442 (N_18442,N_14643,N_14309);
xnor U18443 (N_18443,N_13280,N_14341);
nand U18444 (N_18444,N_11887,N_10130);
xnor U18445 (N_18445,N_14360,N_12529);
nor U18446 (N_18446,N_13140,N_13479);
xnor U18447 (N_18447,N_14919,N_10028);
nor U18448 (N_18448,N_14456,N_10529);
nor U18449 (N_18449,N_10521,N_11840);
xnor U18450 (N_18450,N_11167,N_11255);
and U18451 (N_18451,N_10524,N_14904);
xor U18452 (N_18452,N_14021,N_11637);
xor U18453 (N_18453,N_11903,N_11826);
nor U18454 (N_18454,N_12336,N_11033);
nor U18455 (N_18455,N_13473,N_14282);
or U18456 (N_18456,N_13502,N_10421);
and U18457 (N_18457,N_11386,N_14409);
nor U18458 (N_18458,N_12341,N_10916);
and U18459 (N_18459,N_13759,N_12958);
xor U18460 (N_18460,N_10504,N_10309);
nand U18461 (N_18461,N_10164,N_12329);
and U18462 (N_18462,N_10788,N_13955);
or U18463 (N_18463,N_13004,N_14756);
and U18464 (N_18464,N_14041,N_13021);
nor U18465 (N_18465,N_13275,N_11304);
xnor U18466 (N_18466,N_13917,N_11905);
nand U18467 (N_18467,N_11260,N_14382);
xnor U18468 (N_18468,N_12611,N_11619);
xnor U18469 (N_18469,N_14771,N_13743);
and U18470 (N_18470,N_12735,N_12099);
and U18471 (N_18471,N_10273,N_10869);
xnor U18472 (N_18472,N_12813,N_14674);
nand U18473 (N_18473,N_14103,N_13754);
nor U18474 (N_18474,N_12625,N_13471);
and U18475 (N_18475,N_12531,N_12204);
nand U18476 (N_18476,N_14458,N_13813);
xor U18477 (N_18477,N_14443,N_14381);
or U18478 (N_18478,N_10368,N_12738);
or U18479 (N_18479,N_10529,N_13091);
nor U18480 (N_18480,N_11577,N_14557);
nor U18481 (N_18481,N_14397,N_13801);
nand U18482 (N_18482,N_10485,N_11030);
nor U18483 (N_18483,N_12078,N_12658);
and U18484 (N_18484,N_14711,N_13035);
xnor U18485 (N_18485,N_12900,N_14079);
nand U18486 (N_18486,N_12021,N_11400);
nor U18487 (N_18487,N_13589,N_14095);
nand U18488 (N_18488,N_12475,N_11933);
or U18489 (N_18489,N_11399,N_13839);
or U18490 (N_18490,N_13132,N_11249);
xnor U18491 (N_18491,N_11177,N_12898);
and U18492 (N_18492,N_10598,N_10954);
xnor U18493 (N_18493,N_12793,N_11972);
nor U18494 (N_18494,N_12756,N_14300);
xor U18495 (N_18495,N_11676,N_14608);
nand U18496 (N_18496,N_14319,N_13364);
and U18497 (N_18497,N_14116,N_10025);
and U18498 (N_18498,N_11965,N_10111);
or U18499 (N_18499,N_11294,N_11341);
or U18500 (N_18500,N_11383,N_14301);
nor U18501 (N_18501,N_13182,N_10353);
xor U18502 (N_18502,N_11706,N_11028);
nand U18503 (N_18503,N_13058,N_11823);
nor U18504 (N_18504,N_11289,N_12764);
or U18505 (N_18505,N_11775,N_14241);
nor U18506 (N_18506,N_12433,N_13620);
nor U18507 (N_18507,N_11627,N_11484);
nor U18508 (N_18508,N_10917,N_14710);
nand U18509 (N_18509,N_11096,N_10643);
and U18510 (N_18510,N_13512,N_13575);
nor U18511 (N_18511,N_13082,N_14588);
and U18512 (N_18512,N_14059,N_10118);
and U18513 (N_18513,N_10302,N_12447);
and U18514 (N_18514,N_10610,N_14852);
and U18515 (N_18515,N_13270,N_12938);
nor U18516 (N_18516,N_11951,N_12676);
nand U18517 (N_18517,N_14007,N_13716);
nor U18518 (N_18518,N_12889,N_13999);
or U18519 (N_18519,N_13212,N_10671);
xor U18520 (N_18520,N_13517,N_14497);
nor U18521 (N_18521,N_12407,N_13713);
and U18522 (N_18522,N_12539,N_10065);
nand U18523 (N_18523,N_13547,N_12551);
nor U18524 (N_18524,N_13942,N_12463);
nor U18525 (N_18525,N_13605,N_12672);
or U18526 (N_18526,N_10588,N_12206);
nor U18527 (N_18527,N_14434,N_14048);
nor U18528 (N_18528,N_11574,N_12781);
nor U18529 (N_18529,N_12467,N_14677);
nor U18530 (N_18530,N_11448,N_14592);
or U18531 (N_18531,N_11636,N_12069);
and U18532 (N_18532,N_14925,N_14251);
or U18533 (N_18533,N_12846,N_13771);
nand U18534 (N_18534,N_10273,N_10112);
nor U18535 (N_18535,N_12116,N_12391);
xor U18536 (N_18536,N_10735,N_11260);
nand U18537 (N_18537,N_13287,N_12347);
or U18538 (N_18538,N_12062,N_13682);
nand U18539 (N_18539,N_13514,N_14836);
nand U18540 (N_18540,N_13910,N_11208);
or U18541 (N_18541,N_14874,N_10728);
xnor U18542 (N_18542,N_14813,N_10121);
nor U18543 (N_18543,N_13562,N_13918);
and U18544 (N_18544,N_12951,N_10331);
or U18545 (N_18545,N_14392,N_10495);
nand U18546 (N_18546,N_14957,N_14751);
and U18547 (N_18547,N_13565,N_11886);
nand U18548 (N_18548,N_10075,N_11494);
or U18549 (N_18549,N_14801,N_13952);
nand U18550 (N_18550,N_14412,N_12075);
and U18551 (N_18551,N_14427,N_10585);
or U18552 (N_18552,N_14644,N_14583);
nor U18553 (N_18553,N_14042,N_13474);
xnor U18554 (N_18554,N_14271,N_11221);
xor U18555 (N_18555,N_10086,N_12315);
and U18556 (N_18556,N_12389,N_11935);
or U18557 (N_18557,N_13293,N_12050);
or U18558 (N_18558,N_14693,N_13165);
and U18559 (N_18559,N_12536,N_12892);
or U18560 (N_18560,N_12751,N_10470);
or U18561 (N_18561,N_10716,N_10700);
nor U18562 (N_18562,N_12549,N_12229);
nand U18563 (N_18563,N_14254,N_14530);
and U18564 (N_18564,N_10616,N_11119);
nand U18565 (N_18565,N_14288,N_14749);
or U18566 (N_18566,N_11219,N_11352);
and U18567 (N_18567,N_13068,N_12332);
nor U18568 (N_18568,N_14928,N_14433);
or U18569 (N_18569,N_14355,N_13695);
and U18570 (N_18570,N_10945,N_12434);
nor U18571 (N_18571,N_13544,N_13883);
or U18572 (N_18572,N_12447,N_11336);
or U18573 (N_18573,N_12031,N_12702);
and U18574 (N_18574,N_12771,N_12541);
xnor U18575 (N_18575,N_11764,N_13816);
and U18576 (N_18576,N_11879,N_13134);
xnor U18577 (N_18577,N_12495,N_14737);
xor U18578 (N_18578,N_11096,N_12625);
xor U18579 (N_18579,N_14982,N_10909);
or U18580 (N_18580,N_10885,N_12576);
nand U18581 (N_18581,N_11447,N_14607);
and U18582 (N_18582,N_11237,N_14243);
or U18583 (N_18583,N_12555,N_13869);
nand U18584 (N_18584,N_11956,N_12993);
nor U18585 (N_18585,N_11697,N_10528);
xor U18586 (N_18586,N_13390,N_10886);
and U18587 (N_18587,N_14466,N_14503);
xor U18588 (N_18588,N_10691,N_10298);
or U18589 (N_18589,N_14672,N_14612);
nor U18590 (N_18590,N_13614,N_10422);
nor U18591 (N_18591,N_10513,N_13259);
nand U18592 (N_18592,N_13550,N_12837);
and U18593 (N_18593,N_13931,N_14246);
nand U18594 (N_18594,N_10770,N_10544);
or U18595 (N_18595,N_14482,N_14026);
nor U18596 (N_18596,N_10277,N_14897);
nand U18597 (N_18597,N_10886,N_10681);
xnor U18598 (N_18598,N_13102,N_14426);
nor U18599 (N_18599,N_10802,N_10359);
nand U18600 (N_18600,N_14561,N_12231);
xor U18601 (N_18601,N_10992,N_10687);
and U18602 (N_18602,N_14621,N_11885);
and U18603 (N_18603,N_13784,N_14068);
nor U18604 (N_18604,N_12410,N_12715);
and U18605 (N_18605,N_11132,N_12388);
nand U18606 (N_18606,N_14274,N_11880);
or U18607 (N_18607,N_11515,N_12240);
xor U18608 (N_18608,N_13430,N_11969);
or U18609 (N_18609,N_12924,N_10262);
nor U18610 (N_18610,N_14786,N_11145);
and U18611 (N_18611,N_12779,N_10038);
nor U18612 (N_18612,N_14783,N_11774);
or U18613 (N_18613,N_13563,N_10934);
or U18614 (N_18614,N_12469,N_11352);
or U18615 (N_18615,N_14573,N_10913);
nand U18616 (N_18616,N_11533,N_14574);
and U18617 (N_18617,N_11744,N_14798);
nand U18618 (N_18618,N_11516,N_11465);
xnor U18619 (N_18619,N_11527,N_13757);
nand U18620 (N_18620,N_12712,N_10679);
nor U18621 (N_18621,N_11556,N_14625);
nand U18622 (N_18622,N_11073,N_13914);
nand U18623 (N_18623,N_11321,N_14404);
and U18624 (N_18624,N_10150,N_12310);
and U18625 (N_18625,N_14095,N_11889);
or U18626 (N_18626,N_13981,N_12020);
xnor U18627 (N_18627,N_13294,N_13819);
and U18628 (N_18628,N_12928,N_11241);
and U18629 (N_18629,N_11960,N_12822);
nand U18630 (N_18630,N_11313,N_13963);
nand U18631 (N_18631,N_11073,N_14119);
xor U18632 (N_18632,N_12956,N_14253);
or U18633 (N_18633,N_11454,N_12162);
xor U18634 (N_18634,N_14055,N_14831);
nand U18635 (N_18635,N_12931,N_11165);
nand U18636 (N_18636,N_14388,N_14426);
and U18637 (N_18637,N_11430,N_11017);
and U18638 (N_18638,N_13226,N_12862);
nand U18639 (N_18639,N_13994,N_13259);
nor U18640 (N_18640,N_14404,N_13879);
nor U18641 (N_18641,N_10065,N_11391);
nor U18642 (N_18642,N_10788,N_14409);
and U18643 (N_18643,N_13866,N_10524);
nor U18644 (N_18644,N_12160,N_12705);
xor U18645 (N_18645,N_12172,N_12383);
nand U18646 (N_18646,N_10717,N_11258);
and U18647 (N_18647,N_14242,N_14576);
nor U18648 (N_18648,N_11631,N_10000);
and U18649 (N_18649,N_11592,N_11038);
and U18650 (N_18650,N_13237,N_14160);
nand U18651 (N_18651,N_14626,N_10875);
nand U18652 (N_18652,N_13146,N_14298);
and U18653 (N_18653,N_12945,N_14182);
nand U18654 (N_18654,N_10430,N_11246);
or U18655 (N_18655,N_10795,N_10946);
xnor U18656 (N_18656,N_14332,N_14988);
or U18657 (N_18657,N_13994,N_12819);
nor U18658 (N_18658,N_13083,N_10033);
xor U18659 (N_18659,N_11420,N_10346);
xnor U18660 (N_18660,N_10897,N_12719);
and U18661 (N_18661,N_11257,N_14533);
and U18662 (N_18662,N_13286,N_10724);
nand U18663 (N_18663,N_13745,N_13140);
nor U18664 (N_18664,N_11902,N_10990);
and U18665 (N_18665,N_13842,N_11106);
or U18666 (N_18666,N_12757,N_12185);
xnor U18667 (N_18667,N_10570,N_10502);
nand U18668 (N_18668,N_14764,N_12772);
nand U18669 (N_18669,N_12882,N_10086);
nor U18670 (N_18670,N_10906,N_12894);
or U18671 (N_18671,N_10918,N_11616);
or U18672 (N_18672,N_10459,N_13180);
nand U18673 (N_18673,N_11293,N_13817);
nor U18674 (N_18674,N_11520,N_12119);
and U18675 (N_18675,N_14782,N_11067);
and U18676 (N_18676,N_14201,N_11352);
nand U18677 (N_18677,N_11373,N_10902);
and U18678 (N_18678,N_13682,N_12428);
or U18679 (N_18679,N_14735,N_13529);
and U18680 (N_18680,N_12645,N_12686);
or U18681 (N_18681,N_13982,N_12432);
and U18682 (N_18682,N_14897,N_11608);
nor U18683 (N_18683,N_12703,N_13587);
nand U18684 (N_18684,N_14983,N_12157);
nor U18685 (N_18685,N_10495,N_10853);
nor U18686 (N_18686,N_11761,N_12173);
nand U18687 (N_18687,N_11303,N_10172);
nand U18688 (N_18688,N_10116,N_14844);
nand U18689 (N_18689,N_13068,N_13792);
or U18690 (N_18690,N_12978,N_10738);
xor U18691 (N_18691,N_10314,N_12458);
nand U18692 (N_18692,N_14362,N_11461);
or U18693 (N_18693,N_11495,N_14806);
or U18694 (N_18694,N_14261,N_11210);
or U18695 (N_18695,N_12013,N_14326);
xnor U18696 (N_18696,N_11302,N_12298);
nand U18697 (N_18697,N_14165,N_12346);
nor U18698 (N_18698,N_10950,N_13668);
nor U18699 (N_18699,N_12812,N_14788);
and U18700 (N_18700,N_14812,N_11878);
nor U18701 (N_18701,N_14333,N_10949);
and U18702 (N_18702,N_10830,N_13036);
nor U18703 (N_18703,N_13214,N_11393);
nand U18704 (N_18704,N_12289,N_13424);
nand U18705 (N_18705,N_11586,N_13879);
nor U18706 (N_18706,N_14370,N_11545);
and U18707 (N_18707,N_10847,N_10517);
and U18708 (N_18708,N_11678,N_12046);
nor U18709 (N_18709,N_11429,N_10793);
nor U18710 (N_18710,N_14077,N_12842);
nand U18711 (N_18711,N_13643,N_12539);
xor U18712 (N_18712,N_14431,N_14722);
xor U18713 (N_18713,N_14827,N_13390);
and U18714 (N_18714,N_11134,N_14059);
nor U18715 (N_18715,N_10896,N_14083);
nor U18716 (N_18716,N_10858,N_14451);
or U18717 (N_18717,N_14408,N_14006);
xnor U18718 (N_18718,N_11534,N_10787);
xnor U18719 (N_18719,N_12891,N_13968);
xnor U18720 (N_18720,N_11767,N_11534);
and U18721 (N_18721,N_13318,N_13008);
and U18722 (N_18722,N_10724,N_11891);
or U18723 (N_18723,N_12176,N_14509);
or U18724 (N_18724,N_11211,N_12918);
xnor U18725 (N_18725,N_11689,N_13988);
and U18726 (N_18726,N_11866,N_13066);
and U18727 (N_18727,N_12772,N_10388);
xnor U18728 (N_18728,N_14898,N_11755);
nand U18729 (N_18729,N_14539,N_14924);
nand U18730 (N_18730,N_14219,N_10976);
nor U18731 (N_18731,N_11732,N_12006);
and U18732 (N_18732,N_10429,N_14458);
xnor U18733 (N_18733,N_10010,N_11513);
and U18734 (N_18734,N_10036,N_12862);
nand U18735 (N_18735,N_13657,N_14256);
nand U18736 (N_18736,N_14103,N_11971);
nor U18737 (N_18737,N_10551,N_10667);
or U18738 (N_18738,N_10837,N_10232);
xor U18739 (N_18739,N_10213,N_13306);
nand U18740 (N_18740,N_10291,N_11750);
or U18741 (N_18741,N_12852,N_11878);
or U18742 (N_18742,N_10981,N_11747);
nand U18743 (N_18743,N_12022,N_13737);
nor U18744 (N_18744,N_14929,N_14144);
nand U18745 (N_18745,N_14630,N_10407);
nor U18746 (N_18746,N_12028,N_14759);
or U18747 (N_18747,N_11214,N_14118);
xor U18748 (N_18748,N_12110,N_12366);
and U18749 (N_18749,N_11354,N_14351);
nand U18750 (N_18750,N_12370,N_13720);
nand U18751 (N_18751,N_10893,N_13390);
nand U18752 (N_18752,N_13620,N_13869);
nor U18753 (N_18753,N_14016,N_13212);
and U18754 (N_18754,N_11857,N_11011);
nand U18755 (N_18755,N_13381,N_14593);
nor U18756 (N_18756,N_11028,N_10735);
xnor U18757 (N_18757,N_14828,N_14922);
nor U18758 (N_18758,N_10306,N_12474);
nand U18759 (N_18759,N_13929,N_10217);
or U18760 (N_18760,N_11236,N_14445);
nor U18761 (N_18761,N_14329,N_13501);
and U18762 (N_18762,N_13851,N_11874);
nand U18763 (N_18763,N_13245,N_14592);
nand U18764 (N_18764,N_12814,N_13866);
xnor U18765 (N_18765,N_13052,N_12586);
xnor U18766 (N_18766,N_12098,N_11731);
nor U18767 (N_18767,N_12610,N_11471);
xnor U18768 (N_18768,N_13614,N_12956);
nor U18769 (N_18769,N_13835,N_14432);
nand U18770 (N_18770,N_14883,N_12987);
or U18771 (N_18771,N_13902,N_10830);
nand U18772 (N_18772,N_11973,N_14300);
or U18773 (N_18773,N_10335,N_14623);
nor U18774 (N_18774,N_12845,N_14046);
nand U18775 (N_18775,N_10585,N_13247);
nor U18776 (N_18776,N_12196,N_14310);
nor U18777 (N_18777,N_11893,N_14872);
and U18778 (N_18778,N_14782,N_11833);
and U18779 (N_18779,N_13635,N_11791);
and U18780 (N_18780,N_14842,N_13465);
and U18781 (N_18781,N_10701,N_14239);
and U18782 (N_18782,N_10628,N_13370);
or U18783 (N_18783,N_14797,N_11624);
xnor U18784 (N_18784,N_14720,N_14541);
xor U18785 (N_18785,N_10975,N_13272);
nor U18786 (N_18786,N_11939,N_11629);
nor U18787 (N_18787,N_14445,N_12824);
and U18788 (N_18788,N_11665,N_13640);
or U18789 (N_18789,N_10226,N_11272);
and U18790 (N_18790,N_11824,N_13136);
or U18791 (N_18791,N_11627,N_12888);
nand U18792 (N_18792,N_11997,N_14750);
xnor U18793 (N_18793,N_11270,N_10179);
nand U18794 (N_18794,N_11108,N_11975);
nand U18795 (N_18795,N_13805,N_11897);
nand U18796 (N_18796,N_13694,N_10536);
or U18797 (N_18797,N_10900,N_13787);
and U18798 (N_18798,N_11631,N_13953);
and U18799 (N_18799,N_10171,N_14002);
xnor U18800 (N_18800,N_12523,N_12234);
or U18801 (N_18801,N_12483,N_11429);
and U18802 (N_18802,N_10965,N_12794);
or U18803 (N_18803,N_11183,N_13417);
nor U18804 (N_18804,N_11829,N_12102);
xor U18805 (N_18805,N_13242,N_12921);
nand U18806 (N_18806,N_10772,N_11018);
nor U18807 (N_18807,N_13737,N_14539);
or U18808 (N_18808,N_12416,N_13287);
or U18809 (N_18809,N_11764,N_13237);
nor U18810 (N_18810,N_10857,N_13749);
xor U18811 (N_18811,N_13171,N_10224);
nor U18812 (N_18812,N_13408,N_12963);
xnor U18813 (N_18813,N_14151,N_13354);
or U18814 (N_18814,N_13462,N_11470);
nand U18815 (N_18815,N_12613,N_13282);
or U18816 (N_18816,N_14364,N_13155);
nand U18817 (N_18817,N_14822,N_10649);
nand U18818 (N_18818,N_14017,N_10335);
and U18819 (N_18819,N_10952,N_14681);
nand U18820 (N_18820,N_13070,N_13670);
and U18821 (N_18821,N_11840,N_10981);
nor U18822 (N_18822,N_10561,N_14500);
xnor U18823 (N_18823,N_13190,N_11699);
nand U18824 (N_18824,N_13668,N_10360);
nor U18825 (N_18825,N_14992,N_14787);
xnor U18826 (N_18826,N_11609,N_13867);
nand U18827 (N_18827,N_12215,N_11176);
nand U18828 (N_18828,N_12659,N_11085);
nor U18829 (N_18829,N_14617,N_14149);
or U18830 (N_18830,N_10791,N_13937);
or U18831 (N_18831,N_13400,N_10486);
and U18832 (N_18832,N_14818,N_10861);
or U18833 (N_18833,N_12636,N_13008);
nand U18834 (N_18834,N_13933,N_14871);
and U18835 (N_18835,N_14030,N_10088);
and U18836 (N_18836,N_12385,N_13880);
nand U18837 (N_18837,N_11695,N_10703);
nor U18838 (N_18838,N_12357,N_10278);
xor U18839 (N_18839,N_14891,N_10030);
or U18840 (N_18840,N_10105,N_12404);
or U18841 (N_18841,N_11492,N_13581);
nor U18842 (N_18842,N_12922,N_12603);
nand U18843 (N_18843,N_14752,N_12246);
nor U18844 (N_18844,N_11339,N_11036);
and U18845 (N_18845,N_14639,N_10241);
and U18846 (N_18846,N_12781,N_12473);
nor U18847 (N_18847,N_13225,N_14566);
and U18848 (N_18848,N_13904,N_14877);
and U18849 (N_18849,N_14574,N_13112);
xnor U18850 (N_18850,N_12728,N_10602);
nand U18851 (N_18851,N_11782,N_11148);
xor U18852 (N_18852,N_11452,N_11095);
and U18853 (N_18853,N_14216,N_11756);
nor U18854 (N_18854,N_12613,N_13729);
nand U18855 (N_18855,N_13050,N_11101);
nand U18856 (N_18856,N_10059,N_13907);
nor U18857 (N_18857,N_13744,N_11643);
and U18858 (N_18858,N_14454,N_12302);
or U18859 (N_18859,N_11502,N_10499);
and U18860 (N_18860,N_12959,N_11164);
or U18861 (N_18861,N_13264,N_11425);
nor U18862 (N_18862,N_10618,N_13277);
nand U18863 (N_18863,N_11764,N_10422);
nor U18864 (N_18864,N_13650,N_12394);
nor U18865 (N_18865,N_14757,N_13573);
xor U18866 (N_18866,N_11999,N_12367);
nor U18867 (N_18867,N_14807,N_12128);
nor U18868 (N_18868,N_10278,N_10216);
nor U18869 (N_18869,N_14828,N_14860);
nor U18870 (N_18870,N_13462,N_12449);
nor U18871 (N_18871,N_13327,N_14124);
xor U18872 (N_18872,N_14664,N_13353);
and U18873 (N_18873,N_14541,N_13241);
xnor U18874 (N_18874,N_14271,N_12272);
xnor U18875 (N_18875,N_12928,N_14573);
and U18876 (N_18876,N_11903,N_14568);
and U18877 (N_18877,N_10579,N_11971);
or U18878 (N_18878,N_13964,N_11663);
and U18879 (N_18879,N_11196,N_10390);
or U18880 (N_18880,N_11162,N_12594);
or U18881 (N_18881,N_12166,N_10757);
or U18882 (N_18882,N_12910,N_10286);
and U18883 (N_18883,N_11470,N_12315);
nand U18884 (N_18884,N_13412,N_11621);
or U18885 (N_18885,N_11324,N_14686);
or U18886 (N_18886,N_13955,N_11112);
nor U18887 (N_18887,N_11771,N_10537);
nand U18888 (N_18888,N_11253,N_14592);
xnor U18889 (N_18889,N_14756,N_11326);
nand U18890 (N_18890,N_13891,N_13053);
or U18891 (N_18891,N_14997,N_10531);
nand U18892 (N_18892,N_14175,N_14549);
or U18893 (N_18893,N_10236,N_13373);
or U18894 (N_18894,N_12728,N_13489);
and U18895 (N_18895,N_12207,N_11345);
nor U18896 (N_18896,N_10721,N_13506);
xnor U18897 (N_18897,N_10216,N_11333);
xnor U18898 (N_18898,N_12927,N_14586);
nand U18899 (N_18899,N_14593,N_14988);
and U18900 (N_18900,N_11063,N_12499);
and U18901 (N_18901,N_11884,N_11702);
or U18902 (N_18902,N_12062,N_12426);
and U18903 (N_18903,N_12940,N_13296);
or U18904 (N_18904,N_11174,N_11533);
nor U18905 (N_18905,N_14025,N_11221);
or U18906 (N_18906,N_10724,N_13676);
nand U18907 (N_18907,N_13607,N_10566);
nand U18908 (N_18908,N_14774,N_12843);
nor U18909 (N_18909,N_14772,N_11855);
xor U18910 (N_18910,N_11745,N_13574);
xnor U18911 (N_18911,N_14588,N_10429);
xnor U18912 (N_18912,N_11358,N_10524);
nand U18913 (N_18913,N_13522,N_10715);
nor U18914 (N_18914,N_10102,N_10390);
nor U18915 (N_18915,N_14547,N_13671);
xnor U18916 (N_18916,N_12948,N_11363);
or U18917 (N_18917,N_14542,N_13660);
or U18918 (N_18918,N_14507,N_11683);
and U18919 (N_18919,N_14858,N_14575);
and U18920 (N_18920,N_12962,N_13480);
and U18921 (N_18921,N_14317,N_12272);
xor U18922 (N_18922,N_11087,N_10271);
and U18923 (N_18923,N_14150,N_14499);
nand U18924 (N_18924,N_12555,N_10811);
nor U18925 (N_18925,N_13854,N_11718);
nor U18926 (N_18926,N_10577,N_12777);
nor U18927 (N_18927,N_11762,N_11864);
or U18928 (N_18928,N_12327,N_10490);
nand U18929 (N_18929,N_11392,N_11110);
nand U18930 (N_18930,N_10157,N_14340);
and U18931 (N_18931,N_12487,N_14256);
xnor U18932 (N_18932,N_10644,N_10353);
or U18933 (N_18933,N_13463,N_10045);
nand U18934 (N_18934,N_12446,N_10962);
xor U18935 (N_18935,N_11697,N_14487);
nor U18936 (N_18936,N_12567,N_10666);
and U18937 (N_18937,N_12658,N_12364);
xor U18938 (N_18938,N_12043,N_13789);
nand U18939 (N_18939,N_14305,N_11333);
nor U18940 (N_18940,N_14858,N_11511);
and U18941 (N_18941,N_12530,N_10286);
xor U18942 (N_18942,N_14263,N_12923);
xor U18943 (N_18943,N_10636,N_13040);
and U18944 (N_18944,N_10861,N_14085);
or U18945 (N_18945,N_14005,N_10623);
nand U18946 (N_18946,N_13408,N_12953);
xor U18947 (N_18947,N_12047,N_11643);
or U18948 (N_18948,N_13927,N_11377);
or U18949 (N_18949,N_13669,N_13735);
nor U18950 (N_18950,N_13817,N_13409);
and U18951 (N_18951,N_14309,N_14745);
xnor U18952 (N_18952,N_13466,N_13819);
or U18953 (N_18953,N_14518,N_14393);
nand U18954 (N_18954,N_12393,N_13583);
or U18955 (N_18955,N_11750,N_14620);
xor U18956 (N_18956,N_10735,N_13538);
nand U18957 (N_18957,N_14720,N_14512);
and U18958 (N_18958,N_13812,N_10077);
nor U18959 (N_18959,N_12346,N_13115);
and U18960 (N_18960,N_14495,N_14532);
and U18961 (N_18961,N_12126,N_13153);
xor U18962 (N_18962,N_13617,N_14041);
xor U18963 (N_18963,N_11669,N_11543);
nand U18964 (N_18964,N_10580,N_12016);
or U18965 (N_18965,N_12366,N_11023);
nand U18966 (N_18966,N_10240,N_14438);
xor U18967 (N_18967,N_10377,N_14311);
or U18968 (N_18968,N_11593,N_11245);
and U18969 (N_18969,N_10155,N_11953);
nand U18970 (N_18970,N_10014,N_10612);
nor U18971 (N_18971,N_14419,N_14045);
or U18972 (N_18972,N_12133,N_11578);
nand U18973 (N_18973,N_10933,N_13064);
and U18974 (N_18974,N_14918,N_13381);
xor U18975 (N_18975,N_14849,N_12024);
xor U18976 (N_18976,N_13694,N_10640);
xor U18977 (N_18977,N_13042,N_14689);
or U18978 (N_18978,N_12673,N_14302);
nor U18979 (N_18979,N_12984,N_14053);
xor U18980 (N_18980,N_11931,N_12457);
or U18981 (N_18981,N_12463,N_14890);
nand U18982 (N_18982,N_11575,N_14938);
and U18983 (N_18983,N_14032,N_13969);
or U18984 (N_18984,N_11533,N_11325);
xor U18985 (N_18985,N_11146,N_10497);
nand U18986 (N_18986,N_11517,N_10366);
nand U18987 (N_18987,N_10076,N_11866);
and U18988 (N_18988,N_10540,N_11541);
nand U18989 (N_18989,N_14429,N_14672);
nand U18990 (N_18990,N_12622,N_14601);
xnor U18991 (N_18991,N_10182,N_12827);
and U18992 (N_18992,N_11764,N_11288);
nand U18993 (N_18993,N_11585,N_10414);
nand U18994 (N_18994,N_12112,N_12971);
or U18995 (N_18995,N_12326,N_13506);
xor U18996 (N_18996,N_10883,N_14815);
and U18997 (N_18997,N_11538,N_11505);
nor U18998 (N_18998,N_10972,N_10414);
or U18999 (N_18999,N_13099,N_12238);
nand U19000 (N_19000,N_14600,N_12794);
nor U19001 (N_19001,N_13839,N_12138);
nor U19002 (N_19002,N_12937,N_14085);
nand U19003 (N_19003,N_13185,N_12910);
and U19004 (N_19004,N_14133,N_14645);
and U19005 (N_19005,N_11421,N_12384);
or U19006 (N_19006,N_14245,N_10326);
xnor U19007 (N_19007,N_11156,N_12765);
nor U19008 (N_19008,N_11212,N_13203);
nand U19009 (N_19009,N_13394,N_14389);
and U19010 (N_19010,N_11048,N_13402);
and U19011 (N_19011,N_10721,N_14716);
nand U19012 (N_19012,N_13226,N_13421);
and U19013 (N_19013,N_10039,N_12780);
nand U19014 (N_19014,N_10692,N_14802);
or U19015 (N_19015,N_13041,N_11462);
xor U19016 (N_19016,N_12994,N_13002);
nor U19017 (N_19017,N_14413,N_14307);
nand U19018 (N_19018,N_10674,N_12021);
nand U19019 (N_19019,N_12242,N_12623);
nand U19020 (N_19020,N_10225,N_14257);
and U19021 (N_19021,N_12139,N_11723);
nor U19022 (N_19022,N_14166,N_13267);
nor U19023 (N_19023,N_13937,N_14444);
nand U19024 (N_19024,N_12055,N_14291);
nand U19025 (N_19025,N_11687,N_13168);
or U19026 (N_19026,N_14840,N_12770);
nor U19027 (N_19027,N_14234,N_11056);
nor U19028 (N_19028,N_12250,N_12240);
or U19029 (N_19029,N_14146,N_13381);
nor U19030 (N_19030,N_11685,N_10336);
and U19031 (N_19031,N_11848,N_14035);
nand U19032 (N_19032,N_11891,N_11058);
xnor U19033 (N_19033,N_11585,N_14399);
and U19034 (N_19034,N_12989,N_14383);
xor U19035 (N_19035,N_11746,N_11986);
nand U19036 (N_19036,N_13294,N_13890);
nor U19037 (N_19037,N_12915,N_10235);
and U19038 (N_19038,N_14256,N_13120);
nand U19039 (N_19039,N_14476,N_13587);
xnor U19040 (N_19040,N_10999,N_10273);
and U19041 (N_19041,N_13541,N_12894);
nor U19042 (N_19042,N_11345,N_14283);
xor U19043 (N_19043,N_13461,N_10129);
and U19044 (N_19044,N_14578,N_14560);
xor U19045 (N_19045,N_12339,N_13301);
and U19046 (N_19046,N_10358,N_12189);
and U19047 (N_19047,N_12137,N_13600);
and U19048 (N_19048,N_12368,N_11360);
nand U19049 (N_19049,N_11303,N_14271);
xor U19050 (N_19050,N_10171,N_11529);
xnor U19051 (N_19051,N_11842,N_10270);
nor U19052 (N_19052,N_10614,N_14777);
nor U19053 (N_19053,N_13653,N_11423);
and U19054 (N_19054,N_11886,N_14861);
nand U19055 (N_19055,N_13784,N_10583);
and U19056 (N_19056,N_13213,N_10833);
and U19057 (N_19057,N_12267,N_12034);
and U19058 (N_19058,N_12466,N_14278);
nand U19059 (N_19059,N_14728,N_14758);
xnor U19060 (N_19060,N_14317,N_13729);
nand U19061 (N_19061,N_13004,N_11967);
nor U19062 (N_19062,N_11065,N_12292);
and U19063 (N_19063,N_13928,N_11158);
xnor U19064 (N_19064,N_13638,N_11876);
or U19065 (N_19065,N_13184,N_12240);
or U19066 (N_19066,N_12351,N_13070);
nand U19067 (N_19067,N_11563,N_12741);
and U19068 (N_19068,N_12717,N_10472);
xor U19069 (N_19069,N_10326,N_13932);
xnor U19070 (N_19070,N_12135,N_11533);
xnor U19071 (N_19071,N_14097,N_14336);
nand U19072 (N_19072,N_14945,N_11753);
or U19073 (N_19073,N_13022,N_11731);
or U19074 (N_19074,N_14882,N_10477);
xor U19075 (N_19075,N_14599,N_14930);
or U19076 (N_19076,N_12686,N_14477);
and U19077 (N_19077,N_14494,N_14605);
or U19078 (N_19078,N_13435,N_13680);
or U19079 (N_19079,N_12113,N_11353);
xnor U19080 (N_19080,N_10204,N_12535);
and U19081 (N_19081,N_11363,N_13928);
nor U19082 (N_19082,N_12346,N_10780);
nor U19083 (N_19083,N_10644,N_13159);
nand U19084 (N_19084,N_12251,N_12198);
nor U19085 (N_19085,N_11241,N_10996);
nor U19086 (N_19086,N_14079,N_10102);
nand U19087 (N_19087,N_14524,N_10098);
nor U19088 (N_19088,N_12328,N_11791);
nand U19089 (N_19089,N_13188,N_13587);
or U19090 (N_19090,N_14682,N_13579);
nand U19091 (N_19091,N_12395,N_10266);
nor U19092 (N_19092,N_14138,N_14190);
nor U19093 (N_19093,N_13470,N_11598);
nand U19094 (N_19094,N_10595,N_14368);
or U19095 (N_19095,N_12738,N_11620);
and U19096 (N_19096,N_12476,N_14377);
or U19097 (N_19097,N_14831,N_11201);
nor U19098 (N_19098,N_13141,N_12015);
xnor U19099 (N_19099,N_13897,N_13884);
xnor U19100 (N_19100,N_11334,N_14924);
nand U19101 (N_19101,N_10149,N_13623);
xor U19102 (N_19102,N_14633,N_14024);
nor U19103 (N_19103,N_13648,N_12049);
nand U19104 (N_19104,N_10375,N_13216);
xnor U19105 (N_19105,N_11764,N_11240);
nand U19106 (N_19106,N_10594,N_10399);
and U19107 (N_19107,N_11818,N_14085);
xor U19108 (N_19108,N_13890,N_12389);
xor U19109 (N_19109,N_10988,N_11968);
nand U19110 (N_19110,N_13478,N_12151);
nor U19111 (N_19111,N_12775,N_11471);
nor U19112 (N_19112,N_12928,N_13340);
nand U19113 (N_19113,N_14597,N_13029);
and U19114 (N_19114,N_11966,N_13643);
and U19115 (N_19115,N_12031,N_13300);
nor U19116 (N_19116,N_10961,N_13523);
xor U19117 (N_19117,N_12593,N_10189);
xnor U19118 (N_19118,N_13094,N_13424);
or U19119 (N_19119,N_14581,N_13889);
nor U19120 (N_19120,N_14371,N_13622);
or U19121 (N_19121,N_13717,N_10742);
and U19122 (N_19122,N_12378,N_11977);
and U19123 (N_19123,N_10824,N_10769);
and U19124 (N_19124,N_13557,N_12461);
xor U19125 (N_19125,N_12746,N_14453);
nand U19126 (N_19126,N_13375,N_13796);
or U19127 (N_19127,N_14624,N_11196);
and U19128 (N_19128,N_13360,N_13911);
xnor U19129 (N_19129,N_14079,N_11343);
or U19130 (N_19130,N_13949,N_10134);
nor U19131 (N_19131,N_13203,N_13220);
nand U19132 (N_19132,N_10422,N_11827);
nand U19133 (N_19133,N_13232,N_12795);
xnor U19134 (N_19134,N_12056,N_13920);
xnor U19135 (N_19135,N_12109,N_12591);
or U19136 (N_19136,N_11074,N_10233);
nand U19137 (N_19137,N_13732,N_12073);
xor U19138 (N_19138,N_13093,N_13033);
nand U19139 (N_19139,N_13900,N_13787);
nor U19140 (N_19140,N_12646,N_13290);
or U19141 (N_19141,N_14366,N_14035);
or U19142 (N_19142,N_11509,N_10845);
nor U19143 (N_19143,N_10016,N_10325);
and U19144 (N_19144,N_10747,N_11092);
xnor U19145 (N_19145,N_10664,N_13955);
or U19146 (N_19146,N_10199,N_11985);
or U19147 (N_19147,N_11984,N_13662);
xnor U19148 (N_19148,N_11288,N_10426);
and U19149 (N_19149,N_10184,N_14293);
and U19150 (N_19150,N_14056,N_14976);
or U19151 (N_19151,N_10163,N_10287);
nor U19152 (N_19152,N_13260,N_14002);
and U19153 (N_19153,N_13593,N_12794);
or U19154 (N_19154,N_14071,N_13200);
xnor U19155 (N_19155,N_10181,N_11565);
nand U19156 (N_19156,N_13584,N_12779);
xor U19157 (N_19157,N_13182,N_14460);
and U19158 (N_19158,N_10453,N_11944);
nand U19159 (N_19159,N_12067,N_14649);
xor U19160 (N_19160,N_13595,N_10902);
xnor U19161 (N_19161,N_12729,N_10356);
nor U19162 (N_19162,N_10604,N_12956);
nor U19163 (N_19163,N_11376,N_11513);
nor U19164 (N_19164,N_14933,N_14075);
xor U19165 (N_19165,N_12827,N_13366);
xor U19166 (N_19166,N_11822,N_14270);
xnor U19167 (N_19167,N_12834,N_12351);
nand U19168 (N_19168,N_11688,N_14275);
nor U19169 (N_19169,N_11417,N_13521);
nor U19170 (N_19170,N_14278,N_12485);
xnor U19171 (N_19171,N_12066,N_13761);
nor U19172 (N_19172,N_13269,N_13879);
nand U19173 (N_19173,N_14273,N_14507);
or U19174 (N_19174,N_10852,N_14209);
xor U19175 (N_19175,N_13965,N_12556);
nor U19176 (N_19176,N_10970,N_11149);
xor U19177 (N_19177,N_14270,N_14757);
xnor U19178 (N_19178,N_14000,N_13280);
or U19179 (N_19179,N_13029,N_13091);
nor U19180 (N_19180,N_12492,N_12814);
and U19181 (N_19181,N_13824,N_13473);
nand U19182 (N_19182,N_11058,N_10762);
xor U19183 (N_19183,N_14721,N_13832);
nor U19184 (N_19184,N_12281,N_11831);
xor U19185 (N_19185,N_13130,N_13036);
and U19186 (N_19186,N_13130,N_14719);
xnor U19187 (N_19187,N_14877,N_12325);
nand U19188 (N_19188,N_13202,N_14214);
nand U19189 (N_19189,N_14488,N_12124);
or U19190 (N_19190,N_11429,N_11953);
xnor U19191 (N_19191,N_13220,N_11311);
nor U19192 (N_19192,N_13382,N_13095);
xnor U19193 (N_19193,N_13653,N_11067);
nor U19194 (N_19194,N_14265,N_10414);
or U19195 (N_19195,N_12526,N_12210);
xor U19196 (N_19196,N_10053,N_12272);
nand U19197 (N_19197,N_10263,N_10881);
nor U19198 (N_19198,N_13635,N_10878);
xnor U19199 (N_19199,N_10454,N_14418);
and U19200 (N_19200,N_14465,N_10980);
or U19201 (N_19201,N_10294,N_12529);
and U19202 (N_19202,N_13828,N_10934);
nor U19203 (N_19203,N_11496,N_13654);
and U19204 (N_19204,N_13433,N_11310);
or U19205 (N_19205,N_14026,N_14295);
or U19206 (N_19206,N_10559,N_10706);
and U19207 (N_19207,N_10331,N_14985);
or U19208 (N_19208,N_14858,N_14593);
and U19209 (N_19209,N_13447,N_13394);
nor U19210 (N_19210,N_13191,N_10245);
nand U19211 (N_19211,N_13528,N_10398);
and U19212 (N_19212,N_14460,N_13689);
and U19213 (N_19213,N_12430,N_13768);
or U19214 (N_19214,N_14511,N_12093);
nor U19215 (N_19215,N_13184,N_13139);
or U19216 (N_19216,N_13119,N_11447);
xor U19217 (N_19217,N_11786,N_12121);
nor U19218 (N_19218,N_14064,N_13389);
or U19219 (N_19219,N_14616,N_12480);
and U19220 (N_19220,N_11596,N_10405);
or U19221 (N_19221,N_13264,N_10826);
or U19222 (N_19222,N_14821,N_11375);
nor U19223 (N_19223,N_11658,N_14646);
and U19224 (N_19224,N_10990,N_11986);
or U19225 (N_19225,N_11763,N_13731);
and U19226 (N_19226,N_12725,N_11951);
xor U19227 (N_19227,N_14750,N_14769);
nor U19228 (N_19228,N_13112,N_10076);
or U19229 (N_19229,N_10721,N_10225);
nor U19230 (N_19230,N_10511,N_12309);
nand U19231 (N_19231,N_12596,N_11395);
nor U19232 (N_19232,N_13741,N_10240);
nor U19233 (N_19233,N_13866,N_12393);
nor U19234 (N_19234,N_14521,N_14280);
or U19235 (N_19235,N_13846,N_11717);
or U19236 (N_19236,N_14687,N_10304);
nand U19237 (N_19237,N_13206,N_11434);
or U19238 (N_19238,N_14513,N_12779);
xnor U19239 (N_19239,N_14136,N_14818);
nor U19240 (N_19240,N_11015,N_11770);
or U19241 (N_19241,N_13814,N_14875);
or U19242 (N_19242,N_12761,N_10623);
and U19243 (N_19243,N_13021,N_13192);
or U19244 (N_19244,N_10624,N_11186);
and U19245 (N_19245,N_10046,N_11994);
nor U19246 (N_19246,N_10875,N_13004);
xnor U19247 (N_19247,N_11973,N_10596);
and U19248 (N_19248,N_14416,N_14384);
and U19249 (N_19249,N_12235,N_11816);
xnor U19250 (N_19250,N_13906,N_10903);
nand U19251 (N_19251,N_11516,N_13645);
xor U19252 (N_19252,N_14781,N_11742);
xnor U19253 (N_19253,N_11695,N_10256);
or U19254 (N_19254,N_13476,N_14948);
nor U19255 (N_19255,N_12246,N_13954);
and U19256 (N_19256,N_13994,N_10734);
nor U19257 (N_19257,N_10275,N_10574);
xnor U19258 (N_19258,N_13023,N_10387);
or U19259 (N_19259,N_10811,N_14438);
nor U19260 (N_19260,N_14860,N_11008);
or U19261 (N_19261,N_14492,N_13657);
or U19262 (N_19262,N_14670,N_13244);
and U19263 (N_19263,N_11569,N_11528);
nand U19264 (N_19264,N_11056,N_13217);
and U19265 (N_19265,N_12417,N_14415);
and U19266 (N_19266,N_10337,N_12100);
and U19267 (N_19267,N_11841,N_12379);
nor U19268 (N_19268,N_12817,N_11990);
or U19269 (N_19269,N_10481,N_12217);
or U19270 (N_19270,N_10635,N_11738);
nor U19271 (N_19271,N_13841,N_13314);
xnor U19272 (N_19272,N_12633,N_13566);
or U19273 (N_19273,N_11311,N_12557);
nand U19274 (N_19274,N_11324,N_10243);
xnor U19275 (N_19275,N_10148,N_13200);
or U19276 (N_19276,N_12121,N_10374);
and U19277 (N_19277,N_13910,N_11982);
and U19278 (N_19278,N_13284,N_11087);
nor U19279 (N_19279,N_14054,N_10798);
nor U19280 (N_19280,N_10025,N_11110);
and U19281 (N_19281,N_10129,N_13495);
xnor U19282 (N_19282,N_11189,N_10042);
xor U19283 (N_19283,N_14658,N_11580);
or U19284 (N_19284,N_14376,N_10924);
nand U19285 (N_19285,N_14096,N_10348);
nor U19286 (N_19286,N_14750,N_11947);
nor U19287 (N_19287,N_10453,N_11478);
or U19288 (N_19288,N_10230,N_10319);
and U19289 (N_19289,N_12573,N_11283);
nor U19290 (N_19290,N_11799,N_13294);
or U19291 (N_19291,N_13219,N_12226);
and U19292 (N_19292,N_11512,N_14525);
nand U19293 (N_19293,N_14135,N_13181);
and U19294 (N_19294,N_11038,N_13606);
nand U19295 (N_19295,N_10412,N_11612);
or U19296 (N_19296,N_11024,N_13953);
nor U19297 (N_19297,N_14447,N_14935);
or U19298 (N_19298,N_11113,N_12683);
xnor U19299 (N_19299,N_14335,N_14633);
or U19300 (N_19300,N_12617,N_12036);
xor U19301 (N_19301,N_12550,N_13570);
and U19302 (N_19302,N_14750,N_14164);
nand U19303 (N_19303,N_10768,N_14890);
nor U19304 (N_19304,N_14478,N_13810);
and U19305 (N_19305,N_12952,N_12942);
xor U19306 (N_19306,N_11441,N_10189);
or U19307 (N_19307,N_13461,N_11289);
or U19308 (N_19308,N_14255,N_11930);
nand U19309 (N_19309,N_10622,N_10103);
nor U19310 (N_19310,N_13013,N_13541);
and U19311 (N_19311,N_14140,N_11336);
nor U19312 (N_19312,N_13002,N_14068);
xnor U19313 (N_19313,N_12465,N_11384);
nand U19314 (N_19314,N_10328,N_11191);
or U19315 (N_19315,N_13141,N_10717);
xor U19316 (N_19316,N_12432,N_13676);
and U19317 (N_19317,N_12438,N_13212);
and U19318 (N_19318,N_13817,N_10652);
xor U19319 (N_19319,N_12457,N_11938);
or U19320 (N_19320,N_12575,N_10812);
nand U19321 (N_19321,N_10520,N_13782);
nand U19322 (N_19322,N_12400,N_11260);
nand U19323 (N_19323,N_12871,N_11635);
and U19324 (N_19324,N_14200,N_12651);
xnor U19325 (N_19325,N_11506,N_10500);
nand U19326 (N_19326,N_10429,N_11412);
xor U19327 (N_19327,N_13891,N_14555);
xnor U19328 (N_19328,N_14117,N_14349);
and U19329 (N_19329,N_13204,N_13596);
and U19330 (N_19330,N_10276,N_12724);
and U19331 (N_19331,N_10708,N_14206);
and U19332 (N_19332,N_13338,N_10289);
xor U19333 (N_19333,N_10361,N_14215);
nor U19334 (N_19334,N_12995,N_12038);
xnor U19335 (N_19335,N_13853,N_14881);
or U19336 (N_19336,N_12953,N_12884);
and U19337 (N_19337,N_10793,N_13729);
nand U19338 (N_19338,N_13809,N_10649);
nand U19339 (N_19339,N_13616,N_13730);
and U19340 (N_19340,N_10908,N_11735);
nand U19341 (N_19341,N_12322,N_12551);
nand U19342 (N_19342,N_13797,N_13566);
or U19343 (N_19343,N_10110,N_11655);
and U19344 (N_19344,N_12212,N_10989);
and U19345 (N_19345,N_13265,N_12821);
and U19346 (N_19346,N_13685,N_14127);
and U19347 (N_19347,N_12057,N_11002);
and U19348 (N_19348,N_12397,N_10516);
xnor U19349 (N_19349,N_12955,N_14586);
and U19350 (N_19350,N_10607,N_10308);
xnor U19351 (N_19351,N_12417,N_10334);
xor U19352 (N_19352,N_10224,N_11832);
or U19353 (N_19353,N_13684,N_13130);
or U19354 (N_19354,N_13659,N_12820);
nand U19355 (N_19355,N_13413,N_10521);
nand U19356 (N_19356,N_12341,N_11407);
or U19357 (N_19357,N_12489,N_14977);
nand U19358 (N_19358,N_10776,N_14995);
and U19359 (N_19359,N_13642,N_11581);
or U19360 (N_19360,N_10964,N_13774);
and U19361 (N_19361,N_13620,N_11409);
nor U19362 (N_19362,N_12917,N_11970);
nor U19363 (N_19363,N_14255,N_10308);
nor U19364 (N_19364,N_14360,N_13367);
nand U19365 (N_19365,N_14437,N_11112);
xnor U19366 (N_19366,N_11004,N_10861);
or U19367 (N_19367,N_11091,N_13851);
nor U19368 (N_19368,N_11925,N_11560);
nand U19369 (N_19369,N_11085,N_12689);
xnor U19370 (N_19370,N_12422,N_10399);
xnor U19371 (N_19371,N_11212,N_11278);
nor U19372 (N_19372,N_10226,N_13898);
xor U19373 (N_19373,N_14680,N_14959);
nand U19374 (N_19374,N_10581,N_14829);
nand U19375 (N_19375,N_14688,N_13626);
nand U19376 (N_19376,N_10101,N_10451);
and U19377 (N_19377,N_14488,N_14948);
and U19378 (N_19378,N_14640,N_11330);
and U19379 (N_19379,N_14321,N_11928);
nor U19380 (N_19380,N_13330,N_10648);
or U19381 (N_19381,N_11561,N_10916);
and U19382 (N_19382,N_10120,N_13008);
and U19383 (N_19383,N_11939,N_14201);
xnor U19384 (N_19384,N_12710,N_12201);
or U19385 (N_19385,N_10511,N_11145);
or U19386 (N_19386,N_10373,N_10843);
nand U19387 (N_19387,N_10373,N_12226);
xor U19388 (N_19388,N_11390,N_12116);
nor U19389 (N_19389,N_11293,N_13268);
nor U19390 (N_19390,N_13694,N_14835);
nor U19391 (N_19391,N_12709,N_13586);
nor U19392 (N_19392,N_11631,N_13128);
or U19393 (N_19393,N_14072,N_11396);
nor U19394 (N_19394,N_11659,N_11649);
or U19395 (N_19395,N_14027,N_10519);
or U19396 (N_19396,N_10381,N_14716);
or U19397 (N_19397,N_12708,N_13129);
xor U19398 (N_19398,N_12896,N_10931);
xnor U19399 (N_19399,N_12264,N_14700);
nand U19400 (N_19400,N_11986,N_10972);
or U19401 (N_19401,N_12796,N_13823);
or U19402 (N_19402,N_13097,N_13474);
xor U19403 (N_19403,N_12656,N_12204);
and U19404 (N_19404,N_12191,N_14845);
nor U19405 (N_19405,N_11479,N_14106);
xnor U19406 (N_19406,N_14508,N_14671);
nor U19407 (N_19407,N_12177,N_11489);
and U19408 (N_19408,N_14797,N_12935);
and U19409 (N_19409,N_11801,N_12289);
xnor U19410 (N_19410,N_14695,N_14060);
xnor U19411 (N_19411,N_12337,N_12289);
nand U19412 (N_19412,N_10896,N_13095);
xnor U19413 (N_19413,N_13248,N_12017);
or U19414 (N_19414,N_12432,N_11435);
nor U19415 (N_19415,N_13717,N_13925);
nor U19416 (N_19416,N_13422,N_12100);
nor U19417 (N_19417,N_10263,N_14982);
nor U19418 (N_19418,N_13193,N_11306);
xor U19419 (N_19419,N_14387,N_14746);
nor U19420 (N_19420,N_12291,N_10992);
xor U19421 (N_19421,N_12739,N_14536);
nor U19422 (N_19422,N_10878,N_14517);
xnor U19423 (N_19423,N_11202,N_14708);
nand U19424 (N_19424,N_14013,N_12241);
nand U19425 (N_19425,N_12141,N_14256);
nor U19426 (N_19426,N_11219,N_13057);
and U19427 (N_19427,N_13674,N_14337);
nor U19428 (N_19428,N_13806,N_13630);
and U19429 (N_19429,N_14002,N_12986);
nor U19430 (N_19430,N_11646,N_11001);
nand U19431 (N_19431,N_10155,N_14026);
and U19432 (N_19432,N_13224,N_12302);
nand U19433 (N_19433,N_10623,N_12542);
and U19434 (N_19434,N_12791,N_11418);
nor U19435 (N_19435,N_11808,N_12647);
and U19436 (N_19436,N_10283,N_11646);
nor U19437 (N_19437,N_14165,N_12844);
nor U19438 (N_19438,N_13884,N_13433);
and U19439 (N_19439,N_13203,N_13640);
xnor U19440 (N_19440,N_10027,N_11404);
and U19441 (N_19441,N_14257,N_12598);
or U19442 (N_19442,N_13725,N_13294);
xnor U19443 (N_19443,N_13610,N_13585);
nor U19444 (N_19444,N_10933,N_14078);
nor U19445 (N_19445,N_10077,N_10100);
or U19446 (N_19446,N_10531,N_10275);
nand U19447 (N_19447,N_10465,N_13534);
xnor U19448 (N_19448,N_10718,N_10830);
and U19449 (N_19449,N_11465,N_11997);
or U19450 (N_19450,N_11392,N_14818);
and U19451 (N_19451,N_11678,N_12182);
or U19452 (N_19452,N_13376,N_10884);
xnor U19453 (N_19453,N_12842,N_10331);
and U19454 (N_19454,N_13924,N_12050);
and U19455 (N_19455,N_14586,N_10648);
xor U19456 (N_19456,N_11141,N_12795);
or U19457 (N_19457,N_12008,N_13698);
and U19458 (N_19458,N_13144,N_11056);
and U19459 (N_19459,N_12639,N_12448);
xor U19460 (N_19460,N_13141,N_11532);
nand U19461 (N_19461,N_13139,N_11379);
nand U19462 (N_19462,N_12007,N_13973);
nand U19463 (N_19463,N_10671,N_12570);
xor U19464 (N_19464,N_11926,N_12032);
or U19465 (N_19465,N_11076,N_13126);
or U19466 (N_19466,N_11336,N_10091);
and U19467 (N_19467,N_12234,N_10330);
nor U19468 (N_19468,N_14315,N_13875);
nand U19469 (N_19469,N_14784,N_13668);
nand U19470 (N_19470,N_12155,N_10574);
nor U19471 (N_19471,N_13150,N_14673);
and U19472 (N_19472,N_11120,N_10994);
xnor U19473 (N_19473,N_13364,N_13760);
nand U19474 (N_19474,N_12721,N_13215);
and U19475 (N_19475,N_13163,N_11442);
nand U19476 (N_19476,N_11705,N_12209);
xnor U19477 (N_19477,N_12494,N_10050);
and U19478 (N_19478,N_12674,N_12582);
xnor U19479 (N_19479,N_10677,N_10968);
nor U19480 (N_19480,N_13206,N_11078);
and U19481 (N_19481,N_14989,N_11121);
or U19482 (N_19482,N_12116,N_14082);
nor U19483 (N_19483,N_13061,N_13907);
nand U19484 (N_19484,N_12126,N_11833);
nand U19485 (N_19485,N_12167,N_14701);
and U19486 (N_19486,N_11583,N_14985);
nand U19487 (N_19487,N_11256,N_10088);
and U19488 (N_19488,N_11772,N_12757);
xnor U19489 (N_19489,N_13132,N_13055);
nand U19490 (N_19490,N_12732,N_12862);
xnor U19491 (N_19491,N_13390,N_11881);
xnor U19492 (N_19492,N_12755,N_12490);
and U19493 (N_19493,N_10990,N_13701);
and U19494 (N_19494,N_11575,N_12919);
or U19495 (N_19495,N_10969,N_14461);
nor U19496 (N_19496,N_11026,N_12343);
nand U19497 (N_19497,N_12041,N_14825);
xnor U19498 (N_19498,N_11130,N_14807);
nor U19499 (N_19499,N_11631,N_13470);
nand U19500 (N_19500,N_11243,N_11734);
nor U19501 (N_19501,N_11527,N_14868);
nor U19502 (N_19502,N_14706,N_13322);
and U19503 (N_19503,N_14792,N_10521);
nor U19504 (N_19504,N_12968,N_10970);
nand U19505 (N_19505,N_11653,N_14722);
nand U19506 (N_19506,N_13127,N_13189);
xor U19507 (N_19507,N_14732,N_12498);
or U19508 (N_19508,N_11095,N_13750);
nand U19509 (N_19509,N_14149,N_11598);
nand U19510 (N_19510,N_12833,N_11521);
nor U19511 (N_19511,N_14049,N_11305);
xor U19512 (N_19512,N_11342,N_14986);
and U19513 (N_19513,N_14252,N_14031);
nor U19514 (N_19514,N_12136,N_13365);
xor U19515 (N_19515,N_10911,N_12028);
and U19516 (N_19516,N_14504,N_11644);
nand U19517 (N_19517,N_10713,N_13928);
and U19518 (N_19518,N_11758,N_10993);
nor U19519 (N_19519,N_10571,N_13090);
or U19520 (N_19520,N_10148,N_10535);
or U19521 (N_19521,N_13417,N_14853);
nand U19522 (N_19522,N_12207,N_12319);
or U19523 (N_19523,N_13178,N_14211);
xor U19524 (N_19524,N_12846,N_13861);
xor U19525 (N_19525,N_10781,N_13012);
xor U19526 (N_19526,N_13079,N_12484);
nor U19527 (N_19527,N_13206,N_11906);
xor U19528 (N_19528,N_11212,N_13225);
xnor U19529 (N_19529,N_10085,N_10262);
and U19530 (N_19530,N_10826,N_14595);
nor U19531 (N_19531,N_13382,N_12213);
and U19532 (N_19532,N_10880,N_12043);
xnor U19533 (N_19533,N_12197,N_10262);
and U19534 (N_19534,N_11374,N_13773);
nor U19535 (N_19535,N_12674,N_13047);
or U19536 (N_19536,N_10271,N_14529);
xor U19537 (N_19537,N_10698,N_11680);
nor U19538 (N_19538,N_13807,N_10649);
nand U19539 (N_19539,N_12551,N_11664);
nand U19540 (N_19540,N_10874,N_13344);
and U19541 (N_19541,N_14713,N_11052);
nand U19542 (N_19542,N_10349,N_12869);
or U19543 (N_19543,N_14238,N_13090);
and U19544 (N_19544,N_13949,N_13972);
nor U19545 (N_19545,N_11242,N_13678);
and U19546 (N_19546,N_11054,N_14917);
nand U19547 (N_19547,N_11448,N_13255);
nand U19548 (N_19548,N_10306,N_11407);
nand U19549 (N_19549,N_10856,N_12329);
or U19550 (N_19550,N_14247,N_13067);
nor U19551 (N_19551,N_11743,N_13901);
or U19552 (N_19552,N_14376,N_13336);
nand U19553 (N_19553,N_14257,N_10598);
nand U19554 (N_19554,N_13806,N_14489);
nand U19555 (N_19555,N_10496,N_13350);
xnor U19556 (N_19556,N_14754,N_13041);
nand U19557 (N_19557,N_11522,N_11144);
nand U19558 (N_19558,N_14621,N_12874);
nor U19559 (N_19559,N_14485,N_14528);
nor U19560 (N_19560,N_14164,N_12005);
nand U19561 (N_19561,N_14859,N_14801);
and U19562 (N_19562,N_14415,N_13171);
or U19563 (N_19563,N_14497,N_11406);
nor U19564 (N_19564,N_13639,N_11180);
or U19565 (N_19565,N_11396,N_14403);
nand U19566 (N_19566,N_14068,N_13109);
and U19567 (N_19567,N_12509,N_14003);
nor U19568 (N_19568,N_11839,N_11089);
nand U19569 (N_19569,N_12361,N_13700);
nor U19570 (N_19570,N_14479,N_12360);
or U19571 (N_19571,N_14435,N_14298);
or U19572 (N_19572,N_11648,N_11841);
xor U19573 (N_19573,N_11431,N_12964);
xor U19574 (N_19574,N_11226,N_12333);
xor U19575 (N_19575,N_10208,N_12071);
and U19576 (N_19576,N_10118,N_11526);
or U19577 (N_19577,N_14019,N_12289);
and U19578 (N_19578,N_10384,N_12411);
nor U19579 (N_19579,N_12648,N_11306);
nand U19580 (N_19580,N_13247,N_10783);
and U19581 (N_19581,N_13669,N_10357);
nor U19582 (N_19582,N_14037,N_14902);
nor U19583 (N_19583,N_11883,N_11309);
and U19584 (N_19584,N_14516,N_13478);
nand U19585 (N_19585,N_11344,N_14152);
and U19586 (N_19586,N_13121,N_14093);
and U19587 (N_19587,N_13721,N_10050);
nand U19588 (N_19588,N_13340,N_13091);
and U19589 (N_19589,N_13160,N_14555);
nand U19590 (N_19590,N_13378,N_11694);
nand U19591 (N_19591,N_14887,N_10624);
xnor U19592 (N_19592,N_10163,N_12271);
and U19593 (N_19593,N_10002,N_14651);
nand U19594 (N_19594,N_12928,N_12924);
xor U19595 (N_19595,N_13974,N_12651);
and U19596 (N_19596,N_10566,N_13171);
or U19597 (N_19597,N_14184,N_13002);
nand U19598 (N_19598,N_13217,N_10423);
and U19599 (N_19599,N_10615,N_10024);
nor U19600 (N_19600,N_10911,N_14748);
nor U19601 (N_19601,N_10180,N_14735);
or U19602 (N_19602,N_11312,N_14736);
nand U19603 (N_19603,N_13722,N_10562);
nor U19604 (N_19604,N_13292,N_11410);
and U19605 (N_19605,N_14136,N_13467);
xor U19606 (N_19606,N_12409,N_10370);
nor U19607 (N_19607,N_10054,N_14905);
and U19608 (N_19608,N_12075,N_11996);
xor U19609 (N_19609,N_12792,N_11297);
nor U19610 (N_19610,N_11087,N_12493);
nor U19611 (N_19611,N_12430,N_13779);
or U19612 (N_19612,N_10187,N_10516);
or U19613 (N_19613,N_12015,N_10433);
nor U19614 (N_19614,N_12662,N_14011);
xnor U19615 (N_19615,N_13277,N_12200);
or U19616 (N_19616,N_11142,N_13950);
or U19617 (N_19617,N_10459,N_12819);
and U19618 (N_19618,N_14444,N_10702);
and U19619 (N_19619,N_12037,N_14958);
or U19620 (N_19620,N_14226,N_14805);
nand U19621 (N_19621,N_10781,N_14662);
nand U19622 (N_19622,N_10960,N_13618);
nor U19623 (N_19623,N_13994,N_13861);
or U19624 (N_19624,N_11727,N_11066);
and U19625 (N_19625,N_11811,N_13522);
or U19626 (N_19626,N_13181,N_14926);
xnor U19627 (N_19627,N_13475,N_11432);
nor U19628 (N_19628,N_11166,N_10870);
nor U19629 (N_19629,N_13560,N_10411);
nor U19630 (N_19630,N_14051,N_10571);
and U19631 (N_19631,N_10083,N_14838);
nand U19632 (N_19632,N_10255,N_14840);
xnor U19633 (N_19633,N_11119,N_13196);
nor U19634 (N_19634,N_12585,N_11818);
and U19635 (N_19635,N_12923,N_10417);
xnor U19636 (N_19636,N_12243,N_12025);
and U19637 (N_19637,N_11228,N_10260);
xor U19638 (N_19638,N_11472,N_14021);
and U19639 (N_19639,N_12990,N_11458);
nand U19640 (N_19640,N_13877,N_10823);
nor U19641 (N_19641,N_13203,N_10480);
or U19642 (N_19642,N_12561,N_12759);
nand U19643 (N_19643,N_14364,N_10503);
nor U19644 (N_19644,N_11910,N_13037);
nor U19645 (N_19645,N_12683,N_14862);
and U19646 (N_19646,N_14291,N_14686);
nand U19647 (N_19647,N_14823,N_13763);
nor U19648 (N_19648,N_10458,N_11761);
nor U19649 (N_19649,N_10507,N_10467);
xnor U19650 (N_19650,N_12374,N_11639);
nand U19651 (N_19651,N_12638,N_14207);
and U19652 (N_19652,N_14543,N_11823);
xor U19653 (N_19653,N_12023,N_13689);
or U19654 (N_19654,N_10665,N_13452);
xor U19655 (N_19655,N_11348,N_13985);
or U19656 (N_19656,N_13461,N_12579);
xor U19657 (N_19657,N_14770,N_13539);
nor U19658 (N_19658,N_14326,N_10896);
and U19659 (N_19659,N_10449,N_12762);
or U19660 (N_19660,N_11064,N_13472);
nand U19661 (N_19661,N_13246,N_10539);
or U19662 (N_19662,N_10535,N_12192);
xor U19663 (N_19663,N_10423,N_14781);
nand U19664 (N_19664,N_12453,N_14836);
and U19665 (N_19665,N_11919,N_14145);
and U19666 (N_19666,N_13058,N_12249);
nand U19667 (N_19667,N_12410,N_14299);
and U19668 (N_19668,N_12574,N_10580);
nand U19669 (N_19669,N_13545,N_11904);
and U19670 (N_19670,N_13435,N_10169);
nor U19671 (N_19671,N_14505,N_13781);
nand U19672 (N_19672,N_11294,N_12594);
nor U19673 (N_19673,N_10404,N_11271);
xor U19674 (N_19674,N_10931,N_12526);
nand U19675 (N_19675,N_10517,N_13576);
nand U19676 (N_19676,N_11520,N_12495);
or U19677 (N_19677,N_12197,N_13923);
xor U19678 (N_19678,N_14442,N_12654);
or U19679 (N_19679,N_10731,N_11984);
nand U19680 (N_19680,N_11701,N_12761);
xor U19681 (N_19681,N_12520,N_11317);
and U19682 (N_19682,N_13749,N_12130);
and U19683 (N_19683,N_11434,N_10881);
xor U19684 (N_19684,N_12454,N_13852);
and U19685 (N_19685,N_13571,N_12326);
nor U19686 (N_19686,N_12208,N_13758);
nor U19687 (N_19687,N_13335,N_12756);
nand U19688 (N_19688,N_11378,N_11247);
nand U19689 (N_19689,N_14593,N_11964);
nor U19690 (N_19690,N_14288,N_13540);
and U19691 (N_19691,N_12135,N_12586);
xnor U19692 (N_19692,N_13748,N_13674);
nor U19693 (N_19693,N_14229,N_11505);
nor U19694 (N_19694,N_14109,N_10093);
nand U19695 (N_19695,N_11917,N_11239);
nand U19696 (N_19696,N_12307,N_10279);
nand U19697 (N_19697,N_11605,N_11222);
xor U19698 (N_19698,N_13240,N_13800);
nor U19699 (N_19699,N_11158,N_10447);
nand U19700 (N_19700,N_14318,N_14354);
xor U19701 (N_19701,N_10924,N_14805);
nand U19702 (N_19702,N_13089,N_14971);
nor U19703 (N_19703,N_12058,N_13668);
nand U19704 (N_19704,N_13338,N_14943);
xor U19705 (N_19705,N_10496,N_10967);
xnor U19706 (N_19706,N_10262,N_13963);
xor U19707 (N_19707,N_12220,N_11689);
and U19708 (N_19708,N_13692,N_10859);
nand U19709 (N_19709,N_12544,N_11327);
and U19710 (N_19710,N_12274,N_11308);
or U19711 (N_19711,N_14983,N_14160);
nor U19712 (N_19712,N_12301,N_10487);
or U19713 (N_19713,N_13168,N_14551);
nand U19714 (N_19714,N_10509,N_11193);
xor U19715 (N_19715,N_14010,N_12930);
or U19716 (N_19716,N_13269,N_13244);
nand U19717 (N_19717,N_12710,N_11559);
or U19718 (N_19718,N_10232,N_13641);
xor U19719 (N_19719,N_10566,N_12045);
nor U19720 (N_19720,N_13364,N_10624);
nand U19721 (N_19721,N_14516,N_12539);
nor U19722 (N_19722,N_14293,N_13435);
or U19723 (N_19723,N_12701,N_12049);
and U19724 (N_19724,N_14528,N_14987);
or U19725 (N_19725,N_10798,N_14294);
nor U19726 (N_19726,N_12580,N_11015);
nor U19727 (N_19727,N_11611,N_13274);
nand U19728 (N_19728,N_12006,N_12728);
or U19729 (N_19729,N_13403,N_12468);
nand U19730 (N_19730,N_10707,N_13876);
or U19731 (N_19731,N_12487,N_12859);
or U19732 (N_19732,N_14637,N_14283);
or U19733 (N_19733,N_11145,N_11139);
and U19734 (N_19734,N_14958,N_12767);
nor U19735 (N_19735,N_10545,N_13161);
and U19736 (N_19736,N_11910,N_10760);
xnor U19737 (N_19737,N_10340,N_11161);
xor U19738 (N_19738,N_13083,N_10147);
xnor U19739 (N_19739,N_13957,N_12329);
or U19740 (N_19740,N_10725,N_10135);
or U19741 (N_19741,N_14948,N_12426);
and U19742 (N_19742,N_11886,N_11222);
xnor U19743 (N_19743,N_13673,N_11506);
or U19744 (N_19744,N_12492,N_14364);
xor U19745 (N_19745,N_14190,N_13937);
xor U19746 (N_19746,N_12071,N_10149);
nand U19747 (N_19747,N_10664,N_11202);
xor U19748 (N_19748,N_13582,N_12655);
nand U19749 (N_19749,N_10699,N_11081);
or U19750 (N_19750,N_13365,N_13455);
xnor U19751 (N_19751,N_14983,N_12078);
xor U19752 (N_19752,N_13740,N_12875);
nand U19753 (N_19753,N_11701,N_14757);
nor U19754 (N_19754,N_12477,N_12968);
nand U19755 (N_19755,N_11905,N_13510);
nand U19756 (N_19756,N_12719,N_10866);
or U19757 (N_19757,N_10121,N_13458);
nand U19758 (N_19758,N_11167,N_12702);
xnor U19759 (N_19759,N_12700,N_14577);
nor U19760 (N_19760,N_14539,N_12626);
and U19761 (N_19761,N_11025,N_10935);
nand U19762 (N_19762,N_14805,N_13575);
or U19763 (N_19763,N_13221,N_12711);
and U19764 (N_19764,N_13368,N_10207);
and U19765 (N_19765,N_11144,N_10085);
xor U19766 (N_19766,N_11910,N_12441);
xnor U19767 (N_19767,N_10640,N_14982);
and U19768 (N_19768,N_14402,N_14782);
or U19769 (N_19769,N_13779,N_13449);
nor U19770 (N_19770,N_10544,N_11097);
nand U19771 (N_19771,N_10061,N_13610);
and U19772 (N_19772,N_14772,N_11303);
nand U19773 (N_19773,N_12989,N_10893);
nor U19774 (N_19774,N_13988,N_10917);
xor U19775 (N_19775,N_14677,N_11255);
nand U19776 (N_19776,N_10882,N_13655);
nand U19777 (N_19777,N_12386,N_12122);
nand U19778 (N_19778,N_14387,N_11157);
nor U19779 (N_19779,N_13552,N_11382);
nand U19780 (N_19780,N_14250,N_12381);
and U19781 (N_19781,N_13240,N_13171);
and U19782 (N_19782,N_11328,N_14945);
and U19783 (N_19783,N_13859,N_14780);
xnor U19784 (N_19784,N_14089,N_13519);
nand U19785 (N_19785,N_12072,N_13521);
and U19786 (N_19786,N_10749,N_14901);
xor U19787 (N_19787,N_14435,N_10646);
and U19788 (N_19788,N_13127,N_10658);
nand U19789 (N_19789,N_10127,N_13235);
and U19790 (N_19790,N_10423,N_12836);
xor U19791 (N_19791,N_10097,N_11951);
xnor U19792 (N_19792,N_14213,N_11255);
and U19793 (N_19793,N_10578,N_10720);
or U19794 (N_19794,N_13707,N_12702);
and U19795 (N_19795,N_11674,N_12684);
nand U19796 (N_19796,N_11279,N_10554);
nor U19797 (N_19797,N_11537,N_13877);
and U19798 (N_19798,N_12509,N_10831);
nor U19799 (N_19799,N_11301,N_13122);
or U19800 (N_19800,N_12558,N_13678);
and U19801 (N_19801,N_13502,N_11819);
nor U19802 (N_19802,N_14719,N_12776);
nor U19803 (N_19803,N_12735,N_11916);
xor U19804 (N_19804,N_13018,N_11482);
and U19805 (N_19805,N_10736,N_14843);
or U19806 (N_19806,N_13720,N_12195);
nor U19807 (N_19807,N_10709,N_10503);
nand U19808 (N_19808,N_12408,N_14572);
nor U19809 (N_19809,N_10489,N_13751);
or U19810 (N_19810,N_11724,N_14720);
nand U19811 (N_19811,N_10564,N_12422);
nand U19812 (N_19812,N_10889,N_14296);
xor U19813 (N_19813,N_10281,N_14910);
or U19814 (N_19814,N_13742,N_12448);
nand U19815 (N_19815,N_14815,N_11592);
nand U19816 (N_19816,N_13321,N_13272);
nand U19817 (N_19817,N_12742,N_14751);
or U19818 (N_19818,N_10526,N_10314);
and U19819 (N_19819,N_13076,N_12571);
nor U19820 (N_19820,N_14490,N_11490);
or U19821 (N_19821,N_14553,N_14337);
nand U19822 (N_19822,N_12417,N_11370);
and U19823 (N_19823,N_11613,N_11082);
or U19824 (N_19824,N_12307,N_11000);
xnor U19825 (N_19825,N_14160,N_13002);
and U19826 (N_19826,N_10867,N_12581);
nor U19827 (N_19827,N_14916,N_11766);
xnor U19828 (N_19828,N_14487,N_11492);
or U19829 (N_19829,N_13576,N_11501);
xnor U19830 (N_19830,N_13166,N_13397);
xnor U19831 (N_19831,N_14351,N_11996);
nor U19832 (N_19832,N_10978,N_13857);
or U19833 (N_19833,N_12327,N_11474);
nand U19834 (N_19834,N_13936,N_11475);
and U19835 (N_19835,N_10661,N_10694);
and U19836 (N_19836,N_11770,N_10829);
and U19837 (N_19837,N_14424,N_11784);
and U19838 (N_19838,N_10763,N_13343);
and U19839 (N_19839,N_12229,N_11405);
nor U19840 (N_19840,N_14427,N_12012);
nor U19841 (N_19841,N_11875,N_10435);
nand U19842 (N_19842,N_11104,N_13475);
and U19843 (N_19843,N_11316,N_12883);
xor U19844 (N_19844,N_14932,N_13120);
and U19845 (N_19845,N_14362,N_14672);
or U19846 (N_19846,N_12165,N_11116);
xor U19847 (N_19847,N_13920,N_10298);
xnor U19848 (N_19848,N_13549,N_11069);
nand U19849 (N_19849,N_13836,N_11463);
nor U19850 (N_19850,N_10290,N_14365);
xor U19851 (N_19851,N_12886,N_11609);
and U19852 (N_19852,N_10699,N_10890);
or U19853 (N_19853,N_13478,N_10329);
nor U19854 (N_19854,N_14392,N_13000);
and U19855 (N_19855,N_11400,N_13371);
and U19856 (N_19856,N_14204,N_12237);
nand U19857 (N_19857,N_11875,N_14457);
xor U19858 (N_19858,N_13711,N_11412);
nand U19859 (N_19859,N_12535,N_14796);
nor U19860 (N_19860,N_14754,N_13236);
nand U19861 (N_19861,N_14659,N_14493);
nand U19862 (N_19862,N_10716,N_10277);
or U19863 (N_19863,N_10365,N_13512);
nor U19864 (N_19864,N_11310,N_14181);
or U19865 (N_19865,N_11184,N_10992);
and U19866 (N_19866,N_10799,N_14050);
nand U19867 (N_19867,N_12079,N_10572);
xnor U19868 (N_19868,N_10283,N_14290);
and U19869 (N_19869,N_10037,N_13218);
and U19870 (N_19870,N_10953,N_12502);
nor U19871 (N_19871,N_10548,N_14437);
and U19872 (N_19872,N_11982,N_10917);
nand U19873 (N_19873,N_13121,N_14975);
and U19874 (N_19874,N_14449,N_11352);
xor U19875 (N_19875,N_11070,N_11596);
or U19876 (N_19876,N_14159,N_14323);
xnor U19877 (N_19877,N_10581,N_11582);
nor U19878 (N_19878,N_11940,N_13826);
and U19879 (N_19879,N_10523,N_10066);
xnor U19880 (N_19880,N_11724,N_14413);
nor U19881 (N_19881,N_11961,N_14367);
nor U19882 (N_19882,N_12411,N_12592);
nand U19883 (N_19883,N_11304,N_13933);
nand U19884 (N_19884,N_10054,N_11864);
and U19885 (N_19885,N_13639,N_11382);
nor U19886 (N_19886,N_11975,N_14921);
or U19887 (N_19887,N_12873,N_14942);
nor U19888 (N_19888,N_13777,N_14967);
xor U19889 (N_19889,N_11802,N_14106);
xor U19890 (N_19890,N_13402,N_12693);
or U19891 (N_19891,N_11420,N_14045);
and U19892 (N_19892,N_12334,N_14233);
or U19893 (N_19893,N_14636,N_13234);
nand U19894 (N_19894,N_11665,N_13923);
nand U19895 (N_19895,N_12905,N_13697);
or U19896 (N_19896,N_13097,N_11502);
and U19897 (N_19897,N_12925,N_10502);
nor U19898 (N_19898,N_11400,N_14140);
nand U19899 (N_19899,N_12949,N_13384);
xor U19900 (N_19900,N_11404,N_13550);
and U19901 (N_19901,N_11803,N_13255);
xnor U19902 (N_19902,N_14681,N_13778);
or U19903 (N_19903,N_14874,N_10985);
and U19904 (N_19904,N_10125,N_10568);
or U19905 (N_19905,N_11600,N_10345);
and U19906 (N_19906,N_11723,N_11159);
xnor U19907 (N_19907,N_10093,N_14982);
and U19908 (N_19908,N_12968,N_10824);
or U19909 (N_19909,N_10831,N_13188);
or U19910 (N_19910,N_12282,N_13222);
or U19911 (N_19911,N_10378,N_12149);
or U19912 (N_19912,N_11079,N_13996);
nor U19913 (N_19913,N_13931,N_12152);
xor U19914 (N_19914,N_13439,N_13334);
nand U19915 (N_19915,N_12863,N_11155);
and U19916 (N_19916,N_12841,N_11570);
xor U19917 (N_19917,N_11922,N_11026);
xnor U19918 (N_19918,N_14680,N_11751);
nor U19919 (N_19919,N_10240,N_14913);
and U19920 (N_19920,N_13079,N_12225);
nand U19921 (N_19921,N_11058,N_11816);
or U19922 (N_19922,N_13032,N_10657);
nor U19923 (N_19923,N_10646,N_14206);
nand U19924 (N_19924,N_13178,N_13528);
nor U19925 (N_19925,N_12863,N_12887);
nor U19926 (N_19926,N_14477,N_11818);
or U19927 (N_19927,N_10507,N_11315);
nand U19928 (N_19928,N_13433,N_14714);
nor U19929 (N_19929,N_14273,N_10046);
or U19930 (N_19930,N_13603,N_13370);
nand U19931 (N_19931,N_11785,N_13074);
or U19932 (N_19932,N_11963,N_14066);
and U19933 (N_19933,N_14527,N_12833);
and U19934 (N_19934,N_11060,N_13184);
or U19935 (N_19935,N_13542,N_14408);
and U19936 (N_19936,N_10760,N_14703);
xor U19937 (N_19937,N_11946,N_13738);
nor U19938 (N_19938,N_10494,N_10106);
or U19939 (N_19939,N_14732,N_14983);
or U19940 (N_19940,N_10196,N_12337);
or U19941 (N_19941,N_10077,N_14872);
nand U19942 (N_19942,N_11877,N_12416);
and U19943 (N_19943,N_12780,N_13159);
or U19944 (N_19944,N_12660,N_11000);
or U19945 (N_19945,N_11601,N_12309);
nor U19946 (N_19946,N_13142,N_12428);
or U19947 (N_19947,N_12421,N_10802);
and U19948 (N_19948,N_11475,N_14508);
nand U19949 (N_19949,N_13527,N_10048);
nand U19950 (N_19950,N_12062,N_10836);
and U19951 (N_19951,N_12269,N_11676);
nand U19952 (N_19952,N_14516,N_10173);
or U19953 (N_19953,N_12674,N_12759);
and U19954 (N_19954,N_12642,N_12336);
nand U19955 (N_19955,N_13526,N_10616);
xnor U19956 (N_19956,N_13988,N_10112);
nor U19957 (N_19957,N_14295,N_12507);
and U19958 (N_19958,N_13695,N_10506);
nand U19959 (N_19959,N_13528,N_12167);
xor U19960 (N_19960,N_14983,N_11249);
nand U19961 (N_19961,N_13594,N_13801);
or U19962 (N_19962,N_11436,N_13674);
nor U19963 (N_19963,N_11218,N_10194);
and U19964 (N_19964,N_11787,N_12068);
nand U19965 (N_19965,N_12383,N_14790);
xor U19966 (N_19966,N_13723,N_10121);
and U19967 (N_19967,N_11348,N_13123);
or U19968 (N_19968,N_10359,N_14978);
xnor U19969 (N_19969,N_11270,N_11146);
and U19970 (N_19970,N_12130,N_10280);
nor U19971 (N_19971,N_12951,N_12184);
and U19972 (N_19972,N_13639,N_11023);
and U19973 (N_19973,N_14901,N_12894);
and U19974 (N_19974,N_14278,N_10600);
and U19975 (N_19975,N_10828,N_11375);
or U19976 (N_19976,N_12650,N_14635);
nand U19977 (N_19977,N_12798,N_12177);
nor U19978 (N_19978,N_13107,N_12271);
nor U19979 (N_19979,N_10467,N_12094);
nor U19980 (N_19980,N_11416,N_13938);
or U19981 (N_19981,N_10335,N_10444);
nand U19982 (N_19982,N_10727,N_14193);
nor U19983 (N_19983,N_13497,N_12320);
and U19984 (N_19984,N_12341,N_14337);
or U19985 (N_19985,N_10990,N_12132);
or U19986 (N_19986,N_11878,N_13639);
nor U19987 (N_19987,N_12010,N_10582);
nor U19988 (N_19988,N_14459,N_12457);
nand U19989 (N_19989,N_11390,N_11067);
or U19990 (N_19990,N_13785,N_11670);
or U19991 (N_19991,N_14125,N_14592);
xor U19992 (N_19992,N_13007,N_10620);
or U19993 (N_19993,N_11054,N_14742);
xor U19994 (N_19994,N_11338,N_11899);
or U19995 (N_19995,N_10395,N_13060);
xor U19996 (N_19996,N_10047,N_12242);
xor U19997 (N_19997,N_14547,N_11581);
nand U19998 (N_19998,N_12857,N_14912);
nor U19999 (N_19999,N_11001,N_11085);
nand U20000 (N_20000,N_18386,N_19679);
nand U20001 (N_20001,N_19950,N_18798);
and U20002 (N_20002,N_17330,N_18749);
and U20003 (N_20003,N_17509,N_18033);
xnor U20004 (N_20004,N_16890,N_19220);
and U20005 (N_20005,N_16988,N_19757);
and U20006 (N_20006,N_15622,N_19086);
nor U20007 (N_20007,N_17546,N_19833);
and U20008 (N_20008,N_17858,N_19458);
or U20009 (N_20009,N_18093,N_16628);
and U20010 (N_20010,N_17222,N_16026);
nor U20011 (N_20011,N_16031,N_17852);
or U20012 (N_20012,N_18611,N_15152);
or U20013 (N_20013,N_18905,N_17337);
or U20014 (N_20014,N_17477,N_19977);
and U20015 (N_20015,N_15600,N_17703);
nand U20016 (N_20016,N_18304,N_17817);
or U20017 (N_20017,N_19450,N_15137);
nand U20018 (N_20018,N_15125,N_17368);
nand U20019 (N_20019,N_16286,N_19648);
nor U20020 (N_20020,N_15110,N_15230);
and U20021 (N_20021,N_18312,N_16564);
nor U20022 (N_20022,N_16937,N_16416);
nor U20023 (N_20023,N_19097,N_18384);
and U20024 (N_20024,N_18311,N_18460);
xnor U20025 (N_20025,N_19460,N_17910);
nor U20026 (N_20026,N_15949,N_17680);
xor U20027 (N_20027,N_18595,N_15505);
nor U20028 (N_20028,N_15891,N_19793);
xnor U20029 (N_20029,N_15520,N_19560);
or U20030 (N_20030,N_19138,N_16724);
nor U20031 (N_20031,N_15328,N_18799);
nand U20032 (N_20032,N_16968,N_17804);
xor U20033 (N_20033,N_18725,N_19571);
and U20034 (N_20034,N_17593,N_17156);
and U20035 (N_20035,N_16050,N_17973);
and U20036 (N_20036,N_18796,N_18707);
or U20037 (N_20037,N_15357,N_19468);
nor U20038 (N_20038,N_15160,N_18371);
and U20039 (N_20039,N_17182,N_15626);
xor U20040 (N_20040,N_17310,N_19743);
xnor U20041 (N_20041,N_17980,N_15936);
and U20042 (N_20042,N_17746,N_18824);
and U20043 (N_20043,N_19152,N_19481);
or U20044 (N_20044,N_17913,N_19495);
nor U20045 (N_20045,N_15995,N_17771);
nand U20046 (N_20046,N_17432,N_16986);
and U20047 (N_20047,N_16484,N_16896);
nand U20048 (N_20048,N_17717,N_17170);
xnor U20049 (N_20049,N_15522,N_17054);
and U20050 (N_20050,N_18901,N_18462);
nand U20051 (N_20051,N_17424,N_19062);
or U20052 (N_20052,N_18468,N_18290);
or U20053 (N_20053,N_15890,N_19857);
or U20054 (N_20054,N_15424,N_19299);
or U20055 (N_20055,N_19698,N_19426);
or U20056 (N_20056,N_19213,N_17163);
nor U20057 (N_20057,N_17390,N_15761);
nor U20058 (N_20058,N_19387,N_17334);
nand U20059 (N_20059,N_16612,N_16759);
and U20060 (N_20060,N_15057,N_15299);
or U20061 (N_20061,N_19522,N_16208);
or U20062 (N_20062,N_16225,N_19342);
nor U20063 (N_20063,N_18537,N_19661);
nand U20064 (N_20064,N_16060,N_15694);
or U20065 (N_20065,N_19549,N_17952);
nand U20066 (N_20066,N_18729,N_15143);
or U20067 (N_20067,N_17677,N_17726);
xor U20068 (N_20068,N_19765,N_15275);
nor U20069 (N_20069,N_16247,N_18340);
nand U20070 (N_20070,N_15210,N_16842);
or U20071 (N_20071,N_18333,N_17438);
xor U20072 (N_20072,N_19919,N_18518);
or U20073 (N_20073,N_18098,N_17215);
or U20074 (N_20074,N_19365,N_15216);
xor U20075 (N_20075,N_18286,N_17811);
nand U20076 (N_20076,N_19356,N_18024);
or U20077 (N_20077,N_17954,N_17520);
xor U20078 (N_20078,N_18783,N_15791);
nor U20079 (N_20079,N_17464,N_17266);
and U20080 (N_20080,N_15804,N_18578);
nand U20081 (N_20081,N_17417,N_19845);
nand U20082 (N_20082,N_16695,N_15506);
nand U20083 (N_20083,N_18847,N_19362);
nor U20084 (N_20084,N_17091,N_17890);
nor U20085 (N_20085,N_15387,N_17314);
nor U20086 (N_20086,N_18174,N_17906);
and U20087 (N_20087,N_16337,N_18104);
xor U20088 (N_20088,N_17660,N_17106);
nand U20089 (N_20089,N_18503,N_15266);
or U20090 (N_20090,N_16793,N_19404);
or U20091 (N_20091,N_16142,N_19108);
nor U20092 (N_20092,N_16686,N_19798);
or U20093 (N_20093,N_18586,N_16645);
or U20094 (N_20094,N_19194,N_15453);
and U20095 (N_20095,N_17760,N_19065);
and U20096 (N_20096,N_15236,N_18099);
nand U20097 (N_20097,N_16815,N_18234);
xor U20098 (N_20098,N_15827,N_16336);
and U20099 (N_20099,N_15406,N_16204);
nand U20100 (N_20100,N_16857,N_15774);
and U20101 (N_20101,N_17875,N_18983);
xnor U20102 (N_20102,N_17884,N_18288);
or U20103 (N_20103,N_18778,N_15464);
nand U20104 (N_20104,N_18878,N_18404);
nor U20105 (N_20105,N_16413,N_15831);
nor U20106 (N_20106,N_18950,N_16657);
xnor U20107 (N_20107,N_16807,N_16914);
and U20108 (N_20108,N_19005,N_16453);
nor U20109 (N_20109,N_18722,N_16016);
and U20110 (N_20110,N_16715,N_18270);
and U20111 (N_20111,N_17540,N_19508);
and U20112 (N_20112,N_15183,N_19707);
nor U20113 (N_20113,N_19732,N_18589);
nand U20114 (N_20114,N_16195,N_18125);
nand U20115 (N_20115,N_17622,N_18576);
or U20116 (N_20116,N_16231,N_19116);
and U20117 (N_20117,N_19423,N_16559);
or U20118 (N_20118,N_18599,N_18370);
xor U20119 (N_20119,N_15348,N_17691);
nand U20120 (N_20120,N_16916,N_19266);
nand U20121 (N_20121,N_16278,N_16811);
or U20122 (N_20122,N_16140,N_15544);
xnor U20123 (N_20123,N_17158,N_19318);
and U20124 (N_20124,N_17133,N_15055);
and U20125 (N_20125,N_17402,N_16505);
xor U20126 (N_20126,N_16522,N_18097);
xnor U20127 (N_20127,N_17654,N_17481);
nand U20128 (N_20128,N_18957,N_16718);
nor U20129 (N_20129,N_17358,N_15966);
nor U20130 (N_20130,N_19231,N_17932);
nand U20131 (N_20131,N_19255,N_15799);
and U20132 (N_20132,N_15190,N_19815);
or U20133 (N_20133,N_16828,N_15074);
and U20134 (N_20134,N_18207,N_15740);
nand U20135 (N_20135,N_19120,N_18508);
or U20136 (N_20136,N_19252,N_15240);
xor U20137 (N_20137,N_19650,N_19525);
nor U20138 (N_20138,N_18742,N_16076);
and U20139 (N_20139,N_18861,N_19173);
or U20140 (N_20140,N_17422,N_15434);
nor U20141 (N_20141,N_16917,N_16717);
nor U20142 (N_20142,N_18388,N_16586);
xor U20143 (N_20143,N_17071,N_16949);
xor U20144 (N_20144,N_15498,N_15805);
nor U20145 (N_20145,N_18512,N_18789);
nor U20146 (N_20146,N_19831,N_17284);
and U20147 (N_20147,N_16785,N_15448);
or U20148 (N_20148,N_18377,N_18476);
xor U20149 (N_20149,N_15519,N_16704);
or U20150 (N_20150,N_16602,N_16871);
nor U20151 (N_20151,N_18858,N_17118);
xor U20152 (N_20152,N_15965,N_19951);
and U20153 (N_20153,N_15385,N_18472);
nor U20154 (N_20154,N_16545,N_17398);
nand U20155 (N_20155,N_16116,N_18464);
nand U20156 (N_20156,N_17479,N_19302);
or U20157 (N_20157,N_17192,N_19544);
or U20158 (N_20158,N_18396,N_15900);
and U20159 (N_20159,N_18752,N_15704);
and U20160 (N_20160,N_19205,N_18342);
and U20161 (N_20161,N_16296,N_17434);
and U20162 (N_20162,N_19586,N_15342);
xor U20163 (N_20163,N_16503,N_15010);
and U20164 (N_20164,N_17792,N_15241);
and U20165 (N_20165,N_15497,N_17385);
and U20166 (N_20166,N_19644,N_18059);
nor U20167 (N_20167,N_17372,N_16036);
or U20168 (N_20168,N_17545,N_17309);
xor U20169 (N_20169,N_18680,N_19332);
and U20170 (N_20170,N_18579,N_16452);
nor U20171 (N_20171,N_15693,N_16113);
or U20172 (N_20172,N_15766,N_17474);
or U20173 (N_20173,N_19842,N_17818);
nor U20174 (N_20174,N_15003,N_19367);
nand U20175 (N_20175,N_18320,N_19656);
nor U20176 (N_20176,N_19444,N_18934);
or U20177 (N_20177,N_19841,N_17767);
nand U20178 (N_20178,N_16070,N_18065);
or U20179 (N_20179,N_18960,N_17871);
xor U20180 (N_20180,N_18916,N_17807);
or U20181 (N_20181,N_19888,N_16185);
nand U20182 (N_20182,N_16624,N_16763);
nor U20183 (N_20183,N_18064,N_15352);
xor U20184 (N_20184,N_15122,N_16712);
xor U20185 (N_20185,N_19967,N_18700);
or U20186 (N_20186,N_18378,N_17535);
nand U20187 (N_20187,N_19752,N_19256);
or U20188 (N_20188,N_17532,N_15186);
and U20189 (N_20189,N_18110,N_16633);
and U20190 (N_20190,N_16255,N_15372);
and U20191 (N_20191,N_19093,N_15621);
nand U20192 (N_20192,N_15811,N_15964);
nand U20193 (N_20193,N_17332,N_17510);
xor U20194 (N_20194,N_19337,N_18647);
nor U20195 (N_20195,N_16742,N_16895);
xnor U20196 (N_20196,N_15661,N_15129);
nand U20197 (N_20197,N_17058,N_16782);
or U20198 (N_20198,N_17271,N_19241);
and U20199 (N_20199,N_17525,N_18401);
xor U20200 (N_20200,N_18381,N_16953);
nor U20201 (N_20201,N_19984,N_17078);
nor U20202 (N_20202,N_16262,N_15664);
nor U20203 (N_20203,N_16283,N_15987);
or U20204 (N_20204,N_19368,N_19799);
nand U20205 (N_20205,N_18644,N_15150);
nand U20206 (N_20206,N_18732,N_19452);
and U20207 (N_20207,N_17038,N_16313);
nand U20208 (N_20208,N_15588,N_17748);
xnor U20209 (N_20209,N_17698,N_18146);
xnor U20210 (N_20210,N_17251,N_17589);
nand U20211 (N_20211,N_18527,N_19117);
and U20212 (N_20212,N_17830,N_17763);
nand U20213 (N_20213,N_16762,N_17754);
xor U20214 (N_20214,N_18547,N_18347);
nor U20215 (N_20215,N_15405,N_19176);
nor U20216 (N_20216,N_17781,N_15009);
nand U20217 (N_20217,N_18470,N_16108);
nor U20218 (N_20218,N_18635,N_19464);
nand U20219 (N_20219,N_17802,N_19230);
nand U20220 (N_20220,N_16285,N_19788);
nand U20221 (N_20221,N_16637,N_16274);
and U20222 (N_20222,N_16647,N_18214);
and U20223 (N_20223,N_16956,N_18914);
xnor U20224 (N_20224,N_16123,N_18669);
xnor U20225 (N_20225,N_19838,N_15962);
xor U20226 (N_20226,N_19653,N_17342);
xnor U20227 (N_20227,N_17489,N_16073);
nor U20228 (N_20228,N_16979,N_15617);
or U20229 (N_20229,N_17965,N_18693);
or U20230 (N_20230,N_15543,N_18985);
xor U20231 (N_20231,N_15298,N_17696);
nand U20232 (N_20232,N_16493,N_18826);
nand U20233 (N_20233,N_15111,N_16836);
or U20234 (N_20234,N_15658,N_15744);
xor U20235 (N_20235,N_16355,N_16211);
and U20236 (N_20236,N_16083,N_16611);
nand U20237 (N_20237,N_19132,N_19690);
or U20238 (N_20238,N_15360,N_18170);
nand U20239 (N_20239,N_18874,N_18230);
nor U20240 (N_20240,N_15688,N_17326);
or U20241 (N_20241,N_18860,N_18395);
xnor U20242 (N_20242,N_19575,N_18213);
xnor U20243 (N_20243,N_19882,N_17387);
or U20244 (N_20244,N_19493,N_17943);
or U20245 (N_20245,N_16046,N_17015);
and U20246 (N_20246,N_16374,N_19700);
and U20247 (N_20247,N_19274,N_16034);
nand U20248 (N_20248,N_16386,N_17850);
nor U20249 (N_20249,N_19585,N_18177);
or U20250 (N_20250,N_15164,N_15527);
and U20251 (N_20251,N_15700,N_15772);
or U20252 (N_20252,N_19272,N_19304);
nand U20253 (N_20253,N_15554,N_16054);
or U20254 (N_20254,N_16576,N_19658);
and U20255 (N_20255,N_15451,N_15162);
nor U20256 (N_20256,N_19741,N_19949);
xor U20257 (N_20257,N_19015,N_15848);
or U20258 (N_20258,N_19442,N_15838);
xor U20259 (N_20259,N_18643,N_16351);
nor U20260 (N_20260,N_15353,N_17718);
nor U20261 (N_20261,N_15339,N_17200);
nand U20262 (N_20262,N_16605,N_16965);
nor U20263 (N_20263,N_15018,N_15229);
nand U20264 (N_20264,N_16421,N_17277);
nand U20265 (N_20265,N_16859,N_17995);
xor U20266 (N_20266,N_19987,N_16414);
and U20267 (N_20267,N_16517,N_19758);
or U20268 (N_20268,N_16074,N_16735);
xor U20269 (N_20269,N_18203,N_17216);
or U20270 (N_20270,N_18415,N_19806);
nand U20271 (N_20271,N_18023,N_15728);
nor U20272 (N_20272,N_17824,N_17900);
or U20273 (N_20273,N_19903,N_18695);
nor U20274 (N_20274,N_19580,N_16887);
nand U20275 (N_20275,N_19394,N_16482);
or U20276 (N_20276,N_17421,N_18176);
and U20277 (N_20277,N_16430,N_15188);
nor U20278 (N_20278,N_18372,N_18987);
or U20279 (N_20279,N_16549,N_19001);
and U20280 (N_20280,N_19281,N_17968);
xnor U20281 (N_20281,N_15705,N_18140);
nor U20282 (N_20282,N_16212,N_16062);
xor U20283 (N_20283,N_16569,N_16974);
nand U20284 (N_20284,N_15986,N_16052);
xor U20285 (N_20285,N_18997,N_18086);
or U20286 (N_20286,N_18585,N_16415);
nor U20287 (N_20287,N_18767,N_17352);
and U20288 (N_20288,N_15878,N_17186);
and U20289 (N_20289,N_18921,N_15391);
and U20290 (N_20290,N_17427,N_16180);
or U20291 (N_20291,N_19548,N_15967);
or U20292 (N_20292,N_18947,N_15397);
nand U20293 (N_20293,N_18745,N_16188);
and U20294 (N_20294,N_18686,N_18753);
xor U20295 (N_20295,N_19488,N_15780);
nand U20296 (N_20296,N_19454,N_15564);
nand U20297 (N_20297,N_15749,N_19600);
or U20298 (N_20298,N_18444,N_16981);
xnor U20299 (N_20299,N_19898,N_19466);
or U20300 (N_20300,N_19968,N_16977);
xnor U20301 (N_20301,N_19602,N_17994);
xnor U20302 (N_20302,N_19537,N_19920);
xnor U20303 (N_20303,N_16141,N_18500);
or U20304 (N_20304,N_16338,N_15173);
nor U20305 (N_20305,N_17365,N_17829);
and U20306 (N_20306,N_19290,N_17530);
or U20307 (N_20307,N_16253,N_16470);
xnor U20308 (N_20308,N_15038,N_19325);
nand U20309 (N_20309,N_17490,N_19369);
xor U20310 (N_20310,N_16678,N_17776);
nand U20311 (N_20311,N_18893,N_19383);
nor U20312 (N_20312,N_18497,N_19523);
nor U20313 (N_20313,N_19958,N_15702);
nor U20314 (N_20314,N_19144,N_17144);
or U20315 (N_20315,N_17188,N_15221);
or U20316 (N_20316,N_16086,N_15773);
and U20317 (N_20317,N_18676,N_17895);
nand U20318 (N_20318,N_19469,N_17230);
nand U20319 (N_20319,N_18278,N_17204);
or U20320 (N_20320,N_19209,N_19029);
or U20321 (N_20321,N_15730,N_19701);
or U20322 (N_20322,N_19563,N_15839);
xnor U20323 (N_20323,N_16524,N_15824);
xnor U20324 (N_20324,N_19693,N_16580);
xor U20325 (N_20325,N_15507,N_17713);
or U20326 (N_20326,N_15712,N_18031);
xor U20327 (N_20327,N_18800,N_16494);
nor U20328 (N_20328,N_19007,N_19201);
xor U20329 (N_20329,N_19336,N_18072);
or U20330 (N_20330,N_16547,N_15604);
nor U20331 (N_20331,N_17795,N_17449);
nand U20332 (N_20332,N_17656,N_16197);
nand U20333 (N_20333,N_15721,N_17810);
nand U20334 (N_20334,N_18626,N_19472);
nor U20335 (N_20335,N_19860,N_17847);
or U20336 (N_20336,N_18619,N_16491);
and U20337 (N_20337,N_18991,N_18738);
nor U20338 (N_20338,N_17039,N_18974);
and U20339 (N_20339,N_17280,N_17259);
or U20340 (N_20340,N_15578,N_15073);
nor U20341 (N_20341,N_18632,N_18092);
nor U20342 (N_20342,N_15636,N_16769);
xnor U20343 (N_20343,N_19457,N_15227);
nor U20344 (N_20344,N_16952,N_18910);
nor U20345 (N_20345,N_17350,N_16901);
and U20346 (N_20346,N_16991,N_18667);
or U20347 (N_20347,N_15322,N_18977);
or U20348 (N_20348,N_18353,N_17245);
or U20349 (N_20349,N_17626,N_18556);
nor U20350 (N_20350,N_16248,N_18980);
nor U20351 (N_20351,N_18596,N_19912);
nor U20352 (N_20352,N_19427,N_18489);
xor U20353 (N_20353,N_15668,N_17722);
and U20354 (N_20354,N_16966,N_18906);
nand U20355 (N_20355,N_16287,N_16636);
and U20356 (N_20356,N_17909,N_15889);
or U20357 (N_20357,N_15934,N_15524);
nor U20358 (N_20358,N_19151,N_17956);
or U20359 (N_20359,N_18898,N_15370);
xor U20360 (N_20360,N_15097,N_19333);
or U20361 (N_20361,N_18613,N_19166);
nand U20362 (N_20362,N_19769,N_15202);
nor U20363 (N_20363,N_16693,N_17021);
nor U20364 (N_20364,N_17648,N_19710);
xor U20365 (N_20365,N_17134,N_15760);
and U20366 (N_20366,N_19373,N_15171);
nor U20367 (N_20367,N_18915,N_18041);
xnor U20368 (N_20368,N_16553,N_18535);
nand U20369 (N_20369,N_16063,N_15359);
nor U20370 (N_20370,N_15775,N_16623);
xor U20371 (N_20371,N_18037,N_17731);
nand U20372 (N_20372,N_19699,N_19753);
and U20373 (N_20373,N_18138,N_16428);
nor U20374 (N_20374,N_16927,N_18913);
nor U20375 (N_20375,N_18334,N_15618);
or U20376 (N_20376,N_16906,N_19036);
nand U20377 (N_20377,N_17185,N_16017);
xor U20378 (N_20378,N_18780,N_16816);
nor U20379 (N_20379,N_19978,N_16854);
or U20380 (N_20380,N_19329,N_19663);
xnor U20381 (N_20381,N_17564,N_19676);
nand U20382 (N_20382,N_18869,N_17307);
xor U20383 (N_20383,N_18498,N_19350);
nor U20384 (N_20384,N_16216,N_16822);
and U20385 (N_20385,N_18199,N_18117);
or U20386 (N_20386,N_17666,N_15248);
nand U20387 (N_20387,N_15343,N_19931);
or U20388 (N_20388,N_17503,N_17843);
and U20389 (N_20389,N_19865,N_17552);
and U20390 (N_20390,N_17566,N_15887);
nor U20391 (N_20391,N_19035,N_15457);
nor U20392 (N_20392,N_18782,N_18715);
or U20393 (N_20393,N_15968,N_15809);
nor U20394 (N_20394,N_17247,N_15070);
nand U20395 (N_20395,N_19824,N_15958);
or U20396 (N_20396,N_16349,N_16665);
nand U20397 (N_20397,N_16119,N_16281);
nor U20398 (N_20398,N_15425,N_19591);
nor U20399 (N_20399,N_18516,N_18337);
and U20400 (N_20400,N_16508,N_18422);
or U20401 (N_20401,N_17988,N_15847);
xnor U20402 (N_20402,N_15737,N_15609);
and U20403 (N_20403,N_17032,N_19639);
or U20404 (N_20404,N_19171,N_17712);
nand U20405 (N_20405,N_17793,N_17547);
nor U20406 (N_20406,N_17075,N_19961);
and U20407 (N_20407,N_18307,N_17812);
nor U20408 (N_20408,N_16673,N_19208);
nand U20409 (N_20409,N_19416,N_16124);
and U20410 (N_20410,N_17087,N_16406);
xnor U20411 (N_20411,N_16950,N_18348);
nand U20412 (N_20412,N_15896,N_17563);
xnor U20413 (N_20413,N_18791,N_19502);
nand U20414 (N_20414,N_16347,N_16539);
and U20415 (N_20415,N_15648,N_15284);
and U20416 (N_20416,N_19042,N_15330);
or U20417 (N_20417,N_18225,N_15521);
nor U20418 (N_20418,N_18840,N_19102);
and U20419 (N_20419,N_16679,N_19553);
nor U20420 (N_20420,N_15776,N_15542);
and U20421 (N_20421,N_18238,N_16516);
xnor U20422 (N_20422,N_18820,N_18714);
or U20423 (N_20423,N_15071,N_15858);
nor U20424 (N_20424,N_17672,N_18478);
nor U20425 (N_20425,N_15786,N_16161);
nor U20426 (N_20426,N_16156,N_18706);
nand U20427 (N_20427,N_17012,N_18993);
nor U20428 (N_20428,N_17345,N_17632);
nor U20429 (N_20429,N_15948,N_16346);
or U20430 (N_20430,N_15681,N_19599);
or U20431 (N_20431,N_15751,N_17508);
or U20432 (N_20432,N_18165,N_18267);
nand U20433 (N_20433,N_19101,N_17122);
and U20434 (N_20434,N_16319,N_19545);
xnor U20435 (N_20435,N_19131,N_15392);
or U20436 (N_20436,N_19449,N_18413);
or U20437 (N_20437,N_15881,N_19135);
or U20438 (N_20438,N_18253,N_15136);
and U20439 (N_20439,N_19665,N_15053);
xnor U20440 (N_20440,N_16840,N_15919);
and U20441 (N_20441,N_17550,N_19621);
nand U20442 (N_20442,N_19995,N_16450);
or U20443 (N_20443,N_17789,N_15054);
nand U20444 (N_20444,N_17308,N_15260);
nand U20445 (N_20445,N_15627,N_17000);
xor U20446 (N_20446,N_18246,N_17212);
nand U20447 (N_20447,N_19642,N_15104);
xnor U20448 (N_20448,N_16010,N_16261);
xnor U20449 (N_20449,N_16446,N_15036);
or U20450 (N_20450,N_19418,N_15041);
nand U20451 (N_20451,N_18724,N_18077);
and U20452 (N_20452,N_18151,N_17324);
or U20453 (N_20453,N_15710,N_15174);
nand U20454 (N_20454,N_17082,N_17694);
nor U20455 (N_20455,N_15389,N_17139);
xnor U20456 (N_20456,N_17194,N_15880);
nand U20457 (N_20457,N_15234,N_15195);
or U20458 (N_20458,N_15770,N_19504);
and U20459 (N_20459,N_15043,N_19748);
or U20460 (N_20460,N_19742,N_17609);
or U20461 (N_20461,N_15486,N_15491);
xor U20462 (N_20462,N_16143,N_19654);
or U20463 (N_20463,N_18507,N_18142);
or U20464 (N_20464,N_16269,N_15407);
and U20465 (N_20465,N_19182,N_18393);
and U20466 (N_20466,N_18043,N_17056);
xnor U20467 (N_20467,N_16379,N_15662);
xnor U20468 (N_20468,N_15151,N_15484);
nor U20469 (N_20469,N_17684,N_19960);
nor U20470 (N_20470,N_19110,N_19852);
xnor U20471 (N_20471,N_18245,N_16666);
or U20472 (N_20472,N_15178,N_18575);
nor U20473 (N_20473,N_19186,N_17702);
nor U20474 (N_20474,N_18491,N_19254);
and U20475 (N_20475,N_15114,N_18736);
and U20476 (N_20476,N_17088,N_17831);
or U20477 (N_20477,N_19096,N_15244);
and U20478 (N_20478,N_17458,N_19894);
nor U20479 (N_20479,N_16750,N_19407);
nor U20480 (N_20480,N_19751,N_19360);
or U20481 (N_20481,N_19937,N_18027);
xnor U20482 (N_20482,N_19417,N_18051);
xor U20483 (N_20483,N_15646,N_15825);
nand U20484 (N_20484,N_15495,N_16808);
nor U20485 (N_20485,N_15303,N_17989);
nor U20486 (N_20486,N_15593,N_16318);
or U20487 (N_20487,N_18979,N_18317);
nor U20488 (N_20488,N_19078,N_16440);
xor U20489 (N_20489,N_16946,N_18044);
nand U20490 (N_20490,N_19021,N_18809);
nand U20491 (N_20491,N_15175,N_19780);
or U20492 (N_20492,N_16100,N_17237);
nor U20493 (N_20493,N_17926,N_18255);
xnor U20494 (N_20494,N_15691,N_16169);
nor U20495 (N_20495,N_16529,N_17496);
and U20496 (N_20496,N_19929,N_17420);
nand U20497 (N_20497,N_19538,N_15213);
nor U20498 (N_20498,N_17911,N_17779);
and U20499 (N_20499,N_17026,N_19003);
and U20500 (N_20500,N_18743,N_17400);
and U20501 (N_20501,N_15942,N_17561);
and U20502 (N_20502,N_16870,N_15873);
nand U20503 (N_20503,N_16691,N_16943);
or U20504 (N_20504,N_16701,N_17872);
xnor U20505 (N_20505,N_15572,N_18321);
or U20506 (N_20506,N_19904,N_15226);
nand U20507 (N_20507,N_17914,N_19678);
xnor U20508 (N_20508,N_18520,N_17263);
xnor U20509 (N_20509,N_18305,N_19791);
or U20510 (N_20510,N_19222,N_18972);
or U20511 (N_20511,N_17460,N_16578);
nor U20512 (N_20512,N_15912,N_17556);
and U20513 (N_20513,N_19533,N_17174);
or U20514 (N_20514,N_19669,N_19025);
or U20515 (N_20515,N_18792,N_19060);
nand U20516 (N_20516,N_15085,N_15290);
nand U20517 (N_20517,N_18757,N_17224);
nand U20518 (N_20518,N_19215,N_16537);
nor U20519 (N_20519,N_18935,N_18316);
or U20520 (N_20520,N_18829,N_19348);
nor U20521 (N_20521,N_17130,N_19721);
or U20522 (N_20522,N_19867,N_18868);
nor U20523 (N_20523,N_16994,N_16040);
nor U20524 (N_20524,N_15850,N_15292);
and U20525 (N_20525,N_16656,N_17430);
nand U20526 (N_20526,N_16663,N_16928);
nor U20527 (N_20527,N_18986,N_18387);
or U20528 (N_20528,N_15707,N_16166);
or U20529 (N_20529,N_16596,N_18181);
or U20530 (N_20530,N_16923,N_19090);
and U20531 (N_20531,N_18671,N_15147);
or U20532 (N_20532,N_18149,N_15331);
nand U20533 (N_20533,N_17419,N_15516);
nor U20534 (N_20534,N_18068,N_19534);
nand U20535 (N_20535,N_19146,N_15709);
xor U20536 (N_20536,N_15032,N_15679);
xor U20537 (N_20537,N_18932,N_17634);
or U20538 (N_20538,N_19576,N_16417);
and U20539 (N_20539,N_16312,N_19340);
nor U20540 (N_20540,N_16436,N_16304);
nor U20541 (N_20541,N_17755,N_17511);
nor U20542 (N_20542,N_15559,N_17641);
or U20543 (N_20543,N_19455,N_17868);
nand U20544 (N_20544,N_19516,N_16485);
nand U20545 (N_20545,N_16787,N_18474);
nor U20546 (N_20546,N_17805,N_18897);
and U20547 (N_20547,N_17966,N_17241);
nor U20548 (N_20548,N_18561,N_18625);
xor U20549 (N_20549,N_16555,N_15993);
or U20550 (N_20550,N_18134,N_19687);
xor U20551 (N_20551,N_15026,N_17281);
nor U20552 (N_20552,N_15235,N_19803);
and U20553 (N_20553,N_17492,N_18034);
nor U20554 (N_20554,N_15004,N_15351);
nand U20555 (N_20555,N_19783,N_17775);
or U20556 (N_20556,N_18190,N_17044);
nor U20557 (N_20557,N_16563,N_15577);
nor U20558 (N_20558,N_16186,N_19684);
and U20559 (N_20559,N_16041,N_18713);
nor U20560 (N_20560,N_16758,N_16868);
xor U20561 (N_20561,N_19557,N_15251);
xor U20562 (N_20562,N_19477,N_17762);
and U20563 (N_20563,N_16327,N_15746);
nand U20564 (N_20564,N_15418,N_16467);
nor U20565 (N_20565,N_16232,N_18918);
nor U20566 (N_20566,N_19446,N_17340);
nand U20567 (N_20567,N_18239,N_19613);
nand U20568 (N_20568,N_18654,N_19681);
nand U20569 (N_20569,N_17201,N_19155);
xnor U20570 (N_20570,N_18567,N_16129);
and U20571 (N_20571,N_18206,N_16384);
and U20572 (N_20572,N_16372,N_16130);
nor U20573 (N_20573,N_19972,N_18588);
and U20574 (N_20574,N_15139,N_19197);
nand U20575 (N_20575,N_15079,N_16667);
xnor U20576 (N_20576,N_15722,N_17597);
or U20577 (N_20577,N_18053,N_16146);
nor U20578 (N_20578,N_16955,N_16722);
or U20579 (N_20579,N_16939,N_16909);
or U20580 (N_20580,N_18634,N_17877);
and U20581 (N_20581,N_18017,N_17735);
xor U20582 (N_20582,N_19760,N_18978);
nor U20583 (N_20583,N_19552,N_16675);
xor U20584 (N_20584,N_17199,N_16837);
or U20585 (N_20585,N_17127,N_16094);
nand U20586 (N_20586,N_15365,N_15347);
xor U20587 (N_20587,N_19148,N_15468);
xnor U20588 (N_20588,N_17657,N_17169);
xnor U20589 (N_20589,N_15007,N_15699);
nor U20590 (N_20590,N_15029,N_15449);
nand U20591 (N_20591,N_19611,N_15698);
and U20592 (N_20592,N_19465,N_18964);
and U20593 (N_20593,N_15767,N_15916);
nand U20594 (N_20594,N_16592,N_18359);
or U20595 (N_20595,N_19696,N_16002);
and U20596 (N_20596,N_18526,N_17838);
or U20597 (N_20597,N_17585,N_15337);
nor U20598 (N_20598,N_17764,N_19436);
or U20599 (N_20599,N_19992,N_19280);
nor U20600 (N_20600,N_16179,N_16924);
xor U20601 (N_20601,N_18331,N_16085);
or U20602 (N_20602,N_16886,N_17331);
or U20603 (N_20603,N_15374,N_15906);
or U20604 (N_20604,N_15532,N_15307);
nand U20605 (N_20605,N_17551,N_17171);
and U20606 (N_20606,N_19338,N_19408);
nand U20607 (N_20607,N_19435,N_17592);
and U20608 (N_20608,N_15313,N_19872);
nand U20609 (N_20609,N_16827,N_18196);
nand U20610 (N_20610,N_18175,N_15329);
nand U20611 (N_20611,N_16609,N_15323);
nor U20612 (N_20612,N_18330,N_15595);
nor U20613 (N_20613,N_18651,N_18201);
nand U20614 (N_20614,N_16992,N_19869);
xor U20615 (N_20615,N_15921,N_19295);
nand U20616 (N_20616,N_15403,N_19810);
nor U20617 (N_20617,N_18137,N_18062);
nand U20618 (N_20618,N_19724,N_16132);
xnor U20619 (N_20619,N_15992,N_16621);
xor U20620 (N_20620,N_15820,N_17077);
xor U20621 (N_20621,N_16523,N_17642);
and U20622 (N_20622,N_18570,N_15785);
xnor U20623 (N_20623,N_16266,N_16747);
or U20624 (N_20624,N_17306,N_19402);
xor U20625 (N_20625,N_15118,N_15675);
or U20626 (N_20626,N_16661,N_16477);
nor U20627 (N_20627,N_19768,N_17809);
nand U20628 (N_20628,N_15024,N_18475);
nand U20629 (N_20629,N_17682,N_19812);
nor U20630 (N_20630,N_15534,N_17944);
xor U20631 (N_20631,N_19536,N_19107);
or U20632 (N_20632,N_16342,N_19923);
nand U20633 (N_20633,N_18277,N_15011);
nand U20634 (N_20634,N_18822,N_16213);
xor U20635 (N_20635,N_15282,N_17606);
nand U20636 (N_20636,N_19203,N_15259);
or U20637 (N_20637,N_19345,N_15883);
nor U20638 (N_20638,N_19777,N_19038);
or U20639 (N_20639,N_15754,N_16706);
nor U20640 (N_20640,N_18646,N_19339);
nand U20641 (N_20641,N_17355,N_16454);
xnor U20642 (N_20642,N_15333,N_17343);
nand U20643 (N_20643,N_18078,N_16229);
xnor U20644 (N_20644,N_18723,N_19683);
and U20645 (N_20645,N_17653,N_15708);
nor U20646 (N_20646,N_16552,N_17733);
nand U20647 (N_20647,N_18187,N_17225);
or U20648 (N_20648,N_19214,N_16799);
and U20649 (N_20649,N_15546,N_18139);
xnor U20650 (N_20650,N_16500,N_18652);
and U20651 (N_20651,N_18606,N_17364);
xor U20652 (N_20652,N_18949,N_17670);
xnor U20653 (N_20653,N_15177,N_16672);
nor U20654 (N_20654,N_17074,N_17768);
xor U20655 (N_20655,N_16490,N_16307);
nand U20656 (N_20656,N_17918,N_15739);
nand U20657 (N_20657,N_15817,N_18900);
nand U20658 (N_20658,N_15692,N_19319);
and U20659 (N_20659,N_19264,N_17894);
or U20660 (N_20660,N_19085,N_15575);
xnor U20661 (N_20661,N_18544,N_15872);
and U20662 (N_20662,N_15048,N_16359);
and U20663 (N_20663,N_17783,N_17880);
nor U20664 (N_20664,N_18089,N_15752);
nand U20665 (N_20665,N_19892,N_19519);
nor U20666 (N_20666,N_16059,N_16671);
nand U20667 (N_20667,N_19314,N_16267);
nand U20668 (N_20668,N_15571,N_19705);
and U20669 (N_20669,N_17924,N_19164);
xnor U20670 (N_20670,N_17625,N_18543);
nor U20671 (N_20671,N_18343,N_19928);
or U20672 (N_20672,N_16912,N_15109);
nor U20673 (N_20673,N_16089,N_18339);
xor U20674 (N_20674,N_15953,N_15065);
xor U20675 (N_20675,N_19487,N_15614);
nor U20676 (N_20676,N_17638,N_16389);
and U20677 (N_20677,N_16459,N_18665);
xor U20678 (N_20678,N_15269,N_18908);
xnor U20679 (N_20679,N_18805,N_18283);
or U20680 (N_20680,N_17102,N_16918);
or U20681 (N_20681,N_17689,N_17066);
nand U20682 (N_20682,N_17017,N_19160);
and U20683 (N_20683,N_19730,N_18865);
xor U20684 (N_20684,N_17411,N_18300);
nor U20685 (N_20685,N_16429,N_16931);
and U20686 (N_20686,N_16184,N_15312);
nor U20687 (N_20687,N_15836,N_17317);
nand U20688 (N_20688,N_15349,N_15951);
nand U20689 (N_20689,N_17485,N_18066);
nand U20690 (N_20690,N_17624,N_17298);
nand U20691 (N_20691,N_17366,N_19244);
or U20692 (N_20692,N_16710,N_16772);
nor U20693 (N_20693,N_19326,N_19054);
or U20694 (N_20694,N_15736,N_17276);
and U20695 (N_20695,N_18367,N_17068);
xor U20696 (N_20696,N_17981,N_17957);
nand U20697 (N_20697,N_17905,N_19692);
nor U20698 (N_20698,N_15356,N_19448);
xnor U20699 (N_20699,N_17598,N_17879);
nor U20700 (N_20700,N_15338,N_19680);
or U20701 (N_20701,N_18523,N_18158);
xor U20702 (N_20702,N_15732,N_18296);
and U20703 (N_20703,N_18020,N_16114);
nand U20704 (N_20704,N_19127,N_16541);
or U20705 (N_20705,N_19558,N_17252);
nand U20706 (N_20706,N_17418,N_15763);
nor U20707 (N_20707,N_17189,N_19893);
xor U20708 (N_20708,N_18038,N_18070);
nor U20709 (N_20709,N_16395,N_17720);
or U20710 (N_20710,N_19579,N_17104);
and U20711 (N_20711,N_15131,N_15492);
or U20712 (N_20712,N_19594,N_16748);
or U20713 (N_20713,N_19028,N_18831);
or U20714 (N_20714,N_17289,N_15829);
nor U20715 (N_20715,N_18318,N_19573);
xnor U20716 (N_20716,N_15876,N_17972);
xor U20717 (N_20717,N_18282,N_16565);
nor U20718 (N_20718,N_17958,N_18144);
and U20719 (N_20719,N_18755,N_16370);
and U20720 (N_20720,N_18382,N_18891);
nand U20721 (N_20721,N_18775,N_15005);
xnor U20722 (N_20722,N_17920,N_18917);
xnor U20723 (N_20723,N_16066,N_18892);
nor U20724 (N_20724,N_17013,N_15181);
xnor U20725 (N_20725,N_16356,N_16983);
nor U20726 (N_20726,N_17454,N_15959);
xnor U20727 (N_20727,N_19382,N_19439);
and U20728 (N_20728,N_15354,N_15581);
xor U20729 (N_20729,N_19169,N_18495);
nor U20730 (N_20730,N_16869,N_18962);
nor U20731 (N_20731,N_17045,N_18425);
xnor U20732 (N_20732,N_18683,N_18036);
xor U20733 (N_20733,N_19474,N_17043);
or U20734 (N_20734,N_19380,N_15957);
or U20735 (N_20735,N_18877,N_16098);
and U20736 (N_20736,N_18341,N_18374);
xnor U20737 (N_20737,N_18951,N_16614);
nand U20738 (N_20738,N_19480,N_17322);
nor U20739 (N_20739,N_18030,N_19914);
xnor U20740 (N_20740,N_17399,N_19634);
or U20741 (N_20741,N_17997,N_16813);
and U20742 (N_20742,N_17336,N_18735);
and U20743 (N_20743,N_18319,N_16585);
nor U20744 (N_20744,N_15513,N_16214);
xnor U20745 (N_20745,N_18260,N_15467);
nor U20746 (N_20746,N_19979,N_18047);
xor U20747 (N_20747,N_15545,N_18697);
nor U20748 (N_20748,N_18855,N_18479);
xnor U20749 (N_20749,N_16783,N_19587);
nor U20750 (N_20750,N_18688,N_19822);
nand U20751 (N_20751,N_19184,N_19800);
nor U20752 (N_20752,N_15308,N_18784);
and U20753 (N_20753,N_17413,N_19017);
and U20754 (N_20754,N_19443,N_16455);
nor U20755 (N_20755,N_18484,N_17369);
and U20756 (N_20756,N_15276,N_19514);
and U20757 (N_20757,N_17976,N_17046);
nand U20758 (N_20758,N_19547,N_19217);
or U20759 (N_20759,N_15925,N_15676);
and U20760 (N_20760,N_16222,N_17011);
xnor U20761 (N_20761,N_18217,N_17462);
and U20762 (N_20762,N_19136,N_17933);
and U20763 (N_20763,N_15340,N_15855);
or U20764 (N_20764,N_16855,N_19660);
or U20765 (N_20765,N_16014,N_17260);
and U20766 (N_20766,N_19583,N_17985);
and U20767 (N_20767,N_19069,N_17941);
and U20768 (N_20768,N_15950,N_19353);
and U20769 (N_20769,N_18412,N_16687);
nand U20770 (N_20770,N_17097,N_19111);
nor U20771 (N_20771,N_18630,N_18816);
nand U20772 (N_20772,N_17396,N_15558);
and U20773 (N_20773,N_18009,N_15295);
and U20774 (N_20774,N_16726,N_16850);
and U20775 (N_20775,N_18519,N_19746);
nand U20776 (N_20776,N_18123,N_18154);
xor U20777 (N_20777,N_17294,N_16574);
nand U20778 (N_20778,N_17692,N_15826);
nor U20779 (N_20779,N_15731,N_17255);
xor U20780 (N_20780,N_15750,N_15355);
xnor U20781 (N_20781,N_15196,N_18242);
xor U20782 (N_20782,N_19277,N_17299);
nor U20783 (N_20783,N_18733,N_16652);
xnor U20784 (N_20784,N_19309,N_16498);
nand U20785 (N_20785,N_19638,N_19562);
xor U20786 (N_20786,N_15503,N_16538);
xnor U20787 (N_20787,N_16362,N_19027);
nor U20788 (N_20788,N_18902,N_15841);
or U20789 (N_20789,N_15868,N_16631);
and U20790 (N_20790,N_16601,N_16479);
nand U20791 (N_20791,N_19303,N_19347);
nor U20792 (N_20792,N_16244,N_19016);
nor U20793 (N_20793,N_16823,N_18228);
nand U20794 (N_20794,N_19565,N_15428);
nor U20795 (N_20795,N_19335,N_19113);
nand U20796 (N_20796,N_15087,N_19632);
or U20797 (N_20797,N_17934,N_18163);
nor U20798 (N_20798,N_17353,N_15523);
xnor U20799 (N_20799,N_15533,N_18361);
or U20800 (N_20800,N_17857,N_16651);
and U20801 (N_20801,N_17820,N_15649);
or U20802 (N_20802,N_19566,N_19505);
xor U20803 (N_20803,N_15128,N_17426);
or U20804 (N_20804,N_19055,N_19789);
nor U20805 (N_20805,N_16877,N_19063);
and U20806 (N_20806,N_16151,N_17737);
xnor U20807 (N_20807,N_17785,N_17864);
nor U20808 (N_20808,N_17705,N_16238);
or U20809 (N_20809,N_15155,N_18060);
xor U20810 (N_20810,N_18428,N_19249);
and U20811 (N_20811,N_16334,N_19664);
or U20812 (N_20812,N_16325,N_15462);
xnor U20813 (N_20813,N_15828,N_18383);
or U20814 (N_20814,N_15369,N_19804);
xor U20815 (N_20815,N_15327,N_16134);
and U20816 (N_20816,N_15098,N_18961);
or U20817 (N_20817,N_15366,N_16260);
nor U20818 (N_20818,N_16664,N_16575);
or U20819 (N_20819,N_18766,N_18777);
and U20820 (N_20820,N_18336,N_16293);
and U20821 (N_20821,N_19813,N_18661);
nand U20822 (N_20822,N_15748,N_18045);
xnor U20823 (N_20823,N_16873,N_19647);
nand U20824 (N_20824,N_17062,N_19709);
xnor U20825 (N_20825,N_19805,N_19649);
nand U20826 (N_20826,N_16008,N_15204);
and U20827 (N_20827,N_18039,N_18109);
and U20828 (N_20828,N_16043,N_18366);
or U20829 (N_20829,N_17089,N_16252);
or U20830 (N_20830,N_19020,N_15777);
nand U20831 (N_20831,N_19582,N_18956);
or U20832 (N_20832,N_18682,N_19577);
or U20833 (N_20833,N_17031,N_15771);
nand U20834 (N_20834,N_15557,N_15643);
xnor U20835 (N_20835,N_18555,N_16427);
xor U20836 (N_20836,N_15013,N_15682);
nor U20837 (N_20837,N_16841,N_17152);
and U20838 (N_20838,N_17628,N_17206);
nor U20839 (N_20839,N_15246,N_18008);
or U20840 (N_20840,N_19779,N_18350);
or U20841 (N_20841,N_19947,N_19051);
or U20842 (N_20842,N_17761,N_19341);
xor U20843 (N_20843,N_17586,N_16969);
and U20844 (N_20844,N_19636,N_19677);
and U20845 (N_20845,N_19877,N_17098);
nor U20846 (N_20846,N_17193,N_19306);
or U20847 (N_20847,N_16121,N_19073);
xnor U20848 (N_20848,N_19796,N_16849);
xor U20849 (N_20849,N_16422,N_16273);
and U20850 (N_20850,N_17461,N_17572);
nand U20851 (N_20851,N_17782,N_18449);
or U20852 (N_20852,N_18025,N_17211);
nand U20853 (N_20853,N_19802,N_18673);
or U20854 (N_20854,N_17921,N_15058);
and U20855 (N_20855,N_19425,N_18421);
nor U20856 (N_20856,N_19615,N_19130);
or U20857 (N_20857,N_18452,N_16268);
or U20858 (N_20858,N_18329,N_15642);
or U20859 (N_20859,N_16209,N_18889);
nor U20860 (N_20860,N_17473,N_15112);
nor U20861 (N_20861,N_19253,N_18658);
xnor U20862 (N_20862,N_18241,N_18271);
nand U20863 (N_20863,N_17416,N_15049);
xnor U20864 (N_20864,N_18046,N_19963);
nor U20865 (N_20865,N_17029,N_15040);
nand U20866 (N_20866,N_17856,N_17154);
and U20867 (N_20867,N_15874,N_17569);
nand U20868 (N_20868,N_16390,N_18762);
or U20869 (N_20869,N_16093,N_18256);
nor U20870 (N_20870,N_19736,N_16189);
nor U20871 (N_20871,N_15481,N_17841);
nor U20872 (N_20872,N_18955,N_17470);
and U20873 (N_20873,N_18363,N_16527);
nor U20874 (N_20874,N_16300,N_18456);
nor U20875 (N_20875,N_16597,N_15056);
nor U20876 (N_20876,N_17157,N_18942);
or U20877 (N_20877,N_18014,N_17599);
nand U20878 (N_20878,N_18882,N_18592);
nand U20879 (N_20879,N_16357,N_18390);
and U20880 (N_20880,N_18795,N_18616);
or U20881 (N_20881,N_19031,N_18303);
or U20882 (N_20882,N_17747,N_18872);
or U20883 (N_20883,N_17001,N_15666);
and U20884 (N_20884,N_19957,N_18852);
nand U20885 (N_20885,N_17048,N_15540);
xnor U20886 (N_20886,N_18183,N_15410);
or U20887 (N_20887,N_19061,N_18365);
nand U20888 (N_20888,N_17751,N_16942);
xnor U20889 (N_20889,N_16295,N_16903);
and U20890 (N_20890,N_19374,N_15733);
xor U20891 (N_20891,N_19695,N_19271);
or U20892 (N_20892,N_15562,N_17903);
nand U20893 (N_20893,N_17874,N_17790);
nand U20894 (N_20894,N_17041,N_18845);
nor U20895 (N_20895,N_18954,N_16496);
or U20896 (N_20896,N_19291,N_18549);
nor U20897 (N_20897,N_17951,N_17619);
and U20898 (N_20898,N_15133,N_18719);
or U20899 (N_20899,N_18284,N_16368);
and U20900 (N_20900,N_19974,N_15167);
and U20901 (N_20901,N_15660,N_19324);
and U20902 (N_20902,N_19527,N_17582);
xnor U20903 (N_20903,N_15134,N_18049);
xor U20904 (N_20904,N_18712,N_16879);
xnor U20905 (N_20905,N_15402,N_15943);
xnor U20906 (N_20906,N_15062,N_16398);
and U20907 (N_20907,N_18907,N_18515);
and U20908 (N_20908,N_18802,N_18572);
nor U20909 (N_20909,N_18120,N_15172);
nand U20910 (N_20910,N_19986,N_17899);
or U20911 (N_20911,N_15179,N_16899);
nand U20912 (N_20912,N_15206,N_15127);
nor U20913 (N_20913,N_18672,N_17685);
nor U20914 (N_20914,N_16626,N_19420);
nor U20915 (N_20915,N_18768,N_17925);
xor U20916 (N_20916,N_19776,N_17033);
and U20917 (N_20917,N_17214,N_19593);
and U20918 (N_20918,N_16864,N_17594);
and U20919 (N_20919,N_18657,N_17491);
and U20920 (N_20920,N_19641,N_17190);
and U20921 (N_20921,N_17984,N_19413);
or U20922 (N_20922,N_18010,N_16084);
nand U20923 (N_20923,N_17866,N_15416);
nand U20924 (N_20924,N_18582,N_19901);
or U20925 (N_20925,N_17853,N_19082);
or U20926 (N_20926,N_15877,N_15897);
xnor U20927 (N_20927,N_17833,N_16534);
xnor U20928 (N_20928,N_16629,N_16519);
nor U20929 (N_20929,N_16476,N_19520);
xor U20930 (N_20930,N_18811,N_19041);
nor U20931 (N_20931,N_18458,N_19002);
xnor U20932 (N_20932,N_15264,N_18487);
nor U20933 (N_20933,N_19030,N_19971);
or U20934 (N_20934,N_18557,N_17391);
nor U20935 (N_20935,N_18441,N_17363);
nor U20936 (N_20936,N_18871,N_17686);
and U20937 (N_20937,N_16407,N_18769);
or U20938 (N_20938,N_19207,N_15932);
nand U20939 (N_20939,N_15446,N_19601);
and U20940 (N_20940,N_15724,N_18325);
nor U20941 (N_20941,N_19058,N_16199);
xor U20942 (N_20942,N_18756,N_16270);
nand U20943 (N_20943,N_18801,N_16677);
and U20944 (N_20944,N_16796,N_18804);
or U20945 (N_20945,N_16723,N_16061);
nand U20946 (N_20946,N_18052,N_18689);
nor U20947 (N_20947,N_19119,N_17502);
xnor U20948 (N_20948,N_15570,N_19496);
and U20949 (N_20949,N_19285,N_16289);
nor U20950 (N_20950,N_17415,N_18761);
xor U20951 (N_20951,N_15616,N_16817);
and U20952 (N_20952,N_15411,N_16863);
xnor U20953 (N_20953,N_18886,N_19248);
nor U20954 (N_20954,N_16254,N_18600);
xnor U20955 (N_20955,N_15069,N_17140);
nor U20956 (N_20956,N_19616,N_16299);
or U20957 (N_20957,N_18204,N_17734);
or U20958 (N_20958,N_18191,N_19617);
or U20959 (N_20959,N_16004,N_15937);
nand U20960 (N_20960,N_17602,N_17236);
and U20961 (N_20961,N_15378,N_18710);
nand U20962 (N_20962,N_16022,N_15207);
and U20963 (N_20963,N_17711,N_19227);
or U20964 (N_20964,N_17631,N_15238);
and U20965 (N_20965,N_15999,N_17605);
nor U20966 (N_20966,N_19190,N_19422);
or U20967 (N_20967,N_16550,N_16294);
and U20968 (N_20968,N_19754,N_15001);
nor U20969 (N_20969,N_16556,N_15500);
nand U20970 (N_20970,N_19473,N_15436);
or U20971 (N_20971,N_19969,N_15146);
and U20972 (N_20972,N_19013,N_17887);
and U20973 (N_20973,N_19034,N_19263);
or U20974 (N_20974,N_19744,N_16938);
and U20975 (N_20975,N_15383,N_16716);
xnor U20976 (N_20976,N_15076,N_16761);
nand U20977 (N_20977,N_17668,N_18141);
nor U20978 (N_20978,N_19755,N_15170);
xor U20979 (N_20979,N_16391,N_18656);
nand U20980 (N_20980,N_18442,N_17379);
and U20981 (N_20981,N_17912,N_18063);
nor U20982 (N_20982,N_17103,N_19956);
nor U20983 (N_20983,N_19497,N_16888);
nand U20984 (N_20984,N_17218,N_15603);
or U20985 (N_20985,N_18208,N_16800);
and U20986 (N_20986,N_19725,N_18945);
xnor U20987 (N_20987,N_18410,N_19376);
nor U20988 (N_20988,N_18485,N_19715);
nor U20989 (N_20989,N_16082,N_18326);
or U20990 (N_20990,N_19629,N_15725);
or U20991 (N_20991,N_15294,N_19412);
and U20992 (N_20992,N_17987,N_15989);
nand U20993 (N_20993,N_19478,N_16511);
nand U20994 (N_20994,N_18601,N_19686);
nand U20995 (N_20995,N_15375,N_17652);
and U20996 (N_20996,N_18750,N_17915);
nor U20997 (N_20997,N_18711,N_17205);
nor U20998 (N_20998,N_18645,N_18925);
xor U20999 (N_20999,N_17840,N_18180);
nand U21000 (N_21000,N_15857,N_17495);
or U21001 (N_21001,N_18483,N_19178);
and U21002 (N_21002,N_17745,N_18403);
nand U21003 (N_21003,N_17991,N_19946);
or U21004 (N_21004,N_19500,N_15271);
nand U21005 (N_21005,N_17608,N_15214);
nand U21006 (N_21006,N_16792,N_15086);
and U21007 (N_21007,N_18211,N_18641);
or U21008 (N_21008,N_17161,N_15176);
nand U21009 (N_21009,N_17770,N_16341);
and U21010 (N_21010,N_18623,N_18628);
and U21011 (N_21011,N_15208,N_15671);
or U21012 (N_21012,N_17121,N_17643);
or U21013 (N_21013,N_17960,N_15262);
xor U21014 (N_21014,N_15654,N_15130);
nand U21015 (N_21015,N_16366,N_18617);
nor U21016 (N_21016,N_16566,N_19655);
nand U21017 (N_21017,N_16301,N_15930);
nor U21018 (N_21018,N_17808,N_18240);
nand U21019 (N_21019,N_19083,N_19297);
and U21020 (N_21020,N_19606,N_19328);
and U21021 (N_21021,N_16431,N_16548);
or U21022 (N_21022,N_17659,N_16639);
and U21023 (N_21023,N_18894,N_15211);
nor U21024 (N_21024,N_16893,N_19915);
and U21025 (N_21025,N_16530,N_19389);
xnor U21026 (N_21026,N_17195,N_17837);
nand U21027 (N_21027,N_15019,N_18911);
and U21028 (N_21028,N_16502,N_18807);
nor U21029 (N_21029,N_19044,N_15902);
or U21030 (N_21030,N_16339,N_16641);
and U21031 (N_21031,N_19262,N_19675);
and U21032 (N_21032,N_15050,N_19048);
nand U21033 (N_21033,N_15910,N_18622);
nor U21034 (N_21034,N_17437,N_15981);
and U21035 (N_21035,N_18265,N_16200);
xnor U21036 (N_21036,N_19851,N_16401);
or U21037 (N_21037,N_16045,N_17855);
nor U21038 (N_21038,N_19126,N_19820);
and U21039 (N_21039,N_18076,N_15460);
and U21040 (N_21040,N_19100,N_16540);
nand U21041 (N_21041,N_19670,N_15547);
nand U21042 (N_21042,N_16765,N_17869);
nor U21043 (N_21043,N_17268,N_18844);
nand U21044 (N_21044,N_19870,N_19844);
nand U21045 (N_21045,N_18385,N_16206);
nor U21046 (N_21046,N_17285,N_18113);
and U21047 (N_21047,N_19771,N_16757);
or U21048 (N_21048,N_15105,N_16243);
xnor U21049 (N_21049,N_18450,N_17539);
xor U21050 (N_21050,N_19440,N_16154);
nand U21051 (N_21051,N_15783,N_18391);
nand U21052 (N_21052,N_16081,N_19652);
nor U21053 (N_21053,N_19761,N_19183);
nand U21054 (N_21054,N_17019,N_17518);
xnor U21055 (N_21055,N_18005,N_15442);
xor U21056 (N_21056,N_17356,N_18862);
and U21057 (N_21057,N_16458,N_17640);
nand U21058 (N_21058,N_17695,N_17825);
nand U21059 (N_21059,N_15189,N_16999);
nor U21060 (N_21060,N_17488,N_17208);
nor U21061 (N_21061,N_19188,N_18839);
xnor U21062 (N_21062,N_18224,N_18793);
and U21063 (N_21063,N_17040,N_16352);
or U21064 (N_21064,N_16171,N_17627);
and U21065 (N_21065,N_15090,N_16598);
xnor U21066 (N_21066,N_18414,N_15309);
or U21067 (N_21067,N_15441,N_15153);
nor U21068 (N_21068,N_19592,N_19808);
nor U21069 (N_21069,N_18408,N_18003);
nand U21070 (N_21070,N_17404,N_16448);
xnor U21071 (N_21071,N_15107,N_17125);
xnor U21072 (N_21072,N_17562,N_18409);
and U21073 (N_21073,N_15518,N_19236);
nand U21074 (N_21074,N_19517,N_15399);
xnor U21075 (N_21075,N_18875,N_19917);
nor U21076 (N_21076,N_16126,N_18090);
or U21077 (N_21077,N_17615,N_15267);
xor U21078 (N_21078,N_17620,N_16780);
nor U21079 (N_21079,N_17131,N_18528);
nand U21080 (N_21080,N_15106,N_17565);
or U21081 (N_21081,N_15311,N_19349);
nor U21082 (N_21082,N_19393,N_18108);
and U21083 (N_21083,N_18505,N_17457);
and U21084 (N_21084,N_15461,N_19268);
xnor U21085 (N_21085,N_19792,N_16478);
and U21086 (N_21086,N_18244,N_18832);
nor U21087 (N_21087,N_16018,N_15719);
or U21088 (N_21088,N_16654,N_15165);
and U21089 (N_21089,N_16035,N_18904);
and U21090 (N_21090,N_17445,N_17338);
xor U21091 (N_21091,N_19722,N_16774);
and U21092 (N_21092,N_18035,N_15316);
and U21093 (N_21093,N_15911,N_15539);
xnor U21094 (N_21094,N_16582,N_17573);
xnor U21095 (N_21095,N_16047,N_19728);
or U21096 (N_21096,N_16241,N_19157);
nor U21097 (N_21097,N_18746,N_16791);
xnor U21098 (N_21098,N_15223,N_16510);
and U21099 (N_21099,N_19734,N_15927);
xnor U21100 (N_21100,N_15803,N_17253);
xor U21101 (N_21101,N_16128,N_15899);
and U21102 (N_21102,N_17580,N_16880);
nand U21103 (N_21103,N_17020,N_15376);
and U21104 (N_21104,N_17407,N_15808);
xor U21105 (N_21105,N_17507,N_18727);
or U21106 (N_21106,N_19392,N_17752);
nand U21107 (N_21107,N_16590,N_16858);
nor U21108 (N_21108,N_15788,N_16250);
nand U21109 (N_21109,N_15297,N_15990);
xnor U21110 (N_21110,N_17262,N_16257);
nand U21111 (N_21111,N_16461,N_19067);
nor U21112 (N_21112,N_15923,N_19862);
or U21113 (N_21113,N_19667,N_19467);
nor U21114 (N_21114,N_16913,N_16145);
nand U21115 (N_21115,N_17233,N_16009);
and U21116 (N_21116,N_15296,N_18169);
nand U21117 (N_21117,N_15607,N_19346);
or U21118 (N_21118,N_15250,N_18853);
xor U21119 (N_21119,N_18939,N_17153);
nor U21120 (N_21120,N_16567,N_17493);
nand U21121 (N_21121,N_18827,N_17683);
or U21122 (N_21122,N_16023,N_18111);
and U21123 (N_21123,N_18817,N_16997);
and U21124 (N_21124,N_16079,N_19129);
nor U21125 (N_21125,N_18580,N_17886);
nor U21126 (N_21126,N_17436,N_19814);
or U21127 (N_21127,N_19334,N_15972);
nand U21128 (N_21128,N_19596,N_19922);
nor U21129 (N_21129,N_17816,N_15842);
xnor U21130 (N_21130,N_16889,N_16668);
nor U21131 (N_21131,N_19826,N_16778);
nor U21132 (N_21132,N_18896,N_17714);
nor U21133 (N_21133,N_18699,N_19507);
or U21134 (N_21134,N_16892,N_15908);
nand U21135 (N_21135,N_19218,N_17708);
or U21136 (N_21136,N_15015,N_18262);
nand U21137 (N_21137,N_19907,N_18198);
and U21138 (N_21138,N_17583,N_19727);
and U21139 (N_21139,N_16753,N_19381);
xnor U21140 (N_21140,N_16662,N_16460);
and U21141 (N_21141,N_16297,N_15431);
nor U21142 (N_21142,N_19561,N_16245);
nand U21143 (N_21143,N_17429,N_16642);
nand U21144 (N_21144,N_18298,N_17483);
and U21145 (N_21145,N_18073,N_17160);
nand U21146 (N_21146,N_18797,N_17439);
nand U21147 (N_21147,N_19091,N_17095);
nand U21148 (N_21148,N_19965,N_17543);
or U21149 (N_21149,N_19321,N_18734);
nand U21150 (N_21150,N_15258,N_17528);
nand U21151 (N_21151,N_18739,N_15888);
nand U21152 (N_21152,N_16277,N_19406);
nand U21153 (N_21153,N_19233,N_18621);
or U21154 (N_21154,N_18302,N_18531);
nor U21155 (N_21155,N_18327,N_18577);
nand U21156 (N_21156,N_15640,N_19980);
or U21157 (N_21157,N_19646,N_15194);
xnor U21158 (N_21158,N_17962,N_17749);
and U21159 (N_21159,N_18648,N_18607);
and U21160 (N_21160,N_19982,N_15487);
nand U21161 (N_21161,N_16728,N_18684);
and U21162 (N_21162,N_17209,N_17478);
or U21163 (N_21163,N_18963,N_15849);
nand U21164 (N_21164,N_18268,N_17374);
xnor U21165 (N_21165,N_15582,N_15445);
xor U21166 (N_21166,N_19839,N_17110);
nor U21167 (N_21167,N_16442,N_18221);
xnor U21168 (N_21168,N_15443,N_18215);
xor U21169 (N_21169,N_15798,N_19076);
xnor U21170 (N_21170,N_18927,N_19879);
and U21171 (N_21171,N_16298,N_19795);
or U21172 (N_21172,N_15924,N_15447);
nand U21173 (N_21173,N_16067,N_15851);
or U21174 (N_21174,N_17382,N_15895);
nand U21175 (N_21175,N_19624,N_16311);
nand U21176 (N_21176,N_16520,N_17349);
xnor U21177 (N_21177,N_17548,N_15852);
xnor U21178 (N_21178,N_19486,N_17388);
nand U21179 (N_21179,N_19428,N_15810);
nand U21180 (N_21180,N_17344,N_19187);
and U21181 (N_21181,N_18708,N_18812);
nor U21182 (N_21182,N_15787,N_17758);
nand U21183 (N_21183,N_17371,N_17637);
and U21184 (N_21184,N_15653,N_16802);
or U21185 (N_21185,N_18274,N_16806);
nand U21186 (N_21186,N_17636,N_15680);
and U21187 (N_21187,N_18362,N_17325);
nand U21188 (N_21188,N_15819,N_16444);
nand U21189 (N_21189,N_18291,N_15306);
and U21190 (N_21190,N_15444,N_19518);
nand U21191 (N_21191,N_15490,N_17537);
nor U21192 (N_21192,N_17765,N_19718);
xnor U21193 (N_21193,N_15265,N_19379);
or U21194 (N_21194,N_17992,N_16388);
nor U21195 (N_21195,N_17469,N_18873);
nand U21196 (N_21196,N_18258,N_17178);
or U21197 (N_21197,N_15008,N_19716);
nand U21198 (N_21198,N_19312,N_15476);
nand U21199 (N_21199,N_17955,N_15565);
or U21200 (N_21200,N_15869,N_18629);
nor U21201 (N_21201,N_19975,N_15463);
nor U21202 (N_21202,N_15882,N_17896);
or U21203 (N_21203,N_18006,N_16078);
or U21204 (N_21204,N_16329,N_19836);
nand U21205 (N_21205,N_15718,N_17142);
nand U21206 (N_21206,N_17919,N_16324);
nand U21207 (N_21207,N_18938,N_18846);
or U21208 (N_21208,N_18922,N_18420);
or U21209 (N_21209,N_15969,N_15845);
xnor U21210 (N_21210,N_15344,N_16149);
nand U21211 (N_21211,N_15994,N_19887);
or U21212 (N_21212,N_19905,N_16385);
nor U21213 (N_21213,N_15913,N_17115);
or U21214 (N_21214,N_17693,N_17673);
nand U21215 (N_21215,N_19861,N_17618);
nand U21216 (N_21216,N_15157,N_15456);
nand U21217 (N_21217,N_16465,N_17522);
nand U21218 (N_21218,N_18269,N_17612);
nand U21219 (N_21219,N_15077,N_16021);
xnor U21220 (N_21220,N_17452,N_15781);
or U21221 (N_21221,N_15398,N_18685);
nor U21222 (N_21222,N_15530,N_15892);
xor U21223 (N_21223,N_17347,N_15552);
or U21224 (N_21224,N_18394,N_15432);
or U21225 (N_21225,N_17639,N_18299);
xnor U21226 (N_21226,N_15854,N_19657);
or U21227 (N_21227,N_15059,N_18088);
xor U21228 (N_21228,N_19311,N_16223);
or U21229 (N_21229,N_18322,N_15101);
nor U21230 (N_21230,N_18771,N_18899);
xor U21231 (N_21231,N_18737,N_18958);
nand U21232 (N_21232,N_19759,N_19074);
or U21233 (N_21233,N_17849,N_18019);
nor U21234 (N_21234,N_15126,N_19739);
and U21235 (N_21235,N_17069,N_18454);
xor U21236 (N_21236,N_17105,N_18533);
nand U21237 (N_21237,N_16220,N_16439);
or U21238 (N_21238,N_16705,N_18933);
or U21239 (N_21239,N_16246,N_15064);
nor U21240 (N_21240,N_17982,N_16103);
xor U21241 (N_21241,N_17814,N_17286);
and U21242 (N_21242,N_15573,N_18085);
nor U21243 (N_21243,N_15478,N_17953);
nor U21244 (N_21244,N_18681,N_19876);
nand U21245 (N_21245,N_18222,N_17304);
or U21246 (N_21246,N_15765,N_19619);
and U21247 (N_21247,N_18765,N_18397);
xnor U21248 (N_21248,N_19471,N_19009);
xnor U21249 (N_21249,N_15494,N_19959);
or U21250 (N_21250,N_17109,N_19199);
xnor U21251 (N_21251,N_17137,N_17361);
nand U21252 (N_21252,N_18841,N_15568);
xnor U21253 (N_21253,N_17736,N_19491);
and U21254 (N_21254,N_16344,N_15278);
xor U21255 (N_21255,N_19149,N_15713);
nand U21256 (N_21256,N_19099,N_17293);
nand U21257 (N_21257,N_15067,N_18488);
nor U21258 (N_21258,N_16487,N_19738);
or U21259 (N_21259,N_19551,N_16308);
nand U21260 (N_21260,N_16770,N_17959);
and U21261 (N_21261,N_19745,N_15980);
nor U21262 (N_21262,N_17179,N_16976);
xor U21263 (N_21263,N_15123,N_17081);
nand U21264 (N_21264,N_18920,N_16944);
xnor U21265 (N_21265,N_16127,N_19546);
nor U21266 (N_21266,N_18058,N_17750);
nor U21267 (N_21267,N_16948,N_15541);
xnor U21268 (N_21268,N_17487,N_15068);
nand U21269 (N_21269,N_17145,N_16468);
nor U21270 (N_21270,N_18959,N_19953);
nand U21271 (N_21271,N_17226,N_18975);
nor U21272 (N_21272,N_18332,N_16572);
or U21273 (N_21273,N_18493,N_18659);
and U21274 (N_21274,N_16474,N_18067);
or U21275 (N_21275,N_15116,N_15971);
or U21276 (N_21276,N_17124,N_17848);
xnor U21277 (N_21277,N_16361,N_15321);
nor U21278 (N_21278,N_19717,N_19204);
nand U21279 (N_21279,N_18854,N_19673);
and U21280 (N_21280,N_16940,N_16409);
nand U21281 (N_21281,N_17428,N_15938);
nor U21282 (N_21282,N_17538,N_19554);
nor U21283 (N_21283,N_15983,N_16562);
nor U21284 (N_21284,N_16788,N_15979);
nor U21285 (N_21285,N_18633,N_18287);
nor U21286 (N_21286,N_16648,N_16699);
nor U21287 (N_21287,N_18609,N_19181);
nand U21288 (N_21288,N_16702,N_15674);
nand U21289 (N_21289,N_17644,N_19137);
nand U21290 (N_21290,N_17738,N_16367);
nor U21291 (N_21291,N_19292,N_17394);
nand U21292 (N_21292,N_16731,N_18690);
nand U21293 (N_21293,N_19524,N_19232);
or U21294 (N_21294,N_18794,N_17288);
or U21295 (N_21295,N_15371,N_16434);
nand U21296 (N_21296,N_16321,N_15027);
and U21297 (N_21297,N_18751,N_15758);
and U21298 (N_21298,N_15685,N_17060);
or U21299 (N_21299,N_19433,N_17815);
xnor U21300 (N_21300,N_16058,N_15665);
nand U21301 (N_21301,N_19024,N_15529);
and U21302 (N_21302,N_15420,N_16227);
or U21303 (N_21303,N_19584,N_15509);
xnor U21304 (N_21304,N_19535,N_17946);
or U21305 (N_21305,N_15686,N_19170);
nand U21306 (N_21306,N_15115,N_19840);
nor U21307 (N_21307,N_15859,N_17375);
xor U21308 (N_21308,N_17576,N_19057);
xor U21309 (N_21309,N_17027,N_15567);
nor U21310 (N_21310,N_17055,N_19868);
nand U21311 (N_21311,N_18836,N_19878);
or U21312 (N_21312,N_19322,N_16608);
or U21313 (N_21313,N_18237,N_16584);
and U21314 (N_21314,N_16820,N_16698);
xnor U21315 (N_21315,N_17725,N_19499);
and U21316 (N_21316,N_18772,N_15944);
nand U21317 (N_21317,N_17756,N_18133);
xor U21318 (N_21318,N_16755,N_18890);
xnor U21319 (N_21319,N_19106,N_17587);
nand U21320 (N_21320,N_17287,N_17433);
and U21321 (N_21321,N_17945,N_17531);
and U21322 (N_21322,N_19084,N_17453);
nor U21323 (N_21323,N_17527,N_17384);
nand U21324 (N_21324,N_17658,N_18948);
xnor U21325 (N_21325,N_18563,N_17389);
and U21326 (N_21326,N_16069,N_17063);
nand U21327 (N_21327,N_15280,N_17296);
and U21328 (N_21328,N_15148,N_19095);
nand U21329 (N_21329,N_18368,N_18431);
xnor U21330 (N_21330,N_16709,N_16839);
nand U21331 (N_21331,N_15853,N_15789);
and U21332 (N_21332,N_19610,N_19008);
nand U21333 (N_21333,N_19618,N_15898);
nand U21334 (N_21334,N_17129,N_15970);
or U21335 (N_21335,N_18931,N_15866);
or U21336 (N_21336,N_17406,N_18132);
and U21337 (N_21337,N_19354,N_15239);
xor U21338 (N_21338,N_16573,N_16513);
and U21339 (N_21339,N_18373,N_15415);
nand U21340 (N_21340,N_15946,N_19320);
xor U21341 (N_21341,N_18115,N_16165);
xor U21342 (N_21342,N_16136,N_16499);
nand U21343 (N_21343,N_18157,N_18842);
xor U21344 (N_21344,N_15394,N_15714);
or U21345 (N_21345,N_18021,N_15918);
or U21346 (N_21346,N_17181,N_16322);
nor U21347 (N_21347,N_18481,N_16480);
or U21348 (N_21348,N_18001,N_17177);
nand U21349 (N_21349,N_17440,N_19026);
nor U21350 (N_21350,N_17155,N_16438);
and U21351 (N_21351,N_17272,N_15233);
or U21352 (N_21352,N_16947,N_17893);
or U21353 (N_21353,N_19445,N_19936);
nand U21354 (N_21354,N_19556,N_19772);
and U21355 (N_21355,N_18435,N_17678);
nor U21356 (N_21356,N_15475,N_15219);
xnor U21357 (N_21357,N_19429,N_18880);
nand U21358 (N_21358,N_18285,N_16779);
nand U21359 (N_21359,N_15592,N_15998);
and U21360 (N_21360,N_15501,N_15341);
xnor U21361 (N_21361,N_18522,N_15602);
nor U21362 (N_21362,N_17902,N_19273);
and U21363 (N_21363,N_18721,N_18830);
nor U21364 (N_21364,N_16024,N_15747);
or U21365 (N_21365,N_18223,N_16027);
xor U21366 (N_21366,N_17534,N_18448);
nand U21367 (N_21367,N_16288,N_19589);
or U21368 (N_21368,N_19174,N_18210);
xnor U21369 (N_21369,N_16419,N_19323);
and U21370 (N_21370,N_19871,N_17826);
or U21371 (N_21371,N_18189,N_16387);
nor U21372 (N_21372,N_17794,N_17198);
nor U21373 (N_21373,N_15025,N_17777);
nand U21374 (N_21374,N_19864,N_17769);
and U21375 (N_21375,N_18591,N_19315);
nand U21376 (N_21376,N_15745,N_18257);
nor U21377 (N_21377,N_16961,N_16015);
xnor U21378 (N_21378,N_15400,N_15687);
or U21379 (N_21379,N_17008,N_17030);
xnor U21380 (N_21380,N_16848,N_16056);
xnor U21381 (N_21381,N_18504,N_17512);
or U21382 (N_21382,N_16951,N_15414);
nand U21383 (N_21383,N_16771,N_15386);
and U21384 (N_21384,N_15762,N_16832);
or U21385 (N_21385,N_16375,N_16934);
xnor U21386 (N_21386,N_16638,N_16824);
nand U21387 (N_21387,N_15715,N_19570);
nand U21388 (N_21388,N_15832,N_19890);
nor U21389 (N_21389,N_18813,N_16323);
nor U21390 (N_21390,N_19483,N_19821);
and U21391 (N_21391,N_17065,N_17354);
or U21392 (N_21392,N_18000,N_17929);
and U21393 (N_21393,N_18864,N_19835);
nand U21394 (N_21394,N_16348,N_18748);
nor U21395 (N_21395,N_15304,N_17006);
or U21396 (N_21396,N_19279,N_17397);
xnor U21397 (N_21397,N_19018,N_19874);
and U21398 (N_21398,N_17254,N_19623);
nand U21399 (N_21399,N_15094,N_19909);
xor U21400 (N_21400,N_17904,N_17542);
nor U21401 (N_21401,N_15815,N_18375);
xnor U21402 (N_21402,N_16544,N_18107);
and U21403 (N_21403,N_19847,N_19723);
xor U21404 (N_21404,N_17979,N_15591);
nor U21405 (N_21405,N_16632,N_19990);
nor U21406 (N_21406,N_16560,N_19513);
nand U21407 (N_21407,N_19228,N_19287);
and U21408 (N_21408,N_18194,N_16803);
and U21409 (N_21409,N_15647,N_17053);
or U21410 (N_21410,N_16501,N_16650);
nand U21411 (N_21411,N_19260,N_17865);
or U21412 (N_21412,N_19475,N_19172);
or U21413 (N_21413,N_19103,N_17275);
xor U21414 (N_21414,N_18345,N_18272);
or U21415 (N_21415,N_16526,N_15843);
and U21416 (N_21416,N_16634,N_15093);
or U21417 (N_21417,N_18162,N_16658);
nor U21418 (N_21418,N_18969,N_18398);
nand U21419 (N_21419,N_19668,N_16814);
nor U21420 (N_21420,N_15504,N_16101);
nor U21421 (N_21421,N_15390,N_18232);
or U21422 (N_21422,N_16613,N_17662);
xnor U21423 (N_21423,N_19964,N_15293);
or U21424 (N_21424,N_19177,N_18399);
and U21425 (N_21425,N_18315,N_17588);
nor U21426 (N_21426,N_16053,N_17706);
and U21427 (N_21427,N_16719,N_17085);
or U21428 (N_21428,N_16115,N_17709);
or U21429 (N_21429,N_18568,N_15334);
nand U21430 (N_21430,N_17471,N_16030);
or U21431 (N_21431,N_18248,N_16680);
and U21432 (N_21432,N_19735,N_16786);
and U21433 (N_21433,N_18121,N_15768);
xnor U21434 (N_21434,N_15551,N_18197);
or U21435 (N_21435,N_17318,N_16000);
nor U21436 (N_21436,N_16237,N_17661);
nand U21437 (N_21437,N_15092,N_17862);
nand U21438 (N_21438,N_16481,N_15035);
and U21439 (N_21439,N_19935,N_18338);
nand U21440 (N_21440,N_16907,N_19511);
and U21441 (N_21441,N_19224,N_15586);
nor U21442 (N_21442,N_18740,N_16754);
nand U21443 (N_21443,N_18018,N_16317);
nor U21444 (N_21444,N_16469,N_18276);
xnor U21445 (N_21445,N_16488,N_16998);
nor U21446 (N_21446,N_15120,N_19597);
xor U21447 (N_21447,N_16752,N_16320);
and U21448 (N_21448,N_19039,N_17315);
or U21449 (N_21449,N_17300,N_17861);
nor U21450 (N_21450,N_15528,N_19807);
nand U21451 (N_21451,N_18529,N_16945);
xnor U21452 (N_21452,N_15480,N_15549);
or U21453 (N_21453,N_19158,N_18909);
and U21454 (N_21454,N_17339,N_16805);
nor U21455 (N_21455,N_15185,N_16703);
or U21456 (N_21456,N_15083,N_19391);
and U21457 (N_21457,N_16392,N_15645);
nor U21458 (N_21458,N_17649,N_15837);
nor U21459 (N_21459,N_17835,N_15834);
nand U21460 (N_21460,N_17014,N_17202);
or U21461 (N_21461,N_15884,N_15318);
nor U21462 (N_21462,N_17687,N_17621);
xnor U21463 (N_21463,N_18838,N_16932);
nand U21464 (N_21464,N_16919,N_18251);
xnor U21465 (N_21465,N_16533,N_19607);
nor U21466 (N_21466,N_16383,N_19590);
nor U21467 (N_21467,N_19729,N_19708);
and U21468 (N_21468,N_19010,N_18436);
xnor U21469 (N_21469,N_18823,N_18445);
nor U21470 (N_21470,N_15006,N_15014);
nand U21471 (N_21471,N_16798,N_16133);
nand U21472 (N_21472,N_19385,N_15865);
xnor U21473 (N_21473,N_17431,N_17168);
or U21474 (N_21474,N_15886,N_16568);
and U21475 (N_21475,N_15677,N_16400);
or U21476 (N_21476,N_15598,N_17970);
nand U21477 (N_21477,N_16926,N_18562);
nor U21478 (N_21478,N_15142,N_15291);
nor U21479 (N_21479,N_15922,N_18429);
nand U21480 (N_21480,N_19267,N_15996);
nand U21481 (N_21481,N_18379,N_19490);
and U21482 (N_21482,N_17249,N_15982);
nand U21483 (N_21483,N_15652,N_18558);
xnor U21484 (N_21484,N_16331,N_18764);
or U21485 (N_21485,N_18114,N_15197);
nor U21486 (N_21486,N_18193,N_16640);
or U21487 (N_21487,N_19216,N_19785);
nand U21488 (N_21488,N_16649,N_19572);
xnor U21489 (N_21489,N_17036,N_15117);
or U21490 (N_21490,N_18360,N_19066);
nand U21491 (N_21491,N_18583,N_19569);
and U21492 (N_21492,N_18730,N_17759);
nand U21493 (N_21493,N_16420,N_15159);
nand U21494 (N_21494,N_16236,N_15795);
xor U21495 (N_21495,N_17523,N_15670);
or U21496 (N_21496,N_16411,N_19133);
and U21497 (N_21497,N_19388,N_18357);
nand U21498 (N_21498,N_18953,N_17070);
nor U21499 (N_21499,N_15612,N_17146);
xor U21500 (N_21500,N_15324,N_19794);
or U21501 (N_21501,N_18122,N_16437);
nand U21502 (N_21502,N_18638,N_15790);
xnor U21503 (N_21503,N_19154,N_19633);
nand U21504 (N_21504,N_17229,N_16104);
nor U21505 (N_21505,N_17596,N_17567);
nand U21506 (N_21506,N_17450,N_16571);
xor U21507 (N_21507,N_17579,N_17166);
and U21508 (N_21508,N_16646,N_16029);
nand U21509 (N_21509,N_19550,N_17930);
and U21510 (N_21510,N_16725,N_15755);
xor U21511 (N_21511,N_17993,N_17990);
nand U21512 (N_21512,N_17136,N_15075);
nand U21513 (N_21513,N_16091,N_19294);
xor U21514 (N_21514,N_16643,N_18103);
or U21515 (N_21515,N_17047,N_19626);
or U21516 (N_21516,N_16353,N_18152);
xor U21517 (N_21517,N_15473,N_16688);
nor U21518 (N_21518,N_18704,N_19238);
xor U21519 (N_21519,N_19674,N_16290);
or U21520 (N_21520,N_19682,N_18084);
or U21521 (N_21521,N_18105,N_19259);
nand U21522 (N_21522,N_17141,N_16435);
xor U21523 (N_21523,N_19414,N_15833);
or U21524 (N_21524,N_17560,N_19112);
nand U21525 (N_21525,N_18776,N_15078);
nor U21526 (N_21526,N_16660,N_17571);
nor U21527 (N_21527,N_15956,N_18013);
xor U21528 (N_21528,N_16120,N_18293);
nand U21529 (N_21529,N_15633,N_19424);
nand U21530 (N_21530,N_15835,N_15793);
xnor U21531 (N_21531,N_16258,N_16282);
nor U21532 (N_21532,N_17380,N_18145);
xor U21533 (N_21533,N_15438,N_19773);
nor U21534 (N_21534,N_17715,N_19308);
nor U21535 (N_21535,N_17264,N_18016);
xor U21536 (N_21536,N_16904,N_17348);
or U21537 (N_21537,N_19539,N_17143);
or U21538 (N_21538,N_16201,N_15933);
nand U21539 (N_21539,N_19726,N_17367);
or U21540 (N_21540,N_19161,N_17123);
nand U21541 (N_21541,N_16112,N_15430);
xor U21542 (N_21542,N_15022,N_16990);
or U21543 (N_21543,N_19269,N_16561);
nand U21544 (N_21544,N_18863,N_16885);
or U21545 (N_21545,N_15596,N_16622);
or U21546 (N_21546,N_19837,N_15455);
xor U21547 (N_21547,N_15421,N_18432);
or U21548 (N_21548,N_19014,N_15095);
and U21549 (N_21549,N_17049,N_17037);
and U21550 (N_21550,N_19276,N_18926);
and U21551 (N_21551,N_19219,N_16697);
or U21552 (N_21552,N_18096,N_19358);
or U21553 (N_21553,N_18553,N_19503);
nand U21554 (N_21554,N_15002,N_19122);
xor U21555 (N_21555,N_17442,N_19925);
nand U21556 (N_21556,N_19022,N_17010);
xor U21557 (N_21557,N_16424,N_15335);
xnor U21558 (N_21558,N_15408,N_17513);
or U21559 (N_21559,N_16741,N_16833);
nand U21560 (N_21560,N_16929,N_15039);
nand U21561 (N_21561,N_19283,N_19462);
nand U21562 (N_21562,N_17467,N_17227);
nor U21563 (N_21563,N_15288,N_17938);
and U21564 (N_21564,N_18530,N_18545);
nor U21565 (N_21565,N_16181,N_17557);
nand U21566 (N_21566,N_17269,N_15081);
or U21567 (N_21567,N_19064,N_19854);
nand U21568 (N_21568,N_16335,N_17476);
xnor U21569 (N_21569,N_15684,N_16579);
and U21570 (N_21570,N_17150,N_16958);
xnor U21571 (N_21571,N_18490,N_17798);
nor U21572 (N_21572,N_18879,N_15975);
or U21573 (N_21573,N_19997,N_17119);
nand U21574 (N_21574,N_15792,N_16995);
or U21575 (N_21575,N_19609,N_17908);
xor U21576 (N_21576,N_18702,N_17024);
or U21577 (N_21577,N_15977,N_19456);
xnor U21578 (N_21578,N_15960,N_19767);
nand U21579 (N_21579,N_16708,N_15988);
and U21580 (N_21580,N_18127,N_18660);
and U21581 (N_21581,N_16265,N_16546);
xor U21582 (N_21582,N_15599,N_17664);
nand U21583 (N_21583,N_17359,N_19089);
xnor U21584 (N_21584,N_19714,N_18968);
nand U21585 (N_21585,N_18828,N_17501);
and U21586 (N_21586,N_15237,N_17500);
nor U21587 (N_21587,N_19071,N_19567);
nor U21588 (N_21588,N_18540,N_18992);
and U21589 (N_21589,N_17076,N_18612);
or U21590 (N_21590,N_15696,N_19278);
xnor U21591 (N_21591,N_16908,N_15373);
and U21592 (N_21592,N_19080,N_17312);
or U21593 (N_21593,N_17935,N_18178);
nor U21594 (N_21594,N_19088,N_19976);
xor U21595 (N_21595,N_19240,N_16616);
or U21596 (N_21596,N_15830,N_15945);
nand U21597 (N_21597,N_16272,N_15594);
nand U21598 (N_21598,N_16256,N_19948);
nor U21599 (N_21599,N_15099,N_15191);
xor U21600 (N_21600,N_16105,N_16025);
xor U21601 (N_21601,N_19521,N_16472);
and U21602 (N_21602,N_17107,N_15879);
xor U21603 (N_21603,N_15720,N_16737);
and U21604 (N_21604,N_16240,N_18192);
or U21605 (N_21605,N_19622,N_17357);
nor U21606 (N_21606,N_19529,N_17273);
nand U21607 (N_21607,N_17819,N_19307);
or U21608 (N_21608,N_17854,N_19242);
nor U21609 (N_21609,N_17948,N_17607);
or U21610 (N_21610,N_16233,N_16239);
nor U21611 (N_21611,N_15625,N_15272);
and U21612 (N_21612,N_19770,N_16711);
nor U21613 (N_21613,N_19774,N_16764);
xnor U21614 (N_21614,N_15108,N_19143);
nor U21615 (N_21615,N_16993,N_15096);
and U21616 (N_21616,N_19364,N_16852);
or U21617 (N_21617,N_15846,N_17175);
nand U21618 (N_21618,N_16589,N_17463);
or U21619 (N_21619,N_16593,N_17210);
or U21620 (N_21620,N_17732,N_18538);
or U21621 (N_21621,N_16685,N_17788);
nor U21622 (N_21622,N_17892,N_17922);
nor U21623 (N_21623,N_18640,N_16830);
or U21624 (N_21624,N_19400,N_15072);
xor U21625 (N_21625,N_17863,N_16423);
nand U21626 (N_21626,N_19317,N_16930);
xnor U21627 (N_21627,N_19604,N_19918);
nor U21628 (N_21628,N_19447,N_15844);
and U21629 (N_21629,N_16095,N_17235);
xnor U21630 (N_21630,N_17595,N_17128);
nand U21631 (N_21631,N_16683,N_16224);
or U21632 (N_21632,N_17228,N_19059);
xor U21633 (N_21633,N_16340,N_16271);
or U21634 (N_21634,N_18866,N_19848);
nor U21635 (N_21635,N_17699,N_16462);
nor U21636 (N_21636,N_17290,N_19782);
nand U21637 (N_21637,N_19595,N_19555);
xor U21638 (N_21638,N_17064,N_15051);
nor U21639 (N_21639,N_17191,N_19098);
nor U21640 (N_21640,N_18946,N_19032);
xor U21641 (N_21641,N_17341,N_19463);
or U21642 (N_21642,N_19999,N_17443);
or U21643 (N_21643,N_19114,N_18159);
nand U21644 (N_21644,N_15569,N_18499);
and U21645 (N_21645,N_19501,N_19023);
xor U21646 (N_21646,N_17223,N_19482);
nand U21647 (N_21647,N_17148,N_17700);
or U21648 (N_21648,N_16851,N_19165);
nor U21649 (N_21649,N_15689,N_15030);
nand U21650 (N_21650,N_19121,N_16860);
nor U21651 (N_21651,N_17901,N_19886);
and U21652 (N_21652,N_16463,N_15782);
or U21653 (N_21653,N_18295,N_18728);
nor U21654 (N_21654,N_17766,N_15317);
or U21655 (N_21655,N_15358,N_17373);
and U21656 (N_21656,N_15797,N_19850);
nand U21657 (N_21657,N_16135,N_16518);
and U21658 (N_21658,N_18356,N_18075);
nor U21659 (N_21659,N_16690,N_17244);
xor U21660 (N_21660,N_17544,N_17173);
xnor U21661 (N_21661,N_18324,N_16235);
and U21662 (N_21662,N_18335,N_16456);
and U21663 (N_21663,N_18323,N_18492);
and U21664 (N_21664,N_17093,N_15510);
or U21665 (N_21665,N_16625,N_17963);
xor U21666 (N_21666,N_19401,N_16897);
nand U21667 (N_21667,N_17184,N_15472);
or U21668 (N_21668,N_16554,N_17524);
nor U21669 (N_21669,N_18160,N_18717);
and U21670 (N_21670,N_18881,N_16921);
or U21671 (N_21671,N_16777,N_15020);
nand U21672 (N_21672,N_15274,N_16694);
and U21673 (N_21673,N_15144,N_16876);
nor U21674 (N_21674,N_18405,N_19930);
or U21675 (N_21675,N_18279,N_15812);
and U21676 (N_21676,N_15270,N_17707);
nand U21677 (N_21677,N_16005,N_18787);
and U21678 (N_21678,N_17320,N_16681);
or U21679 (N_21679,N_17159,N_15023);
nor U21680 (N_21680,N_15742,N_19966);
nand U21681 (N_21681,N_19900,N_15286);
xor U21682 (N_21682,N_18602,N_16210);
nor U21683 (N_21683,N_17151,N_19344);
xnor U21684 (N_21684,N_16525,N_16743);
xor U21685 (N_21685,N_16713,N_18128);
nor U21686 (N_21686,N_16875,N_19225);
xnor U21687 (N_21687,N_15488,N_18818);
nand U21688 (N_21688,N_15903,N_15440);
nor U21689 (N_21689,N_15963,N_17321);
nand U21690 (N_21690,N_15978,N_17515);
nand U21691 (N_21691,N_18048,N_18779);
nor U21692 (N_21692,N_15231,N_18463);
nor U21693 (N_21693,N_15885,N_16653);
nand U21694 (N_21694,N_19403,N_18355);
and U21695 (N_21695,N_17799,N_17881);
xor U21696 (N_21696,N_17370,N_16620);
nand U21697 (N_21697,N_19235,N_18814);
xor U21698 (N_21698,N_15469,N_18532);
xor U21699 (N_21699,N_16531,N_16449);
xnor U21700 (N_21700,N_16471,N_15576);
and U21701 (N_21701,N_16404,N_18919);
nand U21702 (N_21702,N_17401,N_15361);
or U21703 (N_21703,N_19434,N_18218);
xnor U21704 (N_21704,N_15187,N_17257);
and U21705 (N_21705,N_17187,N_16845);
nand U21706 (N_21706,N_18392,N_17381);
or U21707 (N_21707,N_17998,N_18354);
nand U21708 (N_21708,N_18608,N_15037);
and U21709 (N_21709,N_17832,N_17034);
nor U21710 (N_21710,N_18079,N_15082);
nor U21711 (N_21711,N_16007,N_19168);
or U21712 (N_21712,N_16328,N_18261);
or U21713 (N_21713,N_19784,N_18662);
xor U21714 (N_21714,N_15778,N_19954);
nand U21715 (N_21715,N_19265,N_18200);
and U21716 (N_21716,N_19072,N_19431);
and U21717 (N_21717,N_15388,N_16825);
nand U21718 (N_21718,N_15818,N_19983);
or U21719 (N_21719,N_15381,N_17149);
and U21720 (N_21720,N_19731,N_18883);
nor U21721 (N_21721,N_19050,N_15560);
nor U21722 (N_21722,N_18220,N_15613);
nand U21723 (N_21723,N_18471,N_18856);
xnor U21724 (N_21724,N_15028,N_18126);
xor U21725 (N_21725,N_19115,N_19685);
nand U21726 (N_21726,N_16975,N_16187);
nand U21727 (N_21727,N_16506,N_17303);
xnor U21728 (N_21728,N_18469,N_16881);
nor U21729 (N_21729,N_17393,N_17558);
xor U21730 (N_21730,N_15526,N_19913);
or U21731 (N_21731,N_18670,N_19781);
nor U21732 (N_21732,N_19703,N_17614);
nand U21733 (N_21733,N_18506,N_19411);
and U21734 (N_21734,N_16006,N_18147);
nand U21735 (N_21735,N_19706,N_15695);
nor U21736 (N_21736,N_15140,N_18185);
and U21737 (N_21737,N_15597,N_18376);
nor U21738 (N_21738,N_16739,N_16846);
xor U21739 (N_21739,N_18430,N_19880);
xor U21740 (N_21740,N_15479,N_15784);
nand U21741 (N_21741,N_16989,N_17311);
and U21742 (N_21742,N_17261,N_17455);
and U21743 (N_21743,N_15289,N_15525);
and U21744 (N_21744,N_16037,N_18012);
nand U21745 (N_21745,N_15100,N_18416);
or U21746 (N_21746,N_18703,N_15154);
nor U21747 (N_21747,N_16219,N_18202);
nor U21748 (N_21748,N_16915,N_15489);
xor U21749 (N_21749,N_17002,N_17822);
nor U21750 (N_21750,N_16610,N_19713);
or U21751 (N_21751,N_17305,N_18212);
and U21752 (N_21752,N_16826,N_19485);
and U21753 (N_21753,N_17633,N_16234);
nor U21754 (N_21754,N_17172,N_17362);
or U21755 (N_21755,N_16202,N_18406);
xnor U21756 (N_21756,N_19939,N_16734);
xnor U21757 (N_21757,N_15396,N_19257);
or U21758 (N_21758,N_18459,N_18678);
xor U21759 (N_21759,N_17577,N_16305);
nor U21760 (N_21760,N_16861,N_17297);
and U21761 (N_21761,N_17497,N_16410);
xor U21762 (N_21762,N_17967,N_17521);
or U21763 (N_21763,N_18136,N_15794);
and U21764 (N_21764,N_17897,N_19377);
nand U21765 (N_21765,N_18597,N_15985);
or U21766 (N_21766,N_15620,N_19141);
nand U21767 (N_21767,N_18466,N_19484);
and U21768 (N_21768,N_15894,N_16512);
nand U21769 (N_21769,N_18346,N_19361);
nor U21770 (N_21770,N_19955,N_16746);
or U21771 (N_21771,N_19778,N_17549);
nor U21772 (N_21772,N_18887,N_18859);
xor U21773 (N_21773,N_15184,N_18888);
and U21774 (N_21774,N_19081,N_16957);
or U21775 (N_21775,N_17234,N_18705);
nor U21776 (N_21776,N_17581,N_18040);
and U21777 (N_21777,N_18790,N_17444);
nor U21778 (N_21778,N_18297,N_19843);
nor U21779 (N_21779,N_18119,N_19398);
nor U21780 (N_21780,N_16866,N_16570);
or U21781 (N_21781,N_19153,N_16102);
nand U21782 (N_21782,N_17292,N_17333);
or U21783 (N_21783,N_15119,N_16489);
nand U21784 (N_21784,N_17059,N_15046);
and U21785 (N_21785,N_16178,N_16077);
xnor U21786 (N_21786,N_19494,N_17651);
or U21787 (N_21787,N_17504,N_17383);
nand U21788 (N_21788,N_15066,N_15285);
nor U21789 (N_21789,N_17741,N_15417);
and U21790 (N_21790,N_19849,N_16603);
nand U21791 (N_21791,N_15412,N_16464);
xor U21792 (N_21792,N_17917,N_19421);
nand U21793 (N_21793,N_18426,N_17061);
and U21794 (N_21794,N_15555,N_18351);
xnor U21795 (N_21795,N_16985,N_15550);
nand U21796 (N_21796,N_16535,N_18639);
xor U21797 (N_21797,N_19004,N_15166);
or U21798 (N_21798,N_16959,N_18250);
xnor U21799 (N_21799,N_15590,N_16168);
nor U21800 (N_21800,N_15232,N_16263);
xor U21801 (N_21801,N_18143,N_19300);
or U21802 (N_21802,N_17971,N_16768);
and U21803 (N_21803,N_19437,N_18884);
or U21804 (N_21804,N_19702,N_18314);
nor U21805 (N_21805,N_16369,N_19386);
xnor U21806 (N_21806,N_17797,N_19875);
xor U21807 (N_21807,N_18843,N_15656);
xnor U21808 (N_21808,N_15384,N_17559);
or U21809 (N_21809,N_15961,N_16330);
or U21810 (N_21810,N_18294,N_16617);
xor U21811 (N_21811,N_16394,N_17050);
and U21812 (N_21812,N_17319,N_17647);
and U21813 (N_21813,N_16399,N_19911);
or U21814 (N_21814,N_15823,N_19637);
nand U21815 (N_21815,N_16607,N_17480);
nor U21816 (N_21816,N_17674,N_18167);
or U21817 (N_21817,N_18292,N_19926);
xnor U21818 (N_21818,N_19817,N_19343);
nand U21819 (N_21819,N_19605,N_19910);
xnor U21820 (N_21820,N_15426,N_17942);
xor U21821 (N_21821,N_16682,N_17787);
nor U21822 (N_21822,N_19438,N_16843);
nor U21823 (N_21823,N_16644,N_17844);
nand U21824 (N_21824,N_15623,N_16721);
nor U21825 (N_21825,N_17410,N_16457);
nor U21826 (N_21826,N_19762,N_19399);
xor U21827 (N_21827,N_19327,N_19927);
xor U21828 (N_21828,N_16898,N_15033);
and U21829 (N_21829,N_16936,N_19737);
xnor U21830 (N_21830,N_15764,N_16064);
and U21831 (N_21831,N_17923,N_17964);
or U21832 (N_21832,N_18564,N_17878);
nor U21833 (N_21833,N_18550,N_17256);
and U21834 (N_21834,N_18687,N_18649);
xor U21835 (N_21835,N_19688,N_19415);
nand U21836 (N_21836,N_18694,N_16096);
nand U21837 (N_21837,N_19202,N_17351);
or U21838 (N_21838,N_15132,N_18423);
and U21839 (N_21839,N_18011,N_18870);
nor U21840 (N_21840,N_17665,N_19614);
xor U21841 (N_21841,N_17090,N_16856);
and U21842 (N_21842,N_19671,N_16441);
nand U21843 (N_21843,N_17167,N_15061);
and U21844 (N_21844,N_16365,N_15580);
and U21845 (N_21845,N_19461,N_18965);
or U21846 (N_21846,N_18744,N_19200);
nand U21847 (N_21847,N_17248,N_16326);
and U21848 (N_21848,N_16099,N_18502);
nand U21849 (N_21849,N_18050,N_16111);
nor U21850 (N_21850,N_16973,N_18815);
and U21851 (N_21851,N_19409,N_19366);
nor U21852 (N_21852,N_15931,N_16676);
nand U21853 (N_21853,N_17898,N_16659);
xnor U21854 (N_21854,N_19543,N_16418);
nor U21855 (N_21855,N_18453,N_15380);
nor U21856 (N_21856,N_16972,N_18785);
nand U21857 (N_21857,N_19645,N_15205);
or U21858 (N_21858,N_16971,N_16905);
nand U21859 (N_21859,N_18943,N_15121);
nor U21860 (N_21860,N_19470,N_19378);
nand U21861 (N_21861,N_17392,N_15367);
xor U21862 (N_21862,N_17669,N_16732);
or U21863 (N_21863,N_17094,N_17377);
nor U21864 (N_21864,N_16378,N_15893);
nor U21865 (N_21865,N_17555,N_18895);
nand U21866 (N_21866,N_16819,N_19630);
nor U21867 (N_21867,N_17213,N_18402);
xor U21868 (N_21868,N_19786,N_15871);
nand U21869 (N_21869,N_19159,N_16148);
xnor U21870 (N_21870,N_15629,N_16065);
nor U21871 (N_21871,N_17635,N_18186);
and U21872 (N_21872,N_18247,N_17092);
and U21873 (N_21873,N_15955,N_16380);
nor U21874 (N_21874,N_18465,N_17221);
nor U21875 (N_21875,N_17667,N_16781);
nand U21876 (N_21876,N_19816,N_18571);
and U21877 (N_21877,N_17505,N_18998);
nor U21878 (N_21878,N_17265,N_19087);
or U21879 (N_21879,N_16377,N_15535);
and U21880 (N_21880,N_19352,N_19247);
nand U21881 (N_21881,N_18542,N_19094);
nor U21882 (N_21882,N_15199,N_16139);
or U21883 (N_21883,N_17079,N_17601);
or U21884 (N_21884,N_17629,N_15587);
nand U21885 (N_21885,N_15201,N_17800);
nand U21886 (N_21886,N_18106,N_18266);
nor U21887 (N_21887,N_18773,N_19863);
and U21888 (N_21888,N_17028,N_16019);
xor U21889 (N_21889,N_15672,N_18615);
nand U21890 (N_21890,N_17451,N_19179);
nor U21891 (N_21891,N_19775,N_15212);
nor U21892 (N_21892,N_18118,N_18056);
nand U21893 (N_21893,N_17744,N_17939);
xnor U21894 (N_21894,N_16473,N_16925);
or U21895 (N_21895,N_17447,N_17514);
or U21896 (N_21896,N_15779,N_18587);
xnor U21897 (N_21897,N_16521,N_15364);
or U21898 (N_21898,N_16773,N_17675);
or U21899 (N_21899,N_18709,N_18184);
xnor U21900 (N_21900,N_15102,N_18912);
xor U21901 (N_21901,N_18674,N_17739);
nor U21902 (N_21902,N_17250,N_15182);
xnor U21903 (N_21903,N_17603,N_19542);
and U21904 (N_21904,N_17784,N_17876);
nand U21905 (N_21905,N_18574,N_16122);
nor U21906 (N_21906,N_15427,N_19105);
nor U21907 (N_21907,N_19895,N_19371);
xnor U21908 (N_21908,N_17937,N_17083);
or U21909 (N_21909,N_18929,N_15741);
xor U21910 (N_21910,N_17086,N_16700);
nand U21911 (N_21911,N_16193,N_15514);
or U21912 (N_21912,N_15729,N_17676);
and U21913 (N_21913,N_17291,N_16627);
xor U21914 (N_21914,N_19261,N_16358);
nand U21915 (N_21915,N_15379,N_15477);
nor U21916 (N_21916,N_18243,N_18593);
xnor U21917 (N_21917,N_16382,N_19515);
xor U21918 (N_21918,N_18227,N_16191);
nand U21919 (N_21919,N_17519,N_18281);
nand U21920 (N_21920,N_19603,N_15044);
xnor U21921 (N_21921,N_18446,N_17435);
or U21922 (N_21922,N_16751,N_18624);
nand U21923 (N_21923,N_16831,N_17710);
nor U21924 (N_21924,N_18620,N_19092);
xnor U21925 (N_21925,N_15531,N_15537);
nand U21926 (N_21926,N_15615,N_16844);
nand U21927 (N_21927,N_18081,N_17828);
or U21928 (N_21928,N_18594,N_17574);
and U21929 (N_21929,N_16028,N_15901);
nor U21930 (N_21930,N_15907,N_19033);
and U21931 (N_21931,N_15813,N_16183);
or U21932 (N_21932,N_18071,N_16376);
nand U21933 (N_21933,N_15021,N_18971);
nand U21934 (N_21934,N_16789,N_17873);
nand U21935 (N_21935,N_18496,N_19298);
nand U21936 (N_21936,N_18833,N_15650);
nor U21937 (N_21937,N_16588,N_19077);
nand U21938 (N_21938,N_15974,N_15563);
xnor U21939 (N_21939,N_16818,N_15512);
and U21940 (N_21940,N_18231,N_19430);
or U21941 (N_21941,N_19855,N_15149);
nor U21942 (N_21942,N_17753,N_17679);
and U21943 (N_21943,N_15320,N_18289);
nand U21944 (N_21944,N_18226,N_16155);
and U21945 (N_21945,N_18928,N_16744);
or U21946 (N_21946,N_17885,N_15935);
nor U21947 (N_21947,N_17126,N_16173);
xor U21948 (N_21948,N_17728,N_16910);
nor U21949 (N_21949,N_17888,N_16736);
or U21950 (N_21950,N_16426,N_19251);
or U21951 (N_21951,N_17859,N_18172);
or U21952 (N_21952,N_17774,N_15806);
or U21953 (N_21953,N_15651,N_15256);
and U21954 (N_21954,N_17003,N_18941);
and U21955 (N_21955,N_16049,N_19355);
nor U21956 (N_21956,N_16106,N_15511);
xor U21957 (N_21957,N_16194,N_17600);
and U21958 (N_21958,N_18741,N_19858);
or U21959 (N_21959,N_15301,N_18161);
nand U21960 (N_21960,N_18438,N_18310);
nor U21961 (N_21961,N_19588,N_18973);
nor U21962 (N_21962,N_15215,N_18473);
xnor U21963 (N_21963,N_16090,N_19286);
and U21964 (N_21964,N_16137,N_17176);
xnor U21965 (N_21965,N_18989,N_16302);
and U21966 (N_21966,N_18720,N_16655);
nor U21967 (N_21967,N_17101,N_17803);
or U21968 (N_21968,N_17729,N_17025);
and U21969 (N_21969,N_16964,N_19764);
nor U21970 (N_21970,N_17196,N_19229);
nor U21971 (N_21971,N_17441,N_15619);
or U21972 (N_21972,N_17983,N_15861);
xor U21973 (N_21973,N_15113,N_19192);
xor U21974 (N_21974,N_17655,N_15161);
and U21975 (N_21975,N_15277,N_18129);
nor U21976 (N_21976,N_18427,N_19934);
nor U21977 (N_21977,N_15242,N_15363);
or U21978 (N_21978,N_18411,N_17845);
nor U21979 (N_21979,N_18080,N_17773);
nor U21980 (N_21980,N_15756,N_15816);
xor U21981 (N_21981,N_18235,N_16396);
and U21982 (N_21982,N_19989,N_19819);
and U21983 (N_21983,N_15624,N_16967);
nand U21984 (N_21984,N_18655,N_16275);
nor U21985 (N_21985,N_19631,N_16619);
and U21986 (N_21986,N_18786,N_18664);
nor U21987 (N_21987,N_16809,N_16509);
nor U21988 (N_21988,N_16900,N_19070);
or U21989 (N_21989,N_16599,N_15659);
or U21990 (N_21990,N_17484,N_18095);
nand U21991 (N_21991,N_17743,N_16615);
and U21992 (N_21992,N_19075,N_17645);
nand U21993 (N_21993,N_18443,N_19395);
and U21994 (N_21994,N_17120,N_15663);
or U21995 (N_21995,N_17591,N_17302);
nand U21996 (N_21996,N_18548,N_16218);
nand U21997 (N_21997,N_19196,N_18233);
xnor U21998 (N_21998,N_17719,N_15875);
xor U21999 (N_21999,N_15326,N_16157);
nand U22000 (N_22000,N_19441,N_16110);
or U22001 (N_22001,N_18754,N_18803);
nand U22002 (N_22002,N_17842,N_15459);
and U22003 (N_22003,N_15914,N_16354);
xnor U22004 (N_22004,N_19310,N_19952);
and U22005 (N_22005,N_18477,N_17220);
nor U22006 (N_22006,N_15017,N_15657);
xor U22007 (N_22007,N_17553,N_17740);
nand U22008 (N_22008,N_16810,N_19985);
or U22009 (N_22009,N_15941,N_17243);
or U22010 (N_22010,N_19883,N_16745);
or U22011 (N_22011,N_18940,N_16109);
or U22012 (N_22012,N_19370,N_17425);
or U22013 (N_22013,N_19053,N_17883);
nor U22014 (N_22014,N_15954,N_18087);
xor U22015 (N_22015,N_15579,N_15047);
xnor U22016 (N_22016,N_17578,N_19012);
nor U22017 (N_22017,N_16153,N_16172);
or U22018 (N_22018,N_15034,N_19834);
nor U22019 (N_22019,N_17408,N_15000);
xnor U22020 (N_22020,N_16962,N_19818);
nor U22021 (N_22021,N_19046,N_19068);
or U22022 (N_22022,N_19357,N_18605);
and U22023 (N_22023,N_15168,N_15485);
xnor U22024 (N_22024,N_16794,N_19635);
nor U22025 (N_22025,N_18726,N_19037);
xor U22026 (N_22026,N_16740,N_15690);
or U22027 (N_22027,N_16164,N_16528);
xnor U22028 (N_22028,N_19921,N_16405);
xnor U22029 (N_22029,N_16894,N_16684);
xnor U22030 (N_22030,N_17283,N_17928);
or U22031 (N_22031,N_16776,N_18590);
xor U22032 (N_22032,N_18455,N_19711);
xnor U22033 (N_22033,N_17806,N_15701);
xor U22034 (N_22034,N_16451,N_17446);
or U22035 (N_22035,N_17316,N_15466);
and U22036 (N_22036,N_17891,N_16514);
xnor U22037 (N_22037,N_18344,N_19363);
or U22038 (N_22038,N_15634,N_18758);
nor U22039 (N_22039,N_19512,N_16350);
nor U22040 (N_22040,N_18536,N_19830);
xnor U22041 (N_22041,N_18517,N_16606);
nand U22042 (N_22042,N_18631,N_18112);
nor U22043 (N_22043,N_18501,N_16847);
and U22044 (N_22044,N_19296,N_19998);
nor U22045 (N_22045,N_19191,N_17630);
nor U22046 (N_22046,N_16475,N_16343);
xnor U22047 (N_22047,N_19243,N_19212);
or U22048 (N_22048,N_19390,N_18252);
and U22049 (N_22049,N_15439,N_15257);
xnor U22050 (N_22050,N_16891,N_18636);
xnor U22051 (N_22051,N_15300,N_17851);
xor U22052 (N_22052,N_17270,N_17724);
and U22053 (N_22053,N_16834,N_17650);
and U22054 (N_22054,N_19962,N_17721);
and U22055 (N_22055,N_19811,N_16707);
and U22056 (N_22056,N_17907,N_18876);
nor U22057 (N_22057,N_15080,N_18451);
xor U22058 (N_22058,N_15553,N_16363);
nor U22059 (N_22059,N_18022,N_19856);
nand U22060 (N_22060,N_16397,N_18439);
and U22061 (N_22061,N_18032,N_19896);
and U22062 (N_22062,N_18603,N_15639);
xor U22063 (N_22063,N_17727,N_18102);
xor U22064 (N_22064,N_16883,N_19245);
and U22065 (N_22065,N_16872,N_18195);
and U22066 (N_22066,N_16131,N_15697);
and U22067 (N_22067,N_16292,N_15928);
nor U22068 (N_22068,N_19823,N_15610);
nand U22069 (N_22069,N_16276,N_15302);
xnor U22070 (N_22070,N_18937,N_16038);
or U22071 (N_22071,N_18565,N_18696);
xor U22072 (N_22072,N_19006,N_19162);
xnor U22073 (N_22073,N_16933,N_19372);
and U22074 (N_22074,N_19142,N_16532);
xnor U22075 (N_22075,N_18627,N_19375);
and U22076 (N_22076,N_15060,N_15608);
xnor U22077 (N_22077,N_15261,N_17466);
nand U22078 (N_22078,N_16720,N_19756);
nand U22079 (N_22079,N_15141,N_17475);
and U22080 (N_22080,N_17616,N_16107);
nand U22081 (N_22081,N_18156,N_16118);
nand U22082 (N_22082,N_15209,N_15637);
nor U22083 (N_22083,N_18074,N_19889);
or U22084 (N_22084,N_17022,N_19719);
and U22085 (N_22085,N_16190,N_17360);
nand U22086 (N_22086,N_15630,N_18994);
and U22087 (N_22087,N_18614,N_15124);
and U22088 (N_22088,N_19689,N_16314);
nor U22089 (N_22089,N_17867,N_15325);
or U22090 (N_22090,N_19250,N_18179);
xor U22091 (N_22091,N_15031,N_17757);
nand U22092 (N_22092,N_19239,N_17323);
xor U22093 (N_22093,N_15556,N_17219);
nand U22094 (N_22094,N_17681,N_17295);
xnor U22095 (N_22095,N_16364,N_18554);
or U22096 (N_22096,N_19118,N_15474);
xor U22097 (N_22097,N_15703,N_16158);
or U22098 (N_22098,N_15203,N_19643);
and U22099 (N_22099,N_17823,N_16600);
xor U22100 (N_22100,N_16167,N_15218);
and U22101 (N_22101,N_19043,N_18264);
and U22102 (N_22102,N_16902,N_17023);
nand U22103 (N_22103,N_19704,N_15281);
or U22104 (N_22104,N_16198,N_16393);
or U22105 (N_22105,N_18028,N_19672);
and U22106 (N_22106,N_18124,N_16486);
or U22107 (N_22107,N_16551,N_18996);
nand U22108 (N_22108,N_16001,N_19853);
and U22109 (N_22109,N_19140,N_17327);
xnor U22110 (N_22110,N_16595,N_17778);
and U22111 (N_22111,N_17821,N_15574);
xor U22112 (N_22112,N_19528,N_18209);
xnor U22113 (N_22113,N_16176,N_18417);
nor U22114 (N_22114,N_19532,N_16221);
nand U22115 (N_22115,N_17986,N_17623);
and U22116 (N_22116,N_18309,N_18358);
xor U22117 (N_22117,N_18524,N_18259);
xnor U22118 (N_22118,N_19124,N_16433);
and U22119 (N_22119,N_18480,N_18434);
or U22120 (N_22120,N_16403,N_18229);
nand U22121 (N_22121,N_15840,N_15734);
nor U22122 (N_22122,N_16284,N_18219);
and U22123 (N_22123,N_17975,N_15433);
and U22124 (N_22124,N_15016,N_15245);
and U22125 (N_22125,N_17801,N_17516);
nor U22126 (N_22126,N_19479,N_15678);
or U22127 (N_22127,N_15283,N_16729);
nor U22128 (N_22128,N_17409,N_16412);
xor U22129 (N_22129,N_18249,N_16020);
nand U22130 (N_22130,N_16483,N_18407);
nand U22131 (N_22131,N_16557,N_15482);
xor U22132 (N_22132,N_19288,N_17405);
and U22133 (N_22133,N_15279,N_17999);
xor U22134 (N_22134,N_15601,N_18718);
nor U22135 (N_22135,N_18806,N_16445);
nand U22136 (N_22136,N_17096,N_18101);
and U22137 (N_22137,N_16012,N_19740);
xnor U22138 (N_22138,N_16230,N_15419);
xnor U22139 (N_22139,N_19432,N_18747);
nand U22140 (N_22140,N_15089,N_19559);
nor U22141 (N_22141,N_15759,N_16251);
or U22142 (N_22142,N_19019,N_18328);
nor U22143 (N_22143,N_17108,N_17663);
xor U22144 (N_22144,N_16670,N_16402);
xor U22145 (N_22145,N_16092,N_15856);
xnor U22146 (N_22146,N_15163,N_16443);
nand U22147 (N_22147,N_15483,N_15909);
xor U22148 (N_22148,N_16954,N_16333);
or U22149 (N_22149,N_19564,N_19897);
nor U22150 (N_22150,N_16838,N_18944);
nand U22151 (N_22151,N_19578,N_18061);
xnor U22152 (N_22152,N_18716,N_18675);
nor U22153 (N_22153,N_15723,N_17328);
or U22154 (N_22154,N_15735,N_16381);
nand U22155 (N_22155,N_15138,N_17541);
or U22156 (N_22156,N_18069,N_16264);
nand U22157 (N_22157,N_15471,N_15465);
nor U22158 (N_22158,N_17860,N_19885);
and U22159 (N_22159,N_17617,N_19938);
and U22160 (N_22160,N_17536,N_18511);
xnor U22161 (N_22161,N_18788,N_15458);
or U22162 (N_22162,N_17839,N_19832);
or U22163 (N_22163,N_17116,N_19206);
xor U22164 (N_22164,N_19608,N_15584);
and U22165 (N_22165,N_17240,N_18810);
nand U22166 (N_22166,N_15362,N_19211);
or U22167 (N_22167,N_15145,N_17004);
or U22168 (N_22168,N_19747,N_17279);
nor U22169 (N_22169,N_16242,N_16730);
nand U22170 (N_22170,N_15929,N_19123);
nand U22171 (N_22171,N_15939,N_19453);
xor U22172 (N_22172,N_16543,N_17969);
xnor U22173 (N_22173,N_18164,N_17996);
xnor U22174 (N_22174,N_19419,N_17827);
and U22175 (N_22175,N_15585,N_16692);
and U22176 (N_22176,N_18015,N_16226);
and U22177 (N_22177,N_17412,N_19809);
and U22178 (N_22178,N_18808,N_18094);
nand U22179 (N_22179,N_18440,N_17448);
nand U22180 (N_22180,N_16497,N_19598);
nand U22181 (N_22181,N_17690,N_19940);
or U22182 (N_22182,N_16862,N_18668);
nand U22183 (N_22183,N_16217,N_16249);
xnor U22184 (N_22184,N_19246,N_18653);
and U22185 (N_22185,N_19226,N_19316);
xnor U22186 (N_22186,N_19991,N_19891);
and U22187 (N_22187,N_15517,N_16138);
and U22188 (N_22188,N_18254,N_15669);
nor U22189 (N_22189,N_16259,N_17376);
and U22190 (N_22190,N_19301,N_18457);
nor U22191 (N_22191,N_17395,N_19906);
xnor U22192 (N_22192,N_16853,N_15496);
and U22193 (N_22193,N_15052,N_19829);
or U22194 (N_22194,N_18552,N_17138);
and U22195 (N_22195,N_16152,N_18834);
xor U22196 (N_22196,N_18148,N_18851);
or U22197 (N_22197,N_19526,N_19787);
xor U22198 (N_22198,N_17057,N_18819);
and U22199 (N_22199,N_19139,N_17704);
xnor U22200 (N_22200,N_19531,N_16635);
or U22201 (N_22201,N_15192,N_19000);
xor U22202 (N_22202,N_15253,N_17080);
nor U22203 (N_22203,N_19924,N_17329);
or U22204 (N_22204,N_16080,N_19944);
xnor U22205 (N_22205,N_19697,N_15905);
xnor U22206 (N_22206,N_16922,N_16587);
nand U22207 (N_22207,N_17697,N_18731);
or U22208 (N_22208,N_19331,N_17506);
or U22209 (N_22209,N_17052,N_16316);
xor U22210 (N_22210,N_16996,N_16775);
or U22211 (N_22211,N_18525,N_18486);
nor U22212 (N_22212,N_16466,N_19981);
xnor U22213 (N_22213,N_15976,N_15263);
or U22214 (N_22214,N_15254,N_15917);
xor U22215 (N_22215,N_18301,N_19384);
and U22216 (N_22216,N_18581,N_18004);
or U22217 (N_22217,N_17117,N_15738);
and U22218 (N_22218,N_17282,N_16756);
xnor U22219 (N_22219,N_15499,N_15135);
or U22220 (N_22220,N_16163,N_16196);
nand U22221 (N_22221,N_15315,N_16408);
and U22222 (N_22222,N_19801,N_16801);
xor U22223 (N_22223,N_17974,N_17936);
or U22224 (N_22224,N_18509,N_16373);
or U22225 (N_22225,N_15437,N_17916);
xor U22226 (N_22226,N_16160,N_15508);
nor U22227 (N_22227,N_18482,N_15583);
nand U22228 (N_22228,N_17346,N_16032);
nor U22229 (N_22229,N_15401,N_19451);
nor U22230 (N_22230,N_18701,N_15012);
and U22231 (N_22231,N_19052,N_16075);
nor U22232 (N_22232,N_19193,N_19866);
and U22233 (N_22233,N_17498,N_19899);
or U22234 (N_22234,N_18566,N_16982);
or U22235 (N_22235,N_15655,N_19234);
xnor U22236 (N_22236,N_16170,N_15538);
and U22237 (N_22237,N_15217,N_15947);
and U22238 (N_22238,N_15088,N_17730);
xnor U22239 (N_22239,N_15225,N_18116);
xor U22240 (N_22240,N_19397,N_15641);
nand U22241 (N_22241,N_15683,N_18966);
xnor U22242 (N_22242,N_19612,N_19125);
nor U22243 (N_22243,N_17889,N_16874);
and U22244 (N_22244,N_19825,N_18698);
xor U22245 (N_22245,N_15822,N_18042);
nand U22246 (N_22246,N_19884,N_16618);
or U22247 (N_22247,N_16790,N_17051);
and U22248 (N_22248,N_16987,N_19859);
nand U22249 (N_22249,N_17499,N_15796);
nand U22250 (N_22250,N_19510,N_19994);
nand U22251 (N_22251,N_18514,N_16714);
nor U22252 (N_22252,N_19766,N_18130);
and U22253 (N_22253,N_19691,N_16669);
and U22254 (N_22254,N_18182,N_16182);
nand U22255 (N_22255,N_18100,N_17786);
xnor U22256 (N_22256,N_15515,N_15632);
xor U22257 (N_22257,N_15470,N_16583);
or U22258 (N_22258,N_16495,N_15870);
xnor U22259 (N_22259,N_17162,N_15973);
xor U22260 (N_22260,N_16515,N_18677);
nand U22261 (N_22261,N_18642,N_15045);
or U22262 (N_22262,N_15561,N_18604);
nor U22263 (N_22263,N_18364,N_17611);
xor U22264 (N_22264,N_15091,N_15450);
or U22265 (N_22265,N_17147,N_18936);
nor U22266 (N_22266,N_19846,N_19574);
nand U22267 (N_22267,N_18995,N_18539);
or U22268 (N_22268,N_19163,N_15991);
and U22269 (N_22269,N_19180,N_15940);
and U22270 (N_22270,N_15382,N_18173);
nor U22271 (N_22271,N_19541,N_18848);
or U22272 (N_22272,N_15502,N_18560);
and U22273 (N_22273,N_16978,N_17791);
xor U22274 (N_22274,N_16767,N_16215);
or U22275 (N_22275,N_18976,N_17882);
or U22276 (N_22276,N_18083,N_19147);
nor U22277 (N_22277,N_17529,N_18923);
nand U22278 (N_22278,N_15589,N_16821);
nor U22279 (N_22279,N_18546,N_17949);
nor U22280 (N_22280,N_17723,N_15395);
xnor U22281 (N_22281,N_18352,N_16345);
xnor U22282 (N_22282,N_17005,N_17836);
and U22283 (N_22283,N_18461,N_17517);
and U22284 (N_22284,N_16920,N_15926);
or U22285 (N_22285,N_18153,N_15769);
and U22286 (N_22286,N_17242,N_15249);
or U22287 (N_22287,N_15673,N_18135);
and U22288 (N_22288,N_17947,N_18168);
or U22289 (N_22289,N_15247,N_18763);
xnor U22290 (N_22290,N_16696,N_17414);
or U22291 (N_22291,N_16003,N_16984);
and U22292 (N_22292,N_19185,N_18573);
and U22293 (N_22293,N_18559,N_16536);
nand U22294 (N_22294,N_18849,N_18349);
or U22295 (N_22295,N_18205,N_18308);
or U22296 (N_22296,N_17135,N_17978);
or U22297 (N_22297,N_19258,N_19134);
and U22298 (N_22298,N_19941,N_19047);
or U22299 (N_22299,N_18263,N_16577);
or U22300 (N_22300,N_17246,N_18610);
or U22301 (N_22301,N_16507,N_16097);
nand U22302 (N_22302,N_17813,N_15862);
xor U22303 (N_22303,N_15743,N_19150);
or U22304 (N_22304,N_18924,N_17568);
xor U22305 (N_22305,N_18280,N_17113);
and U22306 (N_22306,N_16935,N_18885);
and U22307 (N_22307,N_19509,N_16033);
xor U22308 (N_22308,N_15409,N_16310);
nor U22309 (N_22309,N_16057,N_19195);
nand U22310 (N_22310,N_16203,N_19506);
or U22311 (N_22311,N_17465,N_15255);
or U22312 (N_22312,N_17456,N_19568);
or U22313 (N_22313,N_16829,N_18982);
nand U22314 (N_22314,N_16159,N_19750);
and U22315 (N_22315,N_16175,N_16309);
nor U22316 (N_22316,N_17486,N_18007);
xnor U22317 (N_22317,N_17072,N_15273);
or U22318 (N_22318,N_19988,N_19396);
or U22319 (N_22319,N_19662,N_19932);
or U22320 (N_22320,N_19282,N_18216);
nor U22321 (N_22321,N_16048,N_19712);
nand U22322 (N_22322,N_17590,N_15726);
nor U22323 (N_22323,N_16072,N_16044);
xor U22324 (N_22324,N_15867,N_15222);
and U22325 (N_22325,N_18054,N_15198);
or U22326 (N_22326,N_18679,N_15452);
nand U22327 (N_22327,N_17258,N_19797);
nand U22328 (N_22328,N_15435,N_17931);
nor U22329 (N_22329,N_17927,N_17016);
or U22330 (N_22330,N_16970,N_16280);
nand U22331 (N_22331,N_19189,N_17112);
nand U22332 (N_22332,N_17584,N_19873);
nor U22333 (N_22333,N_19045,N_19945);
xnor U22334 (N_22334,N_18903,N_17423);
xor U22335 (N_22335,N_16042,N_17575);
and U22336 (N_22336,N_18082,N_18437);
nand U22337 (N_22337,N_18513,N_18369);
nand U22338 (N_22338,N_17231,N_17780);
and U22339 (N_22339,N_16315,N_18691);
nand U22340 (N_22340,N_18981,N_17238);
nor U22341 (N_22341,N_17042,N_17554);
xor U22342 (N_22342,N_15305,N_15377);
nand U22343 (N_22343,N_19581,N_18618);
nand U22344 (N_22344,N_15863,N_19498);
or U22345 (N_22345,N_16150,N_16087);
or U22346 (N_22346,N_19916,N_17468);
nand U22347 (N_22347,N_15727,N_18825);
or U22348 (N_22348,N_16878,N_16371);
nand U22349 (N_22349,N_18857,N_17073);
and U22350 (N_22350,N_18835,N_17834);
nand U22351 (N_22351,N_16071,N_17084);
xor U22352 (N_22352,N_15243,N_16177);
nand U22353 (N_22353,N_15200,N_18650);
nor U22354 (N_22354,N_16432,N_18521);
or U22355 (N_22355,N_15423,N_18663);
nand U22356 (N_22356,N_15997,N_19237);
nor U22357 (N_22357,N_19530,N_15103);
or U22358 (N_22358,N_16117,N_19109);
and U22359 (N_22359,N_15228,N_15413);
or U22360 (N_22360,N_15801,N_18236);
and U22361 (N_22361,N_19881,N_18999);
nor U22362 (N_22362,N_16727,N_17267);
xor U22363 (N_22363,N_15717,N_17217);
xnor U22364 (N_22364,N_15807,N_17688);
and U22365 (N_22365,N_17183,N_18306);
xnor U22366 (N_22366,N_19270,N_16738);
nand U22367 (N_22367,N_16591,N_17301);
xor U22368 (N_22368,N_19763,N_17526);
nor U22369 (N_22369,N_16749,N_16360);
xor U22370 (N_22370,N_18534,N_19827);
and U22371 (N_22371,N_19210,N_17018);
nand U22372 (N_22372,N_19733,N_19720);
nand U22373 (N_22373,N_16039,N_18002);
nor U22374 (N_22374,N_17570,N_17132);
and U22375 (N_22375,N_18781,N_18759);
nor U22376 (N_22376,N_17114,N_19056);
xnor U22377 (N_22377,N_17274,N_19933);
xor U22378 (N_22378,N_19628,N_15180);
nand U22379 (N_22379,N_15814,N_17180);
and U22380 (N_22380,N_17482,N_17403);
and U22381 (N_22381,N_15711,N_15716);
and U22382 (N_22382,N_18155,N_15904);
and U22383 (N_22383,N_16594,N_17232);
or U22384 (N_22384,N_15346,N_18952);
xnor U22385 (N_22385,N_15158,N_16760);
or U22386 (N_22386,N_15156,N_16835);
or U22387 (N_22387,N_16228,N_17335);
or U22388 (N_22388,N_18494,N_16504);
nand U22389 (N_22389,N_19167,N_17386);
or U22390 (N_22390,N_15169,N_17940);
and U22391 (N_22391,N_19313,N_19284);
xnor U22392 (N_22392,N_15631,N_18166);
nand U22393 (N_22393,N_17472,N_15548);
and U22394 (N_22394,N_16332,N_17278);
xnor U22395 (N_22395,N_16733,N_17378);
or U22396 (N_22396,N_17671,N_15224);
xor U22397 (N_22397,N_16303,N_15800);
and U22398 (N_22398,N_16689,N_15821);
xnor U22399 (N_22399,N_19902,N_15193);
or U22400 (N_22400,N_16192,N_17164);
and U22401 (N_22401,N_15310,N_18131);
or U22402 (N_22402,N_15915,N_16795);
and U22403 (N_22403,N_19079,N_16960);
nand U22404 (N_22404,N_17613,N_17610);
xor U22405 (N_22405,N_16306,N_17533);
or U22406 (N_22406,N_16055,N_19996);
xnor U22407 (N_22407,N_17007,N_19694);
xor U22408 (N_22408,N_18988,N_15605);
or U22409 (N_22409,N_15319,N_16797);
nor U22410 (N_22410,N_19289,N_16784);
or U22411 (N_22411,N_16867,N_19040);
nor U22412 (N_22412,N_18389,N_18770);
xor U22413 (N_22413,N_18837,N_16630);
nand U22414 (N_22414,N_17494,N_18188);
nand U22415 (N_22415,N_15252,N_17067);
nor U22416 (N_22416,N_16963,N_16207);
or U22417 (N_22417,N_18637,N_18055);
or U22418 (N_22418,N_16941,N_16425);
nand U22419 (N_22419,N_16812,N_15706);
or U22420 (N_22420,N_15404,N_16051);
or U22421 (N_22421,N_17197,N_19459);
nor U22422 (N_22422,N_17742,N_19828);
xnor U22423 (N_22423,N_19943,N_17111);
or U22424 (N_22424,N_15063,N_17772);
nor U22425 (N_22425,N_19275,N_15635);
nand U22426 (N_22426,N_18418,N_19405);
and U22427 (N_22427,N_15536,N_18967);
xor U22428 (N_22428,N_18569,N_16279);
or U22429 (N_22429,N_16558,N_15332);
nor U22430 (N_22430,N_15454,N_18026);
nand U22431 (N_22431,N_19351,N_15287);
nor U22432 (N_22432,N_16013,N_17716);
or U22433 (N_22433,N_18091,N_18930);
xor U22434 (N_22434,N_18821,N_17207);
and U22435 (N_22435,N_16068,N_15042);
xor U22436 (N_22436,N_19128,N_19156);
nor U22437 (N_22437,N_18850,N_16147);
and U22438 (N_22438,N_18666,N_18541);
and U22439 (N_22439,N_18774,N_18551);
and U22440 (N_22440,N_19540,N_18467);
or U22441 (N_22441,N_16174,N_17604);
nor U22442 (N_22442,N_15268,N_17099);
nand U22443 (N_22443,N_15393,N_18692);
xnor U22444 (N_22444,N_19221,N_15493);
nor U22445 (N_22445,N_18510,N_19970);
xnor U22446 (N_22446,N_19489,N_15220);
or U22447 (N_22447,N_16205,N_18867);
nand U22448 (N_22448,N_17796,N_17977);
and U22449 (N_22449,N_16804,N_18419);
or U22450 (N_22450,N_18171,N_17165);
nand U22451 (N_22451,N_15802,N_19627);
xnor U22452 (N_22452,N_15606,N_19942);
and U22453 (N_22453,N_18380,N_16447);
xor U22454 (N_22454,N_19993,N_16581);
nand U22455 (N_22455,N_15336,N_16604);
nand U22456 (N_22456,N_19104,N_18584);
or U22457 (N_22457,N_16766,N_17239);
nand U22458 (N_22458,N_15611,N_18273);
and U22459 (N_22459,N_17203,N_18760);
xnor U22460 (N_22460,N_18029,N_15638);
and U22461 (N_22461,N_17646,N_16492);
and U22462 (N_22462,N_15368,N_18447);
and U22463 (N_22463,N_16542,N_19049);
xor U22464 (N_22464,N_18400,N_15753);
and U22465 (N_22465,N_15667,N_19620);
xnor U22466 (N_22466,N_18990,N_16088);
nand U22467 (N_22467,N_19145,N_19410);
nor U22468 (N_22468,N_19659,N_18424);
nand U22469 (N_22469,N_15429,N_16011);
nand U22470 (N_22470,N_19011,N_17961);
nor U22471 (N_22471,N_15314,N_19749);
or U22472 (N_22472,N_19175,N_15628);
xnor U22473 (N_22473,N_17035,N_17100);
or U22474 (N_22474,N_17701,N_17950);
or U22475 (N_22475,N_15345,N_19908);
or U22476 (N_22476,N_19790,N_19305);
nor U22477 (N_22477,N_19223,N_15422);
nor U22478 (N_22478,N_19330,N_15566);
xor U22479 (N_22479,N_17313,N_19651);
nor U22480 (N_22480,N_18057,N_17459);
nand U22481 (N_22481,N_18984,N_16980);
xnor U22482 (N_22482,N_19492,N_18598);
or U22483 (N_22483,N_15952,N_15984);
xnor U22484 (N_22484,N_18150,N_19359);
nand U22485 (N_22485,N_18275,N_16884);
or U22486 (N_22486,N_17846,N_15860);
nor U22487 (N_22487,N_16911,N_16144);
or U22488 (N_22488,N_16674,N_15084);
and U22489 (N_22489,N_19476,N_19625);
nor U22490 (N_22490,N_15350,N_19293);
or U22491 (N_22491,N_16125,N_19640);
xnor U22492 (N_22492,N_16865,N_18970);
or U22493 (N_22493,N_19973,N_17009);
xor U22494 (N_22494,N_15644,N_16291);
and U22495 (N_22495,N_15757,N_19666);
nor U22496 (N_22496,N_15864,N_17870);
and U22497 (N_22497,N_16162,N_15920);
and U22498 (N_22498,N_19198,N_16882);
nand U22499 (N_22499,N_18433,N_18313);
or U22500 (N_22500,N_19058,N_19583);
or U22501 (N_22501,N_18497,N_15748);
nand U22502 (N_22502,N_15981,N_17137);
and U22503 (N_22503,N_17112,N_17950);
nand U22504 (N_22504,N_18575,N_16437);
nor U22505 (N_22505,N_15605,N_18464);
xor U22506 (N_22506,N_17098,N_17882);
nor U22507 (N_22507,N_15300,N_19481);
nand U22508 (N_22508,N_16334,N_18725);
or U22509 (N_22509,N_16020,N_18685);
nor U22510 (N_22510,N_18039,N_18015);
nor U22511 (N_22511,N_15295,N_18834);
and U22512 (N_22512,N_16726,N_16509);
xor U22513 (N_22513,N_18575,N_17999);
nand U22514 (N_22514,N_17584,N_16691);
or U22515 (N_22515,N_15323,N_18522);
and U22516 (N_22516,N_17206,N_15509);
xor U22517 (N_22517,N_18934,N_18363);
or U22518 (N_22518,N_17107,N_19317);
nor U22519 (N_22519,N_17585,N_16272);
and U22520 (N_22520,N_15723,N_18424);
nor U22521 (N_22521,N_16673,N_18634);
nor U22522 (N_22522,N_15880,N_17318);
nand U22523 (N_22523,N_16131,N_19311);
nor U22524 (N_22524,N_15126,N_15307);
and U22525 (N_22525,N_17969,N_15439);
nand U22526 (N_22526,N_17402,N_19027);
nor U22527 (N_22527,N_19306,N_18252);
or U22528 (N_22528,N_17086,N_16089);
xnor U22529 (N_22529,N_16782,N_17371);
or U22530 (N_22530,N_15598,N_17087);
nand U22531 (N_22531,N_16363,N_17411);
xor U22532 (N_22532,N_16705,N_17439);
or U22533 (N_22533,N_16236,N_15896);
nand U22534 (N_22534,N_17334,N_17243);
nand U22535 (N_22535,N_15463,N_15676);
or U22536 (N_22536,N_18876,N_18812);
xnor U22537 (N_22537,N_18354,N_17948);
and U22538 (N_22538,N_17861,N_17375);
nand U22539 (N_22539,N_17119,N_17171);
nor U22540 (N_22540,N_18429,N_16637);
and U22541 (N_22541,N_16528,N_16246);
or U22542 (N_22542,N_15612,N_18409);
and U22543 (N_22543,N_15974,N_16398);
or U22544 (N_22544,N_17385,N_17163);
nor U22545 (N_22545,N_19005,N_19864);
xor U22546 (N_22546,N_19685,N_18299);
nand U22547 (N_22547,N_19024,N_17141);
and U22548 (N_22548,N_16158,N_17850);
xnor U22549 (N_22549,N_18014,N_19746);
or U22550 (N_22550,N_16869,N_19343);
xnor U22551 (N_22551,N_16998,N_16298);
xnor U22552 (N_22552,N_16189,N_19313);
nor U22553 (N_22553,N_19636,N_18815);
nor U22554 (N_22554,N_16009,N_17920);
or U22555 (N_22555,N_17527,N_19518);
and U22556 (N_22556,N_19804,N_16570);
or U22557 (N_22557,N_15214,N_15765);
xor U22558 (N_22558,N_19512,N_19354);
or U22559 (N_22559,N_19990,N_15024);
nand U22560 (N_22560,N_19607,N_18944);
nand U22561 (N_22561,N_18222,N_15759);
xor U22562 (N_22562,N_17047,N_18349);
xor U22563 (N_22563,N_15777,N_16782);
nor U22564 (N_22564,N_16453,N_18578);
or U22565 (N_22565,N_17143,N_19017);
nor U22566 (N_22566,N_17497,N_15780);
xnor U22567 (N_22567,N_18162,N_15973);
and U22568 (N_22568,N_19207,N_17335);
or U22569 (N_22569,N_18258,N_17541);
xor U22570 (N_22570,N_18043,N_15936);
or U22571 (N_22571,N_18402,N_19534);
nor U22572 (N_22572,N_18094,N_18885);
and U22573 (N_22573,N_18024,N_15741);
nor U22574 (N_22574,N_18368,N_19001);
xnor U22575 (N_22575,N_17333,N_17923);
or U22576 (N_22576,N_16209,N_16123);
xnor U22577 (N_22577,N_18327,N_18056);
xor U22578 (N_22578,N_19942,N_16478);
nand U22579 (N_22579,N_19561,N_19329);
or U22580 (N_22580,N_15463,N_19836);
or U22581 (N_22581,N_17392,N_18828);
nor U22582 (N_22582,N_17788,N_17453);
nor U22583 (N_22583,N_18714,N_17815);
nor U22584 (N_22584,N_18749,N_16486);
nand U22585 (N_22585,N_17847,N_17485);
and U22586 (N_22586,N_15460,N_18336);
nor U22587 (N_22587,N_17471,N_15815);
or U22588 (N_22588,N_19972,N_19283);
nand U22589 (N_22589,N_17774,N_18935);
nand U22590 (N_22590,N_18656,N_17468);
nor U22591 (N_22591,N_18792,N_19655);
nor U22592 (N_22592,N_15482,N_17666);
xnor U22593 (N_22593,N_15599,N_15846);
nand U22594 (N_22594,N_17488,N_16611);
xnor U22595 (N_22595,N_18271,N_18136);
xor U22596 (N_22596,N_19675,N_15238);
xor U22597 (N_22597,N_15250,N_19642);
nor U22598 (N_22598,N_18648,N_17236);
and U22599 (N_22599,N_18541,N_18482);
or U22600 (N_22600,N_19295,N_16458);
nand U22601 (N_22601,N_16716,N_18033);
nor U22602 (N_22602,N_18145,N_16762);
nand U22603 (N_22603,N_18567,N_16241);
or U22604 (N_22604,N_19628,N_16879);
or U22605 (N_22605,N_15880,N_15287);
and U22606 (N_22606,N_15364,N_17142);
nor U22607 (N_22607,N_17763,N_18889);
and U22608 (N_22608,N_18565,N_19267);
xor U22609 (N_22609,N_18397,N_16528);
nand U22610 (N_22610,N_19237,N_19493);
and U22611 (N_22611,N_17693,N_16695);
nor U22612 (N_22612,N_16048,N_16392);
or U22613 (N_22613,N_15672,N_15182);
nor U22614 (N_22614,N_18131,N_17520);
nor U22615 (N_22615,N_15692,N_19082);
and U22616 (N_22616,N_17469,N_16828);
xnor U22617 (N_22617,N_16014,N_15623);
nor U22618 (N_22618,N_19741,N_17186);
nand U22619 (N_22619,N_17281,N_15157);
xnor U22620 (N_22620,N_19306,N_15849);
nor U22621 (N_22621,N_17243,N_18295);
and U22622 (N_22622,N_19278,N_15425);
nand U22623 (N_22623,N_18097,N_19780);
and U22624 (N_22624,N_19767,N_17545);
or U22625 (N_22625,N_16434,N_16454);
or U22626 (N_22626,N_16010,N_17790);
xnor U22627 (N_22627,N_17087,N_15043);
nor U22628 (N_22628,N_16624,N_16103);
or U22629 (N_22629,N_18792,N_19455);
nand U22630 (N_22630,N_16275,N_18796);
or U22631 (N_22631,N_18456,N_16167);
xor U22632 (N_22632,N_17823,N_15149);
xor U22633 (N_22633,N_19910,N_18956);
and U22634 (N_22634,N_18448,N_15389);
or U22635 (N_22635,N_19771,N_17570);
or U22636 (N_22636,N_19288,N_17309);
nand U22637 (N_22637,N_17606,N_19761);
nor U22638 (N_22638,N_15180,N_15620);
xor U22639 (N_22639,N_15337,N_15270);
and U22640 (N_22640,N_15163,N_16807);
or U22641 (N_22641,N_18280,N_19766);
or U22642 (N_22642,N_15820,N_16647);
nor U22643 (N_22643,N_17133,N_17105);
nand U22644 (N_22644,N_17185,N_17856);
xnor U22645 (N_22645,N_17252,N_17933);
or U22646 (N_22646,N_17041,N_19833);
xnor U22647 (N_22647,N_19448,N_16938);
and U22648 (N_22648,N_15957,N_16489);
or U22649 (N_22649,N_15097,N_18613);
or U22650 (N_22650,N_16254,N_19418);
nand U22651 (N_22651,N_16818,N_15981);
nor U22652 (N_22652,N_17815,N_17738);
xor U22653 (N_22653,N_17851,N_18859);
or U22654 (N_22654,N_19256,N_18700);
nand U22655 (N_22655,N_16221,N_17054);
and U22656 (N_22656,N_16150,N_16363);
nor U22657 (N_22657,N_16048,N_15900);
nand U22658 (N_22658,N_18408,N_15656);
or U22659 (N_22659,N_16460,N_15231);
nand U22660 (N_22660,N_17948,N_17587);
nand U22661 (N_22661,N_16889,N_15345);
xnor U22662 (N_22662,N_17443,N_19860);
and U22663 (N_22663,N_17313,N_15857);
xor U22664 (N_22664,N_17246,N_17309);
and U22665 (N_22665,N_15150,N_18618);
nand U22666 (N_22666,N_19400,N_15157);
nor U22667 (N_22667,N_16257,N_17710);
nor U22668 (N_22668,N_16354,N_18159);
nor U22669 (N_22669,N_16686,N_15340);
or U22670 (N_22670,N_19626,N_19901);
or U22671 (N_22671,N_16474,N_16707);
xnor U22672 (N_22672,N_17048,N_16150);
nand U22673 (N_22673,N_18468,N_18582);
nor U22674 (N_22674,N_16025,N_19051);
and U22675 (N_22675,N_18277,N_17995);
and U22676 (N_22676,N_18288,N_15954);
xnor U22677 (N_22677,N_18980,N_18000);
nor U22678 (N_22678,N_18316,N_16120);
xor U22679 (N_22679,N_19268,N_16884);
or U22680 (N_22680,N_18625,N_17579);
nor U22681 (N_22681,N_17359,N_15815);
xor U22682 (N_22682,N_16766,N_17831);
nor U22683 (N_22683,N_15640,N_16793);
nand U22684 (N_22684,N_19840,N_17120);
xnor U22685 (N_22685,N_18173,N_19515);
and U22686 (N_22686,N_19347,N_16220);
nand U22687 (N_22687,N_17245,N_19768);
or U22688 (N_22688,N_17423,N_17860);
or U22689 (N_22689,N_19890,N_18606);
nor U22690 (N_22690,N_16171,N_18427);
nand U22691 (N_22691,N_18565,N_15697);
nor U22692 (N_22692,N_18038,N_19252);
and U22693 (N_22693,N_17056,N_16695);
nor U22694 (N_22694,N_16262,N_15796);
nand U22695 (N_22695,N_19859,N_16276);
nor U22696 (N_22696,N_16926,N_18682);
or U22697 (N_22697,N_16604,N_18647);
xor U22698 (N_22698,N_18953,N_18524);
nand U22699 (N_22699,N_19801,N_18378);
xnor U22700 (N_22700,N_16851,N_18974);
nand U22701 (N_22701,N_19004,N_19860);
xor U22702 (N_22702,N_19455,N_15294);
or U22703 (N_22703,N_15786,N_17219);
and U22704 (N_22704,N_17498,N_16968);
or U22705 (N_22705,N_19526,N_19152);
or U22706 (N_22706,N_16239,N_16333);
nand U22707 (N_22707,N_15590,N_15034);
and U22708 (N_22708,N_16231,N_15466);
or U22709 (N_22709,N_15838,N_19586);
and U22710 (N_22710,N_19815,N_15986);
nand U22711 (N_22711,N_17022,N_17866);
nand U22712 (N_22712,N_17324,N_17548);
or U22713 (N_22713,N_19808,N_17025);
or U22714 (N_22714,N_18586,N_19480);
and U22715 (N_22715,N_18739,N_19992);
nor U22716 (N_22716,N_15178,N_15725);
or U22717 (N_22717,N_18714,N_16041);
and U22718 (N_22718,N_17024,N_19961);
and U22719 (N_22719,N_15954,N_19209);
nor U22720 (N_22720,N_17861,N_16741);
xor U22721 (N_22721,N_19405,N_16751);
nor U22722 (N_22722,N_18807,N_16600);
and U22723 (N_22723,N_17148,N_18075);
xor U22724 (N_22724,N_18293,N_17137);
xor U22725 (N_22725,N_19593,N_15750);
or U22726 (N_22726,N_19982,N_19317);
or U22727 (N_22727,N_17199,N_15252);
nand U22728 (N_22728,N_16371,N_15781);
nand U22729 (N_22729,N_16287,N_15990);
and U22730 (N_22730,N_18487,N_18893);
nor U22731 (N_22731,N_16557,N_16459);
and U22732 (N_22732,N_16137,N_15111);
and U22733 (N_22733,N_18920,N_16798);
xnor U22734 (N_22734,N_18371,N_15315);
nand U22735 (N_22735,N_16669,N_18914);
nor U22736 (N_22736,N_19267,N_18836);
and U22737 (N_22737,N_17899,N_19639);
or U22738 (N_22738,N_19179,N_16598);
and U22739 (N_22739,N_15272,N_17802);
nor U22740 (N_22740,N_18637,N_17954);
xor U22741 (N_22741,N_17383,N_15247);
and U22742 (N_22742,N_17385,N_19755);
or U22743 (N_22743,N_18265,N_18080);
xnor U22744 (N_22744,N_15609,N_19424);
xnor U22745 (N_22745,N_19370,N_16832);
or U22746 (N_22746,N_19244,N_19588);
nor U22747 (N_22747,N_18123,N_15819);
nand U22748 (N_22748,N_15287,N_17594);
nand U22749 (N_22749,N_19666,N_19690);
or U22750 (N_22750,N_18260,N_15736);
xor U22751 (N_22751,N_17909,N_17455);
or U22752 (N_22752,N_16345,N_18526);
xnor U22753 (N_22753,N_19551,N_18819);
and U22754 (N_22754,N_18113,N_15961);
nand U22755 (N_22755,N_18457,N_18697);
or U22756 (N_22756,N_17701,N_16640);
or U22757 (N_22757,N_15240,N_18850);
xor U22758 (N_22758,N_19728,N_18650);
or U22759 (N_22759,N_15639,N_17195);
or U22760 (N_22760,N_19673,N_16870);
or U22761 (N_22761,N_17404,N_19439);
or U22762 (N_22762,N_18810,N_17605);
or U22763 (N_22763,N_16193,N_16870);
and U22764 (N_22764,N_15905,N_15609);
nor U22765 (N_22765,N_17225,N_17819);
nand U22766 (N_22766,N_18672,N_16029);
nor U22767 (N_22767,N_15574,N_17429);
and U22768 (N_22768,N_16836,N_17770);
or U22769 (N_22769,N_19372,N_18648);
nand U22770 (N_22770,N_16778,N_19049);
nand U22771 (N_22771,N_18265,N_19285);
xor U22772 (N_22772,N_19305,N_18708);
xnor U22773 (N_22773,N_15668,N_15926);
or U22774 (N_22774,N_15916,N_17551);
xnor U22775 (N_22775,N_16073,N_15898);
nor U22776 (N_22776,N_19267,N_16219);
nand U22777 (N_22777,N_17862,N_19304);
or U22778 (N_22778,N_19294,N_17568);
or U22779 (N_22779,N_19398,N_19310);
and U22780 (N_22780,N_19418,N_17289);
and U22781 (N_22781,N_18883,N_18524);
xnor U22782 (N_22782,N_17155,N_16286);
xnor U22783 (N_22783,N_17725,N_17058);
xor U22784 (N_22784,N_16323,N_16050);
or U22785 (N_22785,N_17072,N_16880);
nor U22786 (N_22786,N_17545,N_18980);
and U22787 (N_22787,N_18759,N_16123);
or U22788 (N_22788,N_19146,N_17176);
xnor U22789 (N_22789,N_17106,N_19491);
and U22790 (N_22790,N_18013,N_18591);
nor U22791 (N_22791,N_19003,N_19511);
or U22792 (N_22792,N_17003,N_19198);
nor U22793 (N_22793,N_18460,N_16090);
and U22794 (N_22794,N_15538,N_18078);
and U22795 (N_22795,N_16777,N_18093);
nor U22796 (N_22796,N_19341,N_19096);
nand U22797 (N_22797,N_16097,N_15976);
or U22798 (N_22798,N_15616,N_17197);
and U22799 (N_22799,N_16613,N_15286);
or U22800 (N_22800,N_16779,N_16791);
or U22801 (N_22801,N_15614,N_17473);
nor U22802 (N_22802,N_19856,N_15273);
and U22803 (N_22803,N_18154,N_15733);
xnor U22804 (N_22804,N_16044,N_16431);
or U22805 (N_22805,N_15044,N_18970);
and U22806 (N_22806,N_16616,N_18747);
or U22807 (N_22807,N_16441,N_18084);
nor U22808 (N_22808,N_17558,N_18216);
xnor U22809 (N_22809,N_15138,N_18577);
or U22810 (N_22810,N_15815,N_18007);
or U22811 (N_22811,N_18478,N_16972);
and U22812 (N_22812,N_16922,N_17261);
nor U22813 (N_22813,N_16150,N_17928);
xor U22814 (N_22814,N_16974,N_16255);
xnor U22815 (N_22815,N_19149,N_15718);
or U22816 (N_22816,N_15231,N_18210);
and U22817 (N_22817,N_17572,N_18480);
xor U22818 (N_22818,N_17554,N_18058);
or U22819 (N_22819,N_19313,N_19132);
xnor U22820 (N_22820,N_18406,N_17995);
or U22821 (N_22821,N_17102,N_19789);
nor U22822 (N_22822,N_15872,N_19202);
and U22823 (N_22823,N_17603,N_17564);
nor U22824 (N_22824,N_16107,N_17401);
xor U22825 (N_22825,N_19167,N_17636);
xor U22826 (N_22826,N_17839,N_17260);
nor U22827 (N_22827,N_18614,N_19052);
xnor U22828 (N_22828,N_15056,N_15368);
and U22829 (N_22829,N_17938,N_19935);
nand U22830 (N_22830,N_18266,N_18030);
xnor U22831 (N_22831,N_15015,N_19033);
or U22832 (N_22832,N_19027,N_19437);
xnor U22833 (N_22833,N_18185,N_19376);
xnor U22834 (N_22834,N_17985,N_16263);
or U22835 (N_22835,N_19442,N_15237);
nand U22836 (N_22836,N_15741,N_15188);
nor U22837 (N_22837,N_17900,N_15980);
or U22838 (N_22838,N_19982,N_17022);
and U22839 (N_22839,N_18926,N_16732);
nor U22840 (N_22840,N_19984,N_15813);
nand U22841 (N_22841,N_17662,N_16061);
or U22842 (N_22842,N_18001,N_15462);
nor U22843 (N_22843,N_18183,N_17364);
or U22844 (N_22844,N_15253,N_16439);
or U22845 (N_22845,N_19342,N_17223);
nand U22846 (N_22846,N_16779,N_18671);
nor U22847 (N_22847,N_18473,N_19245);
nand U22848 (N_22848,N_18801,N_16464);
or U22849 (N_22849,N_17922,N_18352);
and U22850 (N_22850,N_15517,N_19423);
nand U22851 (N_22851,N_16951,N_19667);
or U22852 (N_22852,N_16610,N_19035);
nor U22853 (N_22853,N_15273,N_15885);
nor U22854 (N_22854,N_15456,N_16070);
xor U22855 (N_22855,N_17887,N_18010);
xor U22856 (N_22856,N_19682,N_15359);
nor U22857 (N_22857,N_19646,N_19558);
or U22858 (N_22858,N_18788,N_15121);
or U22859 (N_22859,N_18784,N_16988);
xor U22860 (N_22860,N_18932,N_15140);
nand U22861 (N_22861,N_18163,N_18435);
xnor U22862 (N_22862,N_15353,N_18513);
nor U22863 (N_22863,N_16677,N_18207);
nor U22864 (N_22864,N_17065,N_17842);
xor U22865 (N_22865,N_18191,N_15227);
xnor U22866 (N_22866,N_17114,N_19767);
xor U22867 (N_22867,N_17439,N_18446);
xnor U22868 (N_22868,N_15850,N_16401);
nand U22869 (N_22869,N_17715,N_17781);
and U22870 (N_22870,N_18313,N_15600);
xnor U22871 (N_22871,N_17241,N_18001);
xor U22872 (N_22872,N_19181,N_15297);
nand U22873 (N_22873,N_15471,N_19355);
nor U22874 (N_22874,N_15708,N_16942);
nor U22875 (N_22875,N_17821,N_19086);
nor U22876 (N_22876,N_19384,N_19423);
and U22877 (N_22877,N_16317,N_16674);
or U22878 (N_22878,N_19377,N_15680);
and U22879 (N_22879,N_18736,N_17976);
and U22880 (N_22880,N_16384,N_16582);
nand U22881 (N_22881,N_16635,N_17923);
nor U22882 (N_22882,N_16366,N_15501);
and U22883 (N_22883,N_18894,N_16280);
and U22884 (N_22884,N_16742,N_16236);
nand U22885 (N_22885,N_15297,N_17748);
xor U22886 (N_22886,N_15421,N_19509);
or U22887 (N_22887,N_19742,N_18651);
xor U22888 (N_22888,N_17487,N_16599);
nor U22889 (N_22889,N_19888,N_17856);
xnor U22890 (N_22890,N_17140,N_16622);
or U22891 (N_22891,N_17103,N_15640);
xnor U22892 (N_22892,N_17407,N_17682);
or U22893 (N_22893,N_18521,N_16449);
or U22894 (N_22894,N_17445,N_17435);
xor U22895 (N_22895,N_15546,N_17938);
nor U22896 (N_22896,N_16133,N_17383);
nand U22897 (N_22897,N_19923,N_17684);
nand U22898 (N_22898,N_19998,N_16427);
or U22899 (N_22899,N_15627,N_19059);
or U22900 (N_22900,N_18272,N_15237);
nand U22901 (N_22901,N_19531,N_17395);
nand U22902 (N_22902,N_16615,N_15241);
nor U22903 (N_22903,N_18233,N_19484);
or U22904 (N_22904,N_16186,N_15940);
nand U22905 (N_22905,N_15189,N_19231);
nand U22906 (N_22906,N_19410,N_15329);
or U22907 (N_22907,N_16817,N_19286);
xor U22908 (N_22908,N_19022,N_17080);
nand U22909 (N_22909,N_16737,N_16611);
nand U22910 (N_22910,N_18517,N_18233);
nor U22911 (N_22911,N_16053,N_16112);
nor U22912 (N_22912,N_18027,N_16661);
xnor U22913 (N_22913,N_15695,N_19105);
nor U22914 (N_22914,N_19257,N_15719);
and U22915 (N_22915,N_16173,N_16750);
or U22916 (N_22916,N_18756,N_16940);
nand U22917 (N_22917,N_17856,N_15833);
and U22918 (N_22918,N_17292,N_18540);
or U22919 (N_22919,N_15490,N_18754);
nor U22920 (N_22920,N_16289,N_15777);
xnor U22921 (N_22921,N_18241,N_19444);
nand U22922 (N_22922,N_16439,N_19019);
xnor U22923 (N_22923,N_19603,N_15439);
nand U22924 (N_22924,N_16550,N_16365);
nand U22925 (N_22925,N_16952,N_19846);
or U22926 (N_22926,N_19860,N_18279);
nor U22927 (N_22927,N_16172,N_17072);
xnor U22928 (N_22928,N_18552,N_19135);
and U22929 (N_22929,N_15196,N_15345);
or U22930 (N_22930,N_18038,N_17138);
and U22931 (N_22931,N_17701,N_16314);
xor U22932 (N_22932,N_15732,N_17289);
xnor U22933 (N_22933,N_17544,N_16145);
and U22934 (N_22934,N_17374,N_15944);
xor U22935 (N_22935,N_16338,N_19487);
and U22936 (N_22936,N_17861,N_15846);
or U22937 (N_22937,N_16291,N_18701);
xor U22938 (N_22938,N_17394,N_18124);
nand U22939 (N_22939,N_18677,N_19946);
nor U22940 (N_22940,N_19155,N_19588);
nor U22941 (N_22941,N_17552,N_16604);
xnor U22942 (N_22942,N_19222,N_16044);
nand U22943 (N_22943,N_17755,N_18577);
and U22944 (N_22944,N_18857,N_18799);
or U22945 (N_22945,N_19238,N_19129);
xor U22946 (N_22946,N_16613,N_15716);
nand U22947 (N_22947,N_17978,N_17792);
nor U22948 (N_22948,N_15049,N_15382);
xnor U22949 (N_22949,N_16994,N_18846);
nor U22950 (N_22950,N_16705,N_19448);
xnor U22951 (N_22951,N_15136,N_19200);
nand U22952 (N_22952,N_15422,N_18790);
nor U22953 (N_22953,N_19339,N_19969);
or U22954 (N_22954,N_15031,N_17106);
xor U22955 (N_22955,N_16661,N_17693);
or U22956 (N_22956,N_17918,N_16974);
xor U22957 (N_22957,N_18225,N_19510);
nand U22958 (N_22958,N_18680,N_15022);
xor U22959 (N_22959,N_15233,N_16795);
nand U22960 (N_22960,N_18764,N_17343);
nand U22961 (N_22961,N_19644,N_18282);
or U22962 (N_22962,N_17046,N_15174);
or U22963 (N_22963,N_19747,N_17679);
xor U22964 (N_22964,N_18961,N_18434);
nand U22965 (N_22965,N_15510,N_15828);
or U22966 (N_22966,N_19476,N_16397);
nor U22967 (N_22967,N_17289,N_15364);
nor U22968 (N_22968,N_16144,N_15024);
nor U22969 (N_22969,N_17811,N_19420);
xor U22970 (N_22970,N_17484,N_15727);
or U22971 (N_22971,N_18633,N_18830);
or U22972 (N_22972,N_17119,N_18580);
and U22973 (N_22973,N_19366,N_17105);
nor U22974 (N_22974,N_19277,N_18584);
nor U22975 (N_22975,N_19709,N_17038);
and U22976 (N_22976,N_17010,N_17197);
nor U22977 (N_22977,N_18046,N_19193);
nor U22978 (N_22978,N_15058,N_18162);
or U22979 (N_22979,N_16164,N_18702);
nand U22980 (N_22980,N_19665,N_18752);
nand U22981 (N_22981,N_15437,N_18856);
nor U22982 (N_22982,N_16458,N_18333);
nor U22983 (N_22983,N_18889,N_15032);
or U22984 (N_22984,N_16309,N_17286);
or U22985 (N_22985,N_15738,N_18617);
xnor U22986 (N_22986,N_15214,N_17605);
nand U22987 (N_22987,N_15699,N_18158);
xnor U22988 (N_22988,N_16880,N_15952);
and U22989 (N_22989,N_15338,N_16399);
nand U22990 (N_22990,N_16161,N_18733);
and U22991 (N_22991,N_18029,N_18778);
nand U22992 (N_22992,N_17265,N_19711);
nand U22993 (N_22993,N_15145,N_19599);
and U22994 (N_22994,N_16180,N_17271);
nor U22995 (N_22995,N_19600,N_15533);
or U22996 (N_22996,N_17032,N_19095);
xor U22997 (N_22997,N_15647,N_15209);
nor U22998 (N_22998,N_15526,N_17158);
nor U22999 (N_22999,N_16295,N_17551);
nor U23000 (N_23000,N_15041,N_15455);
nand U23001 (N_23001,N_15869,N_15524);
nor U23002 (N_23002,N_19066,N_19194);
or U23003 (N_23003,N_15699,N_17551);
nor U23004 (N_23004,N_19958,N_16218);
nand U23005 (N_23005,N_15034,N_16319);
xor U23006 (N_23006,N_16744,N_17248);
xnor U23007 (N_23007,N_17470,N_16179);
xnor U23008 (N_23008,N_17744,N_15025);
xnor U23009 (N_23009,N_19961,N_17363);
nor U23010 (N_23010,N_19616,N_17557);
nand U23011 (N_23011,N_19554,N_16015);
xnor U23012 (N_23012,N_15427,N_16015);
nor U23013 (N_23013,N_16268,N_17417);
nand U23014 (N_23014,N_17998,N_15437);
or U23015 (N_23015,N_16555,N_15034);
xnor U23016 (N_23016,N_16994,N_17858);
nand U23017 (N_23017,N_16967,N_16359);
or U23018 (N_23018,N_15000,N_15967);
nor U23019 (N_23019,N_16009,N_18989);
or U23020 (N_23020,N_16054,N_18517);
and U23021 (N_23021,N_15058,N_19336);
and U23022 (N_23022,N_18491,N_19506);
nand U23023 (N_23023,N_16607,N_15822);
or U23024 (N_23024,N_15562,N_15471);
and U23025 (N_23025,N_19614,N_19163);
nand U23026 (N_23026,N_17636,N_16791);
and U23027 (N_23027,N_18819,N_18279);
or U23028 (N_23028,N_18671,N_17836);
and U23029 (N_23029,N_19351,N_16697);
nor U23030 (N_23030,N_18277,N_19184);
nor U23031 (N_23031,N_15632,N_19766);
xor U23032 (N_23032,N_16662,N_15850);
nor U23033 (N_23033,N_17846,N_19726);
nor U23034 (N_23034,N_19388,N_17902);
and U23035 (N_23035,N_17471,N_16920);
xnor U23036 (N_23036,N_16938,N_18207);
nand U23037 (N_23037,N_18761,N_19974);
and U23038 (N_23038,N_19748,N_18908);
nand U23039 (N_23039,N_19051,N_19424);
nand U23040 (N_23040,N_16467,N_17834);
and U23041 (N_23041,N_15974,N_16826);
nand U23042 (N_23042,N_18943,N_15335);
nand U23043 (N_23043,N_17269,N_16063);
nand U23044 (N_23044,N_18499,N_17130);
nor U23045 (N_23045,N_19237,N_19930);
nand U23046 (N_23046,N_19934,N_15294);
xor U23047 (N_23047,N_15678,N_16168);
and U23048 (N_23048,N_17119,N_15294);
nor U23049 (N_23049,N_15668,N_17752);
xor U23050 (N_23050,N_16833,N_15711);
nor U23051 (N_23051,N_16673,N_18512);
nand U23052 (N_23052,N_18100,N_17145);
and U23053 (N_23053,N_18951,N_16733);
xor U23054 (N_23054,N_16560,N_16430);
xnor U23055 (N_23055,N_17564,N_18061);
nor U23056 (N_23056,N_17549,N_15344);
nor U23057 (N_23057,N_16810,N_19140);
xor U23058 (N_23058,N_15731,N_18759);
and U23059 (N_23059,N_18176,N_18430);
nand U23060 (N_23060,N_19874,N_19153);
nor U23061 (N_23061,N_16509,N_15471);
nor U23062 (N_23062,N_15402,N_18310);
and U23063 (N_23063,N_19015,N_17496);
xor U23064 (N_23064,N_17621,N_19134);
xnor U23065 (N_23065,N_19033,N_15006);
nand U23066 (N_23066,N_19400,N_19792);
nand U23067 (N_23067,N_19794,N_16162);
and U23068 (N_23068,N_16712,N_17980);
xor U23069 (N_23069,N_16593,N_15965);
and U23070 (N_23070,N_18653,N_15362);
xnor U23071 (N_23071,N_17610,N_18368);
and U23072 (N_23072,N_16646,N_16269);
or U23073 (N_23073,N_16067,N_16847);
or U23074 (N_23074,N_15391,N_18324);
xor U23075 (N_23075,N_16597,N_17239);
nor U23076 (N_23076,N_15374,N_15207);
xnor U23077 (N_23077,N_15449,N_18110);
xor U23078 (N_23078,N_15118,N_19131);
nor U23079 (N_23079,N_17042,N_18405);
nand U23080 (N_23080,N_15108,N_19188);
nand U23081 (N_23081,N_17773,N_19472);
and U23082 (N_23082,N_19454,N_19908);
nor U23083 (N_23083,N_17939,N_17817);
and U23084 (N_23084,N_17576,N_16442);
nor U23085 (N_23085,N_15354,N_17654);
and U23086 (N_23086,N_18879,N_18213);
nor U23087 (N_23087,N_16677,N_15816);
nand U23088 (N_23088,N_15286,N_19597);
or U23089 (N_23089,N_18983,N_17114);
xnor U23090 (N_23090,N_15573,N_17041);
or U23091 (N_23091,N_19799,N_17555);
and U23092 (N_23092,N_19796,N_18168);
and U23093 (N_23093,N_17667,N_19683);
and U23094 (N_23094,N_16129,N_17142);
nand U23095 (N_23095,N_17570,N_16051);
or U23096 (N_23096,N_16766,N_16972);
xnor U23097 (N_23097,N_17059,N_15308);
or U23098 (N_23098,N_17826,N_17993);
xor U23099 (N_23099,N_15675,N_16941);
nand U23100 (N_23100,N_19215,N_18638);
or U23101 (N_23101,N_16098,N_18608);
nand U23102 (N_23102,N_16337,N_16841);
xnor U23103 (N_23103,N_18999,N_16976);
and U23104 (N_23104,N_18563,N_17555);
nor U23105 (N_23105,N_15093,N_18508);
and U23106 (N_23106,N_17560,N_15088);
nor U23107 (N_23107,N_16372,N_17345);
xor U23108 (N_23108,N_18259,N_16086);
nor U23109 (N_23109,N_19343,N_16489);
xnor U23110 (N_23110,N_18234,N_16168);
xor U23111 (N_23111,N_19704,N_16131);
or U23112 (N_23112,N_16060,N_19405);
nand U23113 (N_23113,N_19878,N_16677);
nor U23114 (N_23114,N_19061,N_19550);
or U23115 (N_23115,N_15478,N_17377);
nand U23116 (N_23116,N_15562,N_17959);
xor U23117 (N_23117,N_19397,N_18082);
and U23118 (N_23118,N_17360,N_17108);
nand U23119 (N_23119,N_19804,N_18271);
nand U23120 (N_23120,N_17227,N_16641);
nand U23121 (N_23121,N_19633,N_19625);
nand U23122 (N_23122,N_16437,N_15313);
or U23123 (N_23123,N_15637,N_18926);
nand U23124 (N_23124,N_19087,N_15922);
nand U23125 (N_23125,N_19019,N_15936);
and U23126 (N_23126,N_16519,N_18016);
nand U23127 (N_23127,N_17980,N_17158);
nor U23128 (N_23128,N_15303,N_15983);
xor U23129 (N_23129,N_15838,N_16932);
and U23130 (N_23130,N_15608,N_19995);
nor U23131 (N_23131,N_18321,N_15155);
or U23132 (N_23132,N_19760,N_16362);
xnor U23133 (N_23133,N_15501,N_16151);
or U23134 (N_23134,N_19915,N_17776);
or U23135 (N_23135,N_17235,N_18588);
or U23136 (N_23136,N_17617,N_18016);
nor U23137 (N_23137,N_17662,N_18838);
nor U23138 (N_23138,N_16321,N_18417);
xnor U23139 (N_23139,N_17628,N_16889);
xor U23140 (N_23140,N_17278,N_17744);
and U23141 (N_23141,N_19668,N_15793);
and U23142 (N_23142,N_16308,N_15703);
and U23143 (N_23143,N_19407,N_16057);
nor U23144 (N_23144,N_18717,N_16058);
xor U23145 (N_23145,N_17437,N_17374);
nand U23146 (N_23146,N_15315,N_19698);
nand U23147 (N_23147,N_15328,N_15077);
nor U23148 (N_23148,N_17182,N_17400);
nor U23149 (N_23149,N_18882,N_17042);
xnor U23150 (N_23150,N_18467,N_19757);
nand U23151 (N_23151,N_17734,N_18989);
nor U23152 (N_23152,N_17614,N_19607);
or U23153 (N_23153,N_19450,N_15862);
or U23154 (N_23154,N_15011,N_18213);
nor U23155 (N_23155,N_15929,N_17412);
nand U23156 (N_23156,N_19790,N_18377);
xnor U23157 (N_23157,N_19085,N_17668);
xnor U23158 (N_23158,N_16349,N_19693);
or U23159 (N_23159,N_15265,N_19868);
or U23160 (N_23160,N_15132,N_18403);
and U23161 (N_23161,N_18173,N_16612);
nand U23162 (N_23162,N_18686,N_17438);
nor U23163 (N_23163,N_19291,N_17964);
xnor U23164 (N_23164,N_16067,N_17357);
xnor U23165 (N_23165,N_18734,N_15134);
xnor U23166 (N_23166,N_15915,N_18378);
xor U23167 (N_23167,N_17410,N_17320);
nand U23168 (N_23168,N_15488,N_16421);
nor U23169 (N_23169,N_15397,N_17517);
nor U23170 (N_23170,N_15493,N_17952);
nor U23171 (N_23171,N_19407,N_16952);
or U23172 (N_23172,N_18682,N_19784);
nand U23173 (N_23173,N_16762,N_19138);
nor U23174 (N_23174,N_19064,N_15215);
and U23175 (N_23175,N_19600,N_16716);
xnor U23176 (N_23176,N_15262,N_15843);
and U23177 (N_23177,N_16143,N_16809);
nand U23178 (N_23178,N_19715,N_18947);
or U23179 (N_23179,N_17271,N_15472);
xor U23180 (N_23180,N_15269,N_16040);
nor U23181 (N_23181,N_16964,N_18800);
or U23182 (N_23182,N_17956,N_15605);
xnor U23183 (N_23183,N_17946,N_18569);
xnor U23184 (N_23184,N_18178,N_16081);
xnor U23185 (N_23185,N_19478,N_15906);
nand U23186 (N_23186,N_16828,N_18981);
xor U23187 (N_23187,N_19785,N_18338);
or U23188 (N_23188,N_17705,N_15770);
or U23189 (N_23189,N_16695,N_19073);
and U23190 (N_23190,N_17173,N_18155);
nor U23191 (N_23191,N_17957,N_19572);
or U23192 (N_23192,N_16139,N_16274);
nand U23193 (N_23193,N_15346,N_18338);
and U23194 (N_23194,N_16300,N_18986);
and U23195 (N_23195,N_17746,N_18437);
xor U23196 (N_23196,N_19684,N_15113);
nand U23197 (N_23197,N_19206,N_15425);
nand U23198 (N_23198,N_17715,N_16470);
or U23199 (N_23199,N_17514,N_17703);
or U23200 (N_23200,N_18740,N_19818);
nand U23201 (N_23201,N_18394,N_15405);
or U23202 (N_23202,N_17579,N_17589);
nand U23203 (N_23203,N_19131,N_15448);
xnor U23204 (N_23204,N_18446,N_17832);
nand U23205 (N_23205,N_19112,N_16234);
and U23206 (N_23206,N_17180,N_15486);
or U23207 (N_23207,N_18881,N_15337);
nand U23208 (N_23208,N_15421,N_18644);
or U23209 (N_23209,N_19284,N_17446);
or U23210 (N_23210,N_19092,N_19040);
and U23211 (N_23211,N_16133,N_16330);
nor U23212 (N_23212,N_15077,N_16861);
and U23213 (N_23213,N_16579,N_16073);
nor U23214 (N_23214,N_16858,N_19275);
xnor U23215 (N_23215,N_17028,N_17155);
and U23216 (N_23216,N_17959,N_15971);
and U23217 (N_23217,N_18086,N_15790);
and U23218 (N_23218,N_18952,N_16049);
nor U23219 (N_23219,N_16094,N_19186);
and U23220 (N_23220,N_19733,N_15897);
nor U23221 (N_23221,N_18436,N_17191);
nand U23222 (N_23222,N_16603,N_15057);
xnor U23223 (N_23223,N_18010,N_17008);
nor U23224 (N_23224,N_15234,N_16993);
and U23225 (N_23225,N_19554,N_16300);
xnor U23226 (N_23226,N_16097,N_19827);
or U23227 (N_23227,N_18325,N_15025);
nand U23228 (N_23228,N_18551,N_19018);
and U23229 (N_23229,N_16192,N_16150);
or U23230 (N_23230,N_15098,N_18946);
nor U23231 (N_23231,N_19269,N_16004);
nor U23232 (N_23232,N_15631,N_19487);
nor U23233 (N_23233,N_18494,N_18339);
and U23234 (N_23234,N_18467,N_19754);
nand U23235 (N_23235,N_18489,N_18607);
nor U23236 (N_23236,N_18663,N_19193);
nor U23237 (N_23237,N_18787,N_19479);
or U23238 (N_23238,N_16718,N_19727);
xor U23239 (N_23239,N_15662,N_15020);
xnor U23240 (N_23240,N_17112,N_19276);
nand U23241 (N_23241,N_16881,N_17956);
and U23242 (N_23242,N_19324,N_17129);
and U23243 (N_23243,N_19140,N_16328);
or U23244 (N_23244,N_15447,N_17370);
xnor U23245 (N_23245,N_15969,N_18667);
or U23246 (N_23246,N_16317,N_16727);
xnor U23247 (N_23247,N_16351,N_15067);
xor U23248 (N_23248,N_17985,N_15310);
nand U23249 (N_23249,N_15195,N_17614);
xor U23250 (N_23250,N_16562,N_16164);
nand U23251 (N_23251,N_15390,N_19815);
nor U23252 (N_23252,N_19090,N_17904);
xnor U23253 (N_23253,N_17992,N_19321);
and U23254 (N_23254,N_15352,N_15942);
xnor U23255 (N_23255,N_17350,N_19846);
and U23256 (N_23256,N_15031,N_17513);
nor U23257 (N_23257,N_15544,N_16417);
or U23258 (N_23258,N_19528,N_19327);
nor U23259 (N_23259,N_15073,N_18011);
xnor U23260 (N_23260,N_17326,N_18413);
and U23261 (N_23261,N_16962,N_17123);
nand U23262 (N_23262,N_15628,N_19220);
nor U23263 (N_23263,N_18261,N_19857);
nand U23264 (N_23264,N_15240,N_17406);
nand U23265 (N_23265,N_16832,N_17383);
and U23266 (N_23266,N_19734,N_19796);
nand U23267 (N_23267,N_19907,N_18212);
nand U23268 (N_23268,N_16369,N_16590);
nor U23269 (N_23269,N_15505,N_19439);
and U23270 (N_23270,N_16954,N_18169);
xor U23271 (N_23271,N_19075,N_16027);
and U23272 (N_23272,N_19084,N_17824);
or U23273 (N_23273,N_19325,N_16817);
nor U23274 (N_23274,N_19368,N_15438);
or U23275 (N_23275,N_18216,N_16635);
or U23276 (N_23276,N_18394,N_15544);
nor U23277 (N_23277,N_16738,N_16922);
nor U23278 (N_23278,N_16333,N_17587);
or U23279 (N_23279,N_15017,N_15621);
xnor U23280 (N_23280,N_15671,N_16543);
nor U23281 (N_23281,N_15146,N_19454);
xor U23282 (N_23282,N_16196,N_18445);
or U23283 (N_23283,N_17382,N_15952);
and U23284 (N_23284,N_18596,N_16304);
and U23285 (N_23285,N_15125,N_16502);
and U23286 (N_23286,N_18957,N_15171);
nor U23287 (N_23287,N_19171,N_19214);
or U23288 (N_23288,N_18527,N_16914);
nand U23289 (N_23289,N_18710,N_17745);
xnor U23290 (N_23290,N_17874,N_16237);
or U23291 (N_23291,N_17409,N_19909);
nor U23292 (N_23292,N_19086,N_16260);
nor U23293 (N_23293,N_18547,N_19870);
xnor U23294 (N_23294,N_15436,N_18200);
or U23295 (N_23295,N_18983,N_18111);
and U23296 (N_23296,N_18869,N_15553);
and U23297 (N_23297,N_16224,N_19496);
nand U23298 (N_23298,N_18218,N_18069);
nand U23299 (N_23299,N_18412,N_19327);
nor U23300 (N_23300,N_19484,N_17050);
nor U23301 (N_23301,N_15233,N_18791);
xor U23302 (N_23302,N_15512,N_19940);
and U23303 (N_23303,N_17228,N_17950);
xnor U23304 (N_23304,N_19362,N_17923);
xnor U23305 (N_23305,N_16701,N_16261);
xnor U23306 (N_23306,N_15413,N_18170);
nor U23307 (N_23307,N_19753,N_16764);
xor U23308 (N_23308,N_19951,N_16894);
nor U23309 (N_23309,N_19931,N_16675);
nand U23310 (N_23310,N_17847,N_18420);
xnor U23311 (N_23311,N_18649,N_16078);
or U23312 (N_23312,N_16527,N_15248);
nor U23313 (N_23313,N_19635,N_15342);
xor U23314 (N_23314,N_15050,N_18366);
nand U23315 (N_23315,N_18803,N_16304);
nor U23316 (N_23316,N_19707,N_19453);
nor U23317 (N_23317,N_18502,N_16223);
nor U23318 (N_23318,N_15315,N_16091);
xnor U23319 (N_23319,N_18215,N_19345);
nand U23320 (N_23320,N_16999,N_15774);
and U23321 (N_23321,N_15870,N_19443);
xnor U23322 (N_23322,N_15385,N_15008);
or U23323 (N_23323,N_16330,N_16518);
xor U23324 (N_23324,N_16969,N_18359);
or U23325 (N_23325,N_15965,N_16679);
nor U23326 (N_23326,N_18066,N_15995);
xnor U23327 (N_23327,N_16726,N_16955);
and U23328 (N_23328,N_16799,N_15592);
or U23329 (N_23329,N_18440,N_19245);
nand U23330 (N_23330,N_17575,N_16907);
nor U23331 (N_23331,N_16197,N_15539);
xnor U23332 (N_23332,N_16181,N_18141);
xnor U23333 (N_23333,N_18682,N_18873);
and U23334 (N_23334,N_19886,N_15834);
nor U23335 (N_23335,N_17644,N_15881);
and U23336 (N_23336,N_19017,N_17384);
and U23337 (N_23337,N_17873,N_17232);
and U23338 (N_23338,N_18775,N_17738);
or U23339 (N_23339,N_18940,N_17112);
and U23340 (N_23340,N_18459,N_15116);
xor U23341 (N_23341,N_17106,N_19832);
or U23342 (N_23342,N_18844,N_15640);
nand U23343 (N_23343,N_15105,N_16298);
xnor U23344 (N_23344,N_16736,N_18424);
nand U23345 (N_23345,N_16315,N_17627);
or U23346 (N_23346,N_18693,N_15219);
and U23347 (N_23347,N_17426,N_16571);
or U23348 (N_23348,N_17568,N_18634);
nand U23349 (N_23349,N_19350,N_19440);
nor U23350 (N_23350,N_18155,N_19359);
and U23351 (N_23351,N_18233,N_19726);
xor U23352 (N_23352,N_17084,N_17676);
xor U23353 (N_23353,N_17863,N_18120);
and U23354 (N_23354,N_17122,N_18855);
and U23355 (N_23355,N_17520,N_19069);
xor U23356 (N_23356,N_17167,N_19651);
or U23357 (N_23357,N_19076,N_19354);
and U23358 (N_23358,N_16586,N_16172);
nand U23359 (N_23359,N_17050,N_19579);
or U23360 (N_23360,N_18113,N_16851);
nor U23361 (N_23361,N_18277,N_17317);
and U23362 (N_23362,N_16523,N_17952);
nor U23363 (N_23363,N_17194,N_15449);
xor U23364 (N_23364,N_18946,N_15661);
xnor U23365 (N_23365,N_18083,N_17567);
or U23366 (N_23366,N_15028,N_19498);
nand U23367 (N_23367,N_16539,N_18061);
xor U23368 (N_23368,N_18408,N_18508);
nand U23369 (N_23369,N_16945,N_17711);
xor U23370 (N_23370,N_15014,N_18972);
xor U23371 (N_23371,N_15274,N_16761);
xnor U23372 (N_23372,N_18475,N_18807);
and U23373 (N_23373,N_18892,N_17019);
xnor U23374 (N_23374,N_16234,N_19004);
xor U23375 (N_23375,N_19439,N_19176);
and U23376 (N_23376,N_16282,N_19503);
nor U23377 (N_23377,N_18164,N_18644);
and U23378 (N_23378,N_18221,N_17182);
nor U23379 (N_23379,N_19449,N_18896);
and U23380 (N_23380,N_15754,N_17800);
nor U23381 (N_23381,N_17394,N_19677);
nand U23382 (N_23382,N_19169,N_16958);
nand U23383 (N_23383,N_15694,N_17565);
and U23384 (N_23384,N_16629,N_19546);
and U23385 (N_23385,N_15155,N_18005);
nand U23386 (N_23386,N_16341,N_16919);
xnor U23387 (N_23387,N_17334,N_17558);
nor U23388 (N_23388,N_18394,N_15096);
or U23389 (N_23389,N_18861,N_17539);
and U23390 (N_23390,N_18407,N_17859);
nand U23391 (N_23391,N_15716,N_15649);
or U23392 (N_23392,N_16531,N_19109);
nand U23393 (N_23393,N_19830,N_17388);
and U23394 (N_23394,N_15005,N_15953);
or U23395 (N_23395,N_18039,N_15831);
or U23396 (N_23396,N_19627,N_18937);
and U23397 (N_23397,N_19328,N_16719);
nand U23398 (N_23398,N_17408,N_15822);
and U23399 (N_23399,N_16594,N_15752);
xnor U23400 (N_23400,N_17065,N_17020);
nor U23401 (N_23401,N_17791,N_15044);
nor U23402 (N_23402,N_15741,N_15291);
nand U23403 (N_23403,N_15502,N_15767);
or U23404 (N_23404,N_17083,N_18880);
or U23405 (N_23405,N_17875,N_19884);
xnor U23406 (N_23406,N_15097,N_19814);
nand U23407 (N_23407,N_16557,N_19029);
nand U23408 (N_23408,N_16013,N_16980);
nor U23409 (N_23409,N_17035,N_17363);
or U23410 (N_23410,N_16501,N_16789);
nor U23411 (N_23411,N_15054,N_18545);
and U23412 (N_23412,N_19266,N_18143);
and U23413 (N_23413,N_18259,N_17541);
or U23414 (N_23414,N_17220,N_18705);
or U23415 (N_23415,N_18404,N_16687);
nor U23416 (N_23416,N_16496,N_17691);
or U23417 (N_23417,N_15970,N_17061);
nand U23418 (N_23418,N_19069,N_17665);
nor U23419 (N_23419,N_18267,N_16776);
or U23420 (N_23420,N_16807,N_19594);
nand U23421 (N_23421,N_15590,N_17193);
or U23422 (N_23422,N_17377,N_17810);
and U23423 (N_23423,N_15210,N_16307);
or U23424 (N_23424,N_17714,N_15340);
or U23425 (N_23425,N_18814,N_17890);
xor U23426 (N_23426,N_18342,N_16090);
nor U23427 (N_23427,N_18236,N_19283);
xnor U23428 (N_23428,N_16338,N_16164);
nor U23429 (N_23429,N_19414,N_18332);
nor U23430 (N_23430,N_17474,N_19831);
nor U23431 (N_23431,N_15475,N_17314);
nand U23432 (N_23432,N_16001,N_16380);
and U23433 (N_23433,N_17065,N_15133);
and U23434 (N_23434,N_17221,N_15355);
xnor U23435 (N_23435,N_17834,N_16658);
nor U23436 (N_23436,N_15806,N_18119);
nand U23437 (N_23437,N_15719,N_16719);
xnor U23438 (N_23438,N_16334,N_19568);
nand U23439 (N_23439,N_16550,N_17563);
nor U23440 (N_23440,N_17758,N_18767);
nor U23441 (N_23441,N_19990,N_18810);
nand U23442 (N_23442,N_19949,N_19883);
nand U23443 (N_23443,N_19507,N_16775);
nand U23444 (N_23444,N_16100,N_15160);
nand U23445 (N_23445,N_17803,N_19348);
nand U23446 (N_23446,N_15653,N_15342);
and U23447 (N_23447,N_15778,N_19270);
nand U23448 (N_23448,N_17792,N_15609);
nor U23449 (N_23449,N_19851,N_17832);
xor U23450 (N_23450,N_19683,N_19425);
and U23451 (N_23451,N_19793,N_16494);
nand U23452 (N_23452,N_17784,N_16787);
and U23453 (N_23453,N_19845,N_15644);
xor U23454 (N_23454,N_15334,N_18507);
nand U23455 (N_23455,N_19226,N_16805);
nand U23456 (N_23456,N_19494,N_19961);
nor U23457 (N_23457,N_15085,N_17402);
nor U23458 (N_23458,N_16467,N_15082);
nor U23459 (N_23459,N_19884,N_15908);
nand U23460 (N_23460,N_19729,N_18163);
nor U23461 (N_23461,N_19717,N_15063);
nor U23462 (N_23462,N_19716,N_19910);
or U23463 (N_23463,N_18246,N_17425);
nor U23464 (N_23464,N_15944,N_15084);
or U23465 (N_23465,N_17435,N_19030);
nand U23466 (N_23466,N_15638,N_19384);
nor U23467 (N_23467,N_16835,N_16482);
nor U23468 (N_23468,N_16681,N_15240);
nor U23469 (N_23469,N_15265,N_16299);
or U23470 (N_23470,N_16484,N_16199);
or U23471 (N_23471,N_18388,N_15319);
or U23472 (N_23472,N_18653,N_17161);
nand U23473 (N_23473,N_15851,N_17532);
nor U23474 (N_23474,N_19426,N_16211);
or U23475 (N_23475,N_17625,N_18618);
and U23476 (N_23476,N_17245,N_15690);
nor U23477 (N_23477,N_17677,N_19501);
nor U23478 (N_23478,N_16699,N_18820);
xor U23479 (N_23479,N_17317,N_18248);
nand U23480 (N_23480,N_19237,N_15497);
xnor U23481 (N_23481,N_16327,N_17805);
nand U23482 (N_23482,N_15102,N_15228);
and U23483 (N_23483,N_18096,N_15978);
or U23484 (N_23484,N_15914,N_19546);
nor U23485 (N_23485,N_17778,N_19258);
and U23486 (N_23486,N_15745,N_18042);
or U23487 (N_23487,N_15076,N_17113);
or U23488 (N_23488,N_18919,N_15219);
xor U23489 (N_23489,N_16230,N_19545);
xor U23490 (N_23490,N_19425,N_16004);
nor U23491 (N_23491,N_18206,N_19365);
nor U23492 (N_23492,N_19392,N_19428);
nand U23493 (N_23493,N_15883,N_19821);
nand U23494 (N_23494,N_18684,N_17591);
xnor U23495 (N_23495,N_19963,N_16057);
nor U23496 (N_23496,N_19275,N_15101);
nor U23497 (N_23497,N_18228,N_19235);
nand U23498 (N_23498,N_15985,N_18098);
nor U23499 (N_23499,N_15439,N_15076);
xor U23500 (N_23500,N_17963,N_18823);
and U23501 (N_23501,N_18771,N_17749);
or U23502 (N_23502,N_19809,N_18602);
or U23503 (N_23503,N_17637,N_18522);
or U23504 (N_23504,N_19328,N_19707);
or U23505 (N_23505,N_16010,N_16504);
nand U23506 (N_23506,N_18535,N_19339);
xnor U23507 (N_23507,N_15886,N_15668);
or U23508 (N_23508,N_15820,N_18924);
nand U23509 (N_23509,N_16446,N_19423);
and U23510 (N_23510,N_18269,N_19608);
or U23511 (N_23511,N_17984,N_17472);
or U23512 (N_23512,N_16439,N_17292);
xnor U23513 (N_23513,N_18024,N_15863);
and U23514 (N_23514,N_16131,N_19691);
nor U23515 (N_23515,N_16435,N_16188);
nand U23516 (N_23516,N_16427,N_18213);
nand U23517 (N_23517,N_15122,N_15108);
nand U23518 (N_23518,N_18795,N_16678);
xnor U23519 (N_23519,N_17450,N_16184);
or U23520 (N_23520,N_17306,N_16526);
xnor U23521 (N_23521,N_17571,N_18189);
or U23522 (N_23522,N_15265,N_17344);
or U23523 (N_23523,N_15513,N_16970);
nand U23524 (N_23524,N_18400,N_16250);
nand U23525 (N_23525,N_18428,N_19267);
nor U23526 (N_23526,N_19491,N_17231);
and U23527 (N_23527,N_17972,N_18210);
nor U23528 (N_23528,N_15606,N_15148);
nor U23529 (N_23529,N_18045,N_19792);
and U23530 (N_23530,N_17054,N_17947);
and U23531 (N_23531,N_17472,N_16151);
or U23532 (N_23532,N_18576,N_17981);
xor U23533 (N_23533,N_17890,N_16959);
and U23534 (N_23534,N_18739,N_18627);
and U23535 (N_23535,N_18955,N_16274);
nand U23536 (N_23536,N_15172,N_15553);
xor U23537 (N_23537,N_16867,N_16436);
xor U23538 (N_23538,N_17564,N_17035);
and U23539 (N_23539,N_15138,N_15425);
nor U23540 (N_23540,N_16390,N_18532);
nand U23541 (N_23541,N_17593,N_17864);
xor U23542 (N_23542,N_17485,N_16464);
nand U23543 (N_23543,N_16745,N_18304);
and U23544 (N_23544,N_19986,N_19050);
nor U23545 (N_23545,N_19072,N_16076);
nor U23546 (N_23546,N_19229,N_19749);
and U23547 (N_23547,N_16449,N_17800);
xnor U23548 (N_23548,N_16875,N_15886);
and U23549 (N_23549,N_19075,N_19372);
nand U23550 (N_23550,N_16012,N_18148);
nand U23551 (N_23551,N_15036,N_17009);
or U23552 (N_23552,N_15843,N_17766);
and U23553 (N_23553,N_19802,N_16582);
xnor U23554 (N_23554,N_19001,N_19730);
xor U23555 (N_23555,N_18018,N_19084);
xnor U23556 (N_23556,N_18427,N_19406);
xnor U23557 (N_23557,N_16897,N_19879);
or U23558 (N_23558,N_15412,N_19152);
or U23559 (N_23559,N_18272,N_18900);
nand U23560 (N_23560,N_15439,N_17693);
and U23561 (N_23561,N_18549,N_18072);
nor U23562 (N_23562,N_15490,N_19696);
and U23563 (N_23563,N_17550,N_18768);
nand U23564 (N_23564,N_16395,N_16861);
xor U23565 (N_23565,N_17806,N_19240);
nor U23566 (N_23566,N_17198,N_17855);
nor U23567 (N_23567,N_17686,N_15056);
nor U23568 (N_23568,N_19386,N_19825);
and U23569 (N_23569,N_16277,N_17780);
nand U23570 (N_23570,N_16785,N_18968);
nor U23571 (N_23571,N_19282,N_17242);
or U23572 (N_23572,N_18833,N_19790);
nand U23573 (N_23573,N_19836,N_19853);
and U23574 (N_23574,N_19723,N_17967);
xor U23575 (N_23575,N_19062,N_19501);
xor U23576 (N_23576,N_18732,N_15892);
and U23577 (N_23577,N_18075,N_19102);
nand U23578 (N_23578,N_15912,N_16017);
xnor U23579 (N_23579,N_15409,N_17763);
and U23580 (N_23580,N_18069,N_17782);
and U23581 (N_23581,N_16210,N_19371);
nor U23582 (N_23582,N_16778,N_15221);
nor U23583 (N_23583,N_16339,N_19405);
nor U23584 (N_23584,N_19469,N_19097);
nor U23585 (N_23585,N_19073,N_18208);
xor U23586 (N_23586,N_17951,N_18251);
nor U23587 (N_23587,N_19153,N_15088);
nand U23588 (N_23588,N_15860,N_19228);
and U23589 (N_23589,N_18814,N_16998);
or U23590 (N_23590,N_18657,N_17312);
xor U23591 (N_23591,N_16135,N_15227);
or U23592 (N_23592,N_15126,N_17043);
nand U23593 (N_23593,N_17823,N_17768);
nor U23594 (N_23594,N_17027,N_19349);
or U23595 (N_23595,N_17758,N_15220);
or U23596 (N_23596,N_19453,N_16937);
xnor U23597 (N_23597,N_17183,N_17244);
and U23598 (N_23598,N_19389,N_16229);
xnor U23599 (N_23599,N_15483,N_16148);
or U23600 (N_23600,N_15144,N_16465);
nand U23601 (N_23601,N_17205,N_15580);
or U23602 (N_23602,N_17199,N_17732);
nor U23603 (N_23603,N_15394,N_15734);
and U23604 (N_23604,N_16541,N_15928);
or U23605 (N_23605,N_19827,N_18356);
or U23606 (N_23606,N_17197,N_18729);
xnor U23607 (N_23607,N_16952,N_16406);
and U23608 (N_23608,N_15272,N_18150);
xor U23609 (N_23609,N_18733,N_17138);
or U23610 (N_23610,N_17374,N_16315);
nor U23611 (N_23611,N_15415,N_16577);
and U23612 (N_23612,N_17543,N_15326);
or U23613 (N_23613,N_18104,N_15816);
xor U23614 (N_23614,N_16215,N_18405);
or U23615 (N_23615,N_15184,N_18839);
or U23616 (N_23616,N_16569,N_17908);
and U23617 (N_23617,N_15673,N_19547);
nand U23618 (N_23618,N_17265,N_16030);
nand U23619 (N_23619,N_16528,N_16150);
xnor U23620 (N_23620,N_16040,N_17033);
nand U23621 (N_23621,N_19333,N_15702);
xor U23622 (N_23622,N_15637,N_17923);
or U23623 (N_23623,N_18898,N_15994);
or U23624 (N_23624,N_15238,N_17842);
xor U23625 (N_23625,N_19810,N_18094);
or U23626 (N_23626,N_18696,N_16011);
or U23627 (N_23627,N_19417,N_15354);
and U23628 (N_23628,N_15684,N_15963);
xnor U23629 (N_23629,N_19040,N_19652);
and U23630 (N_23630,N_16969,N_19188);
nor U23631 (N_23631,N_15959,N_17507);
and U23632 (N_23632,N_16889,N_16405);
xor U23633 (N_23633,N_15536,N_16081);
and U23634 (N_23634,N_17087,N_17532);
nand U23635 (N_23635,N_18659,N_18359);
xnor U23636 (N_23636,N_18646,N_16215);
nor U23637 (N_23637,N_18750,N_16999);
and U23638 (N_23638,N_17090,N_16917);
and U23639 (N_23639,N_15896,N_15833);
nor U23640 (N_23640,N_18156,N_18740);
xnor U23641 (N_23641,N_15792,N_19634);
xnor U23642 (N_23642,N_19247,N_18702);
nor U23643 (N_23643,N_15767,N_16366);
nor U23644 (N_23644,N_16102,N_17836);
nor U23645 (N_23645,N_16628,N_19250);
nor U23646 (N_23646,N_15738,N_18355);
nor U23647 (N_23647,N_17827,N_16382);
nand U23648 (N_23648,N_15731,N_18384);
xor U23649 (N_23649,N_15168,N_15787);
nand U23650 (N_23650,N_18124,N_19605);
nor U23651 (N_23651,N_19171,N_16974);
nor U23652 (N_23652,N_19564,N_17970);
xor U23653 (N_23653,N_17853,N_15834);
or U23654 (N_23654,N_18303,N_18420);
nor U23655 (N_23655,N_18514,N_18486);
or U23656 (N_23656,N_16572,N_19451);
and U23657 (N_23657,N_17597,N_19282);
nand U23658 (N_23658,N_15113,N_15537);
and U23659 (N_23659,N_19878,N_16085);
and U23660 (N_23660,N_16949,N_15091);
and U23661 (N_23661,N_16196,N_16487);
nand U23662 (N_23662,N_18414,N_18326);
nor U23663 (N_23663,N_19347,N_18996);
or U23664 (N_23664,N_18750,N_16480);
nand U23665 (N_23665,N_16387,N_15589);
or U23666 (N_23666,N_15867,N_19175);
nand U23667 (N_23667,N_19969,N_15931);
nor U23668 (N_23668,N_15938,N_18590);
nand U23669 (N_23669,N_19998,N_17399);
xnor U23670 (N_23670,N_19118,N_18384);
xor U23671 (N_23671,N_18975,N_15994);
nand U23672 (N_23672,N_17102,N_19183);
nand U23673 (N_23673,N_17957,N_16427);
nor U23674 (N_23674,N_19071,N_19113);
and U23675 (N_23675,N_16707,N_18988);
and U23676 (N_23676,N_17123,N_19134);
or U23677 (N_23677,N_19321,N_17466);
nand U23678 (N_23678,N_15914,N_16108);
and U23679 (N_23679,N_15718,N_16132);
and U23680 (N_23680,N_16784,N_18705);
xor U23681 (N_23681,N_15022,N_18582);
xor U23682 (N_23682,N_19531,N_17581);
or U23683 (N_23683,N_19347,N_19441);
and U23684 (N_23684,N_16776,N_18303);
nand U23685 (N_23685,N_19152,N_15998);
xnor U23686 (N_23686,N_19263,N_19493);
nor U23687 (N_23687,N_17934,N_19007);
xor U23688 (N_23688,N_19023,N_17464);
or U23689 (N_23689,N_19182,N_19071);
and U23690 (N_23690,N_19899,N_19939);
xnor U23691 (N_23691,N_17554,N_16967);
or U23692 (N_23692,N_18982,N_17080);
nand U23693 (N_23693,N_16676,N_18788);
or U23694 (N_23694,N_18454,N_18867);
xor U23695 (N_23695,N_16117,N_15433);
nor U23696 (N_23696,N_16773,N_19430);
and U23697 (N_23697,N_17367,N_16799);
nand U23698 (N_23698,N_18573,N_17576);
and U23699 (N_23699,N_19460,N_17136);
nand U23700 (N_23700,N_15483,N_19819);
or U23701 (N_23701,N_17765,N_15529);
or U23702 (N_23702,N_19466,N_19294);
nand U23703 (N_23703,N_15241,N_15322);
xor U23704 (N_23704,N_18904,N_18518);
or U23705 (N_23705,N_16668,N_16426);
xnor U23706 (N_23706,N_19587,N_15418);
or U23707 (N_23707,N_16281,N_16667);
nor U23708 (N_23708,N_15833,N_15657);
or U23709 (N_23709,N_18371,N_15894);
nand U23710 (N_23710,N_16553,N_15067);
xnor U23711 (N_23711,N_19102,N_15201);
nor U23712 (N_23712,N_17159,N_15343);
nor U23713 (N_23713,N_15350,N_18759);
nand U23714 (N_23714,N_16778,N_19674);
xor U23715 (N_23715,N_19462,N_19022);
xor U23716 (N_23716,N_17819,N_16067);
nor U23717 (N_23717,N_16030,N_18182);
or U23718 (N_23718,N_15068,N_19197);
and U23719 (N_23719,N_18932,N_17309);
xor U23720 (N_23720,N_17321,N_17972);
or U23721 (N_23721,N_15730,N_17625);
xor U23722 (N_23722,N_19505,N_19985);
nand U23723 (N_23723,N_16186,N_19462);
nand U23724 (N_23724,N_16437,N_18747);
nand U23725 (N_23725,N_19904,N_17790);
and U23726 (N_23726,N_16127,N_15220);
nand U23727 (N_23727,N_16152,N_16455);
xnor U23728 (N_23728,N_16350,N_19938);
and U23729 (N_23729,N_18202,N_15666);
nor U23730 (N_23730,N_18882,N_17581);
nand U23731 (N_23731,N_18742,N_19071);
nor U23732 (N_23732,N_18074,N_17358);
or U23733 (N_23733,N_16065,N_17512);
or U23734 (N_23734,N_15437,N_18382);
or U23735 (N_23735,N_19528,N_19654);
nand U23736 (N_23736,N_18955,N_19167);
or U23737 (N_23737,N_16764,N_15833);
nand U23738 (N_23738,N_18684,N_17740);
nand U23739 (N_23739,N_16660,N_18642);
and U23740 (N_23740,N_19001,N_16916);
or U23741 (N_23741,N_16460,N_17911);
and U23742 (N_23742,N_16026,N_17621);
nand U23743 (N_23743,N_15458,N_15736);
nor U23744 (N_23744,N_19084,N_15111);
and U23745 (N_23745,N_17409,N_15806);
and U23746 (N_23746,N_18611,N_16001);
nor U23747 (N_23747,N_15852,N_19070);
nand U23748 (N_23748,N_16525,N_19190);
or U23749 (N_23749,N_17868,N_19126);
or U23750 (N_23750,N_18881,N_15755);
and U23751 (N_23751,N_18922,N_17262);
xor U23752 (N_23752,N_18348,N_16825);
xnor U23753 (N_23753,N_15717,N_16636);
nor U23754 (N_23754,N_19395,N_19233);
nor U23755 (N_23755,N_15689,N_16111);
xnor U23756 (N_23756,N_18516,N_18477);
or U23757 (N_23757,N_17766,N_17647);
or U23758 (N_23758,N_15366,N_16635);
nor U23759 (N_23759,N_18639,N_19461);
and U23760 (N_23760,N_16104,N_18641);
nor U23761 (N_23761,N_19000,N_18429);
or U23762 (N_23762,N_15184,N_18663);
nand U23763 (N_23763,N_19720,N_15637);
and U23764 (N_23764,N_19553,N_16221);
nand U23765 (N_23765,N_18992,N_15346);
nor U23766 (N_23766,N_18652,N_15279);
xor U23767 (N_23767,N_15549,N_15507);
xnor U23768 (N_23768,N_17175,N_17753);
xor U23769 (N_23769,N_17957,N_19149);
or U23770 (N_23770,N_19232,N_16858);
nor U23771 (N_23771,N_17754,N_18715);
xor U23772 (N_23772,N_19837,N_15762);
nand U23773 (N_23773,N_18381,N_16658);
or U23774 (N_23774,N_18251,N_18901);
and U23775 (N_23775,N_16892,N_16160);
nand U23776 (N_23776,N_17179,N_17459);
and U23777 (N_23777,N_16071,N_17594);
nand U23778 (N_23778,N_19220,N_15244);
nand U23779 (N_23779,N_17682,N_19218);
and U23780 (N_23780,N_16259,N_15435);
or U23781 (N_23781,N_15022,N_16942);
nand U23782 (N_23782,N_17554,N_16882);
or U23783 (N_23783,N_17128,N_16480);
or U23784 (N_23784,N_19382,N_19050);
and U23785 (N_23785,N_18053,N_15996);
nor U23786 (N_23786,N_19020,N_19817);
xnor U23787 (N_23787,N_18463,N_15824);
xor U23788 (N_23788,N_19864,N_16690);
or U23789 (N_23789,N_17561,N_19089);
nor U23790 (N_23790,N_17357,N_16534);
nand U23791 (N_23791,N_16224,N_18617);
nand U23792 (N_23792,N_16958,N_18971);
and U23793 (N_23793,N_15072,N_15723);
xnor U23794 (N_23794,N_18370,N_17197);
or U23795 (N_23795,N_17327,N_15991);
nand U23796 (N_23796,N_17496,N_18260);
xor U23797 (N_23797,N_17899,N_16889);
nand U23798 (N_23798,N_15438,N_19835);
xnor U23799 (N_23799,N_19757,N_16548);
nor U23800 (N_23800,N_15351,N_15649);
or U23801 (N_23801,N_19699,N_15407);
nor U23802 (N_23802,N_15437,N_15094);
nand U23803 (N_23803,N_16713,N_16376);
or U23804 (N_23804,N_19587,N_19287);
nor U23805 (N_23805,N_18923,N_18617);
xnor U23806 (N_23806,N_18629,N_15844);
or U23807 (N_23807,N_17758,N_19799);
nand U23808 (N_23808,N_16002,N_17469);
xor U23809 (N_23809,N_18996,N_16382);
xor U23810 (N_23810,N_18350,N_16597);
and U23811 (N_23811,N_19430,N_18694);
xnor U23812 (N_23812,N_17084,N_15630);
and U23813 (N_23813,N_17375,N_19418);
nor U23814 (N_23814,N_16046,N_18872);
nor U23815 (N_23815,N_16945,N_15890);
or U23816 (N_23816,N_18110,N_15815);
or U23817 (N_23817,N_17446,N_19784);
nor U23818 (N_23818,N_15800,N_17031);
nor U23819 (N_23819,N_15036,N_15444);
nor U23820 (N_23820,N_15711,N_19172);
nand U23821 (N_23821,N_19546,N_15930);
nand U23822 (N_23822,N_17253,N_15662);
nor U23823 (N_23823,N_19109,N_17362);
nor U23824 (N_23824,N_17100,N_17354);
nor U23825 (N_23825,N_19893,N_18125);
nand U23826 (N_23826,N_17200,N_19764);
and U23827 (N_23827,N_19557,N_17629);
or U23828 (N_23828,N_18635,N_17673);
nor U23829 (N_23829,N_16970,N_15782);
or U23830 (N_23830,N_17054,N_17344);
nor U23831 (N_23831,N_16365,N_17042);
or U23832 (N_23832,N_15764,N_15374);
xnor U23833 (N_23833,N_17886,N_18007);
nand U23834 (N_23834,N_19201,N_15132);
xor U23835 (N_23835,N_17388,N_19593);
and U23836 (N_23836,N_19322,N_16301);
and U23837 (N_23837,N_19624,N_16991);
nor U23838 (N_23838,N_16572,N_15475);
or U23839 (N_23839,N_19055,N_16990);
nand U23840 (N_23840,N_17757,N_17107);
or U23841 (N_23841,N_17033,N_17309);
nor U23842 (N_23842,N_18382,N_15609);
xnor U23843 (N_23843,N_16004,N_19060);
nand U23844 (N_23844,N_16805,N_16422);
or U23845 (N_23845,N_15824,N_17607);
nand U23846 (N_23846,N_19111,N_18026);
nand U23847 (N_23847,N_17506,N_15467);
or U23848 (N_23848,N_15788,N_19265);
xor U23849 (N_23849,N_18971,N_18886);
nor U23850 (N_23850,N_17918,N_17861);
or U23851 (N_23851,N_19388,N_17176);
and U23852 (N_23852,N_18586,N_16826);
nand U23853 (N_23853,N_19018,N_17634);
xnor U23854 (N_23854,N_19172,N_18340);
nand U23855 (N_23855,N_15201,N_17097);
and U23856 (N_23856,N_19878,N_19947);
xnor U23857 (N_23857,N_16538,N_19651);
and U23858 (N_23858,N_15307,N_15561);
nor U23859 (N_23859,N_16627,N_15396);
nand U23860 (N_23860,N_17914,N_16574);
and U23861 (N_23861,N_17615,N_16383);
nand U23862 (N_23862,N_18620,N_19006);
or U23863 (N_23863,N_17373,N_16520);
nor U23864 (N_23864,N_19383,N_16596);
nand U23865 (N_23865,N_18444,N_16514);
or U23866 (N_23866,N_15755,N_15463);
nor U23867 (N_23867,N_18886,N_17715);
nand U23868 (N_23868,N_16379,N_18829);
xor U23869 (N_23869,N_19134,N_15853);
or U23870 (N_23870,N_16655,N_18307);
nand U23871 (N_23871,N_18065,N_17337);
and U23872 (N_23872,N_16810,N_19326);
xor U23873 (N_23873,N_17925,N_17097);
xor U23874 (N_23874,N_17384,N_18389);
nand U23875 (N_23875,N_19839,N_19362);
or U23876 (N_23876,N_19264,N_18864);
nand U23877 (N_23877,N_19047,N_17040);
xnor U23878 (N_23878,N_15726,N_17273);
nor U23879 (N_23879,N_17362,N_19463);
nand U23880 (N_23880,N_17804,N_16011);
nor U23881 (N_23881,N_15759,N_19353);
and U23882 (N_23882,N_17898,N_19679);
nor U23883 (N_23883,N_18218,N_18874);
xor U23884 (N_23884,N_17626,N_17522);
nand U23885 (N_23885,N_16499,N_19600);
and U23886 (N_23886,N_16953,N_19864);
and U23887 (N_23887,N_15048,N_16716);
nor U23888 (N_23888,N_16474,N_16992);
nor U23889 (N_23889,N_15486,N_19033);
xor U23890 (N_23890,N_17084,N_18386);
and U23891 (N_23891,N_17141,N_15408);
xor U23892 (N_23892,N_16545,N_15687);
and U23893 (N_23893,N_16354,N_19809);
or U23894 (N_23894,N_18897,N_16799);
nand U23895 (N_23895,N_19856,N_15446);
nand U23896 (N_23896,N_18629,N_17457);
or U23897 (N_23897,N_19655,N_18940);
xor U23898 (N_23898,N_15366,N_16418);
and U23899 (N_23899,N_15192,N_16296);
nand U23900 (N_23900,N_16224,N_15791);
or U23901 (N_23901,N_16445,N_15602);
and U23902 (N_23902,N_15055,N_18876);
xor U23903 (N_23903,N_18884,N_15500);
nand U23904 (N_23904,N_19258,N_19367);
xnor U23905 (N_23905,N_17293,N_16637);
nor U23906 (N_23906,N_17559,N_15515);
xor U23907 (N_23907,N_19094,N_15092);
or U23908 (N_23908,N_17021,N_17497);
xnor U23909 (N_23909,N_16656,N_17992);
nand U23910 (N_23910,N_18849,N_15868);
or U23911 (N_23911,N_19348,N_17281);
or U23912 (N_23912,N_16715,N_15036);
nor U23913 (N_23913,N_18131,N_17898);
nand U23914 (N_23914,N_17155,N_17801);
nand U23915 (N_23915,N_16799,N_18164);
nor U23916 (N_23916,N_18560,N_17823);
xor U23917 (N_23917,N_19245,N_18144);
nand U23918 (N_23918,N_15716,N_18830);
nor U23919 (N_23919,N_16014,N_19410);
nor U23920 (N_23920,N_16886,N_17991);
or U23921 (N_23921,N_16663,N_17339);
nor U23922 (N_23922,N_18132,N_15353);
xor U23923 (N_23923,N_19746,N_17432);
or U23924 (N_23924,N_19090,N_19599);
nand U23925 (N_23925,N_15209,N_15591);
and U23926 (N_23926,N_19544,N_18665);
nor U23927 (N_23927,N_19756,N_15055);
xnor U23928 (N_23928,N_17632,N_15196);
or U23929 (N_23929,N_19685,N_17526);
nand U23930 (N_23930,N_18254,N_18054);
xor U23931 (N_23931,N_17057,N_18405);
and U23932 (N_23932,N_18499,N_15430);
or U23933 (N_23933,N_15893,N_19931);
xnor U23934 (N_23934,N_16264,N_16121);
and U23935 (N_23935,N_16803,N_19641);
nor U23936 (N_23936,N_17693,N_19629);
nor U23937 (N_23937,N_16817,N_16807);
and U23938 (N_23938,N_17578,N_19928);
and U23939 (N_23939,N_17734,N_17031);
nor U23940 (N_23940,N_17494,N_16336);
nor U23941 (N_23941,N_19257,N_15418);
nand U23942 (N_23942,N_19772,N_19633);
nor U23943 (N_23943,N_17521,N_16691);
nor U23944 (N_23944,N_16088,N_15989);
and U23945 (N_23945,N_16658,N_17298);
nand U23946 (N_23946,N_19325,N_18446);
and U23947 (N_23947,N_16065,N_16132);
xnor U23948 (N_23948,N_18369,N_16312);
or U23949 (N_23949,N_19113,N_15851);
xnor U23950 (N_23950,N_16378,N_17394);
nand U23951 (N_23951,N_17590,N_15859);
and U23952 (N_23952,N_16042,N_16821);
nor U23953 (N_23953,N_18835,N_18345);
or U23954 (N_23954,N_18831,N_19762);
or U23955 (N_23955,N_16838,N_17875);
or U23956 (N_23956,N_19067,N_15831);
or U23957 (N_23957,N_16017,N_15961);
nand U23958 (N_23958,N_17010,N_19414);
nor U23959 (N_23959,N_16667,N_15402);
xnor U23960 (N_23960,N_16358,N_17560);
xnor U23961 (N_23961,N_18315,N_16620);
or U23962 (N_23962,N_15558,N_16932);
or U23963 (N_23963,N_17175,N_18822);
or U23964 (N_23964,N_15630,N_19403);
xor U23965 (N_23965,N_15762,N_15498);
nand U23966 (N_23966,N_17665,N_15494);
nor U23967 (N_23967,N_18832,N_15094);
nor U23968 (N_23968,N_17985,N_15323);
and U23969 (N_23969,N_19462,N_18066);
or U23970 (N_23970,N_19036,N_16592);
nand U23971 (N_23971,N_15093,N_17803);
nor U23972 (N_23972,N_16181,N_17876);
nand U23973 (N_23973,N_16297,N_16222);
and U23974 (N_23974,N_18892,N_17723);
nand U23975 (N_23975,N_19179,N_18080);
and U23976 (N_23976,N_19968,N_18531);
xnor U23977 (N_23977,N_16025,N_18333);
or U23978 (N_23978,N_15571,N_18833);
nor U23979 (N_23979,N_19805,N_18305);
xor U23980 (N_23980,N_16835,N_17127);
and U23981 (N_23981,N_19714,N_18915);
nor U23982 (N_23982,N_15768,N_18329);
or U23983 (N_23983,N_15608,N_17390);
nor U23984 (N_23984,N_16643,N_17719);
xnor U23985 (N_23985,N_16819,N_18570);
or U23986 (N_23986,N_15188,N_19764);
nor U23987 (N_23987,N_19191,N_18626);
nor U23988 (N_23988,N_18625,N_17716);
xor U23989 (N_23989,N_18288,N_18512);
nor U23990 (N_23990,N_16951,N_18652);
and U23991 (N_23991,N_17165,N_19701);
xor U23992 (N_23992,N_16865,N_17229);
nand U23993 (N_23993,N_17421,N_16473);
nor U23994 (N_23994,N_15012,N_18572);
xnor U23995 (N_23995,N_15987,N_15851);
nand U23996 (N_23996,N_19922,N_18305);
nor U23997 (N_23997,N_16581,N_18499);
or U23998 (N_23998,N_16799,N_15884);
and U23999 (N_23999,N_15020,N_18048);
nor U24000 (N_24000,N_19736,N_18916);
and U24001 (N_24001,N_18913,N_19467);
or U24002 (N_24002,N_17323,N_18773);
or U24003 (N_24003,N_16021,N_15824);
or U24004 (N_24004,N_18126,N_17082);
nor U24005 (N_24005,N_19387,N_15249);
nor U24006 (N_24006,N_17175,N_16561);
xnor U24007 (N_24007,N_17664,N_18083);
or U24008 (N_24008,N_17485,N_16738);
nand U24009 (N_24009,N_18759,N_15729);
nor U24010 (N_24010,N_18904,N_15321);
and U24011 (N_24011,N_16863,N_15997);
nand U24012 (N_24012,N_19771,N_16587);
and U24013 (N_24013,N_19501,N_18519);
nor U24014 (N_24014,N_15390,N_15503);
xor U24015 (N_24015,N_18196,N_19266);
xor U24016 (N_24016,N_18846,N_17045);
and U24017 (N_24017,N_15043,N_17682);
and U24018 (N_24018,N_17360,N_19810);
or U24019 (N_24019,N_15166,N_17814);
and U24020 (N_24020,N_18629,N_16266);
nor U24021 (N_24021,N_15570,N_19961);
or U24022 (N_24022,N_15326,N_15147);
xnor U24023 (N_24023,N_19102,N_18882);
xor U24024 (N_24024,N_17445,N_19633);
nor U24025 (N_24025,N_19282,N_17668);
nand U24026 (N_24026,N_17809,N_17610);
nand U24027 (N_24027,N_16842,N_17470);
nand U24028 (N_24028,N_18369,N_18118);
nand U24029 (N_24029,N_18323,N_17811);
nor U24030 (N_24030,N_17113,N_19824);
and U24031 (N_24031,N_16326,N_19668);
nand U24032 (N_24032,N_15923,N_15264);
nor U24033 (N_24033,N_16958,N_19439);
and U24034 (N_24034,N_16801,N_19897);
or U24035 (N_24035,N_17176,N_19151);
xor U24036 (N_24036,N_16827,N_15112);
or U24037 (N_24037,N_16696,N_15569);
nand U24038 (N_24038,N_15123,N_16245);
nor U24039 (N_24039,N_15773,N_16699);
and U24040 (N_24040,N_18111,N_15710);
nor U24041 (N_24041,N_18037,N_17393);
and U24042 (N_24042,N_19456,N_19834);
nand U24043 (N_24043,N_18655,N_15216);
and U24044 (N_24044,N_15194,N_17956);
and U24045 (N_24045,N_15772,N_18674);
xor U24046 (N_24046,N_19651,N_15630);
xor U24047 (N_24047,N_17951,N_16115);
xnor U24048 (N_24048,N_19509,N_15667);
xnor U24049 (N_24049,N_19795,N_19407);
and U24050 (N_24050,N_15446,N_19020);
xor U24051 (N_24051,N_19931,N_17421);
xor U24052 (N_24052,N_16613,N_15322);
xnor U24053 (N_24053,N_15651,N_15099);
and U24054 (N_24054,N_18784,N_17322);
xor U24055 (N_24055,N_16792,N_16108);
nand U24056 (N_24056,N_19900,N_18029);
xor U24057 (N_24057,N_18080,N_19044);
nand U24058 (N_24058,N_17168,N_15620);
nor U24059 (N_24059,N_15465,N_17393);
nor U24060 (N_24060,N_19616,N_16946);
and U24061 (N_24061,N_15739,N_17504);
xnor U24062 (N_24062,N_16894,N_18120);
or U24063 (N_24063,N_19053,N_18681);
nor U24064 (N_24064,N_18598,N_19064);
or U24065 (N_24065,N_17836,N_17425);
or U24066 (N_24066,N_15757,N_15493);
nand U24067 (N_24067,N_19967,N_17161);
nor U24068 (N_24068,N_16884,N_19883);
and U24069 (N_24069,N_18370,N_15442);
and U24070 (N_24070,N_15512,N_15332);
or U24071 (N_24071,N_15987,N_17317);
or U24072 (N_24072,N_16448,N_18905);
nand U24073 (N_24073,N_15967,N_19036);
or U24074 (N_24074,N_19916,N_15883);
xnor U24075 (N_24075,N_15802,N_16136);
nor U24076 (N_24076,N_16534,N_17448);
and U24077 (N_24077,N_19987,N_16359);
nor U24078 (N_24078,N_16642,N_15327);
xnor U24079 (N_24079,N_15784,N_16792);
and U24080 (N_24080,N_17960,N_19115);
nor U24081 (N_24081,N_18335,N_16848);
or U24082 (N_24082,N_18290,N_17033);
and U24083 (N_24083,N_15250,N_15180);
or U24084 (N_24084,N_16865,N_18439);
or U24085 (N_24085,N_18487,N_16891);
nor U24086 (N_24086,N_18838,N_16364);
nand U24087 (N_24087,N_15711,N_17701);
and U24088 (N_24088,N_16960,N_16016);
and U24089 (N_24089,N_17164,N_15463);
nor U24090 (N_24090,N_18113,N_19222);
or U24091 (N_24091,N_15689,N_19066);
and U24092 (N_24092,N_17558,N_17026);
xor U24093 (N_24093,N_18607,N_18302);
nand U24094 (N_24094,N_16095,N_17020);
nand U24095 (N_24095,N_16483,N_19206);
xor U24096 (N_24096,N_17542,N_17698);
nor U24097 (N_24097,N_18320,N_16358);
or U24098 (N_24098,N_17020,N_19010);
xor U24099 (N_24099,N_17209,N_17403);
nand U24100 (N_24100,N_17177,N_18401);
or U24101 (N_24101,N_17672,N_16230);
nor U24102 (N_24102,N_17546,N_18944);
nand U24103 (N_24103,N_18969,N_15578);
and U24104 (N_24104,N_18341,N_17541);
xor U24105 (N_24105,N_16387,N_18302);
nand U24106 (N_24106,N_18185,N_18586);
xnor U24107 (N_24107,N_17950,N_18431);
or U24108 (N_24108,N_19546,N_19116);
and U24109 (N_24109,N_16342,N_17270);
xor U24110 (N_24110,N_17419,N_18896);
or U24111 (N_24111,N_19589,N_17892);
or U24112 (N_24112,N_15922,N_19417);
nor U24113 (N_24113,N_16662,N_17132);
xor U24114 (N_24114,N_15731,N_16166);
and U24115 (N_24115,N_15966,N_17505);
nor U24116 (N_24116,N_17717,N_17099);
nand U24117 (N_24117,N_15065,N_17910);
xnor U24118 (N_24118,N_17392,N_18806);
or U24119 (N_24119,N_16338,N_15396);
or U24120 (N_24120,N_15884,N_16779);
xor U24121 (N_24121,N_18770,N_17743);
nor U24122 (N_24122,N_17226,N_15996);
and U24123 (N_24123,N_19468,N_17396);
xnor U24124 (N_24124,N_18947,N_17491);
xnor U24125 (N_24125,N_18385,N_15464);
and U24126 (N_24126,N_16899,N_19276);
nor U24127 (N_24127,N_15929,N_18549);
or U24128 (N_24128,N_16720,N_19474);
xor U24129 (N_24129,N_17162,N_15801);
xor U24130 (N_24130,N_16005,N_17951);
nand U24131 (N_24131,N_16100,N_19963);
or U24132 (N_24132,N_15693,N_18031);
xor U24133 (N_24133,N_19653,N_19639);
nand U24134 (N_24134,N_15752,N_19118);
nand U24135 (N_24135,N_18208,N_19360);
and U24136 (N_24136,N_15844,N_18888);
nand U24137 (N_24137,N_18249,N_15222);
nand U24138 (N_24138,N_18126,N_15595);
nand U24139 (N_24139,N_17383,N_19603);
and U24140 (N_24140,N_16220,N_16551);
xor U24141 (N_24141,N_16638,N_15587);
xnor U24142 (N_24142,N_16786,N_17550);
nand U24143 (N_24143,N_15190,N_18055);
and U24144 (N_24144,N_18675,N_16562);
and U24145 (N_24145,N_16547,N_15886);
or U24146 (N_24146,N_18020,N_17936);
nor U24147 (N_24147,N_16443,N_17455);
xor U24148 (N_24148,N_18369,N_19857);
nand U24149 (N_24149,N_16720,N_18625);
nor U24150 (N_24150,N_15271,N_15011);
or U24151 (N_24151,N_19741,N_17838);
and U24152 (N_24152,N_18133,N_19791);
and U24153 (N_24153,N_17603,N_16268);
and U24154 (N_24154,N_16787,N_18931);
xor U24155 (N_24155,N_17332,N_17913);
and U24156 (N_24156,N_19397,N_19170);
and U24157 (N_24157,N_18907,N_17029);
xnor U24158 (N_24158,N_15903,N_15448);
nand U24159 (N_24159,N_18467,N_19785);
xnor U24160 (N_24160,N_19977,N_15792);
or U24161 (N_24161,N_17844,N_17790);
or U24162 (N_24162,N_17296,N_19852);
and U24163 (N_24163,N_17670,N_17265);
nor U24164 (N_24164,N_18857,N_19493);
or U24165 (N_24165,N_17804,N_15281);
and U24166 (N_24166,N_16940,N_15385);
xor U24167 (N_24167,N_17903,N_16954);
nand U24168 (N_24168,N_18488,N_15629);
nand U24169 (N_24169,N_15233,N_18620);
nor U24170 (N_24170,N_18177,N_15915);
xnor U24171 (N_24171,N_18604,N_19498);
and U24172 (N_24172,N_15471,N_18409);
xnor U24173 (N_24173,N_19952,N_16914);
nor U24174 (N_24174,N_19445,N_19226);
xnor U24175 (N_24175,N_15181,N_17488);
xor U24176 (N_24176,N_18283,N_18990);
nand U24177 (N_24177,N_19006,N_15211);
nand U24178 (N_24178,N_15765,N_16150);
nor U24179 (N_24179,N_17817,N_16491);
and U24180 (N_24180,N_17467,N_16968);
xnor U24181 (N_24181,N_17295,N_18402);
or U24182 (N_24182,N_18143,N_19078);
and U24183 (N_24183,N_18928,N_15049);
and U24184 (N_24184,N_17396,N_17954);
nor U24185 (N_24185,N_19609,N_17261);
and U24186 (N_24186,N_18401,N_18581);
and U24187 (N_24187,N_18377,N_15337);
nor U24188 (N_24188,N_17658,N_16424);
xor U24189 (N_24189,N_17195,N_18826);
and U24190 (N_24190,N_18900,N_19126);
nand U24191 (N_24191,N_18705,N_19648);
xnor U24192 (N_24192,N_18731,N_15423);
nand U24193 (N_24193,N_15336,N_15530);
and U24194 (N_24194,N_19725,N_19911);
and U24195 (N_24195,N_19056,N_17745);
and U24196 (N_24196,N_16731,N_17200);
nor U24197 (N_24197,N_18594,N_19947);
xnor U24198 (N_24198,N_19102,N_19238);
or U24199 (N_24199,N_17601,N_17038);
xnor U24200 (N_24200,N_18327,N_18926);
xnor U24201 (N_24201,N_15234,N_18133);
xor U24202 (N_24202,N_17474,N_18212);
or U24203 (N_24203,N_17498,N_16947);
xor U24204 (N_24204,N_17112,N_16700);
xor U24205 (N_24205,N_16045,N_19860);
nand U24206 (N_24206,N_16241,N_18092);
xor U24207 (N_24207,N_18295,N_16094);
nand U24208 (N_24208,N_15965,N_17860);
nor U24209 (N_24209,N_16241,N_16040);
xnor U24210 (N_24210,N_18542,N_15136);
nand U24211 (N_24211,N_16616,N_19066);
nor U24212 (N_24212,N_19585,N_15381);
or U24213 (N_24213,N_19265,N_15459);
xor U24214 (N_24214,N_19499,N_17050);
xor U24215 (N_24215,N_19976,N_17790);
or U24216 (N_24216,N_17472,N_18355);
and U24217 (N_24217,N_18395,N_17447);
or U24218 (N_24218,N_18435,N_17278);
xor U24219 (N_24219,N_17484,N_16720);
or U24220 (N_24220,N_15983,N_19461);
or U24221 (N_24221,N_19598,N_18338);
nand U24222 (N_24222,N_15009,N_17904);
and U24223 (N_24223,N_17561,N_16878);
nor U24224 (N_24224,N_15705,N_17537);
xor U24225 (N_24225,N_19382,N_15976);
or U24226 (N_24226,N_16020,N_17905);
nor U24227 (N_24227,N_19646,N_19524);
and U24228 (N_24228,N_16756,N_19127);
nor U24229 (N_24229,N_15166,N_19511);
xor U24230 (N_24230,N_16333,N_17140);
or U24231 (N_24231,N_19653,N_19326);
nor U24232 (N_24232,N_15388,N_16909);
nand U24233 (N_24233,N_18478,N_17229);
and U24234 (N_24234,N_16946,N_18200);
nor U24235 (N_24235,N_15375,N_19839);
xnor U24236 (N_24236,N_15034,N_18678);
or U24237 (N_24237,N_17894,N_18406);
nor U24238 (N_24238,N_15467,N_16555);
nand U24239 (N_24239,N_17581,N_19288);
and U24240 (N_24240,N_16842,N_17476);
xnor U24241 (N_24241,N_15798,N_17827);
xnor U24242 (N_24242,N_18815,N_19198);
nor U24243 (N_24243,N_15069,N_15926);
nor U24244 (N_24244,N_18593,N_19055);
nor U24245 (N_24245,N_19293,N_19347);
nand U24246 (N_24246,N_17059,N_17716);
or U24247 (N_24247,N_15615,N_15849);
nand U24248 (N_24248,N_18459,N_17283);
xor U24249 (N_24249,N_17944,N_19980);
xor U24250 (N_24250,N_16272,N_15953);
and U24251 (N_24251,N_17501,N_19429);
or U24252 (N_24252,N_15568,N_17703);
or U24253 (N_24253,N_17272,N_18921);
nand U24254 (N_24254,N_15769,N_17454);
xnor U24255 (N_24255,N_18077,N_18197);
and U24256 (N_24256,N_18122,N_18244);
and U24257 (N_24257,N_16146,N_15478);
xnor U24258 (N_24258,N_18999,N_16684);
nor U24259 (N_24259,N_17748,N_15039);
or U24260 (N_24260,N_15322,N_15351);
nor U24261 (N_24261,N_17495,N_17828);
and U24262 (N_24262,N_17983,N_16325);
or U24263 (N_24263,N_19624,N_15861);
nand U24264 (N_24264,N_18173,N_19286);
or U24265 (N_24265,N_15632,N_15582);
nand U24266 (N_24266,N_16846,N_18955);
xor U24267 (N_24267,N_15109,N_18830);
and U24268 (N_24268,N_15154,N_16668);
nand U24269 (N_24269,N_18112,N_18975);
nor U24270 (N_24270,N_15013,N_15561);
nand U24271 (N_24271,N_16321,N_16487);
and U24272 (N_24272,N_19377,N_17785);
nand U24273 (N_24273,N_15051,N_18315);
nand U24274 (N_24274,N_18222,N_18911);
and U24275 (N_24275,N_18803,N_16628);
nand U24276 (N_24276,N_17763,N_18719);
nand U24277 (N_24277,N_18179,N_18937);
nor U24278 (N_24278,N_16397,N_16723);
xor U24279 (N_24279,N_17178,N_15899);
xor U24280 (N_24280,N_15944,N_18345);
or U24281 (N_24281,N_16826,N_19844);
or U24282 (N_24282,N_17715,N_19697);
or U24283 (N_24283,N_18069,N_19959);
xnor U24284 (N_24284,N_17772,N_15500);
xor U24285 (N_24285,N_18304,N_19668);
nand U24286 (N_24286,N_19172,N_16828);
or U24287 (N_24287,N_18315,N_18461);
and U24288 (N_24288,N_18100,N_15650);
nor U24289 (N_24289,N_17912,N_19206);
nor U24290 (N_24290,N_19468,N_19442);
nor U24291 (N_24291,N_15649,N_18968);
xor U24292 (N_24292,N_18801,N_19292);
and U24293 (N_24293,N_18863,N_17060);
or U24294 (N_24294,N_19513,N_17694);
xnor U24295 (N_24295,N_19341,N_16023);
and U24296 (N_24296,N_19954,N_18096);
and U24297 (N_24297,N_16601,N_17507);
nor U24298 (N_24298,N_18081,N_16056);
nor U24299 (N_24299,N_17461,N_19869);
or U24300 (N_24300,N_19518,N_18956);
nand U24301 (N_24301,N_15636,N_19835);
nor U24302 (N_24302,N_15801,N_18507);
nor U24303 (N_24303,N_17088,N_17604);
xor U24304 (N_24304,N_16982,N_18463);
xnor U24305 (N_24305,N_15623,N_17252);
xnor U24306 (N_24306,N_16758,N_15692);
or U24307 (N_24307,N_19630,N_15756);
xor U24308 (N_24308,N_17814,N_18457);
or U24309 (N_24309,N_18680,N_19050);
or U24310 (N_24310,N_16514,N_17459);
nand U24311 (N_24311,N_16367,N_18284);
or U24312 (N_24312,N_17139,N_19575);
nand U24313 (N_24313,N_19558,N_17657);
xnor U24314 (N_24314,N_18233,N_15863);
nor U24315 (N_24315,N_19238,N_15216);
xor U24316 (N_24316,N_17575,N_18080);
nand U24317 (N_24317,N_17927,N_18976);
or U24318 (N_24318,N_16536,N_17477);
nor U24319 (N_24319,N_16221,N_16982);
and U24320 (N_24320,N_15090,N_17193);
or U24321 (N_24321,N_18744,N_19923);
or U24322 (N_24322,N_15801,N_15088);
nand U24323 (N_24323,N_15114,N_19528);
nand U24324 (N_24324,N_17641,N_18696);
nand U24325 (N_24325,N_17774,N_19398);
nand U24326 (N_24326,N_18894,N_15491);
or U24327 (N_24327,N_16505,N_16792);
xnor U24328 (N_24328,N_17192,N_16560);
xnor U24329 (N_24329,N_15652,N_18394);
nand U24330 (N_24330,N_15616,N_15594);
xor U24331 (N_24331,N_18616,N_16602);
nand U24332 (N_24332,N_17200,N_16761);
nand U24333 (N_24333,N_18953,N_18603);
and U24334 (N_24334,N_17290,N_18357);
and U24335 (N_24335,N_16093,N_18376);
and U24336 (N_24336,N_19582,N_17927);
nor U24337 (N_24337,N_15505,N_18816);
xnor U24338 (N_24338,N_16775,N_18979);
nand U24339 (N_24339,N_18951,N_15544);
or U24340 (N_24340,N_16665,N_17740);
xnor U24341 (N_24341,N_18031,N_18057);
nand U24342 (N_24342,N_16015,N_17681);
nand U24343 (N_24343,N_17323,N_15751);
xnor U24344 (N_24344,N_15367,N_15764);
nor U24345 (N_24345,N_16867,N_17692);
and U24346 (N_24346,N_18890,N_16781);
xor U24347 (N_24347,N_16420,N_15927);
or U24348 (N_24348,N_16855,N_18517);
or U24349 (N_24349,N_15599,N_19902);
nand U24350 (N_24350,N_15703,N_19303);
and U24351 (N_24351,N_18043,N_19249);
xnor U24352 (N_24352,N_19291,N_19854);
and U24353 (N_24353,N_15348,N_17158);
xor U24354 (N_24354,N_16860,N_15330);
or U24355 (N_24355,N_15763,N_17233);
and U24356 (N_24356,N_17343,N_15085);
and U24357 (N_24357,N_17287,N_19136);
nand U24358 (N_24358,N_18426,N_15538);
nor U24359 (N_24359,N_19588,N_18508);
nor U24360 (N_24360,N_19498,N_18491);
or U24361 (N_24361,N_15390,N_17813);
nand U24362 (N_24362,N_18104,N_19309);
nor U24363 (N_24363,N_19080,N_17606);
and U24364 (N_24364,N_19472,N_17430);
xor U24365 (N_24365,N_17457,N_19753);
nand U24366 (N_24366,N_19395,N_19873);
and U24367 (N_24367,N_17263,N_18204);
xor U24368 (N_24368,N_17301,N_19957);
nor U24369 (N_24369,N_15207,N_18893);
nor U24370 (N_24370,N_18893,N_17696);
nand U24371 (N_24371,N_18526,N_16134);
and U24372 (N_24372,N_16409,N_15143);
and U24373 (N_24373,N_17544,N_15208);
xnor U24374 (N_24374,N_15196,N_19423);
nor U24375 (N_24375,N_18154,N_16737);
nand U24376 (N_24376,N_16226,N_19953);
and U24377 (N_24377,N_19668,N_18506);
and U24378 (N_24378,N_18989,N_16093);
nor U24379 (N_24379,N_17596,N_19288);
nor U24380 (N_24380,N_16711,N_18480);
and U24381 (N_24381,N_19256,N_15238);
xnor U24382 (N_24382,N_17599,N_16633);
nor U24383 (N_24383,N_19402,N_19851);
and U24384 (N_24384,N_18935,N_16795);
nand U24385 (N_24385,N_16034,N_16148);
nand U24386 (N_24386,N_17380,N_18151);
nor U24387 (N_24387,N_16691,N_18273);
or U24388 (N_24388,N_18486,N_18121);
and U24389 (N_24389,N_17117,N_17629);
or U24390 (N_24390,N_16832,N_15569);
or U24391 (N_24391,N_15144,N_19829);
xnor U24392 (N_24392,N_19240,N_15076);
and U24393 (N_24393,N_15760,N_19168);
nand U24394 (N_24394,N_15309,N_18499);
nand U24395 (N_24395,N_19846,N_18514);
xnor U24396 (N_24396,N_18539,N_15762);
nor U24397 (N_24397,N_17371,N_19790);
xor U24398 (N_24398,N_18837,N_19338);
nand U24399 (N_24399,N_16448,N_16481);
and U24400 (N_24400,N_18136,N_18265);
and U24401 (N_24401,N_15501,N_15625);
nor U24402 (N_24402,N_19524,N_16180);
nand U24403 (N_24403,N_19611,N_15662);
nand U24404 (N_24404,N_15561,N_17390);
or U24405 (N_24405,N_18230,N_17573);
xnor U24406 (N_24406,N_15477,N_19920);
xor U24407 (N_24407,N_15755,N_16884);
or U24408 (N_24408,N_16626,N_17760);
or U24409 (N_24409,N_18430,N_16850);
xor U24410 (N_24410,N_17365,N_17895);
nand U24411 (N_24411,N_15670,N_18161);
or U24412 (N_24412,N_18952,N_19283);
xor U24413 (N_24413,N_17196,N_16364);
xnor U24414 (N_24414,N_19631,N_16713);
nand U24415 (N_24415,N_15721,N_19947);
xnor U24416 (N_24416,N_16197,N_16204);
xor U24417 (N_24417,N_15415,N_18172);
or U24418 (N_24418,N_15959,N_15191);
nand U24419 (N_24419,N_19139,N_16129);
nor U24420 (N_24420,N_17300,N_18434);
nand U24421 (N_24421,N_18351,N_17329);
nand U24422 (N_24422,N_19582,N_18186);
xnor U24423 (N_24423,N_18677,N_15967);
nor U24424 (N_24424,N_16621,N_17295);
nor U24425 (N_24425,N_16740,N_16776);
xor U24426 (N_24426,N_19940,N_19322);
and U24427 (N_24427,N_15227,N_15334);
nor U24428 (N_24428,N_16010,N_17090);
xnor U24429 (N_24429,N_16212,N_17050);
nor U24430 (N_24430,N_15882,N_17122);
and U24431 (N_24431,N_19461,N_17360);
nor U24432 (N_24432,N_17135,N_19449);
nor U24433 (N_24433,N_16873,N_19946);
or U24434 (N_24434,N_18636,N_18866);
and U24435 (N_24435,N_19614,N_15930);
or U24436 (N_24436,N_15801,N_18264);
nand U24437 (N_24437,N_18278,N_17041);
and U24438 (N_24438,N_18880,N_19357);
nand U24439 (N_24439,N_16472,N_18150);
nand U24440 (N_24440,N_15150,N_19090);
nor U24441 (N_24441,N_19166,N_18358);
and U24442 (N_24442,N_18790,N_15736);
nand U24443 (N_24443,N_17835,N_16913);
xor U24444 (N_24444,N_19436,N_16999);
xor U24445 (N_24445,N_18788,N_15930);
xor U24446 (N_24446,N_19303,N_16425);
and U24447 (N_24447,N_18066,N_17811);
nor U24448 (N_24448,N_18593,N_17188);
nor U24449 (N_24449,N_18683,N_15019);
and U24450 (N_24450,N_17014,N_18615);
xor U24451 (N_24451,N_19575,N_16496);
and U24452 (N_24452,N_19851,N_17463);
nor U24453 (N_24453,N_18492,N_17966);
nor U24454 (N_24454,N_15487,N_16284);
nor U24455 (N_24455,N_16959,N_16145);
nand U24456 (N_24456,N_17877,N_18715);
or U24457 (N_24457,N_16164,N_15404);
and U24458 (N_24458,N_18770,N_17617);
xnor U24459 (N_24459,N_16240,N_17472);
xnor U24460 (N_24460,N_15185,N_15841);
and U24461 (N_24461,N_17715,N_17008);
xor U24462 (N_24462,N_19048,N_17313);
or U24463 (N_24463,N_15636,N_17497);
nand U24464 (N_24464,N_15782,N_15453);
and U24465 (N_24465,N_18037,N_18823);
or U24466 (N_24466,N_17261,N_18858);
and U24467 (N_24467,N_19196,N_17484);
nor U24468 (N_24468,N_18799,N_18953);
nor U24469 (N_24469,N_17673,N_16430);
or U24470 (N_24470,N_18035,N_15487);
nor U24471 (N_24471,N_15798,N_17291);
nor U24472 (N_24472,N_17848,N_15313);
xor U24473 (N_24473,N_15454,N_18846);
xor U24474 (N_24474,N_19296,N_18347);
nor U24475 (N_24475,N_17264,N_18939);
nor U24476 (N_24476,N_16384,N_19823);
or U24477 (N_24477,N_17357,N_19889);
nand U24478 (N_24478,N_18164,N_19301);
xnor U24479 (N_24479,N_16947,N_15605);
nand U24480 (N_24480,N_15861,N_17160);
or U24481 (N_24481,N_19371,N_19805);
nor U24482 (N_24482,N_18233,N_18821);
nor U24483 (N_24483,N_19262,N_16302);
nand U24484 (N_24484,N_17504,N_19007);
and U24485 (N_24485,N_18149,N_16161);
nand U24486 (N_24486,N_15040,N_15206);
and U24487 (N_24487,N_15695,N_18388);
and U24488 (N_24488,N_18521,N_15383);
and U24489 (N_24489,N_17463,N_19275);
and U24490 (N_24490,N_16250,N_15791);
and U24491 (N_24491,N_16749,N_19069);
nand U24492 (N_24492,N_16571,N_17755);
xor U24493 (N_24493,N_15276,N_19700);
or U24494 (N_24494,N_19595,N_15220);
xor U24495 (N_24495,N_18644,N_16084);
or U24496 (N_24496,N_16055,N_18554);
xnor U24497 (N_24497,N_15354,N_19101);
xor U24498 (N_24498,N_17637,N_18559);
nor U24499 (N_24499,N_15575,N_18823);
nand U24500 (N_24500,N_18626,N_17002);
or U24501 (N_24501,N_17708,N_17232);
nand U24502 (N_24502,N_17873,N_16500);
nor U24503 (N_24503,N_19857,N_16010);
xnor U24504 (N_24504,N_15065,N_16139);
nand U24505 (N_24505,N_18876,N_16096);
xnor U24506 (N_24506,N_16705,N_16518);
nor U24507 (N_24507,N_18109,N_16994);
and U24508 (N_24508,N_15917,N_17547);
and U24509 (N_24509,N_15068,N_17597);
nor U24510 (N_24510,N_15334,N_17370);
nor U24511 (N_24511,N_15373,N_18143);
xnor U24512 (N_24512,N_18155,N_17424);
nor U24513 (N_24513,N_17478,N_18159);
nand U24514 (N_24514,N_17285,N_16282);
nand U24515 (N_24515,N_18299,N_18921);
nor U24516 (N_24516,N_18374,N_16676);
nand U24517 (N_24517,N_16093,N_16417);
xor U24518 (N_24518,N_17764,N_17802);
nand U24519 (N_24519,N_17925,N_19561);
xor U24520 (N_24520,N_16584,N_15910);
or U24521 (N_24521,N_15172,N_18270);
nand U24522 (N_24522,N_19742,N_17569);
nand U24523 (N_24523,N_17852,N_18894);
and U24524 (N_24524,N_16114,N_18906);
nand U24525 (N_24525,N_15282,N_18165);
xor U24526 (N_24526,N_16756,N_16602);
and U24527 (N_24527,N_19627,N_16044);
or U24528 (N_24528,N_16874,N_19145);
nand U24529 (N_24529,N_18758,N_16186);
or U24530 (N_24530,N_19517,N_18953);
and U24531 (N_24531,N_19596,N_16677);
nor U24532 (N_24532,N_17649,N_16416);
xor U24533 (N_24533,N_15042,N_15332);
nand U24534 (N_24534,N_17268,N_19352);
nor U24535 (N_24535,N_16635,N_19043);
xor U24536 (N_24536,N_17539,N_16006);
or U24537 (N_24537,N_16322,N_15419);
or U24538 (N_24538,N_16331,N_15465);
and U24539 (N_24539,N_17301,N_18240);
xor U24540 (N_24540,N_15765,N_15443);
xor U24541 (N_24541,N_19177,N_16332);
nor U24542 (N_24542,N_16540,N_17856);
nand U24543 (N_24543,N_16954,N_19477);
xor U24544 (N_24544,N_19133,N_19898);
or U24545 (N_24545,N_16935,N_16341);
or U24546 (N_24546,N_16708,N_18990);
nand U24547 (N_24547,N_15625,N_15949);
nor U24548 (N_24548,N_15432,N_17451);
xor U24549 (N_24549,N_15988,N_18485);
nand U24550 (N_24550,N_18068,N_17072);
xnor U24551 (N_24551,N_17168,N_15722);
nor U24552 (N_24552,N_15126,N_19166);
xor U24553 (N_24553,N_18503,N_15878);
nand U24554 (N_24554,N_16640,N_15485);
or U24555 (N_24555,N_15260,N_17169);
and U24556 (N_24556,N_18512,N_19463);
and U24557 (N_24557,N_17311,N_15729);
xnor U24558 (N_24558,N_18208,N_19363);
xor U24559 (N_24559,N_15216,N_15980);
and U24560 (N_24560,N_16928,N_18563);
nand U24561 (N_24561,N_17940,N_17911);
or U24562 (N_24562,N_15956,N_16914);
nor U24563 (N_24563,N_18079,N_18574);
and U24564 (N_24564,N_17317,N_16451);
nor U24565 (N_24565,N_17094,N_18046);
and U24566 (N_24566,N_16578,N_19290);
or U24567 (N_24567,N_17275,N_15194);
and U24568 (N_24568,N_18786,N_17544);
nor U24569 (N_24569,N_15131,N_17793);
or U24570 (N_24570,N_16388,N_19264);
and U24571 (N_24571,N_17827,N_17563);
nor U24572 (N_24572,N_15157,N_15538);
nand U24573 (N_24573,N_18462,N_18131);
nor U24574 (N_24574,N_18343,N_15912);
nand U24575 (N_24575,N_18781,N_16671);
nand U24576 (N_24576,N_18217,N_19283);
and U24577 (N_24577,N_15797,N_17237);
and U24578 (N_24578,N_15505,N_17872);
and U24579 (N_24579,N_18274,N_18501);
and U24580 (N_24580,N_19547,N_15465);
or U24581 (N_24581,N_18527,N_19222);
or U24582 (N_24582,N_19514,N_17317);
and U24583 (N_24583,N_18872,N_15064);
or U24584 (N_24584,N_15079,N_16322);
xnor U24585 (N_24585,N_17808,N_15645);
nor U24586 (N_24586,N_17233,N_19278);
nor U24587 (N_24587,N_17106,N_15668);
and U24588 (N_24588,N_15457,N_16463);
xor U24589 (N_24589,N_18247,N_18048);
xor U24590 (N_24590,N_19651,N_15278);
xnor U24591 (N_24591,N_17223,N_15551);
and U24592 (N_24592,N_15547,N_19273);
nor U24593 (N_24593,N_16500,N_18157);
nand U24594 (N_24594,N_18471,N_15063);
nand U24595 (N_24595,N_15874,N_18003);
xor U24596 (N_24596,N_18912,N_16221);
nor U24597 (N_24597,N_19849,N_16293);
nor U24598 (N_24598,N_18533,N_16365);
or U24599 (N_24599,N_17523,N_19905);
xnor U24600 (N_24600,N_19644,N_16548);
xnor U24601 (N_24601,N_17805,N_17668);
nor U24602 (N_24602,N_19634,N_15288);
nor U24603 (N_24603,N_16504,N_18627);
nor U24604 (N_24604,N_15508,N_17933);
nand U24605 (N_24605,N_15817,N_19879);
and U24606 (N_24606,N_18073,N_16044);
or U24607 (N_24607,N_16402,N_15948);
nor U24608 (N_24608,N_15503,N_17600);
nor U24609 (N_24609,N_19986,N_17574);
and U24610 (N_24610,N_16656,N_16883);
nand U24611 (N_24611,N_16653,N_17203);
or U24612 (N_24612,N_16062,N_16206);
xnor U24613 (N_24613,N_15550,N_19271);
or U24614 (N_24614,N_19747,N_17844);
nor U24615 (N_24615,N_15708,N_15079);
and U24616 (N_24616,N_17841,N_15109);
nand U24617 (N_24617,N_15635,N_15135);
and U24618 (N_24618,N_15235,N_15426);
xnor U24619 (N_24619,N_17159,N_18557);
or U24620 (N_24620,N_16399,N_19198);
or U24621 (N_24621,N_17496,N_17540);
xor U24622 (N_24622,N_17392,N_16277);
and U24623 (N_24623,N_16311,N_15709);
nor U24624 (N_24624,N_16861,N_19522);
and U24625 (N_24625,N_18563,N_15040);
and U24626 (N_24626,N_15604,N_15018);
and U24627 (N_24627,N_18084,N_16897);
nor U24628 (N_24628,N_17832,N_19376);
xor U24629 (N_24629,N_18606,N_19910);
nor U24630 (N_24630,N_17586,N_17044);
xnor U24631 (N_24631,N_15902,N_19554);
nand U24632 (N_24632,N_19337,N_16521);
nor U24633 (N_24633,N_19732,N_17577);
nor U24634 (N_24634,N_18477,N_19545);
xnor U24635 (N_24635,N_18067,N_15730);
nor U24636 (N_24636,N_17100,N_18002);
xor U24637 (N_24637,N_15598,N_17322);
or U24638 (N_24638,N_17611,N_18598);
and U24639 (N_24639,N_15096,N_16712);
and U24640 (N_24640,N_15551,N_16749);
xnor U24641 (N_24641,N_18322,N_19367);
nand U24642 (N_24642,N_17777,N_19874);
or U24643 (N_24643,N_18932,N_15675);
nor U24644 (N_24644,N_18982,N_19812);
xor U24645 (N_24645,N_17010,N_18793);
nand U24646 (N_24646,N_19776,N_16705);
xor U24647 (N_24647,N_18551,N_18990);
and U24648 (N_24648,N_15700,N_15326);
nor U24649 (N_24649,N_17923,N_18235);
xor U24650 (N_24650,N_17860,N_17818);
and U24651 (N_24651,N_15658,N_16318);
xnor U24652 (N_24652,N_15838,N_18057);
nand U24653 (N_24653,N_16330,N_19005);
nor U24654 (N_24654,N_16569,N_16745);
xor U24655 (N_24655,N_17269,N_18196);
or U24656 (N_24656,N_17004,N_17839);
xnor U24657 (N_24657,N_18377,N_19010);
nand U24658 (N_24658,N_17718,N_18679);
nor U24659 (N_24659,N_17645,N_16689);
nor U24660 (N_24660,N_15381,N_19420);
nor U24661 (N_24661,N_16476,N_16121);
and U24662 (N_24662,N_15857,N_16187);
xnor U24663 (N_24663,N_17323,N_19977);
or U24664 (N_24664,N_19246,N_15973);
or U24665 (N_24665,N_15480,N_19951);
nor U24666 (N_24666,N_19597,N_17189);
or U24667 (N_24667,N_15552,N_19320);
xor U24668 (N_24668,N_19406,N_19309);
nor U24669 (N_24669,N_15756,N_16231);
xnor U24670 (N_24670,N_15408,N_19167);
nand U24671 (N_24671,N_17408,N_19460);
and U24672 (N_24672,N_18661,N_19850);
nor U24673 (N_24673,N_18408,N_17308);
xnor U24674 (N_24674,N_16499,N_17118);
nor U24675 (N_24675,N_19656,N_18492);
or U24676 (N_24676,N_19673,N_18662);
nand U24677 (N_24677,N_19353,N_15593);
or U24678 (N_24678,N_19508,N_16462);
or U24679 (N_24679,N_19481,N_16156);
nor U24680 (N_24680,N_15388,N_17191);
or U24681 (N_24681,N_16857,N_19701);
xor U24682 (N_24682,N_19537,N_19035);
nand U24683 (N_24683,N_18112,N_16283);
nor U24684 (N_24684,N_16129,N_19700);
and U24685 (N_24685,N_18199,N_15145);
nor U24686 (N_24686,N_18478,N_16674);
xor U24687 (N_24687,N_17843,N_18468);
and U24688 (N_24688,N_18197,N_19934);
xor U24689 (N_24689,N_17590,N_18263);
nor U24690 (N_24690,N_19226,N_15325);
nor U24691 (N_24691,N_17899,N_15658);
nor U24692 (N_24692,N_19360,N_16346);
xnor U24693 (N_24693,N_16645,N_15490);
or U24694 (N_24694,N_16443,N_18356);
xnor U24695 (N_24695,N_15653,N_19832);
and U24696 (N_24696,N_18846,N_17971);
and U24697 (N_24697,N_16075,N_17816);
nand U24698 (N_24698,N_18651,N_19160);
nand U24699 (N_24699,N_19401,N_15395);
and U24700 (N_24700,N_18642,N_18286);
or U24701 (N_24701,N_19347,N_18858);
and U24702 (N_24702,N_15114,N_17050);
xor U24703 (N_24703,N_16044,N_17643);
nor U24704 (N_24704,N_18291,N_15059);
xor U24705 (N_24705,N_16590,N_19615);
or U24706 (N_24706,N_19070,N_17953);
and U24707 (N_24707,N_16630,N_15029);
nand U24708 (N_24708,N_17688,N_18654);
and U24709 (N_24709,N_16365,N_19820);
xnor U24710 (N_24710,N_19818,N_17192);
or U24711 (N_24711,N_19341,N_16651);
xnor U24712 (N_24712,N_17650,N_15031);
xnor U24713 (N_24713,N_17489,N_18484);
nand U24714 (N_24714,N_17723,N_19680);
xor U24715 (N_24715,N_17134,N_16962);
xor U24716 (N_24716,N_15834,N_16943);
nor U24717 (N_24717,N_17917,N_16677);
and U24718 (N_24718,N_18226,N_15030);
and U24719 (N_24719,N_17760,N_15233);
xor U24720 (N_24720,N_18276,N_17552);
nand U24721 (N_24721,N_15320,N_17379);
or U24722 (N_24722,N_18917,N_16647);
nand U24723 (N_24723,N_15465,N_17288);
or U24724 (N_24724,N_15280,N_16438);
nor U24725 (N_24725,N_19561,N_16099);
or U24726 (N_24726,N_17754,N_18734);
nor U24727 (N_24727,N_18724,N_16299);
xnor U24728 (N_24728,N_17751,N_17852);
xor U24729 (N_24729,N_15630,N_18639);
or U24730 (N_24730,N_15798,N_18971);
or U24731 (N_24731,N_18799,N_17188);
and U24732 (N_24732,N_19566,N_17673);
nand U24733 (N_24733,N_16321,N_18465);
nand U24734 (N_24734,N_17524,N_15631);
nor U24735 (N_24735,N_17474,N_17764);
and U24736 (N_24736,N_17587,N_18279);
or U24737 (N_24737,N_15721,N_18371);
and U24738 (N_24738,N_18453,N_17683);
and U24739 (N_24739,N_19432,N_15382);
nand U24740 (N_24740,N_17042,N_15849);
nand U24741 (N_24741,N_16509,N_15431);
and U24742 (N_24742,N_18784,N_15699);
xor U24743 (N_24743,N_19040,N_19322);
and U24744 (N_24744,N_17092,N_16265);
nand U24745 (N_24745,N_15466,N_19351);
or U24746 (N_24746,N_18548,N_19541);
xnor U24747 (N_24747,N_16358,N_17189);
and U24748 (N_24748,N_17923,N_17548);
and U24749 (N_24749,N_19946,N_15557);
and U24750 (N_24750,N_15631,N_15857);
nand U24751 (N_24751,N_17850,N_15876);
xor U24752 (N_24752,N_17508,N_19856);
and U24753 (N_24753,N_19393,N_19106);
xnor U24754 (N_24754,N_15913,N_19720);
nor U24755 (N_24755,N_15476,N_16816);
nand U24756 (N_24756,N_18180,N_17426);
and U24757 (N_24757,N_18543,N_15284);
and U24758 (N_24758,N_19436,N_16611);
xor U24759 (N_24759,N_17538,N_18824);
nor U24760 (N_24760,N_17412,N_19795);
nand U24761 (N_24761,N_18156,N_18204);
xnor U24762 (N_24762,N_16425,N_19245);
nor U24763 (N_24763,N_16291,N_19819);
and U24764 (N_24764,N_19140,N_19374);
nand U24765 (N_24765,N_15085,N_19949);
nor U24766 (N_24766,N_15800,N_16499);
nand U24767 (N_24767,N_18472,N_15175);
and U24768 (N_24768,N_18482,N_17693);
nand U24769 (N_24769,N_15558,N_17799);
or U24770 (N_24770,N_19231,N_19754);
xor U24771 (N_24771,N_17833,N_19891);
and U24772 (N_24772,N_17662,N_18671);
or U24773 (N_24773,N_19047,N_18865);
nor U24774 (N_24774,N_19683,N_18955);
xnor U24775 (N_24775,N_17987,N_19574);
nand U24776 (N_24776,N_16936,N_16485);
nand U24777 (N_24777,N_18324,N_17647);
and U24778 (N_24778,N_19394,N_17605);
xor U24779 (N_24779,N_16783,N_19594);
xnor U24780 (N_24780,N_17553,N_16101);
nor U24781 (N_24781,N_17193,N_17834);
nor U24782 (N_24782,N_18687,N_18554);
xor U24783 (N_24783,N_18635,N_17287);
xor U24784 (N_24784,N_15560,N_15609);
nor U24785 (N_24785,N_15003,N_18441);
nor U24786 (N_24786,N_15050,N_15807);
nor U24787 (N_24787,N_15252,N_16479);
or U24788 (N_24788,N_16863,N_16356);
nor U24789 (N_24789,N_18308,N_19993);
nand U24790 (N_24790,N_19208,N_19473);
nor U24791 (N_24791,N_16280,N_16212);
or U24792 (N_24792,N_15972,N_16586);
or U24793 (N_24793,N_16529,N_18195);
and U24794 (N_24794,N_17018,N_17571);
nand U24795 (N_24795,N_19767,N_15238);
nor U24796 (N_24796,N_19291,N_18594);
nor U24797 (N_24797,N_17484,N_18453);
or U24798 (N_24798,N_16234,N_15390);
nand U24799 (N_24799,N_16118,N_19564);
nor U24800 (N_24800,N_16204,N_15425);
or U24801 (N_24801,N_15474,N_18897);
nor U24802 (N_24802,N_15320,N_17429);
nor U24803 (N_24803,N_19539,N_17757);
and U24804 (N_24804,N_16645,N_15128);
or U24805 (N_24805,N_18276,N_17134);
or U24806 (N_24806,N_16728,N_19389);
or U24807 (N_24807,N_16802,N_18387);
nor U24808 (N_24808,N_17119,N_19866);
nand U24809 (N_24809,N_15188,N_17062);
nor U24810 (N_24810,N_15299,N_18577);
and U24811 (N_24811,N_15784,N_19241);
and U24812 (N_24812,N_15472,N_16097);
nor U24813 (N_24813,N_17356,N_15158);
nor U24814 (N_24814,N_15346,N_17311);
nor U24815 (N_24815,N_15953,N_15173);
nor U24816 (N_24816,N_16225,N_16058);
and U24817 (N_24817,N_19805,N_19898);
or U24818 (N_24818,N_18820,N_15831);
nand U24819 (N_24819,N_16304,N_17354);
xor U24820 (N_24820,N_16349,N_18733);
nor U24821 (N_24821,N_17411,N_17400);
xor U24822 (N_24822,N_15126,N_17362);
xor U24823 (N_24823,N_18991,N_19742);
nand U24824 (N_24824,N_16317,N_15580);
or U24825 (N_24825,N_19812,N_17275);
and U24826 (N_24826,N_16468,N_18263);
nand U24827 (N_24827,N_17900,N_18296);
xnor U24828 (N_24828,N_17102,N_15554);
or U24829 (N_24829,N_18458,N_16905);
and U24830 (N_24830,N_16006,N_18447);
nand U24831 (N_24831,N_15447,N_18018);
and U24832 (N_24832,N_17109,N_17698);
nand U24833 (N_24833,N_18636,N_18152);
and U24834 (N_24834,N_18671,N_16798);
xor U24835 (N_24835,N_17632,N_16206);
nand U24836 (N_24836,N_17155,N_15198);
xnor U24837 (N_24837,N_18745,N_15457);
and U24838 (N_24838,N_19489,N_18102);
and U24839 (N_24839,N_19537,N_15910);
nand U24840 (N_24840,N_19015,N_17533);
nor U24841 (N_24841,N_19150,N_19770);
nor U24842 (N_24842,N_18361,N_19501);
or U24843 (N_24843,N_16882,N_16834);
and U24844 (N_24844,N_19097,N_15085);
and U24845 (N_24845,N_19303,N_17075);
or U24846 (N_24846,N_18986,N_15814);
xnor U24847 (N_24847,N_18788,N_15160);
and U24848 (N_24848,N_15313,N_19780);
or U24849 (N_24849,N_18394,N_17363);
or U24850 (N_24850,N_16415,N_19897);
nand U24851 (N_24851,N_17053,N_19544);
and U24852 (N_24852,N_15956,N_18494);
nand U24853 (N_24853,N_18081,N_19347);
nor U24854 (N_24854,N_16644,N_17435);
xor U24855 (N_24855,N_15423,N_16679);
xnor U24856 (N_24856,N_16487,N_15319);
xnor U24857 (N_24857,N_17657,N_19346);
or U24858 (N_24858,N_15010,N_16933);
or U24859 (N_24859,N_17184,N_16271);
xor U24860 (N_24860,N_16131,N_15060);
and U24861 (N_24861,N_17508,N_18771);
xor U24862 (N_24862,N_18749,N_16120);
or U24863 (N_24863,N_19621,N_18533);
nand U24864 (N_24864,N_18781,N_19434);
nor U24865 (N_24865,N_18346,N_17635);
or U24866 (N_24866,N_19081,N_17767);
or U24867 (N_24867,N_17133,N_15349);
xor U24868 (N_24868,N_17907,N_18920);
xor U24869 (N_24869,N_18115,N_17697);
or U24870 (N_24870,N_19057,N_19579);
and U24871 (N_24871,N_18882,N_16541);
and U24872 (N_24872,N_19058,N_18753);
nand U24873 (N_24873,N_19360,N_16244);
nor U24874 (N_24874,N_18183,N_19659);
nor U24875 (N_24875,N_18947,N_16590);
or U24876 (N_24876,N_18705,N_17193);
nor U24877 (N_24877,N_15758,N_15163);
nor U24878 (N_24878,N_19414,N_15460);
or U24879 (N_24879,N_16526,N_19854);
nand U24880 (N_24880,N_18093,N_15577);
nand U24881 (N_24881,N_16322,N_15628);
nor U24882 (N_24882,N_15416,N_18264);
xor U24883 (N_24883,N_16362,N_18251);
nand U24884 (N_24884,N_17619,N_19676);
nand U24885 (N_24885,N_16109,N_17701);
and U24886 (N_24886,N_15397,N_18038);
nand U24887 (N_24887,N_16265,N_18033);
and U24888 (N_24888,N_15166,N_18748);
and U24889 (N_24889,N_15278,N_16149);
nor U24890 (N_24890,N_15928,N_16305);
xnor U24891 (N_24891,N_18249,N_16749);
and U24892 (N_24892,N_17854,N_19939);
and U24893 (N_24893,N_16844,N_19977);
nor U24894 (N_24894,N_15485,N_18078);
nand U24895 (N_24895,N_18994,N_17621);
or U24896 (N_24896,N_16098,N_17398);
and U24897 (N_24897,N_15574,N_17432);
xnor U24898 (N_24898,N_17463,N_15655);
xor U24899 (N_24899,N_18200,N_15916);
xnor U24900 (N_24900,N_16120,N_19579);
nand U24901 (N_24901,N_18183,N_19044);
nand U24902 (N_24902,N_15042,N_19318);
and U24903 (N_24903,N_15767,N_15189);
nor U24904 (N_24904,N_15771,N_16051);
xnor U24905 (N_24905,N_17952,N_17658);
and U24906 (N_24906,N_19804,N_15893);
nor U24907 (N_24907,N_17451,N_18771);
nor U24908 (N_24908,N_19447,N_15027);
nor U24909 (N_24909,N_18434,N_18101);
and U24910 (N_24910,N_17274,N_15888);
nand U24911 (N_24911,N_19991,N_19183);
nor U24912 (N_24912,N_16322,N_19191);
nand U24913 (N_24913,N_18902,N_17408);
and U24914 (N_24914,N_16190,N_15646);
nand U24915 (N_24915,N_15640,N_17425);
xor U24916 (N_24916,N_19472,N_16375);
or U24917 (N_24917,N_16407,N_19289);
nand U24918 (N_24918,N_18541,N_19512);
nor U24919 (N_24919,N_17407,N_19425);
or U24920 (N_24920,N_18473,N_18530);
and U24921 (N_24921,N_18016,N_15853);
or U24922 (N_24922,N_19700,N_19922);
nor U24923 (N_24923,N_18020,N_18817);
nor U24924 (N_24924,N_15484,N_16715);
or U24925 (N_24925,N_17813,N_18870);
and U24926 (N_24926,N_17087,N_17571);
or U24927 (N_24927,N_16655,N_16548);
nor U24928 (N_24928,N_19171,N_16287);
or U24929 (N_24929,N_18113,N_17793);
and U24930 (N_24930,N_19704,N_19782);
and U24931 (N_24931,N_19497,N_19008);
or U24932 (N_24932,N_18250,N_18858);
and U24933 (N_24933,N_16445,N_15005);
nor U24934 (N_24934,N_17676,N_16954);
and U24935 (N_24935,N_18862,N_15152);
or U24936 (N_24936,N_18970,N_18056);
xor U24937 (N_24937,N_19339,N_18003);
xnor U24938 (N_24938,N_16720,N_16830);
nand U24939 (N_24939,N_17616,N_19361);
nor U24940 (N_24940,N_17842,N_19130);
xor U24941 (N_24941,N_15560,N_18374);
or U24942 (N_24942,N_19785,N_16999);
nor U24943 (N_24943,N_17449,N_19555);
or U24944 (N_24944,N_19802,N_16669);
or U24945 (N_24945,N_18037,N_16396);
or U24946 (N_24946,N_16723,N_16087);
xor U24947 (N_24947,N_15116,N_18859);
or U24948 (N_24948,N_17622,N_17799);
and U24949 (N_24949,N_18744,N_15293);
nor U24950 (N_24950,N_18843,N_18199);
or U24951 (N_24951,N_15486,N_15860);
xor U24952 (N_24952,N_18417,N_16807);
xnor U24953 (N_24953,N_18802,N_16164);
xnor U24954 (N_24954,N_17243,N_15877);
nand U24955 (N_24955,N_16369,N_16788);
xnor U24956 (N_24956,N_19269,N_16695);
nor U24957 (N_24957,N_17511,N_18160);
xor U24958 (N_24958,N_19042,N_17417);
and U24959 (N_24959,N_17354,N_15849);
nor U24960 (N_24960,N_18885,N_17978);
or U24961 (N_24961,N_19661,N_16055);
nor U24962 (N_24962,N_17899,N_15477);
or U24963 (N_24963,N_16368,N_19754);
or U24964 (N_24964,N_16607,N_18640);
and U24965 (N_24965,N_19770,N_19925);
and U24966 (N_24966,N_17475,N_16398);
nor U24967 (N_24967,N_19944,N_16747);
or U24968 (N_24968,N_19092,N_17255);
nor U24969 (N_24969,N_17290,N_17451);
xnor U24970 (N_24970,N_17221,N_18273);
nand U24971 (N_24971,N_18761,N_15391);
xor U24972 (N_24972,N_17605,N_19465);
and U24973 (N_24973,N_18245,N_18590);
nor U24974 (N_24974,N_18295,N_17645);
nand U24975 (N_24975,N_15654,N_18688);
or U24976 (N_24976,N_16514,N_17234);
nand U24977 (N_24977,N_17143,N_19989);
nor U24978 (N_24978,N_16221,N_17187);
nor U24979 (N_24979,N_16832,N_18786);
nand U24980 (N_24980,N_18464,N_15870);
nand U24981 (N_24981,N_17824,N_19974);
and U24982 (N_24982,N_19374,N_19323);
xor U24983 (N_24983,N_18503,N_15808);
or U24984 (N_24984,N_19379,N_19652);
and U24985 (N_24985,N_18915,N_17415);
and U24986 (N_24986,N_19138,N_18028);
nand U24987 (N_24987,N_19371,N_15371);
xor U24988 (N_24988,N_17335,N_15750);
and U24989 (N_24989,N_19643,N_15294);
and U24990 (N_24990,N_17110,N_16747);
nor U24991 (N_24991,N_15321,N_16140);
nor U24992 (N_24992,N_15351,N_16499);
or U24993 (N_24993,N_19123,N_16768);
and U24994 (N_24994,N_17278,N_15626);
and U24995 (N_24995,N_16767,N_15834);
nand U24996 (N_24996,N_16163,N_15794);
nand U24997 (N_24997,N_17604,N_17315);
or U24998 (N_24998,N_15463,N_16808);
nand U24999 (N_24999,N_16134,N_19882);
and U25000 (N_25000,N_22102,N_20511);
nor U25001 (N_25001,N_24854,N_23585);
nor U25002 (N_25002,N_21388,N_22440);
xor U25003 (N_25003,N_22633,N_24760);
xnor U25004 (N_25004,N_22457,N_21542);
xnor U25005 (N_25005,N_20648,N_21769);
nand U25006 (N_25006,N_23801,N_21141);
xnor U25007 (N_25007,N_20010,N_22044);
xnor U25008 (N_25008,N_24010,N_21168);
nor U25009 (N_25009,N_24465,N_22798);
nor U25010 (N_25010,N_21371,N_20689);
or U25011 (N_25011,N_21875,N_24041);
xnor U25012 (N_25012,N_20722,N_23796);
nand U25013 (N_25013,N_22425,N_24392);
xnor U25014 (N_25014,N_24403,N_23149);
nand U25015 (N_25015,N_21179,N_23010);
nand U25016 (N_25016,N_21585,N_22038);
and U25017 (N_25017,N_21402,N_20543);
xnor U25018 (N_25018,N_24697,N_24445);
or U25019 (N_25019,N_21060,N_21240);
or U25020 (N_25020,N_24668,N_22476);
xor U25021 (N_25021,N_24990,N_24607);
and U25022 (N_25022,N_23685,N_23275);
nand U25023 (N_25023,N_24974,N_21939);
and U25024 (N_25024,N_24147,N_20277);
xnor U25025 (N_25025,N_22692,N_24785);
nor U25026 (N_25026,N_20681,N_20774);
and U25027 (N_25027,N_22793,N_24376);
or U25028 (N_25028,N_23199,N_23688);
and U25029 (N_25029,N_20215,N_22853);
and U25030 (N_25030,N_24433,N_22138);
and U25031 (N_25031,N_24837,N_20286);
nor U25032 (N_25032,N_20747,N_21699);
nand U25033 (N_25033,N_22687,N_24282);
nand U25034 (N_25034,N_23881,N_20849);
xor U25035 (N_25035,N_24371,N_22372);
nor U25036 (N_25036,N_23743,N_21719);
nor U25037 (N_25037,N_21811,N_22471);
xor U25038 (N_25038,N_24358,N_23464);
nor U25039 (N_25039,N_21018,N_22479);
and U25040 (N_25040,N_23193,N_24917);
or U25041 (N_25041,N_20516,N_20556);
nand U25042 (N_25042,N_22599,N_22929);
nor U25043 (N_25043,N_24339,N_20090);
xor U25044 (N_25044,N_23011,N_23327);
nor U25045 (N_25045,N_20453,N_22645);
and U25046 (N_25046,N_22041,N_23963);
or U25047 (N_25047,N_24763,N_21029);
nand U25048 (N_25048,N_20779,N_22486);
nand U25049 (N_25049,N_23217,N_20864);
xor U25050 (N_25050,N_21352,N_20848);
nand U25051 (N_25051,N_20466,N_22828);
and U25052 (N_25052,N_20268,N_20824);
and U25053 (N_25053,N_22606,N_22611);
nand U25054 (N_25054,N_23650,N_22814);
nor U25055 (N_25055,N_22467,N_20524);
nor U25056 (N_25056,N_21039,N_22781);
xnor U25057 (N_25057,N_20762,N_24477);
or U25058 (N_25058,N_22621,N_20623);
nor U25059 (N_25059,N_22261,N_23039);
nand U25060 (N_25060,N_23959,N_24300);
and U25061 (N_25061,N_21904,N_24152);
or U25062 (N_25062,N_23960,N_20222);
nor U25063 (N_25063,N_20121,N_20248);
or U25064 (N_25064,N_22080,N_21895);
and U25065 (N_25065,N_22332,N_24245);
nand U25066 (N_25066,N_21080,N_24635);
nand U25067 (N_25067,N_22343,N_21826);
xor U25068 (N_25068,N_21510,N_22089);
and U25069 (N_25069,N_20674,N_22048);
nor U25070 (N_25070,N_20479,N_24175);
or U25071 (N_25071,N_22040,N_20252);
nand U25072 (N_25072,N_20083,N_22160);
nor U25073 (N_25073,N_21047,N_20744);
xor U25074 (N_25074,N_24968,N_21279);
nor U25075 (N_25075,N_23416,N_24157);
or U25076 (N_25076,N_24159,N_20782);
and U25077 (N_25077,N_21357,N_24484);
xnor U25078 (N_25078,N_20423,N_23883);
nor U25079 (N_25079,N_21022,N_22030);
nand U25080 (N_25080,N_24643,N_22029);
and U25081 (N_25081,N_24215,N_20814);
or U25082 (N_25082,N_20509,N_24323);
and U25083 (N_25083,N_22151,N_20442);
xor U25084 (N_25084,N_23675,N_24609);
nand U25085 (N_25085,N_23103,N_23172);
and U25086 (N_25086,N_23350,N_21052);
or U25087 (N_25087,N_24564,N_24324);
and U25088 (N_25088,N_24318,N_22171);
and U25089 (N_25089,N_23474,N_21833);
and U25090 (N_25090,N_20783,N_24584);
xnor U25091 (N_25091,N_22974,N_21564);
or U25092 (N_25092,N_20520,N_24751);
nor U25093 (N_25093,N_20743,N_24040);
and U25094 (N_25094,N_23091,N_20703);
nand U25095 (N_25095,N_23244,N_21554);
xnor U25096 (N_25096,N_20660,N_21944);
or U25097 (N_25097,N_24512,N_23588);
xor U25098 (N_25098,N_21553,N_24450);
or U25099 (N_25099,N_24641,N_22386);
xor U25100 (N_25100,N_24123,N_20195);
nor U25101 (N_25101,N_22414,N_20209);
xor U25102 (N_25102,N_24954,N_20335);
nor U25103 (N_25103,N_23578,N_21199);
nand U25104 (N_25104,N_20649,N_24464);
xnor U25105 (N_25105,N_24741,N_22627);
nand U25106 (N_25106,N_24991,N_22843);
or U25107 (N_25107,N_20030,N_23660);
nand U25108 (N_25108,N_21577,N_20294);
or U25109 (N_25109,N_21429,N_23053);
nand U25110 (N_25110,N_21433,N_22805);
xor U25111 (N_25111,N_20568,N_20351);
or U25112 (N_25112,N_21410,N_20273);
nand U25113 (N_25113,N_24335,N_20013);
nor U25114 (N_25114,N_20019,N_22802);
or U25115 (N_25115,N_24349,N_22218);
xor U25116 (N_25116,N_23750,N_24574);
nand U25117 (N_25117,N_22406,N_22537);
nand U25118 (N_25118,N_24171,N_23526);
or U25119 (N_25119,N_20807,N_20684);
and U25120 (N_25120,N_22765,N_23107);
nor U25121 (N_25121,N_21097,N_21445);
and U25122 (N_25122,N_21846,N_22310);
or U25123 (N_25123,N_22842,N_23223);
xor U25124 (N_25124,N_22348,N_23191);
xnor U25125 (N_25125,N_20656,N_23468);
nor U25126 (N_25126,N_20203,N_24458);
nand U25127 (N_25127,N_20915,N_23569);
nor U25128 (N_25128,N_22717,N_20735);
and U25129 (N_25129,N_23098,N_23171);
and U25130 (N_25130,N_21658,N_20666);
nor U25131 (N_25131,N_22932,N_24727);
nand U25132 (N_25132,N_20866,N_24983);
or U25133 (N_25133,N_20282,N_22921);
and U25134 (N_25134,N_22439,N_20455);
nor U25135 (N_25135,N_22838,N_23269);
xnor U25136 (N_25136,N_24317,N_22540);
nor U25137 (N_25137,N_21837,N_24939);
and U25138 (N_25138,N_20820,N_24435);
xor U25139 (N_25139,N_21398,N_24193);
xor U25140 (N_25140,N_24481,N_21691);
or U25141 (N_25141,N_22973,N_24679);
nor U25142 (N_25142,N_22356,N_21803);
and U25143 (N_25143,N_22416,N_24439);
xnor U25144 (N_25144,N_23980,N_21479);
or U25145 (N_25145,N_22259,N_24720);
xnor U25146 (N_25146,N_22472,N_24253);
xor U25147 (N_25147,N_24006,N_23558);
xor U25148 (N_25148,N_23900,N_22474);
and U25149 (N_25149,N_21382,N_22679);
nand U25150 (N_25150,N_22980,N_22329);
and U25151 (N_25151,N_20211,N_20719);
xor U25152 (N_25152,N_22544,N_23934);
xnor U25153 (N_25153,N_22039,N_23167);
nand U25154 (N_25154,N_21105,N_24996);
and U25155 (N_25155,N_20596,N_23168);
and U25156 (N_25156,N_23078,N_20150);
xnor U25157 (N_25157,N_20132,N_21633);
or U25158 (N_25158,N_22168,N_24614);
xor U25159 (N_25159,N_20122,N_24091);
nand U25160 (N_25160,N_24242,N_24347);
xnor U25161 (N_25161,N_23469,N_20078);
nand U25162 (N_25162,N_20522,N_23631);
nand U25163 (N_25163,N_22588,N_23953);
nor U25164 (N_25164,N_21346,N_23337);
xnor U25165 (N_25165,N_22668,N_21967);
nand U25166 (N_25166,N_21061,N_22661);
nand U25167 (N_25167,N_23236,N_24148);
xor U25168 (N_25168,N_24408,N_23164);
nand U25169 (N_25169,N_22441,N_24849);
nand U25170 (N_25170,N_24912,N_24921);
nor U25171 (N_25171,N_24674,N_22804);
or U25172 (N_25172,N_22268,N_23728);
or U25173 (N_25173,N_20004,N_23289);
and U25174 (N_25174,N_20134,N_20514);
nor U25175 (N_25175,N_21348,N_20289);
xor U25176 (N_25176,N_24548,N_24831);
nand U25177 (N_25177,N_23245,N_21465);
xnor U25178 (N_25178,N_24438,N_21931);
or U25179 (N_25179,N_22004,N_24892);
xor U25180 (N_25180,N_23067,N_22159);
and U25181 (N_25181,N_24361,N_24087);
nor U25182 (N_25182,N_22622,N_21857);
xnor U25183 (N_25183,N_24287,N_23060);
or U25184 (N_25184,N_22714,N_23659);
or U25185 (N_25185,N_22702,N_21014);
xnor U25186 (N_25186,N_20686,N_21372);
and U25187 (N_25187,N_23476,N_21184);
and U25188 (N_25188,N_20699,N_22641);
nand U25189 (N_25189,N_21159,N_21471);
or U25190 (N_25190,N_24841,N_22150);
and U25191 (N_25191,N_20680,N_24448);
or U25192 (N_25192,N_24493,N_24172);
nor U25193 (N_25193,N_20859,N_22629);
and U25194 (N_25194,N_22423,N_22610);
or U25195 (N_25195,N_22002,N_20067);
and U25196 (N_25196,N_23777,N_23919);
nor U25197 (N_25197,N_24305,N_21792);
xor U25198 (N_25198,N_24688,N_20549);
nand U25199 (N_25199,N_21870,N_24441);
nand U25200 (N_25200,N_21661,N_20233);
or U25201 (N_25201,N_23707,N_21458);
xnor U25202 (N_25202,N_20652,N_21472);
and U25203 (N_25203,N_22947,N_21683);
xor U25204 (N_25204,N_24090,N_22945);
and U25205 (N_25205,N_22255,N_23910);
and U25206 (N_25206,N_21729,N_20169);
nor U25207 (N_25207,N_23681,N_24829);
nor U25208 (N_25208,N_22164,N_24001);
xnor U25209 (N_25209,N_20764,N_21981);
or U25210 (N_25210,N_23853,N_22407);
nand U25211 (N_25211,N_23366,N_24116);
xnor U25212 (N_25212,N_24330,N_21293);
nand U25213 (N_25213,N_20749,N_21524);
nor U25214 (N_25214,N_23694,N_21761);
nor U25215 (N_25215,N_23930,N_21893);
nor U25216 (N_25216,N_22354,N_21140);
nor U25217 (N_25217,N_23291,N_23979);
and U25218 (N_25218,N_23705,N_21541);
nand U25219 (N_25219,N_23874,N_21274);
nor U25220 (N_25220,N_20197,N_22927);
nand U25221 (N_25221,N_24633,N_24234);
or U25222 (N_25222,N_23412,N_24186);
and U25223 (N_25223,N_22018,N_24197);
nand U25224 (N_25224,N_22716,N_23518);
or U25225 (N_25225,N_21982,N_20531);
xnor U25226 (N_25226,N_24748,N_22013);
nor U25227 (N_25227,N_22052,N_22235);
nand U25228 (N_25228,N_20658,N_20357);
nand U25229 (N_25229,N_24813,N_23991);
and U25230 (N_25230,N_24025,N_22491);
and U25231 (N_25231,N_21273,N_22938);
nor U25232 (N_25232,N_24079,N_24073);
nor U25233 (N_25233,N_23006,N_24124);
xor U25234 (N_25234,N_23297,N_24350);
nor U25235 (N_25235,N_23523,N_20044);
nand U25236 (N_25236,N_20785,N_20109);
nand U25237 (N_25237,N_23741,N_23886);
and U25238 (N_25238,N_22788,N_20627);
nor U25239 (N_25239,N_22459,N_20712);
and U25240 (N_25240,N_21209,N_22667);
and U25241 (N_25241,N_23003,N_21071);
and U25242 (N_25242,N_21839,N_21180);
or U25243 (N_25243,N_24729,N_22025);
nor U25244 (N_25244,N_24104,N_22446);
nor U25245 (N_25245,N_21501,N_22819);
nand U25246 (N_25246,N_20042,N_20281);
nand U25247 (N_25247,N_24292,N_22107);
and U25248 (N_25248,N_23386,N_20962);
nand U25249 (N_25249,N_22353,N_24606);
nand U25250 (N_25250,N_24936,N_21587);
and U25251 (N_25251,N_20668,N_20716);
nor U25252 (N_25252,N_21758,N_22922);
and U25253 (N_25253,N_22597,N_24065);
xnor U25254 (N_25254,N_23661,N_20733);
nand U25255 (N_25255,N_21696,N_22291);
xor U25256 (N_25256,N_22670,N_22122);
or U25257 (N_25257,N_22460,N_23633);
nor U25258 (N_25258,N_24012,N_21092);
nand U25259 (N_25259,N_23068,N_23996);
or U25260 (N_25260,N_23725,N_21546);
and U25261 (N_25261,N_21918,N_24738);
or U25262 (N_25262,N_23671,N_20945);
or U25263 (N_25263,N_23268,N_23485);
xor U25264 (N_25264,N_22120,N_22241);
nand U25265 (N_25265,N_21930,N_24084);
xor U25266 (N_25266,N_24691,N_22663);
and U25267 (N_25267,N_21131,N_22444);
or U25268 (N_25268,N_24033,N_21225);
or U25269 (N_25269,N_24610,N_21389);
xnor U25270 (N_25270,N_21772,N_23112);
nor U25271 (N_25271,N_23057,N_21584);
and U25272 (N_25272,N_22276,N_22596);
nor U25273 (N_25273,N_20934,N_21778);
nand U25274 (N_25274,N_21394,N_21948);
or U25275 (N_25275,N_22345,N_22834);
nand U25276 (N_25276,N_24999,N_24074);
xnor U25277 (N_25277,N_24655,N_21597);
nand U25278 (N_25278,N_21117,N_23530);
xnor U25279 (N_25279,N_24102,N_20539);
xnor U25280 (N_25280,N_24961,N_23494);
nand U25281 (N_25281,N_21639,N_23888);
or U25282 (N_25282,N_23463,N_21521);
nor U25283 (N_25283,N_20626,N_21093);
xnor U25284 (N_25284,N_22427,N_20752);
and U25285 (N_25285,N_22761,N_24900);
xor U25286 (N_25286,N_22361,N_23591);
nand U25287 (N_25287,N_24836,N_22735);
nand U25288 (N_25288,N_22698,N_22121);
nand U25289 (N_25289,N_20170,N_21203);
nand U25290 (N_25290,N_24583,N_21721);
xnor U25291 (N_25291,N_21886,N_23737);
or U25292 (N_25292,N_24495,N_23047);
xor U25293 (N_25293,N_23403,N_21237);
or U25294 (N_25294,N_24931,N_22127);
and U25295 (N_25295,N_21783,N_20550);
nor U25296 (N_25296,N_20307,N_23389);
nand U25297 (N_25297,N_24334,N_22538);
xnor U25298 (N_25298,N_22650,N_22779);
nand U25299 (N_25299,N_21387,N_22986);
or U25300 (N_25300,N_22753,N_22078);
or U25301 (N_25301,N_23013,N_20465);
nand U25302 (N_25302,N_24711,N_22910);
xnor U25303 (N_25303,N_21636,N_23148);
nor U25304 (N_25304,N_20165,N_23839);
and U25305 (N_25305,N_20299,N_23879);
xnor U25306 (N_25306,N_21135,N_23449);
nor U25307 (N_25307,N_24331,N_21088);
and U25308 (N_25308,N_21077,N_24953);
nand U25309 (N_25309,N_23108,N_23473);
xnor U25310 (N_25310,N_20430,N_23880);
nor U25311 (N_25311,N_21120,N_24206);
xor U25312 (N_25312,N_20481,N_20742);
xnor U25313 (N_25313,N_20504,N_20841);
nor U25314 (N_25314,N_24558,N_20471);
xor U25315 (N_25315,N_24018,N_23678);
xnor U25316 (N_25316,N_22939,N_22950);
and U25317 (N_25317,N_21303,N_24381);
nor U25318 (N_25318,N_21867,N_21017);
nand U25319 (N_25319,N_23308,N_24935);
nor U25320 (N_25320,N_23362,N_22520);
xnor U25321 (N_25321,N_24756,N_24276);
nor U25322 (N_25322,N_23890,N_23165);
nand U25323 (N_25323,N_23064,N_22585);
or U25324 (N_25324,N_23495,N_23752);
nand U25325 (N_25325,N_20376,N_20646);
nand U25326 (N_25326,N_24718,N_20208);
xor U25327 (N_25327,N_22536,N_21208);
nor U25328 (N_25328,N_20932,N_24375);
nand U25329 (N_25329,N_21216,N_24250);
nand U25330 (N_25330,N_22971,N_23797);
or U25331 (N_25331,N_22614,N_21064);
or U25332 (N_25332,N_21058,N_23851);
xor U25333 (N_25333,N_22638,N_20336);
nor U25334 (N_25334,N_22415,N_22059);
or U25335 (N_25335,N_22174,N_22082);
or U25336 (N_25336,N_20055,N_21278);
or U25337 (N_25337,N_22914,N_23998);
xnor U25338 (N_25338,N_21828,N_22857);
and U25339 (N_25339,N_23351,N_22706);
or U25340 (N_25340,N_20464,N_21298);
and U25341 (N_25341,N_23400,N_20914);
and U25342 (N_25342,N_20768,N_21333);
nand U25343 (N_25343,N_21155,N_21157);
xor U25344 (N_25344,N_22675,N_23524);
nor U25345 (N_25345,N_21320,N_21438);
xnor U25346 (N_25346,N_21046,N_23312);
nand U25347 (N_25347,N_23342,N_22820);
and U25348 (N_25348,N_24274,N_20757);
xor U25349 (N_25349,N_22870,N_20463);
or U25350 (N_25350,N_23535,N_21724);
nand U25351 (N_25351,N_20799,N_21752);
and U25352 (N_25352,N_20959,N_24780);
nand U25353 (N_25353,N_21879,N_20338);
or U25354 (N_25354,N_20535,N_21032);
xor U25355 (N_25355,N_20979,N_21201);
or U25356 (N_25356,N_23085,N_20234);
nand U25357 (N_25357,N_21789,N_20189);
and U25358 (N_25358,N_21884,N_24218);
xnor U25359 (N_25359,N_22649,N_21376);
or U25360 (N_25360,N_21625,N_23527);
nor U25361 (N_25361,N_22877,N_22222);
nor U25362 (N_25362,N_22823,N_22286);
or U25363 (N_25363,N_22132,N_23136);
and U25364 (N_25364,N_24951,N_22336);
or U25365 (N_25365,N_21858,N_22024);
xnor U25366 (N_25366,N_24184,N_21367);
xnor U25367 (N_25367,N_20889,N_21455);
xor U25368 (N_25368,N_20918,N_24007);
and U25369 (N_25369,N_20987,N_22527);
nor U25370 (N_25370,N_22841,N_22426);
and U25371 (N_25371,N_23071,N_21243);
or U25372 (N_25372,N_24766,N_23153);
nor U25373 (N_25373,N_21806,N_24835);
or U25374 (N_25374,N_22253,N_21171);
and U25375 (N_25375,N_22751,N_20451);
and U25376 (N_25376,N_21233,N_24115);
or U25377 (N_25377,N_24008,N_23932);
nand U25378 (N_25378,N_24264,N_23477);
or U25379 (N_25379,N_21463,N_23490);
or U25380 (N_25380,N_22135,N_21748);
nor U25381 (N_25381,N_21812,N_23027);
or U25382 (N_25382,N_20232,N_21148);
nor U25383 (N_25383,N_23509,N_23925);
or U25384 (N_25384,N_23307,N_20500);
nor U25385 (N_25385,N_20781,N_24907);
nor U25386 (N_25386,N_22274,N_24267);
xor U25387 (N_25387,N_20425,N_22478);
nand U25388 (N_25388,N_21666,N_21145);
nand U25389 (N_25389,N_24733,N_24386);
or U25390 (N_25390,N_21128,N_21414);
nand U25391 (N_25391,N_24686,N_20225);
nand U25392 (N_25392,N_20198,N_24830);
xor U25393 (N_25393,N_22434,N_23697);
xnor U25394 (N_25394,N_24340,N_23024);
and U25395 (N_25395,N_24265,N_20727);
nor U25396 (N_25396,N_22287,N_22840);
nor U25397 (N_25397,N_22170,N_23882);
or U25398 (N_25398,N_24745,N_21673);
or U25399 (N_25399,N_22110,N_23134);
or U25400 (N_25400,N_21503,N_23042);
nor U25401 (N_25401,N_22143,N_20943);
nand U25402 (N_25402,N_22999,N_22505);
or U25403 (N_25403,N_23332,N_24731);
and U25404 (N_25404,N_20912,N_23231);
nand U25405 (N_25405,N_24322,N_20851);
nand U25406 (N_25406,N_23138,N_22182);
nand U25407 (N_25407,N_24112,N_24811);
nor U25408 (N_25408,N_24979,N_24129);
or U25409 (N_25409,N_22352,N_21063);
xor U25410 (N_25410,N_24035,N_21449);
and U25411 (N_25411,N_20245,N_20310);
and U25412 (N_25412,N_24522,N_21759);
xor U25413 (N_25413,N_23277,N_24544);
nor U25414 (N_25414,N_24857,N_23966);
nand U25415 (N_25415,N_24950,N_23313);
and U25416 (N_25416,N_23314,N_20045);
and U25417 (N_25417,N_20958,N_20809);
xnor U25418 (N_25418,N_21589,N_20893);
or U25419 (N_25419,N_24158,N_23109);
xnor U25420 (N_25420,N_21112,N_24149);
nor U25421 (N_25421,N_20216,N_23347);
and U25422 (N_25422,N_21207,N_20720);
nor U25423 (N_25423,N_23620,N_21821);
nand U25424 (N_25424,N_23607,N_24572);
and U25425 (N_25425,N_24409,N_22126);
and U25426 (N_25426,N_20828,N_24378);
xnor U25427 (N_25427,N_24949,N_24778);
and U25428 (N_25428,N_24794,N_23118);
xor U25429 (N_25429,N_20012,N_22951);
or U25430 (N_25430,N_21409,N_20382);
xor U25431 (N_25431,N_21249,N_24213);
and U25432 (N_25432,N_22115,N_24325);
and U25433 (N_25433,N_23410,N_23461);
nand U25434 (N_25434,N_23499,N_20347);
and U25435 (N_25435,N_23912,N_21785);
nor U25436 (N_25436,N_24861,N_21775);
or U25437 (N_25437,N_20598,N_22607);
xnor U25438 (N_25438,N_23634,N_21626);
nand U25439 (N_25439,N_21280,N_23187);
or U25440 (N_25440,N_22000,N_20869);
nor U25441 (N_25441,N_23363,N_21880);
xor U25442 (N_25442,N_21989,N_23427);
and U25443 (N_25443,N_24487,N_24314);
nand U25444 (N_25444,N_24556,N_22315);
or U25445 (N_25445,N_21642,N_20452);
or U25446 (N_25446,N_22600,N_24454);
xnor U25447 (N_25447,N_23713,N_21646);
and U25448 (N_25448,N_24881,N_22769);
and U25449 (N_25449,N_20988,N_23050);
nand U25450 (N_25450,N_21798,N_21688);
nand U25451 (N_25451,N_20591,N_23529);
xor U25452 (N_25452,N_20502,N_21481);
xor U25453 (N_25453,N_22424,N_23593);
nor U25454 (N_25454,N_22017,N_22892);
or U25455 (N_25455,N_22007,N_20570);
or U25456 (N_25456,N_23087,N_24475);
xnor U25457 (N_25457,N_22412,N_20131);
and U25458 (N_25458,N_23937,N_24472);
xor U25459 (N_25459,N_20576,N_21245);
nor U25460 (N_25460,N_24480,N_21255);
or U25461 (N_25461,N_23316,N_22992);
nor U25462 (N_25462,N_20533,N_23311);
nand U25463 (N_25463,N_20256,N_20717);
or U25464 (N_25464,N_22443,N_24622);
nand U25465 (N_25465,N_23947,N_22032);
xor U25466 (N_25466,N_20552,N_24747);
and U25467 (N_25467,N_23398,N_20883);
or U25468 (N_25468,N_20790,N_23293);
or U25469 (N_25469,N_20283,N_20021);
or U25470 (N_25470,N_20534,N_23160);
and U25471 (N_25471,N_22382,N_22758);
and U25472 (N_25472,N_24787,N_22789);
or U25473 (N_25473,N_21268,N_21907);
nor U25474 (N_25474,N_23765,N_24737);
and U25475 (N_25475,N_23026,N_20542);
and U25476 (N_25476,N_24395,N_23695);
xnor U25477 (N_25477,N_22481,N_24915);
nand U25478 (N_25478,N_22379,N_21733);
nor U25479 (N_25479,N_24382,N_23667);
and U25480 (N_25480,N_23318,N_20949);
nor U25481 (N_25481,N_24138,N_21277);
nor U25482 (N_25482,N_20194,N_24848);
xnor U25483 (N_25483,N_20243,N_22764);
and U25484 (N_25484,N_23715,N_23417);
nand U25485 (N_25485,N_24078,N_24886);
or U25486 (N_25486,N_24677,N_20476);
nand U25487 (N_25487,N_22550,N_22366);
and U25488 (N_25488,N_24355,N_20578);
nand U25489 (N_25489,N_23982,N_21594);
nand U25490 (N_25490,N_22846,N_23864);
xor U25491 (N_25491,N_23799,N_20951);
and U25492 (N_25492,N_22799,N_21330);
nor U25493 (N_25493,N_20886,N_20345);
and U25494 (N_25494,N_20844,N_20997);
and U25495 (N_25495,N_21345,N_23163);
xnor U25496 (N_25496,N_24183,N_24771);
or U25497 (N_25497,N_22866,N_20415);
nand U25498 (N_25498,N_24427,N_24966);
or U25499 (N_25499,N_21637,N_22507);
nor U25500 (N_25500,N_24095,N_23724);
nor U25501 (N_25501,N_20868,N_23653);
xnor U25502 (N_25502,N_24919,N_21055);
nand U25503 (N_25503,N_24161,N_21911);
xnor U25504 (N_25504,N_24866,N_23969);
xor U25505 (N_25505,N_21364,N_23114);
and U25506 (N_25506,N_20188,N_23748);
nand U25507 (N_25507,N_23742,N_21321);
nor U25508 (N_25508,N_20919,N_24496);
nor U25509 (N_25509,N_23747,N_22496);
and U25510 (N_25510,N_21335,N_23128);
nor U25511 (N_25511,N_20125,N_21177);
xor U25512 (N_25512,N_20220,N_21275);
nand U25513 (N_25513,N_21158,N_24582);
nand U25514 (N_25514,N_21413,N_22177);
nand U25515 (N_25515,N_22749,N_23137);
or U25516 (N_25516,N_22050,N_23823);
nand U25517 (N_25517,N_21189,N_20100);
nor U25518 (N_25518,N_20571,N_21906);
xnor U25519 (N_25519,N_20334,N_22238);
and U25520 (N_25520,N_20101,N_21254);
nor U25521 (N_25521,N_23708,N_20025);
nor U25522 (N_25522,N_23072,N_20892);
nand U25523 (N_25523,N_24401,N_22236);
xor U25524 (N_25524,N_21315,N_21466);
xnor U25525 (N_25525,N_21992,N_20532);
xnor U25526 (N_25526,N_22296,N_24639);
or U25527 (N_25527,N_20510,N_22557);
nand U25528 (N_25528,N_24905,N_23699);
xor U25529 (N_25529,N_20728,N_23986);
or U25530 (N_25530,N_21439,N_21874);
and U25531 (N_25531,N_24880,N_24390);
and U25532 (N_25532,N_21025,N_24793);
xor U25533 (N_25533,N_23958,N_20607);
or U25534 (N_25534,N_21197,N_24177);
or U25535 (N_25535,N_20096,N_23286);
xor U25536 (N_25536,N_23792,N_21072);
xor U25537 (N_25537,N_22806,N_23331);
or U25538 (N_25538,N_23333,N_22699);
nor U25539 (N_25539,N_22608,N_21995);
and U25540 (N_25540,N_24597,N_24667);
nor U25541 (N_25541,N_22239,N_22162);
nand U25542 (N_25542,N_24734,N_22221);
or U25543 (N_25543,N_24970,N_22399);
or U25544 (N_25544,N_21818,N_20050);
nor U25545 (N_25545,N_20745,N_24687);
nand U25546 (N_25546,N_24897,N_22413);
nor U25547 (N_25547,N_22755,N_20046);
xor U25548 (N_25548,N_22376,N_21917);
nor U25549 (N_25549,N_22346,N_21523);
or U25550 (N_25550,N_21400,N_21574);
and U25551 (N_25551,N_21332,N_22319);
xnor U25552 (N_25552,N_22955,N_21825);
xnor U25553 (N_25553,N_20274,N_22726);
nand U25554 (N_25554,N_22700,N_20881);
nand U25555 (N_25555,N_20265,N_21687);
nor U25556 (N_25556,N_22049,N_20996);
nor U25557 (N_25557,N_23406,N_24060);
xor U25558 (N_25558,N_23525,N_24712);
nand U25559 (N_25559,N_22995,N_21246);
and U25560 (N_25560,N_24963,N_24773);
nor U25561 (N_25561,N_21485,N_20141);
or U25562 (N_25562,N_23238,N_24110);
nand U25563 (N_25563,N_21202,N_24945);
and U25564 (N_25564,N_22652,N_23288);
xor U25565 (N_25565,N_23428,N_24997);
or U25566 (N_25566,N_22118,N_21460);
nand U25567 (N_25567,N_23687,N_21425);
or U25568 (N_25568,N_21557,N_20405);
or U25569 (N_25569,N_21099,N_22117);
nand U25570 (N_25570,N_23536,N_21605);
nand U25571 (N_25571,N_22915,N_21955);
nor U25572 (N_25572,N_24136,N_23920);
and U25573 (N_25573,N_24107,N_20346);
and U25574 (N_25574,N_21305,N_22707);
and U25575 (N_25575,N_20173,N_24094);
nor U25576 (N_25576,N_20406,N_22831);
nand U25577 (N_25577,N_21669,N_23329);
nand U25578 (N_25578,N_23898,N_20672);
xnor U25579 (N_25579,N_24089,N_23604);
nor U25580 (N_25580,N_20483,N_23145);
or U25581 (N_25581,N_24590,N_21634);
nand U25582 (N_25582,N_20434,N_23957);
xnor U25583 (N_25583,N_21736,N_20032);
xor U25584 (N_25584,N_22223,N_24550);
nor U25585 (N_25585,N_22084,N_22473);
nand U25586 (N_25586,N_23938,N_21599);
and U25587 (N_25587,N_21535,N_22669);
and U25588 (N_25588,N_20495,N_22494);
nand U25589 (N_25589,N_24993,N_21373);
and U25590 (N_25590,N_23967,N_20595);
nor U25591 (N_25591,N_20091,N_21272);
nor U25592 (N_25592,N_22617,N_20624);
and U25593 (N_25593,N_20037,N_20142);
nor U25594 (N_25594,N_23444,N_22777);
nor U25595 (N_25595,N_22832,N_24329);
nand U25596 (N_25596,N_21657,N_21901);
or U25597 (N_25597,N_20813,N_24150);
or U25598 (N_25598,N_24432,N_24166);
and U25599 (N_25599,N_23646,N_23935);
xnor U25600 (N_25600,N_23868,N_21390);
nand U25601 (N_25601,N_20136,N_24598);
nor U25602 (N_25602,N_20352,N_20592);
xnor U25603 (N_25603,N_22155,N_23405);
nand U25604 (N_25604,N_20810,N_20836);
nand U25605 (N_25605,N_22175,N_24918);
nand U25606 (N_25606,N_21218,N_20072);
nor U25607 (N_25607,N_21889,N_21675);
nor U25608 (N_25608,N_23364,N_21814);
nand U25609 (N_25609,N_22605,N_21533);
or U25610 (N_25610,N_21452,N_22207);
and U25611 (N_25611,N_21572,N_23115);
and U25612 (N_25612,N_22521,N_23790);
nor U25613 (N_25613,N_20437,N_24601);
nor U25614 (N_25614,N_24865,N_22728);
or U25615 (N_25615,N_23774,N_23788);
xnor U25616 (N_25616,N_22598,N_24372);
xnor U25617 (N_25617,N_23349,N_23704);
xor U25618 (N_25618,N_23896,N_21746);
nor U25619 (N_25619,N_21222,N_23856);
nor U25620 (N_25620,N_24587,N_23784);
and U25621 (N_25621,N_24821,N_23306);
xor U25622 (N_25622,N_20020,N_24732);
nand U25623 (N_25623,N_20312,N_24876);
xor U25624 (N_25624,N_24578,N_22784);
nand U25625 (N_25625,N_24194,N_21979);
nand U25626 (N_25626,N_21037,N_24579);
xnor U25627 (N_25627,N_22658,N_21888);
nand U25628 (N_25628,N_24410,N_22936);
and U25629 (N_25629,N_21484,N_22066);
nand U25630 (N_25630,N_23122,N_23968);
and U25631 (N_25631,N_21835,N_20654);
and U25632 (N_25632,N_24055,N_21427);
nand U25633 (N_25633,N_22229,N_21604);
nor U25634 (N_25634,N_22429,N_20725);
nor U25635 (N_25635,N_21779,N_23298);
and U25636 (N_25636,N_24246,N_22815);
xor U25637 (N_25637,N_20454,N_24283);
or U25638 (N_25638,N_24470,N_22906);
xnor U25639 (N_25639,N_23339,N_20073);
nor U25640 (N_25640,N_22519,N_21507);
or U25641 (N_25641,N_23436,N_22584);
nand U25642 (N_25642,N_24806,N_20916);
xnor U25643 (N_25643,N_24229,N_21684);
or U25644 (N_25644,N_22737,N_21693);
nand U25645 (N_25645,N_20818,N_20564);
or U25646 (N_25646,N_24217,N_22033);
and U25647 (N_25647,N_22360,N_23645);
or U25648 (N_25648,N_22514,N_21491);
xor U25649 (N_25649,N_22859,N_24877);
and U25650 (N_25650,N_21469,N_22067);
nor U25651 (N_25651,N_24675,N_23891);
nor U25652 (N_25652,N_23345,N_20158);
nor U25653 (N_25653,N_24934,N_23677);
nand U25654 (N_25654,N_22580,N_23548);
nand U25655 (N_25655,N_24155,N_21059);
or U25656 (N_25656,N_24998,N_21057);
or U25657 (N_25657,N_23305,N_21545);
and U25658 (N_25658,N_23189,N_20760);
or U25659 (N_25659,N_21424,N_20388);
and U25660 (N_25660,N_21436,N_24948);
xnor U25661 (N_25661,N_22047,N_21861);
nor U25662 (N_25662,N_20400,N_24088);
xor U25663 (N_25663,N_20877,N_22742);
xor U25664 (N_25664,N_24910,N_20984);
nand U25665 (N_25665,N_22477,N_21864);
or U25666 (N_25666,N_22586,N_20961);
nand U25667 (N_25667,N_22108,N_20651);
nor U25668 (N_25668,N_22498,N_23544);
nand U25669 (N_25669,N_20171,N_21635);
nor U25670 (N_25670,N_22185,N_23772);
or U25671 (N_25671,N_20385,N_24266);
nand U25672 (N_25672,N_20315,N_20373);
nor U25673 (N_25673,N_24297,N_21614);
or U25674 (N_25674,N_22208,N_20431);
or U25675 (N_25675,N_23599,N_20348);
or U25676 (N_25676,N_24986,N_22776);
nand U25677 (N_25677,N_22458,N_21978);
xor U25678 (N_25678,N_21877,N_23041);
and U25679 (N_25679,N_21717,N_20035);
and U25680 (N_25680,N_20196,N_24642);
nand U25681 (N_25681,N_23034,N_21502);
and U25682 (N_25682,N_23266,N_24781);
xnor U25683 (N_25683,N_20829,N_24977);
and U25684 (N_25684,N_23557,N_23387);
and U25685 (N_25685,N_20600,N_21716);
or U25686 (N_25686,N_24357,N_24559);
or U25687 (N_25687,N_22430,N_20456);
or U25688 (N_25688,N_24384,N_23804);
nand U25689 (N_25689,N_22723,N_22263);
nor U25690 (N_25690,N_20292,N_22060);
xnor U25691 (N_25691,N_24249,N_20512);
xor U25692 (N_25692,N_21020,N_23721);
or U25693 (N_25693,N_24044,N_22901);
xor U25694 (N_25694,N_21797,N_23922);
nand U25695 (N_25695,N_24988,N_24839);
nand U25696 (N_25696,N_22464,N_22368);
or U25697 (N_25697,N_21450,N_22940);
and U25698 (N_25698,N_23690,N_22398);
xnor U25699 (N_25699,N_20432,N_20908);
nand U25700 (N_25700,N_24086,N_20342);
or U25701 (N_25701,N_21896,N_23185);
and U25702 (N_25702,N_20236,N_20705);
xor U25703 (N_25703,N_23271,N_21534);
nor U25704 (N_25704,N_21704,N_23287);
nor U25705 (N_25705,N_20677,N_21961);
nand U25706 (N_25706,N_24746,N_22076);
nor U25707 (N_25707,N_24535,N_24833);
nor U25708 (N_25708,N_20606,N_24510);
nor U25709 (N_25709,N_23512,N_20257);
nor U25710 (N_25710,N_22988,N_20832);
nand U25711 (N_25711,N_21292,N_21920);
or U25712 (N_25712,N_23394,N_24453);
nand U25713 (N_25713,N_21568,N_21187);
xor U25714 (N_25714,N_20427,N_24623);
nand U25715 (N_25715,N_23744,N_24987);
nand U25716 (N_25716,N_24165,N_22845);
or U25717 (N_25717,N_24519,N_23421);
xnor U25718 (N_25718,N_22113,N_24809);
nand U25719 (N_25719,N_22576,N_24776);
nand U25720 (N_25720,N_20748,N_20264);
or U25721 (N_25721,N_21926,N_20350);
and U25722 (N_25722,N_23388,N_23626);
xor U25723 (N_25723,N_24269,N_24626);
nor U25724 (N_25724,N_20602,N_24093);
nor U25725 (N_25725,N_24288,N_24671);
nand U25726 (N_25726,N_20931,N_21086);
nand U25727 (N_25727,N_24872,N_20537);
nand U25728 (N_25728,N_22450,N_21513);
nand U25729 (N_25729,N_24651,N_20276);
or U25730 (N_25730,N_22690,N_20137);
and U25731 (N_25731,N_22384,N_21122);
xnor U25732 (N_25732,N_22981,N_24032);
and U25733 (N_25733,N_22463,N_20187);
nand U25734 (N_25734,N_21496,N_24363);
or U25735 (N_25735,N_23105,N_24462);
and U25736 (N_25736,N_22232,N_21543);
nor U25737 (N_25737,N_21663,N_22277);
or U25738 (N_25738,N_23282,N_23508);
or U25739 (N_25739,N_22313,N_21281);
or U25740 (N_25740,N_23423,N_23859);
or U25741 (N_25741,N_22515,N_24491);
nor U25742 (N_25742,N_23740,N_21351);
or U25743 (N_25743,N_20364,N_23944);
xor U25744 (N_25744,N_23070,N_21963);
nand U25745 (N_25745,N_21476,N_20770);
and U25746 (N_25746,N_20138,N_20111);
xor U25747 (N_25747,N_24352,N_23361);
and U25748 (N_25748,N_22740,N_22480);
and U25749 (N_25749,N_24414,N_24588);
nand U25750 (N_25750,N_22837,N_22680);
nand U25751 (N_25751,N_20320,N_21987);
nor U25752 (N_25752,N_24725,N_21654);
or U25753 (N_25753,N_20062,N_21569);
or U25754 (N_25754,N_23005,N_21223);
xor U25755 (N_25755,N_21668,N_24767);
or U25756 (N_25756,N_21876,N_22531);
or U25757 (N_25757,N_23395,N_22744);
and U25758 (N_25758,N_23903,N_23076);
and U25759 (N_25759,N_20487,N_22856);
or U25760 (N_25760,N_20804,N_20443);
and U25761 (N_25761,N_22523,N_23939);
and U25762 (N_25762,N_21464,N_22293);
or U25763 (N_25763,N_24844,N_24705);
xnor U25764 (N_25764,N_21151,N_24168);
and U25765 (N_25765,N_23770,N_21960);
xnor U25766 (N_25766,N_21527,N_23285);
and U25767 (N_25767,N_24273,N_21591);
and U25768 (N_25768,N_21606,N_23767);
and U25769 (N_25769,N_24198,N_20429);
nor U25770 (N_25770,N_22985,N_21794);
and U25771 (N_25771,N_20695,N_23635);
nor U25772 (N_25772,N_22644,N_24290);
nor U25773 (N_25773,N_23895,N_22326);
nor U25774 (N_25774,N_24415,N_21566);
or U25775 (N_25775,N_21347,N_23182);
nand U25776 (N_25776,N_20489,N_21969);
and U25777 (N_25777,N_21252,N_23452);
xor U25778 (N_25778,N_22747,N_24847);
or U25779 (N_25779,N_20477,N_24777);
nor U25780 (N_25780,N_24436,N_21319);
nor U25781 (N_25781,N_24542,N_22305);
nand U25782 (N_25782,N_20146,N_22193);
or U25783 (N_25783,N_20449,N_23296);
nand U25784 (N_25784,N_20152,N_21079);
nor U25785 (N_25785,N_23322,N_20590);
or U25786 (N_25786,N_22085,N_23120);
or U25787 (N_25787,N_23460,N_21475);
or U25788 (N_25788,N_23514,N_20731);
nor U25789 (N_25789,N_24312,N_22686);
or U25790 (N_25790,N_23429,N_23309);
nor U25791 (N_25791,N_21119,N_22511);
nor U25792 (N_25792,N_24471,N_22701);
nand U25793 (N_25793,N_21681,N_21749);
xnor U25794 (N_25794,N_23970,N_23294);
and U25795 (N_25795,N_22219,N_22240);
nand U25796 (N_25796,N_20693,N_22643);
nand U25797 (N_25797,N_21069,N_20667);
and U25798 (N_25798,N_20129,N_20375);
and U25799 (N_25799,N_21068,N_21765);
xor U25800 (N_25800,N_21065,N_23901);
and U25801 (N_25801,N_21488,N_22803);
or U25802 (N_25802,N_23213,N_22215);
and U25803 (N_25803,N_23663,N_21287);
and U25804 (N_25804,N_23280,N_21049);
xor U25805 (N_25805,N_21970,N_20802);
and U25806 (N_25806,N_22388,N_24644);
xor U25807 (N_25807,N_23012,N_21416);
or U25808 (N_25808,N_21498,N_21732);
xor U25809 (N_25809,N_21461,N_23230);
nor U25810 (N_25810,N_23976,N_20337);
xnor U25811 (N_25811,N_24902,N_22785);
nor U25812 (N_25812,N_23572,N_24170);
or U25813 (N_25813,N_23564,N_24875);
xor U25814 (N_25814,N_21537,N_22028);
nor U25815 (N_25815,N_20436,N_23228);
nor U25816 (N_25816,N_23805,N_20501);
and U25817 (N_25817,N_20358,N_21610);
and U25818 (N_25818,N_24659,N_22883);
and U25819 (N_25819,N_24596,N_23139);
xnor U25820 (N_25820,N_20191,N_23325);
nand U25821 (N_25821,N_22405,N_20653);
nand U25822 (N_25822,N_23424,N_21204);
and U25823 (N_25823,N_24070,N_22878);
and U25824 (N_25824,N_22068,N_22546);
xor U25825 (N_25825,N_24960,N_20581);
xnor U25826 (N_25826,N_24920,N_20031);
nor U25827 (N_25827,N_23008,N_21192);
or U25828 (N_25828,N_21824,N_22210);
xor U25829 (N_25829,N_23791,N_20786);
nor U25830 (N_25830,N_21751,N_20861);
or U25831 (N_25831,N_23926,N_24233);
nand U25832 (N_25832,N_24605,N_22228);
xnor U25833 (N_25833,N_22022,N_20784);
or U25834 (N_25834,N_22849,N_22672);
xor U25835 (N_25835,N_23093,N_23124);
and U25836 (N_25836,N_23430,N_21002);
nand U25837 (N_25837,N_23343,N_20144);
or U25838 (N_25838,N_20765,N_20723);
or U25839 (N_25839,N_21738,N_23310);
nand U25840 (N_25840,N_24113,N_20610);
nand U25841 (N_25841,N_24422,N_23978);
and U25842 (N_25842,N_23251,N_24393);
or U25843 (N_25843,N_21181,N_22651);
or U25844 (N_25844,N_24843,N_23043);
xnor U25845 (N_25845,N_20180,N_20970);
or U25846 (N_25846,N_21745,N_20412);
xnor U25847 (N_25847,N_23655,N_20053);
or U25848 (N_25848,N_20605,N_20904);
or U25849 (N_25849,N_20247,N_23181);
nand U25850 (N_25850,N_23570,N_23703);
nor U25851 (N_25851,N_21403,N_24132);
and U25852 (N_25852,N_23489,N_24338);
xor U25853 (N_25853,N_23510,N_23399);
or U25854 (N_25854,N_23739,N_21643);
xor U25855 (N_25855,N_24816,N_22230);
and U25856 (N_25856,N_20326,N_23905);
nand U25857 (N_25857,N_23158,N_20490);
nor U25858 (N_25858,N_23216,N_22023);
nand U25859 (N_25859,N_22709,N_21713);
nor U25860 (N_25860,N_20496,N_22855);
and U25861 (N_25861,N_23573,N_23372);
xnor U25862 (N_25862,N_22960,N_24072);
and U25863 (N_25863,N_22620,N_23861);
and U25864 (N_25864,N_21823,N_20900);
nand U25865 (N_25865,N_22972,N_22389);
xor U25866 (N_25866,N_23256,N_23504);
xnor U25867 (N_25867,N_21051,N_23007);
or U25868 (N_25868,N_22001,N_24299);
nand U25869 (N_25869,N_21822,N_21924);
nor U25870 (N_25870,N_23004,N_22447);
or U25871 (N_25871,N_20049,N_24379);
nand U25872 (N_25872,N_22318,N_21338);
or U25873 (N_25873,N_23571,N_22816);
nand U25874 (N_25874,N_24853,N_20835);
nand U25875 (N_25875,N_23822,N_24726);
xor U25876 (N_25876,N_23205,N_21518);
nand U25877 (N_25877,N_20633,N_23373);
nand U25878 (N_25878,N_24169,N_21897);
or U25879 (N_25879,N_20640,N_20118);
nor U25880 (N_25880,N_22397,N_23899);
nor U25881 (N_25881,N_22504,N_22926);
nand U25882 (N_25882,N_23407,N_24406);
nor U25883 (N_25883,N_20953,N_24666);
nand U25884 (N_25884,N_23380,N_24391);
xnor U25885 (N_25885,N_24735,N_20058);
nor U25886 (N_25886,N_22428,N_20706);
nor U25887 (N_25887,N_20615,N_21299);
and U25888 (N_25888,N_20395,N_20026);
nand U25889 (N_25889,N_21016,N_20788);
nor U25890 (N_25890,N_20638,N_24710);
and U25891 (N_25891,N_23629,N_21082);
nor U25892 (N_25892,N_20011,N_21408);
nor U25893 (N_25893,N_20029,N_21771);
nand U25894 (N_25894,N_21943,N_21121);
xnor U25895 (N_25895,N_20515,N_24566);
xnor U25896 (N_25896,N_21006,N_21698);
and U25897 (N_25897,N_21677,N_21980);
nand U25898 (N_25898,N_21210,N_21608);
and U25899 (N_25899,N_22298,N_21084);
xnor U25900 (N_25900,N_20936,N_21430);
and U25901 (N_25901,N_21103,N_24758);
and U25902 (N_25902,N_20803,N_23802);
nor U25903 (N_25903,N_22502,N_24370);
nand U25904 (N_25904,N_20426,N_22534);
nor U25905 (N_25905,N_22630,N_20819);
nand U25906 (N_25906,N_24698,N_22952);
or U25907 (N_25907,N_24492,N_20461);
and U25908 (N_25908,N_20942,N_23909);
nor U25909 (N_25909,N_22983,N_21848);
xor U25910 (N_25910,N_23401,N_23471);
nor U25911 (N_25911,N_24511,N_21528);
xnor U25912 (N_25912,N_20644,N_24003);
nand U25913 (N_25913,N_21286,N_24156);
nor U25914 (N_25914,N_22351,N_22530);
nor U25915 (N_25915,N_24621,N_21166);
nor U25916 (N_25916,N_22887,N_21490);
xnor U25917 (N_25917,N_22657,N_23020);
nand U25918 (N_25918,N_24887,N_24940);
and U25919 (N_25919,N_20986,N_21609);
xor U25920 (N_25920,N_23063,N_22172);
or U25921 (N_25921,N_21834,N_23334);
nand U25922 (N_25922,N_24790,N_20290);
xor U25923 (N_25923,N_22325,N_22695);
nand U25924 (N_25924,N_24852,N_22595);
xor U25925 (N_25925,N_24135,N_21631);
xnor U25926 (N_25926,N_20616,N_20271);
nand U25927 (N_25927,N_22711,N_20850);
or U25928 (N_25928,N_22205,N_23871);
and U25929 (N_25929,N_24134,N_21762);
and U25930 (N_25930,N_23290,N_21615);
nor U25931 (N_25931,N_23601,N_21130);
or U25932 (N_25932,N_21627,N_20536);
nor U25933 (N_25933,N_20617,N_21482);
and U25934 (N_25934,N_20139,N_24537);
or U25935 (N_25935,N_21005,N_22260);
xor U25936 (N_25936,N_21788,N_21423);
and U25937 (N_25937,N_21250,N_21289);
or U25938 (N_25938,N_21928,N_20751);
xor U25939 (N_25939,N_22136,N_21573);
nor U25940 (N_25940,N_20244,N_22603);
nand U25941 (N_25941,N_20817,N_21392);
xnor U25942 (N_25942,N_22483,N_20905);
or U25943 (N_25943,N_21563,N_21623);
or U25944 (N_25944,N_23132,N_20940);
nand U25945 (N_25945,N_21318,N_22393);
nand U25946 (N_25946,N_20409,N_21457);
or U25947 (N_25947,N_22555,N_23642);
and U25948 (N_25948,N_22809,N_22817);
nor U25949 (N_25949,N_24281,N_24097);
xor U25950 (N_25950,N_23036,N_21028);
and U25951 (N_25951,N_23204,N_22231);
or U25952 (N_25952,N_23278,N_23889);
xor U25953 (N_25953,N_21150,N_21087);
nor U25954 (N_25954,N_23015,N_24539);
or U25955 (N_25955,N_21827,N_21118);
and U25956 (N_25956,N_20518,N_21971);
or U25957 (N_25957,N_23611,N_20730);
nor U25958 (N_25958,N_23203,N_20399);
nand U25959 (N_25959,N_22619,N_21001);
or U25960 (N_25960,N_20387,N_23755);
nand U25961 (N_25961,N_20924,N_21377);
xnor U25962 (N_25962,N_22694,N_24077);
xnor U25963 (N_25963,N_22736,N_20332);
or U25964 (N_25964,N_23283,N_20998);
or U25965 (N_25965,N_23619,N_22437);
and U25966 (N_25966,N_22646,N_24808);
nor U25967 (N_25967,N_24824,N_23618);
nor U25968 (N_25968,N_21486,N_22129);
or U25969 (N_25969,N_22203,N_22812);
nand U25970 (N_25970,N_22272,N_22380);
and U25971 (N_25971,N_21221,N_23000);
xor U25972 (N_25972,N_20193,N_24430);
or U25973 (N_25973,N_21267,N_21132);
and U25974 (N_25974,N_22909,N_24248);
and U25975 (N_25975,N_21952,N_21363);
nand U25976 (N_25976,N_24270,N_24567);
or U25977 (N_25977,N_22881,N_20991);
xor U25978 (N_25978,N_20950,N_20796);
and U25979 (N_25979,N_22340,N_24827);
nand U25980 (N_25980,N_20446,N_21802);
nand U25981 (N_25981,N_21174,N_21620);
and U25982 (N_25982,N_24573,N_21530);
and U25983 (N_25983,N_22124,N_24611);
and U25984 (N_25984,N_20224,N_24592);
and U25985 (N_25985,N_20267,N_21962);
nor U25986 (N_25986,N_23219,N_22539);
or U25987 (N_25987,N_20682,N_23816);
xnor U25988 (N_25988,N_24042,N_20577);
xor U25989 (N_25989,N_20891,N_24342);
nor U25990 (N_25990,N_23731,N_24786);
or U25991 (N_25991,N_24555,N_24295);
xnor U25992 (N_25992,N_20789,N_22524);
or U25993 (N_25993,N_23069,N_24532);
nand U25994 (N_25994,N_24374,N_22327);
xor U25995 (N_25995,N_21300,N_21454);
nand U25996 (N_25996,N_22257,N_20048);
nor U25997 (N_25997,N_24191,N_22300);
xor U25998 (N_25998,N_24882,N_24618);
xnor U25999 (N_25999,N_22456,N_24978);
xor U26000 (N_26000,N_22065,N_22216);
or U26001 (N_26001,N_21977,N_23807);
or U26002 (N_26002,N_24145,N_20450);
xor U26003 (N_26003,N_20086,N_24775);
and U26004 (N_26004,N_20033,N_23142);
and U26005 (N_26005,N_24879,N_24106);
and U26006 (N_26006,N_21829,N_21517);
xor U26007 (N_26007,N_22891,N_24981);
xor U26008 (N_26008,N_23355,N_24063);
and U26009 (N_26009,N_23102,N_23100);
xor U26010 (N_26010,N_20632,N_24076);
nand U26011 (N_26011,N_24442,N_24715);
or U26012 (N_26012,N_22071,N_22359);
xor U26013 (N_26013,N_21383,N_21480);
or U26014 (N_26014,N_20368,N_23037);
xnor U26015 (N_26015,N_21354,N_22495);
and U26016 (N_26016,N_20439,N_20293);
and U26017 (N_26017,N_23818,N_22292);
nand U26018 (N_26018,N_22482,N_24619);
or U26019 (N_26019,N_24247,N_24856);
or U26020 (N_26020,N_23961,N_22176);
xor U26021 (N_26021,N_21056,N_20763);
and U26022 (N_26022,N_22064,N_20614);
xnor U26023 (N_26023,N_24895,N_21054);
xor U26024 (N_26024,N_23609,N_22894);
nand U26025 (N_26025,N_21253,N_20584);
or U26026 (N_26026,N_20287,N_22528);
nor U26027 (N_26027,N_23664,N_24236);
nand U26028 (N_26028,N_22037,N_20589);
nor U26029 (N_26029,N_23492,N_23587);
and U26030 (N_26030,N_21540,N_20285);
and U26031 (N_26031,N_24092,N_22997);
nor U26032 (N_26032,N_24755,N_23827);
and U26033 (N_26033,N_22969,N_24036);
nor U26034 (N_26034,N_23506,N_22438);
and U26035 (N_26035,N_20513,N_23090);
xor U26036 (N_26036,N_22867,N_22949);
or U26037 (N_26037,N_24826,N_21611);
nor U26038 (N_26038,N_20438,N_21297);
and U26039 (N_26039,N_20305,N_20231);
nor U26040 (N_26040,N_22281,N_22454);
xnor U26041 (N_26041,N_22594,N_24243);
nand U26042 (N_26042,N_21048,N_23328);
or U26043 (N_26043,N_23906,N_23367);
xnor U26044 (N_26044,N_21847,N_22826);
nor U26045 (N_26045,N_21947,N_21694);
nor U26046 (N_26046,N_20675,N_22959);
xor U26047 (N_26047,N_20371,N_21815);
xnor U26048 (N_26048,N_21412,N_20428);
nand U26049 (N_26049,N_23214,N_22289);
nor U26050 (N_26050,N_21737,N_20458);
and U26051 (N_26051,N_21282,N_23402);
or U26052 (N_26052,N_20700,N_22609);
or U26053 (N_26053,N_21638,N_20565);
or U26054 (N_26054,N_22631,N_21126);
nor U26055 (N_26055,N_23858,N_23127);
xnor U26056 (N_26056,N_20729,N_23665);
xor U26057 (N_26057,N_21588,N_24660);
nand U26058 (N_26058,N_22258,N_20186);
or U26059 (N_26059,N_20737,N_22455);
nor U26060 (N_26060,N_21374,N_23088);
and U26061 (N_26061,N_22572,N_24533);
and U26062 (N_26062,N_22178,N_20160);
and U26063 (N_26063,N_23260,N_22485);
and U26064 (N_26064,N_20846,N_23195);
xnor U26065 (N_26065,N_21664,N_21096);
or U26066 (N_26066,N_20775,N_20587);
nor U26067 (N_26067,N_23775,N_22335);
xnor U26068 (N_26068,N_22864,N_20340);
or U26069 (N_26069,N_20099,N_23046);
nand U26070 (N_26070,N_22288,N_23353);
nand U26071 (N_26071,N_22710,N_23051);
nor U26072 (N_26072,N_22743,N_23265);
nor U26073 (N_26073,N_22754,N_24280);
or U26074 (N_26074,N_20469,N_24600);
or U26075 (N_26075,N_21621,N_21817);
nand U26076 (N_26076,N_21940,N_24489);
nand U26077 (N_26077,N_20696,N_21777);
or U26078 (N_26078,N_24828,N_22899);
nor U26079 (N_26079,N_23948,N_21310);
or U26080 (N_26080,N_22908,N_24761);
and U26081 (N_26081,N_20424,N_22752);
or U26082 (N_26082,N_24303,N_21767);
or U26083 (N_26083,N_24719,N_20457);
nand U26084 (N_26084,N_22757,N_21215);
nor U26085 (N_26085,N_23519,N_23106);
xor U26086 (N_26086,N_20523,N_22911);
xnor U26087 (N_26087,N_22251,N_22161);
xnor U26088 (N_26088,N_22010,N_24385);
and U26089 (N_26089,N_22578,N_24005);
xnor U26090 (N_26090,N_22665,N_23445);
or U26091 (N_26091,N_22269,N_23972);
and U26092 (N_26092,N_24992,N_24211);
xnor U26093 (N_26093,N_23885,N_22125);
and U26094 (N_26094,N_24617,N_22920);
nand U26095 (N_26095,N_20858,N_24701);
xnor U26096 (N_26096,N_20753,N_23596);
xnor U26097 (N_26097,N_20095,N_23500);
xor U26098 (N_26098,N_22099,N_21559);
xor U26099 (N_26099,N_20148,N_24649);
xnor U26100 (N_26100,N_21205,N_22556);
xor U26101 (N_26101,N_21000,N_22091);
nor U26102 (N_26102,N_22341,N_23545);
and U26103 (N_26103,N_21645,N_23927);
or U26104 (N_26104,N_24360,N_24825);
nor U26105 (N_26105,N_22526,N_21153);
or U26106 (N_26106,N_23253,N_20906);
and U26107 (N_26107,N_21632,N_20087);
xor U26108 (N_26108,N_20554,N_21434);
xnor U26109 (N_26109,N_22404,N_23657);
nor U26110 (N_26110,N_21972,N_22344);
and U26111 (N_26111,N_20778,N_21081);
xor U26112 (N_26112,N_22671,N_22771);
nand U26113 (N_26113,N_24061,N_20204);
and U26114 (N_26114,N_24637,N_22403);
and U26115 (N_26115,N_23484,N_22676);
nor U26116 (N_26116,N_24764,N_21294);
xor U26117 (N_26117,N_23249,N_24315);
and U26118 (N_26118,N_22822,N_23498);
and U26119 (N_26119,N_20333,N_21314);
nand U26120 (N_26120,N_23360,N_24122);
and U26121 (N_26121,N_20360,N_23369);
or U26122 (N_26122,N_24926,N_23358);
nor U26123 (N_26123,N_21850,N_21707);
nor U26124 (N_26124,N_20922,N_22012);
nor U26125 (N_26125,N_22808,N_21810);
nand U26126 (N_26126,N_20362,N_23981);
and U26127 (N_26127,N_20028,N_23793);
or U26128 (N_26128,N_21796,N_23019);
nor U26129 (N_26129,N_21855,N_20329);
nand U26130 (N_26130,N_21526,N_23789);
nor U26131 (N_26131,N_20179,N_22381);
nor U26132 (N_26132,N_24114,N_23434);
nor U26133 (N_26133,N_24400,N_22321);
nand U26134 (N_26134,N_21786,N_20721);
xor U26135 (N_26135,N_24517,N_23850);
and U26136 (N_26136,N_24111,N_20583);
nand U26137 (N_26137,N_22581,N_22074);
and U26138 (N_26138,N_22739,N_22725);
nor U26139 (N_26139,N_22592,N_20413);
or U26140 (N_26140,N_23516,N_20322);
nor U26141 (N_26141,N_21504,N_21679);
nand U26142 (N_26142,N_23237,N_22035);
xnor U26143 (N_26143,N_24549,N_24027);
and U26144 (N_26144,N_23590,N_23828);
xor U26145 (N_26145,N_23648,N_23104);
nor U26146 (N_26146,N_21231,N_22900);
and U26147 (N_26147,N_24832,N_21095);
and U26148 (N_26148,N_22209,N_23056);
xnor U26149 (N_26149,N_20920,N_23639);
and U26150 (N_26150,N_21370,N_23470);
or U26151 (N_26151,N_24706,N_24878);
xnor U26152 (N_26152,N_20657,N_21859);
xnor U26153 (N_26153,N_24647,N_20175);
xnor U26154 (N_26154,N_22083,N_23875);
and U26155 (N_26155,N_22848,N_20418);
or U26156 (N_26156,N_23089,N_21958);
nor U26157 (N_26157,N_20635,N_21671);
nand U26158 (N_26158,N_22543,N_22790);
and U26159 (N_26159,N_21714,N_20710);
nand U26160 (N_26160,N_24259,N_22244);
or U26161 (N_26161,N_20460,N_23094);
nor U26162 (N_26162,N_23248,N_21914);
and U26163 (N_26163,N_20433,N_20230);
and U26164 (N_26164,N_22863,N_23952);
or U26165 (N_26165,N_23190,N_22889);
or U26166 (N_26166,N_23754,N_22077);
xnor U26167 (N_26167,N_20237,N_23696);
nand U26168 (N_26168,N_23798,N_23315);
and U26169 (N_26169,N_24182,N_24214);
and U26170 (N_26170,N_23528,N_21740);
xnor U26171 (N_26171,N_24142,N_24050);
xnor U26172 (N_26172,N_21327,N_21182);
nor U26173 (N_26173,N_20636,N_21073);
xnor U26174 (N_26174,N_21098,N_22931);
nand U26175 (N_26175,N_20957,N_23955);
nand U26176 (N_26176,N_23735,N_23806);
or U26177 (N_26177,N_23811,N_24515);
and U26178 (N_26178,N_21922,N_23616);
nand U26179 (N_26179,N_23984,N_20930);
nor U26180 (N_26180,N_21782,N_20954);
nand U26181 (N_26181,N_21865,N_21149);
and U26182 (N_26182,N_20304,N_20323);
nor U26183 (N_26183,N_24457,N_23632);
or U26184 (N_26184,N_23456,N_20833);
xor U26185 (N_26185,N_23866,N_21807);
nand U26186 (N_26186,N_20863,N_24670);
nand U26187 (N_26187,N_20842,N_22869);
or U26188 (N_26188,N_20639,N_22797);
and U26189 (N_26189,N_21832,N_20941);
or U26190 (N_26190,N_24576,N_21270);
and U26191 (N_26191,N_23119,N_24031);
nor U26192 (N_26192,N_20065,N_24616);
xnor U26193 (N_26193,N_20059,N_21908);
nand U26194 (N_26194,N_20791,N_21756);
nand U26195 (N_26195,N_22365,N_22086);
and U26196 (N_26196,N_23567,N_20077);
nand U26197 (N_26197,N_24941,N_21735);
nor U26198 (N_26198,N_21706,N_24540);
and U26199 (N_26199,N_21379,N_20075);
or U26200 (N_26200,N_21401,N_22976);
xnor U26201 (N_26201,N_24774,N_23418);
or U26202 (N_26202,N_22861,N_22724);
and U26203 (N_26203,N_24219,N_23159);
or U26204 (N_26204,N_20548,N_22374);
or U26205 (N_26205,N_23029,N_22046);
or U26206 (N_26206,N_24187,N_24612);
nor U26207 (N_26207,N_24570,N_21406);
nand U26208 (N_26208,N_20573,N_21407);
nand U26209 (N_26209,N_23338,N_24680);
and U26210 (N_26210,N_20133,N_20119);
or U26211 (N_26211,N_20545,N_20714);
nor U26212 (N_26212,N_21304,N_24437);
and U26213 (N_26213,N_24004,N_21380);
xor U26214 (N_26214,N_24302,N_22295);
nor U26215 (N_26215,N_20990,N_21162);
or U26216 (N_26216,N_24874,N_22590);
nor U26217 (N_26217,N_21024,N_20572);
nor U26218 (N_26218,N_21266,N_20726);
xor U26219 (N_26219,N_23672,N_21915);
nor U26220 (N_26220,N_22759,N_20394);
or U26221 (N_26221,N_22636,N_23782);
and U26222 (N_26222,N_24923,N_21921);
or U26223 (N_26223,N_22347,N_22014);
and U26224 (N_26224,N_24420,N_21369);
xor U26225 (N_26225,N_24634,N_22516);
xor U26226 (N_26226,N_24418,N_22682);
nand U26227 (N_26227,N_24354,N_20948);
nor U26228 (N_26228,N_21104,N_23876);
xnor U26229 (N_26229,N_22031,N_21841);
xnor U26230 (N_26230,N_21842,N_23150);
or U26231 (N_26231,N_20344,N_21561);
xor U26232 (N_26232,N_21964,N_21008);
or U26233 (N_26233,N_20009,N_22948);
and U26234 (N_26234,N_23956,N_21764);
xnor U26235 (N_26235,N_24389,N_20909);
xnor U26236 (N_26236,N_20377,N_20508);
nand U26237 (N_26237,N_24238,N_23630);
nand U26238 (N_26238,N_21800,N_23247);
nand U26239 (N_26239,N_23561,N_21988);
nor U26240 (N_26240,N_21860,N_21107);
xnor U26241 (N_26241,N_23161,N_21692);
nand U26242 (N_26242,N_20184,N_22862);
and U26243 (N_26243,N_24294,N_21531);
or U26244 (N_26244,N_20856,N_21499);
nor U26245 (N_26245,N_21459,N_21885);
xnor U26246 (N_26246,N_22005,N_22200);
and U26247 (N_26247,N_23819,N_24762);
or U26248 (N_26248,N_20544,N_23194);
xnor U26249 (N_26249,N_21009,N_20135);
xnor U26250 (N_26250,N_20389,N_23264);
and U26251 (N_26251,N_21974,N_23583);
nand U26252 (N_26252,N_21813,N_20361);
xor U26253 (N_26253,N_24930,N_23884);
and U26254 (N_26254,N_24444,N_21739);
nor U26255 (N_26255,N_22821,N_20295);
nand U26256 (N_26256,N_20228,N_20969);
or U26257 (N_26257,N_24700,N_24819);
xnor U26258 (N_26258,N_20562,N_24277);
xnor U26259 (N_26259,N_24534,N_23628);
or U26260 (N_26260,N_23279,N_21446);
or U26261 (N_26261,N_21957,N_23550);
and U26262 (N_26262,N_23592,N_21341);
nor U26263 (N_26263,N_24754,N_23221);
or U26264 (N_26264,N_22254,N_20079);
xor U26265 (N_26265,N_21193,N_21618);
or U26266 (N_26266,N_20944,N_21170);
or U26267 (N_26267,N_22402,N_22184);
nand U26268 (N_26268,N_24321,N_20982);
or U26269 (N_26269,N_20692,N_23224);
and U26270 (N_26270,N_24377,N_21592);
or U26271 (N_26271,N_23641,N_22278);
and U26272 (N_26272,N_22738,N_22935);
and U26273 (N_26273,N_23778,N_21795);
xnor U26274 (N_26274,N_23841,N_20098);
nand U26275 (N_26275,N_20561,N_22522);
nand U26276 (N_26276,N_20057,N_22003);
nand U26277 (N_26277,N_24656,N_23714);
nor U26278 (N_26278,N_22852,N_20308);
xor U26279 (N_26279,N_21529,N_22601);
xor U26280 (N_26280,N_22961,N_23997);
nand U26281 (N_26281,N_22043,N_24176);
xor U26282 (N_26282,N_22506,N_21805);
xor U26283 (N_26283,N_24125,N_22720);
xor U26284 (N_26284,N_23674,N_21793);
and U26285 (N_26285,N_24685,N_22073);
xnor U26286 (N_26286,N_24440,N_20738);
or U26287 (N_26287,N_24309,N_20493);
nor U26288 (N_26288,N_20120,N_20898);
xnor U26289 (N_26289,N_21269,N_23693);
nand U26290 (N_26290,N_20235,N_21556);
nor U26291 (N_26291,N_24591,N_22484);
xor U26292 (N_26292,N_20673,N_22626);
and U26293 (N_26293,N_22963,N_21206);
nor U26294 (N_26294,N_21933,N_24818);
nor U26295 (N_26295,N_24058,N_23295);
xnor U26296 (N_26296,N_24319,N_24478);
nand U26297 (N_26297,N_20391,N_21720);
nor U26298 (N_26298,N_22322,N_20162);
xor U26299 (N_26299,N_22792,N_24388);
nand U26300 (N_26300,N_20153,N_24109);
xnor U26301 (N_26301,N_23916,N_22056);
nand U26302 (N_26302,N_21869,N_21894);
and U26303 (N_26303,N_22391,N_22154);
nor U26304 (N_26304,N_23783,N_24468);
nor U26305 (N_26305,N_23769,N_22625);
nor U26306 (N_26306,N_22879,N_23836);
xnor U26307 (N_26307,N_20155,N_23517);
nor U26308 (N_26308,N_23341,N_22990);
nand U26309 (N_26309,N_20780,N_20043);
nor U26310 (N_26310,N_23113,N_22237);
xor U26311 (N_26311,N_20383,N_20403);
xor U26312 (N_26312,N_21328,N_22666);
or U26313 (N_26313,N_20459,N_22858);
xor U26314 (N_26314,N_20642,N_21936);
nor U26315 (N_26315,N_24119,N_22144);
nand U26316 (N_26316,N_22943,N_23605);
or U26317 (N_26317,N_22501,N_24024);
nor U26318 (N_26318,N_22133,N_22847);
nor U26319 (N_26319,N_20112,N_24969);
nand U26320 (N_26320,N_24098,N_20115);
nand U26321 (N_26321,N_20223,N_24538);
nor U26322 (N_26322,N_23553,N_20407);
xor U26323 (N_26323,N_24118,N_21418);
and U26324 (N_26324,N_20183,N_24387);
or U26325 (N_26325,N_21878,N_21139);
and U26326 (N_26326,N_21808,N_20000);
xor U26327 (N_26327,N_23303,N_21973);
nor U26328 (N_26328,N_22307,N_20965);
xor U26329 (N_26329,N_21133,N_21386);
or U26330 (N_26330,N_20798,N_20907);
or U26331 (N_26331,N_20486,N_23534);
and U26332 (N_26332,N_20369,N_24291);
and U26333 (N_26333,N_24562,N_20447);
nor U26334 (N_26334,N_23537,N_23202);
nand U26335 (N_26335,N_22512,N_22217);
or U26336 (N_26336,N_21743,N_22027);
nor U26337 (N_26337,N_20553,N_20688);
nand U26338 (N_26338,N_23723,N_24049);
and U26339 (N_26339,N_21247,N_22954);
nand U26340 (N_26340,N_20249,N_24085);
nor U26341 (N_26341,N_22323,N_22560);
or U26342 (N_26342,N_24047,N_23586);
xnor U26343 (N_26343,N_23580,N_20178);
and U26344 (N_26344,N_24703,N_23438);
or U26345 (N_26345,N_20880,N_20316);
or U26346 (N_26346,N_23496,N_23924);
nand U26347 (N_26347,N_23263,N_22895);
nor U26348 (N_26348,N_22772,N_20834);
nand U26349 (N_26349,N_24120,N_24268);
xor U26350 (N_26350,N_22541,N_21712);
xnor U26351 (N_26351,N_21212,N_24914);
and U26352 (N_26352,N_23676,N_23276);
nor U26353 (N_26353,N_21021,N_20378);
nor U26354 (N_26354,N_24015,N_21898);
or U26355 (N_26355,N_21198,N_23472);
or U26356 (N_26356,N_24791,N_23654);
xor U26357 (N_26357,N_22390,N_20104);
xnor U26358 (N_26358,N_22026,N_24023);
and U26359 (N_26359,N_22271,N_23581);
and U26360 (N_26360,N_20547,N_21984);
nor U26361 (N_26361,N_20622,N_21050);
xor U26362 (N_26362,N_21173,N_21144);
and U26363 (N_26363,N_21753,N_20521);
nand U26364 (N_26364,N_21090,N_23757);
xor U26365 (N_26365,N_21923,N_22653);
nor U26366 (N_26366,N_22204,N_20618);
or U26367 (N_26367,N_23170,N_21660);
nand U26368 (N_26368,N_20708,N_24000);
xnor U26369 (N_26369,N_24467,N_20973);
nand U26370 (N_26370,N_20670,N_22304);
xnor U26371 (N_26371,N_21887,N_24944);
nor U26372 (N_26372,N_24451,N_21091);
xor U26373 (N_26373,N_24985,N_20935);
or U26374 (N_26374,N_22114,N_23242);
or U26375 (N_26375,N_20300,N_24860);
and U26376 (N_26376,N_20016,N_20445);
nor U26377 (N_26377,N_21183,N_24594);
or U26378 (N_26378,N_21477,N_24100);
and U26379 (N_26379,N_20805,N_22635);
xor U26380 (N_26380,N_23702,N_20163);
xnor U26381 (N_26381,N_23680,N_22249);
nand U26382 (N_26382,N_22552,N_22763);
nor U26383 (N_26383,N_20999,N_24750);
nor U26384 (N_26384,N_21580,N_22349);
nor U26385 (N_26385,N_21396,N_23865);
xnor U26386 (N_26386,N_24221,N_20341);
nand U26387 (N_26387,N_23745,N_24509);
and U26388 (N_26388,N_20955,N_22284);
xnor U26389 (N_26389,N_20082,N_23547);
and U26390 (N_26390,N_24531,N_22312);
and U26391 (N_26391,N_22095,N_22422);
nand U26392 (N_26392,N_23324,N_23196);
or U26393 (N_26393,N_22186,N_22987);
nor U26394 (N_26394,N_24028,N_21652);
nand U26395 (N_26395,N_20637,N_20474);
or U26396 (N_26396,N_22499,N_24783);
nor U26397 (N_26397,N_24547,N_23892);
nor U26398 (N_26398,N_22436,N_23186);
nor U26399 (N_26399,N_22825,N_22767);
xnor U26400 (N_26400,N_20410,N_21228);
and U26401 (N_26401,N_20769,N_24924);
or U26402 (N_26402,N_23709,N_22158);
and U26403 (N_26403,N_21801,N_22748);
nor U26404 (N_26404,N_24336,N_20755);
nor U26405 (N_26405,N_20507,N_22053);
and U26406 (N_26406,N_22098,N_24333);
or U26407 (N_26407,N_21362,N_21612);
or U26408 (N_26408,N_23542,N_21368);
nor U26409 (N_26409,N_22708,N_23301);
and U26410 (N_26410,N_20641,N_22873);
nor U26411 (N_26411,N_23712,N_23670);
or U26412 (N_26412,N_24449,N_24307);
or U26413 (N_26413,N_20258,N_23946);
or U26414 (N_26414,N_20538,N_21680);
nor U26415 (N_26415,N_22206,N_22917);
and U26416 (N_26416,N_20707,N_20484);
and U26417 (N_26417,N_24423,N_23482);
xnor U26418 (N_26418,N_22637,N_24162);
nor U26419 (N_26419,N_20356,N_21892);
or U26420 (N_26420,N_20123,N_23381);
and U26421 (N_26421,N_24933,N_22070);
xnor U26422 (N_26422,N_23348,N_24284);
or U26423 (N_26423,N_21819,N_23097);
nand U26424 (N_26424,N_24308,N_23180);
and U26425 (N_26425,N_24127,N_22109);
nand U26426 (N_26426,N_21844,N_24862);
or U26427 (N_26427,N_21565,N_23435);
nor U26428 (N_26428,N_23079,N_22468);
xnor U26429 (N_26429,N_22647,N_22401);
xor U26430 (N_26430,N_20260,N_23501);
nand U26431 (N_26431,N_24494,N_21953);
nand U26432 (N_26432,N_21340,N_20317);
and U26433 (N_26433,N_24154,N_24530);
xnor U26434 (N_26434,N_21934,N_21570);
and U26435 (N_26435,N_22562,N_22958);
nor U26436 (N_26436,N_21356,N_24525);
nor U26437 (N_26437,N_23475,N_20246);
nor U26438 (N_26438,N_21868,N_23448);
or U26439 (N_26439,N_24224,N_23637);
or U26440 (N_26440,N_24713,N_23235);
nor U26441 (N_26441,N_23808,N_23908);
or U26442 (N_26442,N_22011,N_24405);
nor U26443 (N_26443,N_21838,N_23730);
nand U26444 (N_26444,N_20145,N_24296);
xor U26445 (N_26445,N_20444,N_22419);
and U26446 (N_26446,N_24431,N_21138);
and U26447 (N_26447,N_22152,N_20947);
xnor U26448 (N_26448,N_20201,N_24195);
and U26449 (N_26449,N_20068,N_21143);
xor U26450 (N_26450,N_21571,N_24227);
xnor U26451 (N_26451,N_24524,N_23555);
and U26452 (N_26452,N_21520,N_23129);
nor U26453 (N_26453,N_22884,N_24306);
nand U26454 (N_26454,N_21555,N_23365);
and U26455 (N_26455,N_21667,N_24842);
xor U26456 (N_26456,N_24366,N_21302);
nor U26457 (N_26457,N_22072,N_20266);
xor U26458 (N_26458,N_20517,N_24798);
xor U26459 (N_26459,N_24057,N_23652);
and U26460 (N_26460,N_22824,N_24560);
xnor U26461 (N_26461,N_22140,N_21784);
xnor U26462 (N_26462,N_23867,N_23175);
and U26463 (N_26463,N_24368,N_24608);
nand U26464 (N_26464,N_23409,N_23450);
nor U26465 (N_26465,N_24505,N_22146);
nor U26466 (N_26466,N_22727,N_24938);
and U26467 (N_26467,N_23595,N_20240);
and U26468 (N_26468,N_23382,N_20631);
or U26469 (N_26469,N_20967,N_22563);
and U26470 (N_26470,N_20181,N_22796);
xnor U26471 (N_26471,N_23111,N_20977);
and U26472 (N_26472,N_24364,N_23135);
or U26473 (N_26473,N_22262,N_24131);
xor U26474 (N_26474,N_20665,N_20715);
xnor U26475 (N_26475,N_24716,N_22722);
nand U26476 (N_26476,N_22417,N_20663);
and U26477 (N_26477,N_22854,N_22978);
xnor U26478 (N_26478,N_20586,N_23408);
or U26479 (N_26479,N_21291,N_21820);
nand U26480 (N_26480,N_24650,N_24056);
nor U26481 (N_26481,N_20467,N_22548);
nor U26482 (N_26482,N_23240,N_23844);
xor U26483 (N_26483,N_23207,N_21703);
and U26484 (N_26484,N_21234,N_20968);
and U26485 (N_26485,N_24199,N_23949);
or U26486 (N_26486,N_22882,N_21359);
nor U26487 (N_26487,N_22574,N_22314);
nor U26488 (N_26488,N_23829,N_21102);
nand U26489 (N_26489,N_23226,N_23183);
and U26490 (N_26490,N_23990,N_20374);
nor U26491 (N_26491,N_20541,N_24889);
xor U26492 (N_26492,N_23066,N_20885);
and U26493 (N_26493,N_22612,N_24285);
nand U26494 (N_26494,N_23803,N_22233);
and U26495 (N_26495,N_22252,N_21172);
xnor U26496 (N_26496,N_24479,N_21308);
xnor U26497 (N_26497,N_20094,N_23255);
xor U26498 (N_26498,N_24412,N_22283);
and U26499 (N_26499,N_20650,N_23123);
xor U26500 (N_26500,N_22377,N_22697);
and U26501 (N_26501,N_22242,N_22532);
or U26502 (N_26502,N_20199,N_21331);
and U26503 (N_26503,N_23826,N_23292);
nor U26504 (N_26504,N_22871,N_23130);
xnor U26505 (N_26505,N_20976,N_22525);
xor U26506 (N_26506,N_23764,N_20685);
nor U26507 (N_26507,N_24932,N_24196);
nand U26508 (N_26508,N_20110,N_22116);
and U26509 (N_26509,N_24722,N_21990);
and U26510 (N_26510,N_23951,N_23513);
xor U26511 (N_26511,N_23505,N_20297);
xnor U26512 (N_26512,N_22678,N_21031);
nor U26513 (N_26513,N_22535,N_24160);
xnor U26514 (N_26514,N_22128,N_21856);
or U26515 (N_26515,N_20054,N_20840);
or U26516 (N_26516,N_21397,N_21108);
or U26517 (N_26517,N_23584,N_20192);
xor U26518 (N_26518,N_21560,N_22045);
and U26519 (N_26519,N_24311,N_21431);
xnor U26520 (N_26520,N_20609,N_23458);
and U26521 (N_26521,N_23493,N_21353);
nor U26522 (N_26522,N_20974,N_20105);
or U26523 (N_26523,N_21444,N_22142);
nor U26524 (N_26524,N_24244,N_23300);
or U26525 (N_26525,N_21770,N_23209);
nand U26526 (N_26526,N_24054,N_22079);
nor U26527 (N_26527,N_21323,N_24139);
nor U26528 (N_26528,N_23442,N_21932);
nand U26529 (N_26529,N_24137,N_24424);
or U26530 (N_26530,N_22996,N_20878);
nor U26531 (N_26531,N_20925,N_21226);
and U26532 (N_26532,N_22874,N_21213);
or U26533 (N_26533,N_22583,N_21938);
nor U26534 (N_26534,N_23267,N_23497);
and U26535 (N_26535,N_24971,N_23543);
nand U26536 (N_26536,N_22839,N_23638);
or U26537 (N_26537,N_20017,N_23487);
or U26538 (N_26538,N_22674,N_21919);
xnor U26539 (N_26539,N_22566,N_23999);
nor U26540 (N_26540,N_20800,N_24714);
xnor U26541 (N_26541,N_22273,N_23507);
and U26542 (N_26542,N_21905,N_22616);
or U26543 (N_26543,N_21641,N_20130);
and U26544 (N_26544,N_22421,N_21200);
or U26545 (N_26545,N_20902,N_24128);
and U26546 (N_26546,N_24682,N_21283);
and U26547 (N_26547,N_20985,N_24212);
xnor U26548 (N_26548,N_21116,N_21447);
or U26549 (N_26549,N_22705,N_20718);
nor U26550 (N_26550,N_21468,N_20355);
and U26551 (N_26551,N_20001,N_22904);
and U26552 (N_26552,N_24030,N_23614);
or U26553 (N_26553,N_20182,N_20525);
xnor U26554 (N_26554,N_24034,N_22334);
or U26555 (N_26555,N_22956,N_20772);
and U26556 (N_26556,N_20161,N_24696);
and U26557 (N_26557,N_22165,N_23356);
or U26558 (N_26558,N_21003,N_22970);
or U26559 (N_26559,N_23032,N_20736);
xor U26560 (N_26560,N_20343,N_20643);
or U26561 (N_26561,N_23541,N_20024);
nand U26562 (N_26562,N_22303,N_21110);
or U26563 (N_26563,N_23259,N_21760);
or U26564 (N_26564,N_23038,N_21883);
and U26565 (N_26565,N_21946,N_24858);
or U26566 (N_26566,N_23533,N_23462);
nor U26567 (N_26567,N_23001,N_22642);
nand U26568 (N_26568,N_22775,N_21773);
or U26569 (N_26569,N_22148,N_21263);
xor U26570 (N_26570,N_21125,N_22993);
or U26571 (N_26571,N_20217,N_23973);
and U26572 (N_26572,N_21700,N_22549);
nor U26573 (N_26573,N_22989,N_21242);
nor U26574 (N_26574,N_20879,N_22016);
xor U26575 (N_26575,N_21033,N_22363);
nor U26576 (N_26576,N_23539,N_22865);
nand U26577 (N_26577,N_23651,N_24083);
or U26578 (N_26578,N_21950,N_23840);
or U26579 (N_26579,N_20402,N_21067);
xnor U26580 (N_26580,N_23627,N_21053);
nand U26581 (N_26581,N_23131,N_24501);
xnor U26582 (N_26582,N_22282,N_22962);
nand U26583 (N_26583,N_22338,N_23589);
and U26584 (N_26584,N_22721,N_23873);
or U26585 (N_26585,N_24604,N_22378);
and U26586 (N_26586,N_22104,N_24795);
and U26587 (N_26587,N_20200,N_20263);
nor U26588 (N_26588,N_23061,N_21598);
and U26589 (N_26589,N_22860,N_22941);
nor U26590 (N_26590,N_20081,N_20202);
nand U26591 (N_26591,N_22090,N_21196);
or U26592 (N_26592,N_21702,N_20034);
or U26593 (N_26593,N_23227,N_21012);
nand U26594 (N_26594,N_24463,N_22567);
xor U26595 (N_26595,N_20929,N_23184);
nand U26596 (N_26596,N_24369,N_21900);
or U26597 (N_26597,N_22500,N_21854);
nor U26598 (N_26598,N_24185,N_21672);
or U26599 (N_26599,N_23943,N_21404);
xnor U26600 (N_26600,N_20895,N_21781);
or U26601 (N_26601,N_24789,N_24586);
nand U26602 (N_26602,N_23706,N_21730);
nor U26603 (N_26603,N_22937,N_23560);
nor U26604 (N_26604,N_23393,N_24507);
nand U26605 (N_26605,N_23602,N_23229);
or U26606 (N_26606,N_22198,N_22058);
or U26607 (N_26607,N_24859,N_20076);
nor U26608 (N_26608,N_20601,N_20767);
xor U26609 (N_26609,N_22008,N_22800);
and U26610 (N_26610,N_24230,N_23368);
or U26611 (N_26611,N_22245,N_20575);
nand U26612 (N_26612,N_20151,N_22385);
nand U26613 (N_26613,N_21728,N_20740);
xnor U26614 (N_26614,N_21725,N_24258);
nand U26615 (N_26615,N_24815,N_23258);
xnor U26616 (N_26616,N_21100,N_22975);
and U26617 (N_26617,N_20794,N_20529);
and U26618 (N_26618,N_24972,N_23643);
nor U26619 (N_26619,N_20823,N_23613);
or U26620 (N_26620,N_21271,N_21190);
nor U26621 (N_26621,N_22984,N_23965);
or U26622 (N_26622,N_21881,N_21715);
nand U26623 (N_26623,N_24817,N_23814);
xor U26624 (N_26624,N_24252,N_22051);
nor U26625 (N_26625,N_24792,N_24473);
and U26626 (N_26626,N_24223,N_24476);
or U26627 (N_26627,N_24316,N_23335);
nand U26628 (N_26628,N_20386,N_20370);
xor U26629 (N_26629,N_21567,N_22364);
xor U26630 (N_26630,N_20758,N_23208);
xor U26631 (N_26631,N_24272,N_22718);
nor U26632 (N_26632,N_21276,N_24952);
nor U26633 (N_26633,N_24864,N_20567);
xor U26634 (N_26634,N_21422,N_22375);
nand U26635 (N_26635,N_22100,N_22306);
and U26636 (N_26636,N_24693,N_21023);
or U26637 (N_26637,N_21235,N_23766);
and U26638 (N_26638,N_24709,N_24345);
and U26639 (N_26639,N_22770,N_21945);
xor U26640 (N_26640,N_21787,N_20503);
xor U26641 (N_26641,N_21949,N_23152);
nand U26642 (N_26642,N_24752,N_24955);
xor U26643 (N_26643,N_22432,N_21927);
nand U26644 (N_26644,N_20488,N_22787);
nor U26645 (N_26645,N_24678,N_21035);
nand U26646 (N_26646,N_20093,N_22358);
or U26647 (N_26647,N_20499,N_21603);
xnor U26648 (N_26648,N_22746,N_21094);
xor U26649 (N_26649,N_24906,N_24869);
nor U26650 (N_26650,N_21366,N_20662);
nor U26651 (N_26651,N_23166,N_23546);
nor U26652 (N_26652,N_21544,N_21161);
or U26653 (N_26653,N_21956,N_20210);
or U26654 (N_26654,N_21902,N_21489);
nor U26655 (N_26655,N_20036,N_20070);
xor U26656 (N_26656,N_22112,N_24167);
nand U26657 (N_26657,N_20157,N_20349);
xnor U26658 (N_26658,N_20694,N_24736);
nor U26659 (N_26659,N_20971,N_21831);
xor U26660 (N_26660,N_23666,N_24446);
xor U26661 (N_26661,N_23197,N_23640);
or U26662 (N_26662,N_24838,N_23009);
xor U26663 (N_26663,N_20126,N_21872);
or U26664 (N_26664,N_21996,N_24850);
or U26665 (N_26665,N_23096,N_23030);
or U26666 (N_26666,N_20116,N_24708);
xnor U26667 (N_26667,N_21487,N_23261);
and U26668 (N_26668,N_21891,N_21045);
and U26669 (N_26669,N_20041,N_23658);
nor U26670 (N_26670,N_24946,N_24893);
xor U26671 (N_26671,N_22449,N_21441);
xor U26672 (N_26672,N_21248,N_21343);
xor U26673 (N_26673,N_24967,N_21890);
or U26674 (N_26674,N_21078,N_20229);
and U26675 (N_26675,N_22330,N_23375);
and U26676 (N_26676,N_22681,N_23732);
nor U26677 (N_26677,N_20325,N_24222);
nor U26678 (N_26678,N_24581,N_21194);
xor U26679 (N_26679,N_23147,N_20603);
or U26680 (N_26680,N_23075,N_23845);
or U26681 (N_26681,N_24527,N_22731);
nand U26682 (N_26682,N_21337,N_20540);
xor U26683 (N_26683,N_20379,N_22513);
and U26684 (N_26684,N_23852,N_21983);
or U26685 (N_26685,N_20585,N_24068);
nand U26686 (N_26686,N_23673,N_21257);
and U26687 (N_26687,N_24452,N_20766);
nor U26688 (N_26688,N_24603,N_22055);
xnor U26689 (N_26689,N_22756,N_21741);
or U26690 (N_26690,N_21937,N_20411);
or U26691 (N_26691,N_23340,N_21313);
and U26692 (N_26692,N_21229,N_24202);
nand U26693 (N_26693,N_24867,N_21264);
nor U26694 (N_26694,N_24563,N_21619);
or U26695 (N_26695,N_21062,N_21142);
xnor U26696 (N_26696,N_23556,N_22130);
or U26697 (N_26697,N_22264,N_20724);
or U26698 (N_26698,N_21399,N_20421);
and U26699 (N_26699,N_20422,N_24779);
nand U26700 (N_26700,N_20468,N_22435);
xor U26701 (N_26701,N_21083,N_21649);
xnor U26702 (N_26702,N_20857,N_24062);
nand U26703 (N_26703,N_22850,N_21089);
xor U26704 (N_26704,N_22383,N_22145);
and U26705 (N_26705,N_20903,N_22465);
nor U26706 (N_26706,N_22373,N_24421);
nor U26707 (N_26707,N_21686,N_23317);
nor U26708 (N_26708,N_24396,N_20698);
or U26709 (N_26709,N_20978,N_24067);
or U26710 (N_26710,N_21040,N_20560);
nor U26711 (N_26711,N_20473,N_20995);
nand U26712 (N_26712,N_24891,N_22270);
nand U26713 (N_26713,N_22337,N_21607);
nand U26714 (N_26714,N_23086,N_22062);
and U26715 (N_26715,N_24313,N_22015);
xor U26716 (N_26716,N_23465,N_21986);
or U26717 (N_26717,N_23594,N_22733);
xnor U26718 (N_26718,N_23729,N_23453);
and U26719 (N_26719,N_24046,N_20384);
or U26720 (N_26720,N_24695,N_24689);
nand U26721 (N_26721,N_22683,N_21074);
or U26722 (N_26722,N_22169,N_20367);
xnor U26723 (N_26723,N_22247,N_22191);
xor U26724 (N_26724,N_24275,N_20911);
xnor U26725 (N_26725,N_22794,N_23174);
nand U26726 (N_26726,N_23945,N_22602);
and U26727 (N_26727,N_20822,N_21325);
xor U26728 (N_26728,N_23370,N_20174);
xnor U26729 (N_26729,N_23794,N_24645);
nor U26730 (N_26730,N_23074,N_21665);
nand U26731 (N_26731,N_20398,N_24434);
xor U26732 (N_26732,N_20816,N_23531);
or U26733 (N_26733,N_20928,N_24189);
nor U26734 (N_26734,N_22213,N_23274);
nor U26735 (N_26735,N_22488,N_20993);
and U26736 (N_26736,N_24397,N_21493);
or U26737 (N_26737,N_24293,N_24624);
and U26738 (N_26738,N_20313,N_20579);
and U26739 (N_26739,N_21790,N_24765);
and U26740 (N_26740,N_20103,N_23243);
or U26741 (N_26741,N_20291,N_21004);
nor U26742 (N_26742,N_24654,N_21852);
nor U26743 (N_26743,N_23878,N_21350);
and U26744 (N_26744,N_22250,N_21929);
and U26745 (N_26745,N_24545,N_21440);
nor U26746 (N_26746,N_21214,N_21075);
xnor U26747 (N_26747,N_20852,N_22868);
nor U26748 (N_26748,N_21355,N_23392);
nor U26749 (N_26749,N_23710,N_21290);
and U26750 (N_26750,N_22357,N_21763);
and U26751 (N_26751,N_21682,N_21515);
or U26752 (N_26752,N_23760,N_23756);
or U26753 (N_26753,N_21344,N_23902);
xor U26754 (N_26754,N_23330,N_22924);
or U26755 (N_26755,N_23776,N_20933);
or U26756 (N_26756,N_21508,N_20380);
nor U26757 (N_26757,N_21134,N_23691);
nor U26758 (N_26758,N_23872,N_20619);
xnor U26759 (N_26759,N_21195,N_20008);
xnor U26760 (N_26760,N_23603,N_24753);
nor U26761 (N_26761,N_21509,N_24770);
xnor U26762 (N_26762,N_20628,N_20546);
nand U26763 (N_26763,N_22195,N_21851);
or U26764 (N_26764,N_22021,N_23615);
nand U26765 (N_26765,N_22487,N_22662);
xnor U26766 (N_26766,N_20047,N_20061);
xor U26767 (N_26767,N_23210,N_20594);
nand U26768 (N_26768,N_24683,N_22639);
or U26769 (N_26769,N_24759,N_24037);
and U26770 (N_26770,N_21999,N_23621);
nand U26771 (N_26771,N_23239,N_24051);
nor U26772 (N_26772,N_21419,N_23758);
nor U26773 (N_26773,N_24814,N_21581);
xnor U26774 (N_26774,N_21595,N_23815);
nand U26775 (N_26775,N_22545,N_20420);
nor U26776 (N_26776,N_23121,N_22774);
or U26777 (N_26777,N_21307,N_24497);
nand U26778 (N_26778,N_21136,N_22180);
xnor U26779 (N_26779,N_21262,N_22123);
xnor U26780 (N_26780,N_20330,N_23914);
nor U26781 (N_26781,N_24846,N_24554);
and U26782 (N_26782,N_24958,N_22703);
or U26783 (N_26783,N_22188,N_24419);
nor U26784 (N_26784,N_22020,N_20838);
nand U26785 (N_26785,N_24482,N_24599);
nand U26786 (N_26786,N_22998,N_20440);
nor U26787 (N_26787,N_24568,N_21586);
xor U26788 (N_26788,N_22042,N_22324);
or U26789 (N_26789,N_23257,N_23931);
xnor U26790 (N_26790,N_23763,N_22087);
and U26791 (N_26791,N_24632,N_20321);
and U26792 (N_26792,N_20027,N_22768);
nand U26793 (N_26793,N_22918,N_22559);
nor U26794 (N_26794,N_21127,N_20254);
and U26795 (N_26795,N_23419,N_22579);
or U26796 (N_26796,N_24636,N_20855);
xnor U26797 (N_26797,N_24143,N_21453);
and U26798 (N_26798,N_24404,N_22689);
nand U26799 (N_26799,N_20946,N_24059);
nor U26800 (N_26800,N_24469,N_22370);
nand U26801 (N_26801,N_22331,N_23059);
nor U26802 (N_26802,N_22034,N_22571);
nor U26803 (N_26803,N_24011,N_23077);
and U26804 (N_26804,N_24658,N_21774);
or U26805 (N_26805,N_23049,N_22192);
xor U26806 (N_26806,N_21261,N_21959);
and U26807 (N_26807,N_22729,N_22333);
xor U26808 (N_26808,N_20314,N_23662);
nand U26809 (N_26809,N_20526,N_21106);
nand U26810 (N_26810,N_22827,N_23467);
xor U26811 (N_26811,N_23151,N_24204);
xor U26812 (N_26812,N_21101,N_24661);
or U26813 (N_26813,N_21500,N_23521);
nor U26814 (N_26814,N_20242,N_24181);
nand U26815 (N_26815,N_20069,N_21809);
nor U26816 (N_26816,N_21644,N_21381);
and U26817 (N_26817,N_21265,N_22648);
and U26818 (N_26818,N_21630,N_23846);
or U26819 (N_26819,N_24053,N_20306);
or U26820 (N_26820,N_21395,N_21428);
nand U26821 (N_26821,N_21113,N_22715);
and U26822 (N_26822,N_23549,N_23232);
or U26823 (N_26823,N_21539,N_20939);
or U26824 (N_26824,N_22655,N_24279);
nand U26825 (N_26825,N_21165,N_24108);
nand U26826 (N_26826,N_21871,N_23143);
and U26827 (N_26827,N_21951,N_22554);
xor U26828 (N_26828,N_20901,N_23028);
or U26829 (N_26829,N_20470,N_24426);
nor U26830 (N_26830,N_21227,N_20015);
or U26831 (N_26831,N_24652,N_23252);
or U26832 (N_26832,N_21154,N_24913);
nand U26833 (N_26833,N_22876,N_21478);
xor U26834 (N_26834,N_20860,N_21676);
or U26835 (N_26835,N_24262,N_24174);
nor U26836 (N_26836,N_22811,N_22773);
and U26837 (N_26837,N_22194,N_24289);
nor U26838 (N_26838,N_20298,N_24804);
nor U26839 (N_26839,N_24580,N_23023);
nand U26840 (N_26840,N_21160,N_24894);
and U26841 (N_26841,N_21417,N_20659);
nor U26842 (N_26842,N_21329,N_23443);
or U26843 (N_26843,N_20002,N_24101);
nor U26844 (N_26844,N_22462,N_22836);
nor U26845 (N_26845,N_22187,N_20980);
and U26846 (N_26846,N_22624,N_21994);
and U26847 (N_26847,N_24232,N_23284);
and U26848 (N_26848,N_23413,N_23433);
and U26849 (N_26849,N_23441,N_24117);
nand U26850 (N_26850,N_21780,N_20683);
xor U26851 (N_26851,N_20212,N_21220);
or U26852 (N_26852,N_20671,N_21301);
nand U26853 (N_26853,N_22902,N_24523);
nor U26854 (N_26854,N_23336,N_20897);
and U26855 (N_26855,N_20634,N_23759);
and U26856 (N_26856,N_21448,N_21219);
nand U26857 (N_26857,N_24672,N_24802);
nand U26858 (N_26858,N_23273,N_24982);
or U26859 (N_26859,N_22211,N_24173);
xnor U26860 (N_26860,N_20599,N_24383);
nor U26861 (N_26861,N_23623,N_23781);
and U26862 (N_26862,N_22979,N_20992);
xnor U26863 (N_26863,N_22810,N_20963);
xor U26864 (N_26864,N_21830,N_22807);
nand U26865 (N_26865,N_23133,N_23022);
nand U26866 (N_26866,N_20328,N_20845);
nand U26867 (N_26867,N_24075,N_22189);
or U26868 (N_26868,N_22395,N_21311);
or U26869 (N_26869,N_22408,N_21497);
or U26870 (N_26870,N_23579,N_24964);
or U26871 (N_26871,N_24721,N_24518);
nor U26872 (N_26872,N_21845,N_24490);
and U26873 (N_26873,N_20301,N_21701);
and U26874 (N_26874,N_21903,N_24975);
and U26875 (N_26875,N_20253,N_21656);
xnor U26876 (N_26876,N_20709,N_24048);
or U26877 (N_26877,N_23480,N_24367);
nand U26878 (N_26878,N_22448,N_24020);
nor U26879 (N_26879,N_23928,N_23857);
nor U26880 (N_26880,N_22156,N_20669);
nor U26881 (N_26881,N_21836,N_22903);
and U26882 (N_26882,N_23155,N_23863);
nand U26883 (N_26883,N_23359,N_22654);
xnor U26884 (N_26884,N_22964,N_21312);
and U26885 (N_26885,N_24673,N_20064);
or U26886 (N_26886,N_20821,N_23942);
and U26887 (N_26887,N_22489,N_24320);
nand U26888 (N_26888,N_23140,N_23551);
and U26889 (N_26889,N_23270,N_20185);
nand U26890 (N_26890,N_21866,N_22019);
xnor U26891 (N_26891,N_20697,N_23993);
or U26892 (N_26892,N_23566,N_20853);
nand U26893 (N_26893,N_21288,N_24822);
or U26894 (N_26894,N_21123,N_24989);
and U26895 (N_26895,N_21393,N_23002);
nor U26896 (N_26896,N_20792,N_20555);
or U26897 (N_26897,N_20566,N_22591);
and U26898 (N_26898,N_20921,N_22691);
and U26899 (N_26899,N_23479,N_24873);
nand U26900 (N_26900,N_20366,N_24928);
nor U26901 (N_26901,N_24994,N_23035);
nor U26902 (N_26902,N_21709,N_24466);
and U26903 (N_26903,N_21579,N_24328);
nor U26904 (N_26904,N_23649,N_20756);
and U26905 (N_26905,N_21640,N_22220);
xor U26906 (N_26906,N_24664,N_24133);
xnor U26907 (N_26907,N_24896,N_22968);
xnor U26908 (N_26908,N_20102,N_21622);
nor U26909 (N_26909,N_20994,N_21583);
nor U26910 (N_26910,N_21443,N_24332);
and U26911 (N_26911,N_22656,N_22930);
and U26912 (N_26912,N_23915,N_22320);
xnor U26913 (N_26913,N_21435,N_22885);
or U26914 (N_26914,N_24863,N_23065);
nand U26915 (N_26915,N_23154,N_20416);
and U26916 (N_26916,N_22431,N_22628);
xnor U26917 (N_26917,N_22553,N_23457);
and U26918 (N_26918,N_20611,N_20761);
nor U26919 (N_26919,N_21731,N_22094);
or U26920 (N_26920,N_23390,N_22131);
nor U26921 (N_26921,N_23319,N_21596);
and U26922 (N_26922,N_21648,N_20176);
nor U26923 (N_26923,N_23726,N_23835);
nor U26924 (N_26924,N_20052,N_23141);
and U26925 (N_26925,N_24665,N_21685);
nand U26926 (N_26926,N_20080,N_24730);
or U26927 (N_26927,N_23225,N_21258);
xnor U26928 (N_26928,N_21532,N_21689);
or U26929 (N_26929,N_22750,N_22907);
and U26930 (N_26930,N_24595,N_23683);
xnor U26931 (N_26931,N_23234,N_24190);
nor U26932 (N_26932,N_24898,N_22734);
or U26933 (N_26933,N_21697,N_20899);
xor U26934 (N_26934,N_23800,N_22400);
or U26935 (N_26935,N_22994,N_23212);
nand U26936 (N_26936,N_24743,N_20106);
or U26937 (N_26937,N_20275,N_22897);
xor U26938 (N_26938,N_24021,N_22081);
nand U26939 (N_26939,N_21224,N_20837);
nand U26940 (N_26940,N_24327,N_21754);
nand U26941 (N_26941,N_24528,N_23733);
nor U26942 (N_26942,N_20206,N_24413);
xnor U26943 (N_26943,N_22916,N_22103);
xnor U26944 (N_26944,N_24717,N_24096);
nand U26945 (N_26945,N_24699,N_23600);
and U26946 (N_26946,N_22573,N_21750);
nor U26947 (N_26947,N_24039,N_24995);
nand U26948 (N_26948,N_20419,N_20876);
or U26949 (N_26949,N_24351,N_23950);
or U26950 (N_26950,N_23083,N_21467);
xor U26951 (N_26951,N_23302,N_24871);
and U26952 (N_26952,N_24416,N_24205);
nor U26953 (N_26953,N_23870,N_22147);
nand U26954 (N_26954,N_21991,N_22551);
or U26955 (N_26955,N_20806,N_20088);
nand U26956 (N_26956,N_23684,N_20734);
xor U26957 (N_26957,N_22741,N_20630);
nand U26958 (N_26958,N_22875,N_21506);
nand U26959 (N_26959,N_22664,N_24575);
nor U26960 (N_26960,N_20448,N_21186);
nor U26961 (N_26961,N_24823,N_22006);
or U26962 (N_26962,N_23017,N_22898);
xnor U26963 (N_26963,N_22054,N_23824);
xnor U26964 (N_26964,N_20661,N_21041);
xnor U26965 (N_26965,N_20143,N_20917);
or U26966 (N_26966,N_21011,N_24868);
and U26967 (N_26967,N_22830,N_24080);
or U26968 (N_26968,N_22225,N_24504);
nand U26969 (N_26969,N_20826,N_22290);
xor U26970 (N_26970,N_23786,N_23488);
or U26971 (N_26971,N_23995,N_21451);
nand U26972 (N_26972,N_22890,N_22355);
xor U26973 (N_26973,N_23044,N_24045);
or U26974 (N_26974,N_20797,N_23396);
and U26975 (N_26975,N_20741,N_22688);
xnor U26976 (N_26976,N_24627,N_23377);
or U26977 (N_26977,N_21747,N_23048);
or U26978 (N_26978,N_20793,N_20363);
or U26979 (N_26979,N_20795,N_24071);
nand U26980 (N_26980,N_20167,N_21849);
nand U26981 (N_26981,N_23431,N_24676);
nand U26982 (N_26982,N_24241,N_24690);
or U26983 (N_26983,N_22469,N_24834);
nor U26984 (N_26984,N_24855,N_22953);
nor U26985 (N_26985,N_23045,N_23904);
nand U26986 (N_26986,N_21236,N_21375);
xnor U26987 (N_26987,N_22181,N_21576);
nand U26988 (N_26988,N_23092,N_24411);
and U26989 (N_26989,N_21548,N_24140);
nor U26990 (N_26990,N_23717,N_24684);
nand U26991 (N_26991,N_23821,N_21027);
or U26992 (N_26992,N_22518,N_21365);
and U26993 (N_26993,N_23893,N_21863);
xnor U26994 (N_26994,N_24066,N_22461);
and U26995 (N_26995,N_21306,N_21976);
nand U26996 (N_26996,N_23771,N_21718);
or U26997 (N_26997,N_23062,N_20172);
nand U26998 (N_26998,N_20284,N_23736);
xnor U26999 (N_26999,N_24577,N_23323);
or U27000 (N_27000,N_23842,N_24585);
or U27001 (N_27001,N_20679,N_23716);
or U27002 (N_27002,N_22201,N_23110);
or U27003 (N_27003,N_24014,N_23817);
xor U27004 (N_27004,N_24257,N_20956);
nor U27005 (N_27005,N_21115,N_21734);
and U27006 (N_27006,N_24043,N_22350);
and U27007 (N_27007,N_21137,N_24356);
nand U27008 (N_27008,N_21617,N_21519);
nor U27009 (N_27009,N_22275,N_22575);
nor U27010 (N_27010,N_24017,N_23344);
nor U27011 (N_27011,N_20759,N_22451);
xnor U27012 (N_27012,N_24768,N_21411);
or U27013 (N_27013,N_20435,N_20311);
nand U27014 (N_27014,N_23820,N_23994);
and U27015 (N_27015,N_20739,N_21147);
or U27016 (N_27016,N_23679,N_24820);
xnor U27017 (N_27017,N_24298,N_20862);
xnor U27018 (N_27018,N_20239,N_22212);
or U27019 (N_27019,N_22942,N_22141);
xnor U27020 (N_27020,N_24081,N_21690);
nand U27021 (N_27021,N_23575,N_21309);
xor U27022 (N_27022,N_20114,N_24984);
nand U27023 (N_27023,N_20156,N_20847);
or U27024 (N_27024,N_21998,N_23021);
or U27025 (N_27025,N_22623,N_23720);
nor U27026 (N_27026,N_23656,N_21853);
nor U27027 (N_27027,N_24845,N_21562);
and U27028 (N_27028,N_22409,N_24348);
nor U27029 (N_27029,N_22712,N_23911);
nor U27030 (N_27030,N_22503,N_20888);
nor U27031 (N_27031,N_20645,N_21167);
xnor U27032 (N_27032,N_23869,N_20867);
nor U27033 (N_27033,N_24429,N_23018);
and U27034 (N_27034,N_22394,N_20701);
or U27035 (N_27035,N_23624,N_22234);
xnor U27036 (N_27036,N_23964,N_24163);
and U27037 (N_27037,N_22604,N_22111);
nor U27038 (N_27038,N_21935,N_22833);
xnor U27039 (N_27039,N_22570,N_22096);
nor U27040 (N_27040,N_22279,N_20865);
xnor U27041 (N_27041,N_22433,N_21755);
nor U27042 (N_27042,N_24235,N_24443);
or U27043 (N_27043,N_20972,N_24801);
nand U27044 (N_27044,N_22137,N_20815);
or U27045 (N_27045,N_22299,N_24799);
xnor U27046 (N_27046,N_20251,N_20754);
or U27047 (N_27047,N_21494,N_23200);
nor U27048 (N_27048,N_21176,N_23812);
or U27049 (N_27049,N_23761,N_24344);
nand U27050 (N_27050,N_22101,N_20582);
xor U27051 (N_27051,N_22542,N_20339);
and U27052 (N_27052,N_24629,N_20678);
or U27053 (N_27053,N_24254,N_21432);
nand U27054 (N_27054,N_23478,N_21653);
or U27055 (N_27055,N_20625,N_22967);
or U27056 (N_27056,N_22316,N_22888);
and U27057 (N_27057,N_21942,N_23454);
and U27058 (N_27058,N_24164,N_23215);
xnor U27059 (N_27059,N_23644,N_22673);
or U27060 (N_27060,N_20302,N_23597);
xor U27061 (N_27061,N_20261,N_22088);
and U27062 (N_27062,N_22905,N_21766);
xor U27063 (N_27063,N_24228,N_22369);
or U27064 (N_27064,N_23974,N_24394);
xnor U27065 (N_27065,N_22886,N_21695);
xnor U27066 (N_27066,N_21188,N_20219);
or U27067 (N_27067,N_22934,N_22801);
xnor U27068 (N_27068,N_21651,N_20890);
and U27069 (N_27069,N_24105,N_23917);
or U27070 (N_27070,N_21378,N_20927);
nor U27071 (N_27071,N_22685,N_20319);
or U27072 (N_27072,N_23052,N_24486);
or U27073 (N_27073,N_21655,N_23425);
xnor U27074 (N_27074,N_20676,N_23780);
nor U27075 (N_27075,N_22294,N_23810);
nand U27076 (N_27076,N_24529,N_22912);
or U27077 (N_27077,N_23894,N_20205);
nand U27078 (N_27078,N_24903,N_21013);
nand U27079 (N_27079,N_21217,N_24769);
nor U27080 (N_27080,N_22795,N_20588);
or U27081 (N_27081,N_21109,N_20039);
xor U27082 (N_27082,N_22760,N_23144);
xnor U27083 (N_27083,N_20365,N_20557);
and U27084 (N_27084,N_20280,N_22199);
or U27085 (N_27085,N_21334,N_21768);
or U27086 (N_27086,N_20801,N_24757);
and U27087 (N_27087,N_20226,N_24203);
nand U27088 (N_27088,N_22149,N_23422);
and U27089 (N_27089,N_20983,N_22634);
nand U27090 (N_27090,N_20478,N_21415);
xor U27091 (N_27091,N_22762,N_20241);
nand U27092 (N_27092,N_22410,N_22226);
xor U27093 (N_27093,N_22957,N_23383);
nor U27094 (N_27094,N_20480,N_22923);
and U27095 (N_27095,N_22227,N_24870);
and U27096 (N_27096,N_23834,N_24474);
nor U27097 (N_27097,N_24796,N_24904);
and U27098 (N_27098,N_21317,N_22309);
xor U27099 (N_27099,N_23352,N_21550);
or U27100 (N_27100,N_20702,N_21678);
or U27101 (N_27101,N_22564,N_24146);
nor U27102 (N_27102,N_22075,N_24278);
nand U27103 (N_27103,N_23877,N_24286);
xor U27104 (N_27104,N_21600,N_20690);
nand U27105 (N_27105,N_21152,N_23830);
nor U27106 (N_27106,N_24942,N_24888);
or U27107 (N_27107,N_22265,N_24208);
nand U27108 (N_27108,N_23222,N_20060);
xnor U27109 (N_27109,N_23126,N_21966);
and U27110 (N_27110,N_21776,N_20023);
or U27111 (N_27111,N_21670,N_23854);
or U27112 (N_27112,N_21742,N_23522);
nor U27113 (N_27113,N_22061,N_23082);
xnor U27114 (N_27114,N_21070,N_24638);
or U27115 (N_27115,N_23483,N_20166);
nand U27116 (N_27116,N_22420,N_24002);
xor U27117 (N_27117,N_21862,N_21342);
or U27118 (N_27118,N_23188,N_24909);
or U27119 (N_27119,N_23787,N_23084);
or U27120 (N_27120,N_21360,N_21913);
or U27121 (N_27121,N_24553,N_23156);
nor U27122 (N_27122,N_23439,N_20288);
or U27123 (N_27123,N_23832,N_21230);
nand U27124 (N_27124,N_21442,N_24200);
nand U27125 (N_27125,N_20414,N_23833);
or U27126 (N_27126,N_24460,N_24402);
nor U27127 (N_27127,N_23520,N_24022);
nand U27128 (N_27128,N_23404,N_22093);
xnor U27129 (N_27129,N_20107,N_20875);
or U27130 (N_27130,N_21211,N_20213);
nor U27131 (N_27131,N_20593,N_20066);
xnor U27132 (N_27132,N_20620,N_24251);
nor U27133 (N_27133,N_23749,N_21727);
xnor U27134 (N_27134,N_21316,N_20854);
nand U27135 (N_27135,N_22173,N_24625);
or U27136 (N_27136,N_24929,N_22844);
xor U27137 (N_27137,N_21129,N_24807);
nor U27138 (N_27138,N_20038,N_24669);
nor U27139 (N_27139,N_21659,N_22510);
nand U27140 (N_27140,N_21899,N_22308);
nor U27141 (N_27141,N_23206,N_23988);
or U27142 (N_27142,N_20085,N_23426);
nand U27143 (N_27143,N_23058,N_23532);
nor U27144 (N_27144,N_23734,N_24180);
and U27145 (N_27145,N_21710,N_24151);
nor U27146 (N_27146,N_21178,N_24240);
xor U27147 (N_27147,N_24797,N_21492);
nor U27148 (N_27148,N_20108,N_21010);
xor U27149 (N_27149,N_23080,N_21843);
nor U27150 (N_27150,N_24648,N_23281);
xnor U27151 (N_27151,N_24359,N_24640);
nand U27152 (N_27152,N_24459,N_24179);
nand U27153 (N_27153,N_20612,N_22301);
or U27154 (N_27154,N_23176,N_22492);
xor U27155 (N_27155,N_20558,N_23440);
nor U27156 (N_27156,N_21038,N_23647);
or U27157 (N_27157,N_24657,N_22966);
nor U27158 (N_27158,N_22362,N_22615);
xor U27159 (N_27159,N_24237,N_24885);
nand U27160 (N_27160,N_20117,N_20190);
nand U27161 (N_27161,N_23698,N_23117);
nor U27162 (N_27162,N_20149,N_24261);
nand U27163 (N_27163,N_23272,N_24069);
nor U27164 (N_27164,N_24890,N_21624);
nand U27165 (N_27165,N_23992,N_21985);
nand U27166 (N_27166,N_21662,N_22944);
and U27167 (N_27167,N_22214,N_22593);
nor U27168 (N_27168,N_21295,N_24976);
xnor U27169 (N_27169,N_21804,N_21705);
nand U27170 (N_27170,N_23455,N_24456);
nor U27171 (N_27171,N_22835,N_23486);
xor U27172 (N_27172,N_22713,N_24488);
or U27173 (N_27173,N_22640,N_21616);
nand U27174 (N_27174,N_24803,N_24739);
and U27175 (N_27175,N_20309,N_24901);
or U27176 (N_27176,N_24546,N_22119);
xor U27177 (N_27177,N_22339,N_21164);
or U27178 (N_27178,N_20272,N_20506);
nor U27179 (N_27179,N_20952,N_21030);
nor U27180 (N_27180,N_20894,N_20574);
or U27181 (N_27181,N_21156,N_21514);
and U27182 (N_27182,N_22704,N_22196);
or U27183 (N_27183,N_23933,N_22783);
and U27184 (N_27184,N_20127,N_20270);
nand U27185 (N_27185,N_21968,N_23625);
or U27186 (N_27186,N_24399,N_22157);
nand U27187 (N_27187,N_23598,N_23987);
or U27188 (N_27188,N_24812,N_22517);
and U27189 (N_27189,N_23718,N_20873);
xor U27190 (N_27190,N_23511,N_22280);
xnor U27191 (N_27191,N_22872,N_24304);
nor U27192 (N_27192,N_24646,N_23198);
and U27193 (N_27193,N_23073,N_20485);
xnor U27194 (N_27194,N_23692,N_21285);
or U27195 (N_27195,N_20711,N_20113);
nand U27196 (N_27196,N_24428,N_20221);
or U27197 (N_27197,N_24483,N_20381);
or U27198 (N_27198,N_21547,N_20655);
xor U27199 (N_27199,N_20390,N_23989);
and U27200 (N_27200,N_23921,N_22991);
xnor U27201 (N_27201,N_20505,N_20482);
nand U27202 (N_27202,N_23304,N_24956);
nand U27203 (N_27203,N_23116,N_21043);
nand U27204 (N_27204,N_20214,N_22248);
and U27205 (N_27205,N_22267,N_21552);
nand U27206 (N_27206,N_23162,N_24694);
nor U27207 (N_27207,N_20397,N_24744);
xnor U27208 (N_27208,N_24103,N_23459);
nor U27209 (N_27209,N_23954,N_22105);
or U27210 (N_27210,N_20354,N_23220);
nor U27211 (N_27211,N_21259,N_22097);
xor U27212 (N_27212,N_23577,N_20124);
or U27213 (N_27213,N_20040,N_20168);
nor U27214 (N_27214,N_24141,N_20913);
nand U27215 (N_27215,N_24346,N_21483);
or U27216 (N_27216,N_20003,N_21026);
and U27217 (N_27217,N_20981,N_22613);
xnor U27218 (N_27218,N_22965,N_22893);
nand U27219 (N_27219,N_23825,N_23768);
nor U27220 (N_27220,N_23233,N_24662);
nor U27221 (N_27221,N_21175,N_22925);
nor U27222 (N_27222,N_23025,N_24565);
or U27223 (N_27223,N_24271,N_21726);
or U27224 (N_27224,N_23414,N_22106);
or U27225 (N_27225,N_20392,N_21558);
and U27226 (N_27226,N_21816,N_24508);
or U27227 (N_27227,N_23376,N_22618);
nor U27228 (N_27228,N_22134,N_21163);
or U27229 (N_27229,N_24013,N_24365);
nand U27230 (N_27230,N_20839,N_20128);
nor U27231 (N_27231,N_20989,N_24613);
and U27232 (N_27232,N_20056,N_21473);
and U27233 (N_27233,N_23374,N_20006);
and U27234 (N_27234,N_20071,N_20527);
nor U27235 (N_27235,N_22166,N_23014);
and U27236 (N_27236,N_24255,N_24417);
xnor U27237 (N_27237,N_24301,N_21912);
xor U27238 (N_27238,N_24704,N_22561);
nand U27239 (N_27239,N_20871,N_21744);
nor U27240 (N_27240,N_22092,N_23321);
or U27241 (N_27241,N_22977,N_22786);
nor U27242 (N_27242,N_23218,N_24749);
or U27243 (N_27243,N_24082,N_22285);
nor U27244 (N_27244,N_20519,N_23582);
nand U27245 (N_27245,N_24256,N_24551);
nand U27246 (N_27246,N_20746,N_21650);
xnor U27247 (N_27247,N_20051,N_20472);
and U27248 (N_27248,N_20074,N_21578);
nor U27249 (N_27249,N_21232,N_23962);
or U27250 (N_27250,N_20787,N_22057);
or U27251 (N_27251,N_21965,N_22167);
or U27252 (N_27252,N_21613,N_23689);
xnor U27253 (N_27253,N_22452,N_24499);
xor U27254 (N_27254,N_24947,N_24500);
and U27255 (N_27255,N_22766,N_20491);
and U27256 (N_27256,N_20408,N_22396);
and U27257 (N_27257,N_24805,N_23397);
xor U27258 (N_27258,N_23432,N_24571);
nor U27259 (N_27259,N_22569,N_20296);
and U27260 (N_27260,N_20262,N_24569);
or U27261 (N_27261,N_21708,N_22442);
nor U27262 (N_27262,N_21007,N_23975);
and U27263 (N_27263,N_22782,N_20353);
nand U27264 (N_27264,N_22475,N_24130);
nand U27265 (N_27265,N_23622,N_24506);
nor U27266 (N_27266,N_24937,N_22063);
xnor U27267 (N_27267,N_20608,N_20227);
xor U27268 (N_27268,N_24263,N_24728);
nand U27269 (N_27269,N_20843,N_24052);
and U27270 (N_27270,N_22190,N_22243);
and U27271 (N_27271,N_24447,N_23606);
or U27272 (N_27272,N_21511,N_23923);
and U27273 (N_27273,N_23779,N_24899);
nor U27274 (N_27274,N_24455,N_21405);
xor U27275 (N_27275,N_20966,N_21015);
nor U27276 (N_27276,N_23437,N_22392);
nor U27277 (N_27277,N_20393,N_22371);
and U27278 (N_27278,N_24425,N_22470);
nand U27279 (N_27279,N_24561,N_23738);
or U27280 (N_27280,N_23701,N_21361);
nand U27281 (N_27281,N_24353,N_22558);
and U27282 (N_27282,N_20528,N_24009);
nand U27283 (N_27283,N_24226,N_20827);
and U27284 (N_27284,N_22445,N_20177);
or U27285 (N_27285,N_24260,N_22153);
or U27286 (N_27286,N_20896,N_24225);
and U27287 (N_27287,N_24341,N_21076);
nor U27288 (N_27288,N_22202,N_20580);
nor U27289 (N_27289,N_21882,N_24925);
or U27290 (N_27290,N_20613,N_24602);
and U27291 (N_27291,N_23125,N_23451);
nand U27292 (N_27292,N_23855,N_23559);
nand U27293 (N_27293,N_21336,N_21470);
and U27294 (N_27294,N_24209,N_23719);
xnor U27295 (N_27295,N_20147,N_24723);
and U27296 (N_27296,N_20097,N_23466);
or U27297 (N_27297,N_20559,N_21169);
xor U27298 (N_27298,N_20563,N_21421);
and U27299 (N_27299,N_24231,N_23502);
nor U27300 (N_27300,N_23391,N_24026);
nand U27301 (N_27301,N_24153,N_21954);
and U27302 (N_27302,N_21146,N_22367);
xnor U27303 (N_27303,N_22317,N_23420);
nand U27304 (N_27304,N_20497,N_20089);
nor U27305 (N_27305,N_20359,N_23617);
xnor U27306 (N_27306,N_20597,N_24615);
or U27307 (N_27307,N_24724,N_22791);
and U27308 (N_27308,N_22778,N_20887);
or U27309 (N_27309,N_21916,N_21791);
nor U27310 (N_27310,N_23608,N_21593);
or U27311 (N_27311,N_20063,N_23040);
or U27312 (N_27312,N_23636,N_22302);
or U27313 (N_27313,N_24526,N_23326);
and U27314 (N_27314,N_23246,N_23848);
nor U27315 (N_27315,N_24326,N_20604);
and U27316 (N_27316,N_24310,N_24543);
and U27317 (N_27317,N_21042,N_22818);
nor U27318 (N_27318,N_23250,N_20629);
or U27319 (N_27319,N_23795,N_21757);
and U27320 (N_27320,N_22684,N_22568);
or U27321 (N_27321,N_20372,N_23751);
nand U27322 (N_27322,N_21722,N_20964);
nor U27323 (N_27323,N_24210,N_21324);
xnor U27324 (N_27324,N_21085,N_23700);
xor U27325 (N_27325,N_20530,N_24380);
and U27326 (N_27326,N_21525,N_21385);
and U27327 (N_27327,N_24740,N_21456);
or U27328 (N_27328,N_20808,N_23262);
xnor U27329 (N_27329,N_24943,N_23862);
xnor U27330 (N_27330,N_24126,N_20250);
nand U27331 (N_27331,N_21251,N_21549);
and U27332 (N_27332,N_20154,N_23146);
nand U27333 (N_27333,N_21474,N_21674);
nand U27334 (N_27334,N_20938,N_24772);
and U27335 (N_27335,N_21256,N_21601);
nor U27336 (N_27336,N_23446,N_20830);
nand U27337 (N_27337,N_20569,N_23192);
nor U27338 (N_27338,N_24631,N_24916);
nor U27339 (N_27339,N_23773,N_21993);
xnor U27340 (N_27340,N_24653,N_24239);
xnor U27341 (N_27341,N_22913,N_20462);
or U27342 (N_27342,N_21602,N_24019);
nor U27343 (N_27343,N_21590,N_20825);
nor U27344 (N_27344,N_22466,N_23941);
xor U27345 (N_27345,N_21873,N_24192);
and U27346 (N_27346,N_21551,N_20303);
xor U27347 (N_27347,N_24742,N_23686);
xor U27348 (N_27348,N_22529,N_23887);
and U27349 (N_27349,N_23320,N_21284);
xor U27350 (N_27350,N_23668,N_23354);
nand U27351 (N_27351,N_20492,N_23447);
and U27352 (N_27352,N_24064,N_24513);
nand U27353 (N_27353,N_24485,N_22036);
nand U27354 (N_27354,N_21975,N_24536);
and U27355 (N_27355,N_23299,N_20396);
nor U27356 (N_27356,N_24220,N_24927);
nand U27357 (N_27357,N_20498,N_21941);
or U27358 (N_27358,N_21339,N_21536);
xor U27359 (N_27359,N_24503,N_20910);
xor U27360 (N_27360,N_23831,N_24965);
and U27361 (N_27361,N_21239,N_23095);
nor U27362 (N_27362,N_24343,N_22224);
or U27363 (N_27363,N_22677,N_24188);
xnor U27364 (N_27364,N_21296,N_24800);
or U27365 (N_27365,N_20404,N_24784);
or U27366 (N_27366,N_24707,N_20092);
nand U27367 (N_27367,N_22139,N_21840);
or U27368 (N_27368,N_22453,N_24216);
and U27369 (N_27369,N_22632,N_21044);
or U27370 (N_27370,N_20005,N_20732);
nand U27371 (N_27371,N_22183,N_20773);
nand U27372 (N_27372,N_23491,N_24810);
nand U27373 (N_27373,N_24692,N_20014);
xnor U27374 (N_27374,N_20975,N_20324);
or U27375 (N_27375,N_23241,N_22813);
nor U27376 (N_27376,N_23843,N_23538);
or U27377 (N_27377,N_22009,N_24516);
nand U27378 (N_27378,N_21522,N_24407);
xor U27379 (N_27379,N_20621,N_22497);
and U27380 (N_27380,N_24962,N_23913);
nand U27381 (N_27381,N_24702,N_20687);
nor U27382 (N_27382,N_21185,N_23612);
and U27383 (N_27383,N_21723,N_23809);
or U27384 (N_27384,N_23940,N_22582);
nor U27385 (N_27385,N_20704,N_20923);
and U27386 (N_27386,N_21505,N_24337);
xnor U27387 (N_27387,N_23574,N_21426);
or U27388 (N_27388,N_23178,N_22418);
or U27389 (N_27389,N_20218,N_22163);
nand U27390 (N_27390,N_20691,N_21910);
nor U27391 (N_27391,N_24016,N_20401);
xnor U27392 (N_27392,N_20926,N_23576);
xor U27393 (N_27393,N_20664,N_21019);
nor U27394 (N_27394,N_24922,N_24521);
and U27395 (N_27395,N_24398,N_20022);
nor U27396 (N_27396,N_22547,N_22533);
and U27397 (N_27397,N_21124,N_21538);
and U27398 (N_27398,N_20884,N_21437);
nand U27399 (N_27399,N_22660,N_21711);
or U27400 (N_27400,N_21066,N_23211);
and U27401 (N_27401,N_22069,N_21628);
xnor U27402 (N_27402,N_21799,N_23918);
nand U27403 (N_27403,N_22577,N_20140);
nand U27404 (N_27404,N_22587,N_20777);
xor U27405 (N_27405,N_24911,N_22256);
nand U27406 (N_27406,N_23682,N_24514);
nor U27407 (N_27407,N_22589,N_21384);
xnor U27408 (N_27408,N_24630,N_23411);
and U27409 (N_27409,N_23907,N_20238);
nor U27410 (N_27410,N_23179,N_23540);
and U27411 (N_27411,N_23254,N_24502);
and U27412 (N_27412,N_20007,N_20259);
and U27413 (N_27413,N_20551,N_21925);
nand U27414 (N_27414,N_22297,N_22851);
nor U27415 (N_27415,N_23610,N_22933);
nor U27416 (N_27416,N_22730,N_23033);
and U27417 (N_27417,N_22829,N_23838);
or U27418 (N_27418,N_24099,N_22342);
or U27419 (N_27419,N_21358,N_22719);
or U27420 (N_27420,N_20159,N_20255);
xor U27421 (N_27421,N_22509,N_23099);
xor U27422 (N_27422,N_23562,N_22197);
nor U27423 (N_27423,N_21111,N_24782);
or U27424 (N_27424,N_20713,N_23565);
nor U27425 (N_27425,N_24663,N_20874);
nor U27426 (N_27426,N_23847,N_22693);
and U27427 (N_27427,N_21909,N_20164);
nor U27428 (N_27428,N_24461,N_23554);
nand U27429 (N_27429,N_24884,N_20417);
xor U27430 (N_27430,N_24593,N_23101);
nor U27431 (N_27431,N_20278,N_23722);
nand U27432 (N_27432,N_23379,N_23031);
nand U27433 (N_27433,N_23346,N_24207);
or U27434 (N_27434,N_23481,N_24980);
nand U27435 (N_27435,N_22919,N_23568);
xnor U27436 (N_27436,N_23385,N_20327);
and U27437 (N_27437,N_23727,N_21512);
nand U27438 (N_27438,N_23711,N_23552);
nor U27439 (N_27439,N_20811,N_22493);
and U27440 (N_27440,N_22732,N_20937);
and U27441 (N_27441,N_23762,N_23016);
nand U27442 (N_27442,N_22266,N_22490);
or U27443 (N_27443,N_23977,N_21420);
xor U27444 (N_27444,N_23415,N_23054);
xor U27445 (N_27445,N_22411,N_23201);
xnor U27446 (N_27446,N_24959,N_21582);
nand U27447 (N_27447,N_23371,N_22387);
and U27448 (N_27448,N_20018,N_21629);
nand U27449 (N_27449,N_21260,N_22659);
nand U27450 (N_27450,N_20441,N_24788);
or U27451 (N_27451,N_21997,N_21462);
xnor U27452 (N_27452,N_20084,N_23503);
or U27453 (N_27453,N_22928,N_23785);
nor U27454 (N_27454,N_20960,N_24628);
or U27455 (N_27455,N_23929,N_23357);
xor U27456 (N_27456,N_22946,N_21244);
nand U27457 (N_27457,N_24541,N_20870);
xor U27458 (N_27458,N_22696,N_20771);
nor U27459 (N_27459,N_22246,N_23669);
nand U27460 (N_27460,N_21516,N_20318);
xnor U27461 (N_27461,N_24373,N_23177);
nand U27462 (N_27462,N_24589,N_23055);
or U27463 (N_27463,N_24840,N_24557);
or U27464 (N_27464,N_21036,N_23936);
nor U27465 (N_27465,N_21391,N_21647);
or U27466 (N_27466,N_21238,N_24362);
nand U27467 (N_27467,N_20279,N_21114);
xnor U27468 (N_27468,N_23173,N_23378);
and U27469 (N_27469,N_23169,N_24620);
xnor U27470 (N_27470,N_21241,N_21575);
or U27471 (N_27471,N_20269,N_23971);
or U27472 (N_27472,N_23563,N_22311);
and U27473 (N_27473,N_22982,N_23897);
xor U27474 (N_27474,N_20812,N_24681);
and U27475 (N_27475,N_23515,N_23157);
and U27476 (N_27476,N_20831,N_20647);
nand U27477 (N_27477,N_21322,N_24201);
nand U27478 (N_27478,N_22508,N_24144);
nor U27479 (N_27479,N_24908,N_23384);
or U27480 (N_27480,N_22780,N_24520);
and U27481 (N_27481,N_24883,N_21191);
nand U27482 (N_27482,N_20882,N_23813);
nand U27483 (N_27483,N_22745,N_22328);
and U27484 (N_27484,N_21495,N_20207);
nor U27485 (N_27485,N_20872,N_24552);
xnor U27486 (N_27486,N_20776,N_20750);
xor U27487 (N_27487,N_22179,N_21326);
and U27488 (N_27488,N_24973,N_23983);
nand U27489 (N_27489,N_22880,N_24178);
nand U27490 (N_27490,N_24121,N_23985);
and U27491 (N_27491,N_24498,N_23860);
or U27492 (N_27492,N_20494,N_23837);
nand U27493 (N_27493,N_20331,N_23746);
nor U27494 (N_27494,N_23753,N_23081);
nor U27495 (N_27495,N_21349,N_21034);
and U27496 (N_27496,N_24851,N_20475);
xor U27497 (N_27497,N_22896,N_22565);
nor U27498 (N_27498,N_24029,N_24038);
or U27499 (N_27499,N_24957,N_23849);
nor U27500 (N_27500,N_22593,N_24385);
or U27501 (N_27501,N_23847,N_22477);
or U27502 (N_27502,N_22639,N_20765);
xnor U27503 (N_27503,N_23595,N_21123);
or U27504 (N_27504,N_23885,N_20695);
xor U27505 (N_27505,N_22785,N_23134);
nor U27506 (N_27506,N_24231,N_23215);
nor U27507 (N_27507,N_22591,N_24104);
xnor U27508 (N_27508,N_24953,N_23441);
xor U27509 (N_27509,N_22143,N_24335);
nand U27510 (N_27510,N_23606,N_22796);
and U27511 (N_27511,N_23827,N_20552);
nor U27512 (N_27512,N_24372,N_23806);
nand U27513 (N_27513,N_24680,N_22029);
and U27514 (N_27514,N_22336,N_24703);
xor U27515 (N_27515,N_20665,N_24693);
xor U27516 (N_27516,N_23823,N_21283);
and U27517 (N_27517,N_23188,N_20162);
nand U27518 (N_27518,N_24601,N_22206);
and U27519 (N_27519,N_20723,N_23369);
or U27520 (N_27520,N_22562,N_24344);
xnor U27521 (N_27521,N_22196,N_20162);
and U27522 (N_27522,N_24715,N_24739);
nor U27523 (N_27523,N_21991,N_23414);
nor U27524 (N_27524,N_23394,N_23583);
and U27525 (N_27525,N_24701,N_21562);
nand U27526 (N_27526,N_20408,N_24687);
nor U27527 (N_27527,N_24516,N_24734);
or U27528 (N_27528,N_21344,N_24692);
xnor U27529 (N_27529,N_21488,N_24613);
nand U27530 (N_27530,N_21356,N_21747);
nor U27531 (N_27531,N_22654,N_24578);
or U27532 (N_27532,N_23973,N_24697);
nor U27533 (N_27533,N_22575,N_24784);
nor U27534 (N_27534,N_21386,N_22287);
and U27535 (N_27535,N_23797,N_23985);
nand U27536 (N_27536,N_22660,N_21915);
and U27537 (N_27537,N_24687,N_22842);
nand U27538 (N_27538,N_24499,N_24235);
xor U27539 (N_27539,N_23234,N_20365);
and U27540 (N_27540,N_23873,N_21506);
nand U27541 (N_27541,N_20324,N_24932);
nand U27542 (N_27542,N_22974,N_23356);
nand U27543 (N_27543,N_21257,N_20525);
and U27544 (N_27544,N_22301,N_21934);
xor U27545 (N_27545,N_22860,N_21003);
or U27546 (N_27546,N_22051,N_22114);
and U27547 (N_27547,N_23513,N_23392);
nand U27548 (N_27548,N_20428,N_20734);
nor U27549 (N_27549,N_21896,N_20430);
nor U27550 (N_27550,N_22409,N_24719);
nor U27551 (N_27551,N_23701,N_21116);
nor U27552 (N_27552,N_23481,N_22166);
nor U27553 (N_27553,N_23759,N_22380);
xor U27554 (N_27554,N_23256,N_22439);
and U27555 (N_27555,N_23689,N_23421);
or U27556 (N_27556,N_20743,N_22374);
nand U27557 (N_27557,N_20153,N_21156);
xnor U27558 (N_27558,N_22259,N_20147);
nand U27559 (N_27559,N_20583,N_22532);
or U27560 (N_27560,N_20621,N_24331);
and U27561 (N_27561,N_21238,N_21176);
nor U27562 (N_27562,N_21297,N_24839);
nand U27563 (N_27563,N_24755,N_23316);
xor U27564 (N_27564,N_21440,N_24592);
nand U27565 (N_27565,N_20319,N_23152);
xnor U27566 (N_27566,N_21721,N_24269);
and U27567 (N_27567,N_21717,N_24783);
nand U27568 (N_27568,N_23619,N_23648);
xor U27569 (N_27569,N_24325,N_21787);
xnor U27570 (N_27570,N_20616,N_21650);
nand U27571 (N_27571,N_23353,N_22336);
nand U27572 (N_27572,N_20625,N_21087);
or U27573 (N_27573,N_22139,N_22073);
and U27574 (N_27574,N_24051,N_20287);
and U27575 (N_27575,N_23228,N_20783);
and U27576 (N_27576,N_20715,N_23384);
xor U27577 (N_27577,N_22210,N_21866);
and U27578 (N_27578,N_24329,N_24371);
nor U27579 (N_27579,N_21966,N_20636);
xor U27580 (N_27580,N_24656,N_22372);
nor U27581 (N_27581,N_22347,N_24457);
xor U27582 (N_27582,N_21295,N_22605);
nor U27583 (N_27583,N_21621,N_20836);
nor U27584 (N_27584,N_21420,N_20434);
xor U27585 (N_27585,N_20945,N_24977);
nand U27586 (N_27586,N_23450,N_24322);
xnor U27587 (N_27587,N_22679,N_24698);
nor U27588 (N_27588,N_22649,N_20708);
or U27589 (N_27589,N_23768,N_22597);
nand U27590 (N_27590,N_22989,N_21841);
and U27591 (N_27591,N_22025,N_20706);
nand U27592 (N_27592,N_24936,N_20540);
and U27593 (N_27593,N_20510,N_24660);
nand U27594 (N_27594,N_24651,N_24950);
xor U27595 (N_27595,N_22462,N_23980);
nor U27596 (N_27596,N_24775,N_21207);
nor U27597 (N_27597,N_22416,N_20469);
nor U27598 (N_27598,N_20094,N_22414);
nand U27599 (N_27599,N_24774,N_24104);
xnor U27600 (N_27600,N_24155,N_20689);
or U27601 (N_27601,N_21558,N_22335);
nand U27602 (N_27602,N_21230,N_23732);
nor U27603 (N_27603,N_22463,N_20824);
and U27604 (N_27604,N_20190,N_21508);
xor U27605 (N_27605,N_20945,N_20069);
nor U27606 (N_27606,N_21035,N_22686);
nand U27607 (N_27607,N_24466,N_21838);
or U27608 (N_27608,N_21885,N_20903);
or U27609 (N_27609,N_22726,N_21122);
and U27610 (N_27610,N_20124,N_24313);
nand U27611 (N_27611,N_22785,N_22137);
xor U27612 (N_27612,N_24152,N_22783);
nand U27613 (N_27613,N_22080,N_24805);
or U27614 (N_27614,N_24978,N_24411);
and U27615 (N_27615,N_24407,N_22568);
and U27616 (N_27616,N_21660,N_22570);
nor U27617 (N_27617,N_24902,N_22811);
nand U27618 (N_27618,N_22921,N_23594);
nand U27619 (N_27619,N_22805,N_22196);
or U27620 (N_27620,N_21182,N_20108);
and U27621 (N_27621,N_24311,N_24643);
xor U27622 (N_27622,N_23881,N_24498);
or U27623 (N_27623,N_23531,N_23324);
and U27624 (N_27624,N_23792,N_21801);
nand U27625 (N_27625,N_21562,N_22855);
xnor U27626 (N_27626,N_21548,N_22887);
and U27627 (N_27627,N_21323,N_21680);
and U27628 (N_27628,N_21760,N_20893);
or U27629 (N_27629,N_24413,N_22896);
and U27630 (N_27630,N_23750,N_24146);
and U27631 (N_27631,N_23191,N_23945);
nand U27632 (N_27632,N_23457,N_21295);
and U27633 (N_27633,N_21335,N_24113);
xor U27634 (N_27634,N_23687,N_24020);
nor U27635 (N_27635,N_20336,N_21011);
and U27636 (N_27636,N_22706,N_23812);
or U27637 (N_27637,N_23923,N_22719);
and U27638 (N_27638,N_22040,N_23419);
or U27639 (N_27639,N_23815,N_24568);
or U27640 (N_27640,N_21637,N_22963);
or U27641 (N_27641,N_23688,N_23047);
or U27642 (N_27642,N_21124,N_21143);
xor U27643 (N_27643,N_24377,N_20534);
or U27644 (N_27644,N_20535,N_23467);
and U27645 (N_27645,N_21851,N_23876);
or U27646 (N_27646,N_20088,N_23219);
and U27647 (N_27647,N_24999,N_22542);
nand U27648 (N_27648,N_22713,N_24626);
nor U27649 (N_27649,N_23004,N_20367);
or U27650 (N_27650,N_24553,N_24009);
nor U27651 (N_27651,N_22052,N_21324);
or U27652 (N_27652,N_22544,N_23853);
and U27653 (N_27653,N_21624,N_24945);
xnor U27654 (N_27654,N_21600,N_21500);
or U27655 (N_27655,N_20961,N_24479);
xor U27656 (N_27656,N_24824,N_21999);
and U27657 (N_27657,N_23840,N_20514);
or U27658 (N_27658,N_22422,N_23286);
xnor U27659 (N_27659,N_21089,N_24962);
nor U27660 (N_27660,N_20884,N_23014);
or U27661 (N_27661,N_22265,N_22954);
or U27662 (N_27662,N_22327,N_23419);
nor U27663 (N_27663,N_22814,N_24962);
and U27664 (N_27664,N_21243,N_24492);
xor U27665 (N_27665,N_20704,N_22383);
xor U27666 (N_27666,N_23886,N_24068);
xor U27667 (N_27667,N_23675,N_23822);
nor U27668 (N_27668,N_23854,N_21124);
nor U27669 (N_27669,N_23443,N_23765);
nor U27670 (N_27670,N_20435,N_20116);
nor U27671 (N_27671,N_24520,N_21058);
and U27672 (N_27672,N_22665,N_24214);
or U27673 (N_27673,N_20543,N_24380);
nor U27674 (N_27674,N_22267,N_20464);
nand U27675 (N_27675,N_20971,N_21999);
and U27676 (N_27676,N_24351,N_24969);
nand U27677 (N_27677,N_24218,N_24802);
nor U27678 (N_27678,N_23030,N_24996);
nor U27679 (N_27679,N_24734,N_21134);
nand U27680 (N_27680,N_24651,N_24814);
xnor U27681 (N_27681,N_24844,N_23559);
and U27682 (N_27682,N_23511,N_23385);
and U27683 (N_27683,N_24748,N_22741);
or U27684 (N_27684,N_24518,N_21210);
nand U27685 (N_27685,N_20238,N_24216);
or U27686 (N_27686,N_23899,N_21758);
nand U27687 (N_27687,N_24431,N_21477);
nand U27688 (N_27688,N_21035,N_21250);
and U27689 (N_27689,N_20627,N_23106);
xor U27690 (N_27690,N_20756,N_22396);
and U27691 (N_27691,N_21912,N_20269);
xnor U27692 (N_27692,N_21490,N_22795);
nand U27693 (N_27693,N_23462,N_21906);
nand U27694 (N_27694,N_24540,N_23745);
nand U27695 (N_27695,N_20441,N_22789);
nand U27696 (N_27696,N_21422,N_22789);
nor U27697 (N_27697,N_21797,N_24542);
or U27698 (N_27698,N_23370,N_24355);
xnor U27699 (N_27699,N_24524,N_20408);
nand U27700 (N_27700,N_22495,N_23313);
xnor U27701 (N_27701,N_21569,N_23491);
xor U27702 (N_27702,N_20424,N_23047);
or U27703 (N_27703,N_22581,N_21750);
and U27704 (N_27704,N_20214,N_24416);
nor U27705 (N_27705,N_21326,N_20580);
and U27706 (N_27706,N_23665,N_21134);
or U27707 (N_27707,N_23743,N_23949);
nor U27708 (N_27708,N_24906,N_23223);
or U27709 (N_27709,N_21465,N_24754);
nor U27710 (N_27710,N_20384,N_22319);
nand U27711 (N_27711,N_24542,N_22401);
or U27712 (N_27712,N_24471,N_24642);
xnor U27713 (N_27713,N_21746,N_24522);
and U27714 (N_27714,N_22462,N_22636);
xnor U27715 (N_27715,N_24064,N_23556);
xor U27716 (N_27716,N_22074,N_23559);
and U27717 (N_27717,N_21209,N_21526);
xor U27718 (N_27718,N_24675,N_23227);
or U27719 (N_27719,N_24600,N_22129);
xor U27720 (N_27720,N_22817,N_20613);
xnor U27721 (N_27721,N_24147,N_21130);
or U27722 (N_27722,N_24291,N_23504);
or U27723 (N_27723,N_20065,N_23736);
xor U27724 (N_27724,N_24379,N_21869);
xnor U27725 (N_27725,N_24117,N_24555);
or U27726 (N_27726,N_22928,N_24778);
xor U27727 (N_27727,N_23281,N_22409);
and U27728 (N_27728,N_22120,N_22541);
nor U27729 (N_27729,N_24981,N_20426);
nor U27730 (N_27730,N_22239,N_22123);
or U27731 (N_27731,N_24970,N_23161);
or U27732 (N_27732,N_21672,N_21233);
nor U27733 (N_27733,N_22280,N_20254);
xnor U27734 (N_27734,N_24221,N_20051);
nand U27735 (N_27735,N_21184,N_24020);
or U27736 (N_27736,N_24348,N_24529);
xor U27737 (N_27737,N_20244,N_20678);
nand U27738 (N_27738,N_24096,N_21088);
and U27739 (N_27739,N_20494,N_22973);
xor U27740 (N_27740,N_21442,N_22982);
or U27741 (N_27741,N_23949,N_23563);
or U27742 (N_27742,N_24730,N_23567);
and U27743 (N_27743,N_21038,N_20594);
and U27744 (N_27744,N_22441,N_21584);
nand U27745 (N_27745,N_22716,N_21510);
nor U27746 (N_27746,N_20714,N_20327);
nand U27747 (N_27747,N_22661,N_22901);
and U27748 (N_27748,N_20737,N_24730);
nand U27749 (N_27749,N_23389,N_23963);
nand U27750 (N_27750,N_22662,N_20777);
and U27751 (N_27751,N_24001,N_24152);
nand U27752 (N_27752,N_22827,N_22148);
nand U27753 (N_27753,N_23030,N_20923);
xnor U27754 (N_27754,N_20724,N_21680);
and U27755 (N_27755,N_23679,N_23584);
nand U27756 (N_27756,N_21712,N_21681);
xnor U27757 (N_27757,N_23069,N_23789);
nor U27758 (N_27758,N_20851,N_20498);
xor U27759 (N_27759,N_20827,N_20980);
nor U27760 (N_27760,N_20552,N_20823);
nand U27761 (N_27761,N_22089,N_23725);
nor U27762 (N_27762,N_20911,N_24720);
and U27763 (N_27763,N_20139,N_21423);
xnor U27764 (N_27764,N_22636,N_21018);
or U27765 (N_27765,N_22572,N_23560);
xor U27766 (N_27766,N_20199,N_22532);
and U27767 (N_27767,N_22786,N_22587);
and U27768 (N_27768,N_21823,N_23898);
nor U27769 (N_27769,N_24766,N_23384);
nand U27770 (N_27770,N_22149,N_22675);
or U27771 (N_27771,N_24752,N_22882);
and U27772 (N_27772,N_20041,N_23979);
nor U27773 (N_27773,N_24736,N_21990);
or U27774 (N_27774,N_20693,N_23417);
nor U27775 (N_27775,N_21031,N_24625);
nor U27776 (N_27776,N_23234,N_21217);
or U27777 (N_27777,N_22856,N_22284);
and U27778 (N_27778,N_21913,N_22904);
and U27779 (N_27779,N_23920,N_24320);
nor U27780 (N_27780,N_21401,N_23698);
nor U27781 (N_27781,N_20770,N_20395);
xor U27782 (N_27782,N_22964,N_20207);
nor U27783 (N_27783,N_22726,N_20120);
or U27784 (N_27784,N_23227,N_24066);
nand U27785 (N_27785,N_21648,N_20964);
xnor U27786 (N_27786,N_24957,N_22521);
nand U27787 (N_27787,N_22680,N_22601);
xnor U27788 (N_27788,N_24458,N_24824);
nor U27789 (N_27789,N_24061,N_24605);
nand U27790 (N_27790,N_20310,N_23852);
or U27791 (N_27791,N_24271,N_20471);
nand U27792 (N_27792,N_23755,N_21986);
and U27793 (N_27793,N_23024,N_20509);
xnor U27794 (N_27794,N_20040,N_20787);
nand U27795 (N_27795,N_23923,N_20757);
and U27796 (N_27796,N_23865,N_20419);
nor U27797 (N_27797,N_20725,N_23348);
nor U27798 (N_27798,N_21238,N_20323);
xor U27799 (N_27799,N_23300,N_20297);
or U27800 (N_27800,N_24241,N_24229);
nand U27801 (N_27801,N_22754,N_21380);
and U27802 (N_27802,N_20575,N_23422);
xor U27803 (N_27803,N_20427,N_21872);
xnor U27804 (N_27804,N_21632,N_20063);
or U27805 (N_27805,N_21396,N_21950);
nand U27806 (N_27806,N_22984,N_23275);
nor U27807 (N_27807,N_20543,N_22380);
and U27808 (N_27808,N_23304,N_20101);
nor U27809 (N_27809,N_24017,N_22618);
or U27810 (N_27810,N_22266,N_23199);
xnor U27811 (N_27811,N_23128,N_22311);
nor U27812 (N_27812,N_24692,N_20054);
xor U27813 (N_27813,N_24525,N_23278);
xnor U27814 (N_27814,N_23988,N_21149);
nor U27815 (N_27815,N_20928,N_24845);
xor U27816 (N_27816,N_21209,N_20408);
nor U27817 (N_27817,N_20609,N_21304);
nand U27818 (N_27818,N_21396,N_24659);
nor U27819 (N_27819,N_23496,N_22997);
or U27820 (N_27820,N_22243,N_23759);
xor U27821 (N_27821,N_20144,N_20098);
nand U27822 (N_27822,N_21357,N_22071);
xnor U27823 (N_27823,N_20924,N_23158);
xnor U27824 (N_27824,N_24109,N_22074);
and U27825 (N_27825,N_20355,N_20663);
xor U27826 (N_27826,N_24383,N_22047);
xor U27827 (N_27827,N_24902,N_21181);
nor U27828 (N_27828,N_20420,N_22980);
and U27829 (N_27829,N_22381,N_23406);
nor U27830 (N_27830,N_22613,N_23214);
and U27831 (N_27831,N_20180,N_22832);
nand U27832 (N_27832,N_23613,N_21120);
or U27833 (N_27833,N_22459,N_22858);
nand U27834 (N_27834,N_21158,N_20991);
nor U27835 (N_27835,N_22049,N_24787);
xor U27836 (N_27836,N_20216,N_20859);
nand U27837 (N_27837,N_23273,N_24123);
nor U27838 (N_27838,N_22509,N_20667);
nor U27839 (N_27839,N_21503,N_24668);
nand U27840 (N_27840,N_24818,N_21751);
nor U27841 (N_27841,N_20838,N_20654);
nand U27842 (N_27842,N_20097,N_23396);
xor U27843 (N_27843,N_23724,N_22588);
or U27844 (N_27844,N_22976,N_22093);
nand U27845 (N_27845,N_20765,N_22783);
and U27846 (N_27846,N_22108,N_23641);
and U27847 (N_27847,N_23895,N_23359);
xnor U27848 (N_27848,N_22969,N_24615);
nor U27849 (N_27849,N_23434,N_23373);
and U27850 (N_27850,N_23213,N_23445);
or U27851 (N_27851,N_22566,N_24691);
nor U27852 (N_27852,N_21041,N_20846);
nand U27853 (N_27853,N_20956,N_20163);
nor U27854 (N_27854,N_21784,N_24548);
nor U27855 (N_27855,N_24431,N_20315);
nor U27856 (N_27856,N_24651,N_20256);
nor U27857 (N_27857,N_24797,N_21720);
and U27858 (N_27858,N_20447,N_20432);
nor U27859 (N_27859,N_20551,N_22943);
and U27860 (N_27860,N_22953,N_21205);
and U27861 (N_27861,N_21148,N_23684);
nor U27862 (N_27862,N_24362,N_21020);
xor U27863 (N_27863,N_22002,N_24372);
and U27864 (N_27864,N_23816,N_20787);
nand U27865 (N_27865,N_24640,N_21088);
and U27866 (N_27866,N_23908,N_21956);
xor U27867 (N_27867,N_21267,N_21379);
or U27868 (N_27868,N_23416,N_22681);
or U27869 (N_27869,N_23185,N_22581);
nand U27870 (N_27870,N_20988,N_20193);
and U27871 (N_27871,N_21086,N_21893);
xor U27872 (N_27872,N_24115,N_24317);
nor U27873 (N_27873,N_24879,N_21601);
nor U27874 (N_27874,N_20223,N_21113);
and U27875 (N_27875,N_22170,N_24490);
nor U27876 (N_27876,N_22677,N_21139);
nand U27877 (N_27877,N_23676,N_20320);
nor U27878 (N_27878,N_20235,N_22963);
and U27879 (N_27879,N_23586,N_22681);
xor U27880 (N_27880,N_21109,N_22048);
nand U27881 (N_27881,N_23288,N_22689);
or U27882 (N_27882,N_20198,N_23114);
xor U27883 (N_27883,N_20723,N_21397);
or U27884 (N_27884,N_20916,N_21074);
xnor U27885 (N_27885,N_24699,N_23083);
nor U27886 (N_27886,N_24966,N_24207);
and U27887 (N_27887,N_24484,N_22736);
or U27888 (N_27888,N_24203,N_20056);
xor U27889 (N_27889,N_21754,N_24873);
nor U27890 (N_27890,N_22133,N_20475);
xor U27891 (N_27891,N_21237,N_23174);
or U27892 (N_27892,N_20698,N_20925);
nand U27893 (N_27893,N_21930,N_22753);
xor U27894 (N_27894,N_24641,N_21734);
xnor U27895 (N_27895,N_24064,N_21786);
xor U27896 (N_27896,N_23892,N_23177);
xnor U27897 (N_27897,N_20704,N_21081);
nand U27898 (N_27898,N_22359,N_22297);
xor U27899 (N_27899,N_24976,N_20624);
nand U27900 (N_27900,N_20359,N_24672);
xor U27901 (N_27901,N_21912,N_20820);
xor U27902 (N_27902,N_24989,N_23547);
xnor U27903 (N_27903,N_22428,N_23269);
or U27904 (N_27904,N_21749,N_23610);
xnor U27905 (N_27905,N_22770,N_21317);
nand U27906 (N_27906,N_23894,N_23933);
or U27907 (N_27907,N_24999,N_20585);
nand U27908 (N_27908,N_24341,N_24073);
and U27909 (N_27909,N_21604,N_20502);
xnor U27910 (N_27910,N_22752,N_23446);
xnor U27911 (N_27911,N_23656,N_22739);
nand U27912 (N_27912,N_20159,N_24472);
xnor U27913 (N_27913,N_23756,N_23842);
nand U27914 (N_27914,N_22746,N_24424);
xor U27915 (N_27915,N_21763,N_24220);
or U27916 (N_27916,N_23004,N_21187);
xor U27917 (N_27917,N_23097,N_22748);
xnor U27918 (N_27918,N_20529,N_23232);
and U27919 (N_27919,N_21971,N_21932);
nor U27920 (N_27920,N_21369,N_24197);
nor U27921 (N_27921,N_23039,N_21376);
or U27922 (N_27922,N_23778,N_23161);
nand U27923 (N_27923,N_23306,N_24320);
nor U27924 (N_27924,N_23921,N_21503);
xor U27925 (N_27925,N_22816,N_23656);
xor U27926 (N_27926,N_24801,N_22959);
and U27927 (N_27927,N_20269,N_24500);
and U27928 (N_27928,N_23157,N_20688);
and U27929 (N_27929,N_21038,N_24901);
xnor U27930 (N_27930,N_20176,N_22306);
nor U27931 (N_27931,N_22572,N_22021);
nor U27932 (N_27932,N_20907,N_22913);
nor U27933 (N_27933,N_23880,N_22001);
and U27934 (N_27934,N_23084,N_22259);
nor U27935 (N_27935,N_24451,N_23609);
and U27936 (N_27936,N_22816,N_21624);
and U27937 (N_27937,N_24651,N_20822);
nor U27938 (N_27938,N_20701,N_20576);
and U27939 (N_27939,N_20463,N_21978);
and U27940 (N_27940,N_21388,N_24564);
nand U27941 (N_27941,N_21469,N_22745);
and U27942 (N_27942,N_22800,N_23910);
or U27943 (N_27943,N_20069,N_21061);
nor U27944 (N_27944,N_24050,N_21018);
nor U27945 (N_27945,N_21432,N_23823);
nand U27946 (N_27946,N_20597,N_20933);
nand U27947 (N_27947,N_21262,N_21992);
nor U27948 (N_27948,N_24075,N_23571);
nand U27949 (N_27949,N_23195,N_20576);
or U27950 (N_27950,N_21713,N_23328);
or U27951 (N_27951,N_21752,N_21482);
and U27952 (N_27952,N_21359,N_20680);
or U27953 (N_27953,N_21583,N_24560);
xnor U27954 (N_27954,N_20977,N_20325);
nand U27955 (N_27955,N_20236,N_22115);
or U27956 (N_27956,N_22593,N_22040);
nand U27957 (N_27957,N_21905,N_22163);
and U27958 (N_27958,N_24394,N_20237);
nor U27959 (N_27959,N_22017,N_21749);
or U27960 (N_27960,N_23268,N_20598);
or U27961 (N_27961,N_20548,N_20499);
or U27962 (N_27962,N_23806,N_22625);
nand U27963 (N_27963,N_20686,N_22130);
xnor U27964 (N_27964,N_22224,N_20553);
nor U27965 (N_27965,N_21115,N_23401);
and U27966 (N_27966,N_20934,N_20757);
xnor U27967 (N_27967,N_22740,N_20755);
nand U27968 (N_27968,N_23087,N_22334);
and U27969 (N_27969,N_24855,N_24121);
xor U27970 (N_27970,N_24565,N_20089);
nor U27971 (N_27971,N_20589,N_23632);
nor U27972 (N_27972,N_23778,N_20853);
nor U27973 (N_27973,N_24471,N_23026);
nand U27974 (N_27974,N_24110,N_21406);
nand U27975 (N_27975,N_20981,N_24217);
or U27976 (N_27976,N_23852,N_20176);
and U27977 (N_27977,N_22493,N_23398);
and U27978 (N_27978,N_24170,N_20551);
and U27979 (N_27979,N_21809,N_24881);
xnor U27980 (N_27980,N_21538,N_24811);
xnor U27981 (N_27981,N_23814,N_21872);
or U27982 (N_27982,N_22204,N_24415);
nand U27983 (N_27983,N_20544,N_22063);
xnor U27984 (N_27984,N_20549,N_22561);
nand U27985 (N_27985,N_23918,N_23544);
or U27986 (N_27986,N_22304,N_21320);
or U27987 (N_27987,N_24362,N_20274);
or U27988 (N_27988,N_21830,N_21619);
nor U27989 (N_27989,N_21416,N_23132);
nor U27990 (N_27990,N_21689,N_20560);
or U27991 (N_27991,N_23687,N_21046);
nor U27992 (N_27992,N_23971,N_23477);
and U27993 (N_27993,N_24502,N_22309);
xnor U27994 (N_27994,N_24857,N_24650);
nor U27995 (N_27995,N_20027,N_20427);
nor U27996 (N_27996,N_23318,N_23520);
or U27997 (N_27997,N_22485,N_24115);
nor U27998 (N_27998,N_20250,N_21315);
and U27999 (N_27999,N_20921,N_21705);
nand U28000 (N_28000,N_20693,N_24882);
nand U28001 (N_28001,N_23684,N_21555);
or U28002 (N_28002,N_20884,N_21854);
xnor U28003 (N_28003,N_23534,N_21958);
nand U28004 (N_28004,N_24214,N_23401);
or U28005 (N_28005,N_20680,N_24927);
nand U28006 (N_28006,N_21055,N_22555);
nor U28007 (N_28007,N_21225,N_23515);
and U28008 (N_28008,N_24179,N_23713);
nand U28009 (N_28009,N_24081,N_24708);
or U28010 (N_28010,N_24541,N_23085);
or U28011 (N_28011,N_21658,N_24837);
nor U28012 (N_28012,N_22203,N_21292);
and U28013 (N_28013,N_21581,N_21781);
nor U28014 (N_28014,N_23599,N_23535);
xor U28015 (N_28015,N_22947,N_23882);
nand U28016 (N_28016,N_24085,N_22256);
or U28017 (N_28017,N_21439,N_22843);
nor U28018 (N_28018,N_21879,N_20266);
and U28019 (N_28019,N_22771,N_23822);
nor U28020 (N_28020,N_24150,N_21120);
nand U28021 (N_28021,N_23648,N_24329);
xnor U28022 (N_28022,N_24656,N_24727);
or U28023 (N_28023,N_24523,N_21578);
xnor U28024 (N_28024,N_21875,N_21382);
nand U28025 (N_28025,N_23099,N_23133);
or U28026 (N_28026,N_23230,N_23759);
nor U28027 (N_28027,N_20157,N_21184);
nor U28028 (N_28028,N_21318,N_24259);
and U28029 (N_28029,N_21898,N_24292);
or U28030 (N_28030,N_20033,N_20918);
xnor U28031 (N_28031,N_22199,N_23742);
nor U28032 (N_28032,N_20249,N_21575);
xor U28033 (N_28033,N_22494,N_24545);
nor U28034 (N_28034,N_23947,N_24244);
xor U28035 (N_28035,N_20869,N_22317);
nand U28036 (N_28036,N_23233,N_21801);
nor U28037 (N_28037,N_24489,N_24251);
xnor U28038 (N_28038,N_21719,N_24636);
or U28039 (N_28039,N_21477,N_20651);
or U28040 (N_28040,N_22505,N_21631);
and U28041 (N_28041,N_24557,N_24174);
and U28042 (N_28042,N_20069,N_21583);
and U28043 (N_28043,N_22798,N_22693);
nor U28044 (N_28044,N_22549,N_23814);
xor U28045 (N_28045,N_20453,N_21311);
and U28046 (N_28046,N_24732,N_22811);
nor U28047 (N_28047,N_22464,N_23236);
or U28048 (N_28048,N_24407,N_20324);
xor U28049 (N_28049,N_20031,N_23721);
and U28050 (N_28050,N_24612,N_24757);
nor U28051 (N_28051,N_24222,N_23918);
nor U28052 (N_28052,N_24341,N_24590);
xor U28053 (N_28053,N_24793,N_21384);
nand U28054 (N_28054,N_24595,N_23447);
nor U28055 (N_28055,N_23710,N_24423);
xor U28056 (N_28056,N_23186,N_22374);
xor U28057 (N_28057,N_21306,N_21120);
nand U28058 (N_28058,N_23540,N_24775);
or U28059 (N_28059,N_22379,N_23188);
and U28060 (N_28060,N_21586,N_23716);
nand U28061 (N_28061,N_23092,N_23511);
nor U28062 (N_28062,N_23492,N_22696);
xor U28063 (N_28063,N_23768,N_23859);
nor U28064 (N_28064,N_20612,N_20942);
or U28065 (N_28065,N_24332,N_21449);
or U28066 (N_28066,N_22966,N_22500);
or U28067 (N_28067,N_24885,N_21990);
or U28068 (N_28068,N_22069,N_20761);
nor U28069 (N_28069,N_23054,N_22319);
or U28070 (N_28070,N_23904,N_20424);
xnor U28071 (N_28071,N_24202,N_24781);
xnor U28072 (N_28072,N_23964,N_22516);
nor U28073 (N_28073,N_23829,N_22411);
or U28074 (N_28074,N_24679,N_21932);
xor U28075 (N_28075,N_20019,N_22568);
xnor U28076 (N_28076,N_21231,N_23322);
or U28077 (N_28077,N_20125,N_21826);
and U28078 (N_28078,N_24256,N_20497);
nand U28079 (N_28079,N_23216,N_20000);
or U28080 (N_28080,N_20013,N_23242);
or U28081 (N_28081,N_21413,N_23580);
and U28082 (N_28082,N_21684,N_23289);
xor U28083 (N_28083,N_23213,N_22667);
xnor U28084 (N_28084,N_24130,N_21430);
nand U28085 (N_28085,N_20868,N_22593);
nand U28086 (N_28086,N_22142,N_23739);
nand U28087 (N_28087,N_24051,N_22591);
nor U28088 (N_28088,N_24276,N_24308);
xnor U28089 (N_28089,N_21609,N_22325);
xnor U28090 (N_28090,N_20741,N_24673);
xor U28091 (N_28091,N_24899,N_24884);
nor U28092 (N_28092,N_24679,N_24686);
nor U28093 (N_28093,N_21645,N_23056);
or U28094 (N_28094,N_24031,N_24150);
or U28095 (N_28095,N_24956,N_20008);
nand U28096 (N_28096,N_21658,N_22363);
xnor U28097 (N_28097,N_23068,N_21739);
or U28098 (N_28098,N_24427,N_24318);
nand U28099 (N_28099,N_24526,N_20664);
xor U28100 (N_28100,N_22462,N_23632);
or U28101 (N_28101,N_24962,N_21565);
xnor U28102 (N_28102,N_23204,N_23953);
nand U28103 (N_28103,N_23000,N_24602);
nand U28104 (N_28104,N_22075,N_23393);
or U28105 (N_28105,N_21903,N_20440);
or U28106 (N_28106,N_22754,N_23533);
or U28107 (N_28107,N_22638,N_21859);
xnor U28108 (N_28108,N_20979,N_21438);
nand U28109 (N_28109,N_21569,N_24216);
or U28110 (N_28110,N_21244,N_24808);
or U28111 (N_28111,N_24261,N_24938);
xnor U28112 (N_28112,N_20913,N_24677);
and U28113 (N_28113,N_23162,N_22638);
xnor U28114 (N_28114,N_22402,N_24415);
and U28115 (N_28115,N_23528,N_23677);
nand U28116 (N_28116,N_23842,N_21724);
xnor U28117 (N_28117,N_23553,N_21079);
nor U28118 (N_28118,N_23867,N_24649);
or U28119 (N_28119,N_24442,N_23471);
nor U28120 (N_28120,N_21784,N_20294);
or U28121 (N_28121,N_24438,N_23821);
nor U28122 (N_28122,N_21904,N_24884);
nand U28123 (N_28123,N_23414,N_20253);
or U28124 (N_28124,N_23004,N_23510);
nor U28125 (N_28125,N_21661,N_24843);
xor U28126 (N_28126,N_24473,N_20597);
and U28127 (N_28127,N_22156,N_23517);
xnor U28128 (N_28128,N_24787,N_24816);
xor U28129 (N_28129,N_23637,N_24158);
nand U28130 (N_28130,N_22853,N_22078);
nand U28131 (N_28131,N_20007,N_24950);
or U28132 (N_28132,N_21750,N_24321);
nand U28133 (N_28133,N_21416,N_21358);
nor U28134 (N_28134,N_23630,N_21239);
and U28135 (N_28135,N_24504,N_20103);
and U28136 (N_28136,N_20635,N_20240);
and U28137 (N_28137,N_23119,N_21391);
and U28138 (N_28138,N_21638,N_21617);
nand U28139 (N_28139,N_22430,N_20831);
or U28140 (N_28140,N_22046,N_21219);
and U28141 (N_28141,N_24053,N_24261);
nand U28142 (N_28142,N_24742,N_22640);
xor U28143 (N_28143,N_21359,N_23614);
or U28144 (N_28144,N_23584,N_22024);
nand U28145 (N_28145,N_22894,N_20711);
nand U28146 (N_28146,N_21240,N_23430);
nand U28147 (N_28147,N_23805,N_23969);
xor U28148 (N_28148,N_21264,N_21207);
and U28149 (N_28149,N_21459,N_23084);
nand U28150 (N_28150,N_23032,N_20196);
nor U28151 (N_28151,N_23765,N_20794);
and U28152 (N_28152,N_23449,N_20580);
or U28153 (N_28153,N_23997,N_24554);
xnor U28154 (N_28154,N_20186,N_20031);
xor U28155 (N_28155,N_24821,N_20892);
xnor U28156 (N_28156,N_24545,N_23416);
nand U28157 (N_28157,N_23067,N_23586);
or U28158 (N_28158,N_23270,N_20574);
or U28159 (N_28159,N_22204,N_24707);
xnor U28160 (N_28160,N_24474,N_20253);
or U28161 (N_28161,N_21429,N_22289);
nand U28162 (N_28162,N_20985,N_24393);
nand U28163 (N_28163,N_22591,N_23019);
nand U28164 (N_28164,N_20052,N_22861);
or U28165 (N_28165,N_24804,N_20338);
nor U28166 (N_28166,N_21370,N_21398);
nand U28167 (N_28167,N_24645,N_22825);
xor U28168 (N_28168,N_23025,N_20574);
nor U28169 (N_28169,N_23113,N_21441);
xor U28170 (N_28170,N_23094,N_24346);
nand U28171 (N_28171,N_23063,N_24835);
or U28172 (N_28172,N_23670,N_24351);
or U28173 (N_28173,N_22423,N_24333);
xnor U28174 (N_28174,N_23172,N_23008);
and U28175 (N_28175,N_20253,N_22124);
xor U28176 (N_28176,N_23757,N_20149);
or U28177 (N_28177,N_22060,N_23531);
or U28178 (N_28178,N_21349,N_24557);
xnor U28179 (N_28179,N_23615,N_24493);
xnor U28180 (N_28180,N_21423,N_20209);
nand U28181 (N_28181,N_22108,N_20461);
and U28182 (N_28182,N_20195,N_24279);
or U28183 (N_28183,N_20905,N_20270);
or U28184 (N_28184,N_24159,N_24654);
nand U28185 (N_28185,N_21167,N_23203);
or U28186 (N_28186,N_24955,N_21087);
xor U28187 (N_28187,N_23517,N_20401);
nor U28188 (N_28188,N_24935,N_23606);
or U28189 (N_28189,N_21232,N_23237);
nor U28190 (N_28190,N_20878,N_22527);
or U28191 (N_28191,N_21887,N_22340);
or U28192 (N_28192,N_20210,N_22876);
xor U28193 (N_28193,N_21286,N_23250);
and U28194 (N_28194,N_24845,N_23510);
xor U28195 (N_28195,N_22457,N_20852);
nand U28196 (N_28196,N_21747,N_22252);
xnor U28197 (N_28197,N_22085,N_24683);
nor U28198 (N_28198,N_20274,N_20995);
nor U28199 (N_28199,N_23954,N_21301);
xor U28200 (N_28200,N_20504,N_21717);
xnor U28201 (N_28201,N_22181,N_22191);
or U28202 (N_28202,N_23989,N_20941);
and U28203 (N_28203,N_23675,N_21380);
nor U28204 (N_28204,N_22217,N_20424);
nor U28205 (N_28205,N_20379,N_22100);
or U28206 (N_28206,N_24320,N_20771);
xor U28207 (N_28207,N_20613,N_24885);
nand U28208 (N_28208,N_22471,N_21892);
nand U28209 (N_28209,N_24255,N_24891);
and U28210 (N_28210,N_21312,N_24457);
xor U28211 (N_28211,N_20329,N_20902);
nand U28212 (N_28212,N_21471,N_21199);
and U28213 (N_28213,N_21446,N_22174);
nor U28214 (N_28214,N_24455,N_20437);
nor U28215 (N_28215,N_20606,N_20008);
or U28216 (N_28216,N_20936,N_20182);
xor U28217 (N_28217,N_22540,N_22075);
nor U28218 (N_28218,N_23032,N_23021);
or U28219 (N_28219,N_20654,N_21930);
or U28220 (N_28220,N_20162,N_22314);
xnor U28221 (N_28221,N_20635,N_24807);
and U28222 (N_28222,N_24603,N_24982);
nor U28223 (N_28223,N_21001,N_22927);
nor U28224 (N_28224,N_22281,N_20783);
xnor U28225 (N_28225,N_23233,N_23293);
and U28226 (N_28226,N_21132,N_22307);
xor U28227 (N_28227,N_23255,N_22213);
or U28228 (N_28228,N_23183,N_22815);
and U28229 (N_28229,N_20804,N_21414);
nor U28230 (N_28230,N_22130,N_23899);
and U28231 (N_28231,N_20164,N_23802);
xnor U28232 (N_28232,N_23270,N_21265);
or U28233 (N_28233,N_24561,N_21741);
nand U28234 (N_28234,N_21564,N_21825);
xnor U28235 (N_28235,N_21169,N_20512);
xor U28236 (N_28236,N_21186,N_23092);
nor U28237 (N_28237,N_21014,N_23868);
xor U28238 (N_28238,N_23171,N_24806);
or U28239 (N_28239,N_23124,N_24914);
or U28240 (N_28240,N_24527,N_23492);
or U28241 (N_28241,N_22406,N_24020);
and U28242 (N_28242,N_20015,N_23233);
nor U28243 (N_28243,N_21910,N_22329);
nor U28244 (N_28244,N_21950,N_24257);
nor U28245 (N_28245,N_23604,N_24826);
and U28246 (N_28246,N_22394,N_22418);
and U28247 (N_28247,N_20888,N_21814);
or U28248 (N_28248,N_21629,N_21893);
and U28249 (N_28249,N_20998,N_20421);
nand U28250 (N_28250,N_24685,N_21922);
or U28251 (N_28251,N_20323,N_23022);
and U28252 (N_28252,N_21429,N_24539);
and U28253 (N_28253,N_23339,N_20131);
nand U28254 (N_28254,N_23562,N_21093);
nand U28255 (N_28255,N_24832,N_24196);
xnor U28256 (N_28256,N_24044,N_24040);
or U28257 (N_28257,N_24404,N_23264);
and U28258 (N_28258,N_21999,N_21341);
nand U28259 (N_28259,N_20372,N_23253);
xnor U28260 (N_28260,N_21619,N_20662);
nor U28261 (N_28261,N_24641,N_21846);
nand U28262 (N_28262,N_22723,N_20211);
xor U28263 (N_28263,N_22820,N_20972);
nand U28264 (N_28264,N_22595,N_22838);
nand U28265 (N_28265,N_22221,N_22716);
nor U28266 (N_28266,N_24006,N_23362);
and U28267 (N_28267,N_24683,N_21753);
or U28268 (N_28268,N_22221,N_23034);
and U28269 (N_28269,N_24339,N_24096);
nor U28270 (N_28270,N_22906,N_23311);
nand U28271 (N_28271,N_24634,N_21417);
or U28272 (N_28272,N_23136,N_20297);
nor U28273 (N_28273,N_21544,N_20143);
nor U28274 (N_28274,N_22882,N_23841);
and U28275 (N_28275,N_20638,N_20676);
nand U28276 (N_28276,N_24794,N_23084);
nand U28277 (N_28277,N_23846,N_22922);
xor U28278 (N_28278,N_22268,N_23508);
nand U28279 (N_28279,N_21144,N_20532);
nand U28280 (N_28280,N_24451,N_20031);
or U28281 (N_28281,N_21616,N_20561);
nor U28282 (N_28282,N_24624,N_23706);
nor U28283 (N_28283,N_21009,N_23261);
xnor U28284 (N_28284,N_20720,N_20837);
nand U28285 (N_28285,N_20052,N_21620);
nor U28286 (N_28286,N_20813,N_23018);
and U28287 (N_28287,N_24893,N_20018);
or U28288 (N_28288,N_24257,N_21131);
nor U28289 (N_28289,N_22103,N_20964);
or U28290 (N_28290,N_21092,N_21471);
and U28291 (N_28291,N_20938,N_24408);
xor U28292 (N_28292,N_24581,N_21799);
nand U28293 (N_28293,N_22255,N_21628);
xnor U28294 (N_28294,N_22160,N_21812);
and U28295 (N_28295,N_22787,N_20354);
and U28296 (N_28296,N_22272,N_24982);
nand U28297 (N_28297,N_24312,N_22810);
nor U28298 (N_28298,N_24158,N_21939);
or U28299 (N_28299,N_24672,N_24978);
nand U28300 (N_28300,N_20906,N_20067);
or U28301 (N_28301,N_21474,N_20665);
xor U28302 (N_28302,N_23541,N_21815);
nor U28303 (N_28303,N_20950,N_22705);
and U28304 (N_28304,N_24921,N_22515);
xor U28305 (N_28305,N_21659,N_22832);
xnor U28306 (N_28306,N_20553,N_23116);
nand U28307 (N_28307,N_24855,N_20787);
or U28308 (N_28308,N_21398,N_23235);
nor U28309 (N_28309,N_22877,N_22092);
and U28310 (N_28310,N_22295,N_23890);
and U28311 (N_28311,N_23299,N_24258);
nand U28312 (N_28312,N_20333,N_21366);
nand U28313 (N_28313,N_21259,N_23417);
or U28314 (N_28314,N_23378,N_22942);
nand U28315 (N_28315,N_24938,N_23585);
and U28316 (N_28316,N_22744,N_23795);
and U28317 (N_28317,N_24600,N_21034);
or U28318 (N_28318,N_24616,N_21734);
nor U28319 (N_28319,N_24575,N_20515);
xnor U28320 (N_28320,N_23545,N_22903);
and U28321 (N_28321,N_24037,N_24927);
nor U28322 (N_28322,N_23715,N_24856);
nor U28323 (N_28323,N_23580,N_22532);
xor U28324 (N_28324,N_24577,N_21635);
nor U28325 (N_28325,N_20544,N_20676);
or U28326 (N_28326,N_24958,N_20286);
nand U28327 (N_28327,N_23519,N_20816);
and U28328 (N_28328,N_23070,N_24648);
or U28329 (N_28329,N_20323,N_20070);
and U28330 (N_28330,N_24765,N_20646);
or U28331 (N_28331,N_20479,N_22888);
nand U28332 (N_28332,N_24631,N_20641);
or U28333 (N_28333,N_20470,N_23209);
xnor U28334 (N_28334,N_20347,N_20810);
and U28335 (N_28335,N_22135,N_21876);
nor U28336 (N_28336,N_20818,N_24887);
xor U28337 (N_28337,N_23846,N_23794);
xor U28338 (N_28338,N_23432,N_23823);
xnor U28339 (N_28339,N_21872,N_20161);
or U28340 (N_28340,N_21443,N_21455);
nor U28341 (N_28341,N_20654,N_22412);
nand U28342 (N_28342,N_20971,N_20356);
nand U28343 (N_28343,N_23122,N_21679);
nand U28344 (N_28344,N_21201,N_21903);
or U28345 (N_28345,N_21295,N_20745);
nor U28346 (N_28346,N_23169,N_22945);
and U28347 (N_28347,N_22202,N_20876);
nand U28348 (N_28348,N_23631,N_24047);
nor U28349 (N_28349,N_21290,N_24699);
nand U28350 (N_28350,N_23764,N_20796);
and U28351 (N_28351,N_22390,N_22185);
nor U28352 (N_28352,N_22266,N_24036);
and U28353 (N_28353,N_21678,N_21532);
nor U28354 (N_28354,N_23322,N_21693);
and U28355 (N_28355,N_20289,N_22834);
xnor U28356 (N_28356,N_20632,N_23595);
xor U28357 (N_28357,N_24620,N_22844);
xor U28358 (N_28358,N_24525,N_22962);
or U28359 (N_28359,N_21264,N_21800);
xor U28360 (N_28360,N_23279,N_23542);
or U28361 (N_28361,N_22644,N_22336);
and U28362 (N_28362,N_23704,N_20338);
xor U28363 (N_28363,N_20242,N_20286);
nor U28364 (N_28364,N_24961,N_23340);
nor U28365 (N_28365,N_21360,N_23692);
and U28366 (N_28366,N_22379,N_20690);
and U28367 (N_28367,N_21498,N_21290);
nand U28368 (N_28368,N_23697,N_23525);
nand U28369 (N_28369,N_24114,N_20269);
xor U28370 (N_28370,N_24135,N_20803);
nand U28371 (N_28371,N_20557,N_21598);
and U28372 (N_28372,N_23420,N_23711);
xnor U28373 (N_28373,N_21789,N_23610);
nand U28374 (N_28374,N_23052,N_20408);
xor U28375 (N_28375,N_24128,N_20635);
xnor U28376 (N_28376,N_24526,N_22817);
or U28377 (N_28377,N_21104,N_23066);
nor U28378 (N_28378,N_24201,N_24576);
nand U28379 (N_28379,N_20030,N_20578);
nand U28380 (N_28380,N_20421,N_22535);
xor U28381 (N_28381,N_22421,N_23784);
or U28382 (N_28382,N_24844,N_21391);
nor U28383 (N_28383,N_21417,N_24519);
nor U28384 (N_28384,N_21223,N_22369);
and U28385 (N_28385,N_24677,N_21105);
or U28386 (N_28386,N_23276,N_21693);
or U28387 (N_28387,N_21456,N_24837);
or U28388 (N_28388,N_23206,N_21369);
and U28389 (N_28389,N_23481,N_21191);
or U28390 (N_28390,N_23059,N_21936);
xnor U28391 (N_28391,N_23499,N_24960);
nor U28392 (N_28392,N_21154,N_23341);
nor U28393 (N_28393,N_20819,N_24179);
nand U28394 (N_28394,N_23429,N_21400);
or U28395 (N_28395,N_22897,N_22474);
nor U28396 (N_28396,N_23619,N_22393);
nand U28397 (N_28397,N_20061,N_22842);
nand U28398 (N_28398,N_22774,N_23812);
or U28399 (N_28399,N_22669,N_20902);
nor U28400 (N_28400,N_22478,N_22002);
and U28401 (N_28401,N_22179,N_23810);
nand U28402 (N_28402,N_22153,N_24200);
nor U28403 (N_28403,N_23858,N_22591);
or U28404 (N_28404,N_20921,N_21092);
nand U28405 (N_28405,N_22367,N_21605);
xnor U28406 (N_28406,N_24909,N_24243);
or U28407 (N_28407,N_23544,N_21709);
or U28408 (N_28408,N_21751,N_24536);
and U28409 (N_28409,N_23343,N_23053);
nor U28410 (N_28410,N_21972,N_20784);
nor U28411 (N_28411,N_21016,N_23243);
nor U28412 (N_28412,N_22458,N_21478);
or U28413 (N_28413,N_24229,N_23263);
or U28414 (N_28414,N_24922,N_22602);
and U28415 (N_28415,N_24418,N_21392);
xor U28416 (N_28416,N_21909,N_23593);
nand U28417 (N_28417,N_24502,N_21712);
and U28418 (N_28418,N_23434,N_22501);
and U28419 (N_28419,N_21622,N_22040);
and U28420 (N_28420,N_21203,N_21814);
nor U28421 (N_28421,N_20514,N_20310);
and U28422 (N_28422,N_20235,N_22184);
nor U28423 (N_28423,N_24840,N_23691);
nand U28424 (N_28424,N_24743,N_24326);
xnor U28425 (N_28425,N_24775,N_24475);
or U28426 (N_28426,N_21776,N_23594);
nand U28427 (N_28427,N_23656,N_22107);
xnor U28428 (N_28428,N_24963,N_21699);
and U28429 (N_28429,N_23406,N_20694);
xor U28430 (N_28430,N_24694,N_21123);
and U28431 (N_28431,N_21858,N_24940);
and U28432 (N_28432,N_24170,N_23457);
nor U28433 (N_28433,N_24096,N_20155);
or U28434 (N_28434,N_23714,N_21631);
xnor U28435 (N_28435,N_20209,N_23659);
and U28436 (N_28436,N_22389,N_24359);
xnor U28437 (N_28437,N_23758,N_22691);
xnor U28438 (N_28438,N_24596,N_22159);
or U28439 (N_28439,N_20856,N_20351);
nor U28440 (N_28440,N_23820,N_23810);
and U28441 (N_28441,N_20955,N_21302);
nand U28442 (N_28442,N_24401,N_21100);
xor U28443 (N_28443,N_21630,N_22599);
xor U28444 (N_28444,N_23698,N_23794);
and U28445 (N_28445,N_20005,N_21287);
nand U28446 (N_28446,N_23045,N_20224);
nand U28447 (N_28447,N_22998,N_23390);
nand U28448 (N_28448,N_21763,N_23012);
or U28449 (N_28449,N_23179,N_23424);
and U28450 (N_28450,N_20609,N_21867);
or U28451 (N_28451,N_23810,N_24621);
nor U28452 (N_28452,N_21259,N_20552);
xnor U28453 (N_28453,N_24027,N_20001);
and U28454 (N_28454,N_23618,N_24020);
or U28455 (N_28455,N_24074,N_24233);
or U28456 (N_28456,N_20104,N_20140);
xnor U28457 (N_28457,N_24937,N_20361);
xor U28458 (N_28458,N_24064,N_21151);
or U28459 (N_28459,N_20166,N_20585);
nor U28460 (N_28460,N_20551,N_20073);
and U28461 (N_28461,N_21598,N_24062);
or U28462 (N_28462,N_22134,N_24884);
or U28463 (N_28463,N_23071,N_24422);
or U28464 (N_28464,N_22268,N_23945);
xnor U28465 (N_28465,N_23037,N_22760);
xor U28466 (N_28466,N_21754,N_23923);
xnor U28467 (N_28467,N_20121,N_21714);
xnor U28468 (N_28468,N_24960,N_24137);
nand U28469 (N_28469,N_21739,N_20174);
or U28470 (N_28470,N_24218,N_20902);
xnor U28471 (N_28471,N_23300,N_20902);
xor U28472 (N_28472,N_23523,N_21671);
or U28473 (N_28473,N_24261,N_21712);
and U28474 (N_28474,N_23943,N_24923);
nor U28475 (N_28475,N_24240,N_24342);
xnor U28476 (N_28476,N_24076,N_22006);
or U28477 (N_28477,N_20877,N_22677);
xor U28478 (N_28478,N_22589,N_24650);
xnor U28479 (N_28479,N_20925,N_22917);
and U28480 (N_28480,N_20486,N_21203);
nand U28481 (N_28481,N_24012,N_23399);
xnor U28482 (N_28482,N_24997,N_21115);
or U28483 (N_28483,N_20257,N_22557);
nand U28484 (N_28484,N_23084,N_24111);
nand U28485 (N_28485,N_22254,N_23002);
and U28486 (N_28486,N_24643,N_22670);
nand U28487 (N_28487,N_23207,N_24857);
xor U28488 (N_28488,N_21341,N_23648);
or U28489 (N_28489,N_21622,N_21012);
xnor U28490 (N_28490,N_21085,N_21803);
xnor U28491 (N_28491,N_24509,N_23589);
xor U28492 (N_28492,N_24156,N_22982);
and U28493 (N_28493,N_21017,N_22338);
xnor U28494 (N_28494,N_23004,N_21534);
and U28495 (N_28495,N_22027,N_20021);
and U28496 (N_28496,N_23217,N_23975);
xnor U28497 (N_28497,N_23940,N_24182);
and U28498 (N_28498,N_24947,N_22430);
nand U28499 (N_28499,N_24748,N_20349);
or U28500 (N_28500,N_23670,N_23086);
nor U28501 (N_28501,N_23004,N_22306);
xnor U28502 (N_28502,N_21397,N_23596);
or U28503 (N_28503,N_21612,N_20857);
and U28504 (N_28504,N_23708,N_20260);
and U28505 (N_28505,N_21405,N_23575);
or U28506 (N_28506,N_24210,N_20010);
and U28507 (N_28507,N_22367,N_23623);
nand U28508 (N_28508,N_23598,N_21029);
xnor U28509 (N_28509,N_21419,N_22320);
nor U28510 (N_28510,N_20025,N_22180);
nor U28511 (N_28511,N_24133,N_23608);
or U28512 (N_28512,N_22489,N_21560);
xor U28513 (N_28513,N_22289,N_20196);
or U28514 (N_28514,N_24884,N_24794);
xor U28515 (N_28515,N_21625,N_20939);
nand U28516 (N_28516,N_24269,N_24853);
nand U28517 (N_28517,N_24918,N_21126);
and U28518 (N_28518,N_20977,N_21307);
xor U28519 (N_28519,N_21716,N_20296);
nand U28520 (N_28520,N_20976,N_23054);
and U28521 (N_28521,N_22293,N_23077);
and U28522 (N_28522,N_20202,N_23981);
or U28523 (N_28523,N_24624,N_22112);
nor U28524 (N_28524,N_23829,N_24560);
nor U28525 (N_28525,N_22415,N_21597);
and U28526 (N_28526,N_24871,N_24252);
and U28527 (N_28527,N_21346,N_23941);
nor U28528 (N_28528,N_22555,N_22983);
xnor U28529 (N_28529,N_24417,N_24517);
xor U28530 (N_28530,N_24078,N_22950);
nand U28531 (N_28531,N_23253,N_24399);
nor U28532 (N_28532,N_22526,N_23033);
nor U28533 (N_28533,N_23495,N_20074);
nand U28534 (N_28534,N_20366,N_24122);
and U28535 (N_28535,N_21968,N_24659);
xnor U28536 (N_28536,N_21652,N_21183);
or U28537 (N_28537,N_24502,N_24967);
nand U28538 (N_28538,N_24894,N_20384);
xnor U28539 (N_28539,N_21716,N_20271);
nand U28540 (N_28540,N_20746,N_23791);
xor U28541 (N_28541,N_22095,N_20023);
nor U28542 (N_28542,N_23336,N_22099);
or U28543 (N_28543,N_22497,N_21957);
xnor U28544 (N_28544,N_20432,N_23144);
xnor U28545 (N_28545,N_23185,N_22986);
nor U28546 (N_28546,N_21252,N_23255);
or U28547 (N_28547,N_24038,N_21007);
xor U28548 (N_28548,N_24965,N_20786);
xor U28549 (N_28549,N_20180,N_23998);
or U28550 (N_28550,N_22990,N_24661);
nor U28551 (N_28551,N_21304,N_20948);
nor U28552 (N_28552,N_22511,N_23940);
xor U28553 (N_28553,N_23056,N_24077);
xnor U28554 (N_28554,N_23264,N_24174);
and U28555 (N_28555,N_24042,N_21388);
and U28556 (N_28556,N_24927,N_23853);
and U28557 (N_28557,N_23774,N_22672);
or U28558 (N_28558,N_23190,N_21532);
and U28559 (N_28559,N_24014,N_21900);
xnor U28560 (N_28560,N_22241,N_24140);
xnor U28561 (N_28561,N_20958,N_23854);
or U28562 (N_28562,N_24948,N_22632);
nor U28563 (N_28563,N_21719,N_23325);
xnor U28564 (N_28564,N_21624,N_20662);
nor U28565 (N_28565,N_20508,N_22346);
xor U28566 (N_28566,N_24440,N_22098);
or U28567 (N_28567,N_20874,N_20469);
and U28568 (N_28568,N_20879,N_23899);
nor U28569 (N_28569,N_24847,N_22956);
or U28570 (N_28570,N_24796,N_22299);
or U28571 (N_28571,N_21956,N_20827);
or U28572 (N_28572,N_23666,N_21368);
or U28573 (N_28573,N_21992,N_21604);
nor U28574 (N_28574,N_23795,N_22073);
nand U28575 (N_28575,N_24778,N_24119);
nand U28576 (N_28576,N_23437,N_21237);
xnor U28577 (N_28577,N_21393,N_21998);
xnor U28578 (N_28578,N_20572,N_24443);
xnor U28579 (N_28579,N_21638,N_20664);
xnor U28580 (N_28580,N_21566,N_20089);
nor U28581 (N_28581,N_21254,N_24012);
and U28582 (N_28582,N_21186,N_24667);
xnor U28583 (N_28583,N_23064,N_22133);
xnor U28584 (N_28584,N_23865,N_22229);
and U28585 (N_28585,N_22592,N_22488);
nand U28586 (N_28586,N_23080,N_20882);
xor U28587 (N_28587,N_22459,N_23268);
or U28588 (N_28588,N_22164,N_23861);
xor U28589 (N_28589,N_23926,N_20807);
or U28590 (N_28590,N_22671,N_21115);
or U28591 (N_28591,N_20520,N_23916);
and U28592 (N_28592,N_24669,N_23252);
and U28593 (N_28593,N_24580,N_20354);
nand U28594 (N_28594,N_22895,N_23925);
or U28595 (N_28595,N_21868,N_24777);
nor U28596 (N_28596,N_20286,N_24892);
xnor U28597 (N_28597,N_24968,N_24463);
or U28598 (N_28598,N_22337,N_21809);
nor U28599 (N_28599,N_22492,N_23502);
xor U28600 (N_28600,N_22831,N_21568);
xnor U28601 (N_28601,N_20374,N_24414);
or U28602 (N_28602,N_23060,N_24333);
xnor U28603 (N_28603,N_22170,N_20039);
or U28604 (N_28604,N_22778,N_23588);
and U28605 (N_28605,N_22492,N_23016);
nor U28606 (N_28606,N_21684,N_24026);
xor U28607 (N_28607,N_21536,N_24120);
or U28608 (N_28608,N_21625,N_21835);
and U28609 (N_28609,N_20259,N_24311);
or U28610 (N_28610,N_22033,N_22796);
nor U28611 (N_28611,N_22136,N_22507);
nor U28612 (N_28612,N_20038,N_22016);
and U28613 (N_28613,N_22221,N_21950);
xor U28614 (N_28614,N_23782,N_20605);
nand U28615 (N_28615,N_20675,N_21991);
and U28616 (N_28616,N_21792,N_24746);
or U28617 (N_28617,N_24954,N_20086);
xor U28618 (N_28618,N_23145,N_24724);
nor U28619 (N_28619,N_21357,N_22769);
and U28620 (N_28620,N_21027,N_21915);
or U28621 (N_28621,N_22497,N_23507);
and U28622 (N_28622,N_21426,N_21032);
or U28623 (N_28623,N_21368,N_24213);
and U28624 (N_28624,N_20219,N_23858);
and U28625 (N_28625,N_20791,N_24895);
nor U28626 (N_28626,N_20623,N_20470);
and U28627 (N_28627,N_23369,N_24337);
nor U28628 (N_28628,N_20789,N_20592);
or U28629 (N_28629,N_20638,N_21504);
nand U28630 (N_28630,N_23730,N_21726);
or U28631 (N_28631,N_21489,N_21896);
nand U28632 (N_28632,N_22011,N_22640);
nor U28633 (N_28633,N_24499,N_23148);
nand U28634 (N_28634,N_22426,N_22787);
nand U28635 (N_28635,N_22942,N_23839);
nor U28636 (N_28636,N_20129,N_21506);
xnor U28637 (N_28637,N_24385,N_20000);
and U28638 (N_28638,N_20099,N_24919);
nand U28639 (N_28639,N_22616,N_23784);
xnor U28640 (N_28640,N_23745,N_23139);
xnor U28641 (N_28641,N_23393,N_24785);
or U28642 (N_28642,N_21021,N_23557);
or U28643 (N_28643,N_22921,N_23571);
or U28644 (N_28644,N_20355,N_21543);
xor U28645 (N_28645,N_23119,N_24195);
xnor U28646 (N_28646,N_20710,N_20189);
or U28647 (N_28647,N_23278,N_21060);
and U28648 (N_28648,N_20742,N_20659);
or U28649 (N_28649,N_20952,N_23430);
and U28650 (N_28650,N_24468,N_21135);
or U28651 (N_28651,N_24676,N_22290);
or U28652 (N_28652,N_21034,N_24615);
nand U28653 (N_28653,N_22484,N_23320);
nor U28654 (N_28654,N_21677,N_21589);
nand U28655 (N_28655,N_20222,N_21317);
nand U28656 (N_28656,N_21666,N_20810);
xnor U28657 (N_28657,N_20091,N_20098);
nand U28658 (N_28658,N_24646,N_21921);
or U28659 (N_28659,N_24516,N_22405);
or U28660 (N_28660,N_22870,N_22834);
xor U28661 (N_28661,N_22957,N_22877);
nor U28662 (N_28662,N_20828,N_22047);
and U28663 (N_28663,N_20528,N_20853);
and U28664 (N_28664,N_21339,N_22329);
and U28665 (N_28665,N_20289,N_24510);
and U28666 (N_28666,N_24909,N_22076);
or U28667 (N_28667,N_24512,N_21124);
nor U28668 (N_28668,N_21936,N_23638);
and U28669 (N_28669,N_23594,N_20403);
and U28670 (N_28670,N_20689,N_23167);
or U28671 (N_28671,N_24106,N_21194);
nor U28672 (N_28672,N_21809,N_24922);
xnor U28673 (N_28673,N_22359,N_21399);
or U28674 (N_28674,N_21186,N_21388);
xor U28675 (N_28675,N_23185,N_21201);
nand U28676 (N_28676,N_24110,N_22619);
and U28677 (N_28677,N_22232,N_21974);
xor U28678 (N_28678,N_22734,N_22597);
nand U28679 (N_28679,N_22417,N_20262);
nor U28680 (N_28680,N_24123,N_24161);
and U28681 (N_28681,N_20874,N_21910);
and U28682 (N_28682,N_22018,N_22055);
and U28683 (N_28683,N_20588,N_20515);
xnor U28684 (N_28684,N_22006,N_22254);
nor U28685 (N_28685,N_23314,N_22248);
nor U28686 (N_28686,N_22580,N_20611);
and U28687 (N_28687,N_23568,N_21057);
and U28688 (N_28688,N_24420,N_22968);
xor U28689 (N_28689,N_22499,N_24281);
nand U28690 (N_28690,N_23363,N_24731);
and U28691 (N_28691,N_20547,N_23486);
or U28692 (N_28692,N_22397,N_24083);
nor U28693 (N_28693,N_20115,N_24741);
nor U28694 (N_28694,N_24691,N_23338);
nor U28695 (N_28695,N_20595,N_24068);
xor U28696 (N_28696,N_24233,N_24217);
nand U28697 (N_28697,N_24497,N_24631);
nand U28698 (N_28698,N_20226,N_22990);
and U28699 (N_28699,N_24670,N_24612);
nand U28700 (N_28700,N_23430,N_22653);
xnor U28701 (N_28701,N_24567,N_23149);
nand U28702 (N_28702,N_21183,N_21522);
or U28703 (N_28703,N_24957,N_24802);
xor U28704 (N_28704,N_20240,N_24857);
xor U28705 (N_28705,N_21010,N_24604);
nand U28706 (N_28706,N_20287,N_23444);
or U28707 (N_28707,N_23731,N_23904);
xor U28708 (N_28708,N_22222,N_23427);
xnor U28709 (N_28709,N_21093,N_20551);
nor U28710 (N_28710,N_23347,N_24291);
xnor U28711 (N_28711,N_22166,N_22493);
and U28712 (N_28712,N_24477,N_22283);
nor U28713 (N_28713,N_24883,N_22067);
xnor U28714 (N_28714,N_24526,N_23245);
nor U28715 (N_28715,N_23385,N_22032);
nor U28716 (N_28716,N_22894,N_23272);
xnor U28717 (N_28717,N_21755,N_21054);
nand U28718 (N_28718,N_22641,N_21492);
nand U28719 (N_28719,N_20899,N_21149);
or U28720 (N_28720,N_22484,N_23722);
or U28721 (N_28721,N_23192,N_24380);
and U28722 (N_28722,N_22706,N_24974);
nand U28723 (N_28723,N_22467,N_23813);
nand U28724 (N_28724,N_24268,N_20126);
and U28725 (N_28725,N_21973,N_24924);
and U28726 (N_28726,N_21541,N_21003);
and U28727 (N_28727,N_23738,N_22864);
xor U28728 (N_28728,N_20755,N_24550);
xor U28729 (N_28729,N_24504,N_24783);
nor U28730 (N_28730,N_23312,N_24988);
or U28731 (N_28731,N_20270,N_22570);
or U28732 (N_28732,N_22428,N_21548);
xnor U28733 (N_28733,N_21748,N_24201);
and U28734 (N_28734,N_20668,N_22587);
nor U28735 (N_28735,N_24087,N_23419);
nor U28736 (N_28736,N_24940,N_23294);
or U28737 (N_28737,N_23071,N_22646);
and U28738 (N_28738,N_20845,N_23026);
and U28739 (N_28739,N_23414,N_24192);
or U28740 (N_28740,N_21765,N_22497);
and U28741 (N_28741,N_23526,N_23408);
xor U28742 (N_28742,N_24769,N_22510);
xor U28743 (N_28743,N_20604,N_20678);
nor U28744 (N_28744,N_21407,N_21721);
and U28745 (N_28745,N_20363,N_21461);
xor U28746 (N_28746,N_24061,N_20997);
and U28747 (N_28747,N_20805,N_21383);
or U28748 (N_28748,N_24480,N_22297);
nand U28749 (N_28749,N_23193,N_24978);
nand U28750 (N_28750,N_23116,N_21640);
and U28751 (N_28751,N_23484,N_22884);
nand U28752 (N_28752,N_20012,N_22640);
nor U28753 (N_28753,N_24871,N_21199);
nor U28754 (N_28754,N_21483,N_20264);
xor U28755 (N_28755,N_24931,N_22505);
xnor U28756 (N_28756,N_22940,N_20811);
or U28757 (N_28757,N_24639,N_23020);
nand U28758 (N_28758,N_23898,N_24377);
nor U28759 (N_28759,N_24660,N_21210);
xor U28760 (N_28760,N_20471,N_22441);
nor U28761 (N_28761,N_20436,N_20026);
and U28762 (N_28762,N_20782,N_23499);
nand U28763 (N_28763,N_24484,N_23309);
xnor U28764 (N_28764,N_20992,N_21866);
nand U28765 (N_28765,N_20452,N_23066);
xor U28766 (N_28766,N_22412,N_20162);
nand U28767 (N_28767,N_21026,N_22710);
nand U28768 (N_28768,N_23790,N_21089);
nand U28769 (N_28769,N_24537,N_23721);
or U28770 (N_28770,N_21436,N_24524);
nand U28771 (N_28771,N_21166,N_23103);
xnor U28772 (N_28772,N_24185,N_20940);
nand U28773 (N_28773,N_24875,N_20182);
or U28774 (N_28774,N_21773,N_22736);
nor U28775 (N_28775,N_23785,N_21595);
and U28776 (N_28776,N_24018,N_24229);
nor U28777 (N_28777,N_20929,N_20091);
nor U28778 (N_28778,N_23083,N_24583);
xor U28779 (N_28779,N_21459,N_22629);
nor U28780 (N_28780,N_23260,N_23315);
or U28781 (N_28781,N_21992,N_24282);
xnor U28782 (N_28782,N_21701,N_21323);
or U28783 (N_28783,N_22703,N_22335);
and U28784 (N_28784,N_23005,N_24223);
or U28785 (N_28785,N_22376,N_20288);
or U28786 (N_28786,N_21754,N_21746);
nand U28787 (N_28787,N_24677,N_22164);
and U28788 (N_28788,N_21823,N_22261);
nand U28789 (N_28789,N_20891,N_20099);
and U28790 (N_28790,N_20499,N_20059);
nor U28791 (N_28791,N_24051,N_23359);
nand U28792 (N_28792,N_21582,N_22628);
and U28793 (N_28793,N_20959,N_22067);
or U28794 (N_28794,N_23077,N_22791);
nor U28795 (N_28795,N_22043,N_23215);
and U28796 (N_28796,N_21454,N_20844);
xnor U28797 (N_28797,N_24619,N_24139);
and U28798 (N_28798,N_21580,N_22728);
nor U28799 (N_28799,N_21853,N_24720);
xor U28800 (N_28800,N_24897,N_24973);
nor U28801 (N_28801,N_21646,N_22886);
or U28802 (N_28802,N_24218,N_24457);
xnor U28803 (N_28803,N_22206,N_20454);
nor U28804 (N_28804,N_20616,N_22009);
or U28805 (N_28805,N_23382,N_24127);
and U28806 (N_28806,N_21753,N_24733);
nor U28807 (N_28807,N_21716,N_24928);
or U28808 (N_28808,N_21187,N_23697);
and U28809 (N_28809,N_21653,N_21146);
nor U28810 (N_28810,N_23415,N_22977);
xnor U28811 (N_28811,N_20431,N_21859);
and U28812 (N_28812,N_24769,N_21454);
or U28813 (N_28813,N_22758,N_23851);
and U28814 (N_28814,N_20565,N_20300);
nand U28815 (N_28815,N_21863,N_23933);
xor U28816 (N_28816,N_24660,N_21216);
nor U28817 (N_28817,N_23478,N_22557);
xor U28818 (N_28818,N_21489,N_23349);
nor U28819 (N_28819,N_22094,N_21093);
xnor U28820 (N_28820,N_20757,N_24353);
xor U28821 (N_28821,N_23822,N_22990);
nor U28822 (N_28822,N_21314,N_21398);
and U28823 (N_28823,N_20730,N_24474);
or U28824 (N_28824,N_22283,N_20340);
or U28825 (N_28825,N_21114,N_21630);
nand U28826 (N_28826,N_20944,N_24835);
or U28827 (N_28827,N_22412,N_21121);
and U28828 (N_28828,N_20273,N_20190);
nand U28829 (N_28829,N_21299,N_21508);
xnor U28830 (N_28830,N_22761,N_23293);
and U28831 (N_28831,N_22230,N_24366);
and U28832 (N_28832,N_24825,N_20307);
nor U28833 (N_28833,N_22045,N_24931);
xnor U28834 (N_28834,N_20464,N_20787);
and U28835 (N_28835,N_24631,N_21396);
and U28836 (N_28836,N_20244,N_21137);
and U28837 (N_28837,N_24818,N_20822);
and U28838 (N_28838,N_23168,N_23746);
xor U28839 (N_28839,N_24661,N_20136);
or U28840 (N_28840,N_21529,N_22285);
nand U28841 (N_28841,N_21209,N_22835);
and U28842 (N_28842,N_23247,N_23964);
xnor U28843 (N_28843,N_24081,N_21700);
nand U28844 (N_28844,N_20738,N_22601);
nor U28845 (N_28845,N_21295,N_23355);
or U28846 (N_28846,N_24835,N_22420);
nor U28847 (N_28847,N_21491,N_22853);
xnor U28848 (N_28848,N_20358,N_23619);
nor U28849 (N_28849,N_23443,N_22969);
nand U28850 (N_28850,N_21722,N_22287);
or U28851 (N_28851,N_22022,N_20408);
nand U28852 (N_28852,N_23072,N_21908);
nand U28853 (N_28853,N_24371,N_24478);
or U28854 (N_28854,N_22368,N_20373);
xor U28855 (N_28855,N_23370,N_20589);
or U28856 (N_28856,N_21981,N_23677);
xor U28857 (N_28857,N_22513,N_21759);
nand U28858 (N_28858,N_24419,N_20267);
xor U28859 (N_28859,N_22016,N_20155);
and U28860 (N_28860,N_20348,N_23977);
or U28861 (N_28861,N_21638,N_20893);
nand U28862 (N_28862,N_20137,N_23601);
xnor U28863 (N_28863,N_21115,N_22322);
or U28864 (N_28864,N_20266,N_21898);
xnor U28865 (N_28865,N_21667,N_22434);
xor U28866 (N_28866,N_23381,N_20261);
xnor U28867 (N_28867,N_20030,N_23509);
xor U28868 (N_28868,N_21220,N_21239);
xor U28869 (N_28869,N_20344,N_22978);
xnor U28870 (N_28870,N_24149,N_23519);
xnor U28871 (N_28871,N_22530,N_20342);
or U28872 (N_28872,N_22987,N_20119);
and U28873 (N_28873,N_23691,N_23830);
and U28874 (N_28874,N_23201,N_22599);
and U28875 (N_28875,N_24654,N_22787);
or U28876 (N_28876,N_23365,N_23997);
nor U28877 (N_28877,N_20057,N_24224);
nor U28878 (N_28878,N_23669,N_23945);
and U28879 (N_28879,N_21040,N_23336);
nor U28880 (N_28880,N_22216,N_21523);
or U28881 (N_28881,N_23386,N_24354);
or U28882 (N_28882,N_21302,N_20314);
xnor U28883 (N_28883,N_21430,N_21982);
nor U28884 (N_28884,N_22545,N_23817);
nor U28885 (N_28885,N_24769,N_24722);
xor U28886 (N_28886,N_21223,N_24227);
or U28887 (N_28887,N_22371,N_22950);
nand U28888 (N_28888,N_24181,N_23699);
and U28889 (N_28889,N_21616,N_24987);
nand U28890 (N_28890,N_22234,N_24352);
nand U28891 (N_28891,N_22598,N_20892);
xnor U28892 (N_28892,N_20264,N_21493);
nor U28893 (N_28893,N_24792,N_24190);
nor U28894 (N_28894,N_23403,N_22830);
or U28895 (N_28895,N_23797,N_22685);
nand U28896 (N_28896,N_21305,N_23348);
and U28897 (N_28897,N_20007,N_23179);
xnor U28898 (N_28898,N_21246,N_20785);
and U28899 (N_28899,N_23772,N_20057);
nor U28900 (N_28900,N_21509,N_21239);
nor U28901 (N_28901,N_21838,N_20573);
nor U28902 (N_28902,N_21789,N_24671);
and U28903 (N_28903,N_21130,N_24272);
xor U28904 (N_28904,N_21316,N_20885);
or U28905 (N_28905,N_20561,N_21200);
or U28906 (N_28906,N_22926,N_22270);
nor U28907 (N_28907,N_24350,N_21074);
nand U28908 (N_28908,N_24000,N_22718);
xnor U28909 (N_28909,N_24749,N_20419);
nor U28910 (N_28910,N_22472,N_24485);
nor U28911 (N_28911,N_21562,N_20593);
and U28912 (N_28912,N_20369,N_22887);
nor U28913 (N_28913,N_22271,N_22543);
xnor U28914 (N_28914,N_21579,N_24911);
xor U28915 (N_28915,N_24526,N_21494);
or U28916 (N_28916,N_22082,N_21112);
or U28917 (N_28917,N_23208,N_20426);
or U28918 (N_28918,N_21105,N_24422);
nor U28919 (N_28919,N_23750,N_20131);
nand U28920 (N_28920,N_21233,N_20974);
nand U28921 (N_28921,N_21115,N_23586);
or U28922 (N_28922,N_20883,N_22602);
and U28923 (N_28923,N_23419,N_21976);
nor U28924 (N_28924,N_21626,N_22763);
nand U28925 (N_28925,N_21176,N_20924);
nor U28926 (N_28926,N_20354,N_23202);
nor U28927 (N_28927,N_22416,N_21549);
or U28928 (N_28928,N_20218,N_20760);
nor U28929 (N_28929,N_24300,N_20458);
or U28930 (N_28930,N_20488,N_22968);
nor U28931 (N_28931,N_24078,N_20846);
and U28932 (N_28932,N_22676,N_21896);
and U28933 (N_28933,N_20986,N_20647);
nor U28934 (N_28934,N_23697,N_21865);
and U28935 (N_28935,N_20711,N_20715);
or U28936 (N_28936,N_21668,N_23493);
nand U28937 (N_28937,N_22964,N_23993);
and U28938 (N_28938,N_21028,N_20597);
nor U28939 (N_28939,N_23000,N_22900);
and U28940 (N_28940,N_23165,N_23419);
or U28941 (N_28941,N_22019,N_21124);
xnor U28942 (N_28942,N_20557,N_21292);
or U28943 (N_28943,N_20722,N_24216);
or U28944 (N_28944,N_20762,N_20875);
or U28945 (N_28945,N_21870,N_20383);
xnor U28946 (N_28946,N_22173,N_24760);
nand U28947 (N_28947,N_21362,N_23892);
xnor U28948 (N_28948,N_20042,N_22942);
xor U28949 (N_28949,N_21311,N_23286);
xnor U28950 (N_28950,N_23176,N_21431);
xor U28951 (N_28951,N_20955,N_22418);
nor U28952 (N_28952,N_23444,N_23903);
or U28953 (N_28953,N_23666,N_23571);
nor U28954 (N_28954,N_23633,N_20108);
xor U28955 (N_28955,N_21932,N_22881);
and U28956 (N_28956,N_23412,N_20006);
xor U28957 (N_28957,N_24937,N_24189);
nor U28958 (N_28958,N_24300,N_24897);
or U28959 (N_28959,N_21113,N_24716);
xor U28960 (N_28960,N_23335,N_20271);
xor U28961 (N_28961,N_23376,N_21529);
and U28962 (N_28962,N_24868,N_20871);
and U28963 (N_28963,N_24542,N_23901);
nor U28964 (N_28964,N_21831,N_23863);
or U28965 (N_28965,N_22918,N_21726);
xnor U28966 (N_28966,N_23953,N_20897);
nand U28967 (N_28967,N_20845,N_20722);
xor U28968 (N_28968,N_22671,N_21259);
nor U28969 (N_28969,N_23979,N_22930);
nor U28970 (N_28970,N_24109,N_22786);
nand U28971 (N_28971,N_21189,N_23462);
nor U28972 (N_28972,N_23871,N_22659);
nor U28973 (N_28973,N_20404,N_21852);
and U28974 (N_28974,N_21428,N_20862);
nor U28975 (N_28975,N_21538,N_20421);
nand U28976 (N_28976,N_20456,N_20049);
and U28977 (N_28977,N_23393,N_21407);
nor U28978 (N_28978,N_20951,N_23792);
or U28979 (N_28979,N_23818,N_21034);
and U28980 (N_28980,N_23000,N_20079);
or U28981 (N_28981,N_21923,N_23324);
xnor U28982 (N_28982,N_23308,N_20637);
or U28983 (N_28983,N_21306,N_20797);
xor U28984 (N_28984,N_23072,N_22977);
nor U28985 (N_28985,N_22363,N_23972);
nor U28986 (N_28986,N_21947,N_21600);
or U28987 (N_28987,N_24650,N_20154);
xor U28988 (N_28988,N_24310,N_22847);
or U28989 (N_28989,N_21690,N_23170);
and U28990 (N_28990,N_22363,N_21788);
or U28991 (N_28991,N_22973,N_23728);
nand U28992 (N_28992,N_22907,N_23580);
nand U28993 (N_28993,N_24386,N_20102);
and U28994 (N_28994,N_24940,N_20439);
xor U28995 (N_28995,N_24222,N_22962);
nand U28996 (N_28996,N_24088,N_23443);
and U28997 (N_28997,N_22861,N_24521);
or U28998 (N_28998,N_22439,N_23864);
xnor U28999 (N_28999,N_20426,N_21796);
nor U29000 (N_29000,N_20515,N_21678);
and U29001 (N_29001,N_22983,N_24567);
nand U29002 (N_29002,N_20442,N_24584);
nand U29003 (N_29003,N_23987,N_24499);
nand U29004 (N_29004,N_22563,N_24611);
xnor U29005 (N_29005,N_22560,N_20876);
and U29006 (N_29006,N_20562,N_20956);
and U29007 (N_29007,N_23703,N_20763);
xor U29008 (N_29008,N_22993,N_21788);
xnor U29009 (N_29009,N_21519,N_24818);
nor U29010 (N_29010,N_21034,N_24585);
or U29011 (N_29011,N_21103,N_22957);
nor U29012 (N_29012,N_22304,N_20268);
and U29013 (N_29013,N_23750,N_22019);
xnor U29014 (N_29014,N_20715,N_23811);
xor U29015 (N_29015,N_22790,N_23039);
nor U29016 (N_29016,N_24160,N_22563);
and U29017 (N_29017,N_23434,N_22188);
or U29018 (N_29018,N_21121,N_24232);
nand U29019 (N_29019,N_21510,N_20721);
xnor U29020 (N_29020,N_23162,N_21272);
xnor U29021 (N_29021,N_22970,N_21691);
and U29022 (N_29022,N_20686,N_24571);
or U29023 (N_29023,N_21928,N_20842);
nor U29024 (N_29024,N_23136,N_24765);
xnor U29025 (N_29025,N_20021,N_24849);
or U29026 (N_29026,N_23811,N_22907);
xnor U29027 (N_29027,N_22367,N_24207);
nor U29028 (N_29028,N_21986,N_22464);
and U29029 (N_29029,N_21314,N_23314);
nand U29030 (N_29030,N_24603,N_24840);
nor U29031 (N_29031,N_21689,N_22650);
nor U29032 (N_29032,N_20461,N_23573);
nand U29033 (N_29033,N_20594,N_20348);
and U29034 (N_29034,N_22114,N_24384);
xnor U29035 (N_29035,N_22650,N_24657);
nand U29036 (N_29036,N_21337,N_24888);
nand U29037 (N_29037,N_21906,N_22239);
xor U29038 (N_29038,N_22434,N_23082);
or U29039 (N_29039,N_20279,N_24079);
nor U29040 (N_29040,N_23669,N_20530);
nand U29041 (N_29041,N_23883,N_24352);
nor U29042 (N_29042,N_24045,N_20615);
and U29043 (N_29043,N_21509,N_20373);
or U29044 (N_29044,N_20343,N_23325);
nor U29045 (N_29045,N_22273,N_20020);
and U29046 (N_29046,N_20263,N_21149);
or U29047 (N_29047,N_23594,N_23718);
nand U29048 (N_29048,N_21643,N_24478);
or U29049 (N_29049,N_22792,N_20217);
xnor U29050 (N_29050,N_22819,N_21257);
and U29051 (N_29051,N_23768,N_22204);
nand U29052 (N_29052,N_22030,N_23356);
xor U29053 (N_29053,N_21007,N_23048);
nor U29054 (N_29054,N_20105,N_22976);
nand U29055 (N_29055,N_22735,N_20815);
nand U29056 (N_29056,N_21345,N_22528);
and U29057 (N_29057,N_21634,N_20284);
nor U29058 (N_29058,N_23898,N_24884);
or U29059 (N_29059,N_24748,N_23327);
and U29060 (N_29060,N_21157,N_21831);
nor U29061 (N_29061,N_23510,N_21545);
nor U29062 (N_29062,N_24936,N_24506);
xnor U29063 (N_29063,N_23608,N_22462);
nand U29064 (N_29064,N_23086,N_20216);
nand U29065 (N_29065,N_23751,N_24646);
nand U29066 (N_29066,N_20001,N_24028);
and U29067 (N_29067,N_21284,N_22165);
and U29068 (N_29068,N_24372,N_24245);
and U29069 (N_29069,N_21909,N_22155);
nor U29070 (N_29070,N_21013,N_22178);
nor U29071 (N_29071,N_22722,N_23800);
nand U29072 (N_29072,N_23817,N_24224);
nor U29073 (N_29073,N_20332,N_20233);
nand U29074 (N_29074,N_22215,N_23926);
or U29075 (N_29075,N_22447,N_21649);
nand U29076 (N_29076,N_22446,N_20563);
or U29077 (N_29077,N_24585,N_24388);
nor U29078 (N_29078,N_23458,N_21624);
or U29079 (N_29079,N_22317,N_24833);
xor U29080 (N_29080,N_24053,N_21781);
xnor U29081 (N_29081,N_23009,N_21496);
and U29082 (N_29082,N_23346,N_24051);
or U29083 (N_29083,N_24493,N_21275);
xor U29084 (N_29084,N_23616,N_20536);
xor U29085 (N_29085,N_22913,N_23391);
nand U29086 (N_29086,N_22999,N_20731);
xnor U29087 (N_29087,N_24090,N_24064);
and U29088 (N_29088,N_21734,N_22699);
nor U29089 (N_29089,N_21390,N_24808);
nor U29090 (N_29090,N_21467,N_21426);
nor U29091 (N_29091,N_20858,N_24951);
xnor U29092 (N_29092,N_20768,N_23898);
and U29093 (N_29093,N_22093,N_22619);
nor U29094 (N_29094,N_22814,N_21189);
nor U29095 (N_29095,N_22621,N_22609);
nand U29096 (N_29096,N_22523,N_21436);
nor U29097 (N_29097,N_21914,N_21060);
nand U29098 (N_29098,N_24779,N_20456);
xor U29099 (N_29099,N_24889,N_24034);
nand U29100 (N_29100,N_24555,N_20318);
xnor U29101 (N_29101,N_23540,N_21431);
or U29102 (N_29102,N_22915,N_21450);
and U29103 (N_29103,N_20737,N_20596);
and U29104 (N_29104,N_23619,N_22774);
xor U29105 (N_29105,N_20887,N_21788);
nor U29106 (N_29106,N_20956,N_20732);
and U29107 (N_29107,N_20470,N_24357);
nor U29108 (N_29108,N_21528,N_20021);
xnor U29109 (N_29109,N_21890,N_24716);
and U29110 (N_29110,N_23081,N_20796);
and U29111 (N_29111,N_24641,N_23238);
nor U29112 (N_29112,N_20524,N_24350);
xnor U29113 (N_29113,N_23501,N_24778);
and U29114 (N_29114,N_20814,N_23479);
or U29115 (N_29115,N_24008,N_24545);
nand U29116 (N_29116,N_20976,N_20478);
nor U29117 (N_29117,N_23861,N_23978);
nand U29118 (N_29118,N_22495,N_20168);
or U29119 (N_29119,N_23660,N_24290);
and U29120 (N_29120,N_24204,N_21424);
and U29121 (N_29121,N_24889,N_23452);
xor U29122 (N_29122,N_22615,N_23752);
xor U29123 (N_29123,N_24531,N_22033);
xnor U29124 (N_29124,N_21598,N_21298);
xor U29125 (N_29125,N_23833,N_20853);
or U29126 (N_29126,N_22149,N_24470);
and U29127 (N_29127,N_23755,N_21393);
nand U29128 (N_29128,N_23992,N_23132);
and U29129 (N_29129,N_22459,N_22350);
nor U29130 (N_29130,N_24239,N_22523);
nand U29131 (N_29131,N_20651,N_24667);
xnor U29132 (N_29132,N_20189,N_22745);
nor U29133 (N_29133,N_20701,N_22364);
or U29134 (N_29134,N_20120,N_20271);
or U29135 (N_29135,N_20110,N_24883);
or U29136 (N_29136,N_23485,N_20782);
or U29137 (N_29137,N_24488,N_23719);
xor U29138 (N_29138,N_24104,N_23054);
and U29139 (N_29139,N_22811,N_22382);
xor U29140 (N_29140,N_24356,N_22259);
or U29141 (N_29141,N_23817,N_21984);
or U29142 (N_29142,N_22822,N_24488);
nor U29143 (N_29143,N_21267,N_21561);
or U29144 (N_29144,N_24328,N_21555);
or U29145 (N_29145,N_24256,N_21866);
nand U29146 (N_29146,N_22917,N_23824);
nand U29147 (N_29147,N_23768,N_20200);
nand U29148 (N_29148,N_21717,N_22414);
nand U29149 (N_29149,N_21728,N_24140);
nor U29150 (N_29150,N_23496,N_20033);
xor U29151 (N_29151,N_24478,N_24406);
nor U29152 (N_29152,N_22029,N_20550);
xor U29153 (N_29153,N_24326,N_22764);
or U29154 (N_29154,N_24159,N_21972);
xor U29155 (N_29155,N_20103,N_23312);
and U29156 (N_29156,N_21123,N_21511);
nor U29157 (N_29157,N_21584,N_24826);
xnor U29158 (N_29158,N_22694,N_21626);
nand U29159 (N_29159,N_23348,N_20463);
or U29160 (N_29160,N_23953,N_23419);
xnor U29161 (N_29161,N_20198,N_21893);
xor U29162 (N_29162,N_24492,N_20290);
or U29163 (N_29163,N_20570,N_24288);
nand U29164 (N_29164,N_22384,N_22171);
xnor U29165 (N_29165,N_24904,N_21951);
nor U29166 (N_29166,N_23287,N_24345);
nand U29167 (N_29167,N_24512,N_21533);
nor U29168 (N_29168,N_24467,N_24226);
xor U29169 (N_29169,N_23505,N_24644);
nor U29170 (N_29170,N_22986,N_24998);
nand U29171 (N_29171,N_20320,N_24130);
and U29172 (N_29172,N_20749,N_20820);
nand U29173 (N_29173,N_23716,N_20675);
xnor U29174 (N_29174,N_20007,N_24797);
or U29175 (N_29175,N_24811,N_20640);
nor U29176 (N_29176,N_21180,N_23911);
or U29177 (N_29177,N_24582,N_24473);
and U29178 (N_29178,N_22516,N_23306);
and U29179 (N_29179,N_20228,N_22215);
and U29180 (N_29180,N_22479,N_22429);
xnor U29181 (N_29181,N_22897,N_20230);
xor U29182 (N_29182,N_21246,N_23011);
or U29183 (N_29183,N_22923,N_21999);
nor U29184 (N_29184,N_21295,N_23976);
nor U29185 (N_29185,N_23969,N_21931);
nor U29186 (N_29186,N_24733,N_22553);
and U29187 (N_29187,N_21483,N_22835);
or U29188 (N_29188,N_21129,N_22057);
nor U29189 (N_29189,N_20963,N_23709);
nand U29190 (N_29190,N_22576,N_23884);
or U29191 (N_29191,N_24992,N_21895);
and U29192 (N_29192,N_20160,N_20416);
or U29193 (N_29193,N_20503,N_22840);
xnor U29194 (N_29194,N_24984,N_22765);
nor U29195 (N_29195,N_22345,N_21839);
and U29196 (N_29196,N_24881,N_24418);
and U29197 (N_29197,N_23822,N_24533);
nor U29198 (N_29198,N_21278,N_21248);
or U29199 (N_29199,N_21369,N_24061);
nand U29200 (N_29200,N_24724,N_22210);
nand U29201 (N_29201,N_22226,N_23033);
or U29202 (N_29202,N_21274,N_22386);
nand U29203 (N_29203,N_21347,N_20016);
nor U29204 (N_29204,N_22427,N_23669);
xor U29205 (N_29205,N_20851,N_23663);
and U29206 (N_29206,N_20971,N_24571);
nand U29207 (N_29207,N_20098,N_20474);
and U29208 (N_29208,N_21678,N_21644);
nor U29209 (N_29209,N_23726,N_22269);
and U29210 (N_29210,N_20952,N_24595);
nor U29211 (N_29211,N_23137,N_20879);
and U29212 (N_29212,N_23680,N_22111);
nand U29213 (N_29213,N_20645,N_21976);
xnor U29214 (N_29214,N_22767,N_20666);
nand U29215 (N_29215,N_24770,N_20160);
nor U29216 (N_29216,N_23024,N_24901);
or U29217 (N_29217,N_22711,N_23350);
and U29218 (N_29218,N_24351,N_20447);
xor U29219 (N_29219,N_20291,N_24794);
nand U29220 (N_29220,N_23981,N_23139);
nor U29221 (N_29221,N_21801,N_22638);
nor U29222 (N_29222,N_23789,N_20152);
and U29223 (N_29223,N_23977,N_22078);
or U29224 (N_29224,N_24516,N_23260);
nor U29225 (N_29225,N_24677,N_21922);
or U29226 (N_29226,N_20167,N_23485);
nor U29227 (N_29227,N_20742,N_20001);
nand U29228 (N_29228,N_24373,N_20653);
or U29229 (N_29229,N_20829,N_21171);
xor U29230 (N_29230,N_24362,N_22039);
or U29231 (N_29231,N_20989,N_23422);
or U29232 (N_29232,N_20478,N_24889);
xor U29233 (N_29233,N_24174,N_23945);
and U29234 (N_29234,N_20228,N_22242);
and U29235 (N_29235,N_20348,N_21585);
or U29236 (N_29236,N_22545,N_21721);
nand U29237 (N_29237,N_23862,N_22715);
nand U29238 (N_29238,N_22207,N_24644);
or U29239 (N_29239,N_24340,N_22046);
xnor U29240 (N_29240,N_23667,N_20627);
nor U29241 (N_29241,N_20396,N_20646);
and U29242 (N_29242,N_24577,N_24061);
or U29243 (N_29243,N_20140,N_22163);
nand U29244 (N_29244,N_23703,N_21971);
xnor U29245 (N_29245,N_20455,N_22955);
xor U29246 (N_29246,N_20192,N_24561);
and U29247 (N_29247,N_20026,N_21417);
nand U29248 (N_29248,N_22447,N_21985);
xor U29249 (N_29249,N_22163,N_22970);
nor U29250 (N_29250,N_24995,N_20273);
nand U29251 (N_29251,N_22546,N_21315);
nor U29252 (N_29252,N_24927,N_22328);
nand U29253 (N_29253,N_24064,N_20848);
or U29254 (N_29254,N_24817,N_23450);
nor U29255 (N_29255,N_21184,N_21360);
or U29256 (N_29256,N_20838,N_23192);
xnor U29257 (N_29257,N_21109,N_23415);
nor U29258 (N_29258,N_24780,N_21640);
xor U29259 (N_29259,N_22909,N_24797);
and U29260 (N_29260,N_22392,N_22201);
nand U29261 (N_29261,N_21978,N_20988);
or U29262 (N_29262,N_20845,N_24915);
and U29263 (N_29263,N_21048,N_21816);
nand U29264 (N_29264,N_24998,N_23736);
nand U29265 (N_29265,N_24291,N_22380);
and U29266 (N_29266,N_20191,N_24914);
nor U29267 (N_29267,N_21473,N_22408);
xor U29268 (N_29268,N_24878,N_22887);
nand U29269 (N_29269,N_24962,N_23350);
nand U29270 (N_29270,N_22362,N_21348);
nand U29271 (N_29271,N_21460,N_20433);
nand U29272 (N_29272,N_21714,N_23492);
nand U29273 (N_29273,N_22774,N_21811);
nor U29274 (N_29274,N_24293,N_22438);
nor U29275 (N_29275,N_24559,N_22191);
xnor U29276 (N_29276,N_23878,N_21062);
nand U29277 (N_29277,N_20975,N_24271);
nand U29278 (N_29278,N_24241,N_24899);
nor U29279 (N_29279,N_20690,N_20914);
xor U29280 (N_29280,N_24852,N_22532);
and U29281 (N_29281,N_24045,N_21384);
nor U29282 (N_29282,N_22557,N_23164);
xor U29283 (N_29283,N_21399,N_23175);
and U29284 (N_29284,N_24854,N_22214);
and U29285 (N_29285,N_24389,N_24931);
or U29286 (N_29286,N_24314,N_24321);
nand U29287 (N_29287,N_22468,N_20136);
or U29288 (N_29288,N_20190,N_21219);
nand U29289 (N_29289,N_22929,N_22640);
and U29290 (N_29290,N_24265,N_22673);
nor U29291 (N_29291,N_24365,N_23025);
or U29292 (N_29292,N_24577,N_22238);
nand U29293 (N_29293,N_21293,N_24403);
and U29294 (N_29294,N_21850,N_23866);
nor U29295 (N_29295,N_20811,N_22279);
nand U29296 (N_29296,N_23484,N_24803);
nand U29297 (N_29297,N_23414,N_21248);
nand U29298 (N_29298,N_24165,N_20290);
or U29299 (N_29299,N_23835,N_21536);
nand U29300 (N_29300,N_22676,N_20165);
or U29301 (N_29301,N_20807,N_22115);
xor U29302 (N_29302,N_23309,N_20067);
xor U29303 (N_29303,N_22702,N_24901);
xor U29304 (N_29304,N_20910,N_24802);
xnor U29305 (N_29305,N_24911,N_21245);
or U29306 (N_29306,N_20167,N_21327);
or U29307 (N_29307,N_23970,N_23920);
nor U29308 (N_29308,N_21827,N_24987);
or U29309 (N_29309,N_24184,N_24673);
nor U29310 (N_29310,N_22351,N_21536);
nor U29311 (N_29311,N_23767,N_22069);
or U29312 (N_29312,N_21758,N_23166);
nor U29313 (N_29313,N_22733,N_23271);
or U29314 (N_29314,N_23785,N_23240);
xor U29315 (N_29315,N_24440,N_24965);
nand U29316 (N_29316,N_22545,N_20416);
or U29317 (N_29317,N_24042,N_22436);
and U29318 (N_29318,N_22249,N_23294);
and U29319 (N_29319,N_21366,N_24668);
nand U29320 (N_29320,N_24737,N_22881);
and U29321 (N_29321,N_20945,N_24205);
nand U29322 (N_29322,N_22649,N_20237);
and U29323 (N_29323,N_22323,N_22320);
xor U29324 (N_29324,N_20450,N_21983);
and U29325 (N_29325,N_20333,N_21431);
xor U29326 (N_29326,N_22596,N_22564);
nor U29327 (N_29327,N_21309,N_23894);
or U29328 (N_29328,N_23847,N_24542);
and U29329 (N_29329,N_23207,N_24863);
or U29330 (N_29330,N_23457,N_22317);
nor U29331 (N_29331,N_21838,N_21904);
nor U29332 (N_29332,N_22777,N_24780);
nor U29333 (N_29333,N_21448,N_21384);
or U29334 (N_29334,N_21086,N_23583);
or U29335 (N_29335,N_20728,N_24217);
xnor U29336 (N_29336,N_20003,N_20951);
xor U29337 (N_29337,N_20480,N_22068);
or U29338 (N_29338,N_21899,N_24976);
or U29339 (N_29339,N_21092,N_23911);
xnor U29340 (N_29340,N_24872,N_21253);
xnor U29341 (N_29341,N_24182,N_23167);
nand U29342 (N_29342,N_23600,N_24378);
nor U29343 (N_29343,N_24534,N_22550);
xor U29344 (N_29344,N_22964,N_24274);
nor U29345 (N_29345,N_22165,N_24038);
and U29346 (N_29346,N_20195,N_21336);
nor U29347 (N_29347,N_23481,N_22583);
or U29348 (N_29348,N_20637,N_21744);
or U29349 (N_29349,N_21620,N_24940);
or U29350 (N_29350,N_24928,N_23293);
or U29351 (N_29351,N_20227,N_22948);
nand U29352 (N_29352,N_21163,N_24519);
nand U29353 (N_29353,N_22124,N_23527);
and U29354 (N_29354,N_22369,N_21903);
or U29355 (N_29355,N_22971,N_23895);
xor U29356 (N_29356,N_22377,N_23562);
xnor U29357 (N_29357,N_24466,N_24448);
nor U29358 (N_29358,N_24414,N_23474);
or U29359 (N_29359,N_24618,N_22595);
xor U29360 (N_29360,N_24424,N_23212);
and U29361 (N_29361,N_21983,N_21776);
and U29362 (N_29362,N_21365,N_20026);
xor U29363 (N_29363,N_24151,N_20340);
nor U29364 (N_29364,N_23632,N_21519);
or U29365 (N_29365,N_21839,N_24349);
xnor U29366 (N_29366,N_24942,N_23328);
and U29367 (N_29367,N_23799,N_20645);
or U29368 (N_29368,N_24024,N_24648);
nand U29369 (N_29369,N_20081,N_24802);
and U29370 (N_29370,N_24334,N_22987);
nor U29371 (N_29371,N_20395,N_20003);
and U29372 (N_29372,N_21163,N_21762);
nand U29373 (N_29373,N_22610,N_24264);
nor U29374 (N_29374,N_20826,N_23456);
xor U29375 (N_29375,N_23191,N_20815);
nor U29376 (N_29376,N_23884,N_21799);
nand U29377 (N_29377,N_20952,N_23243);
nand U29378 (N_29378,N_22609,N_22692);
and U29379 (N_29379,N_20275,N_22048);
nand U29380 (N_29380,N_22864,N_21582);
or U29381 (N_29381,N_24060,N_24669);
and U29382 (N_29382,N_23511,N_20883);
and U29383 (N_29383,N_20050,N_22602);
nand U29384 (N_29384,N_20300,N_21844);
nor U29385 (N_29385,N_20428,N_23653);
nor U29386 (N_29386,N_24718,N_22494);
xor U29387 (N_29387,N_24286,N_24470);
nand U29388 (N_29388,N_23768,N_24043);
nand U29389 (N_29389,N_20594,N_23509);
nor U29390 (N_29390,N_24938,N_23048);
and U29391 (N_29391,N_21160,N_22904);
nor U29392 (N_29392,N_22954,N_24639);
and U29393 (N_29393,N_20139,N_22688);
nand U29394 (N_29394,N_20238,N_22854);
or U29395 (N_29395,N_22260,N_24412);
nand U29396 (N_29396,N_22492,N_23752);
xnor U29397 (N_29397,N_22130,N_24181);
nor U29398 (N_29398,N_22983,N_21789);
nand U29399 (N_29399,N_24422,N_23143);
and U29400 (N_29400,N_20684,N_22526);
nor U29401 (N_29401,N_21184,N_23843);
and U29402 (N_29402,N_24780,N_22514);
xnor U29403 (N_29403,N_24653,N_23648);
xnor U29404 (N_29404,N_22451,N_24140);
xnor U29405 (N_29405,N_24546,N_22614);
or U29406 (N_29406,N_21959,N_22877);
xor U29407 (N_29407,N_24186,N_20484);
xnor U29408 (N_29408,N_21715,N_24456);
and U29409 (N_29409,N_21720,N_24671);
xor U29410 (N_29410,N_22065,N_22963);
or U29411 (N_29411,N_24468,N_20244);
nor U29412 (N_29412,N_24771,N_20266);
nand U29413 (N_29413,N_22198,N_24086);
and U29414 (N_29414,N_21789,N_23837);
xor U29415 (N_29415,N_20112,N_23561);
or U29416 (N_29416,N_21409,N_21807);
and U29417 (N_29417,N_23862,N_23489);
nand U29418 (N_29418,N_24317,N_21021);
nor U29419 (N_29419,N_22331,N_20191);
xnor U29420 (N_29420,N_21157,N_21207);
nor U29421 (N_29421,N_22490,N_21555);
nand U29422 (N_29422,N_24941,N_20173);
nand U29423 (N_29423,N_24074,N_24750);
nand U29424 (N_29424,N_21414,N_22206);
nor U29425 (N_29425,N_24231,N_23169);
and U29426 (N_29426,N_20902,N_24759);
and U29427 (N_29427,N_21438,N_24969);
nand U29428 (N_29428,N_23872,N_24147);
xor U29429 (N_29429,N_21002,N_22226);
and U29430 (N_29430,N_20791,N_21482);
xor U29431 (N_29431,N_21569,N_23024);
nor U29432 (N_29432,N_22218,N_20149);
xor U29433 (N_29433,N_22526,N_20513);
nor U29434 (N_29434,N_24059,N_24341);
nand U29435 (N_29435,N_22625,N_20614);
nor U29436 (N_29436,N_20596,N_23392);
and U29437 (N_29437,N_22982,N_21510);
and U29438 (N_29438,N_20360,N_22084);
nor U29439 (N_29439,N_21753,N_22077);
and U29440 (N_29440,N_22612,N_24031);
nand U29441 (N_29441,N_22817,N_22185);
or U29442 (N_29442,N_23624,N_21527);
and U29443 (N_29443,N_23836,N_20315);
or U29444 (N_29444,N_22842,N_23685);
nand U29445 (N_29445,N_20645,N_23128);
nor U29446 (N_29446,N_20982,N_22960);
or U29447 (N_29447,N_23186,N_22745);
or U29448 (N_29448,N_24855,N_21206);
xnor U29449 (N_29449,N_22990,N_22139);
nor U29450 (N_29450,N_23322,N_22692);
xnor U29451 (N_29451,N_22661,N_23231);
xor U29452 (N_29452,N_23835,N_21085);
nand U29453 (N_29453,N_21045,N_23634);
and U29454 (N_29454,N_24856,N_23523);
or U29455 (N_29455,N_20948,N_23119);
nor U29456 (N_29456,N_21365,N_21089);
or U29457 (N_29457,N_24888,N_24338);
nand U29458 (N_29458,N_22561,N_20841);
nand U29459 (N_29459,N_20835,N_22580);
and U29460 (N_29460,N_21262,N_22271);
nor U29461 (N_29461,N_24731,N_24779);
xnor U29462 (N_29462,N_22891,N_22118);
or U29463 (N_29463,N_23681,N_23492);
or U29464 (N_29464,N_23207,N_24329);
nand U29465 (N_29465,N_23965,N_20631);
nand U29466 (N_29466,N_22131,N_24055);
nor U29467 (N_29467,N_20306,N_21659);
nand U29468 (N_29468,N_24796,N_20011);
nor U29469 (N_29469,N_22385,N_21140);
and U29470 (N_29470,N_23220,N_23429);
nor U29471 (N_29471,N_21750,N_21870);
nor U29472 (N_29472,N_23500,N_21518);
or U29473 (N_29473,N_21133,N_23409);
and U29474 (N_29474,N_24098,N_24643);
or U29475 (N_29475,N_20482,N_21416);
nand U29476 (N_29476,N_24903,N_21655);
nor U29477 (N_29477,N_22626,N_21770);
and U29478 (N_29478,N_22518,N_21009);
nor U29479 (N_29479,N_24088,N_22123);
and U29480 (N_29480,N_22285,N_21763);
nor U29481 (N_29481,N_24823,N_24052);
nor U29482 (N_29482,N_24579,N_24569);
and U29483 (N_29483,N_23000,N_21382);
nor U29484 (N_29484,N_22015,N_21412);
nor U29485 (N_29485,N_24793,N_22992);
or U29486 (N_29486,N_24218,N_21745);
nor U29487 (N_29487,N_23928,N_22208);
nor U29488 (N_29488,N_20234,N_20808);
xor U29489 (N_29489,N_22288,N_23102);
xnor U29490 (N_29490,N_23865,N_24291);
xor U29491 (N_29491,N_24737,N_21696);
or U29492 (N_29492,N_20998,N_22015);
or U29493 (N_29493,N_20570,N_24363);
xor U29494 (N_29494,N_21533,N_22966);
and U29495 (N_29495,N_22319,N_24960);
nor U29496 (N_29496,N_22310,N_21660);
nand U29497 (N_29497,N_21804,N_23327);
nor U29498 (N_29498,N_20736,N_24498);
xnor U29499 (N_29499,N_20338,N_22324);
nor U29500 (N_29500,N_20512,N_23602);
nand U29501 (N_29501,N_21229,N_24291);
nand U29502 (N_29502,N_21930,N_23935);
xnor U29503 (N_29503,N_20728,N_24051);
xor U29504 (N_29504,N_24915,N_21502);
nor U29505 (N_29505,N_24696,N_24371);
nand U29506 (N_29506,N_22994,N_24263);
or U29507 (N_29507,N_22351,N_22922);
or U29508 (N_29508,N_20506,N_22965);
nor U29509 (N_29509,N_20213,N_22586);
nor U29510 (N_29510,N_20133,N_22424);
xnor U29511 (N_29511,N_22771,N_23096);
nand U29512 (N_29512,N_24661,N_24840);
or U29513 (N_29513,N_21624,N_23957);
nor U29514 (N_29514,N_22648,N_24927);
and U29515 (N_29515,N_21577,N_23674);
or U29516 (N_29516,N_24167,N_22133);
nand U29517 (N_29517,N_21143,N_24464);
or U29518 (N_29518,N_22286,N_22360);
and U29519 (N_29519,N_21182,N_20601);
or U29520 (N_29520,N_24782,N_23680);
or U29521 (N_29521,N_24255,N_20530);
nand U29522 (N_29522,N_22312,N_21005);
and U29523 (N_29523,N_23772,N_21839);
nor U29524 (N_29524,N_22644,N_21887);
and U29525 (N_29525,N_21013,N_22205);
or U29526 (N_29526,N_24991,N_22079);
and U29527 (N_29527,N_20032,N_21838);
and U29528 (N_29528,N_21795,N_23453);
xnor U29529 (N_29529,N_21718,N_21048);
nor U29530 (N_29530,N_24572,N_20048);
nand U29531 (N_29531,N_22867,N_24125);
nor U29532 (N_29532,N_21795,N_24240);
or U29533 (N_29533,N_24476,N_23524);
and U29534 (N_29534,N_23555,N_23908);
and U29535 (N_29535,N_23505,N_20653);
or U29536 (N_29536,N_23542,N_23244);
nand U29537 (N_29537,N_22645,N_24734);
xnor U29538 (N_29538,N_23182,N_24443);
and U29539 (N_29539,N_22513,N_24759);
and U29540 (N_29540,N_24551,N_22125);
or U29541 (N_29541,N_24830,N_24757);
or U29542 (N_29542,N_23068,N_21910);
xnor U29543 (N_29543,N_20057,N_24260);
and U29544 (N_29544,N_22348,N_22643);
nand U29545 (N_29545,N_21099,N_21491);
nor U29546 (N_29546,N_21330,N_22374);
xor U29547 (N_29547,N_23458,N_22657);
nand U29548 (N_29548,N_21185,N_23386);
nor U29549 (N_29549,N_21070,N_23232);
nor U29550 (N_29550,N_20161,N_21668);
xnor U29551 (N_29551,N_22661,N_23382);
xor U29552 (N_29552,N_24680,N_20146);
xor U29553 (N_29553,N_21165,N_24531);
nand U29554 (N_29554,N_21215,N_23699);
nand U29555 (N_29555,N_24343,N_24906);
xnor U29556 (N_29556,N_20398,N_24834);
and U29557 (N_29557,N_24882,N_22545);
and U29558 (N_29558,N_21224,N_21429);
or U29559 (N_29559,N_20292,N_21504);
and U29560 (N_29560,N_21196,N_24698);
nand U29561 (N_29561,N_22715,N_21882);
and U29562 (N_29562,N_20213,N_23262);
and U29563 (N_29563,N_20303,N_20807);
and U29564 (N_29564,N_21703,N_22185);
or U29565 (N_29565,N_24842,N_23701);
xnor U29566 (N_29566,N_24686,N_22983);
nor U29567 (N_29567,N_24685,N_23244);
nand U29568 (N_29568,N_23672,N_23298);
xor U29569 (N_29569,N_23482,N_21196);
nand U29570 (N_29570,N_22912,N_24351);
or U29571 (N_29571,N_24730,N_21594);
nand U29572 (N_29572,N_20261,N_21581);
nor U29573 (N_29573,N_20128,N_21002);
or U29574 (N_29574,N_24592,N_24971);
and U29575 (N_29575,N_23106,N_20566);
nand U29576 (N_29576,N_24014,N_23379);
xor U29577 (N_29577,N_23085,N_23088);
nor U29578 (N_29578,N_24628,N_20875);
and U29579 (N_29579,N_22405,N_24470);
nor U29580 (N_29580,N_20340,N_23191);
nand U29581 (N_29581,N_22648,N_21843);
nor U29582 (N_29582,N_21854,N_22352);
nand U29583 (N_29583,N_21696,N_24404);
xor U29584 (N_29584,N_20670,N_23497);
xor U29585 (N_29585,N_20114,N_21759);
and U29586 (N_29586,N_20633,N_20501);
nand U29587 (N_29587,N_21074,N_21891);
or U29588 (N_29588,N_24730,N_22475);
or U29589 (N_29589,N_22725,N_21328);
nand U29590 (N_29590,N_22273,N_22804);
and U29591 (N_29591,N_23605,N_23224);
or U29592 (N_29592,N_24106,N_21078);
nand U29593 (N_29593,N_20025,N_20784);
nand U29594 (N_29594,N_21593,N_21993);
or U29595 (N_29595,N_24660,N_22424);
and U29596 (N_29596,N_20042,N_24199);
nor U29597 (N_29597,N_22593,N_23200);
or U29598 (N_29598,N_21752,N_24801);
or U29599 (N_29599,N_21820,N_22538);
and U29600 (N_29600,N_24222,N_22277);
nand U29601 (N_29601,N_23623,N_23937);
nor U29602 (N_29602,N_23125,N_20283);
nor U29603 (N_29603,N_22124,N_21919);
nand U29604 (N_29604,N_21388,N_21165);
nand U29605 (N_29605,N_22613,N_22750);
nor U29606 (N_29606,N_21898,N_21996);
or U29607 (N_29607,N_22787,N_20108);
and U29608 (N_29608,N_24142,N_20248);
nor U29609 (N_29609,N_22918,N_20422);
or U29610 (N_29610,N_22338,N_21276);
or U29611 (N_29611,N_21346,N_20165);
nor U29612 (N_29612,N_24755,N_24640);
nand U29613 (N_29613,N_24714,N_21863);
nor U29614 (N_29614,N_20941,N_22181);
or U29615 (N_29615,N_23570,N_23942);
and U29616 (N_29616,N_23864,N_24652);
nand U29617 (N_29617,N_21898,N_21297);
nand U29618 (N_29618,N_24351,N_24588);
nor U29619 (N_29619,N_21380,N_20791);
nor U29620 (N_29620,N_23980,N_24692);
xor U29621 (N_29621,N_24643,N_24733);
nand U29622 (N_29622,N_24019,N_22723);
nand U29623 (N_29623,N_23972,N_22906);
xnor U29624 (N_29624,N_23276,N_22128);
xor U29625 (N_29625,N_24647,N_23988);
nand U29626 (N_29626,N_22455,N_23014);
or U29627 (N_29627,N_20618,N_21232);
nand U29628 (N_29628,N_22460,N_21332);
nor U29629 (N_29629,N_22878,N_22853);
or U29630 (N_29630,N_23745,N_23061);
nand U29631 (N_29631,N_20798,N_22178);
nand U29632 (N_29632,N_23061,N_21723);
or U29633 (N_29633,N_24736,N_23353);
nor U29634 (N_29634,N_22376,N_21429);
and U29635 (N_29635,N_20977,N_20625);
or U29636 (N_29636,N_20858,N_20236);
and U29637 (N_29637,N_21922,N_23514);
nand U29638 (N_29638,N_22494,N_20575);
xnor U29639 (N_29639,N_24141,N_20514);
xor U29640 (N_29640,N_20148,N_23680);
or U29641 (N_29641,N_23897,N_23380);
nor U29642 (N_29642,N_23789,N_23495);
and U29643 (N_29643,N_23660,N_24442);
or U29644 (N_29644,N_24493,N_20545);
and U29645 (N_29645,N_23584,N_20359);
xor U29646 (N_29646,N_21334,N_24230);
xor U29647 (N_29647,N_24124,N_20792);
xor U29648 (N_29648,N_23583,N_20130);
nand U29649 (N_29649,N_24832,N_24336);
nor U29650 (N_29650,N_24055,N_24401);
or U29651 (N_29651,N_23038,N_23932);
nor U29652 (N_29652,N_20904,N_23525);
xor U29653 (N_29653,N_24435,N_21483);
nand U29654 (N_29654,N_24235,N_21833);
nand U29655 (N_29655,N_24737,N_24394);
nand U29656 (N_29656,N_24754,N_23918);
nor U29657 (N_29657,N_20468,N_21491);
nand U29658 (N_29658,N_22638,N_20748);
or U29659 (N_29659,N_24687,N_22666);
nor U29660 (N_29660,N_22841,N_20843);
nand U29661 (N_29661,N_20119,N_23855);
xor U29662 (N_29662,N_23493,N_21392);
or U29663 (N_29663,N_20314,N_20929);
nor U29664 (N_29664,N_23281,N_24525);
nor U29665 (N_29665,N_23128,N_24169);
and U29666 (N_29666,N_20741,N_24542);
xnor U29667 (N_29667,N_24146,N_24202);
xnor U29668 (N_29668,N_22864,N_23614);
nand U29669 (N_29669,N_22025,N_20225);
or U29670 (N_29670,N_24914,N_22615);
xnor U29671 (N_29671,N_23455,N_21679);
and U29672 (N_29672,N_24752,N_21813);
or U29673 (N_29673,N_22879,N_21814);
xor U29674 (N_29674,N_20639,N_21350);
or U29675 (N_29675,N_24640,N_20910);
nand U29676 (N_29676,N_24065,N_20334);
or U29677 (N_29677,N_20850,N_21344);
or U29678 (N_29678,N_24443,N_20322);
and U29679 (N_29679,N_21350,N_22064);
xnor U29680 (N_29680,N_23282,N_24583);
nand U29681 (N_29681,N_20832,N_21213);
nand U29682 (N_29682,N_24418,N_22148);
and U29683 (N_29683,N_22126,N_22976);
nand U29684 (N_29684,N_22139,N_20197);
nand U29685 (N_29685,N_23717,N_21177);
xor U29686 (N_29686,N_23460,N_21453);
xnor U29687 (N_29687,N_20675,N_21704);
and U29688 (N_29688,N_24754,N_20944);
or U29689 (N_29689,N_21685,N_24390);
xor U29690 (N_29690,N_21122,N_21793);
nand U29691 (N_29691,N_24052,N_21633);
nand U29692 (N_29692,N_22841,N_20679);
or U29693 (N_29693,N_24793,N_21439);
xnor U29694 (N_29694,N_20531,N_22328);
xnor U29695 (N_29695,N_20505,N_21454);
nor U29696 (N_29696,N_23296,N_20167);
nand U29697 (N_29697,N_21856,N_22923);
nand U29698 (N_29698,N_24102,N_24840);
nand U29699 (N_29699,N_22368,N_24642);
nand U29700 (N_29700,N_23380,N_24960);
and U29701 (N_29701,N_23500,N_24648);
nand U29702 (N_29702,N_21887,N_24103);
and U29703 (N_29703,N_21523,N_22827);
and U29704 (N_29704,N_22777,N_21953);
or U29705 (N_29705,N_22456,N_20871);
and U29706 (N_29706,N_20960,N_22070);
nand U29707 (N_29707,N_24755,N_23097);
or U29708 (N_29708,N_20533,N_22697);
nor U29709 (N_29709,N_22981,N_22480);
nor U29710 (N_29710,N_22866,N_20164);
or U29711 (N_29711,N_24066,N_21966);
or U29712 (N_29712,N_21152,N_23165);
nor U29713 (N_29713,N_20008,N_21296);
and U29714 (N_29714,N_20027,N_24438);
nand U29715 (N_29715,N_20006,N_22591);
xor U29716 (N_29716,N_23835,N_20897);
xnor U29717 (N_29717,N_23605,N_22678);
nand U29718 (N_29718,N_23202,N_22349);
xnor U29719 (N_29719,N_20266,N_22017);
nor U29720 (N_29720,N_22191,N_21312);
nor U29721 (N_29721,N_24802,N_23271);
and U29722 (N_29722,N_20987,N_22794);
nand U29723 (N_29723,N_21950,N_23768);
nand U29724 (N_29724,N_20106,N_22928);
nand U29725 (N_29725,N_23663,N_21903);
xor U29726 (N_29726,N_22899,N_23547);
nand U29727 (N_29727,N_24617,N_24046);
and U29728 (N_29728,N_24157,N_20625);
and U29729 (N_29729,N_20190,N_24591);
or U29730 (N_29730,N_21917,N_21784);
nand U29731 (N_29731,N_21707,N_24254);
or U29732 (N_29732,N_22483,N_24091);
and U29733 (N_29733,N_20436,N_21901);
nor U29734 (N_29734,N_24527,N_21558);
or U29735 (N_29735,N_22785,N_21916);
xnor U29736 (N_29736,N_20868,N_20598);
or U29737 (N_29737,N_24165,N_20035);
xor U29738 (N_29738,N_20707,N_22942);
xor U29739 (N_29739,N_24094,N_24598);
xor U29740 (N_29740,N_20213,N_24719);
xor U29741 (N_29741,N_21161,N_20061);
xnor U29742 (N_29742,N_20692,N_24806);
and U29743 (N_29743,N_20288,N_23699);
nor U29744 (N_29744,N_22428,N_23044);
or U29745 (N_29745,N_23661,N_20015);
or U29746 (N_29746,N_22023,N_20117);
nand U29747 (N_29747,N_24831,N_24696);
nand U29748 (N_29748,N_23832,N_22145);
nor U29749 (N_29749,N_23692,N_21827);
nor U29750 (N_29750,N_23332,N_22126);
and U29751 (N_29751,N_21547,N_24359);
nand U29752 (N_29752,N_24013,N_24121);
xnor U29753 (N_29753,N_22765,N_22597);
xnor U29754 (N_29754,N_20471,N_22680);
or U29755 (N_29755,N_24215,N_23163);
nand U29756 (N_29756,N_22334,N_24495);
or U29757 (N_29757,N_23832,N_24220);
nor U29758 (N_29758,N_24441,N_22693);
xnor U29759 (N_29759,N_23338,N_21762);
nor U29760 (N_29760,N_24365,N_24844);
and U29761 (N_29761,N_22418,N_24169);
and U29762 (N_29762,N_21543,N_23172);
and U29763 (N_29763,N_24308,N_23782);
or U29764 (N_29764,N_22452,N_24941);
and U29765 (N_29765,N_20727,N_24057);
nor U29766 (N_29766,N_24395,N_21987);
or U29767 (N_29767,N_21866,N_22377);
and U29768 (N_29768,N_21365,N_23529);
or U29769 (N_29769,N_22121,N_20109);
and U29770 (N_29770,N_24220,N_23461);
nand U29771 (N_29771,N_21589,N_23065);
or U29772 (N_29772,N_21911,N_23509);
and U29773 (N_29773,N_24403,N_24037);
and U29774 (N_29774,N_20151,N_21267);
xnor U29775 (N_29775,N_21585,N_22978);
xor U29776 (N_29776,N_20412,N_23846);
and U29777 (N_29777,N_20415,N_24585);
nand U29778 (N_29778,N_24152,N_22951);
or U29779 (N_29779,N_24680,N_20887);
or U29780 (N_29780,N_24953,N_23960);
nand U29781 (N_29781,N_21690,N_22517);
or U29782 (N_29782,N_23956,N_21525);
and U29783 (N_29783,N_20102,N_22808);
and U29784 (N_29784,N_20537,N_23559);
nand U29785 (N_29785,N_20489,N_20208);
xnor U29786 (N_29786,N_24271,N_24994);
nand U29787 (N_29787,N_24713,N_24649);
nor U29788 (N_29788,N_22794,N_21693);
nand U29789 (N_29789,N_20587,N_24092);
nor U29790 (N_29790,N_22254,N_24603);
nand U29791 (N_29791,N_20867,N_24280);
and U29792 (N_29792,N_24589,N_20382);
or U29793 (N_29793,N_20823,N_24952);
or U29794 (N_29794,N_21309,N_24332);
nor U29795 (N_29795,N_24619,N_22608);
nor U29796 (N_29796,N_21831,N_23463);
nand U29797 (N_29797,N_22683,N_23461);
nand U29798 (N_29798,N_20682,N_22996);
or U29799 (N_29799,N_23983,N_23541);
nor U29800 (N_29800,N_24561,N_24796);
or U29801 (N_29801,N_22861,N_24184);
and U29802 (N_29802,N_22175,N_20413);
and U29803 (N_29803,N_24071,N_23390);
nor U29804 (N_29804,N_24994,N_24403);
nand U29805 (N_29805,N_22812,N_20071);
and U29806 (N_29806,N_23827,N_20491);
nand U29807 (N_29807,N_24707,N_24827);
nand U29808 (N_29808,N_22499,N_21527);
xor U29809 (N_29809,N_20433,N_22516);
xnor U29810 (N_29810,N_22850,N_23212);
xnor U29811 (N_29811,N_24702,N_23723);
xnor U29812 (N_29812,N_23039,N_20298);
nor U29813 (N_29813,N_21102,N_20644);
and U29814 (N_29814,N_23714,N_21636);
nand U29815 (N_29815,N_22407,N_21081);
or U29816 (N_29816,N_24615,N_20377);
nor U29817 (N_29817,N_21391,N_24917);
nor U29818 (N_29818,N_21525,N_22368);
nor U29819 (N_29819,N_20896,N_22977);
or U29820 (N_29820,N_24893,N_23820);
nor U29821 (N_29821,N_22331,N_20850);
xnor U29822 (N_29822,N_20038,N_21193);
or U29823 (N_29823,N_23276,N_23549);
or U29824 (N_29824,N_23740,N_23835);
nand U29825 (N_29825,N_24913,N_21514);
nand U29826 (N_29826,N_24032,N_23428);
nand U29827 (N_29827,N_24098,N_22637);
and U29828 (N_29828,N_23083,N_24494);
xor U29829 (N_29829,N_20805,N_22190);
or U29830 (N_29830,N_20104,N_23244);
nor U29831 (N_29831,N_23517,N_22997);
or U29832 (N_29832,N_21635,N_21862);
nor U29833 (N_29833,N_21132,N_24411);
nor U29834 (N_29834,N_20977,N_22679);
nor U29835 (N_29835,N_23950,N_22345);
nand U29836 (N_29836,N_24208,N_23814);
or U29837 (N_29837,N_20127,N_21830);
and U29838 (N_29838,N_24858,N_20996);
or U29839 (N_29839,N_23968,N_22216);
or U29840 (N_29840,N_24463,N_20436);
xor U29841 (N_29841,N_24538,N_20642);
and U29842 (N_29842,N_24264,N_23793);
or U29843 (N_29843,N_22842,N_20611);
xnor U29844 (N_29844,N_20477,N_24658);
or U29845 (N_29845,N_21492,N_22827);
or U29846 (N_29846,N_22768,N_24819);
nor U29847 (N_29847,N_22340,N_21568);
and U29848 (N_29848,N_21011,N_24974);
nor U29849 (N_29849,N_22369,N_21413);
xnor U29850 (N_29850,N_22722,N_20661);
nand U29851 (N_29851,N_23021,N_20849);
or U29852 (N_29852,N_21302,N_21334);
nand U29853 (N_29853,N_22288,N_21123);
nand U29854 (N_29854,N_20842,N_21580);
nand U29855 (N_29855,N_20158,N_23951);
xnor U29856 (N_29856,N_22382,N_22012);
nor U29857 (N_29857,N_21708,N_20742);
nand U29858 (N_29858,N_20191,N_21964);
or U29859 (N_29859,N_21522,N_24499);
and U29860 (N_29860,N_20717,N_24832);
nor U29861 (N_29861,N_20614,N_20535);
or U29862 (N_29862,N_24303,N_24680);
nand U29863 (N_29863,N_22967,N_22956);
or U29864 (N_29864,N_23136,N_24457);
or U29865 (N_29865,N_20072,N_22089);
nor U29866 (N_29866,N_20285,N_24177);
nand U29867 (N_29867,N_24741,N_20333);
and U29868 (N_29868,N_24111,N_20415);
nor U29869 (N_29869,N_24343,N_22378);
nor U29870 (N_29870,N_23348,N_22441);
nor U29871 (N_29871,N_21939,N_22049);
nor U29872 (N_29872,N_21757,N_20687);
or U29873 (N_29873,N_21909,N_22599);
xnor U29874 (N_29874,N_22866,N_20849);
and U29875 (N_29875,N_22864,N_21557);
nand U29876 (N_29876,N_22986,N_23731);
nor U29877 (N_29877,N_21438,N_21194);
and U29878 (N_29878,N_23825,N_23392);
and U29879 (N_29879,N_22456,N_23406);
xor U29880 (N_29880,N_21260,N_21021);
nand U29881 (N_29881,N_24724,N_24495);
or U29882 (N_29882,N_20926,N_24183);
and U29883 (N_29883,N_23382,N_22694);
xor U29884 (N_29884,N_22051,N_24370);
nand U29885 (N_29885,N_23507,N_21661);
or U29886 (N_29886,N_22285,N_20861);
nand U29887 (N_29887,N_23484,N_20545);
and U29888 (N_29888,N_24518,N_23797);
nor U29889 (N_29889,N_21630,N_24445);
nand U29890 (N_29890,N_20301,N_23199);
and U29891 (N_29891,N_20245,N_21572);
and U29892 (N_29892,N_20071,N_21860);
nand U29893 (N_29893,N_21207,N_22456);
xnor U29894 (N_29894,N_23277,N_23851);
and U29895 (N_29895,N_23563,N_24559);
or U29896 (N_29896,N_22407,N_24649);
nand U29897 (N_29897,N_22289,N_21294);
xor U29898 (N_29898,N_20064,N_22196);
xor U29899 (N_29899,N_23880,N_21283);
xnor U29900 (N_29900,N_22221,N_20290);
xor U29901 (N_29901,N_22319,N_23451);
nor U29902 (N_29902,N_21890,N_21691);
or U29903 (N_29903,N_24031,N_24483);
or U29904 (N_29904,N_22599,N_24306);
xnor U29905 (N_29905,N_21888,N_24466);
nor U29906 (N_29906,N_21008,N_22647);
and U29907 (N_29907,N_24790,N_24546);
or U29908 (N_29908,N_22165,N_21448);
nor U29909 (N_29909,N_23527,N_20451);
nand U29910 (N_29910,N_23390,N_21143);
or U29911 (N_29911,N_20503,N_22771);
nor U29912 (N_29912,N_20536,N_21228);
or U29913 (N_29913,N_21753,N_23598);
and U29914 (N_29914,N_23165,N_24140);
xnor U29915 (N_29915,N_21425,N_24236);
xor U29916 (N_29916,N_24597,N_20321);
nor U29917 (N_29917,N_24935,N_23529);
nor U29918 (N_29918,N_23863,N_20085);
and U29919 (N_29919,N_24554,N_23161);
xnor U29920 (N_29920,N_24208,N_23045);
or U29921 (N_29921,N_21682,N_20129);
or U29922 (N_29922,N_20216,N_21487);
nand U29923 (N_29923,N_21848,N_23657);
nor U29924 (N_29924,N_22489,N_20457);
xor U29925 (N_29925,N_22853,N_20057);
or U29926 (N_29926,N_22347,N_21027);
xor U29927 (N_29927,N_21280,N_23823);
xor U29928 (N_29928,N_23243,N_21584);
or U29929 (N_29929,N_23987,N_24898);
nor U29930 (N_29930,N_24426,N_22313);
xor U29931 (N_29931,N_21629,N_21707);
xnor U29932 (N_29932,N_20662,N_24495);
and U29933 (N_29933,N_23933,N_22177);
or U29934 (N_29934,N_20702,N_24454);
nor U29935 (N_29935,N_21828,N_23713);
xnor U29936 (N_29936,N_22718,N_23114);
and U29937 (N_29937,N_24297,N_22385);
nand U29938 (N_29938,N_24422,N_22018);
nor U29939 (N_29939,N_24991,N_20246);
or U29940 (N_29940,N_21490,N_24698);
nor U29941 (N_29941,N_20555,N_20449);
and U29942 (N_29942,N_23131,N_24474);
nand U29943 (N_29943,N_21516,N_22652);
and U29944 (N_29944,N_24869,N_22790);
nand U29945 (N_29945,N_20946,N_21079);
nand U29946 (N_29946,N_21106,N_21519);
xor U29947 (N_29947,N_23649,N_21894);
nand U29948 (N_29948,N_20103,N_20825);
nor U29949 (N_29949,N_22183,N_20042);
nand U29950 (N_29950,N_24372,N_21100);
xnor U29951 (N_29951,N_23048,N_20652);
nor U29952 (N_29952,N_21266,N_23472);
or U29953 (N_29953,N_23436,N_20565);
nand U29954 (N_29954,N_24428,N_22160);
and U29955 (N_29955,N_23650,N_21622);
and U29956 (N_29956,N_23578,N_23952);
nor U29957 (N_29957,N_20194,N_23698);
nor U29958 (N_29958,N_21163,N_22041);
or U29959 (N_29959,N_23989,N_22704);
xnor U29960 (N_29960,N_24999,N_22164);
nand U29961 (N_29961,N_24037,N_21604);
nor U29962 (N_29962,N_21724,N_24480);
xnor U29963 (N_29963,N_24764,N_22050);
nor U29964 (N_29964,N_22163,N_23146);
xnor U29965 (N_29965,N_24206,N_22469);
nor U29966 (N_29966,N_23946,N_22751);
nor U29967 (N_29967,N_24010,N_23147);
or U29968 (N_29968,N_24810,N_21454);
or U29969 (N_29969,N_24065,N_22988);
xor U29970 (N_29970,N_22502,N_21147);
xor U29971 (N_29971,N_20229,N_20529);
and U29972 (N_29972,N_24296,N_21542);
nand U29973 (N_29973,N_23204,N_21165);
or U29974 (N_29974,N_24254,N_21011);
or U29975 (N_29975,N_22883,N_20102);
xor U29976 (N_29976,N_24591,N_21877);
xor U29977 (N_29977,N_24112,N_21705);
or U29978 (N_29978,N_23354,N_21778);
nand U29979 (N_29979,N_21387,N_21659);
xor U29980 (N_29980,N_24637,N_20169);
xor U29981 (N_29981,N_24703,N_22046);
xnor U29982 (N_29982,N_20381,N_24535);
nor U29983 (N_29983,N_21940,N_20902);
and U29984 (N_29984,N_24571,N_22091);
nand U29985 (N_29985,N_23756,N_23997);
nand U29986 (N_29986,N_24651,N_21283);
nor U29987 (N_29987,N_20425,N_23452);
nand U29988 (N_29988,N_22406,N_23067);
nor U29989 (N_29989,N_20145,N_21336);
and U29990 (N_29990,N_24530,N_24510);
nand U29991 (N_29991,N_22646,N_24045);
nor U29992 (N_29992,N_21177,N_20598);
xor U29993 (N_29993,N_21076,N_24400);
or U29994 (N_29994,N_22495,N_24178);
or U29995 (N_29995,N_21319,N_23118);
xor U29996 (N_29996,N_20316,N_23642);
nand U29997 (N_29997,N_22238,N_20330);
xnor U29998 (N_29998,N_21232,N_24884);
xor U29999 (N_29999,N_21776,N_24977);
and U30000 (N_30000,N_29260,N_27304);
or U30001 (N_30001,N_29817,N_26880);
xnor U30002 (N_30002,N_29488,N_27743);
nor U30003 (N_30003,N_29111,N_26315);
and U30004 (N_30004,N_26760,N_29615);
xnor U30005 (N_30005,N_27133,N_29469);
xor U30006 (N_30006,N_28176,N_29419);
or U30007 (N_30007,N_29002,N_27604);
and U30008 (N_30008,N_29290,N_27835);
nand U30009 (N_30009,N_27961,N_28254);
or U30010 (N_30010,N_29439,N_27605);
and U30011 (N_30011,N_27795,N_29377);
and U30012 (N_30012,N_26106,N_28087);
xnor U30013 (N_30013,N_26447,N_28285);
and U30014 (N_30014,N_27053,N_25549);
and U30015 (N_30015,N_27817,N_27325);
nand U30016 (N_30016,N_26318,N_25037);
or U30017 (N_30017,N_25003,N_29974);
nor U30018 (N_30018,N_25820,N_27942);
xor U30019 (N_30019,N_28315,N_27348);
and U30020 (N_30020,N_29385,N_27326);
nor U30021 (N_30021,N_25294,N_28999);
or U30022 (N_30022,N_29578,N_26790);
or U30023 (N_30023,N_28183,N_26301);
and U30024 (N_30024,N_29356,N_27566);
or U30025 (N_30025,N_29969,N_25725);
and U30026 (N_30026,N_26319,N_29534);
xor U30027 (N_30027,N_27969,N_25778);
or U30028 (N_30028,N_27346,N_27812);
nor U30029 (N_30029,N_27054,N_29651);
or U30030 (N_30030,N_29941,N_28495);
nor U30031 (N_30031,N_26683,N_26486);
xnor U30032 (N_30032,N_25584,N_25144);
and U30033 (N_30033,N_29898,N_29593);
nor U30034 (N_30034,N_28415,N_25284);
nor U30035 (N_30035,N_25949,N_29727);
and U30036 (N_30036,N_29850,N_28963);
nand U30037 (N_30037,N_26182,N_27366);
nand U30038 (N_30038,N_29499,N_29863);
or U30039 (N_30039,N_29884,N_27957);
or U30040 (N_30040,N_26293,N_25127);
nor U30041 (N_30041,N_25086,N_27117);
nand U30042 (N_30042,N_28652,N_26172);
and U30043 (N_30043,N_26767,N_29476);
nor U30044 (N_30044,N_27824,N_25557);
and U30045 (N_30045,N_26498,N_26845);
xnor U30046 (N_30046,N_25743,N_29920);
nand U30047 (N_30047,N_29177,N_26809);
or U30048 (N_30048,N_26402,N_28655);
nor U30049 (N_30049,N_28420,N_27268);
nand U30050 (N_30050,N_26549,N_27241);
nand U30051 (N_30051,N_26739,N_26704);
xor U30052 (N_30052,N_26951,N_28596);
nand U30053 (N_30053,N_26735,N_28128);
and U30054 (N_30054,N_27678,N_27970);
xor U30055 (N_30055,N_25221,N_27912);
nor U30056 (N_30056,N_26088,N_27881);
or U30057 (N_30057,N_27293,N_25385);
nor U30058 (N_30058,N_25435,N_26964);
and U30059 (N_30059,N_27676,N_25984);
nand U30060 (N_30060,N_28390,N_27918);
xnor U30061 (N_30061,N_25645,N_27659);
xor U30062 (N_30062,N_28160,N_27550);
xor U30063 (N_30063,N_29066,N_26371);
or U30064 (N_30064,N_27525,N_26522);
or U30065 (N_30065,N_25338,N_25030);
nand U30066 (N_30066,N_28123,N_26677);
xor U30067 (N_30067,N_26868,N_27426);
nor U30068 (N_30068,N_29130,N_29880);
or U30069 (N_30069,N_27548,N_25275);
or U30070 (N_30070,N_29720,N_26632);
and U30071 (N_30071,N_29360,N_25678);
xor U30072 (N_30072,N_25696,N_27224);
nand U30073 (N_30073,N_27171,N_25379);
nor U30074 (N_30074,N_27438,N_26574);
nand U30075 (N_30075,N_25561,N_27288);
nand U30076 (N_30076,N_29473,N_28565);
nand U30077 (N_30077,N_28671,N_27768);
xor U30078 (N_30078,N_26703,N_26785);
nor U30079 (N_30079,N_29363,N_28525);
nor U30080 (N_30080,N_25912,N_28832);
and U30081 (N_30081,N_26456,N_26882);
nor U30082 (N_30082,N_29313,N_29565);
or U30083 (N_30083,N_28981,N_29386);
and U30084 (N_30084,N_27492,N_28593);
nor U30085 (N_30085,N_26600,N_26277);
and U30086 (N_30086,N_28738,N_28580);
or U30087 (N_30087,N_29885,N_29187);
nor U30088 (N_30088,N_25403,N_25100);
and U30089 (N_30089,N_29163,N_25257);
or U30090 (N_30090,N_26709,N_25384);
xnor U30091 (N_30091,N_25703,N_27526);
and U30092 (N_30092,N_28629,N_25442);
nor U30093 (N_30093,N_27986,N_29082);
or U30094 (N_30094,N_29086,N_28098);
nor U30095 (N_30095,N_29547,N_28897);
nand U30096 (N_30096,N_28196,N_29027);
nand U30097 (N_30097,N_26359,N_25859);
and U30098 (N_30098,N_26786,N_28812);
xnor U30099 (N_30099,N_26637,N_26471);
and U30100 (N_30100,N_26516,N_26733);
and U30101 (N_30101,N_27593,N_27352);
nor U30102 (N_30102,N_27746,N_29459);
nand U30103 (N_30103,N_27946,N_26451);
or U30104 (N_30104,N_26343,N_29810);
nor U30105 (N_30105,N_29116,N_28319);
nor U30106 (N_30106,N_27156,N_26997);
and U30107 (N_30107,N_28635,N_27335);
nand U30108 (N_30108,N_27757,N_25963);
nor U30109 (N_30109,N_29460,N_25489);
and U30110 (N_30110,N_29512,N_27359);
and U30111 (N_30111,N_29814,N_26240);
or U30112 (N_30112,N_26808,N_29945);
and U30113 (N_30113,N_26353,N_26229);
nor U30114 (N_30114,N_28190,N_29596);
or U30115 (N_30115,N_27370,N_29126);
and U30116 (N_30116,N_28186,N_29959);
nand U30117 (N_30117,N_28218,N_29550);
xor U30118 (N_30118,N_26261,N_29120);
xor U30119 (N_30119,N_27447,N_28006);
nor U30120 (N_30120,N_27238,N_28450);
nand U30121 (N_30121,N_26089,N_27916);
nor U30122 (N_30122,N_26420,N_28851);
nand U30123 (N_30123,N_27523,N_27564);
or U30124 (N_30124,N_29014,N_27032);
or U30125 (N_30125,N_28368,N_28025);
nor U30126 (N_30126,N_27497,N_28120);
nor U30127 (N_30127,N_29455,N_25755);
and U30128 (N_30128,N_29140,N_26365);
or U30129 (N_30129,N_25594,N_25835);
or U30130 (N_30130,N_28866,N_28181);
and U30131 (N_30131,N_25577,N_27882);
or U30132 (N_30132,N_28735,N_28797);
and U30133 (N_30133,N_27384,N_25461);
or U30134 (N_30134,N_26598,N_25791);
nor U30135 (N_30135,N_26531,N_26769);
xor U30136 (N_30136,N_29859,N_29673);
and U30137 (N_30137,N_25234,N_26025);
and U30138 (N_30138,N_27730,N_26814);
nor U30139 (N_30139,N_25992,N_25097);
and U30140 (N_30140,N_25323,N_26092);
and U30141 (N_30141,N_27467,N_28037);
and U30142 (N_30142,N_29607,N_29680);
nor U30143 (N_30143,N_25058,N_26164);
and U30144 (N_30144,N_26244,N_29368);
or U30145 (N_30145,N_28323,N_28017);
xor U30146 (N_30146,N_27199,N_29235);
nand U30147 (N_30147,N_27189,N_28592);
nand U30148 (N_30148,N_27388,N_29504);
or U30149 (N_30149,N_29211,N_27994);
nand U30150 (N_30150,N_28284,N_27381);
xor U30151 (N_30151,N_25299,N_26864);
nand U30152 (N_30152,N_29277,N_27985);
nand U30153 (N_30153,N_28957,N_25940);
nand U30154 (N_30154,N_29824,N_29767);
and U30155 (N_30155,N_26298,N_25776);
and U30156 (N_30156,N_25015,N_28211);
and U30157 (N_30157,N_26855,N_25140);
nand U30158 (N_30158,N_26362,N_27483);
or U30159 (N_30159,N_27434,N_25961);
or U30160 (N_30160,N_29761,N_29675);
nor U30161 (N_30161,N_25865,N_29273);
or U30162 (N_30162,N_27193,N_29521);
xor U30163 (N_30163,N_26278,N_25125);
xnor U30164 (N_30164,N_29792,N_29339);
nand U30165 (N_30165,N_28949,N_26387);
xor U30166 (N_30166,N_29876,N_26995);
nor U30167 (N_30167,N_27614,N_27377);
or U30168 (N_30168,N_26994,N_25325);
and U30169 (N_30169,N_26428,N_29015);
nand U30170 (N_30170,N_28551,N_25064);
nand U30171 (N_30171,N_29878,N_29097);
or U30172 (N_30172,N_28440,N_25170);
xnor U30173 (N_30173,N_26552,N_27867);
nor U30174 (N_30174,N_25602,N_26701);
nand U30175 (N_30175,N_28153,N_28443);
nand U30176 (N_30176,N_25295,N_26884);
and U30177 (N_30177,N_28760,N_27580);
nor U30178 (N_30178,N_29394,N_29216);
nand U30179 (N_30179,N_25191,N_25365);
or U30180 (N_30180,N_27670,N_27724);
nand U30181 (N_30181,N_27919,N_29156);
xor U30182 (N_30182,N_25981,N_26817);
nand U30183 (N_30183,N_29361,N_26504);
nor U30184 (N_30184,N_25516,N_27302);
nor U30185 (N_30185,N_28562,N_25884);
nor U30186 (N_30186,N_28118,N_25406);
xor U30187 (N_30187,N_25334,N_28626);
nand U30188 (N_30188,N_27488,N_29838);
or U30189 (N_30189,N_25149,N_29653);
or U30190 (N_30190,N_27265,N_27131);
and U30191 (N_30191,N_28257,N_25027);
nand U30192 (N_30192,N_26251,N_29826);
and U30193 (N_30193,N_28387,N_26573);
or U30194 (N_30194,N_26751,N_29463);
nand U30195 (N_30195,N_25559,N_27274);
xor U30196 (N_30196,N_27926,N_28825);
or U30197 (N_30197,N_29400,N_29695);
nand U30198 (N_30198,N_26840,N_29319);
xnor U30199 (N_30199,N_29533,N_25508);
and U30200 (N_30200,N_28479,N_25157);
nand U30201 (N_30201,N_29042,N_29035);
and U30202 (N_30202,N_26892,N_25563);
and U30203 (N_30203,N_27530,N_25651);
nor U30204 (N_30204,N_25395,N_28732);
nand U30205 (N_30205,N_26539,N_26140);
nor U30206 (N_30206,N_26779,N_25335);
and U30207 (N_30207,N_25415,N_25288);
or U30208 (N_30208,N_27841,N_28520);
xnor U30209 (N_30209,N_27857,N_29248);
xor U30210 (N_30210,N_26485,N_28365);
and U30211 (N_30211,N_26466,N_25811);
nor U30212 (N_30212,N_25239,N_29839);
and U30213 (N_30213,N_25204,N_27754);
or U30214 (N_30214,N_29404,N_29094);
and U30215 (N_30215,N_26437,N_28276);
and U30216 (N_30216,N_29879,N_29167);
or U30217 (N_30217,N_26519,N_26288);
nand U30218 (N_30218,N_26854,N_28436);
xnor U30219 (N_30219,N_29435,N_26233);
and U30220 (N_30220,N_26592,N_27071);
xor U30221 (N_30221,N_27365,N_25950);
nand U30222 (N_30222,N_25908,N_25095);
or U30223 (N_30223,N_25844,N_25034);
nor U30224 (N_30224,N_29833,N_25972);
nand U30225 (N_30225,N_28528,N_28513);
nor U30226 (N_30226,N_27278,N_29636);
xor U30227 (N_30227,N_25736,N_26440);
xor U30228 (N_30228,N_27613,N_27983);
or U30229 (N_30229,N_28489,N_27889);
or U30230 (N_30230,N_28873,N_28517);
or U30231 (N_30231,N_29338,N_26688);
nor U30232 (N_30232,N_28704,N_27089);
and U30233 (N_30233,N_25219,N_26405);
nor U30234 (N_30234,N_29519,N_27267);
xnor U30235 (N_30235,N_29152,N_25405);
nor U30236 (N_30236,N_28032,N_27554);
xor U30237 (N_30237,N_25619,N_29217);
xor U30238 (N_30238,N_26044,N_25002);
and U30239 (N_30239,N_27603,N_29413);
nand U30240 (N_30240,N_29182,N_28954);
xor U30241 (N_30241,N_28739,N_29209);
xor U30242 (N_30242,N_28793,N_28928);
nand U30243 (N_30243,N_29933,N_29210);
nand U30244 (N_30244,N_28158,N_28516);
or U30245 (N_30245,N_28075,N_27173);
and U30246 (N_30246,N_28480,N_29129);
nor U30247 (N_30247,N_25026,N_27151);
xor U30248 (N_30248,N_27445,N_26642);
nor U30249 (N_30249,N_29552,N_28983);
xor U30250 (N_30250,N_28984,N_25139);
xnor U30251 (N_30251,N_28103,N_28129);
nor U30252 (N_30252,N_29784,N_26918);
nand U30253 (N_30253,N_28990,N_26943);
and U30254 (N_30254,N_25888,N_29026);
and U30255 (N_30255,N_27466,N_26321);
and U30256 (N_30256,N_29171,N_28830);
nor U30257 (N_30257,N_25142,N_27818);
nand U30258 (N_30258,N_26793,N_26538);
or U30259 (N_30259,N_27684,N_29666);
xor U30260 (N_30260,N_29223,N_25331);
and U30261 (N_30261,N_27831,N_26056);
or U30262 (N_30262,N_28358,N_28795);
xnor U30263 (N_30263,N_29490,N_28690);
nor U30264 (N_30264,N_26376,N_27674);
or U30265 (N_30265,N_27935,N_27209);
nand U30266 (N_30266,N_27367,N_28498);
or U30267 (N_30267,N_26650,N_28349);
xnor U30268 (N_30268,N_27132,N_27476);
xnor U30269 (N_30269,N_27414,N_25350);
xor U30270 (N_30270,N_27010,N_29643);
nand U30271 (N_30271,N_27030,N_27908);
or U30272 (N_30272,N_28581,N_25396);
nor U30273 (N_30273,N_29697,N_28058);
and U30274 (N_30274,N_29254,N_26046);
nor U30275 (N_30275,N_27056,N_26936);
or U30276 (N_30276,N_27699,N_29527);
nor U30277 (N_30277,N_25803,N_29748);
and U30278 (N_30278,N_28270,N_27886);
and U30279 (N_30279,N_28606,N_29844);
xnor U30280 (N_30280,N_28609,N_25378);
nand U30281 (N_30281,N_28717,N_26924);
nand U30282 (N_30282,N_28320,N_27937);
or U30283 (N_30283,N_26896,N_25935);
nand U30284 (N_30284,N_29205,N_26553);
xor U30285 (N_30285,N_27707,N_26163);
nand U30286 (N_30286,N_28291,N_29203);
nand U30287 (N_30287,N_25550,N_26983);
nand U30288 (N_30288,N_29269,N_28012);
or U30289 (N_30289,N_25287,N_27727);
nand U30290 (N_30290,N_25460,N_27379);
nor U30291 (N_30291,N_28545,N_27158);
or U30292 (N_30292,N_26827,N_27877);
nor U30293 (N_30293,N_28624,N_28891);
xor U30294 (N_30294,N_26273,N_25737);
xor U30295 (N_30295,N_26459,N_28326);
nand U30296 (N_30296,N_27529,N_28945);
and U30297 (N_30297,N_29682,N_28811);
nand U30298 (N_30298,N_29757,N_28071);
xor U30299 (N_30299,N_25988,N_28406);
nor U30300 (N_30300,N_27277,N_26074);
and U30301 (N_30301,N_26883,N_28288);
and U30302 (N_30302,N_29153,N_26360);
nand U30303 (N_30303,N_28824,N_25428);
or U30304 (N_30304,N_29548,N_25391);
or U30305 (N_30305,N_26079,N_29347);
xnor U30306 (N_30306,N_27160,N_25271);
nor U30307 (N_30307,N_28680,N_26407);
xnor U30308 (N_30308,N_26004,N_29608);
and U30309 (N_30309,N_29921,N_26127);
nor U30310 (N_30310,N_26794,N_28558);
nand U30311 (N_30311,N_25478,N_29219);
and U30312 (N_30312,N_29856,N_26999);
xnor U30313 (N_30313,N_27111,N_25667);
xor U30314 (N_30314,N_26181,N_28715);
xnor U30315 (N_30315,N_28563,N_25790);
nand U30316 (N_30316,N_29637,N_25429);
nor U30317 (N_30317,N_27792,N_26467);
xor U30318 (N_30318,N_27082,N_27606);
nor U30319 (N_30319,N_28328,N_27140);
and U30320 (N_30320,N_28678,N_29780);
xnor U30321 (N_30321,N_26078,N_26851);
and U30322 (N_30322,N_25497,N_27034);
xor U30323 (N_30323,N_25728,N_26804);
and U30324 (N_30324,N_26116,N_28266);
and U30325 (N_30325,N_28858,N_29718);
nor U30326 (N_30326,N_29935,N_27696);
or U30327 (N_30327,N_27509,N_26661);
or U30328 (N_30328,N_27516,N_27883);
and U30329 (N_30329,N_26805,N_27294);
nand U30330 (N_30330,N_29827,N_29583);
xor U30331 (N_30331,N_28935,N_28378);
nor U30332 (N_30332,N_29947,N_29968);
xnor U30333 (N_30333,N_26155,N_26582);
xor U30334 (N_30334,N_26908,N_26307);
or U30335 (N_30335,N_29312,N_27654);
nand U30336 (N_30336,N_25475,N_26175);
and U30337 (N_30337,N_26641,N_29450);
and U30338 (N_30338,N_29261,N_27441);
nor U30339 (N_30339,N_29713,N_26558);
nor U30340 (N_30340,N_29772,N_27996);
nand U30341 (N_30341,N_28357,N_29174);
or U30342 (N_30342,N_27124,N_25321);
xor U30343 (N_30343,N_26841,N_29364);
nor U30344 (N_30344,N_25023,N_28177);
xnor U30345 (N_30345,N_27729,N_29468);
nand U30346 (N_30346,N_25094,N_26449);
nor U30347 (N_30347,N_28927,N_25909);
nand U30348 (N_30348,N_28082,N_25727);
nor U30349 (N_30349,N_25782,N_29457);
nor U30350 (N_30350,N_26103,N_29756);
nand U30351 (N_30351,N_25996,N_26835);
xor U30352 (N_30352,N_25181,N_25020);
and U30353 (N_30353,N_27280,N_25409);
or U30354 (N_30354,N_28537,N_26073);
or U30355 (N_30355,N_29796,N_29458);
and U30356 (N_30356,N_26057,N_25154);
or U30357 (N_30357,N_28380,N_27577);
nor U30358 (N_30358,N_27793,N_25322);
nor U30359 (N_30359,N_26055,N_28065);
nor U30360 (N_30360,N_28850,N_25845);
xnor U30361 (N_30361,N_27259,N_27100);
nand U30362 (N_30362,N_26090,N_26408);
nor U30363 (N_30363,N_29836,N_27971);
nand U30364 (N_30364,N_28608,N_25087);
nor U30365 (N_30365,N_28305,N_28772);
nor U30366 (N_30366,N_27805,N_28345);
nand U30367 (N_30367,N_27952,N_28731);
nor U30368 (N_30368,N_27594,N_27977);
nor U30369 (N_30369,N_27596,N_29915);
nand U30370 (N_30370,N_28461,N_26961);
nand U30371 (N_30371,N_25311,N_29694);
xnor U30372 (N_30372,N_27997,N_29809);
and U30373 (N_30373,N_26596,N_25664);
nand U30374 (N_30374,N_28800,N_29985);
nor U30375 (N_30375,N_27298,N_26570);
nand U30376 (N_30376,N_26564,N_27104);
xnor U30377 (N_30377,N_25065,N_29399);
or U30378 (N_30378,N_28615,N_28505);
and U30379 (N_30379,N_29275,N_28660);
or U30380 (N_30380,N_27430,N_26967);
nor U30381 (N_30381,N_25343,N_28556);
or U30382 (N_30382,N_27266,N_25259);
xor U30383 (N_30383,N_29415,N_27862);
or U30384 (N_30384,N_26929,N_26061);
nor U30385 (N_30385,N_27648,N_29229);
and U30386 (N_30386,N_29664,N_27907);
xor U30387 (N_30387,N_28969,N_27584);
and U30388 (N_30388,N_27582,N_25307);
nor U30389 (N_30389,N_26130,N_25432);
or U30390 (N_30390,N_26873,N_27610);
nor U30391 (N_30391,N_29284,N_28634);
xnor U30392 (N_30392,N_27092,N_28251);
nor U30393 (N_30393,N_27153,N_25357);
or U30394 (N_30394,N_25407,N_25910);
nand U30395 (N_30395,N_27642,N_29812);
nor U30396 (N_30396,N_25630,N_26458);
or U30397 (N_30397,N_25326,N_28508);
nor U30398 (N_30398,N_28669,N_28653);
or U30399 (N_30399,N_26174,N_26614);
nand U30400 (N_30400,N_29157,N_29401);
nor U30401 (N_30401,N_28370,N_27940);
or U30402 (N_30402,N_27551,N_26267);
nor U30403 (N_30403,N_26334,N_28588);
xor U30404 (N_30404,N_28217,N_26361);
nand U30405 (N_30405,N_27949,N_28676);
and U30406 (N_30406,N_25680,N_28057);
nor U30407 (N_30407,N_28256,N_29541);
xor U30408 (N_30408,N_25172,N_25555);
or U30409 (N_30409,N_26966,N_28597);
or U30410 (N_30410,N_26064,N_28777);
xor U30411 (N_30411,N_27787,N_26118);
xor U30412 (N_30412,N_27407,N_27130);
or U30413 (N_30413,N_26603,N_28815);
nor U30414 (N_30414,N_27894,N_26971);
and U30415 (N_30415,N_26448,N_29145);
nor U30416 (N_30416,N_26724,N_25768);
nor U30417 (N_30417,N_29891,N_26210);
or U30418 (N_30418,N_25558,N_28363);
nand U30419 (N_30419,N_27592,N_27932);
xnor U30420 (N_30420,N_26563,N_27500);
and U30421 (N_30421,N_29994,N_28548);
or U30422 (N_30422,N_25241,N_27892);
nand U30423 (N_30423,N_29782,N_28024);
and U30424 (N_30424,N_29676,N_27436);
nand U30425 (N_30425,N_26935,N_26262);
and U30426 (N_30426,N_28388,N_26673);
nand U30427 (N_30427,N_25861,N_26374);
xor U30428 (N_30428,N_26129,N_28268);
or U30429 (N_30429,N_26492,N_28549);
nor U30430 (N_30430,N_28998,N_27214);
or U30431 (N_30431,N_29585,N_28195);
nor U30432 (N_30432,N_27195,N_27533);
xor U30433 (N_30433,N_28574,N_25634);
xor U30434 (N_30434,N_28808,N_27815);
xor U30435 (N_30435,N_26207,N_28754);
or U30436 (N_30436,N_28023,N_25383);
nor U30437 (N_30437,N_26132,N_27044);
xnor U30438 (N_30438,N_28837,N_29904);
xnor U30439 (N_30439,N_25767,N_25423);
nand U30440 (N_30440,N_29924,N_27187);
xnor U30441 (N_30441,N_25059,N_28646);
xnor U30442 (N_30442,N_28881,N_25898);
and U30443 (N_30443,N_29158,N_29592);
and U30444 (N_30444,N_29494,N_28198);
and U30445 (N_30445,N_28852,N_25040);
and U30446 (N_30446,N_28670,N_26173);
or U30447 (N_30447,N_25240,N_27095);
nand U30448 (N_30448,N_25248,N_29428);
nor U30449 (N_30449,N_26822,N_29916);
nand U30450 (N_30450,N_26148,N_25138);
nor U30451 (N_30451,N_26748,N_28369);
nor U30452 (N_30452,N_25209,N_27383);
nand U30453 (N_30453,N_26975,N_28148);
and U30454 (N_30454,N_25991,N_28589);
or U30455 (N_30455,N_25956,N_25573);
nand U30456 (N_30456,N_25397,N_26388);
nor U30457 (N_30457,N_25067,N_28985);
nand U30458 (N_30458,N_26444,N_29906);
and U30459 (N_30459,N_25860,N_27588);
nand U30460 (N_30460,N_27682,N_28599);
xor U30461 (N_30461,N_25413,N_29530);
and U30462 (N_30462,N_25883,N_29083);
or U30463 (N_30463,N_26300,N_29305);
nor U30464 (N_30464,N_26452,N_27917);
xor U30465 (N_30465,N_29049,N_25580);
and U30466 (N_30466,N_25480,N_27735);
nor U30467 (N_30467,N_28453,N_26601);
nand U30468 (N_30468,N_28993,N_26477);
or U30469 (N_30469,N_26279,N_26100);
and U30470 (N_30470,N_27012,N_26397);
and U30471 (N_30471,N_26871,N_27794);
or U30472 (N_30472,N_26224,N_25185);
and U30473 (N_30473,N_26714,N_26096);
or U30474 (N_30474,N_25458,N_29344);
nor U30475 (N_30475,N_29293,N_25684);
nand U30476 (N_30476,N_27826,N_28847);
or U30477 (N_30477,N_26065,N_26686);
nand U30478 (N_30478,N_25608,N_27349);
xor U30479 (N_30479,N_29526,N_28447);
and U30480 (N_30480,N_25960,N_26234);
or U30481 (N_30481,N_26803,N_28767);
or U30482 (N_30482,N_27148,N_27777);
and U30483 (N_30483,N_26655,N_28871);
xor U30484 (N_30484,N_28952,N_29332);
nand U30485 (N_30485,N_25532,N_26685);
nand U30486 (N_30486,N_25669,N_29783);
and U30487 (N_30487,N_25711,N_25032);
nor U30488 (N_30488,N_27215,N_28745);
xor U30489 (N_30489,N_25151,N_29255);
and U30490 (N_30490,N_28070,N_28296);
and U30491 (N_30491,N_25527,N_26204);
and U30492 (N_30492,N_27116,N_28314);
nand U30493 (N_30493,N_29257,N_28448);
and U30494 (N_30494,N_26950,N_29725);
and U30495 (N_30495,N_28155,N_25869);
nor U30496 (N_30496,N_27261,N_25652);
xor U30497 (N_30497,N_27184,N_29687);
xnor U30498 (N_30498,N_26815,N_28689);
nand U30499 (N_30499,N_26345,N_25775);
nand U30500 (N_30500,N_27518,N_25110);
nor U30501 (N_30501,N_28553,N_29853);
and U30502 (N_30502,N_29088,N_26742);
xnor U30503 (N_30503,N_29506,N_28383);
nor U30504 (N_30504,N_26400,N_29979);
and U30505 (N_30505,N_26186,N_25253);
nor U30506 (N_30506,N_29711,N_28978);
or U30507 (N_30507,N_25566,N_25153);
nand U30508 (N_30508,N_26310,N_27600);
nor U30509 (N_30509,N_29851,N_29078);
nor U30510 (N_30510,N_28668,N_26501);
nor U30511 (N_30511,N_29905,N_27360);
xnor U30512 (N_30512,N_25313,N_28429);
and U30513 (N_30513,N_29604,N_25493);
and U30514 (N_30514,N_29102,N_27301);
xnor U30515 (N_30515,N_26659,N_25875);
and U30516 (N_30516,N_28583,N_25841);
nor U30517 (N_30517,N_28780,N_28061);
nor U30518 (N_30518,N_28557,N_26844);
or U30519 (N_30519,N_26750,N_25529);
xnor U30520 (N_30520,N_28507,N_27402);
nand U30521 (N_30521,N_29848,N_29346);
or U30522 (N_30522,N_28262,N_25606);
xnor U30523 (N_30523,N_26780,N_29251);
and U30524 (N_30524,N_27000,N_27789);
or U30525 (N_30525,N_29194,N_26797);
or U30526 (N_30526,N_27234,N_26493);
nor U30527 (N_30527,N_29840,N_27322);
nand U30528 (N_30528,N_28085,N_27495);
nand U30529 (N_30529,N_25408,N_26216);
nor U30530 (N_30530,N_28267,N_25611);
nor U30531 (N_30531,N_25045,N_26008);
nor U30532 (N_30532,N_28996,N_29333);
or U30533 (N_30533,N_27066,N_26670);
nor U30534 (N_30534,N_26001,N_26721);
nand U30535 (N_30535,N_29298,N_28527);
xor U30536 (N_30536,N_26542,N_25425);
xnor U30537 (N_30537,N_29908,N_29829);
nor U30538 (N_30538,N_28351,N_25591);
xnor U30539 (N_30539,N_25999,N_29580);
or U30540 (N_30540,N_25366,N_27972);
nand U30541 (N_30541,N_25691,N_25846);
xor U30542 (N_30542,N_25312,N_26922);
and U30543 (N_30543,N_29497,N_26366);
or U30544 (N_30544,N_27845,N_27945);
xor U30545 (N_30545,N_26612,N_29072);
and U30546 (N_30546,N_27329,N_25158);
or U30547 (N_30547,N_26023,N_27073);
nand U30548 (N_30548,N_27762,N_26465);
xnor U30549 (N_30549,N_27571,N_27599);
nand U30550 (N_30550,N_29523,N_27097);
nor U30551 (N_30551,N_28665,N_26220);
xor U30552 (N_30552,N_27305,N_25496);
nor U30553 (N_30553,N_27897,N_29150);
xnor U30554 (N_30554,N_28108,N_26027);
or U30555 (N_30555,N_27236,N_25601);
nand U30556 (N_30556,N_26607,N_28201);
nand U30557 (N_30557,N_25818,N_26135);
nand U30558 (N_30558,N_26617,N_27105);
xor U30559 (N_30559,N_26520,N_25672);
nand U30560 (N_30560,N_25482,N_26575);
and U30561 (N_30561,N_27121,N_28471);
and U30562 (N_30562,N_27216,N_29820);
nor U30563 (N_30563,N_25523,N_28199);
nor U30564 (N_30564,N_27967,N_25666);
nand U30565 (N_30565,N_26347,N_28602);
and U30566 (N_30566,N_28274,N_27773);
or U30567 (N_30567,N_27611,N_27966);
xor U30568 (N_30568,N_26215,N_28342);
xor U30569 (N_30569,N_25873,N_26047);
nor U30570 (N_30570,N_27753,N_27890);
and U30571 (N_30571,N_29096,N_25661);
xnor U30572 (N_30572,N_26996,N_26707);
nand U30573 (N_30573,N_25746,N_29927);
or U30574 (N_30574,N_28473,N_26656);
nor U30575 (N_30575,N_26867,N_29418);
xor U30576 (N_30576,N_25538,N_29751);
xor U30577 (N_30577,N_29327,N_26770);
nand U30578 (N_30578,N_26972,N_29128);
or U30579 (N_30579,N_25215,N_27312);
nor U30580 (N_30580,N_25380,N_27046);
xnor U30581 (N_30581,N_26333,N_25359);
and U30582 (N_30582,N_28788,N_25747);
xor U30583 (N_30583,N_25824,N_26968);
and U30584 (N_30584,N_28442,N_26898);
and U30585 (N_30585,N_25188,N_28905);
or U30586 (N_30586,N_26990,N_26393);
and U30587 (N_30587,N_25534,N_25685);
and U30588 (N_30588,N_25556,N_25565);
or U30589 (N_30589,N_26080,N_29503);
nand U30590 (N_30590,N_26398,N_26532);
nand U30591 (N_30591,N_29091,N_29614);
nor U30592 (N_30592,N_25255,N_27418);
xnor U30593 (N_30593,N_25544,N_25887);
nand U30594 (N_30594,N_25089,N_29487);
or U30595 (N_30595,N_26853,N_29054);
or U30596 (N_30596,N_25226,N_28360);
nand U30597 (N_30597,N_27213,N_26663);
or U30598 (N_30598,N_29553,N_26285);
and U30599 (N_30599,N_28801,N_26305);
or U30600 (N_30600,N_28004,N_26599);
xor U30601 (N_30601,N_28189,N_29232);
or U30602 (N_30602,N_28864,N_29029);
xnor U30603 (N_30603,N_27799,N_26392);
nand U30604 (N_30604,N_27231,N_29502);
nor U30605 (N_30605,N_25076,N_29073);
nand U30606 (N_30606,N_29272,N_28216);
and U30607 (N_30607,N_28988,N_26594);
nand U30608 (N_30608,N_26336,N_27398);
or U30609 (N_30609,N_27651,N_27417);
xnor U30610 (N_30610,N_27247,N_25620);
nand U30611 (N_30611,N_25128,N_28906);
nand U30612 (N_30612,N_27314,N_26513);
xnor U30613 (N_30613,N_28253,N_25631);
and U30614 (N_30614,N_29791,N_26988);
and U30615 (N_30615,N_27113,N_27263);
and U30616 (N_30616,N_29663,N_26926);
and U30617 (N_30617,N_29004,N_26734);
xnor U30618 (N_30618,N_27300,N_26317);
and U30619 (N_30619,N_27512,N_26053);
nand U30620 (N_30620,N_26264,N_26455);
or U30621 (N_30621,N_28080,N_26416);
nor U30622 (N_30622,N_27602,N_28884);
and U30623 (N_30623,N_25539,N_27775);
and U30624 (N_30624,N_28311,N_26114);
nor U30625 (N_30625,N_28675,N_29491);
and U30626 (N_30626,N_27175,N_29890);
xor U30627 (N_30627,N_28465,N_28894);
and U30628 (N_30628,N_26856,N_25175);
nor U30629 (N_30629,N_27120,N_28531);
or U30630 (N_30630,N_28003,N_26923);
nor U30631 (N_30631,N_26208,N_29017);
nor U30632 (N_30632,N_28535,N_27490);
and U30633 (N_30633,N_28681,N_26694);
nand U30634 (N_30634,N_28720,N_25261);
nand U30635 (N_30635,N_26529,N_25289);
xor U30636 (N_30636,N_29074,N_28965);
and U30637 (N_30637,N_29719,N_26113);
nor U30638 (N_30638,N_25880,N_28992);
nor U30639 (N_30639,N_26941,N_29892);
nor U30640 (N_30640,N_26094,N_27226);
nand U30641 (N_30641,N_29041,N_27258);
xnor U30642 (N_30642,N_25134,N_25707);
xor U30643 (N_30643,N_28295,N_28041);
xor U30644 (N_30644,N_29240,N_26133);
and U30645 (N_30645,N_25132,N_27103);
nor U30646 (N_30646,N_26011,N_29870);
or U30647 (N_30647,N_29749,N_27196);
nand U30648 (N_30648,N_25062,N_29331);
nand U30649 (N_30649,N_26778,N_29655);
xnor U30650 (N_30650,N_26009,N_27455);
nand U30651 (N_30651,N_26789,N_29062);
or U30652 (N_30652,N_29709,N_26891);
xnor U30653 (N_30653,N_27567,N_27416);
and U30654 (N_30654,N_25269,N_28333);
xnor U30655 (N_30655,N_29934,N_26245);
and U30656 (N_30656,N_26123,N_27166);
or U30657 (N_30657,N_29610,N_28810);
or U30658 (N_30658,N_27507,N_29508);
and U30659 (N_30659,N_28445,N_28247);
nand U30660 (N_30660,N_27064,N_27403);
nand U30661 (N_30661,N_29345,N_28605);
and U30662 (N_30662,N_28289,N_28050);
and U30663 (N_30663,N_28245,N_29103);
or U30664 (N_30664,N_25048,N_29044);
or U30665 (N_30665,N_25280,N_28174);
xnor U30666 (N_30666,N_27976,N_29942);
xnor U30667 (N_30667,N_25638,N_29500);
nor U30668 (N_30668,N_27098,N_28974);
and U30669 (N_30669,N_27115,N_29160);
xnor U30670 (N_30670,N_28923,N_26810);
xor U30671 (N_30671,N_29040,N_29141);
nand U30672 (N_30672,N_27825,N_25740);
or U30673 (N_30673,N_29980,N_29657);
and U30674 (N_30674,N_28916,N_26509);
xor U30675 (N_30675,N_27420,N_29656);
and U30676 (N_30676,N_27096,N_27802);
xnor U30677 (N_30677,N_28230,N_26881);
and U30678 (N_30678,N_28768,N_27311);
and U30679 (N_30679,N_26417,N_27313);
nor U30680 (N_30680,N_25804,N_27002);
and U30681 (N_30681,N_27778,N_27578);
xor U30682 (N_30682,N_25986,N_27528);
nand U30683 (N_30683,N_29125,N_26666);
or U30684 (N_30684,N_27452,N_29180);
xor U30685 (N_30685,N_28997,N_28178);
xnor U30686 (N_30686,N_27419,N_29540);
and U30687 (N_30687,N_27040,N_28914);
and U30688 (N_30688,N_26263,N_29444);
nor U30689 (N_30689,N_27478,N_25068);
nand U30690 (N_30690,N_29603,N_26671);
nor U30691 (N_30691,N_29314,N_28481);
nor U30692 (N_30692,N_27559,N_25230);
xor U30693 (N_30693,N_25498,N_28700);
nand U30694 (N_30694,N_25987,N_25892);
or U30695 (N_30695,N_29638,N_28457);
and U30696 (N_30696,N_26953,N_25354);
nor U30697 (N_30697,N_27943,N_29896);
nand U30698 (N_30698,N_26120,N_29938);
xor U30699 (N_30699,N_27558,N_29431);
or U30700 (N_30700,N_26668,N_28968);
and U30701 (N_30701,N_27842,N_27820);
xor U30702 (N_30702,N_27431,N_25655);
xnor U30703 (N_30703,N_29265,N_28640);
xnor U30704 (N_30704,N_26352,N_25410);
nand U30705 (N_30705,N_26145,N_26109);
nand U30706 (N_30706,N_25454,N_26672);
xor U30707 (N_30707,N_27433,N_26657);
or U30708 (N_30708,N_29253,N_25842);
and U30709 (N_30709,N_27328,N_29901);
nor U30710 (N_30710,N_26121,N_29005);
nor U30711 (N_30711,N_28209,N_25080);
and U30712 (N_30712,N_28422,N_29970);
or U30713 (N_30713,N_27369,N_25693);
xor U30714 (N_30714,N_26441,N_27585);
nor U30715 (N_30715,N_27801,N_29352);
and U30716 (N_30716,N_27245,N_28092);
or U30717 (N_30717,N_29242,N_26715);
nand U30718 (N_30718,N_27468,N_26954);
nand U30719 (N_30719,N_27016,N_25078);
and U30720 (N_30720,N_26698,N_29279);
xnor U30721 (N_30721,N_25794,N_26630);
nor U30722 (N_30722,N_28764,N_25070);
or U30723 (N_30723,N_27832,N_26108);
or U30724 (N_30724,N_27168,N_27444);
nand U30725 (N_30725,N_27786,N_29480);
xnor U30726 (N_30726,N_25646,N_28727);
nand U30727 (N_30727,N_26753,N_28707);
and U30728 (N_30728,N_29790,N_26342);
nand U30729 (N_30729,N_26877,N_25192);
nand U30730 (N_30730,N_25159,N_26198);
or U30731 (N_30731,N_25492,N_25969);
and U30732 (N_30732,N_27726,N_27790);
nand U30733 (N_30733,N_26725,N_28679);
and U30734 (N_30734,N_29423,N_27545);
and U30735 (N_30735,N_25739,N_27864);
xor U30736 (N_30736,N_29278,N_27134);
nand U30737 (N_30737,N_27738,N_25381);
and U30738 (N_30738,N_27879,N_28401);
and U30739 (N_30739,N_28775,N_28115);
nor U30740 (N_30740,N_28877,N_29750);
xnor U30741 (N_30741,N_25011,N_25164);
nor U30742 (N_30742,N_28031,N_26272);
nand U30743 (N_30743,N_28982,N_28663);
and U30744 (N_30744,N_26052,N_29665);
xor U30745 (N_30745,N_29815,N_25985);
or U30746 (N_30746,N_29292,N_29561);
nand U30747 (N_30747,N_28439,N_27342);
and U30748 (N_30748,N_26606,N_26691);
or U30749 (N_30749,N_26411,N_25600);
xor U30750 (N_30750,N_29025,N_25201);
or U30751 (N_30751,N_26476,N_27249);
nand U30752 (N_30752,N_29215,N_28008);
and U30753 (N_30753,N_25522,N_29395);
or U30754 (N_30754,N_25013,N_25826);
nand U30755 (N_30755,N_29645,N_26231);
xnor U30756 (N_30756,N_29625,N_28643);
xor U30757 (N_30757,N_29763,N_27843);
nor U30758 (N_30758,N_28550,N_27448);
or U30759 (N_30759,N_29958,N_28170);
xnor U30760 (N_30760,N_29700,N_29123);
nand U30761 (N_30761,N_27732,N_27072);
and U30762 (N_30762,N_27978,N_29619);
nor U30763 (N_30763,N_29971,N_29776);
nand U30764 (N_30764,N_28054,N_26593);
nor U30765 (N_30765,N_25605,N_28695);
nor U30766 (N_30766,N_25855,N_28343);
nand U30767 (N_30767,N_27728,N_29847);
nand U30768 (N_30768,N_27650,N_29631);
xor U30769 (N_30769,N_28475,N_29357);
xor U30770 (N_30770,N_27681,N_29823);
or U30771 (N_30771,N_26619,N_26430);
or U30772 (N_30772,N_27376,N_26043);
xor U30773 (N_30773,N_26653,N_26389);
nor U30774 (N_30774,N_27462,N_27479);
nand U30775 (N_30775,N_25622,N_29124);
nor U30776 (N_30776,N_26350,N_26550);
and U30777 (N_30777,N_29159,N_28282);
xor U30778 (N_30778,N_25196,N_26743);
and U30779 (N_30779,N_26740,N_29562);
nor U30780 (N_30780,N_26354,N_28590);
xnor U30781 (N_30781,N_29997,N_26499);
and U30782 (N_30782,N_25194,N_29291);
nand U30783 (N_30783,N_25543,N_28977);
and U30784 (N_30784,N_25968,N_25947);
or U30785 (N_30785,N_29982,N_25422);
and U30786 (N_30786,N_29623,N_26076);
xnor U30787 (N_30787,N_26717,N_25750);
xor U30788 (N_30788,N_27138,N_26211);
nand U30789 (N_30789,N_29518,N_29398);
nand U30790 (N_30790,N_28753,N_29118);
xor U30791 (N_30791,N_28833,N_25839);
nand U30792 (N_30792,N_26021,N_26017);
nand U30793 (N_30793,N_25697,N_27992);
or U30794 (N_30794,N_28645,N_28278);
xnor U30795 (N_30795,N_28892,N_27903);
nand U30796 (N_30796,N_25051,N_25233);
or U30797 (N_30797,N_28946,N_26620);
nand U30798 (N_30798,N_29429,N_28509);
and U30799 (N_30799,N_27619,N_28301);
xor U30800 (N_30800,N_27690,N_25731);
nand U30801 (N_30801,N_28741,N_25109);
or U30802 (N_30802,N_27915,N_27355);
xnor U30803 (N_30803,N_29006,N_29405);
or U30804 (N_30804,N_26372,N_28664);
and U30805 (N_30805,N_26003,N_26829);
xnor U30806 (N_30806,N_25806,N_27137);
nor U30807 (N_30807,N_29023,N_29649);
nor U30808 (N_30808,N_27099,N_25936);
or U30809 (N_30809,N_25787,N_29397);
or U30810 (N_30810,N_26662,N_26335);
xor U30811 (N_30811,N_29139,N_26187);
nand U30812 (N_30812,N_28778,N_27715);
xor U30813 (N_30813,N_29846,N_25617);
nand U30814 (N_30814,N_26227,N_26149);
nand U30815 (N_30815,N_25714,N_29351);
or U30816 (N_30816,N_27540,N_28379);
or U30817 (N_30817,N_25162,N_26338);
nor U30818 (N_30818,N_26247,N_28861);
or U30819 (N_30819,N_27442,N_25733);
xnor U30820 (N_30820,N_26275,N_25942);
or U30821 (N_30821,N_27722,N_28114);
xnor U30822 (N_30822,N_29926,N_26839);
and U30823 (N_30823,N_27413,N_29542);
nand U30824 (N_30824,N_25821,N_27206);
or U30825 (N_30825,N_25741,N_29043);
and U30826 (N_30826,N_28299,N_27125);
nand U30827 (N_30827,N_27921,N_27008);
or U30828 (N_30828,N_26085,N_27371);
or U30829 (N_30829,N_29246,N_29268);
xnor U30830 (N_30830,N_25105,N_26138);
xor U30831 (N_30831,N_29195,N_28241);
nor U30832 (N_30832,N_26569,N_25033);
or U30833 (N_30833,N_25208,N_29181);
nand U30834 (N_30834,N_29213,N_27617);
or U30835 (N_30835,N_28416,N_27107);
nand U30836 (N_30836,N_25304,N_25868);
and U30837 (N_30837,N_26910,N_28093);
or U30838 (N_30838,N_25290,N_29372);
and U30839 (N_30839,N_26368,N_29698);
and U30840 (N_30840,N_26987,N_28133);
nor U30841 (N_30841,N_28856,N_28161);
xnor U30842 (N_30842,N_27876,N_29525);
nor U30843 (N_30843,N_26206,N_26562);
and U30844 (N_30844,N_27269,N_26540);
xnor U30845 (N_30845,N_25430,N_28536);
nand U30846 (N_30846,N_29391,N_28470);
or U30847 (N_30847,N_26024,N_25994);
nand U30848 (N_30848,N_29818,N_27271);
xor U30849 (N_30849,N_29449,N_26747);
nand U30850 (N_30850,N_28718,N_26314);
nor U30851 (N_30851,N_26093,N_27338);
nand U30852 (N_30852,N_28749,N_29795);
xor U30853 (N_30853,N_29498,N_27084);
xnor U30854 (N_30854,N_29175,N_25609);
or U30855 (N_30855,N_28272,N_25075);
or U30856 (N_30856,N_26885,N_27804);
and U30857 (N_30857,N_27884,N_26475);
xnor U30858 (N_30858,N_25476,N_25604);
nor U30859 (N_30859,N_26035,N_26287);
and U30860 (N_30860,N_25073,N_25464);
xnor U30861 (N_30861,N_25665,N_29729);
nor U30862 (N_30862,N_27701,N_29742);
xor U30863 (N_30863,N_27505,N_28246);
xor U30864 (N_30864,N_29316,N_29559);
nand U30865 (N_30865,N_27608,N_25511);
or U30866 (N_30866,N_26117,N_27159);
and U30867 (N_30867,N_27780,N_29535);
or U30868 (N_30868,N_26836,N_25849);
nor U30869 (N_30869,N_25890,N_28163);
nand U30870 (N_30870,N_29822,N_28229);
nor U30871 (N_30871,N_29009,N_29031);
nand U30872 (N_30872,N_26800,N_27450);
nand U30873 (N_30873,N_26433,N_27458);
or U30874 (N_30874,N_29101,N_25973);
nand U30875 (N_30875,N_27643,N_25500);
nor U30876 (N_30876,N_26410,N_29831);
nor U30877 (N_30877,N_29806,N_27859);
nand U30878 (N_30878,N_26112,N_28400);
xnor U30879 (N_30879,N_28642,N_26689);
nand U30880 (N_30880,N_27027,N_27620);
xor U30881 (N_30881,N_29155,N_26727);
and U30882 (N_30882,N_25347,N_27637);
or U30883 (N_30883,N_26308,N_29913);
and U30884 (N_30884,N_28444,N_29324);
xnor U30885 (N_30885,N_28269,N_27244);
nand U30886 (N_30886,N_26254,N_29537);
nor U30887 (N_30887,N_25627,N_27597);
or U30888 (N_30888,N_25624,N_28399);
xnor U30889 (N_30889,N_29237,N_25928);
nor U30890 (N_30890,N_26784,N_28920);
or U30891 (N_30891,N_28986,N_27933);
nand U30892 (N_30892,N_26584,N_28631);
xnor U30893 (N_30893,N_26622,N_25843);
xnor U30894 (N_30894,N_27340,N_27474);
xor U30895 (N_30895,N_27310,N_29059);
or U30896 (N_30896,N_27955,N_26857);
and U30897 (N_30897,N_28842,N_28970);
xor U30898 (N_30898,N_29212,N_29871);
and U30899 (N_30899,N_29154,N_27772);
or U30900 (N_30900,N_29425,N_25904);
or U30901 (N_30901,N_25852,N_27989);
nor U30902 (N_30902,N_29794,N_27101);
nor U30903 (N_30903,N_26915,N_28244);
xnor U30904 (N_30904,N_28740,N_26179);
and U30905 (N_30905,N_25676,N_27683);
and U30906 (N_30906,N_28325,N_26107);
or U30907 (N_30907,N_28192,N_28102);
nor U30908 (N_30908,N_26018,N_29485);
and U30909 (N_30909,N_25463,N_29532);
xor U30910 (N_30910,N_28971,N_26414);
or U30911 (N_30911,N_28392,N_25171);
or U30912 (N_30912,N_27929,N_28694);
nand U30913 (N_30913,N_27705,N_28944);
and U30914 (N_30914,N_26484,N_25473);
or U30915 (N_30915,N_25586,N_27191);
nor U30916 (N_30916,N_28373,N_28747);
xnor U30917 (N_30917,N_26978,N_26432);
or U30918 (N_30918,N_26849,N_27062);
and U30919 (N_30919,N_27556,N_27211);
and U30920 (N_30920,N_27248,N_25468);
nand U30921 (N_30921,N_26777,N_29303);
xor U30922 (N_30922,N_28649,N_26159);
nor U30923 (N_30923,N_29320,N_28332);
xnor U30924 (N_30924,N_29873,N_27653);
or U30925 (N_30925,N_25176,N_27482);
xnor U30926 (N_30926,N_28567,N_25583);
nand U30927 (N_30927,N_26869,N_25878);
xor U30928 (N_30928,N_27170,N_25404);
nor U30929 (N_30929,N_27289,N_29658);
and U30930 (N_30930,N_25317,N_27586);
xnor U30931 (N_30931,N_25723,N_26745);
nor U30932 (N_30932,N_27058,N_26510);
and U30933 (N_30933,N_25174,N_28555);
nand U30934 (N_30934,N_28693,N_29600);
xnor U30935 (N_30935,N_29301,N_28249);
nand U30936 (N_30936,N_28048,N_28899);
nor U30937 (N_30937,N_27647,N_28350);
or U30938 (N_30938,N_29754,N_29288);
nand U30939 (N_30939,N_29925,N_27185);
xor U30940 (N_30940,N_29371,N_29317);
nand U30941 (N_30941,N_26167,N_26299);
xor U30942 (N_30942,N_27618,N_29672);
nor U30943 (N_30943,N_25553,N_25462);
nor U30944 (N_30944,N_28613,N_27079);
nor U30945 (N_30945,N_25781,N_28488);
or U30946 (N_30946,N_29515,N_25721);
xnor U30947 (N_30947,N_29402,N_26478);
and U30948 (N_30948,N_29668,N_29986);
nand U30949 (N_30949,N_26435,N_25877);
xnor U30950 (N_30950,N_28168,N_27901);
and U30951 (N_30951,N_28397,N_25145);
nor U30952 (N_30952,N_27612,N_28184);
and U30953 (N_30953,N_29477,N_28433);
xor U30954 (N_30954,N_26992,N_26775);
and U30955 (N_30955,N_27055,N_29354);
nand U30956 (N_30956,N_29337,N_25938);
nand U30957 (N_30957,N_25933,N_26576);
and U30958 (N_30958,N_29520,N_27405);
and U30959 (N_30959,N_28449,N_28105);
nor U30960 (N_30960,N_25146,N_26022);
and U30961 (N_30961,N_25434,N_27373);
nand U30962 (N_30962,N_25303,N_27925);
nand U30963 (N_30963,N_28290,N_26664);
nand U30964 (N_30964,N_29864,N_28474);
or U30965 (N_30965,N_28530,N_27295);
nand U30966 (N_30966,N_28673,N_28225);
and U30967 (N_30967,N_26912,N_27406);
xor U30968 (N_30968,N_25970,N_28144);
nand U30969 (N_30969,N_25035,N_27404);
or U30970 (N_30970,N_29568,N_29081);
or U30971 (N_30971,N_29621,N_26241);
xor U30972 (N_30972,N_28402,N_26032);
nor U30973 (N_30973,N_26917,N_26843);
and U30974 (N_30974,N_25957,N_27380);
xnor U30975 (N_30975,N_25632,N_25393);
and U30976 (N_30976,N_25548,N_28213);
nand U30977 (N_30977,N_25546,N_29243);
and U30978 (N_30978,N_26976,N_29432);
nand U30979 (N_30979,N_25281,N_25486);
nor U30980 (N_30980,N_26618,N_25019);
nor U30981 (N_30981,N_29961,N_28142);
or U30982 (N_30982,N_25438,N_29929);
or U30983 (N_30983,N_27731,N_29085);
nand U30984 (N_30984,N_29902,N_25744);
nand U30985 (N_30985,N_29960,N_27741);
nor U30986 (N_30986,N_26772,N_25472);
nand U30987 (N_30987,N_28396,N_27024);
xor U30988 (N_30988,N_27909,N_27109);
nand U30989 (N_30989,N_25989,N_29065);
nand U30990 (N_30990,N_29617,N_27747);
xnor U30991 (N_30991,N_28014,N_28650);
or U30992 (N_30992,N_27327,N_28964);
nand U30993 (N_30993,N_25394,N_26136);
and U30994 (N_30994,N_29602,N_28621);
xnor U30995 (N_30995,N_26984,N_26421);
xor U30996 (N_30996,N_25792,N_27595);
and U30997 (N_30997,N_27863,N_27337);
nor U30998 (N_30998,N_27106,N_26453);
and U30999 (N_30999,N_28958,N_25926);
nor U31000 (N_31000,N_29434,N_25751);
and U31001 (N_31001,N_28662,N_29652);
nand U31002 (N_31002,N_28836,N_28542);
and U31003 (N_31003,N_25474,N_25823);
xor U31004 (N_31004,N_26472,N_29283);
nor U31005 (N_31005,N_25223,N_25310);
nor U31006 (N_31006,N_29406,N_26756);
nor U31007 (N_31007,N_26015,N_25610);
and U31008 (N_31008,N_25578,N_26621);
or U31009 (N_31009,N_29055,N_25929);
and U31010 (N_31010,N_25738,N_27838);
and U31011 (N_31011,N_28564,N_25962);
nor U31012 (N_31012,N_28099,N_27562);
nand U31013 (N_31013,N_29696,N_25867);
nor U31014 (N_31014,N_26615,N_25426);
and U31015 (N_31015,N_25593,N_29570);
nand U31016 (N_31016,N_29708,N_25944);
nand U31017 (N_31017,N_25545,N_28595);
and U31018 (N_31018,N_25931,N_29001);
or U31019 (N_31019,N_27830,N_25491);
nand U31020 (N_31020,N_28816,N_29678);
and U31021 (N_31021,N_28306,N_28936);
nor U31022 (N_31022,N_29207,N_28434);
or U31023 (N_31023,N_27993,N_29736);
and U31024 (N_31024,N_26674,N_29930);
nand U31025 (N_31025,N_28648,N_25427);
and U31026 (N_31026,N_29104,N_28283);
xnor U31027 (N_31027,N_26212,N_25871);
or U31028 (N_31028,N_28711,N_26693);
or U31029 (N_31029,N_25306,N_26633);
nor U31030 (N_31030,N_27816,N_27858);
nor U31031 (N_31031,N_27671,N_27749);
xnor U31032 (N_31032,N_29861,N_28275);
xor U31033 (N_31033,N_29860,N_25705);
nor U31034 (N_31034,N_27640,N_29470);
and U31035 (N_31035,N_25623,N_28149);
or U31036 (N_31036,N_25017,N_28521);
and U31037 (N_31037,N_29882,N_25816);
xnor U31038 (N_31038,N_26364,N_29147);
nand U31039 (N_31039,N_26063,N_27878);
nand U31040 (N_31040,N_27285,N_26517);
nor U31041 (N_31041,N_29740,N_28632);
and U31042 (N_31042,N_25554,N_26282);
xnor U31043 (N_31043,N_29057,N_28034);
nor U31044 (N_31044,N_29546,N_25152);
and U31045 (N_31045,N_28883,N_28582);
nand U31046 (N_31046,N_25796,N_28552);
nand U31047 (N_31047,N_27672,N_27253);
or U31048 (N_31048,N_29013,N_26556);
xnor U31049 (N_31049,N_25585,N_27086);
nor U31050 (N_31050,N_25050,N_29185);
and U31051 (N_31051,N_28431,N_29862);
or U31052 (N_31052,N_28208,N_27622);
and U31053 (N_31053,N_28364,N_27771);
nor U31054 (N_31054,N_27437,N_26050);
nor U31055 (N_31055,N_27609,N_26528);
nand U31056 (N_31056,N_29747,N_29379);
nor U31057 (N_31057,N_29403,N_25641);
nand U31058 (N_31058,N_26859,N_28478);
xor U31059 (N_31059,N_28467,N_26716);
xnor U31060 (N_31060,N_25266,N_29721);
and U31061 (N_31061,N_25418,N_26705);
xor U31062 (N_31062,N_26382,N_26695);
or U31063 (N_31063,N_28169,N_25683);
nor U31064 (N_31064,N_25507,N_29654);
or U31065 (N_31065,N_28814,N_29918);
or U31066 (N_31066,N_27350,N_27944);
xnor U31067 (N_31067,N_29575,N_28500);
or U31068 (N_31068,N_25467,N_26385);
or U31069 (N_31069,N_25211,N_25302);
nor U31070 (N_31070,N_26491,N_26266);
or U31071 (N_31071,N_25590,N_29202);
xnor U31072 (N_31072,N_26862,N_27856);
and U31073 (N_31073,N_29365,N_29825);
nor U31074 (N_31074,N_28925,N_27708);
nand U31075 (N_31075,N_28140,N_26949);
and U31076 (N_31076,N_26788,N_28375);
nand U31077 (N_31077,N_27013,N_25975);
and U31078 (N_31078,N_25997,N_27628);
and U31079 (N_31079,N_28339,N_26386);
nor U31080 (N_31080,N_29000,N_26363);
and U31081 (N_31081,N_25766,N_27547);
and U31082 (N_31082,N_28499,N_27704);
nand U31083 (N_31083,N_27979,N_29193);
nor U31084 (N_31084,N_28322,N_27020);
or U31085 (N_31085,N_26137,N_29226);
and U31086 (N_31086,N_28395,N_27228);
nor U31087 (N_31087,N_27347,N_25165);
nor U31088 (N_31088,N_25903,N_25424);
xor U31089 (N_31089,N_26071,N_26682);
xor U31090 (N_31090,N_28705,N_26738);
and U31091 (N_31091,N_29131,N_27221);
nor U31092 (N_31092,N_28038,N_27833);
or U31093 (N_31093,N_25345,N_27292);
nor U31094 (N_31094,N_28865,N_29108);
and U31095 (N_31095,N_25330,N_26895);
or U31096 (N_31096,N_27691,N_28569);
nand U31097 (N_31097,N_25649,N_27286);
nor U31098 (N_31098,N_29990,N_28682);
nand U31099 (N_31099,N_27641,N_26945);
nand U31100 (N_31100,N_27454,N_28458);
xor U31101 (N_31101,N_29380,N_29735);
nor U31102 (N_31102,N_25710,N_29730);
or U31103 (N_31103,N_27677,N_29135);
or U31104 (N_31104,N_28255,N_26783);
nand U31105 (N_31105,N_26861,N_25071);
or U31106 (N_31106,N_27201,N_28455);
nand U31107 (N_31107,N_25983,N_26316);
and U31108 (N_31108,N_28335,N_27813);
xnor U31109 (N_31109,N_28503,N_29106);
or U31110 (N_31110,N_26257,N_26223);
xnor U31111 (N_31111,N_28391,N_25180);
nand U31112 (N_31112,N_29594,N_25572);
xnor U31113 (N_31113,N_27698,N_26812);
and U31114 (N_31114,N_28723,N_27808);
nor U31115 (N_31115,N_25131,N_29755);
or U31116 (N_31116,N_27767,N_27669);
or U31117 (N_31117,N_26201,N_28506);
nand U31118 (N_31118,N_28644,N_29886);
xnor U31119 (N_31119,N_28888,N_26557);
or U31120 (N_31120,N_27893,N_25689);
nand U31121 (N_31121,N_28737,N_29359);
and U31122 (N_31122,N_25038,N_26796);
xor U31123 (N_31123,N_28622,N_28021);
nor U31124 (N_31124,N_29923,N_27088);
xnor U31125 (N_31125,N_29038,N_25760);
nand U31126 (N_31126,N_29121,N_27069);
or U31127 (N_31127,N_25090,N_28994);
nor U31128 (N_31128,N_29366,N_26425);
or U31129 (N_31129,N_25595,N_25267);
xnor U31130 (N_31130,N_27385,N_29084);
and U31131 (N_31131,N_25709,N_27139);
or U31132 (N_31132,N_29739,N_28469);
xnor U31133 (N_31133,N_26731,N_28781);
or U31134 (N_31134,N_27639,N_29536);
nor U31135 (N_31135,N_28132,N_26887);
nand U31136 (N_31136,N_28878,N_29944);
xnor U31137 (N_31137,N_27145,N_26156);
nor U31138 (N_31138,N_26111,N_28334);
nand U31139 (N_31139,N_26378,N_29574);
nor U31140 (N_31140,N_27958,N_28911);
and U31141 (N_31141,N_29648,N_28112);
xor U31142 (N_31142,N_27865,N_28750);
nor U31143 (N_31143,N_26720,N_28435);
nor U31144 (N_31144,N_26900,N_25025);
and U31145 (N_31145,N_27320,N_27822);
and U31146 (N_31146,N_25607,N_25582);
and U31147 (N_31147,N_27081,N_26205);
and U31148 (N_31148,N_27784,N_28838);
xor U31149 (N_31149,N_27321,N_27663);
and U31150 (N_31150,N_29011,N_27553);
nor U31151 (N_31151,N_28831,N_29775);
or U31152 (N_31152,N_28293,N_28529);
xnor U31153 (N_31153,N_28976,N_26237);
nor U31154 (N_31154,N_28687,N_25547);
or U31155 (N_31155,N_28684,N_27718);
nand U31156 (N_31156,N_25773,N_25574);
nor U31157 (N_31157,N_25977,N_29341);
or U31158 (N_31158,N_26938,N_29289);
and U31159 (N_31159,N_26309,N_26604);
or U31160 (N_31160,N_26991,N_27393);
and U31161 (N_31161,N_28191,N_26409);
or U31162 (N_31162,N_27141,N_26914);
xor U31163 (N_31163,N_26141,N_28575);
or U31164 (N_31164,N_27235,N_26587);
xnor U31165 (N_31165,N_26443,N_28658);
nand U31166 (N_31166,N_29909,N_27885);
nand U31167 (N_31167,N_29233,N_26281);
xnor U31168 (N_31168,N_27555,N_27811);
or U31169 (N_31169,N_25135,N_25798);
xnor U31170 (N_31170,N_26985,N_26981);
nand U31171 (N_31171,N_25487,N_26955);
xnor U31172 (N_31172,N_25367,N_26426);
nand U31173 (N_31173,N_27809,N_26489);
and U31174 (N_31174,N_27023,N_25112);
nand U31175 (N_31175,N_25771,N_29109);
xor U31176 (N_31176,N_29967,N_26326);
or U31177 (N_31177,N_26060,N_28843);
xnor U31178 (N_31178,N_28263,N_26344);
and U31179 (N_31179,N_28234,N_26508);
and U31180 (N_31180,N_28374,N_25270);
and U31181 (N_31181,N_28889,N_27242);
and U31182 (N_31182,N_26190,N_27119);
or U31183 (N_31183,N_29447,N_26469);
and U31184 (N_31184,N_28367,N_27481);
or U31185 (N_31185,N_27896,N_25198);
xor U31186 (N_31186,N_26799,N_29482);
xnor U31187 (N_31187,N_26087,N_28614);
nand U31188 (N_31188,N_29981,N_25119);
nor U31189 (N_31189,N_27673,N_26166);
nor U31190 (N_31190,N_29582,N_25735);
and U31191 (N_31191,N_26442,N_25136);
nand U31192 (N_31192,N_26640,N_28821);
nand U31193 (N_31193,N_25836,N_27358);
nor U31194 (N_31194,N_25900,N_28022);
nand U31195 (N_31195,N_26858,N_27232);
xor U31196 (N_31196,N_28096,N_26280);
nand U31197 (N_31197,N_27695,N_29801);
nor U31198 (N_31198,N_28743,N_25485);
and U31199 (N_31199,N_26627,N_28820);
and U31200 (N_31200,N_28459,N_28734);
or U31201 (N_31201,N_27415,N_25995);
xnor U31202 (N_31202,N_25390,N_27829);
nor U31203 (N_31203,N_27208,N_28651);
xnor U31204 (N_31204,N_26901,N_25848);
and U31205 (N_31205,N_29601,N_27233);
or U31206 (N_31206,N_27888,N_29516);
xnor U31207 (N_31207,N_26296,N_26312);
or U31208 (N_31208,N_25291,N_27998);
and U31209 (N_31209,N_26367,N_28237);
xnor U31210 (N_31210,N_25274,N_27742);
nand U31211 (N_31211,N_29461,N_29489);
nor U31212 (N_31212,N_27623,N_28011);
and U31213 (N_31213,N_28205,N_25854);
or U31214 (N_31214,N_28016,N_29953);
or U31215 (N_31215,N_28933,N_25392);
and U31216 (N_31216,N_26958,N_27987);
nor U31217 (N_31217,N_28867,N_28410);
nand U31218 (N_31218,N_25490,N_25862);
and U31219 (N_31219,N_26034,N_27076);
nand U31220 (N_31220,N_27575,N_28919);
nand U31221 (N_31221,N_26890,N_28421);
and U31222 (N_31222,N_25300,N_26652);
xnor U31223 (N_31223,N_26608,N_29179);
nor U31224 (N_31224,N_29070,N_29414);
and U31225 (N_31225,N_28763,N_29462);
nand U31226 (N_31226,N_29010,N_26128);
xor U31227 (N_31227,N_27839,N_25681);
and U31228 (N_31228,N_29433,N_25057);
xnor U31229 (N_31229,N_28915,N_28046);
nand U31230 (N_31230,N_28064,N_25190);
nand U31231 (N_31231,N_29445,N_26959);
nand U31232 (N_31232,N_28125,N_29270);
or U31233 (N_31233,N_29674,N_28490);
and U31234 (N_31234,N_25772,N_28854);
xnor U31235 (N_31235,N_25373,N_26993);
xor U31236 (N_31236,N_25742,N_26828);
xnor U31237 (N_31237,N_29329,N_27535);
xnor U31238 (N_31238,N_29807,N_28951);
and U31239 (N_31239,N_26651,N_28424);
or U31240 (N_31240,N_25111,N_27309);
nor U31241 (N_31241,N_25980,N_25085);
nor U31242 (N_31242,N_26948,N_27220);
xnor U31243 (N_31243,N_25530,N_27714);
or U31244 (N_31244,N_25858,N_28779);
and U31245 (N_31245,N_29572,N_25830);
nand U31246 (N_31246,N_28755,N_26147);
xnor U31247 (N_31247,N_25449,N_28044);
and U31248 (N_31248,N_25251,N_26962);
or U31249 (N_31249,N_29710,N_29699);
nand U31250 (N_31250,N_25955,N_25990);
or U31251 (N_31251,N_29800,N_26837);
and U31252 (N_31252,N_27872,N_26580);
and U31253 (N_31253,N_26848,N_29382);
nor U31254 (N_31254,N_25722,N_25613);
or U31255 (N_31255,N_29496,N_28000);
nand U31256 (N_31256,N_29164,N_25047);
xnor U31257 (N_31257,N_29420,N_26534);
nand U31258 (N_31258,N_27750,N_28215);
nor U31259 (N_31259,N_26801,N_25431);
nand U31260 (N_31260,N_25036,N_29895);
nand U31261 (N_31261,N_25206,N_27065);
xnor U31262 (N_31262,N_28930,N_26219);
or U31263 (N_31263,N_25370,N_26083);
or U31264 (N_31264,N_25264,N_29858);
nor U31265 (N_31265,N_29693,N_28572);
and U31266 (N_31266,N_28300,N_29326);
or U31267 (N_31267,N_29881,N_28260);
or U31268 (N_31268,N_28538,N_26973);
and U31269 (N_31269,N_28491,N_27290);
nand U31270 (N_31270,N_25452,N_26157);
nand U31271 (N_31271,N_29148,N_29962);
and U31272 (N_31272,N_29143,N_27264);
nor U31273 (N_31273,N_25436,N_29191);
nand U31274 (N_31274,N_26541,N_25402);
or U31275 (N_31275,N_29745,N_26676);
nand U31276 (N_31276,N_27378,N_25121);
xor U31277 (N_31277,N_28493,N_28403);
nor U31278 (N_31278,N_26286,N_26625);
and U31279 (N_31279,N_28104,N_26629);
and U31280 (N_31280,N_25749,N_28336);
xor U31281 (N_31281,N_27093,N_28806);
and U31282 (N_31282,N_26170,N_27449);
xor U31283 (N_31283,N_27770,N_29517);
xnor U31284 (N_31284,N_27797,N_25029);
nand U31285 (N_31285,N_25952,N_25361);
nand U31286 (N_31286,N_28043,N_28187);
xor U31287 (N_31287,N_26178,N_26464);
nand U31288 (N_31288,N_29162,N_28688);
or U31289 (N_31289,N_28456,N_26690);
xor U31290 (N_31290,N_27372,N_25469);
or U31291 (N_31291,N_27527,N_28641);
nand U31292 (N_31292,N_26304,N_29244);
nor U31293 (N_31293,N_25375,N_26185);
or U31294 (N_31294,N_26537,N_26872);
and U31295 (N_31295,N_26931,N_25807);
nor U31296 (N_31296,N_27887,N_28156);
xor U31297 (N_31297,N_27959,N_26124);
or U31298 (N_31298,N_29501,N_29340);
and U31299 (N_31299,N_25455,N_26904);
nand U31300 (N_31300,N_29021,N_26548);
or U31301 (N_31301,N_28725,N_27531);
nor U31302 (N_31302,N_26249,N_26171);
and U31303 (N_31303,N_27260,N_29008);
or U31304 (N_31304,N_27306,N_26379);
xnor U31305 (N_31305,N_27256,N_25795);
and U31306 (N_31306,N_29234,N_27487);
or U31307 (N_31307,N_28113,N_29723);
nor U31308 (N_31308,N_27283,N_25276);
nand U31309 (N_31309,N_25588,N_27356);
and U31310 (N_31310,N_29047,N_26832);
and U31311 (N_31311,N_28303,N_26700);
nor U31312 (N_31312,N_28007,N_27217);
nor U31313 (N_31313,N_29306,N_26903);
nor U31314 (N_31314,N_25202,N_25881);
and U31315 (N_31315,N_28036,N_27060);
nand U31316 (N_31316,N_25297,N_27973);
or U31317 (N_31317,N_28307,N_26099);
nand U31318 (N_31318,N_25183,N_28261);
xor U31319 (N_31319,N_29119,N_25976);
nand U31320 (N_31320,N_25077,N_27542);
or U31321 (N_31321,N_28313,N_25780);
and U31322 (N_31322,N_26101,N_25688);
nor U31323 (N_31323,N_27634,N_27067);
and U31324 (N_31324,N_25690,N_27200);
and U31325 (N_31325,N_29639,N_29022);
xor U31326 (N_31326,N_26422,N_26875);
nand U31327 (N_31327,N_26758,N_25179);
or U31328 (N_31328,N_28338,N_25277);
or U31329 (N_31329,N_26547,N_29644);
or U31330 (N_31330,N_25213,N_26097);
nand U31331 (N_31331,N_25369,N_26183);
or U31332 (N_31332,N_26986,N_28752);
and U31333 (N_31333,N_26346,N_26028);
or U31334 (N_31334,N_26963,N_27520);
xnor U31335 (N_31335,N_27656,N_25007);
nand U31336 (N_31336,N_28405,N_27999);
xor U31337 (N_31337,N_27868,N_26511);
and U31338 (N_31338,N_29686,N_28139);
nor U31339 (N_31339,N_28348,N_25817);
nor U31340 (N_31340,N_25000,N_25177);
xnor U31341 (N_31341,N_29883,N_25320);
and U31342 (N_31342,N_27210,N_29894);
xor U31343 (N_31343,N_27710,N_28286);
xor U31344 (N_31344,N_25168,N_26768);
nand U31345 (N_31345,N_28955,N_27129);
xor U31346 (N_31346,N_26110,N_28487);
and U31347 (N_31347,N_26524,N_29731);
nor U31348 (N_31348,N_27499,N_26031);
nand U31349 (N_31349,N_28352,N_29770);
nor U31350 (N_31350,N_26699,N_29545);
xor U31351 (N_31351,N_29707,N_28302);
and U31352 (N_31352,N_28586,N_27974);
or U31353 (N_31353,N_25123,N_28404);
or U31354 (N_31354,N_29943,N_27389);
nand U31355 (N_31355,N_29992,N_26438);
xnor U31356 (N_31356,N_27143,N_25319);
nand U31357 (N_31357,N_25626,N_26373);
or U31358 (N_31358,N_27279,N_28953);
nand U31359 (N_31359,N_26045,N_29704);
nand U31360 (N_31360,N_27194,N_29765);
xnor U31361 (N_31361,N_28264,N_28067);
xnor U31362 (N_31362,N_28111,N_29310);
xor U31363 (N_31363,N_26913,N_26082);
or U31364 (N_31364,N_27764,N_26536);
and U31365 (N_31365,N_29922,N_28460);
nor U31366 (N_31366,N_26611,N_26667);
xnor U31367 (N_31367,N_26259,N_26980);
xnor U31368 (N_31368,N_26483,N_25921);
xnor U31369 (N_31369,N_27755,N_28496);
nand U31370 (N_31370,N_26680,N_25451);
and U31371 (N_31371,N_27029,N_28376);
nand U31372 (N_31372,N_28869,N_28308);
nor U31373 (N_31373,N_27692,N_28094);
nand U31374 (N_31374,N_27849,N_27118);
xor U31375 (N_31375,N_27543,N_26105);
nor U31376 (N_31376,N_26678,N_29214);
or U31377 (N_31377,N_27428,N_25301);
nor U31378 (N_31378,N_25371,N_26927);
nand U31379 (N_31379,N_28829,N_29702);
or U31380 (N_31380,N_27765,N_28227);
or U31381 (N_31381,N_26391,N_26010);
and U31382 (N_31382,N_29586,N_25083);
nand U31383 (N_31383,N_29505,N_26243);
and U31384 (N_31384,N_26194,N_27583);
xnor U31385 (N_31385,N_29322,N_28386);
nor U31386 (N_31386,N_27598,N_27172);
nor U31387 (N_31387,N_26635,N_25133);
nor U31388 (N_31388,N_28494,N_27374);
nand U31389 (N_31389,N_29144,N_29390);
nor U31390 (N_31390,N_26403,N_29358);
or U31391 (N_31391,N_25694,N_25906);
xor U31392 (N_31392,N_29308,N_29453);
and U31393 (N_31393,N_25847,N_28020);
nand U31394 (N_31394,N_28666,N_28381);
nand U31395 (N_31395,N_25098,N_26723);
xor U31396 (N_31396,N_26228,N_28647);
or U31397 (N_31397,N_29832,N_29424);
and U31398 (N_31398,N_25318,N_29691);
or U31399 (N_31399,N_29733,N_28240);
xnor U31400 (N_31400,N_29077,N_25242);
nor U31401 (N_31401,N_26773,N_28522);
nor U31402 (N_31402,N_26737,N_29051);
or U31403 (N_31403,N_29087,N_28875);
or U31404 (N_31404,N_29868,N_29640);
xor U31405 (N_31405,N_25420,N_25229);
nand U31406 (N_31406,N_27203,N_25210);
or U31407 (N_31407,N_29875,N_29630);
or U31408 (N_31408,N_27964,N_25712);
or U31409 (N_31409,N_28853,N_25520);
xnor U31410 (N_31410,N_26706,N_27686);
xor U31411 (N_31411,N_28576,N_25074);
and U31412 (N_31412,N_27900,N_26176);
or U31413 (N_31413,N_28868,N_28756);
nor U31414 (N_31414,N_27601,N_26795);
or U31415 (N_31415,N_25053,N_25599);
nor U31416 (N_31416,N_28656,N_27751);
or U31417 (N_31417,N_26533,N_26623);
nand U31418 (N_31418,N_27425,N_26370);
and U31419 (N_31419,N_29095,N_28880);
nor U31420 (N_31420,N_26578,N_25692);
xnor U31421 (N_31421,N_29053,N_29577);
and U31422 (N_31422,N_25060,N_28887);
or U31423 (N_31423,N_29221,N_25184);
nand U31424 (N_31424,N_25673,N_29939);
nand U31425 (N_31425,N_28761,N_29151);
nand U31426 (N_31426,N_26708,N_27716);
xor U31427 (N_31427,N_26571,N_29889);
nor U31428 (N_31428,N_25758,N_29451);
nand U31429 (N_31429,N_25913,N_29897);
or U31430 (N_31430,N_28298,N_25012);
nor U31431 (N_31431,N_26681,N_25005);
and U31432 (N_31432,N_29343,N_29113);
xnor U31433 (N_31433,N_27239,N_27638);
xor U31434 (N_31434,N_27988,N_27204);
nor U31435 (N_31435,N_28483,N_28207);
or U31436 (N_31436,N_29588,N_28762);
xnor U31437 (N_31437,N_25647,N_25894);
or U31438 (N_31438,N_25789,N_26787);
nand U31439 (N_31439,N_25825,N_26643);
nor U31440 (N_31440,N_26470,N_29281);
nor U31441 (N_31441,N_29294,N_26158);
nand U31442 (N_31442,N_28519,N_29903);
or U31443 (N_31443,N_26605,N_26406);
and U31444 (N_31444,N_29061,N_25216);
nand U31445 (N_31445,N_25911,N_25953);
nand U31446 (N_31446,N_29549,N_25389);
or U31447 (N_31447,N_25979,N_28250);
or U31448 (N_31448,N_27004,N_28015);
xnor U31449 (N_31449,N_25512,N_27721);
xnor U31450 (N_31450,N_27333,N_27758);
or U31451 (N_31451,N_25967,N_29646);
or U31452 (N_31452,N_29975,N_25363);
nand U31453 (N_31453,N_25456,N_26648);
xnor U31454 (N_31454,N_27962,N_28130);
and U31455 (N_31455,N_28882,N_28309);
nand U31456 (N_31456,N_28116,N_26989);
or U31457 (N_31457,N_25231,N_27934);
nor U31458 (N_31458,N_25237,N_29900);
nand U31459 (N_31459,N_27779,N_27563);
nand U31460 (N_31460,N_27756,N_29389);
nor U31461 (N_31461,N_29612,N_28691);
xor U31462 (N_31462,N_26526,N_26255);
or U31463 (N_31463,N_28771,N_29259);
and U31464 (N_31464,N_28716,N_29262);
or U31465 (N_31465,N_29753,N_29857);
nor U31466 (N_31466,N_29620,N_26098);
nand U31467 (N_31467,N_25124,N_29276);
nand U31468 (N_31468,N_29661,N_25374);
xor U31469 (N_31469,N_28773,N_26150);
and U31470 (N_31470,N_27823,N_25238);
nand U31471 (N_31471,N_28124,N_26122);
nor U31472 (N_31472,N_29307,N_25250);
and U31473 (N_31473,N_29957,N_29183);
nor U31474 (N_31474,N_29107,N_27078);
nand U31475 (N_31475,N_27982,N_28792);
nor U31476 (N_31476,N_26030,N_27739);
and U31477 (N_31477,N_28874,N_28010);
and U31478 (N_31478,N_28152,N_26591);
nor U31479 (N_31479,N_28126,N_25143);
nor U31480 (N_31480,N_29075,N_27182);
or U31481 (N_31481,N_28776,N_26146);
nor U31482 (N_31482,N_26000,N_29146);
xnor U31483 (N_31483,N_26191,N_25113);
nand U31484 (N_31484,N_26070,N_27251);
nand U31485 (N_31485,N_27480,N_28758);
xor U31486 (N_31486,N_28219,N_25031);
nor U31487 (N_31487,N_25116,N_27591);
nor U31488 (N_31488,N_27703,N_29556);
nand U31489 (N_31489,N_27905,N_29679);
xor U31490 (N_31490,N_29437,N_28956);
or U31491 (N_31491,N_28297,N_28212);
nor U31492 (N_31492,N_27538,N_28876);
xor U31493 (N_31493,N_27766,N_28890);
or U31494 (N_31494,N_27629,N_25745);
nor U31495 (N_31495,N_28623,N_28147);
nor U31496 (N_31496,N_25099,N_28089);
nor U31497 (N_31497,N_28073,N_29427);
or U31498 (N_31498,N_27465,N_28157);
xor U31499 (N_31499,N_25246,N_28973);
and U31500 (N_31500,N_28510,N_28389);
and U31501 (N_31501,N_29983,N_28787);
or U31502 (N_31502,N_27399,N_26846);
xnor U31503 (N_31503,N_25419,N_26741);
or U31504 (N_31504,N_25212,N_26218);
and U31505 (N_31505,N_27094,N_27353);
xnor U31506 (N_31506,N_25092,N_28107);
xor U31507 (N_31507,N_28009,N_26256);
or U31508 (N_31508,N_29252,N_25937);
and U31509 (N_31509,N_29802,N_27560);
nor U31510 (N_31510,N_26479,N_27343);
xor U31511 (N_31511,N_26020,N_29483);
xnor U31512 (N_31512,N_27506,N_26222);
nor U31513 (N_31513,N_25525,N_25042);
xnor U31514 (N_31514,N_27362,N_26248);
and U31515 (N_31515,N_26059,N_26265);
or U31516 (N_31516,N_26969,N_29030);
and U31517 (N_31517,N_26250,N_29626);
xor U31518 (N_31518,N_27375,N_28917);
or U31519 (N_31519,N_25576,N_25082);
and U31520 (N_31520,N_25899,N_27091);
xnor U31521 (N_31521,N_27579,N_27491);
nor U31522 (N_31522,N_27227,N_25598);
or U31523 (N_31523,N_28164,N_27572);
nor U31524 (N_31524,N_25734,N_26463);
xnor U31525 (N_31525,N_25568,N_25650);
and U31526 (N_31526,N_25564,N_27939);
and U31527 (N_31527,N_25337,N_25897);
nor U31528 (N_31528,N_28579,N_28438);
nand U31529 (N_31529,N_27687,N_29576);
and U31530 (N_31530,N_26104,N_29869);
and U31531 (N_31531,N_25901,N_26193);
xnor U31532 (N_31532,N_25695,N_25272);
nor U31533 (N_31533,N_26752,N_27180);
nor U31534 (N_31534,N_28233,N_25853);
and U31535 (N_31535,N_28937,N_29874);
and U31536 (N_31536,N_29703,N_29068);
xnor U31537 (N_31537,N_29835,N_27009);
xor U31538 (N_31538,N_28819,N_28317);
or U31539 (N_31539,N_28577,N_29893);
nand U31540 (N_31540,N_27776,N_27035);
xor U31541 (N_31541,N_26507,N_26500);
or U31542 (N_31542,N_25108,N_25930);
and U31543 (N_31543,N_26940,N_26340);
xnor U31544 (N_31544,N_28929,N_26732);
nand U31545 (N_31545,N_28587,N_26866);
xnor U31546 (N_31546,N_27984,N_29768);
nand U31547 (N_31547,N_25096,N_26893);
and U31548 (N_31548,N_28040,N_26647);
and U31549 (N_31549,N_29039,N_29230);
xnor U31550 (N_31550,N_25414,N_27630);
or U31551 (N_31551,N_29093,N_28484);
nand U31552 (N_31552,N_29816,N_28685);
and U31553 (N_31553,N_25150,N_27461);
or U31554 (N_31554,N_25833,N_29019);
or U31555 (N_31555,N_28179,N_27412);
and U31556 (N_31556,N_28273,N_28714);
nor U31557 (N_31557,N_28501,N_27162);
nand U31558 (N_31558,N_26457,N_29865);
xor U31559 (N_31559,N_28979,N_27510);
or U31560 (N_31560,N_26383,N_26879);
nand U31561 (N_31561,N_27068,N_28607);
and U31562 (N_31562,N_27401,N_28796);
and U31563 (N_31563,N_25115,N_25360);
and U31564 (N_31564,N_29495,N_29701);
xnor U31565 (N_31565,N_28846,N_29774);
and U31566 (N_31566,N_27521,N_26755);
nor U31567 (N_31567,N_29335,N_27626);
xnor U31568 (N_31568,N_25635,N_28612);
nand U31569 (N_31569,N_29479,N_25537);
or U31570 (N_31570,N_25851,N_26358);
xor U31571 (N_31571,N_29849,N_27223);
and U31572 (N_31572,N_28948,N_29033);
and U31573 (N_31573,N_28699,N_25528);
nand U31574 (N_31574,N_27819,N_25401);
xnor U31575 (N_31575,N_27652,N_25644);
xor U31576 (N_31576,N_26369,N_29613);
xor U31577 (N_31577,N_27469,N_25448);
nand U31578 (N_31578,N_26816,N_26665);
or U31579 (N_31579,N_25107,N_25876);
xnor U31580 (N_31580,N_29977,N_26736);
and U31581 (N_31581,N_27336,N_29797);
or U31582 (N_31582,N_27005,N_26427);
nand U31583 (N_31583,N_25948,N_29828);
or U31584 (N_31584,N_29309,N_25022);
xnor U31585 (N_31585,N_29441,N_25774);
or U31586 (N_31586,N_28941,N_29627);
xor U31587 (N_31587,N_28226,N_28742);
nand U31588 (N_31588,N_25959,N_26572);
xor U31589 (N_31589,N_26581,N_29635);
xnor U31590 (N_31590,N_26454,N_27427);
xor U31591 (N_31591,N_26377,N_29681);
xnor U31592 (N_31592,N_28095,N_29258);
nor U31593 (N_31593,N_25514,N_25063);
nor U31594 (N_31594,N_28137,N_29841);
nand U31595 (N_31595,N_28995,N_28464);
nor U31596 (N_31596,N_26067,N_28733);
and U31597 (N_31597,N_25660,N_25857);
nor U31598 (N_31598,N_29964,N_25364);
nor U31599 (N_31599,N_27387,N_25596);
or U31600 (N_31600,N_28922,N_26774);
or U31601 (N_31601,N_28062,N_25236);
xor U31602 (N_31602,N_29486,N_27922);
xnor U31603 (N_31603,N_29311,N_27827);
nor U31604 (N_31604,N_25800,N_25286);
nand U31605 (N_31605,N_25724,N_27051);
nand U31606 (N_31606,N_27011,N_29845);
and U31607 (N_31607,N_25674,N_25341);
and U31608 (N_31608,N_29743,N_27860);
or U31609 (N_31609,N_28304,N_26956);
and U31610 (N_31610,N_29003,N_26236);
and U31611 (N_31611,N_28841,N_27759);
nand U31612 (N_31612,N_29528,N_25256);
and U31613 (N_31613,N_27331,N_29045);
xnor U31614 (N_31614,N_27549,N_27057);
or U31615 (N_31615,N_27382,N_25220);
and U31616 (N_31616,N_26481,N_26322);
and U31617 (N_31617,N_29374,N_29362);
or U31618 (N_31618,N_27873,N_27960);
nor U31619 (N_31619,N_29837,N_27503);
and U31620 (N_31620,N_25642,N_25916);
or U31621 (N_31621,N_25958,N_25433);
nor U31622 (N_31622,N_25864,N_26197);
and U31623 (N_31623,N_26819,N_28677);
and U31624 (N_31624,N_25120,N_29471);
or U31625 (N_31625,N_27001,N_25283);
xor U31626 (N_31626,N_25197,N_25470);
nand U31627 (N_31627,N_25579,N_27821);
nand U31628 (N_31628,N_26002,N_28667);
xnor U31629 (N_31629,N_29954,N_29788);
and U31630 (N_31630,N_29551,N_28585);
nor U31631 (N_31631,N_27494,N_27544);
nand U31632 (N_31632,N_25506,N_29566);
xor U31633 (N_31633,N_25488,N_29683);
xnor U31634 (N_31634,N_26151,N_25784);
or U31635 (N_31635,N_25207,N_25515);
and U31636 (N_31636,N_25777,N_27891);
or U31637 (N_31637,N_28141,N_29539);
or U31638 (N_31638,N_29282,N_27270);
nand U31639 (N_31639,N_29716,N_26115);
or U31640 (N_31640,N_25822,N_25260);
nor U31641 (N_31641,N_27898,N_26496);
xnor U31642 (N_31642,N_25103,N_25524);
nor U31643 (N_31643,N_29024,N_28069);
and U31644 (N_31644,N_27539,N_26654);
or U31645 (N_31645,N_25923,N_29811);
nand U31646 (N_31646,N_28859,N_27854);
and U31647 (N_31647,N_27590,N_26792);
xor U31648 (N_31648,N_27075,N_26894);
xnor U31649 (N_31649,N_27904,N_26274);
xor U31650 (N_31650,N_25265,N_27152);
nand U31651 (N_31651,N_28242,N_25417);
nand U31652 (N_31652,N_25021,N_28409);
and U31653 (N_31653,N_29706,N_26330);
xnor U31654 (N_31654,N_25346,N_26332);
nand U31655 (N_31655,N_28610,N_28524);
nor U31656 (N_31656,N_27511,N_27390);
or U31657 (N_31657,N_26631,N_27666);
or U31658 (N_31658,N_25387,N_28683);
or U31659 (N_31659,N_27411,N_28277);
xnor U31660 (N_31660,N_29940,N_26401);
xnor U31661 (N_31661,N_28523,N_28947);
xor U31662 (N_31662,N_28512,N_27752);
nor U31663 (N_31663,N_26823,N_28101);
xnor U31664 (N_31664,N_25889,N_25376);
or U31665 (N_31665,N_26075,N_29611);
xnor U31666 (N_31666,N_25328,N_26561);
and U31667 (N_31667,N_28789,N_25358);
or U31668 (N_31668,N_27645,N_25575);
nor U31669 (N_31669,N_29726,N_26860);
xnor U31670 (N_31670,N_27083,N_27906);
nor U31671 (N_31671,N_27036,N_29225);
and U31672 (N_31672,N_28940,N_26431);
xor U31673 (N_31673,N_26543,N_29381);
xnor U31674 (N_31674,N_29080,N_29854);
nor U31675 (N_31675,N_28633,N_27504);
xnor U31676 (N_31676,N_29274,N_25757);
or U31677 (N_31677,N_26776,N_29599);
and U31678 (N_31678,N_28967,N_28657);
and U31679 (N_31679,N_27806,N_28862);
and U31680 (N_31680,N_25759,N_25510);
or U31681 (N_31681,N_28477,N_27649);
or U31682 (N_31682,N_25333,N_29513);
nand U31683 (N_31683,N_26276,N_25446);
nor U31684 (N_31684,N_27205,N_26697);
xor U31685 (N_31685,N_28001,N_25314);
and U31686 (N_31686,N_26942,N_26798);
or U31687 (N_31687,N_25597,N_25344);
and U31688 (N_31688,N_26049,N_29855);
nand U31689 (N_31689,N_27565,N_25732);
nand U31690 (N_31690,N_29378,N_27453);
or U31691 (N_31691,N_28818,N_28584);
xor U31692 (N_31692,N_25730,N_25951);
nor U31693 (N_31693,N_28280,N_26646);
nand U31694 (N_31694,N_27954,N_27963);
nand U31695 (N_31695,N_25440,N_27246);
or U31696 (N_31696,N_29247,N_29587);
or U31697 (N_31697,N_27514,N_29036);
xor U31698 (N_31698,N_26911,N_25895);
nand U31699 (N_31699,N_27616,N_29529);
xnor U31700 (N_31700,N_27709,N_28910);
nand U31701 (N_31701,N_29336,N_29208);
nor U31702 (N_31702,N_25671,N_26357);
nand U31703 (N_31703,N_25812,N_27685);
and U31704 (N_31704,N_25130,N_28571);
or U31705 (N_31705,N_27112,N_27050);
nor U31706 (N_31706,N_26590,N_28287);
nand U31707 (N_31707,N_26418,N_28318);
or U31708 (N_31708,N_27022,N_29115);
or U31709 (N_31709,N_28769,N_26579);
nor U31710 (N_31710,N_26937,N_27869);
xor U31711 (N_31711,N_29409,N_28354);
or U31712 (N_31712,N_27275,N_29328);
nor U31713 (N_31713,N_25235,N_27052);
and U31714 (N_31714,N_25203,N_29079);
xnor U31715 (N_31715,N_28560,N_27783);
nor U31716 (N_31716,N_25802,N_26051);
and U31717 (N_31717,N_28200,N_29712);
nand U31718 (N_31718,N_29178,N_29771);
or U31719 (N_31719,N_25398,N_28407);
xor U31720 (N_31720,N_26095,N_29012);
or U31721 (N_31721,N_28194,N_28202);
and U31722 (N_31722,N_25495,N_27070);
nand U31723 (N_31723,N_29777,N_27568);
nand U31724 (N_31724,N_25629,N_29973);
nor U31725 (N_31725,N_25943,N_29421);
and U31726 (N_31726,N_25966,N_25893);
xor U31727 (N_31727,N_28543,N_26899);
or U31728 (N_31728,N_29280,N_26530);
xnor U31729 (N_31729,N_25258,N_28119);
and U31730 (N_31730,N_28224,N_27828);
nand U31731 (N_31731,N_28989,N_25041);
xnor U31732 (N_31732,N_28398,N_25081);
xor U31733 (N_31733,N_26042,N_27948);
xnor U31734 (N_31734,N_26644,N_29286);
nand U31735 (N_31735,N_29323,N_25055);
nand U31736 (N_31736,N_26850,N_27532);
and U31737 (N_31737,N_25659,N_25919);
or U31738 (N_31738,N_29250,N_28828);
or U31739 (N_31739,N_27658,N_27911);
nor U31740 (N_31740,N_28620,N_29342);
nor U31741 (N_31741,N_27697,N_26944);
nand U31742 (N_31742,N_29117,N_27968);
nand U31743 (N_31743,N_29122,N_26268);
nand U31744 (N_31744,N_29936,N_27850);
or U31745 (N_31745,N_25770,N_27409);
nor U31746 (N_31746,N_27303,N_26450);
and U31747 (N_31747,N_29567,N_29955);
xor U31748 (N_31748,N_25633,N_29132);
or U31749 (N_31749,N_28310,N_25137);
or U31750 (N_31750,N_29475,N_28166);
nand U31751 (N_31751,N_25009,N_27344);
nor U31752 (N_31752,N_25499,N_26506);
and U31753 (N_31753,N_25682,N_29465);
and U31754 (N_31754,N_25069,N_28604);
xnor U31755 (N_31755,N_26610,N_28088);
nand U31756 (N_31756,N_27769,N_26351);
nor U31757 (N_31757,N_28347,N_28056);
nand U31758 (N_31758,N_25118,N_25762);
nand U31759 (N_31759,N_26660,N_27174);
nand U31760 (N_31760,N_28901,N_27627);
nand U31761 (N_31761,N_29367,N_27031);
nor U31762 (N_31762,N_27561,N_27126);
nor U31763 (N_31763,N_29590,N_25799);
nor U31764 (N_31764,N_25706,N_27324);
nand U31765 (N_31765,N_28131,N_28939);
nand U31766 (N_31766,N_28063,N_28807);
and U31767 (N_31767,N_25308,N_27207);
and U31768 (N_31768,N_28185,N_27287);
nand U31769 (N_31769,N_28252,N_28428);
nor U31770 (N_31770,N_25637,N_27899);
nand U31771 (N_31771,N_25850,N_28091);
or U31772 (N_31772,N_27435,N_28188);
or U31773 (N_31773,N_26131,N_26012);
nor U31774 (N_31774,N_27524,N_28346);
xnor U31775 (N_31775,N_26192,N_27363);
or U31776 (N_31776,N_29692,N_28258);
or U31777 (N_31777,N_29789,N_28281);
nor U31778 (N_31778,N_25939,N_28573);
nor U31779 (N_31779,N_29412,N_29677);
nand U31780 (N_31780,N_25072,N_25914);
xor U31781 (N_31781,N_27537,N_25412);
nor U31782 (N_31782,N_28214,N_26331);
nor U31783 (N_31783,N_25831,N_28802);
or U31784 (N_31784,N_29714,N_29738);
nand U31785 (N_31785,N_25971,N_25715);
xor U31786 (N_31786,N_25708,N_27163);
xor U31787 (N_31787,N_27589,N_28411);
nand U31788 (N_31788,N_27880,N_26639);
nand U31789 (N_31789,N_27318,N_27719);
nand U31790 (N_31790,N_28872,N_29099);
or U31791 (N_31791,N_29737,N_28719);
xnor U31792 (N_31792,N_29524,N_28029);
nor U31793 (N_31793,N_27956,N_26826);
nor U31794 (N_31794,N_26294,N_26238);
or U31795 (N_31795,N_28248,N_27457);
or U31796 (N_31796,N_28617,N_26081);
nor U31797 (N_31797,N_25797,N_29218);
xnor U31798 (N_31798,N_29996,N_27803);
xnor U31799 (N_31799,N_26283,N_26302);
nor U31800 (N_31800,N_25570,N_29628);
xnor U31801 (N_31801,N_28972,N_27852);
nor U31802 (N_31802,N_28729,N_25298);
or U31803 (N_31803,N_28931,N_26154);
nand U31804 (N_31804,N_26763,N_27178);
nand U31805 (N_31805,N_27446,N_25227);
xor U31806 (N_31806,N_26066,N_27541);
or U31807 (N_31807,N_26831,N_29353);
or U31808 (N_31808,N_27688,N_26806);
or U31809 (N_31809,N_25061,N_26473);
xnor U31810 (N_31810,N_26039,N_27222);
and U31811 (N_31811,N_27165,N_26482);
and U31812 (N_31812,N_28026,N_28430);
xor U31813 (N_31813,N_26270,N_29297);
or U31814 (N_31814,N_29722,N_29197);
and U31815 (N_31815,N_29650,N_29669);
and U31816 (N_31816,N_25421,N_27587);
or U31817 (N_31817,N_25698,N_29173);
nand U31818 (N_31818,N_29978,N_28966);
or U31819 (N_31819,N_28637,N_27225);
and U31820 (N_31820,N_26876,N_28774);
xnor U31821 (N_31821,N_25827,N_27814);
nand U31822 (N_31822,N_28486,N_29759);
and U31823 (N_31823,N_26878,N_28794);
nand U31824 (N_31824,N_27489,N_26626);
and U31825 (N_31825,N_25640,N_27774);
and U31826 (N_31826,N_27451,N_27950);
and U31827 (N_31827,N_28591,N_28987);
nand U31828 (N_31828,N_29522,N_26902);
nor U31829 (N_31829,N_29633,N_26084);
nor U31830 (N_31830,N_26341,N_27334);
or U31831 (N_31831,N_29067,N_25815);
or U31832 (N_31832,N_26947,N_27493);
nor U31833 (N_31833,N_25519,N_28625);
and U31834 (N_31834,N_27361,N_28540);
xnor U31835 (N_31835,N_29110,N_27102);
or U31836 (N_31836,N_25753,N_27713);
nor U31837 (N_31837,N_26203,N_28636);
and U31838 (N_31838,N_29100,N_27136);
nand U31839 (N_31839,N_26349,N_29127);
nand U31840 (N_31840,N_25643,N_28047);
nor U31841 (N_31841,N_26920,N_27733);
nand U31842 (N_31842,N_29952,N_27846);
xnor U31843 (N_31843,N_26933,N_25189);
nor U31844 (N_31844,N_25332,N_27033);
nand U31845 (N_31845,N_28135,N_26221);
and U31846 (N_31846,N_27644,N_25268);
nor U31847 (N_31847,N_26649,N_27368);
or U31848 (N_31848,N_26058,N_25141);
nand U31849 (N_31849,N_28243,N_27085);
or U31850 (N_31850,N_29597,N_27219);
nor U31851 (N_31851,N_28451,N_25713);
nor U31852 (N_31852,N_29660,N_27041);
xor U31853 (N_31853,N_27748,N_25205);
nand U31854 (N_31854,N_28702,N_29689);
or U31855 (N_31855,N_29204,N_29137);
or U31856 (N_31856,N_25927,N_25675);
nor U31857 (N_31857,N_25809,N_28709);
xnor U31858 (N_31858,N_28146,N_29058);
and U31859 (N_31859,N_27870,N_27254);
nor U31860 (N_31860,N_29670,N_27202);
nand U31861 (N_31861,N_26068,N_27049);
nand U31862 (N_31862,N_27477,N_28697);
xnor U31863 (N_31863,N_28809,N_26863);
or U31864 (N_31864,N_28059,N_25214);
nand U31865 (N_31865,N_27679,N_28090);
nor U31866 (N_31866,N_28611,N_25801);
xnor U31867 (N_31867,N_27074,N_29688);
xnor U31868 (N_31868,N_29299,N_26636);
and U31869 (N_31869,N_26497,N_26559);
nor U31870 (N_31870,N_28159,N_29912);
nor U31871 (N_31871,N_25126,N_28924);
nor U31872 (N_31872,N_26525,N_29999);
xnor U31873 (N_31873,N_27513,N_26415);
nand U31874 (N_31874,N_28900,N_28857);
nor U31875 (N_31875,N_27484,N_27570);
or U31876 (N_31876,N_29032,N_29222);
and U31877 (N_31877,N_28382,N_28950);
or U31878 (N_31878,N_28959,N_28086);
nor U31879 (N_31879,N_29375,N_27573);
nand U31880 (N_31880,N_28639,N_29417);
nor U31881 (N_31881,N_27127,N_25793);
and U31882 (N_31882,N_27164,N_26957);
or U31883 (N_31883,N_28839,N_26729);
nand U31884 (N_31884,N_29910,N_25618);
or U31885 (N_31885,N_25122,N_28427);
and U31886 (N_31886,N_25459,N_28546);
nand U31887 (N_31887,N_29430,N_25001);
nand U31888 (N_31888,N_29325,N_29370);
nand U31889 (N_31889,N_28744,N_25217);
nor U31890 (N_31890,N_27319,N_27108);
xor U31891 (N_31891,N_28898,N_27422);
xor U31892 (N_31892,N_25155,N_27930);
and U31893 (N_31893,N_28121,N_28045);
and U31894 (N_31894,N_28030,N_26495);
nand U31895 (N_31895,N_28027,N_28566);
nand U31896 (N_31896,N_29172,N_26687);
nand U31897 (N_31897,N_26970,N_29376);
nand U31898 (N_31898,N_26502,N_28228);
nand U31899 (N_31899,N_29016,N_29052);
and U31900 (N_31900,N_26830,N_27460);
and U31901 (N_31901,N_26337,N_26413);
or U31902 (N_31902,N_26461,N_26284);
nand U31903 (N_31903,N_29966,N_26645);
and U31904 (N_31904,N_26544,N_28236);
nand U31905 (N_31905,N_29766,N_29581);
xor U31906 (N_31906,N_25400,N_28316);
nand U31907 (N_31907,N_29076,N_28934);
or U31908 (N_31908,N_29888,N_27176);
xor U31909 (N_31909,N_26551,N_25657);
or U31910 (N_31910,N_29161,N_25503);
or U31911 (N_31911,N_29662,N_26490);
nand U31912 (N_31912,N_28393,N_25084);
nor U31913 (N_31913,N_26554,N_28603);
and U31914 (N_31914,N_27218,N_27043);
nand U31915 (N_31915,N_29238,N_26870);
or U31916 (N_31916,N_28532,N_25466);
or U31917 (N_31917,N_29914,N_28618);
nand U31918 (N_31918,N_29514,N_27664);
or U31919 (N_31919,N_25786,N_28791);
nand U31920 (N_31920,N_26160,N_25998);
nor U31921 (N_31921,N_29507,N_27042);
or U31922 (N_31922,N_29393,N_29987);
xnor U31923 (N_31923,N_27761,N_27272);
and U31924 (N_31924,N_29852,N_25114);
or U31925 (N_31925,N_27144,N_25569);
and U31926 (N_31926,N_27760,N_29369);
xor U31927 (N_31927,N_28408,N_29227);
xnor U31928 (N_31928,N_28554,N_25915);
and U31929 (N_31929,N_26907,N_28630);
or U31930 (N_31930,N_26820,N_27432);
nand U31931 (N_31931,N_25885,N_25351);
xnor U31932 (N_31932,N_25589,N_27902);
or U31933 (N_31933,N_28220,N_26036);
nand U31934 (N_31934,N_29492,N_25362);
and U31935 (N_31935,N_26180,N_26960);
xor U31936 (N_31936,N_28568,N_29724);
nor U31937 (N_31937,N_25329,N_26134);
nor U31938 (N_31938,N_28728,N_29778);
xor U31939 (N_31939,N_28790,N_25562);
or U31940 (N_31940,N_26290,N_27077);
and U31941 (N_31941,N_27498,N_27791);
and U31942 (N_31942,N_28083,N_29060);
nand U31943 (N_31943,N_28172,N_28619);
or U31944 (N_31944,N_27840,N_26679);
xnor U31945 (N_31945,N_29196,N_28692);
and U31946 (N_31946,N_29170,N_29872);
xnor U31947 (N_31947,N_27660,N_25526);
and U31948 (N_31948,N_26177,N_26834);
xor U31949 (N_31949,N_27423,N_26535);
nand U31950 (N_31950,N_26889,N_26802);
or U31951 (N_31951,N_26930,N_27910);
and U31952 (N_31952,N_29595,N_25004);
and U31953 (N_31953,N_28466,N_25148);
xnor U31954 (N_31954,N_28425,N_27440);
nand U31955 (N_31955,N_26246,N_28661);
nand U31956 (N_31956,N_27308,N_25769);
nand U31957 (N_31957,N_28600,N_29911);
and U31958 (N_31958,N_29819,N_26545);
nand U31959 (N_31959,N_27546,N_25819);
nor U31960 (N_31960,N_29734,N_29830);
xor U31961 (N_31961,N_27146,N_25719);
nor U31962 (N_31962,N_29098,N_27250);
xor U31963 (N_31963,N_25879,N_27788);
nor U31964 (N_31964,N_25411,N_28476);
nor U31965 (N_31965,N_28730,N_27569);
or U31966 (N_31966,N_29138,N_29467);
nor U31967 (N_31967,N_25010,N_26436);
xor U31968 (N_31968,N_27003,N_26934);
nand U31969 (N_31969,N_25355,N_26199);
and U31970 (N_31970,N_27665,N_25232);
nand U31971 (N_31971,N_25886,N_26054);
or U31972 (N_31972,N_26909,N_29558);
nand U31973 (N_31973,N_25518,N_28879);
or U31974 (N_31974,N_28895,N_25779);
nand U31975 (N_31975,N_25982,N_25870);
and U31976 (N_31976,N_27655,N_29271);
and U31977 (N_31977,N_28860,N_25810);
and U31978 (N_31978,N_26825,N_27345);
and U31979 (N_31979,N_27015,N_25533);
or U31980 (N_31980,N_28076,N_27895);
nor U31981 (N_31981,N_27037,N_28921);
or U31982 (N_31982,N_26675,N_25918);
or U31983 (N_31983,N_28039,N_26390);
nor U31984 (N_31984,N_28204,N_26977);
or U31985 (N_31985,N_29972,N_25785);
nand U31986 (N_31986,N_26381,N_26196);
nand U31987 (N_31987,N_28765,N_27400);
and U31988 (N_31988,N_28541,N_26033);
nor U31989 (N_31989,N_28175,N_28173);
nand U31990 (N_31990,N_27212,N_28377);
nand U31991 (N_31991,N_26494,N_29798);
xor U31992 (N_31992,N_28849,N_28659);
or U31993 (N_31993,N_29555,N_26026);
nand U31994 (N_31994,N_29168,N_26852);
and U31995 (N_31995,N_26586,N_25296);
nor U31996 (N_31996,N_25765,N_29538);
nand U31997 (N_31997,N_28813,N_25437);
or U31998 (N_31998,N_29188,N_25178);
nand U31999 (N_31999,N_28942,N_29899);
and U32000 (N_32000,N_25457,N_29928);
xor U32001 (N_32001,N_28292,N_26232);
xnor U32002 (N_32002,N_27646,N_25187);
nor U32003 (N_32003,N_26375,N_27135);
and U32004 (N_32004,N_25091,N_28844);
nand U32005 (N_32005,N_26169,N_26565);
xor U32006 (N_32006,N_25279,N_25218);
and U32007 (N_32007,N_28598,N_29442);
xor U32008 (N_32008,N_29267,N_29231);
or U32009 (N_32009,N_25336,N_27394);
or U32010 (N_32010,N_28472,N_28785);
or U32011 (N_32011,N_28441,N_29543);
xnor U32012 (N_32012,N_29705,N_25603);
or U32013 (N_32013,N_27931,N_28713);
or U32014 (N_32014,N_29509,N_27273);
nor U32015 (N_32015,N_27463,N_27315);
nand U32016 (N_32016,N_29263,N_27157);
nor U32017 (N_32017,N_28259,N_28018);
and U32018 (N_32018,N_29407,N_28559);
nand U32019 (N_32019,N_27576,N_28331);
nor U32020 (N_32020,N_26905,N_28013);
or U32021 (N_32021,N_26424,N_27847);
xor U32022 (N_32022,N_25102,N_26921);
or U32023 (N_32023,N_26226,N_29618);
nor U32024 (N_32024,N_26567,N_25677);
and U32025 (N_32025,N_25702,N_28822);
or U32026 (N_32026,N_26029,N_26468);
nand U32027 (N_32027,N_25840,N_28783);
nor U32028 (N_32028,N_29624,N_25245);
or U32029 (N_32029,N_25838,N_26628);
xnor U32030 (N_32030,N_28616,N_26289);
xor U32031 (N_32031,N_26013,N_25439);
nor U32032 (N_32032,N_26474,N_29166);
nor U32033 (N_32033,N_28863,N_28722);
nand U32034 (N_32034,N_29192,N_29018);
xor U32035 (N_32035,N_27662,N_29064);
nor U32036 (N_32036,N_28848,N_27243);
nor U32037 (N_32037,N_27923,N_28804);
xor U32038 (N_32038,N_29112,N_25224);
and U32039 (N_32039,N_29287,N_25039);
nand U32040 (N_32040,N_27161,N_26589);
or U32041 (N_32041,N_28203,N_26069);
nand U32042 (N_32042,N_25477,N_25834);
and U32043 (N_32043,N_27920,N_26791);
or U32044 (N_32044,N_26125,N_28570);
and U32045 (N_32045,N_28932,N_29037);
and U32046 (N_32046,N_27192,N_27928);
or U32047 (N_32047,N_29785,N_25225);
or U32048 (N_32048,N_28912,N_25163);
and U32049 (N_32049,N_29984,N_29348);
xor U32050 (N_32050,N_29020,N_25752);
xnor U32051 (N_32051,N_26439,N_25872);
nand U32052 (N_32052,N_29573,N_29976);
nand U32053 (N_32053,N_26152,N_27517);
or U32054 (N_32054,N_28845,N_26555);
and U32055 (N_32055,N_28913,N_28127);
xnor U32056 (N_32056,N_26585,N_29200);
or U32057 (N_32057,N_26005,N_27853);
nor U32058 (N_32058,N_27007,N_26728);
nand U32059 (N_32059,N_26722,N_27114);
nor U32060 (N_32060,N_25907,N_25173);
or U32061 (N_32061,N_28902,N_28533);
and U32062 (N_32062,N_28356,N_28696);
and U32063 (N_32063,N_27429,N_26928);
nor U32064 (N_32064,N_25471,N_29493);
or U32065 (N_32065,N_28206,N_27025);
and U32066 (N_32066,N_29149,N_26916);
nand U32067 (N_32067,N_25621,N_25718);
and U32068 (N_32068,N_25044,N_27252);
nor U32069 (N_32069,N_25228,N_25941);
or U32070 (N_32070,N_27875,N_28145);
and U32071 (N_32071,N_29948,N_29622);
nor U32072 (N_32072,N_28366,N_26323);
and U32073 (N_32073,N_27090,N_28385);
or U32074 (N_32074,N_25540,N_25079);
and U32075 (N_32075,N_27456,N_26339);
nand U32076 (N_32076,N_27782,N_29206);
or U32077 (N_32077,N_28182,N_25501);
xnor U32078 (N_32078,N_28896,N_28235);
xor U32079 (N_32079,N_29963,N_26434);
xor U32080 (N_32080,N_25388,N_27947);
xor U32081 (N_32081,N_29034,N_28805);
xor U32082 (N_32082,N_26781,N_27924);
nor U32083 (N_32083,N_28827,N_28991);
or U32084 (N_32084,N_25156,N_28384);
nand U32085 (N_32085,N_28578,N_25716);
xor U32086 (N_32086,N_25182,N_29136);
or U32087 (N_32087,N_27047,N_26462);
xor U32088 (N_32088,N_27155,N_26214);
and U32089 (N_32089,N_26546,N_28412);
nor U32090 (N_32090,N_25717,N_26713);
nand U32091 (N_32091,N_27014,N_26200);
and U32092 (N_32092,N_28736,N_28423);
nor U32093 (N_32093,N_29732,N_28418);
and U32094 (N_32094,N_29752,N_29481);
and U32095 (N_32095,N_26518,N_26271);
nor U32096 (N_32096,N_27763,N_29092);
or U32097 (N_32097,N_28294,N_29224);
nand U32098 (N_32098,N_25701,N_28154);
nand U32099 (N_32099,N_26765,N_26165);
nand U32100 (N_32100,N_25484,N_25016);
and U32101 (N_32101,N_29186,N_27299);
or U32102 (N_32102,N_26771,N_26888);
xnor U32103 (N_32103,N_25509,N_28654);
nand U32104 (N_32104,N_25293,N_26399);
and U32105 (N_32105,N_29474,N_28055);
and U32106 (N_32106,N_29388,N_29184);
nor U32107 (N_32107,N_25093,N_27496);
and U32108 (N_32108,N_27607,N_25316);
and U32109 (N_32109,N_25639,N_25541);
or U32110 (N_32110,N_29690,N_27486);
nand U32111 (N_32111,N_27635,N_26252);
nand U32112 (N_32112,N_25252,N_26560);
or U32113 (N_32113,N_27392,N_28962);
or U32114 (N_32114,N_27475,N_29866);
and U32115 (N_32115,N_29769,N_25054);
or U32116 (N_32116,N_29989,N_29411);
nor U32117 (N_32117,N_27621,N_27038);
or U32118 (N_32118,N_29510,N_26213);
or U32119 (N_32119,N_26306,N_29028);
and U32120 (N_32120,N_28909,N_25964);
or U32121 (N_32121,N_29383,N_29440);
or U32122 (N_32122,N_28628,N_25521);
or U32123 (N_32123,N_27661,N_27386);
nor U32124 (N_32124,N_26514,N_29741);
and U32125 (N_32125,N_28231,N_25531);
nor U32126 (N_32126,N_25222,N_27059);
nand U32127 (N_32127,N_25587,N_28638);
nor U32128 (N_32128,N_25896,N_25542);
nand U32129 (N_32129,N_27522,N_27332);
nand U32130 (N_32130,N_28005,N_28515);
or U32131 (N_32131,N_25254,N_26217);
xor U32132 (N_32132,N_28706,N_29808);
and U32133 (N_32133,N_26311,N_25882);
nor U32134 (N_32134,N_29241,N_28165);
nand U32135 (N_32135,N_29746,N_27229);
and U32136 (N_32136,N_25169,N_29464);
nor U32137 (N_32137,N_28834,N_25934);
or U32138 (N_32138,N_26162,N_27914);
nor U32139 (N_32139,N_29165,N_26429);
nand U32140 (N_32140,N_29355,N_25891);
nor U32141 (N_32141,N_25249,N_27351);
nor U32142 (N_32142,N_29199,N_28053);
and U32143 (N_32143,N_29907,N_27364);
and U32144 (N_32144,N_26269,N_28701);
xor U32145 (N_32145,N_28068,N_25147);
or U32146 (N_32146,N_28504,N_26932);
xor U32147 (N_32147,N_25679,N_28721);
xor U32148 (N_32148,N_29634,N_25046);
xnor U32149 (N_32149,N_25008,N_26952);
nand U32150 (N_32150,N_28066,N_29949);
or U32151 (N_32151,N_25479,N_25720);
and U32152 (N_32152,N_27552,N_28049);
nand U32153 (N_32153,N_25263,N_27680);
nand U32154 (N_32154,N_25920,N_29684);
nand U32155 (N_32155,N_27169,N_25788);
nand U32156 (N_32156,N_26297,N_26811);
nor U32157 (N_32157,N_29813,N_29887);
xnor U32158 (N_32158,N_25443,N_25754);
nor U32159 (N_32159,N_26974,N_27006);
nor U32160 (N_32160,N_26568,N_28419);
nor U32161 (N_32161,N_25024,N_26692);
xnor U32162 (N_32162,N_27866,N_29300);
nand U32163 (N_32163,N_25856,N_27181);
or U32164 (N_32164,N_27861,N_28698);
nand U32165 (N_32165,N_26168,N_29190);
xnor U32166 (N_32166,N_28594,N_27391);
nand U32167 (N_32167,N_28485,N_26503);
xnor U32168 (N_32168,N_25560,N_27339);
xnor U32169 (N_32169,N_25273,N_27723);
or U32170 (N_32170,N_25748,N_28446);
and U32171 (N_32171,N_26260,N_25199);
nand U32172 (N_32172,N_25243,N_26423);
or U32173 (N_32173,N_28886,N_28770);
or U32174 (N_32174,N_26419,N_29937);
xor U32175 (N_32175,N_29589,N_29598);
xnor U32176 (N_32176,N_28885,N_29443);
and U32177 (N_32177,N_28394,N_26014);
xor U32178 (N_32178,N_29744,N_29478);
nand U32179 (N_32179,N_27744,N_26824);
xnor U32180 (N_32180,N_29063,N_26412);
and U32181 (N_32181,N_26588,N_27061);
xor U32182 (N_32182,N_26062,N_25056);
xnor U32183 (N_32183,N_27408,N_29189);
or U32184 (N_32184,N_28341,N_27615);
xnor U32185 (N_32185,N_28903,N_27291);
xor U32186 (N_32186,N_27631,N_29133);
nand U32187 (N_32187,N_26658,N_29315);
or U32188 (N_32188,N_29834,N_28060);
and U32189 (N_32189,N_29349,N_25104);
and U32190 (N_32190,N_27357,N_25483);
or U32191 (N_32191,N_28327,N_26624);
xor U32192 (N_32192,N_26833,N_26303);
and U32193 (N_32193,N_28759,N_26295);
xnor U32194 (N_32194,N_28035,N_29007);
or U32195 (N_32195,N_25552,N_25726);
nor U32196 (N_32196,N_28904,N_29321);
xnor U32197 (N_32197,N_25704,N_25049);
or U32198 (N_32198,N_26119,N_25922);
and U32199 (N_32199,N_29220,N_27323);
nand U32200 (N_32200,N_29605,N_28340);
or U32201 (N_32201,N_27781,N_27980);
xor U32202 (N_32202,N_29410,N_28052);
and U32203 (N_32203,N_28817,N_25372);
or U32204 (N_32204,N_29781,N_26521);
or U32205 (N_32205,N_25699,N_27844);
nor U32206 (N_32206,N_28482,N_25066);
and U32207 (N_32207,N_25186,N_28514);
and U32208 (N_32208,N_28463,N_26384);
or U32209 (N_32209,N_29764,N_28312);
nor U32210 (N_32210,N_27515,N_27785);
xor U32211 (N_32211,N_25494,N_27700);
and U32212 (N_32212,N_27142,N_27177);
and U32213 (N_32213,N_28078,N_26007);
nand U32214 (N_32214,N_25327,N_27740);
nor U32215 (N_32215,N_28561,N_26764);
or U32216 (N_32216,N_26329,N_29867);
xor U32217 (N_32217,N_25902,N_26684);
xnor U32218 (N_32218,N_28534,N_29799);
nand U32219 (N_32219,N_25399,N_29456);
nand U32220 (N_32220,N_29805,N_27039);
xor U32221 (N_32221,N_25028,N_28918);
or U32222 (N_32222,N_27534,N_29988);
nor U32223 (N_32223,N_29387,N_27443);
nor U32224 (N_32224,N_25465,N_25628);
nor U32225 (N_32225,N_29632,N_26609);
or U32226 (N_32226,N_29416,N_28372);
nand U32227 (N_32227,N_27834,N_25829);
or U32228 (N_32228,N_29758,N_27745);
or U32229 (N_32229,N_25993,N_28077);
and U32230 (N_32230,N_28232,N_29804);
or U32231 (N_32231,N_28324,N_29114);
and U32232 (N_32232,N_28355,N_28162);
nor U32233 (N_32233,N_29965,N_26325);
nand U32234 (N_32234,N_28426,N_29931);
nor U32235 (N_32235,N_25160,N_29408);
nand U32236 (N_32236,N_29198,N_27995);
nand U32237 (N_32237,N_25166,N_29671);
xor U32238 (N_32238,N_26638,N_27317);
nand U32239 (N_32239,N_26239,N_28042);
or U32240 (N_32240,N_28072,N_27048);
and U32241 (N_32241,N_26998,N_27871);
and U32242 (N_32242,N_27395,N_25504);
and U32243 (N_32243,N_25247,N_26038);
nor U32244 (N_32244,N_28238,N_29048);
and U32245 (N_32245,N_25656,N_27800);
nand U32246 (N_32246,N_25342,N_25447);
nand U32247 (N_32247,N_25663,N_27150);
nor U32248 (N_32248,N_29302,N_27810);
or U32249 (N_32249,N_26006,N_27281);
nand U32250 (N_32250,N_26126,N_26480);
nor U32251 (N_32251,N_26404,N_27154);
and U32252 (N_32252,N_29803,N_28726);
or U32253 (N_32253,N_27836,N_28526);
and U32254 (N_32254,N_28180,N_25416);
xor U32255 (N_32255,N_25502,N_29071);
or U32256 (N_32256,N_26712,N_26488);
and U32257 (N_32257,N_25453,N_25129);
or U32258 (N_32258,N_26041,N_29239);
xnor U32259 (N_32259,N_29330,N_25450);
or U32260 (N_32260,N_29571,N_26577);
or U32261 (N_32261,N_28171,N_26965);
and U32262 (N_32262,N_29105,N_25805);
and U32263 (N_32263,N_29392,N_29396);
nand U32264 (N_32264,N_27951,N_25763);
nand U32265 (N_32265,N_26048,N_26842);
or U32266 (N_32266,N_26086,N_27668);
or U32267 (N_32267,N_26979,N_28492);
nand U32268 (N_32268,N_27625,N_28782);
and U32269 (N_32269,N_29373,N_25932);
and U32270 (N_32270,N_26766,N_28601);
xor U32271 (N_32271,N_28766,N_26394);
nor U32272 (N_32272,N_28117,N_29318);
xor U32273 (N_32273,N_29560,N_29569);
and U32274 (N_32274,N_26209,N_29616);
or U32275 (N_32275,N_27737,N_25954);
and U32276 (N_32276,N_29201,N_25444);
nor U32277 (N_32277,N_25863,N_27284);
xor U32278 (N_32278,N_25571,N_28674);
nor U32279 (N_32279,N_25729,N_26711);
nand U32280 (N_32280,N_25837,N_29296);
and U32281 (N_32281,N_26847,N_26925);
xnor U32282 (N_32282,N_27080,N_29334);
xor U32283 (N_32283,N_27028,N_25386);
and U32284 (N_32284,N_25813,N_25536);
xnor U32285 (N_32285,N_29557,N_28330);
nand U32286 (N_32286,N_26762,N_26328);
nand U32287 (N_32287,N_27632,N_27424);
nor U32288 (N_32288,N_27026,N_26072);
nand U32289 (N_32289,N_27021,N_27633);
nand U32290 (N_32290,N_27508,N_28870);
xor U32291 (N_32291,N_27557,N_28826);
nor U32292 (N_32292,N_28547,N_25088);
xor U32293 (N_32293,N_27855,N_25978);
xor U32294 (N_32294,N_25382,N_27396);
xnor U32295 (N_32295,N_28002,N_27953);
and U32296 (N_32296,N_25167,N_26091);
nand U32297 (N_32297,N_28497,N_26634);
nand U32298 (N_32298,N_29448,N_26291);
and U32299 (N_32299,N_26669,N_27197);
and U32300 (N_32300,N_28353,N_27667);
nor U32301 (N_32301,N_26077,N_26602);
nand U32302 (N_32302,N_26396,N_25195);
and U32303 (N_32303,N_27341,N_29606);
or U32304 (N_32304,N_26292,N_28097);
xor U32305 (N_32305,N_27255,N_26037);
xnor U32306 (N_32306,N_28337,N_27473);
or U32307 (N_32307,N_29786,N_25285);
xor U32308 (N_32308,N_29728,N_26919);
and U32309 (N_32309,N_25117,N_27183);
xor U32310 (N_32310,N_27410,N_27019);
or U32311 (N_32311,N_26946,N_27198);
xor U32312 (N_32312,N_29998,N_27581);
nand U32313 (N_32313,N_28893,N_27711);
nor U32314 (N_32314,N_28980,N_28362);
xor U32315 (N_32315,N_29950,N_29050);
xor U32316 (N_32316,N_25339,N_29426);
or U32317 (N_32317,N_27624,N_26019);
nand U32318 (N_32318,N_27837,N_25756);
and U32319 (N_32319,N_25481,N_28136);
or U32320 (N_32320,N_27693,N_25616);
nor U32321 (N_32321,N_27307,N_28432);
xnor U32322 (N_32322,N_25615,N_26702);
nand U32323 (N_32323,N_29285,N_27262);
xor U32324 (N_32324,N_27990,N_25352);
or U32325 (N_32325,N_29991,N_28134);
xor U32326 (N_32326,N_28321,N_29659);
nand U32327 (N_32327,N_25006,N_26897);
nor U32328 (N_32328,N_27712,N_25161);
nand U32329 (N_32329,N_25309,N_25832);
xnor U32330 (N_32330,N_29762,N_29176);
nand U32331 (N_32331,N_28746,N_26348);
and U32332 (N_32332,N_27519,N_25700);
and U32333 (N_32333,N_25668,N_27045);
xnor U32334 (N_32334,N_26195,N_29877);
and U32335 (N_32335,N_26616,N_26746);
nand U32336 (N_32336,N_29715,N_28686);
and U32337 (N_32337,N_27470,N_29544);
and U32338 (N_32338,N_25924,N_26813);
nand U32339 (N_32339,N_27128,N_28167);
and U32340 (N_32340,N_26982,N_26512);
nand U32341 (N_32341,N_29350,N_27689);
and U32342 (N_32342,N_25783,N_26505);
nor U32343 (N_32343,N_26446,N_26710);
and U32344 (N_32344,N_27276,N_25014);
nand U32345 (N_32345,N_25517,N_25445);
and U32346 (N_32346,N_28106,N_28033);
and U32347 (N_32347,N_28271,N_26613);
or U32348 (N_32348,N_29069,N_26202);
and U32349 (N_32349,N_28371,N_28414);
or U32350 (N_32350,N_26730,N_29842);
xor U32351 (N_32351,N_26189,N_26807);
xnor U32352 (N_32352,N_25592,N_29236);
nor U32353 (N_32353,N_26726,N_26143);
nor U32354 (N_32354,N_29787,N_29609);
and U32355 (N_32355,N_29667,N_26523);
or U32356 (N_32356,N_28855,N_29554);
or U32357 (N_32357,N_26445,N_28786);
xnor U32358 (N_32358,N_25687,N_25535);
xnor U32359 (N_32359,N_26188,N_25262);
nor U32360 (N_32360,N_28193,N_26719);
or U32361 (N_32361,N_25106,N_27725);
and U32362 (N_32362,N_25377,N_28511);
nor U32363 (N_32363,N_26324,N_29438);
xor U32364 (N_32364,N_26597,N_28961);
and U32365 (N_32365,N_29454,N_27851);
xnor U32366 (N_32366,N_29773,N_29779);
nor U32367 (N_32367,N_29579,N_25551);
xor U32368 (N_32368,N_27702,N_27330);
nand U32369 (N_32369,N_29089,N_29591);
xnor U32370 (N_32370,N_26818,N_27296);
and U32371 (N_32371,N_26395,N_29295);
or U32372 (N_32372,N_28143,N_26320);
xor U32373 (N_32373,N_28926,N_25874);
xnor U32374 (N_32374,N_27675,N_26225);
nor U32375 (N_32375,N_28110,N_28938);
and U32376 (N_32376,N_27981,N_27149);
or U32377 (N_32377,N_28975,N_26184);
nor U32378 (N_32378,N_28452,N_29956);
nand U32379 (N_32379,N_26782,N_25567);
or U32380 (N_32380,N_28122,N_28028);
nand U32381 (N_32381,N_25356,N_29584);
and U32382 (N_32382,N_27485,N_27991);
nor U32383 (N_32383,N_29629,N_28943);
nand U32384 (N_32384,N_28751,N_25658);
and U32385 (N_32385,N_26139,N_27807);
nor U32386 (N_32386,N_26040,N_27848);
nor U32387 (N_32387,N_26144,N_27439);
xnor U32388 (N_32388,N_27913,N_29056);
and U32389 (N_32389,N_28835,N_27796);
and U32390 (N_32390,N_29249,N_29946);
and U32391 (N_32391,N_25340,N_29685);
or U32392 (N_32392,N_25654,N_26759);
nand U32393 (N_32393,N_28712,N_28502);
or U32394 (N_32394,N_27421,N_29564);
nor U32395 (N_32395,N_27706,N_25866);
or U32396 (N_32396,N_28708,N_25581);
and U32397 (N_32397,N_25101,N_26313);
or U32398 (N_32398,N_28019,N_28960);
and U32399 (N_32399,N_25925,N_28462);
and U32400 (N_32400,N_28803,N_26355);
or U32401 (N_32401,N_27122,N_26527);
and U32402 (N_32402,N_27936,N_28544);
nor U32403 (N_32403,N_27147,N_29446);
nor U32404 (N_32404,N_25653,N_26886);
xnor U32405 (N_32405,N_28223,N_28798);
nor U32406 (N_32406,N_26242,N_27736);
nand U32407 (N_32407,N_29264,N_26939);
and U32408 (N_32408,N_25441,N_25043);
or U32409 (N_32409,N_28724,N_28840);
and U32410 (N_32410,N_29563,N_29142);
or U32411 (N_32411,N_25662,N_29647);
and U32412 (N_32412,N_25278,N_25670);
nand U32413 (N_32413,N_26460,N_27167);
xor U32414 (N_32414,N_26327,N_27282);
or U32415 (N_32415,N_27063,N_26487);
nand U32416 (N_32416,N_27574,N_28799);
or U32417 (N_32417,N_29995,N_29452);
xor U32418 (N_32418,N_25349,N_26515);
and U32419 (N_32419,N_27927,N_26153);
nor U32420 (N_32420,N_28907,N_26142);
nor U32421 (N_32421,N_29484,N_28265);
nor U32422 (N_32422,N_28329,N_28210);
or U32423 (N_32423,N_27941,N_28784);
nand U32424 (N_32424,N_28138,N_28081);
nand U32425 (N_32425,N_27190,N_29760);
nand U32426 (N_32426,N_28151,N_27874);
xnor U32427 (N_32427,N_25764,N_28518);
nor U32428 (N_32428,N_28109,N_26696);
or U32429 (N_32429,N_28757,N_26566);
nor U32430 (N_32430,N_25305,N_27018);
and U32431 (N_32431,N_28539,N_25368);
nand U32432 (N_32432,N_25292,N_25324);
or U32433 (N_32433,N_27354,N_26744);
nor U32434 (N_32434,N_28468,N_27798);
nor U32435 (N_32435,N_27459,N_26258);
xnor U32436 (N_32436,N_25200,N_25018);
and U32437 (N_32437,N_26838,N_27938);
and U32438 (N_32438,N_28748,N_27087);
or U32439 (N_32439,N_29266,N_28197);
nand U32440 (N_32440,N_25945,N_25828);
or U32441 (N_32441,N_26874,N_25513);
or U32442 (N_32442,N_29256,N_28908);
nand U32443 (N_32443,N_29384,N_29090);
nand U32444 (N_32444,N_25974,N_25808);
and U32445 (N_32445,N_25614,N_29642);
or U32446 (N_32446,N_27502,N_27230);
xor U32447 (N_32447,N_27717,N_28703);
and U32448 (N_32448,N_25348,N_27110);
nand U32449 (N_32449,N_28279,N_27297);
or U32450 (N_32450,N_27397,N_26754);
and U32451 (N_32451,N_29821,N_25505);
nor U32452 (N_32452,N_25052,N_27017);
and U32453 (N_32453,N_28710,N_27186);
nor U32454 (N_32454,N_29304,N_28823);
xor U32455 (N_32455,N_28079,N_26230);
xnor U32456 (N_32456,N_27694,N_29436);
xor U32457 (N_32457,N_28221,N_29134);
nand U32458 (N_32458,N_26906,N_29793);
nor U32459 (N_32459,N_29717,N_28672);
nand U32460 (N_32460,N_29472,N_26380);
nor U32461 (N_32461,N_28051,N_29046);
nor U32462 (N_32462,N_29466,N_27179);
xor U32463 (N_32463,N_26718,N_27975);
or U32464 (N_32464,N_28150,N_29993);
nor U32465 (N_32465,N_25612,N_28437);
and U32466 (N_32466,N_25965,N_26595);
or U32467 (N_32467,N_29169,N_29932);
nor U32468 (N_32468,N_27734,N_28417);
or U32469 (N_32469,N_29511,N_27636);
xor U32470 (N_32470,N_28454,N_29919);
nor U32471 (N_32471,N_29917,N_25686);
nand U32472 (N_32472,N_28359,N_26253);
nand U32473 (N_32473,N_27257,N_28084);
nand U32474 (N_32474,N_25625,N_28627);
xnor U32475 (N_32475,N_27464,N_28344);
nand U32476 (N_32476,N_25946,N_27965);
and U32477 (N_32477,N_27536,N_25648);
or U32478 (N_32478,N_27471,N_29228);
nor U32479 (N_32479,N_25814,N_25353);
nand U32480 (N_32480,N_26761,N_25193);
nor U32481 (N_32481,N_26016,N_27188);
and U32482 (N_32482,N_29245,N_26583);
and U32483 (N_32483,N_27240,N_29531);
and U32484 (N_32484,N_26356,N_27501);
and U32485 (N_32485,N_28239,N_26102);
or U32486 (N_32486,N_26821,N_25905);
nor U32487 (N_32487,N_26757,N_27316);
xnor U32488 (N_32488,N_28074,N_27237);
nand U32489 (N_32489,N_28413,N_27657);
xnor U32490 (N_32490,N_29843,N_25315);
or U32491 (N_32491,N_26865,N_28100);
or U32492 (N_32492,N_26161,N_25917);
xor U32493 (N_32493,N_25282,N_27720);
nor U32494 (N_32494,N_28222,N_27123);
xor U32495 (N_32495,N_28361,N_29951);
xor U32496 (N_32496,N_29422,N_25244);
and U32497 (N_32497,N_29641,N_26235);
nor U32498 (N_32498,N_25636,N_26749);
or U32499 (N_32499,N_27472,N_25761);
xnor U32500 (N_32500,N_25512,N_26180);
nor U32501 (N_32501,N_26809,N_27416);
or U32502 (N_32502,N_29003,N_26849);
and U32503 (N_32503,N_29749,N_26888);
nor U32504 (N_32504,N_26032,N_29832);
nor U32505 (N_32505,N_28793,N_28725);
xor U32506 (N_32506,N_26685,N_26622);
and U32507 (N_32507,N_29950,N_26333);
xnor U32508 (N_32508,N_28642,N_25511);
xnor U32509 (N_32509,N_29131,N_25103);
and U32510 (N_32510,N_25703,N_26330);
or U32511 (N_32511,N_26360,N_27547);
nor U32512 (N_32512,N_28642,N_28009);
or U32513 (N_32513,N_27182,N_29880);
nand U32514 (N_32514,N_28026,N_26188);
nor U32515 (N_32515,N_29705,N_27855);
or U32516 (N_32516,N_29627,N_25728);
xor U32517 (N_32517,N_26457,N_29608);
and U32518 (N_32518,N_28762,N_27029);
xor U32519 (N_32519,N_28927,N_28523);
nand U32520 (N_32520,N_25970,N_27015);
and U32521 (N_32521,N_26520,N_29691);
or U32522 (N_32522,N_26317,N_27193);
or U32523 (N_32523,N_28188,N_27249);
and U32524 (N_32524,N_25882,N_26631);
xor U32525 (N_32525,N_29668,N_29651);
and U32526 (N_32526,N_25219,N_26692);
and U32527 (N_32527,N_26076,N_29803);
xor U32528 (N_32528,N_27957,N_25850);
xnor U32529 (N_32529,N_26537,N_27766);
nor U32530 (N_32530,N_26577,N_26931);
xor U32531 (N_32531,N_29424,N_28904);
nor U32532 (N_32532,N_26573,N_25853);
and U32533 (N_32533,N_28724,N_29289);
or U32534 (N_32534,N_28416,N_26622);
nor U32535 (N_32535,N_29629,N_26388);
nand U32536 (N_32536,N_29306,N_26370);
xnor U32537 (N_32537,N_28416,N_28982);
nor U32538 (N_32538,N_28843,N_26095);
nand U32539 (N_32539,N_25083,N_27656);
nand U32540 (N_32540,N_25866,N_26090);
and U32541 (N_32541,N_25270,N_28415);
nand U32542 (N_32542,N_27991,N_29784);
and U32543 (N_32543,N_28828,N_25609);
or U32544 (N_32544,N_27971,N_28711);
nor U32545 (N_32545,N_26532,N_26745);
xor U32546 (N_32546,N_27115,N_29885);
nor U32547 (N_32547,N_25508,N_29217);
nand U32548 (N_32548,N_26975,N_25690);
or U32549 (N_32549,N_28182,N_27824);
nand U32550 (N_32550,N_28827,N_27827);
nand U32551 (N_32551,N_27747,N_29245);
nand U32552 (N_32552,N_25539,N_26625);
nor U32553 (N_32553,N_29518,N_29249);
nand U32554 (N_32554,N_28100,N_25187);
nor U32555 (N_32555,N_25500,N_27574);
or U32556 (N_32556,N_27511,N_28557);
nor U32557 (N_32557,N_26297,N_26415);
or U32558 (N_32558,N_27437,N_28227);
and U32559 (N_32559,N_28400,N_29029);
nor U32560 (N_32560,N_29379,N_27994);
and U32561 (N_32561,N_28358,N_25488);
or U32562 (N_32562,N_27968,N_25549);
and U32563 (N_32563,N_25650,N_27059);
or U32564 (N_32564,N_28924,N_29792);
or U32565 (N_32565,N_25642,N_25531);
nand U32566 (N_32566,N_28407,N_29825);
nand U32567 (N_32567,N_28374,N_25553);
xnor U32568 (N_32568,N_27890,N_25656);
or U32569 (N_32569,N_29801,N_25305);
xor U32570 (N_32570,N_28412,N_28151);
xor U32571 (N_32571,N_26075,N_25814);
or U32572 (N_32572,N_26077,N_28104);
or U32573 (N_32573,N_27752,N_25088);
nand U32574 (N_32574,N_29529,N_25460);
nor U32575 (N_32575,N_29129,N_28242);
xor U32576 (N_32576,N_27092,N_25415);
nor U32577 (N_32577,N_27582,N_26491);
nand U32578 (N_32578,N_26501,N_26039);
nor U32579 (N_32579,N_28895,N_29758);
xnor U32580 (N_32580,N_26298,N_27038);
xor U32581 (N_32581,N_25397,N_29772);
nand U32582 (N_32582,N_27002,N_25422);
xor U32583 (N_32583,N_26507,N_29999);
and U32584 (N_32584,N_26176,N_25836);
or U32585 (N_32585,N_25174,N_25212);
xor U32586 (N_32586,N_29663,N_29448);
nand U32587 (N_32587,N_27781,N_25245);
or U32588 (N_32588,N_25655,N_28158);
or U32589 (N_32589,N_27406,N_29470);
nand U32590 (N_32590,N_26098,N_28723);
and U32591 (N_32591,N_26052,N_27510);
nor U32592 (N_32592,N_25722,N_29122);
xnor U32593 (N_32593,N_25237,N_25705);
nor U32594 (N_32594,N_25865,N_28259);
or U32595 (N_32595,N_27545,N_25123);
nor U32596 (N_32596,N_26331,N_28352);
and U32597 (N_32597,N_28198,N_26722);
nor U32598 (N_32598,N_29457,N_25590);
and U32599 (N_32599,N_29599,N_29448);
xnor U32600 (N_32600,N_26484,N_26178);
nand U32601 (N_32601,N_28491,N_28025);
nor U32602 (N_32602,N_25852,N_28043);
nand U32603 (N_32603,N_29470,N_27226);
nand U32604 (N_32604,N_29574,N_28718);
xnor U32605 (N_32605,N_27677,N_26869);
or U32606 (N_32606,N_29185,N_27018);
xnor U32607 (N_32607,N_25810,N_27397);
xnor U32608 (N_32608,N_28749,N_28831);
xnor U32609 (N_32609,N_26669,N_28629);
or U32610 (N_32610,N_25689,N_27805);
and U32611 (N_32611,N_27161,N_29237);
xnor U32612 (N_32612,N_26151,N_29963);
nand U32613 (N_32613,N_25105,N_28256);
nand U32614 (N_32614,N_25202,N_25985);
nor U32615 (N_32615,N_28133,N_29935);
or U32616 (N_32616,N_28453,N_28658);
nor U32617 (N_32617,N_27484,N_29926);
nor U32618 (N_32618,N_28243,N_27906);
xor U32619 (N_32619,N_27109,N_28232);
nand U32620 (N_32620,N_26759,N_26006);
or U32621 (N_32621,N_27087,N_27627);
nor U32622 (N_32622,N_29649,N_27299);
nand U32623 (N_32623,N_25889,N_26835);
xor U32624 (N_32624,N_28338,N_28718);
xor U32625 (N_32625,N_29530,N_25266);
and U32626 (N_32626,N_28079,N_25113);
nor U32627 (N_32627,N_28739,N_28557);
or U32628 (N_32628,N_27531,N_27932);
nor U32629 (N_32629,N_29043,N_26012);
or U32630 (N_32630,N_26029,N_27513);
xnor U32631 (N_32631,N_26020,N_25049);
nor U32632 (N_32632,N_26079,N_25398);
xnor U32633 (N_32633,N_26522,N_29658);
nand U32634 (N_32634,N_26041,N_25894);
and U32635 (N_32635,N_25927,N_28420);
and U32636 (N_32636,N_28344,N_28226);
and U32637 (N_32637,N_28601,N_25607);
xor U32638 (N_32638,N_26239,N_26171);
or U32639 (N_32639,N_28078,N_27091);
or U32640 (N_32640,N_26209,N_26332);
nand U32641 (N_32641,N_25288,N_27484);
nand U32642 (N_32642,N_27221,N_26804);
nor U32643 (N_32643,N_29897,N_25380);
xnor U32644 (N_32644,N_25709,N_29103);
or U32645 (N_32645,N_28791,N_28317);
or U32646 (N_32646,N_26969,N_27004);
or U32647 (N_32647,N_29258,N_27563);
nand U32648 (N_32648,N_29298,N_26555);
nor U32649 (N_32649,N_25852,N_28061);
nand U32650 (N_32650,N_29000,N_28772);
xnor U32651 (N_32651,N_26483,N_29616);
nor U32652 (N_32652,N_25410,N_27008);
nor U32653 (N_32653,N_29173,N_29132);
nor U32654 (N_32654,N_26639,N_27644);
nand U32655 (N_32655,N_25573,N_29762);
or U32656 (N_32656,N_27099,N_28362);
and U32657 (N_32657,N_25030,N_29635);
or U32658 (N_32658,N_27176,N_27499);
xnor U32659 (N_32659,N_26011,N_25476);
and U32660 (N_32660,N_29544,N_27738);
xnor U32661 (N_32661,N_25581,N_28017);
nand U32662 (N_32662,N_29271,N_29946);
xnor U32663 (N_32663,N_27831,N_26943);
or U32664 (N_32664,N_27504,N_29378);
xor U32665 (N_32665,N_26873,N_27919);
nand U32666 (N_32666,N_28771,N_29823);
and U32667 (N_32667,N_26420,N_25079);
and U32668 (N_32668,N_26584,N_29708);
nand U32669 (N_32669,N_27649,N_25565);
and U32670 (N_32670,N_26507,N_28057);
nor U32671 (N_32671,N_25413,N_26814);
xnor U32672 (N_32672,N_26948,N_28904);
xor U32673 (N_32673,N_27162,N_28332);
or U32674 (N_32674,N_29793,N_29400);
xnor U32675 (N_32675,N_28830,N_26051);
and U32676 (N_32676,N_28808,N_26876);
nor U32677 (N_32677,N_27941,N_28757);
nor U32678 (N_32678,N_27825,N_28579);
or U32679 (N_32679,N_27330,N_25828);
xor U32680 (N_32680,N_25127,N_28824);
xnor U32681 (N_32681,N_26698,N_28453);
or U32682 (N_32682,N_29982,N_29133);
xor U32683 (N_32683,N_26009,N_25397);
or U32684 (N_32684,N_25926,N_25673);
and U32685 (N_32685,N_26277,N_25454);
and U32686 (N_32686,N_26897,N_29481);
or U32687 (N_32687,N_28080,N_25590);
and U32688 (N_32688,N_26238,N_25804);
nor U32689 (N_32689,N_28283,N_28795);
nor U32690 (N_32690,N_27041,N_28444);
and U32691 (N_32691,N_25089,N_28043);
xnor U32692 (N_32692,N_28498,N_27243);
nor U32693 (N_32693,N_29543,N_26487);
nand U32694 (N_32694,N_27512,N_26238);
xor U32695 (N_32695,N_29543,N_27234);
nor U32696 (N_32696,N_29117,N_25988);
nand U32697 (N_32697,N_25263,N_28675);
and U32698 (N_32698,N_28839,N_29786);
nor U32699 (N_32699,N_25099,N_27291);
nand U32700 (N_32700,N_27334,N_28654);
nand U32701 (N_32701,N_28453,N_25259);
nor U32702 (N_32702,N_25536,N_28570);
nand U32703 (N_32703,N_25954,N_28289);
or U32704 (N_32704,N_25961,N_25520);
nand U32705 (N_32705,N_27506,N_25090);
and U32706 (N_32706,N_26946,N_25497);
nor U32707 (N_32707,N_25259,N_25013);
nor U32708 (N_32708,N_28128,N_25160);
nor U32709 (N_32709,N_28054,N_27445);
nand U32710 (N_32710,N_29204,N_25163);
nand U32711 (N_32711,N_25747,N_25562);
nor U32712 (N_32712,N_28833,N_25744);
nor U32713 (N_32713,N_29203,N_27488);
xor U32714 (N_32714,N_28638,N_28209);
xnor U32715 (N_32715,N_29577,N_25153);
or U32716 (N_32716,N_26275,N_25115);
nor U32717 (N_32717,N_26405,N_29511);
or U32718 (N_32718,N_25310,N_28192);
xor U32719 (N_32719,N_27791,N_29677);
xnor U32720 (N_32720,N_26720,N_29963);
nor U32721 (N_32721,N_25311,N_29294);
nand U32722 (N_32722,N_28071,N_26316);
or U32723 (N_32723,N_25639,N_28897);
and U32724 (N_32724,N_25261,N_27642);
nand U32725 (N_32725,N_27841,N_27353);
xor U32726 (N_32726,N_28504,N_26553);
or U32727 (N_32727,N_29347,N_27588);
nand U32728 (N_32728,N_27683,N_25234);
nor U32729 (N_32729,N_28978,N_29659);
or U32730 (N_32730,N_27797,N_25466);
xnor U32731 (N_32731,N_29875,N_29356);
xor U32732 (N_32732,N_29599,N_27424);
or U32733 (N_32733,N_25208,N_27212);
or U32734 (N_32734,N_25513,N_28728);
and U32735 (N_32735,N_27611,N_28348);
xor U32736 (N_32736,N_26321,N_29563);
nor U32737 (N_32737,N_26584,N_26984);
and U32738 (N_32738,N_29548,N_29154);
and U32739 (N_32739,N_28712,N_29759);
and U32740 (N_32740,N_25933,N_26830);
nor U32741 (N_32741,N_25536,N_28599);
nor U32742 (N_32742,N_27817,N_28533);
or U32743 (N_32743,N_28886,N_28456);
nor U32744 (N_32744,N_29565,N_29972);
xnor U32745 (N_32745,N_28037,N_28378);
and U32746 (N_32746,N_28922,N_27680);
nand U32747 (N_32747,N_26472,N_27168);
and U32748 (N_32748,N_27991,N_27495);
xor U32749 (N_32749,N_26189,N_26685);
xnor U32750 (N_32750,N_28729,N_25699);
or U32751 (N_32751,N_28127,N_29681);
xnor U32752 (N_32752,N_29025,N_26346);
xor U32753 (N_32753,N_28429,N_26905);
or U32754 (N_32754,N_25087,N_25502);
nand U32755 (N_32755,N_28244,N_26407);
or U32756 (N_32756,N_26940,N_26273);
and U32757 (N_32757,N_25500,N_27142);
nand U32758 (N_32758,N_25963,N_29865);
or U32759 (N_32759,N_27777,N_28176);
nor U32760 (N_32760,N_27705,N_29129);
or U32761 (N_32761,N_29983,N_27628);
and U32762 (N_32762,N_25648,N_25366);
nand U32763 (N_32763,N_27138,N_26556);
xnor U32764 (N_32764,N_27977,N_29634);
nand U32765 (N_32765,N_26225,N_26450);
xor U32766 (N_32766,N_25155,N_29830);
nand U32767 (N_32767,N_28588,N_29666);
or U32768 (N_32768,N_27949,N_28214);
and U32769 (N_32769,N_26969,N_28385);
xnor U32770 (N_32770,N_27497,N_26055);
nand U32771 (N_32771,N_29207,N_27918);
or U32772 (N_32772,N_27054,N_27101);
xor U32773 (N_32773,N_28556,N_29587);
nor U32774 (N_32774,N_25119,N_29427);
nor U32775 (N_32775,N_25830,N_28978);
nand U32776 (N_32776,N_28463,N_29035);
nand U32777 (N_32777,N_25840,N_28345);
or U32778 (N_32778,N_25241,N_26493);
nand U32779 (N_32779,N_29585,N_26597);
nand U32780 (N_32780,N_26481,N_27076);
and U32781 (N_32781,N_26892,N_28319);
nand U32782 (N_32782,N_25632,N_27125);
or U32783 (N_32783,N_25973,N_29178);
xor U32784 (N_32784,N_26049,N_25083);
nand U32785 (N_32785,N_26987,N_25421);
nor U32786 (N_32786,N_27678,N_25621);
xnor U32787 (N_32787,N_25469,N_29357);
or U32788 (N_32788,N_26613,N_29884);
nor U32789 (N_32789,N_26383,N_27124);
nand U32790 (N_32790,N_29105,N_28321);
nand U32791 (N_32791,N_25854,N_28709);
xor U32792 (N_32792,N_27409,N_26365);
or U32793 (N_32793,N_26168,N_25095);
or U32794 (N_32794,N_25841,N_26508);
nor U32795 (N_32795,N_26561,N_26305);
nor U32796 (N_32796,N_25105,N_27561);
and U32797 (N_32797,N_27107,N_28381);
nand U32798 (N_32798,N_26673,N_25883);
xnor U32799 (N_32799,N_26401,N_29255);
or U32800 (N_32800,N_28224,N_26145);
and U32801 (N_32801,N_27582,N_25636);
and U32802 (N_32802,N_26427,N_26972);
or U32803 (N_32803,N_25249,N_28457);
nand U32804 (N_32804,N_25741,N_28778);
nor U32805 (N_32805,N_28712,N_27809);
nand U32806 (N_32806,N_28427,N_27938);
or U32807 (N_32807,N_27215,N_25671);
xor U32808 (N_32808,N_27053,N_28501);
nor U32809 (N_32809,N_28784,N_28588);
nor U32810 (N_32810,N_27548,N_28077);
or U32811 (N_32811,N_27435,N_29676);
nor U32812 (N_32812,N_28875,N_27185);
and U32813 (N_32813,N_29286,N_28552);
xnor U32814 (N_32814,N_26900,N_25470);
nor U32815 (N_32815,N_29901,N_26078);
or U32816 (N_32816,N_29382,N_27742);
nor U32817 (N_32817,N_25105,N_25855);
nand U32818 (N_32818,N_29041,N_25135);
xor U32819 (N_32819,N_28691,N_29784);
nor U32820 (N_32820,N_29940,N_28616);
and U32821 (N_32821,N_28200,N_26320);
and U32822 (N_32822,N_25868,N_28573);
and U32823 (N_32823,N_28041,N_26726);
xnor U32824 (N_32824,N_26791,N_26928);
xnor U32825 (N_32825,N_29731,N_27823);
nand U32826 (N_32826,N_28648,N_26813);
or U32827 (N_32827,N_29993,N_27425);
or U32828 (N_32828,N_26507,N_29638);
nor U32829 (N_32829,N_27387,N_28279);
or U32830 (N_32830,N_29376,N_27981);
nor U32831 (N_32831,N_26803,N_29269);
nor U32832 (N_32832,N_29791,N_28805);
nor U32833 (N_32833,N_25250,N_26304);
nand U32834 (N_32834,N_29524,N_25903);
nand U32835 (N_32835,N_26417,N_28658);
nor U32836 (N_32836,N_27467,N_28226);
and U32837 (N_32837,N_28675,N_27156);
nand U32838 (N_32838,N_27874,N_27285);
and U32839 (N_32839,N_25806,N_29008);
nand U32840 (N_32840,N_25457,N_28984);
xnor U32841 (N_32841,N_26495,N_29607);
nor U32842 (N_32842,N_26792,N_29976);
and U32843 (N_32843,N_25261,N_27221);
nor U32844 (N_32844,N_26564,N_29052);
or U32845 (N_32845,N_25805,N_28098);
or U32846 (N_32846,N_28686,N_28757);
or U32847 (N_32847,N_27954,N_27410);
xor U32848 (N_32848,N_26113,N_27264);
nor U32849 (N_32849,N_25843,N_25909);
and U32850 (N_32850,N_26774,N_28842);
and U32851 (N_32851,N_28143,N_25453);
xnor U32852 (N_32852,N_28271,N_25197);
and U32853 (N_32853,N_28272,N_28244);
nand U32854 (N_32854,N_26782,N_26041);
nand U32855 (N_32855,N_26054,N_28461);
xor U32856 (N_32856,N_29769,N_28853);
xor U32857 (N_32857,N_27366,N_26380);
or U32858 (N_32858,N_25018,N_27366);
nor U32859 (N_32859,N_25211,N_26700);
and U32860 (N_32860,N_28936,N_25152);
xor U32861 (N_32861,N_29634,N_28163);
nor U32862 (N_32862,N_29513,N_29541);
or U32863 (N_32863,N_25108,N_27090);
xor U32864 (N_32864,N_29545,N_29980);
or U32865 (N_32865,N_29399,N_28605);
nand U32866 (N_32866,N_28569,N_25929);
or U32867 (N_32867,N_28081,N_27400);
nand U32868 (N_32868,N_28143,N_29331);
nor U32869 (N_32869,N_29579,N_29207);
xnor U32870 (N_32870,N_29036,N_28117);
xnor U32871 (N_32871,N_29052,N_28042);
or U32872 (N_32872,N_26594,N_25004);
nand U32873 (N_32873,N_26523,N_26354);
nor U32874 (N_32874,N_29991,N_29974);
xnor U32875 (N_32875,N_25299,N_25673);
and U32876 (N_32876,N_26445,N_28795);
nor U32877 (N_32877,N_29240,N_25275);
xor U32878 (N_32878,N_25373,N_25033);
nor U32879 (N_32879,N_28704,N_25566);
and U32880 (N_32880,N_25809,N_27212);
nand U32881 (N_32881,N_27257,N_28268);
xnor U32882 (N_32882,N_26139,N_28230);
and U32883 (N_32883,N_29503,N_29688);
or U32884 (N_32884,N_29153,N_29761);
or U32885 (N_32885,N_28025,N_27522);
nor U32886 (N_32886,N_28426,N_28315);
or U32887 (N_32887,N_28593,N_27311);
nand U32888 (N_32888,N_26364,N_25823);
and U32889 (N_32889,N_25754,N_25106);
xnor U32890 (N_32890,N_27677,N_25161);
nor U32891 (N_32891,N_27205,N_25271);
nor U32892 (N_32892,N_27131,N_29236);
or U32893 (N_32893,N_28647,N_26366);
nand U32894 (N_32894,N_26425,N_25189);
nand U32895 (N_32895,N_26991,N_29617);
xnor U32896 (N_32896,N_29174,N_26731);
xor U32897 (N_32897,N_26429,N_26769);
nor U32898 (N_32898,N_29261,N_26614);
or U32899 (N_32899,N_28908,N_28198);
nand U32900 (N_32900,N_28271,N_28707);
xor U32901 (N_32901,N_26891,N_26904);
and U32902 (N_32902,N_29355,N_28821);
or U32903 (N_32903,N_27454,N_29104);
and U32904 (N_32904,N_25847,N_29374);
xor U32905 (N_32905,N_28842,N_28010);
nor U32906 (N_32906,N_26288,N_29020);
or U32907 (N_32907,N_25111,N_25609);
xnor U32908 (N_32908,N_26954,N_28093);
or U32909 (N_32909,N_29014,N_28408);
or U32910 (N_32910,N_28906,N_28356);
nand U32911 (N_32911,N_27224,N_25170);
or U32912 (N_32912,N_25084,N_27865);
xor U32913 (N_32913,N_26975,N_25110);
or U32914 (N_32914,N_29503,N_29259);
or U32915 (N_32915,N_26498,N_27786);
nand U32916 (N_32916,N_27289,N_26920);
nand U32917 (N_32917,N_25249,N_25882);
nand U32918 (N_32918,N_27024,N_27638);
xor U32919 (N_32919,N_27434,N_27849);
and U32920 (N_32920,N_26379,N_28590);
nand U32921 (N_32921,N_28223,N_25616);
nor U32922 (N_32922,N_25233,N_26517);
nand U32923 (N_32923,N_27032,N_25919);
and U32924 (N_32924,N_29413,N_25352);
and U32925 (N_32925,N_27115,N_28700);
nor U32926 (N_32926,N_29731,N_27001);
and U32927 (N_32927,N_28451,N_26176);
and U32928 (N_32928,N_29963,N_25016);
or U32929 (N_32929,N_27514,N_29547);
and U32930 (N_32930,N_25520,N_26069);
nor U32931 (N_32931,N_26852,N_29285);
nand U32932 (N_32932,N_28505,N_29158);
and U32933 (N_32933,N_29379,N_28423);
or U32934 (N_32934,N_28501,N_26302);
nand U32935 (N_32935,N_25390,N_26308);
and U32936 (N_32936,N_25162,N_29137);
nand U32937 (N_32937,N_28091,N_29695);
xor U32938 (N_32938,N_25262,N_25170);
or U32939 (N_32939,N_29668,N_29119);
nor U32940 (N_32940,N_26408,N_27344);
or U32941 (N_32941,N_26405,N_26339);
or U32942 (N_32942,N_29349,N_25416);
nand U32943 (N_32943,N_27646,N_29232);
and U32944 (N_32944,N_27979,N_28078);
nand U32945 (N_32945,N_27124,N_26054);
nand U32946 (N_32946,N_28964,N_28911);
or U32947 (N_32947,N_26229,N_29040);
xor U32948 (N_32948,N_25449,N_29661);
nor U32949 (N_32949,N_28974,N_27884);
and U32950 (N_32950,N_28420,N_27904);
nand U32951 (N_32951,N_26146,N_26861);
or U32952 (N_32952,N_29899,N_27381);
nand U32953 (N_32953,N_28497,N_25291);
nand U32954 (N_32954,N_29092,N_27631);
xnor U32955 (N_32955,N_26461,N_27541);
nand U32956 (N_32956,N_28066,N_26224);
xnor U32957 (N_32957,N_26996,N_29793);
nand U32958 (N_32958,N_27134,N_25625);
nor U32959 (N_32959,N_25155,N_26216);
nand U32960 (N_32960,N_29832,N_29405);
and U32961 (N_32961,N_27720,N_29035);
or U32962 (N_32962,N_26916,N_29381);
nor U32963 (N_32963,N_25971,N_29898);
nand U32964 (N_32964,N_27997,N_26446);
nand U32965 (N_32965,N_25075,N_26262);
xnor U32966 (N_32966,N_25548,N_26825);
and U32967 (N_32967,N_25687,N_29390);
nand U32968 (N_32968,N_25269,N_27874);
nor U32969 (N_32969,N_26855,N_25615);
nor U32970 (N_32970,N_28946,N_26026);
or U32971 (N_32971,N_28821,N_29477);
nor U32972 (N_32972,N_29735,N_27365);
xnor U32973 (N_32973,N_29113,N_25781);
or U32974 (N_32974,N_26001,N_27166);
xnor U32975 (N_32975,N_27984,N_26727);
nand U32976 (N_32976,N_27709,N_29768);
xor U32977 (N_32977,N_25237,N_25885);
or U32978 (N_32978,N_26856,N_25953);
nand U32979 (N_32979,N_26973,N_28120);
and U32980 (N_32980,N_29478,N_28747);
and U32981 (N_32981,N_28941,N_29846);
nor U32982 (N_32982,N_28885,N_26009);
and U32983 (N_32983,N_29754,N_26236);
nand U32984 (N_32984,N_27699,N_27518);
or U32985 (N_32985,N_27588,N_28192);
xnor U32986 (N_32986,N_28575,N_27976);
or U32987 (N_32987,N_27871,N_29931);
and U32988 (N_32988,N_25233,N_25487);
and U32989 (N_32989,N_28059,N_28729);
or U32990 (N_32990,N_26300,N_25618);
xor U32991 (N_32991,N_25592,N_28976);
xnor U32992 (N_32992,N_29503,N_28127);
xnor U32993 (N_32993,N_27114,N_28431);
nor U32994 (N_32994,N_29779,N_27876);
or U32995 (N_32995,N_27006,N_27681);
or U32996 (N_32996,N_28246,N_26187);
xnor U32997 (N_32997,N_25484,N_26282);
xor U32998 (N_32998,N_29920,N_25148);
and U32999 (N_32999,N_29015,N_25845);
nor U33000 (N_33000,N_28971,N_28254);
and U33001 (N_33001,N_26840,N_26100);
xor U33002 (N_33002,N_25194,N_27430);
xor U33003 (N_33003,N_26375,N_25520);
nand U33004 (N_33004,N_27745,N_25203);
and U33005 (N_33005,N_26032,N_27601);
or U33006 (N_33006,N_26358,N_29315);
nor U33007 (N_33007,N_27956,N_28054);
nor U33008 (N_33008,N_26715,N_28342);
xor U33009 (N_33009,N_29591,N_28057);
nor U33010 (N_33010,N_25551,N_25786);
xnor U33011 (N_33011,N_27136,N_26117);
and U33012 (N_33012,N_28305,N_29088);
nand U33013 (N_33013,N_28755,N_26341);
nand U33014 (N_33014,N_25176,N_29104);
nor U33015 (N_33015,N_26052,N_28789);
nor U33016 (N_33016,N_29594,N_26895);
and U33017 (N_33017,N_25545,N_26670);
and U33018 (N_33018,N_26441,N_29144);
or U33019 (N_33019,N_29336,N_25989);
nand U33020 (N_33020,N_27539,N_25552);
or U33021 (N_33021,N_27043,N_28106);
nand U33022 (N_33022,N_25168,N_27619);
or U33023 (N_33023,N_25666,N_25857);
nor U33024 (N_33024,N_28471,N_27622);
nor U33025 (N_33025,N_26945,N_25263);
nand U33026 (N_33026,N_25529,N_28577);
nor U33027 (N_33027,N_25954,N_25751);
or U33028 (N_33028,N_27202,N_26749);
nor U33029 (N_33029,N_26585,N_25786);
nand U33030 (N_33030,N_28496,N_29929);
xor U33031 (N_33031,N_27035,N_28255);
and U33032 (N_33032,N_26328,N_29619);
and U33033 (N_33033,N_28380,N_26928);
nand U33034 (N_33034,N_28537,N_25520);
and U33035 (N_33035,N_27480,N_27849);
nor U33036 (N_33036,N_26775,N_29813);
nand U33037 (N_33037,N_26954,N_26725);
or U33038 (N_33038,N_28353,N_28990);
and U33039 (N_33039,N_27453,N_26630);
xor U33040 (N_33040,N_28411,N_29924);
or U33041 (N_33041,N_27109,N_27643);
nor U33042 (N_33042,N_28810,N_25240);
and U33043 (N_33043,N_26262,N_27446);
nand U33044 (N_33044,N_29545,N_28981);
and U33045 (N_33045,N_27859,N_25904);
xnor U33046 (N_33046,N_28117,N_28057);
nor U33047 (N_33047,N_26311,N_29911);
and U33048 (N_33048,N_27929,N_28632);
or U33049 (N_33049,N_28215,N_28544);
xor U33050 (N_33050,N_27390,N_29017);
nand U33051 (N_33051,N_28724,N_29234);
and U33052 (N_33052,N_29328,N_28569);
xnor U33053 (N_33053,N_26365,N_25437);
nand U33054 (N_33054,N_27938,N_29396);
nand U33055 (N_33055,N_29795,N_27967);
nor U33056 (N_33056,N_25816,N_29281);
xnor U33057 (N_33057,N_25229,N_26736);
xnor U33058 (N_33058,N_29194,N_27053);
and U33059 (N_33059,N_26124,N_27566);
or U33060 (N_33060,N_26745,N_25803);
nand U33061 (N_33061,N_27671,N_25214);
or U33062 (N_33062,N_26355,N_27139);
or U33063 (N_33063,N_28755,N_29523);
nand U33064 (N_33064,N_25114,N_28062);
nand U33065 (N_33065,N_27336,N_29411);
xnor U33066 (N_33066,N_25315,N_25009);
or U33067 (N_33067,N_27016,N_28653);
nand U33068 (N_33068,N_29257,N_25832);
nand U33069 (N_33069,N_25591,N_26105);
nor U33070 (N_33070,N_26000,N_28636);
nor U33071 (N_33071,N_25843,N_25697);
or U33072 (N_33072,N_29783,N_27770);
xnor U33073 (N_33073,N_26785,N_25786);
xnor U33074 (N_33074,N_26114,N_29829);
nor U33075 (N_33075,N_27001,N_25088);
and U33076 (N_33076,N_25195,N_26641);
nor U33077 (N_33077,N_29700,N_27640);
or U33078 (N_33078,N_26653,N_25708);
nor U33079 (N_33079,N_27875,N_26153);
nand U33080 (N_33080,N_26625,N_28427);
nor U33081 (N_33081,N_29570,N_29938);
nand U33082 (N_33082,N_25054,N_27999);
nor U33083 (N_33083,N_25342,N_28612);
nand U33084 (N_33084,N_26613,N_28214);
nand U33085 (N_33085,N_26858,N_29481);
nand U33086 (N_33086,N_26433,N_29133);
nand U33087 (N_33087,N_27158,N_27485);
xor U33088 (N_33088,N_29848,N_29723);
and U33089 (N_33089,N_28722,N_27131);
nand U33090 (N_33090,N_27985,N_28497);
xor U33091 (N_33091,N_28961,N_25064);
nand U33092 (N_33092,N_26287,N_28837);
and U33093 (N_33093,N_27466,N_28289);
and U33094 (N_33094,N_25289,N_25972);
and U33095 (N_33095,N_29137,N_28211);
or U33096 (N_33096,N_29390,N_28726);
and U33097 (N_33097,N_25044,N_28095);
nand U33098 (N_33098,N_28592,N_29380);
nor U33099 (N_33099,N_29561,N_28390);
nand U33100 (N_33100,N_26640,N_25802);
nand U33101 (N_33101,N_26733,N_25446);
and U33102 (N_33102,N_27929,N_27637);
nand U33103 (N_33103,N_29054,N_26132);
nor U33104 (N_33104,N_26247,N_27402);
xor U33105 (N_33105,N_29862,N_27431);
and U33106 (N_33106,N_25421,N_27716);
or U33107 (N_33107,N_25569,N_29160);
nor U33108 (N_33108,N_28157,N_25335);
nor U33109 (N_33109,N_26832,N_28131);
nand U33110 (N_33110,N_26096,N_29729);
or U33111 (N_33111,N_28192,N_28639);
nand U33112 (N_33112,N_25767,N_29210);
and U33113 (N_33113,N_27027,N_29813);
nand U33114 (N_33114,N_27969,N_28108);
nor U33115 (N_33115,N_27671,N_27707);
nor U33116 (N_33116,N_26973,N_29563);
xnor U33117 (N_33117,N_26290,N_28335);
xor U33118 (N_33118,N_25860,N_27598);
and U33119 (N_33119,N_27534,N_26003);
and U33120 (N_33120,N_25743,N_25209);
nand U33121 (N_33121,N_28522,N_26133);
or U33122 (N_33122,N_27488,N_29513);
and U33123 (N_33123,N_25418,N_29924);
nor U33124 (N_33124,N_26411,N_25720);
or U33125 (N_33125,N_26445,N_29313);
nor U33126 (N_33126,N_25941,N_25137);
or U33127 (N_33127,N_25495,N_29330);
nor U33128 (N_33128,N_29904,N_28629);
nand U33129 (N_33129,N_26351,N_29082);
and U33130 (N_33130,N_28402,N_25906);
xor U33131 (N_33131,N_28013,N_26090);
nand U33132 (N_33132,N_29775,N_26058);
or U33133 (N_33133,N_26115,N_28323);
nand U33134 (N_33134,N_26597,N_27159);
and U33135 (N_33135,N_26039,N_28933);
nand U33136 (N_33136,N_29733,N_28681);
xor U33137 (N_33137,N_27453,N_25834);
xor U33138 (N_33138,N_28607,N_26477);
nand U33139 (N_33139,N_26719,N_28230);
and U33140 (N_33140,N_29068,N_27808);
nor U33141 (N_33141,N_29545,N_25586);
and U33142 (N_33142,N_25686,N_25853);
and U33143 (N_33143,N_29399,N_26715);
nand U33144 (N_33144,N_26531,N_25017);
and U33145 (N_33145,N_25275,N_28729);
nor U33146 (N_33146,N_29143,N_28745);
and U33147 (N_33147,N_26129,N_28698);
or U33148 (N_33148,N_29144,N_27786);
or U33149 (N_33149,N_25557,N_26566);
nand U33150 (N_33150,N_25977,N_29052);
and U33151 (N_33151,N_29919,N_26837);
nor U33152 (N_33152,N_28348,N_26308);
nand U33153 (N_33153,N_28824,N_27098);
nand U33154 (N_33154,N_29332,N_27764);
and U33155 (N_33155,N_27411,N_29765);
or U33156 (N_33156,N_27833,N_27361);
nor U33157 (N_33157,N_26512,N_26932);
or U33158 (N_33158,N_28011,N_25538);
nand U33159 (N_33159,N_27743,N_28728);
and U33160 (N_33160,N_28343,N_29706);
nor U33161 (N_33161,N_25345,N_27944);
or U33162 (N_33162,N_29873,N_26325);
or U33163 (N_33163,N_27124,N_26442);
and U33164 (N_33164,N_28988,N_25571);
nor U33165 (N_33165,N_28643,N_25830);
xnor U33166 (N_33166,N_25408,N_28079);
nand U33167 (N_33167,N_27516,N_28892);
and U33168 (N_33168,N_26591,N_29077);
or U33169 (N_33169,N_29281,N_27160);
and U33170 (N_33170,N_25970,N_26306);
xor U33171 (N_33171,N_26278,N_25078);
nor U33172 (N_33172,N_26030,N_26543);
xnor U33173 (N_33173,N_26783,N_29229);
nand U33174 (N_33174,N_27517,N_29755);
and U33175 (N_33175,N_25945,N_28568);
nand U33176 (N_33176,N_25138,N_29334);
and U33177 (N_33177,N_26511,N_26919);
or U33178 (N_33178,N_27271,N_28765);
xor U33179 (N_33179,N_26645,N_28945);
nor U33180 (N_33180,N_25514,N_28205);
xor U33181 (N_33181,N_27088,N_28548);
nand U33182 (N_33182,N_26775,N_26031);
nand U33183 (N_33183,N_29874,N_28566);
and U33184 (N_33184,N_29176,N_25828);
and U33185 (N_33185,N_28890,N_25244);
nand U33186 (N_33186,N_28950,N_29811);
nand U33187 (N_33187,N_29862,N_26950);
nand U33188 (N_33188,N_25483,N_27441);
or U33189 (N_33189,N_28789,N_25611);
xnor U33190 (N_33190,N_27197,N_25977);
nor U33191 (N_33191,N_27502,N_27474);
nand U33192 (N_33192,N_25446,N_26045);
nand U33193 (N_33193,N_25660,N_26260);
or U33194 (N_33194,N_25371,N_28213);
and U33195 (N_33195,N_26446,N_29165);
or U33196 (N_33196,N_29971,N_29855);
nor U33197 (N_33197,N_26124,N_26610);
nor U33198 (N_33198,N_28201,N_25464);
and U33199 (N_33199,N_26554,N_28278);
or U33200 (N_33200,N_29588,N_29222);
nor U33201 (N_33201,N_25482,N_28472);
nor U33202 (N_33202,N_29437,N_27597);
xor U33203 (N_33203,N_29827,N_27988);
or U33204 (N_33204,N_26246,N_28448);
xnor U33205 (N_33205,N_28354,N_28496);
nand U33206 (N_33206,N_29445,N_28734);
and U33207 (N_33207,N_28704,N_25655);
xor U33208 (N_33208,N_29441,N_29324);
xnor U33209 (N_33209,N_28177,N_27457);
and U33210 (N_33210,N_25850,N_25895);
nand U33211 (N_33211,N_25648,N_29749);
nand U33212 (N_33212,N_29415,N_25691);
and U33213 (N_33213,N_26521,N_25784);
xnor U33214 (N_33214,N_28240,N_25417);
nand U33215 (N_33215,N_28402,N_28186);
xnor U33216 (N_33216,N_29492,N_27695);
nor U33217 (N_33217,N_25914,N_26843);
nor U33218 (N_33218,N_26382,N_27721);
xnor U33219 (N_33219,N_26965,N_29887);
nand U33220 (N_33220,N_29559,N_27606);
and U33221 (N_33221,N_26263,N_29676);
or U33222 (N_33222,N_27981,N_29045);
xor U33223 (N_33223,N_27506,N_25922);
or U33224 (N_33224,N_26120,N_26110);
or U33225 (N_33225,N_28171,N_29297);
and U33226 (N_33226,N_27712,N_28985);
and U33227 (N_33227,N_25713,N_25262);
xor U33228 (N_33228,N_26838,N_29531);
xor U33229 (N_33229,N_29822,N_25333);
xnor U33230 (N_33230,N_28822,N_25080);
or U33231 (N_33231,N_25498,N_26511);
or U33232 (N_33232,N_25939,N_29188);
or U33233 (N_33233,N_28682,N_29169);
or U33234 (N_33234,N_29637,N_25069);
nor U33235 (N_33235,N_28862,N_28925);
and U33236 (N_33236,N_26913,N_26952);
xnor U33237 (N_33237,N_29745,N_25592);
and U33238 (N_33238,N_29279,N_29354);
and U33239 (N_33239,N_28936,N_29247);
nor U33240 (N_33240,N_27994,N_27135);
and U33241 (N_33241,N_27965,N_29345);
xnor U33242 (N_33242,N_29627,N_29520);
xor U33243 (N_33243,N_25063,N_25319);
nor U33244 (N_33244,N_29405,N_29896);
and U33245 (N_33245,N_27325,N_29407);
nor U33246 (N_33246,N_26315,N_27263);
nor U33247 (N_33247,N_27015,N_26108);
nor U33248 (N_33248,N_28315,N_29789);
xnor U33249 (N_33249,N_25648,N_26514);
or U33250 (N_33250,N_25960,N_25570);
or U33251 (N_33251,N_26109,N_28398);
nor U33252 (N_33252,N_26027,N_29489);
or U33253 (N_33253,N_29459,N_28580);
nor U33254 (N_33254,N_28704,N_29997);
nand U33255 (N_33255,N_29815,N_25182);
and U33256 (N_33256,N_27253,N_29700);
xor U33257 (N_33257,N_25747,N_25050);
xnor U33258 (N_33258,N_26382,N_27836);
and U33259 (N_33259,N_29046,N_26272);
and U33260 (N_33260,N_27194,N_26062);
or U33261 (N_33261,N_26655,N_27218);
or U33262 (N_33262,N_27570,N_29848);
or U33263 (N_33263,N_26409,N_27693);
and U33264 (N_33264,N_29258,N_26543);
nor U33265 (N_33265,N_27642,N_29165);
nor U33266 (N_33266,N_25374,N_28166);
nor U33267 (N_33267,N_29292,N_25560);
and U33268 (N_33268,N_26080,N_28807);
nor U33269 (N_33269,N_28559,N_28314);
xnor U33270 (N_33270,N_29049,N_27089);
or U33271 (N_33271,N_28565,N_28094);
xnor U33272 (N_33272,N_29912,N_28829);
or U33273 (N_33273,N_29041,N_29944);
or U33274 (N_33274,N_28365,N_25642);
nand U33275 (N_33275,N_25541,N_28527);
nand U33276 (N_33276,N_27643,N_28903);
xor U33277 (N_33277,N_29577,N_28334);
nand U33278 (N_33278,N_26259,N_25398);
or U33279 (N_33279,N_28051,N_28700);
or U33280 (N_33280,N_26865,N_28079);
nor U33281 (N_33281,N_29066,N_26906);
or U33282 (N_33282,N_27866,N_27020);
and U33283 (N_33283,N_28812,N_27935);
and U33284 (N_33284,N_26883,N_28143);
or U33285 (N_33285,N_29381,N_27603);
nand U33286 (N_33286,N_26486,N_25618);
xnor U33287 (N_33287,N_28083,N_26240);
xnor U33288 (N_33288,N_25757,N_29377);
and U33289 (N_33289,N_29085,N_27597);
nor U33290 (N_33290,N_28541,N_28534);
nand U33291 (N_33291,N_29635,N_26047);
xnor U33292 (N_33292,N_26361,N_29935);
xnor U33293 (N_33293,N_28252,N_25440);
or U33294 (N_33294,N_29854,N_27730);
nor U33295 (N_33295,N_26171,N_29508);
nor U33296 (N_33296,N_25258,N_28703);
and U33297 (N_33297,N_28847,N_27382);
nor U33298 (N_33298,N_26804,N_26610);
nor U33299 (N_33299,N_29092,N_27078);
and U33300 (N_33300,N_28151,N_25109);
and U33301 (N_33301,N_26805,N_29030);
or U33302 (N_33302,N_25092,N_28145);
and U33303 (N_33303,N_27981,N_26480);
xnor U33304 (N_33304,N_25093,N_29282);
nor U33305 (N_33305,N_26589,N_28033);
and U33306 (N_33306,N_29384,N_25074);
or U33307 (N_33307,N_25950,N_25397);
and U33308 (N_33308,N_28728,N_29671);
xor U33309 (N_33309,N_25536,N_25223);
nor U33310 (N_33310,N_29214,N_28528);
and U33311 (N_33311,N_29053,N_26890);
nor U33312 (N_33312,N_25991,N_27954);
nor U33313 (N_33313,N_28102,N_28419);
and U33314 (N_33314,N_25859,N_29088);
nor U33315 (N_33315,N_26055,N_25733);
xnor U33316 (N_33316,N_26567,N_29599);
and U33317 (N_33317,N_27208,N_26200);
xor U33318 (N_33318,N_28515,N_29587);
or U33319 (N_33319,N_27980,N_28505);
xnor U33320 (N_33320,N_26042,N_29633);
and U33321 (N_33321,N_27273,N_29040);
xor U33322 (N_33322,N_25612,N_26064);
xnor U33323 (N_33323,N_25784,N_29739);
xnor U33324 (N_33324,N_29666,N_26551);
nand U33325 (N_33325,N_28564,N_28242);
or U33326 (N_33326,N_28770,N_28282);
or U33327 (N_33327,N_26950,N_29789);
nand U33328 (N_33328,N_26782,N_28999);
nor U33329 (N_33329,N_26670,N_28377);
nor U33330 (N_33330,N_27305,N_26112);
nor U33331 (N_33331,N_28555,N_26479);
nor U33332 (N_33332,N_28877,N_26097);
or U33333 (N_33333,N_28102,N_26427);
xor U33334 (N_33334,N_28421,N_27037);
and U33335 (N_33335,N_29377,N_28516);
nand U33336 (N_33336,N_28563,N_29952);
nor U33337 (N_33337,N_28937,N_25272);
or U33338 (N_33338,N_25025,N_29103);
nor U33339 (N_33339,N_27355,N_29978);
or U33340 (N_33340,N_29123,N_28474);
nor U33341 (N_33341,N_27994,N_25894);
nand U33342 (N_33342,N_27337,N_28369);
nor U33343 (N_33343,N_28432,N_29629);
and U33344 (N_33344,N_29236,N_26862);
xnor U33345 (N_33345,N_27797,N_29989);
or U33346 (N_33346,N_25316,N_28502);
and U33347 (N_33347,N_28962,N_25320);
and U33348 (N_33348,N_25351,N_28340);
xnor U33349 (N_33349,N_26011,N_29252);
or U33350 (N_33350,N_25923,N_25974);
nor U33351 (N_33351,N_28615,N_28277);
xnor U33352 (N_33352,N_29895,N_28565);
nand U33353 (N_33353,N_28584,N_25461);
nand U33354 (N_33354,N_27692,N_28835);
and U33355 (N_33355,N_27534,N_28344);
xor U33356 (N_33356,N_25609,N_26230);
nand U33357 (N_33357,N_29041,N_28778);
nand U33358 (N_33358,N_26700,N_29650);
xnor U33359 (N_33359,N_27601,N_28968);
nor U33360 (N_33360,N_25106,N_27911);
nor U33361 (N_33361,N_29122,N_25253);
nand U33362 (N_33362,N_25697,N_27834);
nor U33363 (N_33363,N_26811,N_29796);
nor U33364 (N_33364,N_27752,N_28344);
or U33365 (N_33365,N_26397,N_28653);
xor U33366 (N_33366,N_26546,N_29452);
xnor U33367 (N_33367,N_28868,N_29403);
nand U33368 (N_33368,N_26341,N_27798);
nor U33369 (N_33369,N_25967,N_27496);
xnor U33370 (N_33370,N_29120,N_29682);
or U33371 (N_33371,N_29992,N_25538);
nor U33372 (N_33372,N_27389,N_25941);
xor U33373 (N_33373,N_29845,N_25222);
xor U33374 (N_33374,N_29275,N_28001);
and U33375 (N_33375,N_25214,N_26865);
xor U33376 (N_33376,N_29524,N_25651);
nand U33377 (N_33377,N_26173,N_25837);
or U33378 (N_33378,N_26396,N_28448);
or U33379 (N_33379,N_26140,N_27370);
nand U33380 (N_33380,N_25466,N_26876);
xor U33381 (N_33381,N_25094,N_26564);
and U33382 (N_33382,N_26793,N_26242);
or U33383 (N_33383,N_28478,N_28928);
or U33384 (N_33384,N_28668,N_29989);
nor U33385 (N_33385,N_27707,N_28782);
xnor U33386 (N_33386,N_26765,N_29141);
xor U33387 (N_33387,N_28519,N_26786);
xor U33388 (N_33388,N_29184,N_27611);
nor U33389 (N_33389,N_26173,N_26359);
and U33390 (N_33390,N_29429,N_27675);
and U33391 (N_33391,N_26393,N_26973);
and U33392 (N_33392,N_26044,N_26203);
or U33393 (N_33393,N_27633,N_26574);
nor U33394 (N_33394,N_25692,N_28244);
or U33395 (N_33395,N_28504,N_27098);
and U33396 (N_33396,N_26503,N_26938);
nor U33397 (N_33397,N_27415,N_29497);
xnor U33398 (N_33398,N_25294,N_26825);
xnor U33399 (N_33399,N_26240,N_25341);
or U33400 (N_33400,N_28304,N_28857);
nand U33401 (N_33401,N_26667,N_26714);
and U33402 (N_33402,N_28539,N_28469);
nor U33403 (N_33403,N_27375,N_25117);
nand U33404 (N_33404,N_26883,N_29607);
nand U33405 (N_33405,N_29855,N_27636);
nand U33406 (N_33406,N_26551,N_25785);
or U33407 (N_33407,N_26331,N_29799);
nand U33408 (N_33408,N_28342,N_28574);
xnor U33409 (N_33409,N_27740,N_26151);
or U33410 (N_33410,N_26895,N_28679);
nor U33411 (N_33411,N_25976,N_27440);
and U33412 (N_33412,N_25357,N_28526);
or U33413 (N_33413,N_27013,N_27208);
nand U33414 (N_33414,N_28075,N_28760);
nand U33415 (N_33415,N_29128,N_25679);
nor U33416 (N_33416,N_25196,N_25599);
nand U33417 (N_33417,N_27532,N_25270);
nand U33418 (N_33418,N_27781,N_26142);
or U33419 (N_33419,N_29453,N_28823);
or U33420 (N_33420,N_28257,N_27253);
nor U33421 (N_33421,N_25987,N_26675);
and U33422 (N_33422,N_28920,N_28122);
or U33423 (N_33423,N_28423,N_26456);
or U33424 (N_33424,N_25408,N_27317);
or U33425 (N_33425,N_25816,N_26170);
nor U33426 (N_33426,N_29112,N_27408);
or U33427 (N_33427,N_25852,N_29550);
and U33428 (N_33428,N_27612,N_29789);
nor U33429 (N_33429,N_26394,N_28230);
nand U33430 (N_33430,N_28083,N_28310);
nor U33431 (N_33431,N_27349,N_25885);
and U33432 (N_33432,N_25575,N_28271);
and U33433 (N_33433,N_28780,N_26420);
nor U33434 (N_33434,N_27061,N_29581);
xnor U33435 (N_33435,N_26809,N_26429);
nand U33436 (N_33436,N_26392,N_29934);
and U33437 (N_33437,N_25560,N_25930);
or U33438 (N_33438,N_27555,N_26515);
nor U33439 (N_33439,N_28793,N_27163);
and U33440 (N_33440,N_28231,N_25643);
xor U33441 (N_33441,N_27717,N_26294);
or U33442 (N_33442,N_28952,N_29429);
nand U33443 (N_33443,N_25493,N_29348);
nand U33444 (N_33444,N_25210,N_25611);
nand U33445 (N_33445,N_27165,N_28220);
xnor U33446 (N_33446,N_28984,N_26935);
or U33447 (N_33447,N_29554,N_27612);
xnor U33448 (N_33448,N_25024,N_27675);
nor U33449 (N_33449,N_26729,N_25361);
xnor U33450 (N_33450,N_26892,N_27932);
and U33451 (N_33451,N_29513,N_25627);
or U33452 (N_33452,N_26322,N_27233);
and U33453 (N_33453,N_27233,N_26795);
and U33454 (N_33454,N_26057,N_25735);
xnor U33455 (N_33455,N_26080,N_27682);
nand U33456 (N_33456,N_27321,N_26939);
or U33457 (N_33457,N_25149,N_29415);
or U33458 (N_33458,N_27100,N_26470);
nand U33459 (N_33459,N_26416,N_28594);
and U33460 (N_33460,N_27977,N_27938);
xnor U33461 (N_33461,N_26667,N_26166);
and U33462 (N_33462,N_29784,N_26773);
or U33463 (N_33463,N_27268,N_26304);
or U33464 (N_33464,N_28589,N_26869);
nor U33465 (N_33465,N_25017,N_25683);
or U33466 (N_33466,N_29027,N_27780);
and U33467 (N_33467,N_29037,N_27901);
nand U33468 (N_33468,N_27433,N_28588);
nand U33469 (N_33469,N_25998,N_28829);
and U33470 (N_33470,N_25580,N_28131);
xor U33471 (N_33471,N_27379,N_26388);
and U33472 (N_33472,N_29198,N_28630);
nand U33473 (N_33473,N_26510,N_29200);
and U33474 (N_33474,N_25199,N_26624);
and U33475 (N_33475,N_26781,N_25200);
or U33476 (N_33476,N_27213,N_28880);
and U33477 (N_33477,N_25734,N_28635);
xor U33478 (N_33478,N_25287,N_26308);
or U33479 (N_33479,N_25730,N_27620);
nand U33480 (N_33480,N_27233,N_25228);
nor U33481 (N_33481,N_29472,N_27950);
or U33482 (N_33482,N_25796,N_28347);
and U33483 (N_33483,N_26084,N_27362);
nand U33484 (N_33484,N_26000,N_25758);
and U33485 (N_33485,N_25142,N_26604);
nor U33486 (N_33486,N_27642,N_29166);
nor U33487 (N_33487,N_28004,N_27233);
nand U33488 (N_33488,N_25376,N_27653);
xnor U33489 (N_33489,N_28165,N_28355);
xnor U33490 (N_33490,N_27469,N_28437);
xnor U33491 (N_33491,N_28278,N_29949);
and U33492 (N_33492,N_27398,N_28741);
and U33493 (N_33493,N_25732,N_25219);
or U33494 (N_33494,N_25379,N_28506);
xnor U33495 (N_33495,N_29242,N_28971);
nand U33496 (N_33496,N_26561,N_27873);
nor U33497 (N_33497,N_28898,N_27605);
nor U33498 (N_33498,N_27587,N_29161);
and U33499 (N_33499,N_25257,N_29725);
or U33500 (N_33500,N_27102,N_29988);
or U33501 (N_33501,N_26031,N_27081);
nand U33502 (N_33502,N_29659,N_26036);
nand U33503 (N_33503,N_25674,N_27668);
nand U33504 (N_33504,N_29235,N_25103);
xnor U33505 (N_33505,N_26727,N_28709);
xnor U33506 (N_33506,N_25386,N_25576);
nor U33507 (N_33507,N_26576,N_25017);
xor U33508 (N_33508,N_25100,N_27476);
nor U33509 (N_33509,N_25981,N_29632);
and U33510 (N_33510,N_29699,N_27848);
and U33511 (N_33511,N_25434,N_25134);
and U33512 (N_33512,N_29510,N_28995);
nand U33513 (N_33513,N_28237,N_26482);
or U33514 (N_33514,N_29965,N_29198);
and U33515 (N_33515,N_27649,N_25494);
xor U33516 (N_33516,N_26701,N_28922);
xor U33517 (N_33517,N_25254,N_29574);
xnor U33518 (N_33518,N_27792,N_27715);
nand U33519 (N_33519,N_26040,N_25050);
xor U33520 (N_33520,N_28071,N_27229);
and U33521 (N_33521,N_28626,N_29867);
nor U33522 (N_33522,N_29100,N_25071);
xnor U33523 (N_33523,N_27063,N_29436);
and U33524 (N_33524,N_29560,N_29459);
xnor U33525 (N_33525,N_27290,N_28606);
nor U33526 (N_33526,N_29444,N_26060);
nor U33527 (N_33527,N_25666,N_25333);
or U33528 (N_33528,N_28442,N_29382);
xnor U33529 (N_33529,N_26439,N_26259);
or U33530 (N_33530,N_25018,N_29016);
nand U33531 (N_33531,N_25137,N_29006);
and U33532 (N_33532,N_27922,N_26222);
nor U33533 (N_33533,N_28731,N_29065);
xor U33534 (N_33534,N_25012,N_28145);
nor U33535 (N_33535,N_28118,N_25242);
and U33536 (N_33536,N_25456,N_27977);
nor U33537 (N_33537,N_28340,N_29738);
or U33538 (N_33538,N_29707,N_26801);
nand U33539 (N_33539,N_28348,N_25632);
nand U33540 (N_33540,N_25467,N_27510);
xor U33541 (N_33541,N_27547,N_27670);
xnor U33542 (N_33542,N_29401,N_27325);
or U33543 (N_33543,N_26704,N_27789);
nor U33544 (N_33544,N_26285,N_28228);
and U33545 (N_33545,N_26625,N_29580);
xor U33546 (N_33546,N_26458,N_25754);
and U33547 (N_33547,N_25700,N_25125);
or U33548 (N_33548,N_29423,N_28816);
xnor U33549 (N_33549,N_26849,N_25149);
xnor U33550 (N_33550,N_29588,N_26496);
and U33551 (N_33551,N_26424,N_27058);
and U33552 (N_33552,N_27690,N_26470);
xnor U33553 (N_33553,N_29112,N_27982);
nand U33554 (N_33554,N_28872,N_28425);
or U33555 (N_33555,N_27733,N_29723);
nor U33556 (N_33556,N_28973,N_25678);
nand U33557 (N_33557,N_25921,N_27822);
and U33558 (N_33558,N_27601,N_29921);
nor U33559 (N_33559,N_27442,N_28603);
or U33560 (N_33560,N_28388,N_28512);
or U33561 (N_33561,N_28705,N_25202);
nor U33562 (N_33562,N_28548,N_25800);
nand U33563 (N_33563,N_29762,N_26506);
xnor U33564 (N_33564,N_29268,N_28755);
nand U33565 (N_33565,N_25415,N_28472);
nand U33566 (N_33566,N_28211,N_28995);
or U33567 (N_33567,N_28249,N_25149);
or U33568 (N_33568,N_29525,N_25588);
nor U33569 (N_33569,N_28360,N_29971);
or U33570 (N_33570,N_26267,N_26641);
xnor U33571 (N_33571,N_28303,N_28354);
nand U33572 (N_33572,N_25163,N_25567);
xnor U33573 (N_33573,N_25757,N_27123);
nor U33574 (N_33574,N_25270,N_27760);
xor U33575 (N_33575,N_25750,N_25963);
nor U33576 (N_33576,N_29333,N_26864);
nor U33577 (N_33577,N_27923,N_25917);
nand U33578 (N_33578,N_26965,N_26650);
or U33579 (N_33579,N_27046,N_26109);
and U33580 (N_33580,N_27601,N_28239);
or U33581 (N_33581,N_28568,N_29445);
xor U33582 (N_33582,N_26544,N_28133);
or U33583 (N_33583,N_27767,N_26048);
xor U33584 (N_33584,N_26317,N_28184);
and U33585 (N_33585,N_26839,N_27016);
or U33586 (N_33586,N_29596,N_28545);
nand U33587 (N_33587,N_26431,N_28201);
nand U33588 (N_33588,N_27193,N_25316);
nand U33589 (N_33589,N_25228,N_29166);
or U33590 (N_33590,N_29688,N_28923);
xnor U33591 (N_33591,N_25845,N_27352);
xor U33592 (N_33592,N_27259,N_25397);
and U33593 (N_33593,N_26550,N_28273);
xnor U33594 (N_33594,N_25641,N_28665);
or U33595 (N_33595,N_29832,N_25728);
nor U33596 (N_33596,N_26908,N_27831);
xnor U33597 (N_33597,N_28072,N_28495);
and U33598 (N_33598,N_28726,N_26773);
nand U33599 (N_33599,N_26548,N_29003);
nor U33600 (N_33600,N_25514,N_26227);
nand U33601 (N_33601,N_29487,N_29854);
xor U33602 (N_33602,N_25906,N_27321);
nor U33603 (N_33603,N_25339,N_28767);
and U33604 (N_33604,N_28517,N_25391);
nor U33605 (N_33605,N_26927,N_29190);
or U33606 (N_33606,N_25557,N_28203);
nand U33607 (N_33607,N_27745,N_25762);
xor U33608 (N_33608,N_29097,N_26113);
and U33609 (N_33609,N_25870,N_28201);
or U33610 (N_33610,N_27501,N_26080);
nor U33611 (N_33611,N_26071,N_29022);
or U33612 (N_33612,N_28814,N_25092);
nor U33613 (N_33613,N_27149,N_25956);
and U33614 (N_33614,N_25912,N_28902);
nor U33615 (N_33615,N_29360,N_29290);
nor U33616 (N_33616,N_26993,N_27802);
nand U33617 (N_33617,N_27239,N_27583);
xor U33618 (N_33618,N_25894,N_28873);
nand U33619 (N_33619,N_29040,N_27199);
or U33620 (N_33620,N_29529,N_26979);
and U33621 (N_33621,N_27704,N_28819);
xnor U33622 (N_33622,N_29316,N_29712);
and U33623 (N_33623,N_26715,N_28547);
nand U33624 (N_33624,N_29974,N_26489);
and U33625 (N_33625,N_25218,N_27701);
or U33626 (N_33626,N_26967,N_25654);
or U33627 (N_33627,N_27672,N_26636);
nand U33628 (N_33628,N_25251,N_29893);
nand U33629 (N_33629,N_29577,N_25782);
or U33630 (N_33630,N_26271,N_28720);
xnor U33631 (N_33631,N_29353,N_27146);
nor U33632 (N_33632,N_29298,N_26021);
nand U33633 (N_33633,N_26685,N_29143);
and U33634 (N_33634,N_28355,N_27195);
nand U33635 (N_33635,N_25990,N_28397);
and U33636 (N_33636,N_27056,N_26021);
or U33637 (N_33637,N_25276,N_27850);
nand U33638 (N_33638,N_26985,N_29466);
xor U33639 (N_33639,N_25127,N_27062);
nand U33640 (N_33640,N_27494,N_27236);
or U33641 (N_33641,N_29761,N_25146);
and U33642 (N_33642,N_25474,N_26984);
or U33643 (N_33643,N_28592,N_29259);
nand U33644 (N_33644,N_29264,N_29292);
xor U33645 (N_33645,N_25103,N_25823);
and U33646 (N_33646,N_26606,N_25308);
and U33647 (N_33647,N_26170,N_29607);
nand U33648 (N_33648,N_28554,N_29135);
nand U33649 (N_33649,N_25060,N_25984);
nand U33650 (N_33650,N_28873,N_27066);
nand U33651 (N_33651,N_28616,N_25333);
or U33652 (N_33652,N_25051,N_25709);
nand U33653 (N_33653,N_27279,N_25018);
or U33654 (N_33654,N_25825,N_26983);
and U33655 (N_33655,N_28573,N_28977);
nor U33656 (N_33656,N_26222,N_28533);
or U33657 (N_33657,N_27867,N_27984);
or U33658 (N_33658,N_25021,N_27614);
or U33659 (N_33659,N_26558,N_26894);
or U33660 (N_33660,N_26211,N_29031);
nor U33661 (N_33661,N_27539,N_26752);
or U33662 (N_33662,N_28354,N_25739);
nand U33663 (N_33663,N_25370,N_28560);
nor U33664 (N_33664,N_27325,N_28833);
and U33665 (N_33665,N_28478,N_29086);
and U33666 (N_33666,N_25255,N_25343);
nor U33667 (N_33667,N_28035,N_26869);
and U33668 (N_33668,N_26545,N_29788);
and U33669 (N_33669,N_27838,N_27028);
or U33670 (N_33670,N_27833,N_25009);
or U33671 (N_33671,N_28421,N_28395);
xnor U33672 (N_33672,N_25562,N_29631);
or U33673 (N_33673,N_29675,N_26298);
xnor U33674 (N_33674,N_25011,N_28614);
and U33675 (N_33675,N_28508,N_26660);
and U33676 (N_33676,N_29515,N_27829);
or U33677 (N_33677,N_26842,N_27715);
or U33678 (N_33678,N_26596,N_27578);
and U33679 (N_33679,N_28549,N_29604);
and U33680 (N_33680,N_28004,N_26168);
xor U33681 (N_33681,N_25090,N_25225);
nand U33682 (N_33682,N_29001,N_26806);
and U33683 (N_33683,N_26497,N_25431);
nor U33684 (N_33684,N_25217,N_26267);
nand U33685 (N_33685,N_29795,N_27379);
and U33686 (N_33686,N_27090,N_29726);
or U33687 (N_33687,N_25726,N_29205);
nand U33688 (N_33688,N_27601,N_26918);
nor U33689 (N_33689,N_29667,N_28265);
and U33690 (N_33690,N_29698,N_29088);
nor U33691 (N_33691,N_29207,N_25419);
or U33692 (N_33692,N_28281,N_25190);
nand U33693 (N_33693,N_29720,N_27811);
nor U33694 (N_33694,N_25755,N_26235);
or U33695 (N_33695,N_26314,N_29500);
nor U33696 (N_33696,N_26581,N_28591);
nand U33697 (N_33697,N_26613,N_28822);
xnor U33698 (N_33698,N_25563,N_29174);
or U33699 (N_33699,N_25246,N_25558);
nand U33700 (N_33700,N_28041,N_26549);
xnor U33701 (N_33701,N_29829,N_27730);
nand U33702 (N_33702,N_26179,N_29605);
xor U33703 (N_33703,N_29625,N_25289);
nand U33704 (N_33704,N_28368,N_26870);
nor U33705 (N_33705,N_28629,N_26848);
or U33706 (N_33706,N_27776,N_28860);
nor U33707 (N_33707,N_27280,N_25178);
nand U33708 (N_33708,N_27957,N_25175);
nand U33709 (N_33709,N_27722,N_27921);
and U33710 (N_33710,N_25183,N_26684);
nor U33711 (N_33711,N_25119,N_25367);
xor U33712 (N_33712,N_29054,N_26165);
or U33713 (N_33713,N_28256,N_25552);
nand U33714 (N_33714,N_25264,N_27517);
nor U33715 (N_33715,N_25591,N_25330);
nor U33716 (N_33716,N_26324,N_28374);
or U33717 (N_33717,N_26496,N_26256);
xnor U33718 (N_33718,N_28866,N_25766);
or U33719 (N_33719,N_29045,N_27248);
xnor U33720 (N_33720,N_27161,N_27271);
and U33721 (N_33721,N_28588,N_27440);
or U33722 (N_33722,N_27863,N_28240);
xor U33723 (N_33723,N_25370,N_26783);
and U33724 (N_33724,N_25275,N_25589);
and U33725 (N_33725,N_25013,N_26435);
nor U33726 (N_33726,N_27376,N_28030);
or U33727 (N_33727,N_29926,N_29692);
nor U33728 (N_33728,N_25839,N_25939);
xor U33729 (N_33729,N_25704,N_27473);
nand U33730 (N_33730,N_28564,N_26947);
nand U33731 (N_33731,N_28532,N_29760);
nor U33732 (N_33732,N_29967,N_28166);
nor U33733 (N_33733,N_25190,N_25545);
or U33734 (N_33734,N_27425,N_29520);
and U33735 (N_33735,N_27012,N_29298);
xnor U33736 (N_33736,N_26599,N_27602);
nand U33737 (N_33737,N_28926,N_27242);
xnor U33738 (N_33738,N_25265,N_29172);
nor U33739 (N_33739,N_25991,N_29627);
nand U33740 (N_33740,N_27487,N_27923);
xor U33741 (N_33741,N_28898,N_26749);
nand U33742 (N_33742,N_28237,N_28670);
nor U33743 (N_33743,N_26770,N_27440);
xor U33744 (N_33744,N_26219,N_25719);
and U33745 (N_33745,N_29937,N_27916);
xor U33746 (N_33746,N_28678,N_27808);
nor U33747 (N_33747,N_29857,N_27958);
nand U33748 (N_33748,N_26661,N_27546);
or U33749 (N_33749,N_27267,N_29628);
and U33750 (N_33750,N_28550,N_26954);
or U33751 (N_33751,N_29135,N_25494);
xor U33752 (N_33752,N_25597,N_28858);
xnor U33753 (N_33753,N_28625,N_25553);
and U33754 (N_33754,N_25916,N_29325);
and U33755 (N_33755,N_29195,N_28752);
and U33756 (N_33756,N_26536,N_26912);
nor U33757 (N_33757,N_26895,N_29800);
or U33758 (N_33758,N_25754,N_28261);
nand U33759 (N_33759,N_25455,N_27183);
nor U33760 (N_33760,N_27858,N_25729);
or U33761 (N_33761,N_29421,N_27696);
nand U33762 (N_33762,N_29725,N_27246);
and U33763 (N_33763,N_27424,N_27492);
or U33764 (N_33764,N_28766,N_25745);
and U33765 (N_33765,N_28223,N_28471);
and U33766 (N_33766,N_27866,N_28254);
xnor U33767 (N_33767,N_26692,N_26008);
or U33768 (N_33768,N_27935,N_26789);
nor U33769 (N_33769,N_28755,N_26155);
and U33770 (N_33770,N_28348,N_29968);
nand U33771 (N_33771,N_27837,N_28374);
nand U33772 (N_33772,N_29736,N_26308);
nand U33773 (N_33773,N_28279,N_28095);
nor U33774 (N_33774,N_29910,N_25155);
xor U33775 (N_33775,N_28393,N_27364);
or U33776 (N_33776,N_28586,N_28030);
nand U33777 (N_33777,N_25141,N_25230);
or U33778 (N_33778,N_28484,N_25006);
xnor U33779 (N_33779,N_25990,N_25317);
nor U33780 (N_33780,N_26926,N_26180);
and U33781 (N_33781,N_27212,N_29313);
nand U33782 (N_33782,N_29541,N_25495);
xor U33783 (N_33783,N_26717,N_25407);
and U33784 (N_33784,N_25153,N_29940);
nand U33785 (N_33785,N_29220,N_28336);
xnor U33786 (N_33786,N_29814,N_27097);
and U33787 (N_33787,N_29740,N_28271);
or U33788 (N_33788,N_26382,N_28603);
nor U33789 (N_33789,N_28960,N_26939);
or U33790 (N_33790,N_26809,N_28728);
xor U33791 (N_33791,N_27250,N_29212);
xnor U33792 (N_33792,N_28080,N_27596);
nand U33793 (N_33793,N_26294,N_29917);
and U33794 (N_33794,N_29324,N_27564);
xor U33795 (N_33795,N_27554,N_28969);
nand U33796 (N_33796,N_29611,N_26841);
nor U33797 (N_33797,N_25894,N_28059);
nor U33798 (N_33798,N_27606,N_26389);
or U33799 (N_33799,N_26627,N_25810);
or U33800 (N_33800,N_26389,N_25601);
and U33801 (N_33801,N_27966,N_28516);
nand U33802 (N_33802,N_25459,N_28173);
or U33803 (N_33803,N_26815,N_26562);
nand U33804 (N_33804,N_25863,N_29265);
nand U33805 (N_33805,N_28485,N_28893);
or U33806 (N_33806,N_25320,N_25847);
and U33807 (N_33807,N_29572,N_25440);
xor U33808 (N_33808,N_25656,N_27573);
xnor U33809 (N_33809,N_25446,N_25966);
nor U33810 (N_33810,N_28059,N_28275);
xor U33811 (N_33811,N_25905,N_29191);
xor U33812 (N_33812,N_25809,N_25646);
or U33813 (N_33813,N_28490,N_26705);
nand U33814 (N_33814,N_27175,N_27831);
nand U33815 (N_33815,N_26969,N_27535);
or U33816 (N_33816,N_27935,N_28018);
and U33817 (N_33817,N_25330,N_29899);
nor U33818 (N_33818,N_25859,N_28267);
nor U33819 (N_33819,N_27928,N_28145);
or U33820 (N_33820,N_26865,N_25981);
and U33821 (N_33821,N_26958,N_27445);
and U33822 (N_33822,N_29175,N_28888);
or U33823 (N_33823,N_26586,N_25189);
and U33824 (N_33824,N_26096,N_27492);
or U33825 (N_33825,N_28253,N_25441);
nor U33826 (N_33826,N_25905,N_28428);
and U33827 (N_33827,N_26579,N_25138);
nand U33828 (N_33828,N_28605,N_26768);
nor U33829 (N_33829,N_26593,N_25871);
and U33830 (N_33830,N_26824,N_28979);
and U33831 (N_33831,N_26617,N_28849);
or U33832 (N_33832,N_26904,N_25316);
nor U33833 (N_33833,N_26036,N_29818);
nor U33834 (N_33834,N_28911,N_29337);
or U33835 (N_33835,N_29823,N_26502);
xnor U33836 (N_33836,N_26259,N_29547);
xor U33837 (N_33837,N_29788,N_29316);
nand U33838 (N_33838,N_29728,N_25604);
and U33839 (N_33839,N_28650,N_28346);
and U33840 (N_33840,N_28627,N_28272);
xor U33841 (N_33841,N_26191,N_27423);
or U33842 (N_33842,N_29503,N_26129);
nand U33843 (N_33843,N_25986,N_26347);
xnor U33844 (N_33844,N_27286,N_26576);
nand U33845 (N_33845,N_29668,N_29318);
or U33846 (N_33846,N_27645,N_25013);
nor U33847 (N_33847,N_25053,N_29629);
and U33848 (N_33848,N_29045,N_28643);
xor U33849 (N_33849,N_29376,N_29144);
nor U33850 (N_33850,N_29397,N_27500);
xnor U33851 (N_33851,N_28157,N_26774);
and U33852 (N_33852,N_25312,N_28717);
nand U33853 (N_33853,N_27800,N_26497);
or U33854 (N_33854,N_27807,N_25983);
or U33855 (N_33855,N_27104,N_25921);
xor U33856 (N_33856,N_29678,N_28330);
nor U33857 (N_33857,N_27992,N_29816);
nand U33858 (N_33858,N_29214,N_29055);
xnor U33859 (N_33859,N_25067,N_26472);
xor U33860 (N_33860,N_29750,N_25915);
nor U33861 (N_33861,N_27258,N_26278);
nand U33862 (N_33862,N_28001,N_26349);
and U33863 (N_33863,N_25478,N_25246);
nor U33864 (N_33864,N_28616,N_27863);
and U33865 (N_33865,N_29934,N_27138);
or U33866 (N_33866,N_29033,N_26491);
nor U33867 (N_33867,N_25547,N_25179);
nor U33868 (N_33868,N_27560,N_28240);
xor U33869 (N_33869,N_26676,N_25495);
nand U33870 (N_33870,N_27698,N_28899);
nor U33871 (N_33871,N_27952,N_27673);
or U33872 (N_33872,N_27726,N_27972);
nand U33873 (N_33873,N_27539,N_28868);
xnor U33874 (N_33874,N_26626,N_28912);
nand U33875 (N_33875,N_29094,N_29915);
xnor U33876 (N_33876,N_27072,N_27715);
xnor U33877 (N_33877,N_27395,N_27689);
and U33878 (N_33878,N_27903,N_28630);
xor U33879 (N_33879,N_29300,N_25564);
xnor U33880 (N_33880,N_28105,N_29868);
nand U33881 (N_33881,N_25923,N_29650);
xnor U33882 (N_33882,N_29048,N_26610);
xnor U33883 (N_33883,N_25275,N_28041);
and U33884 (N_33884,N_26736,N_27346);
or U33885 (N_33885,N_25327,N_26304);
and U33886 (N_33886,N_28376,N_26841);
nor U33887 (N_33887,N_27275,N_26210);
or U33888 (N_33888,N_29183,N_29914);
and U33889 (N_33889,N_28800,N_25726);
and U33890 (N_33890,N_28000,N_29916);
xnor U33891 (N_33891,N_28181,N_29586);
or U33892 (N_33892,N_27939,N_28331);
nand U33893 (N_33893,N_25106,N_27901);
nor U33894 (N_33894,N_29828,N_26702);
and U33895 (N_33895,N_27998,N_25813);
xor U33896 (N_33896,N_26992,N_29505);
or U33897 (N_33897,N_28533,N_25154);
or U33898 (N_33898,N_27412,N_26057);
xor U33899 (N_33899,N_27439,N_29717);
nor U33900 (N_33900,N_29823,N_29555);
xnor U33901 (N_33901,N_25864,N_26812);
or U33902 (N_33902,N_27155,N_28934);
nor U33903 (N_33903,N_27773,N_29839);
and U33904 (N_33904,N_26879,N_25242);
and U33905 (N_33905,N_26418,N_25291);
nor U33906 (N_33906,N_27739,N_27432);
xnor U33907 (N_33907,N_25284,N_29837);
xor U33908 (N_33908,N_28332,N_29704);
nor U33909 (N_33909,N_27156,N_29278);
nor U33910 (N_33910,N_26103,N_25734);
nor U33911 (N_33911,N_26947,N_29614);
nand U33912 (N_33912,N_25850,N_28404);
and U33913 (N_33913,N_25637,N_27551);
and U33914 (N_33914,N_26379,N_28501);
or U33915 (N_33915,N_26811,N_26642);
and U33916 (N_33916,N_25026,N_29266);
xor U33917 (N_33917,N_28915,N_26244);
nand U33918 (N_33918,N_29181,N_25422);
and U33919 (N_33919,N_28529,N_29974);
and U33920 (N_33920,N_26818,N_28843);
xnor U33921 (N_33921,N_27095,N_26523);
and U33922 (N_33922,N_26416,N_28607);
nand U33923 (N_33923,N_25750,N_26118);
nor U33924 (N_33924,N_28561,N_28857);
xnor U33925 (N_33925,N_25374,N_25242);
nor U33926 (N_33926,N_29558,N_27403);
or U33927 (N_33927,N_25094,N_26459);
or U33928 (N_33928,N_25080,N_27081);
or U33929 (N_33929,N_29420,N_28018);
and U33930 (N_33930,N_25248,N_25523);
nand U33931 (N_33931,N_29236,N_29905);
nand U33932 (N_33932,N_29358,N_25039);
or U33933 (N_33933,N_26671,N_26020);
and U33934 (N_33934,N_25867,N_27496);
and U33935 (N_33935,N_28489,N_27178);
nor U33936 (N_33936,N_27090,N_28547);
xnor U33937 (N_33937,N_29347,N_28946);
nor U33938 (N_33938,N_25208,N_29559);
or U33939 (N_33939,N_29055,N_26388);
and U33940 (N_33940,N_26510,N_27901);
nand U33941 (N_33941,N_29277,N_28343);
nor U33942 (N_33942,N_27253,N_29154);
and U33943 (N_33943,N_28953,N_27091);
nor U33944 (N_33944,N_25800,N_27343);
or U33945 (N_33945,N_27168,N_28761);
xor U33946 (N_33946,N_29584,N_27902);
xor U33947 (N_33947,N_26025,N_27489);
or U33948 (N_33948,N_27386,N_27414);
xor U33949 (N_33949,N_25442,N_29484);
xor U33950 (N_33950,N_26511,N_28685);
or U33951 (N_33951,N_29659,N_27967);
nor U33952 (N_33952,N_25034,N_29378);
nor U33953 (N_33953,N_25030,N_29012);
xnor U33954 (N_33954,N_25923,N_29099);
xor U33955 (N_33955,N_29712,N_25958);
or U33956 (N_33956,N_29313,N_27400);
or U33957 (N_33957,N_25396,N_27515);
and U33958 (N_33958,N_26121,N_28203);
nor U33959 (N_33959,N_26901,N_26062);
nand U33960 (N_33960,N_29649,N_26352);
nand U33961 (N_33961,N_25757,N_29043);
or U33962 (N_33962,N_29395,N_25765);
and U33963 (N_33963,N_25527,N_29092);
xor U33964 (N_33964,N_27612,N_27347);
xor U33965 (N_33965,N_26848,N_27247);
and U33966 (N_33966,N_25301,N_29182);
and U33967 (N_33967,N_28141,N_27695);
xor U33968 (N_33968,N_26680,N_28702);
xor U33969 (N_33969,N_27730,N_27185);
or U33970 (N_33970,N_28318,N_28784);
nand U33971 (N_33971,N_27011,N_25641);
nand U33972 (N_33972,N_28364,N_25426);
xnor U33973 (N_33973,N_29703,N_25693);
xnor U33974 (N_33974,N_29262,N_26286);
and U33975 (N_33975,N_27223,N_28092);
or U33976 (N_33976,N_29231,N_26587);
and U33977 (N_33977,N_28658,N_28183);
or U33978 (N_33978,N_28309,N_26967);
nor U33979 (N_33979,N_29484,N_29643);
xor U33980 (N_33980,N_25072,N_26758);
or U33981 (N_33981,N_28789,N_29307);
or U33982 (N_33982,N_26076,N_25451);
and U33983 (N_33983,N_26432,N_29660);
nor U33984 (N_33984,N_26216,N_29230);
nand U33985 (N_33985,N_29038,N_27670);
and U33986 (N_33986,N_29526,N_25219);
or U33987 (N_33987,N_25863,N_29365);
and U33988 (N_33988,N_28230,N_25919);
nand U33989 (N_33989,N_28406,N_29240);
xor U33990 (N_33990,N_29105,N_27579);
nand U33991 (N_33991,N_29481,N_27864);
nand U33992 (N_33992,N_27296,N_29798);
or U33993 (N_33993,N_28354,N_27244);
nand U33994 (N_33994,N_27432,N_29193);
and U33995 (N_33995,N_29362,N_29539);
xnor U33996 (N_33996,N_28454,N_25680);
nand U33997 (N_33997,N_28183,N_27925);
or U33998 (N_33998,N_29377,N_25048);
nor U33999 (N_33999,N_29442,N_26225);
xor U34000 (N_34000,N_26550,N_28624);
xor U34001 (N_34001,N_25267,N_27706);
nor U34002 (N_34002,N_29027,N_28416);
xor U34003 (N_34003,N_25624,N_25206);
xnor U34004 (N_34004,N_29765,N_27844);
or U34005 (N_34005,N_25372,N_28631);
or U34006 (N_34006,N_26131,N_26543);
nand U34007 (N_34007,N_26872,N_28357);
or U34008 (N_34008,N_29549,N_25254);
or U34009 (N_34009,N_27735,N_25557);
and U34010 (N_34010,N_25099,N_25329);
nand U34011 (N_34011,N_28644,N_25482);
or U34012 (N_34012,N_25602,N_27677);
nand U34013 (N_34013,N_28380,N_29837);
nand U34014 (N_34014,N_26951,N_27338);
xnor U34015 (N_34015,N_28415,N_29174);
xnor U34016 (N_34016,N_28981,N_29563);
and U34017 (N_34017,N_26684,N_29167);
nor U34018 (N_34018,N_28017,N_25733);
xnor U34019 (N_34019,N_29561,N_29498);
or U34020 (N_34020,N_29127,N_25924);
xor U34021 (N_34021,N_27039,N_26544);
nor U34022 (N_34022,N_28339,N_26111);
or U34023 (N_34023,N_25340,N_28708);
nand U34024 (N_34024,N_26451,N_26695);
and U34025 (N_34025,N_26399,N_29968);
nand U34026 (N_34026,N_27827,N_26478);
nor U34027 (N_34027,N_27863,N_26712);
or U34028 (N_34028,N_27259,N_26321);
or U34029 (N_34029,N_25072,N_25449);
and U34030 (N_34030,N_26442,N_26149);
and U34031 (N_34031,N_25537,N_27497);
or U34032 (N_34032,N_27198,N_27019);
or U34033 (N_34033,N_28380,N_28785);
nor U34034 (N_34034,N_29205,N_27139);
or U34035 (N_34035,N_25942,N_26694);
xnor U34036 (N_34036,N_25672,N_29127);
xor U34037 (N_34037,N_29624,N_29197);
xnor U34038 (N_34038,N_25029,N_28897);
nor U34039 (N_34039,N_27190,N_25524);
or U34040 (N_34040,N_27721,N_25974);
nand U34041 (N_34041,N_27506,N_29854);
or U34042 (N_34042,N_29583,N_25163);
nor U34043 (N_34043,N_28489,N_28514);
or U34044 (N_34044,N_29940,N_25627);
or U34045 (N_34045,N_27218,N_28087);
and U34046 (N_34046,N_27687,N_28300);
nor U34047 (N_34047,N_27457,N_29756);
or U34048 (N_34048,N_25322,N_25885);
or U34049 (N_34049,N_25438,N_29873);
or U34050 (N_34050,N_28258,N_29493);
nor U34051 (N_34051,N_26436,N_28302);
and U34052 (N_34052,N_27559,N_27953);
nor U34053 (N_34053,N_29629,N_25590);
nand U34054 (N_34054,N_27250,N_29684);
and U34055 (N_34055,N_27953,N_25877);
xor U34056 (N_34056,N_29480,N_25911);
nor U34057 (N_34057,N_25930,N_26223);
and U34058 (N_34058,N_29769,N_25056);
nor U34059 (N_34059,N_28089,N_26249);
xnor U34060 (N_34060,N_28055,N_27771);
nand U34061 (N_34061,N_25263,N_27807);
and U34062 (N_34062,N_28846,N_28417);
nor U34063 (N_34063,N_26326,N_29210);
or U34064 (N_34064,N_29427,N_28685);
nor U34065 (N_34065,N_26330,N_25899);
nor U34066 (N_34066,N_25764,N_27339);
or U34067 (N_34067,N_25473,N_28478);
or U34068 (N_34068,N_29461,N_28945);
xor U34069 (N_34069,N_28787,N_27932);
and U34070 (N_34070,N_26062,N_28467);
or U34071 (N_34071,N_29561,N_28901);
xor U34072 (N_34072,N_26691,N_29501);
nor U34073 (N_34073,N_29273,N_25025);
xor U34074 (N_34074,N_25096,N_26216);
nand U34075 (N_34075,N_29889,N_28292);
nor U34076 (N_34076,N_26607,N_26829);
nor U34077 (N_34077,N_26482,N_27861);
and U34078 (N_34078,N_26190,N_27128);
nand U34079 (N_34079,N_27125,N_27565);
nand U34080 (N_34080,N_29249,N_26625);
nand U34081 (N_34081,N_28962,N_25906);
xnor U34082 (N_34082,N_27831,N_25287);
nand U34083 (N_34083,N_28673,N_28334);
nor U34084 (N_34084,N_27615,N_27808);
nand U34085 (N_34085,N_27560,N_26516);
and U34086 (N_34086,N_26644,N_28277);
and U34087 (N_34087,N_27813,N_25194);
or U34088 (N_34088,N_25773,N_28318);
xor U34089 (N_34089,N_29007,N_26471);
nor U34090 (N_34090,N_26072,N_26407);
or U34091 (N_34091,N_25038,N_28631);
xnor U34092 (N_34092,N_27140,N_25351);
nand U34093 (N_34093,N_26664,N_27985);
nand U34094 (N_34094,N_28876,N_29858);
and U34095 (N_34095,N_26516,N_28149);
xor U34096 (N_34096,N_28101,N_26282);
or U34097 (N_34097,N_25617,N_25248);
and U34098 (N_34098,N_27369,N_29785);
nand U34099 (N_34099,N_25513,N_28446);
xnor U34100 (N_34100,N_28645,N_25850);
or U34101 (N_34101,N_27797,N_25155);
nand U34102 (N_34102,N_28405,N_27446);
xor U34103 (N_34103,N_25834,N_25980);
nor U34104 (N_34104,N_25160,N_27252);
nor U34105 (N_34105,N_25185,N_26883);
and U34106 (N_34106,N_26597,N_28671);
nor U34107 (N_34107,N_27170,N_28262);
nor U34108 (N_34108,N_29036,N_25562);
nand U34109 (N_34109,N_25153,N_29210);
or U34110 (N_34110,N_26298,N_28934);
or U34111 (N_34111,N_25581,N_26215);
nand U34112 (N_34112,N_29499,N_29498);
xor U34113 (N_34113,N_25182,N_26978);
and U34114 (N_34114,N_25676,N_25160);
xnor U34115 (N_34115,N_28939,N_26308);
or U34116 (N_34116,N_28763,N_29542);
nor U34117 (N_34117,N_25900,N_26422);
and U34118 (N_34118,N_29490,N_26063);
or U34119 (N_34119,N_26937,N_27377);
nand U34120 (N_34120,N_28883,N_28473);
xor U34121 (N_34121,N_29175,N_29571);
and U34122 (N_34122,N_26018,N_29586);
and U34123 (N_34123,N_25346,N_26776);
and U34124 (N_34124,N_25593,N_25266);
nand U34125 (N_34125,N_29489,N_29868);
xor U34126 (N_34126,N_28778,N_28763);
nor U34127 (N_34127,N_27160,N_25605);
nor U34128 (N_34128,N_29164,N_28308);
and U34129 (N_34129,N_27557,N_28273);
nand U34130 (N_34130,N_25898,N_26496);
nand U34131 (N_34131,N_29279,N_26428);
and U34132 (N_34132,N_25397,N_25790);
nor U34133 (N_34133,N_25698,N_29021);
xor U34134 (N_34134,N_25957,N_28434);
or U34135 (N_34135,N_25170,N_27303);
or U34136 (N_34136,N_26953,N_28722);
nor U34137 (N_34137,N_28078,N_26996);
nand U34138 (N_34138,N_27722,N_29792);
or U34139 (N_34139,N_27527,N_27369);
or U34140 (N_34140,N_29742,N_26168);
and U34141 (N_34141,N_25588,N_28684);
nor U34142 (N_34142,N_26572,N_29847);
nor U34143 (N_34143,N_25102,N_25345);
xor U34144 (N_34144,N_28909,N_27820);
xor U34145 (N_34145,N_29503,N_29146);
nor U34146 (N_34146,N_29906,N_28650);
nor U34147 (N_34147,N_27440,N_25618);
and U34148 (N_34148,N_25781,N_25525);
and U34149 (N_34149,N_29147,N_27140);
nor U34150 (N_34150,N_28675,N_29848);
nand U34151 (N_34151,N_26510,N_26383);
xor U34152 (N_34152,N_26064,N_29587);
nor U34153 (N_34153,N_27046,N_28780);
and U34154 (N_34154,N_27851,N_29589);
or U34155 (N_34155,N_29411,N_29833);
and U34156 (N_34156,N_28953,N_29297);
xor U34157 (N_34157,N_25399,N_25842);
or U34158 (N_34158,N_25857,N_27767);
nand U34159 (N_34159,N_26608,N_29480);
or U34160 (N_34160,N_29572,N_28541);
nor U34161 (N_34161,N_29278,N_27146);
and U34162 (N_34162,N_26073,N_25331);
nand U34163 (N_34163,N_27605,N_29043);
nand U34164 (N_34164,N_28167,N_25892);
xor U34165 (N_34165,N_25895,N_29105);
nand U34166 (N_34166,N_25437,N_28283);
nor U34167 (N_34167,N_29314,N_27080);
and U34168 (N_34168,N_25985,N_26466);
and U34169 (N_34169,N_28039,N_26549);
or U34170 (N_34170,N_29260,N_27339);
or U34171 (N_34171,N_28096,N_29692);
or U34172 (N_34172,N_26459,N_26160);
and U34173 (N_34173,N_26620,N_26192);
or U34174 (N_34174,N_27062,N_29358);
nand U34175 (N_34175,N_27171,N_27097);
xnor U34176 (N_34176,N_28735,N_29225);
nand U34177 (N_34177,N_27965,N_25880);
xnor U34178 (N_34178,N_28253,N_27982);
or U34179 (N_34179,N_29445,N_27435);
nor U34180 (N_34180,N_29217,N_28631);
or U34181 (N_34181,N_26726,N_25452);
nor U34182 (N_34182,N_25065,N_27558);
and U34183 (N_34183,N_27198,N_26550);
xor U34184 (N_34184,N_25016,N_29575);
or U34185 (N_34185,N_28885,N_25317);
or U34186 (N_34186,N_28638,N_27355);
and U34187 (N_34187,N_28139,N_26408);
or U34188 (N_34188,N_28023,N_25582);
or U34189 (N_34189,N_29863,N_29697);
or U34190 (N_34190,N_29786,N_27295);
xor U34191 (N_34191,N_26612,N_25518);
or U34192 (N_34192,N_28068,N_29850);
nand U34193 (N_34193,N_28300,N_29844);
and U34194 (N_34194,N_27764,N_26234);
nor U34195 (N_34195,N_28456,N_26404);
xnor U34196 (N_34196,N_29445,N_26683);
or U34197 (N_34197,N_25800,N_25662);
nor U34198 (N_34198,N_27283,N_29655);
xor U34199 (N_34199,N_29008,N_29150);
or U34200 (N_34200,N_27437,N_27371);
xor U34201 (N_34201,N_27036,N_25067);
nand U34202 (N_34202,N_27865,N_28063);
nand U34203 (N_34203,N_28326,N_25004);
and U34204 (N_34204,N_26437,N_26783);
and U34205 (N_34205,N_26879,N_25407);
xnor U34206 (N_34206,N_26894,N_29619);
or U34207 (N_34207,N_25477,N_28799);
or U34208 (N_34208,N_27571,N_27084);
nand U34209 (N_34209,N_28418,N_26285);
and U34210 (N_34210,N_26591,N_26084);
and U34211 (N_34211,N_25033,N_29397);
nand U34212 (N_34212,N_25357,N_27475);
and U34213 (N_34213,N_26912,N_26633);
or U34214 (N_34214,N_27303,N_25541);
or U34215 (N_34215,N_26175,N_26225);
xnor U34216 (N_34216,N_28340,N_25727);
nor U34217 (N_34217,N_29763,N_27100);
xnor U34218 (N_34218,N_25751,N_28935);
nand U34219 (N_34219,N_27364,N_27485);
and U34220 (N_34220,N_27644,N_29355);
nand U34221 (N_34221,N_25313,N_27590);
xor U34222 (N_34222,N_29558,N_29259);
or U34223 (N_34223,N_28021,N_26847);
xor U34224 (N_34224,N_28171,N_26598);
or U34225 (N_34225,N_27604,N_27863);
xnor U34226 (N_34226,N_25523,N_27098);
nand U34227 (N_34227,N_26535,N_29512);
and U34228 (N_34228,N_28528,N_29074);
and U34229 (N_34229,N_27936,N_28771);
and U34230 (N_34230,N_29107,N_27388);
nand U34231 (N_34231,N_26035,N_29059);
or U34232 (N_34232,N_25044,N_27368);
or U34233 (N_34233,N_29438,N_29782);
nor U34234 (N_34234,N_26747,N_29043);
xnor U34235 (N_34235,N_27787,N_26733);
or U34236 (N_34236,N_29187,N_28056);
nor U34237 (N_34237,N_26352,N_29335);
or U34238 (N_34238,N_27931,N_27007);
or U34239 (N_34239,N_27973,N_28432);
xor U34240 (N_34240,N_26759,N_28441);
nor U34241 (N_34241,N_25526,N_29578);
and U34242 (N_34242,N_27441,N_25389);
or U34243 (N_34243,N_26663,N_28927);
and U34244 (N_34244,N_28806,N_25802);
nand U34245 (N_34245,N_26364,N_25997);
or U34246 (N_34246,N_26141,N_25256);
and U34247 (N_34247,N_25826,N_28957);
xor U34248 (N_34248,N_29386,N_27377);
xor U34249 (N_34249,N_29004,N_26530);
xnor U34250 (N_34250,N_28754,N_26230);
and U34251 (N_34251,N_27658,N_26344);
or U34252 (N_34252,N_26735,N_27972);
and U34253 (N_34253,N_29047,N_27928);
xor U34254 (N_34254,N_25068,N_28194);
nand U34255 (N_34255,N_27927,N_26387);
and U34256 (N_34256,N_29504,N_27900);
nand U34257 (N_34257,N_25817,N_26170);
nor U34258 (N_34258,N_28497,N_25000);
nor U34259 (N_34259,N_29646,N_29310);
xor U34260 (N_34260,N_28589,N_27389);
or U34261 (N_34261,N_29148,N_27769);
xor U34262 (N_34262,N_26118,N_26445);
or U34263 (N_34263,N_28204,N_26920);
and U34264 (N_34264,N_27474,N_27413);
xor U34265 (N_34265,N_25378,N_28511);
xor U34266 (N_34266,N_27315,N_29683);
and U34267 (N_34267,N_25474,N_28741);
nor U34268 (N_34268,N_27184,N_28471);
or U34269 (N_34269,N_28380,N_27094);
nand U34270 (N_34270,N_25659,N_27369);
and U34271 (N_34271,N_29474,N_25589);
and U34272 (N_34272,N_27352,N_26375);
nor U34273 (N_34273,N_27438,N_27334);
nand U34274 (N_34274,N_29328,N_26287);
or U34275 (N_34275,N_29463,N_29035);
xor U34276 (N_34276,N_27357,N_25236);
or U34277 (N_34277,N_27032,N_28049);
xnor U34278 (N_34278,N_27175,N_25149);
or U34279 (N_34279,N_26664,N_26505);
or U34280 (N_34280,N_26823,N_29824);
xor U34281 (N_34281,N_29738,N_27656);
nand U34282 (N_34282,N_25365,N_27041);
and U34283 (N_34283,N_25787,N_29167);
or U34284 (N_34284,N_25973,N_29125);
or U34285 (N_34285,N_28664,N_29115);
and U34286 (N_34286,N_26792,N_26829);
nor U34287 (N_34287,N_27436,N_26428);
nand U34288 (N_34288,N_29603,N_29508);
or U34289 (N_34289,N_29803,N_27591);
and U34290 (N_34290,N_29856,N_29811);
nor U34291 (N_34291,N_25224,N_29884);
and U34292 (N_34292,N_27303,N_27631);
nand U34293 (N_34293,N_26237,N_28975);
and U34294 (N_34294,N_29166,N_26934);
xnor U34295 (N_34295,N_28848,N_25551);
and U34296 (N_34296,N_28924,N_26566);
nand U34297 (N_34297,N_29711,N_26422);
nor U34298 (N_34298,N_28409,N_28323);
xor U34299 (N_34299,N_25319,N_27174);
nand U34300 (N_34300,N_25526,N_28975);
nor U34301 (N_34301,N_29801,N_29937);
or U34302 (N_34302,N_28608,N_28781);
nor U34303 (N_34303,N_29414,N_26806);
nand U34304 (N_34304,N_28054,N_28700);
and U34305 (N_34305,N_29636,N_26235);
or U34306 (N_34306,N_29655,N_29463);
nand U34307 (N_34307,N_25359,N_25277);
or U34308 (N_34308,N_28451,N_27286);
nand U34309 (N_34309,N_28702,N_27836);
and U34310 (N_34310,N_26404,N_28978);
xor U34311 (N_34311,N_29064,N_25723);
and U34312 (N_34312,N_25358,N_29606);
and U34313 (N_34313,N_26237,N_28239);
xnor U34314 (N_34314,N_29934,N_26708);
nor U34315 (N_34315,N_28878,N_29021);
nor U34316 (N_34316,N_29944,N_26898);
nor U34317 (N_34317,N_28244,N_29375);
nand U34318 (N_34318,N_25619,N_27040);
or U34319 (N_34319,N_28473,N_29489);
xor U34320 (N_34320,N_27552,N_26630);
and U34321 (N_34321,N_25917,N_28366);
xnor U34322 (N_34322,N_28203,N_27075);
nor U34323 (N_34323,N_26391,N_29679);
nor U34324 (N_34324,N_27397,N_26495);
xor U34325 (N_34325,N_29716,N_28154);
or U34326 (N_34326,N_27650,N_27503);
nor U34327 (N_34327,N_26058,N_27877);
and U34328 (N_34328,N_26437,N_26045);
and U34329 (N_34329,N_25748,N_28107);
nand U34330 (N_34330,N_25948,N_25645);
and U34331 (N_34331,N_29987,N_26965);
xnor U34332 (N_34332,N_25913,N_26622);
and U34333 (N_34333,N_25875,N_26461);
nor U34334 (N_34334,N_29523,N_28056);
or U34335 (N_34335,N_29842,N_29963);
or U34336 (N_34336,N_28173,N_27786);
xor U34337 (N_34337,N_27379,N_29654);
nor U34338 (N_34338,N_29169,N_29627);
nand U34339 (N_34339,N_26269,N_28925);
and U34340 (N_34340,N_28796,N_25167);
nor U34341 (N_34341,N_27408,N_27603);
or U34342 (N_34342,N_28919,N_25402);
and U34343 (N_34343,N_29077,N_26827);
nand U34344 (N_34344,N_28398,N_27648);
or U34345 (N_34345,N_26638,N_29061);
nand U34346 (N_34346,N_26618,N_25831);
nand U34347 (N_34347,N_29754,N_28905);
nor U34348 (N_34348,N_28321,N_25182);
and U34349 (N_34349,N_29068,N_25220);
nand U34350 (N_34350,N_25359,N_29831);
nor U34351 (N_34351,N_25601,N_28115);
nor U34352 (N_34352,N_26999,N_26369);
nor U34353 (N_34353,N_25441,N_28539);
or U34354 (N_34354,N_26052,N_28792);
xor U34355 (N_34355,N_25784,N_29228);
nor U34356 (N_34356,N_25091,N_25834);
and U34357 (N_34357,N_26539,N_29766);
or U34358 (N_34358,N_25060,N_27323);
or U34359 (N_34359,N_26562,N_28582);
nand U34360 (N_34360,N_29569,N_26939);
or U34361 (N_34361,N_28303,N_27414);
and U34362 (N_34362,N_26867,N_25055);
nand U34363 (N_34363,N_25891,N_25017);
or U34364 (N_34364,N_29890,N_25419);
or U34365 (N_34365,N_26500,N_28600);
or U34366 (N_34366,N_25708,N_26507);
nand U34367 (N_34367,N_25728,N_26342);
xor U34368 (N_34368,N_25592,N_29628);
and U34369 (N_34369,N_29151,N_27232);
xor U34370 (N_34370,N_27709,N_25130);
nor U34371 (N_34371,N_29815,N_28442);
or U34372 (N_34372,N_25280,N_28561);
and U34373 (N_34373,N_26743,N_27905);
nor U34374 (N_34374,N_25214,N_26839);
nor U34375 (N_34375,N_28115,N_29849);
xnor U34376 (N_34376,N_26849,N_28319);
or U34377 (N_34377,N_25657,N_28741);
nand U34378 (N_34378,N_26067,N_27443);
or U34379 (N_34379,N_25664,N_26638);
xor U34380 (N_34380,N_26526,N_28271);
nor U34381 (N_34381,N_25227,N_29142);
and U34382 (N_34382,N_29719,N_28932);
nor U34383 (N_34383,N_28461,N_26070);
nor U34384 (N_34384,N_25174,N_28588);
xor U34385 (N_34385,N_29452,N_25023);
or U34386 (N_34386,N_26514,N_29368);
xor U34387 (N_34387,N_28649,N_28359);
nand U34388 (N_34388,N_28476,N_29694);
or U34389 (N_34389,N_28159,N_27221);
and U34390 (N_34390,N_28128,N_28475);
nor U34391 (N_34391,N_29319,N_25081);
or U34392 (N_34392,N_25959,N_27036);
or U34393 (N_34393,N_26424,N_29477);
or U34394 (N_34394,N_25805,N_25057);
xor U34395 (N_34395,N_27894,N_28783);
nand U34396 (N_34396,N_25009,N_27151);
xor U34397 (N_34397,N_28115,N_27254);
or U34398 (N_34398,N_27238,N_29833);
nand U34399 (N_34399,N_28607,N_25717);
or U34400 (N_34400,N_26298,N_28903);
nor U34401 (N_34401,N_25981,N_29503);
and U34402 (N_34402,N_29232,N_26958);
or U34403 (N_34403,N_25668,N_27582);
or U34404 (N_34404,N_28554,N_29817);
nand U34405 (N_34405,N_25121,N_27569);
nor U34406 (N_34406,N_26809,N_26219);
xnor U34407 (N_34407,N_26394,N_27968);
nor U34408 (N_34408,N_26689,N_25198);
and U34409 (N_34409,N_25904,N_28201);
nand U34410 (N_34410,N_29642,N_26241);
nor U34411 (N_34411,N_26221,N_27250);
nor U34412 (N_34412,N_25830,N_29207);
nor U34413 (N_34413,N_27185,N_28194);
nor U34414 (N_34414,N_25290,N_27911);
or U34415 (N_34415,N_25383,N_27320);
xnor U34416 (N_34416,N_28492,N_29158);
xnor U34417 (N_34417,N_29882,N_27881);
xnor U34418 (N_34418,N_29423,N_29680);
nand U34419 (N_34419,N_26580,N_28982);
nor U34420 (N_34420,N_28135,N_25539);
xor U34421 (N_34421,N_25328,N_26979);
or U34422 (N_34422,N_27895,N_28551);
and U34423 (N_34423,N_27785,N_25197);
nor U34424 (N_34424,N_26315,N_28910);
or U34425 (N_34425,N_27103,N_27441);
xor U34426 (N_34426,N_27373,N_28599);
nor U34427 (N_34427,N_26835,N_29473);
xnor U34428 (N_34428,N_25998,N_29487);
and U34429 (N_34429,N_29420,N_29133);
xnor U34430 (N_34430,N_27971,N_28956);
nor U34431 (N_34431,N_29554,N_27474);
nand U34432 (N_34432,N_28510,N_29743);
nand U34433 (N_34433,N_26537,N_28576);
xnor U34434 (N_34434,N_27417,N_25829);
and U34435 (N_34435,N_27894,N_25133);
or U34436 (N_34436,N_26990,N_25301);
and U34437 (N_34437,N_26264,N_25787);
nand U34438 (N_34438,N_27950,N_29081);
xor U34439 (N_34439,N_29219,N_29214);
nand U34440 (N_34440,N_28672,N_29230);
or U34441 (N_34441,N_29111,N_28703);
or U34442 (N_34442,N_26468,N_25206);
xnor U34443 (N_34443,N_27828,N_27401);
and U34444 (N_34444,N_26164,N_28018);
xor U34445 (N_34445,N_26667,N_27112);
xor U34446 (N_34446,N_27935,N_27318);
xor U34447 (N_34447,N_25670,N_29825);
and U34448 (N_34448,N_25525,N_27849);
xor U34449 (N_34449,N_25146,N_25421);
nor U34450 (N_34450,N_27771,N_25311);
xor U34451 (N_34451,N_27085,N_28198);
or U34452 (N_34452,N_26388,N_28855);
xnor U34453 (N_34453,N_26441,N_29639);
nor U34454 (N_34454,N_27528,N_26230);
nor U34455 (N_34455,N_27177,N_25686);
nand U34456 (N_34456,N_29662,N_25927);
nor U34457 (N_34457,N_26166,N_27958);
or U34458 (N_34458,N_27447,N_27654);
nor U34459 (N_34459,N_25918,N_25197);
and U34460 (N_34460,N_29096,N_28309);
and U34461 (N_34461,N_27319,N_26987);
nor U34462 (N_34462,N_29178,N_26659);
and U34463 (N_34463,N_28505,N_29958);
and U34464 (N_34464,N_25169,N_26697);
nor U34465 (N_34465,N_29689,N_26861);
nand U34466 (N_34466,N_29015,N_28457);
or U34467 (N_34467,N_28956,N_28038);
nor U34468 (N_34468,N_25701,N_29920);
nor U34469 (N_34469,N_28978,N_26187);
xnor U34470 (N_34470,N_29865,N_28604);
xnor U34471 (N_34471,N_29124,N_26515);
or U34472 (N_34472,N_25757,N_28910);
or U34473 (N_34473,N_28291,N_25753);
or U34474 (N_34474,N_25851,N_29289);
and U34475 (N_34475,N_29093,N_27987);
nor U34476 (N_34476,N_28140,N_25902);
xnor U34477 (N_34477,N_27758,N_29541);
nor U34478 (N_34478,N_26833,N_26229);
or U34479 (N_34479,N_28672,N_27122);
xor U34480 (N_34480,N_26869,N_28152);
xnor U34481 (N_34481,N_29292,N_27370);
nor U34482 (N_34482,N_29185,N_28983);
and U34483 (N_34483,N_27495,N_29606);
xnor U34484 (N_34484,N_26538,N_26862);
or U34485 (N_34485,N_26306,N_26509);
and U34486 (N_34486,N_25628,N_27474);
and U34487 (N_34487,N_25742,N_28362);
nand U34488 (N_34488,N_25348,N_25724);
nand U34489 (N_34489,N_27244,N_25026);
nor U34490 (N_34490,N_28261,N_25424);
and U34491 (N_34491,N_28396,N_28792);
nor U34492 (N_34492,N_29624,N_26999);
and U34493 (N_34493,N_25899,N_28313);
or U34494 (N_34494,N_26756,N_26488);
xnor U34495 (N_34495,N_28453,N_26633);
or U34496 (N_34496,N_28964,N_27102);
nor U34497 (N_34497,N_26890,N_27591);
or U34498 (N_34498,N_25066,N_28095);
nor U34499 (N_34499,N_26889,N_28323);
and U34500 (N_34500,N_27336,N_29173);
nor U34501 (N_34501,N_25199,N_25213);
or U34502 (N_34502,N_29960,N_25597);
or U34503 (N_34503,N_26189,N_26035);
nor U34504 (N_34504,N_26732,N_25723);
or U34505 (N_34505,N_28596,N_27397);
nor U34506 (N_34506,N_25218,N_29479);
xor U34507 (N_34507,N_28053,N_28424);
nand U34508 (N_34508,N_29011,N_29611);
or U34509 (N_34509,N_27586,N_25805);
or U34510 (N_34510,N_25594,N_26366);
nand U34511 (N_34511,N_28236,N_26878);
or U34512 (N_34512,N_27227,N_25463);
nand U34513 (N_34513,N_26300,N_26735);
xor U34514 (N_34514,N_27360,N_28968);
or U34515 (N_34515,N_25645,N_27305);
xor U34516 (N_34516,N_27183,N_27489);
and U34517 (N_34517,N_27356,N_26229);
or U34518 (N_34518,N_26630,N_26998);
nand U34519 (N_34519,N_29927,N_28783);
or U34520 (N_34520,N_29246,N_26198);
xnor U34521 (N_34521,N_27621,N_27212);
xnor U34522 (N_34522,N_27091,N_25890);
nor U34523 (N_34523,N_27090,N_29720);
xnor U34524 (N_34524,N_27638,N_27600);
nor U34525 (N_34525,N_28246,N_25837);
nor U34526 (N_34526,N_26089,N_25187);
nand U34527 (N_34527,N_28962,N_27328);
nor U34528 (N_34528,N_26764,N_27053);
nand U34529 (N_34529,N_28470,N_27232);
nor U34530 (N_34530,N_25570,N_26299);
and U34531 (N_34531,N_26059,N_27143);
nand U34532 (N_34532,N_26586,N_28440);
nor U34533 (N_34533,N_29348,N_29738);
or U34534 (N_34534,N_28358,N_27915);
or U34535 (N_34535,N_26238,N_27704);
xor U34536 (N_34536,N_25517,N_26623);
xnor U34537 (N_34537,N_27438,N_25456);
xnor U34538 (N_34538,N_27984,N_26607);
or U34539 (N_34539,N_26112,N_28710);
or U34540 (N_34540,N_26821,N_29570);
xor U34541 (N_34541,N_26255,N_29213);
nand U34542 (N_34542,N_25796,N_29074);
and U34543 (N_34543,N_25833,N_27696);
or U34544 (N_34544,N_27044,N_26176);
nor U34545 (N_34545,N_27638,N_25896);
or U34546 (N_34546,N_29168,N_25449);
nor U34547 (N_34547,N_26987,N_29260);
nand U34548 (N_34548,N_28012,N_29074);
and U34549 (N_34549,N_28464,N_27613);
xor U34550 (N_34550,N_28206,N_29994);
nor U34551 (N_34551,N_29297,N_26428);
nor U34552 (N_34552,N_25602,N_29710);
xor U34553 (N_34553,N_28394,N_27229);
nor U34554 (N_34554,N_25609,N_25414);
and U34555 (N_34555,N_29466,N_25054);
nor U34556 (N_34556,N_26397,N_25015);
xnor U34557 (N_34557,N_28123,N_28062);
or U34558 (N_34558,N_25026,N_26685);
nand U34559 (N_34559,N_25281,N_28352);
nand U34560 (N_34560,N_28787,N_27112);
nand U34561 (N_34561,N_26552,N_25488);
or U34562 (N_34562,N_27345,N_28723);
xor U34563 (N_34563,N_28096,N_27633);
and U34564 (N_34564,N_26389,N_27730);
xnor U34565 (N_34565,N_26609,N_25167);
or U34566 (N_34566,N_28414,N_27848);
nand U34567 (N_34567,N_27093,N_29448);
or U34568 (N_34568,N_27705,N_28451);
or U34569 (N_34569,N_29055,N_27634);
and U34570 (N_34570,N_28740,N_25935);
or U34571 (N_34571,N_27182,N_25472);
xor U34572 (N_34572,N_29941,N_25736);
xor U34573 (N_34573,N_29006,N_27590);
and U34574 (N_34574,N_26431,N_29811);
xor U34575 (N_34575,N_25759,N_27768);
nor U34576 (N_34576,N_27075,N_29366);
nor U34577 (N_34577,N_26827,N_29344);
nor U34578 (N_34578,N_25956,N_27033);
nand U34579 (N_34579,N_29707,N_28360);
and U34580 (N_34580,N_28996,N_26893);
xor U34581 (N_34581,N_28500,N_26731);
xor U34582 (N_34582,N_26109,N_25303);
or U34583 (N_34583,N_28573,N_29378);
nand U34584 (N_34584,N_28222,N_27163);
nor U34585 (N_34585,N_28810,N_25927);
xor U34586 (N_34586,N_28452,N_28060);
nor U34587 (N_34587,N_26102,N_27025);
nor U34588 (N_34588,N_25373,N_26033);
nand U34589 (N_34589,N_26086,N_26392);
nor U34590 (N_34590,N_27246,N_28720);
or U34591 (N_34591,N_26912,N_29599);
nor U34592 (N_34592,N_25712,N_28344);
or U34593 (N_34593,N_25418,N_29385);
or U34594 (N_34594,N_29096,N_28678);
nor U34595 (N_34595,N_26612,N_25366);
xnor U34596 (N_34596,N_25802,N_29338);
nor U34597 (N_34597,N_29387,N_26610);
and U34598 (N_34598,N_28842,N_25741);
nand U34599 (N_34599,N_25421,N_29836);
or U34600 (N_34600,N_29110,N_29820);
nand U34601 (N_34601,N_28795,N_26965);
and U34602 (N_34602,N_26459,N_29555);
xor U34603 (N_34603,N_28426,N_26647);
nand U34604 (N_34604,N_26679,N_27937);
nor U34605 (N_34605,N_27086,N_28775);
nand U34606 (N_34606,N_29014,N_26798);
nor U34607 (N_34607,N_29084,N_27514);
nand U34608 (N_34608,N_28278,N_29571);
nor U34609 (N_34609,N_28453,N_27813);
nand U34610 (N_34610,N_27960,N_28719);
nor U34611 (N_34611,N_29364,N_25777);
nor U34612 (N_34612,N_27785,N_28685);
xor U34613 (N_34613,N_25917,N_29686);
xor U34614 (N_34614,N_25968,N_27664);
nor U34615 (N_34615,N_27058,N_29973);
nand U34616 (N_34616,N_27170,N_26084);
nor U34617 (N_34617,N_25995,N_29871);
and U34618 (N_34618,N_27412,N_26576);
xor U34619 (N_34619,N_27082,N_28728);
nor U34620 (N_34620,N_25616,N_27773);
nand U34621 (N_34621,N_27505,N_28738);
or U34622 (N_34622,N_25553,N_29653);
nand U34623 (N_34623,N_26729,N_28697);
and U34624 (N_34624,N_28842,N_26810);
and U34625 (N_34625,N_26577,N_28197);
or U34626 (N_34626,N_27023,N_28763);
xnor U34627 (N_34627,N_28575,N_25861);
nor U34628 (N_34628,N_26591,N_27934);
nand U34629 (N_34629,N_28325,N_25578);
nand U34630 (N_34630,N_29088,N_25749);
or U34631 (N_34631,N_25992,N_28103);
or U34632 (N_34632,N_26409,N_25615);
xnor U34633 (N_34633,N_25864,N_25740);
or U34634 (N_34634,N_26066,N_28200);
nand U34635 (N_34635,N_25719,N_26494);
nor U34636 (N_34636,N_28297,N_27689);
xor U34637 (N_34637,N_28478,N_26477);
and U34638 (N_34638,N_27480,N_29271);
xnor U34639 (N_34639,N_27477,N_26343);
or U34640 (N_34640,N_25683,N_26613);
or U34641 (N_34641,N_25626,N_27498);
or U34642 (N_34642,N_25287,N_28195);
nor U34643 (N_34643,N_28552,N_26118);
xnor U34644 (N_34644,N_27098,N_28351);
and U34645 (N_34645,N_27222,N_29229);
xnor U34646 (N_34646,N_25993,N_26360);
and U34647 (N_34647,N_29173,N_29711);
xor U34648 (N_34648,N_29161,N_28262);
and U34649 (N_34649,N_27684,N_26411);
or U34650 (N_34650,N_29016,N_28005);
or U34651 (N_34651,N_25620,N_29516);
nand U34652 (N_34652,N_27618,N_28421);
nor U34653 (N_34653,N_29054,N_27064);
or U34654 (N_34654,N_29443,N_26065);
nor U34655 (N_34655,N_26504,N_29921);
nor U34656 (N_34656,N_25471,N_26109);
and U34657 (N_34657,N_28111,N_28993);
or U34658 (N_34658,N_26274,N_29688);
nor U34659 (N_34659,N_26172,N_28431);
nor U34660 (N_34660,N_27236,N_25703);
and U34661 (N_34661,N_26305,N_25905);
and U34662 (N_34662,N_25091,N_28241);
nor U34663 (N_34663,N_27106,N_28399);
nor U34664 (N_34664,N_25766,N_29873);
or U34665 (N_34665,N_27027,N_25865);
or U34666 (N_34666,N_28596,N_29262);
nor U34667 (N_34667,N_25122,N_26788);
and U34668 (N_34668,N_28821,N_27452);
nor U34669 (N_34669,N_27351,N_28897);
nor U34670 (N_34670,N_26447,N_27751);
xor U34671 (N_34671,N_28455,N_25537);
nand U34672 (N_34672,N_27783,N_28801);
nor U34673 (N_34673,N_28492,N_28302);
or U34674 (N_34674,N_29784,N_25098);
and U34675 (N_34675,N_28463,N_28299);
and U34676 (N_34676,N_26388,N_29217);
or U34677 (N_34677,N_26193,N_28128);
nand U34678 (N_34678,N_29947,N_29246);
nor U34679 (N_34679,N_29498,N_26326);
and U34680 (N_34680,N_27135,N_29993);
xnor U34681 (N_34681,N_28880,N_29663);
nor U34682 (N_34682,N_26419,N_27510);
and U34683 (N_34683,N_28819,N_27134);
or U34684 (N_34684,N_25858,N_27826);
or U34685 (N_34685,N_29036,N_26251);
or U34686 (N_34686,N_26952,N_26035);
nor U34687 (N_34687,N_25301,N_27877);
nor U34688 (N_34688,N_27017,N_27898);
nor U34689 (N_34689,N_25564,N_29140);
or U34690 (N_34690,N_27438,N_27640);
xnor U34691 (N_34691,N_27086,N_25500);
or U34692 (N_34692,N_27037,N_25667);
nand U34693 (N_34693,N_25277,N_26714);
and U34694 (N_34694,N_29765,N_29423);
xor U34695 (N_34695,N_25504,N_25012);
nor U34696 (N_34696,N_26139,N_29366);
and U34697 (N_34697,N_25777,N_25467);
and U34698 (N_34698,N_25481,N_27147);
xnor U34699 (N_34699,N_25031,N_28167);
and U34700 (N_34700,N_29993,N_29795);
nor U34701 (N_34701,N_26537,N_26190);
and U34702 (N_34702,N_28508,N_29537);
or U34703 (N_34703,N_25747,N_27168);
xnor U34704 (N_34704,N_27392,N_25603);
xor U34705 (N_34705,N_28713,N_25475);
nor U34706 (N_34706,N_25900,N_28517);
nand U34707 (N_34707,N_27636,N_26523);
xnor U34708 (N_34708,N_28708,N_26650);
and U34709 (N_34709,N_29716,N_28630);
nand U34710 (N_34710,N_27157,N_26073);
nor U34711 (N_34711,N_27812,N_25378);
or U34712 (N_34712,N_25148,N_26674);
xnor U34713 (N_34713,N_26927,N_28808);
or U34714 (N_34714,N_28756,N_25593);
nand U34715 (N_34715,N_26410,N_29184);
nor U34716 (N_34716,N_26566,N_27834);
nand U34717 (N_34717,N_27420,N_27461);
nand U34718 (N_34718,N_28182,N_26984);
or U34719 (N_34719,N_25876,N_26433);
nor U34720 (N_34720,N_26992,N_26852);
and U34721 (N_34721,N_25588,N_29071);
or U34722 (N_34722,N_29125,N_29994);
nand U34723 (N_34723,N_29719,N_27698);
or U34724 (N_34724,N_28875,N_26780);
xnor U34725 (N_34725,N_29053,N_26554);
nor U34726 (N_34726,N_28378,N_25760);
nand U34727 (N_34727,N_27766,N_25815);
nand U34728 (N_34728,N_25021,N_29608);
nor U34729 (N_34729,N_28445,N_26849);
or U34730 (N_34730,N_29998,N_25711);
or U34731 (N_34731,N_26295,N_29235);
and U34732 (N_34732,N_29139,N_29818);
and U34733 (N_34733,N_25517,N_25996);
or U34734 (N_34734,N_27382,N_27669);
nor U34735 (N_34735,N_26024,N_29015);
or U34736 (N_34736,N_26899,N_25355);
xor U34737 (N_34737,N_29462,N_28172);
nand U34738 (N_34738,N_29491,N_25016);
or U34739 (N_34739,N_29123,N_25086);
nor U34740 (N_34740,N_29817,N_28387);
or U34741 (N_34741,N_29833,N_26315);
nor U34742 (N_34742,N_27767,N_29955);
or U34743 (N_34743,N_25612,N_27792);
xor U34744 (N_34744,N_28487,N_26182);
or U34745 (N_34745,N_26407,N_27704);
nand U34746 (N_34746,N_26420,N_28840);
and U34747 (N_34747,N_29977,N_29737);
or U34748 (N_34748,N_26608,N_28362);
and U34749 (N_34749,N_27167,N_26750);
and U34750 (N_34750,N_29832,N_26680);
and U34751 (N_34751,N_26199,N_26068);
xor U34752 (N_34752,N_27133,N_26014);
and U34753 (N_34753,N_27521,N_26037);
nor U34754 (N_34754,N_25259,N_28588);
or U34755 (N_34755,N_25582,N_27686);
or U34756 (N_34756,N_28345,N_29879);
and U34757 (N_34757,N_29327,N_29783);
xnor U34758 (N_34758,N_27604,N_27680);
xor U34759 (N_34759,N_26566,N_26559);
and U34760 (N_34760,N_28142,N_26755);
or U34761 (N_34761,N_26558,N_25745);
nand U34762 (N_34762,N_29960,N_26927);
nand U34763 (N_34763,N_28218,N_29987);
and U34764 (N_34764,N_26294,N_25419);
nand U34765 (N_34765,N_28536,N_29303);
and U34766 (N_34766,N_25912,N_27821);
or U34767 (N_34767,N_29395,N_28684);
or U34768 (N_34768,N_25537,N_29378);
and U34769 (N_34769,N_26234,N_28977);
and U34770 (N_34770,N_29387,N_28449);
and U34771 (N_34771,N_27241,N_28946);
and U34772 (N_34772,N_26688,N_26609);
and U34773 (N_34773,N_27303,N_28775);
nand U34774 (N_34774,N_25615,N_28877);
nor U34775 (N_34775,N_29203,N_29306);
nor U34776 (N_34776,N_27796,N_25331);
nor U34777 (N_34777,N_27246,N_26975);
nand U34778 (N_34778,N_26316,N_25213);
nand U34779 (N_34779,N_26441,N_25025);
and U34780 (N_34780,N_28745,N_29510);
nor U34781 (N_34781,N_26576,N_28747);
nand U34782 (N_34782,N_27412,N_28743);
nor U34783 (N_34783,N_26069,N_29494);
or U34784 (N_34784,N_27626,N_28330);
or U34785 (N_34785,N_26477,N_26868);
nand U34786 (N_34786,N_28442,N_29712);
nand U34787 (N_34787,N_29232,N_25805);
xnor U34788 (N_34788,N_27688,N_25515);
or U34789 (N_34789,N_25010,N_27493);
or U34790 (N_34790,N_27264,N_29071);
nor U34791 (N_34791,N_25312,N_25384);
nand U34792 (N_34792,N_28575,N_25390);
nand U34793 (N_34793,N_29692,N_28684);
or U34794 (N_34794,N_29420,N_26055);
nand U34795 (N_34795,N_28041,N_28436);
nand U34796 (N_34796,N_26614,N_29621);
nand U34797 (N_34797,N_25193,N_28594);
and U34798 (N_34798,N_26222,N_26270);
and U34799 (N_34799,N_26161,N_28258);
or U34800 (N_34800,N_26169,N_25814);
nor U34801 (N_34801,N_27221,N_27528);
xor U34802 (N_34802,N_27342,N_27614);
xnor U34803 (N_34803,N_27931,N_27700);
nand U34804 (N_34804,N_29065,N_29696);
nor U34805 (N_34805,N_25760,N_26065);
xnor U34806 (N_34806,N_25924,N_28002);
nor U34807 (N_34807,N_28742,N_29966);
nand U34808 (N_34808,N_27852,N_26994);
nor U34809 (N_34809,N_25408,N_26953);
or U34810 (N_34810,N_27898,N_25914);
nand U34811 (N_34811,N_27556,N_29054);
or U34812 (N_34812,N_25642,N_29794);
or U34813 (N_34813,N_29671,N_26931);
nand U34814 (N_34814,N_28213,N_26598);
xnor U34815 (N_34815,N_27044,N_29571);
and U34816 (N_34816,N_25261,N_27187);
nand U34817 (N_34817,N_26160,N_26655);
or U34818 (N_34818,N_29586,N_27291);
and U34819 (N_34819,N_27432,N_29655);
nand U34820 (N_34820,N_27784,N_27915);
nor U34821 (N_34821,N_28026,N_29493);
and U34822 (N_34822,N_28509,N_26214);
nand U34823 (N_34823,N_27697,N_28898);
and U34824 (N_34824,N_25384,N_29553);
xor U34825 (N_34825,N_29073,N_28167);
nor U34826 (N_34826,N_26958,N_25049);
nor U34827 (N_34827,N_25197,N_26023);
and U34828 (N_34828,N_29343,N_25035);
nor U34829 (N_34829,N_29869,N_26836);
xnor U34830 (N_34830,N_25113,N_29859);
nand U34831 (N_34831,N_26743,N_26805);
and U34832 (N_34832,N_25547,N_29680);
nand U34833 (N_34833,N_25908,N_26839);
xnor U34834 (N_34834,N_26792,N_29335);
xor U34835 (N_34835,N_25550,N_29513);
or U34836 (N_34836,N_26508,N_26582);
nor U34837 (N_34837,N_28434,N_25310);
and U34838 (N_34838,N_25729,N_27793);
nor U34839 (N_34839,N_26677,N_26404);
or U34840 (N_34840,N_29636,N_28617);
and U34841 (N_34841,N_27807,N_25978);
nand U34842 (N_34842,N_25001,N_28758);
nor U34843 (N_34843,N_27934,N_28640);
nor U34844 (N_34844,N_27131,N_26514);
or U34845 (N_34845,N_26758,N_26481);
nand U34846 (N_34846,N_26068,N_25481);
xnor U34847 (N_34847,N_25721,N_27200);
and U34848 (N_34848,N_27147,N_26272);
and U34849 (N_34849,N_25007,N_29291);
and U34850 (N_34850,N_25698,N_25936);
nor U34851 (N_34851,N_29529,N_27710);
nor U34852 (N_34852,N_29839,N_27172);
nor U34853 (N_34853,N_27251,N_26096);
nor U34854 (N_34854,N_28127,N_25761);
and U34855 (N_34855,N_25786,N_26040);
xor U34856 (N_34856,N_26271,N_28250);
xnor U34857 (N_34857,N_27998,N_28463);
or U34858 (N_34858,N_29733,N_26473);
nand U34859 (N_34859,N_29174,N_27303);
xor U34860 (N_34860,N_29244,N_26809);
or U34861 (N_34861,N_29717,N_27347);
nand U34862 (N_34862,N_28125,N_27709);
xnor U34863 (N_34863,N_27551,N_26067);
nand U34864 (N_34864,N_28380,N_29819);
xnor U34865 (N_34865,N_27192,N_26922);
or U34866 (N_34866,N_27144,N_26391);
and U34867 (N_34867,N_27914,N_28059);
nand U34868 (N_34868,N_29400,N_26139);
and U34869 (N_34869,N_26989,N_26297);
nand U34870 (N_34870,N_28763,N_26142);
nor U34871 (N_34871,N_25998,N_25174);
xnor U34872 (N_34872,N_25880,N_29541);
and U34873 (N_34873,N_28125,N_29946);
or U34874 (N_34874,N_27695,N_29103);
xor U34875 (N_34875,N_25664,N_28043);
and U34876 (N_34876,N_28710,N_29930);
nand U34877 (N_34877,N_27488,N_29147);
nor U34878 (N_34878,N_27619,N_28466);
or U34879 (N_34879,N_29251,N_27283);
and U34880 (N_34880,N_29013,N_28958);
and U34881 (N_34881,N_28900,N_27632);
xor U34882 (N_34882,N_28652,N_25569);
nor U34883 (N_34883,N_26789,N_27850);
and U34884 (N_34884,N_28596,N_25929);
and U34885 (N_34885,N_27786,N_26324);
and U34886 (N_34886,N_28628,N_26736);
nand U34887 (N_34887,N_25280,N_29793);
and U34888 (N_34888,N_25313,N_27808);
nor U34889 (N_34889,N_29800,N_28150);
nand U34890 (N_34890,N_28799,N_28825);
nand U34891 (N_34891,N_25185,N_25005);
nand U34892 (N_34892,N_29940,N_29927);
nor U34893 (N_34893,N_29549,N_25549);
xnor U34894 (N_34894,N_29399,N_25451);
nand U34895 (N_34895,N_26077,N_26831);
or U34896 (N_34896,N_27150,N_27369);
or U34897 (N_34897,N_27716,N_28804);
nand U34898 (N_34898,N_26145,N_28807);
nor U34899 (N_34899,N_27250,N_26712);
xnor U34900 (N_34900,N_28419,N_26475);
nor U34901 (N_34901,N_26273,N_26313);
or U34902 (N_34902,N_26035,N_28134);
and U34903 (N_34903,N_26171,N_28897);
nand U34904 (N_34904,N_27624,N_27394);
nor U34905 (N_34905,N_29693,N_26842);
and U34906 (N_34906,N_25605,N_26510);
nand U34907 (N_34907,N_29279,N_25226);
nor U34908 (N_34908,N_25839,N_28834);
nand U34909 (N_34909,N_28759,N_29032);
nor U34910 (N_34910,N_27240,N_26571);
nor U34911 (N_34911,N_27507,N_27424);
and U34912 (N_34912,N_27934,N_28889);
xnor U34913 (N_34913,N_28671,N_29299);
xor U34914 (N_34914,N_26800,N_26462);
and U34915 (N_34915,N_27712,N_29766);
xor U34916 (N_34916,N_27977,N_26382);
xor U34917 (N_34917,N_26957,N_28582);
nor U34918 (N_34918,N_27208,N_28846);
or U34919 (N_34919,N_25588,N_29553);
nor U34920 (N_34920,N_28699,N_27054);
nand U34921 (N_34921,N_29598,N_25544);
or U34922 (N_34922,N_28525,N_25721);
and U34923 (N_34923,N_27418,N_28201);
and U34924 (N_34924,N_28984,N_25486);
nand U34925 (N_34925,N_28030,N_28686);
and U34926 (N_34926,N_27676,N_29067);
and U34927 (N_34927,N_25539,N_26998);
nand U34928 (N_34928,N_29434,N_25313);
and U34929 (N_34929,N_28474,N_29538);
nor U34930 (N_34930,N_26648,N_29283);
nand U34931 (N_34931,N_25354,N_27830);
nor U34932 (N_34932,N_27048,N_27442);
nand U34933 (N_34933,N_28554,N_26730);
nand U34934 (N_34934,N_28530,N_27174);
xor U34935 (N_34935,N_29870,N_28644);
and U34936 (N_34936,N_28389,N_26725);
or U34937 (N_34937,N_25120,N_26439);
xnor U34938 (N_34938,N_27212,N_29078);
nand U34939 (N_34939,N_29986,N_27285);
nor U34940 (N_34940,N_28149,N_27200);
and U34941 (N_34941,N_27317,N_29758);
nor U34942 (N_34942,N_28322,N_26037);
and U34943 (N_34943,N_28529,N_29600);
nor U34944 (N_34944,N_27940,N_25824);
nand U34945 (N_34945,N_29013,N_28663);
xnor U34946 (N_34946,N_25679,N_27492);
nand U34947 (N_34947,N_28510,N_27994);
or U34948 (N_34948,N_28293,N_25820);
nand U34949 (N_34949,N_26979,N_29159);
and U34950 (N_34950,N_27930,N_29469);
nor U34951 (N_34951,N_26126,N_26783);
and U34952 (N_34952,N_25985,N_25499);
nor U34953 (N_34953,N_27695,N_26550);
nor U34954 (N_34954,N_29513,N_26047);
nor U34955 (N_34955,N_26142,N_29428);
nand U34956 (N_34956,N_26240,N_28058);
or U34957 (N_34957,N_27171,N_26579);
nor U34958 (N_34958,N_26398,N_29289);
nor U34959 (N_34959,N_25441,N_26457);
and U34960 (N_34960,N_26483,N_27999);
nand U34961 (N_34961,N_25194,N_26565);
or U34962 (N_34962,N_28044,N_25367);
or U34963 (N_34963,N_29379,N_27850);
and U34964 (N_34964,N_25230,N_26658);
nor U34965 (N_34965,N_28033,N_26021);
nand U34966 (N_34966,N_27685,N_25514);
or U34967 (N_34967,N_29560,N_27453);
nand U34968 (N_34968,N_27279,N_28267);
or U34969 (N_34969,N_26072,N_29066);
nor U34970 (N_34970,N_28423,N_29404);
or U34971 (N_34971,N_26926,N_27045);
nor U34972 (N_34972,N_25130,N_26614);
or U34973 (N_34973,N_25537,N_28041);
and U34974 (N_34974,N_27012,N_27306);
and U34975 (N_34975,N_29469,N_28583);
nand U34976 (N_34976,N_29139,N_27453);
nor U34977 (N_34977,N_25419,N_29903);
nand U34978 (N_34978,N_27751,N_28617);
nor U34979 (N_34979,N_26323,N_28203);
nor U34980 (N_34980,N_26266,N_25413);
nand U34981 (N_34981,N_29840,N_28701);
nor U34982 (N_34982,N_27165,N_29906);
nor U34983 (N_34983,N_26938,N_29047);
nor U34984 (N_34984,N_25464,N_29502);
xnor U34985 (N_34985,N_27704,N_29259);
xor U34986 (N_34986,N_25136,N_26923);
or U34987 (N_34987,N_25832,N_28117);
xor U34988 (N_34988,N_27058,N_27277);
and U34989 (N_34989,N_25116,N_28411);
nand U34990 (N_34990,N_26060,N_27863);
nor U34991 (N_34991,N_28815,N_26401);
xnor U34992 (N_34992,N_29805,N_26590);
or U34993 (N_34993,N_25196,N_28794);
or U34994 (N_34994,N_28586,N_29043);
nor U34995 (N_34995,N_28231,N_28363);
and U34996 (N_34996,N_28238,N_28208);
and U34997 (N_34997,N_29226,N_29765);
and U34998 (N_34998,N_29001,N_28891);
nor U34999 (N_34999,N_27701,N_25169);
nor U35000 (N_35000,N_33487,N_34781);
or U35001 (N_35001,N_32491,N_33935);
and U35002 (N_35002,N_33477,N_33529);
or U35003 (N_35003,N_34010,N_32121);
xnor U35004 (N_35004,N_30177,N_34114);
nand U35005 (N_35005,N_31402,N_30979);
and U35006 (N_35006,N_31460,N_34386);
xnor U35007 (N_35007,N_33343,N_33733);
nor U35008 (N_35008,N_30175,N_34275);
nand U35009 (N_35009,N_33514,N_32253);
nor U35010 (N_35010,N_30704,N_32228);
and U35011 (N_35011,N_31513,N_30949);
nor U35012 (N_35012,N_34039,N_32544);
xor U35013 (N_35013,N_30315,N_34589);
xor U35014 (N_35014,N_31614,N_32799);
nor U35015 (N_35015,N_32440,N_32419);
nand U35016 (N_35016,N_31338,N_34471);
or U35017 (N_35017,N_31933,N_32294);
nand U35018 (N_35018,N_30489,N_31824);
or U35019 (N_35019,N_33555,N_32211);
xnor U35020 (N_35020,N_31068,N_33114);
nor U35021 (N_35021,N_34168,N_30098);
or U35022 (N_35022,N_31527,N_30256);
xnor U35023 (N_35023,N_32263,N_34080);
nor U35024 (N_35024,N_31094,N_33246);
or U35025 (N_35025,N_31605,N_30673);
nand U35026 (N_35026,N_31406,N_31167);
or U35027 (N_35027,N_30061,N_30806);
and U35028 (N_35028,N_32155,N_33568);
xor U35029 (N_35029,N_33040,N_30487);
nor U35030 (N_35030,N_32282,N_32423);
nor U35031 (N_35031,N_32171,N_31198);
nand U35032 (N_35032,N_30263,N_32026);
xnor U35033 (N_35033,N_34561,N_34276);
or U35034 (N_35034,N_31316,N_31024);
nor U35035 (N_35035,N_30616,N_34366);
nor U35036 (N_35036,N_33738,N_33802);
xnor U35037 (N_35037,N_31514,N_31496);
or U35038 (N_35038,N_32050,N_34250);
and U35039 (N_35039,N_34164,N_31874);
and U35040 (N_35040,N_31903,N_30261);
nand U35041 (N_35041,N_32901,N_33362);
nand U35042 (N_35042,N_32929,N_32495);
or U35043 (N_35043,N_32378,N_31948);
nor U35044 (N_35044,N_32967,N_30351);
nor U35045 (N_35045,N_34880,N_32140);
xnor U35046 (N_35046,N_32503,N_31458);
xnor U35047 (N_35047,N_33181,N_34462);
or U35048 (N_35048,N_31571,N_34488);
and U35049 (N_35049,N_34290,N_34450);
or U35050 (N_35050,N_32324,N_30355);
and U35051 (N_35051,N_34554,N_33298);
and U35052 (N_35052,N_33843,N_30820);
xnor U35053 (N_35053,N_32173,N_30571);
nand U35054 (N_35054,N_33563,N_33744);
and U35055 (N_35055,N_30938,N_31967);
and U35056 (N_35056,N_33020,N_30448);
nor U35057 (N_35057,N_31492,N_31588);
nor U35058 (N_35058,N_34515,N_33695);
nand U35059 (N_35059,N_34750,N_32974);
and U35060 (N_35060,N_32911,N_32906);
xor U35061 (N_35061,N_30718,N_30206);
and U35062 (N_35062,N_31585,N_31825);
or U35063 (N_35063,N_30857,N_32604);
nand U35064 (N_35064,N_30409,N_32592);
nor U35065 (N_35065,N_31762,N_34329);
xor U35066 (N_35066,N_33168,N_32156);
and U35067 (N_35067,N_33091,N_33082);
and U35068 (N_35068,N_32972,N_32144);
nor U35069 (N_35069,N_32307,N_30877);
or U35070 (N_35070,N_34459,N_30163);
nor U35071 (N_35071,N_34719,N_31976);
xnor U35072 (N_35072,N_30179,N_34659);
xor U35073 (N_35073,N_33857,N_32420);
or U35074 (N_35074,N_34716,N_33513);
nand U35075 (N_35075,N_31204,N_32267);
nand U35076 (N_35076,N_33814,N_30278);
xor U35077 (N_35077,N_31386,N_32855);
xor U35078 (N_35078,N_31367,N_31147);
xor U35079 (N_35079,N_34444,N_32193);
xnor U35080 (N_35080,N_31251,N_34272);
nand U35081 (N_35081,N_30195,N_33894);
nor U35082 (N_35082,N_33560,N_31922);
nand U35083 (N_35083,N_31802,N_31589);
nand U35084 (N_35084,N_31451,N_34738);
nor U35085 (N_35085,N_32329,N_32347);
or U35086 (N_35086,N_32470,N_31784);
or U35087 (N_35087,N_30425,N_32997);
xnor U35088 (N_35088,N_31454,N_32196);
nor U35089 (N_35089,N_31950,N_30491);
or U35090 (N_35090,N_33888,N_33337);
and U35091 (N_35091,N_31593,N_30105);
nand U35092 (N_35092,N_30659,N_34348);
or U35093 (N_35093,N_31273,N_33134);
or U35094 (N_35094,N_31708,N_33724);
xnor U35095 (N_35095,N_30400,N_32838);
nand U35096 (N_35096,N_33904,N_30481);
nor U35097 (N_35097,N_33103,N_31537);
xnor U35098 (N_35098,N_31243,N_30010);
xor U35099 (N_35099,N_34063,N_33579);
or U35100 (N_35100,N_34306,N_33628);
or U35101 (N_35101,N_33455,N_31403);
and U35102 (N_35102,N_34445,N_31932);
nor U35103 (N_35103,N_32526,N_30232);
or U35104 (N_35104,N_30238,N_30744);
nor U35105 (N_35105,N_30672,N_32444);
or U35106 (N_35106,N_31020,N_33086);
xnor U35107 (N_35107,N_33672,N_31072);
nand U35108 (N_35108,N_30036,N_31782);
and U35109 (N_35109,N_30260,N_30053);
xor U35110 (N_35110,N_33898,N_32953);
and U35111 (N_35111,N_33216,N_30348);
or U35112 (N_35112,N_33361,N_31547);
or U35113 (N_35113,N_32414,N_33196);
or U35114 (N_35114,N_31796,N_33536);
nor U35115 (N_35115,N_32142,N_31392);
or U35116 (N_35116,N_30711,N_32475);
or U35117 (N_35117,N_34551,N_30589);
nand U35118 (N_35118,N_33413,N_33075);
nand U35119 (N_35119,N_34820,N_32868);
nand U35120 (N_35120,N_30468,N_30911);
or U35121 (N_35121,N_34709,N_32587);
nand U35122 (N_35122,N_30313,N_33318);
nand U35123 (N_35123,N_30986,N_30189);
nor U35124 (N_35124,N_32884,N_34902);
or U35125 (N_35125,N_30936,N_31448);
nand U35126 (N_35126,N_30068,N_31792);
nand U35127 (N_35127,N_34642,N_33851);
and U35128 (N_35128,N_30784,N_34676);
and U35129 (N_35129,N_31469,N_32878);
xnor U35130 (N_35130,N_30650,N_33808);
xnor U35131 (N_35131,N_32702,N_32918);
nand U35132 (N_35132,N_30977,N_33528);
xnor U35133 (N_35133,N_33000,N_32331);
xnor U35134 (N_35134,N_31621,N_31028);
nand U35135 (N_35135,N_33971,N_34298);
or U35136 (N_35136,N_33129,N_34252);
xnor U35137 (N_35137,N_30631,N_32369);
xnor U35138 (N_35138,N_31050,N_34209);
nand U35139 (N_35139,N_32639,N_31764);
xor U35140 (N_35140,N_32080,N_30378);
nand U35141 (N_35141,N_32797,N_34950);
and U35142 (N_35142,N_32984,N_31123);
xnor U35143 (N_35143,N_30187,N_30634);
and U35144 (N_35144,N_33301,N_31687);
nand U35145 (N_35145,N_33770,N_33444);
or U35146 (N_35146,N_32839,N_32805);
and U35147 (N_35147,N_32472,N_30029);
and U35148 (N_35148,N_30221,N_32585);
or U35149 (N_35149,N_30696,N_33753);
nand U35150 (N_35150,N_34162,N_34184);
or U35151 (N_35151,N_33677,N_31297);
xor U35152 (N_35152,N_30214,N_33475);
or U35153 (N_35153,N_33306,N_34767);
or U35154 (N_35154,N_31336,N_32708);
or U35155 (N_35155,N_33104,N_31564);
or U35156 (N_35156,N_30734,N_34893);
and U35157 (N_35157,N_34837,N_32127);
xor U35158 (N_35158,N_30758,N_33972);
xnor U35159 (N_35159,N_31405,N_33264);
or U35160 (N_35160,N_33407,N_31868);
nand U35161 (N_35161,N_31407,N_32023);
or U35162 (N_35162,N_32864,N_33784);
xnor U35163 (N_35163,N_30445,N_32771);
or U35164 (N_35164,N_31644,N_30379);
xor U35165 (N_35165,N_33488,N_32922);
nand U35166 (N_35166,N_32819,N_34940);
xor U35167 (N_35167,N_33047,N_31332);
nand U35168 (N_35168,N_34864,N_32482);
xor U35169 (N_35169,N_31816,N_33393);
nor U35170 (N_35170,N_31998,N_33558);
or U35171 (N_35171,N_34267,N_30080);
or U35172 (N_35172,N_34783,N_34100);
xor U35173 (N_35173,N_30022,N_34196);
and U35174 (N_35174,N_33192,N_30761);
nand U35175 (N_35175,N_33304,N_33583);
nand U35176 (N_35176,N_31766,N_32596);
or U35177 (N_35177,N_30963,N_34001);
nand U35178 (N_35178,N_31793,N_31550);
nor U35179 (N_35179,N_32737,N_34511);
nor U35180 (N_35180,N_30203,N_31786);
or U35181 (N_35181,N_31143,N_32373);
and U35182 (N_35182,N_31928,N_32002);
nor U35183 (N_35183,N_34970,N_32870);
and U35184 (N_35184,N_31634,N_30897);
nand U35185 (N_35185,N_32856,N_30747);
and U35186 (N_35186,N_30019,N_34021);
nand U35187 (N_35187,N_33658,N_33063);
xnor U35188 (N_35188,N_30783,N_30895);
or U35189 (N_35189,N_30507,N_33533);
nand U35190 (N_35190,N_31920,N_32595);
nor U35191 (N_35191,N_34916,N_33542);
or U35192 (N_35192,N_34336,N_32493);
xnor U35193 (N_35193,N_33279,N_34534);
nor U35194 (N_35194,N_33885,N_34317);
and U35195 (N_35195,N_30884,N_32890);
xnor U35196 (N_35196,N_33421,N_34455);
and U35197 (N_35197,N_30852,N_33675);
or U35198 (N_35198,N_34628,N_32866);
and U35199 (N_35199,N_32532,N_30930);
or U35200 (N_35200,N_31076,N_32116);
and U35201 (N_35201,N_30652,N_33406);
xnor U35202 (N_35202,N_32417,N_31670);
nor U35203 (N_35203,N_30989,N_33130);
nor U35204 (N_35204,N_32340,N_33616);
nor U35205 (N_35205,N_33397,N_30833);
or U35206 (N_35206,N_32098,N_34959);
and U35207 (N_35207,N_32599,N_30241);
nor U35208 (N_35208,N_33813,N_30474);
and U35209 (N_35209,N_33938,N_31822);
and U35210 (N_35210,N_30398,N_33254);
and U35211 (N_35211,N_34265,N_34850);
and U35212 (N_35212,N_31226,N_33995);
or U35213 (N_35213,N_30858,N_30300);
and U35214 (N_35214,N_33605,N_30359);
nor U35215 (N_35215,N_34897,N_34542);
xnor U35216 (N_35216,N_33175,N_33067);
nand U35217 (N_35217,N_30051,N_34403);
or U35218 (N_35218,N_32951,N_33769);
or U35219 (N_35219,N_31936,N_32060);
nor U35220 (N_35220,N_31775,N_30692);
and U35221 (N_35221,N_30843,N_32118);
nand U35222 (N_35222,N_31196,N_34907);
xnor U35223 (N_35223,N_30967,N_34286);
and U35224 (N_35224,N_30559,N_34169);
nor U35225 (N_35225,N_32486,N_31445);
nor U35226 (N_35226,N_32876,N_34310);
nor U35227 (N_35227,N_30308,N_34125);
nor U35228 (N_35228,N_34102,N_30918);
nor U35229 (N_35229,N_30234,N_30575);
and U35230 (N_35230,N_31057,N_34091);
nor U35231 (N_35231,N_34634,N_30772);
xor U35232 (N_35232,N_33066,N_32808);
nand U35233 (N_35233,N_33746,N_33050);
nand U35234 (N_35234,N_32888,N_34247);
nand U35235 (N_35235,N_34821,N_30129);
nor U35236 (N_35236,N_32490,N_30140);
xor U35237 (N_35237,N_34120,N_32416);
xor U35238 (N_35238,N_31947,N_31579);
nor U35239 (N_35239,N_32966,N_31215);
nand U35240 (N_35240,N_31075,N_34407);
nor U35241 (N_35241,N_33841,N_34846);
or U35242 (N_35242,N_32637,N_34771);
nor U35243 (N_35243,N_34612,N_34811);
nand U35244 (N_35244,N_33131,N_34373);
xor U35245 (N_35245,N_33053,N_34389);
nand U35246 (N_35246,N_33056,N_31554);
nand U35247 (N_35247,N_34325,N_30705);
and U35248 (N_35248,N_32628,N_33564);
and U35249 (N_35249,N_32111,N_33269);
and U35250 (N_35250,N_32728,N_33910);
nand U35251 (N_35251,N_31872,N_33044);
nor U35252 (N_35252,N_32500,N_31744);
nor U35253 (N_35253,N_33895,N_30681);
xor U35254 (N_35254,N_34240,N_31770);
nor U35255 (N_35255,N_33042,N_31522);
or U35256 (N_35256,N_32137,N_31778);
and U35257 (N_35257,N_31271,N_31939);
and U35258 (N_35258,N_30371,N_30220);
nand U35259 (N_35259,N_34580,N_30084);
xnor U35260 (N_35260,N_30531,N_33300);
nand U35261 (N_35261,N_34223,N_33256);
nand U35262 (N_35262,N_33190,N_33966);
xnor U35263 (N_35263,N_33354,N_32941);
or U35264 (N_35264,N_32858,N_34136);
and U35265 (N_35265,N_32843,N_32082);
and U35266 (N_35266,N_31037,N_31968);
nand U35267 (N_35267,N_33427,N_33509);
xnor U35268 (N_35268,N_31819,N_31736);
or U35269 (N_35269,N_32505,N_34974);
nor U35270 (N_35270,N_31552,N_31815);
nand U35271 (N_35271,N_32697,N_32935);
and U35272 (N_35272,N_31688,N_30708);
or U35273 (N_35273,N_34935,N_34068);
and U35274 (N_35274,N_32853,N_33987);
or U35275 (N_35275,N_34978,N_31329);
xnor U35276 (N_35276,N_30410,N_33835);
or U35277 (N_35277,N_30823,N_31388);
nand U35278 (N_35278,N_32234,N_32304);
xor U35279 (N_35279,N_32977,N_33574);
nor U35280 (N_35280,N_32147,N_32131);
nor U35281 (N_35281,N_32208,N_34024);
nand U35282 (N_35282,N_33526,N_31570);
and U35283 (N_35283,N_34242,N_33442);
xnor U35284 (N_35284,N_34280,N_31877);
xor U35285 (N_35285,N_30419,N_32293);
xnor U35286 (N_35286,N_32372,N_33153);
and U35287 (N_35287,N_32363,N_34721);
and U35288 (N_35288,N_33227,N_32593);
nor U35289 (N_35289,N_34383,N_34422);
nor U35290 (N_35290,N_34076,N_32698);
or U35291 (N_35291,N_33676,N_34505);
nor U35292 (N_35292,N_30978,N_33473);
nor U35293 (N_35293,N_34409,N_33919);
nor U35294 (N_35294,N_33357,N_34013);
nor U35295 (N_35295,N_30506,N_34074);
nand U35296 (N_35296,N_34191,N_34591);
and U35297 (N_35297,N_30018,N_31987);
nand U35298 (N_35298,N_34677,N_33668);
xor U35299 (N_35299,N_32004,N_32035);
nand U35300 (N_35300,N_33646,N_31389);
nor U35301 (N_35301,N_33683,N_31598);
or U35302 (N_35302,N_32914,N_32638);
nand U35303 (N_35303,N_34367,N_30274);
and U35304 (N_35304,N_34127,N_34456);
xor U35305 (N_35305,N_33960,N_31043);
or U35306 (N_35306,N_34270,N_34322);
and U35307 (N_35307,N_30725,N_30600);
or U35308 (N_35308,N_33140,N_30985);
or U35309 (N_35309,N_31021,N_31119);
nand U35310 (N_35310,N_30257,N_32995);
nand U35311 (N_35311,N_33145,N_31826);
and U35312 (N_35312,N_31098,N_32921);
nor U35313 (N_35313,N_30372,N_33467);
nor U35314 (N_35314,N_31875,N_32114);
nor U35315 (N_35315,N_30367,N_33637);
and U35316 (N_35316,N_30045,N_34857);
or U35317 (N_35317,N_30908,N_31066);
and U35318 (N_35318,N_34464,N_33556);
xnor U35319 (N_35319,N_34675,N_34947);
and U35320 (N_35320,N_31342,N_32383);
nand U35321 (N_35321,N_33505,N_33871);
nor U35322 (N_35322,N_34453,N_30388);
xnor U35323 (N_35323,N_33554,N_31398);
nor U35324 (N_35324,N_33693,N_34773);
and U35325 (N_35325,N_32660,N_31091);
and U35326 (N_35326,N_34029,N_33284);
and U35327 (N_35327,N_33088,N_30500);
nand U35328 (N_35328,N_30605,N_34860);
nand U35329 (N_35329,N_31650,N_32243);
nor U35330 (N_35330,N_33241,N_30697);
nand U35331 (N_35331,N_34954,N_34083);
and U35332 (N_35332,N_34160,N_34666);
xor U35333 (N_35333,N_33598,N_30988);
nand U35334 (N_35334,N_31070,N_33117);
and U35335 (N_35335,N_34865,N_31907);
or U35336 (N_35336,N_31452,N_30594);
nor U35337 (N_35337,N_33619,N_32865);
xor U35338 (N_35338,N_31333,N_30484);
nor U35339 (N_35339,N_33211,N_34898);
xor U35340 (N_35340,N_32540,N_30752);
and U35341 (N_35341,N_31781,N_33365);
and U35342 (N_35342,N_32397,N_33029);
nor U35343 (N_35343,N_31195,N_32546);
nor U35344 (N_35344,N_30317,N_34206);
or U35345 (N_35345,N_31664,N_32844);
or U35346 (N_35346,N_31121,N_30389);
or U35347 (N_35347,N_32527,N_30164);
and U35348 (N_35348,N_34299,N_32045);
xor U35349 (N_35349,N_32820,N_30866);
nor U35350 (N_35350,N_33661,N_34578);
nor U35351 (N_35351,N_32762,N_32092);
nand U35352 (N_35352,N_33584,N_32852);
and U35353 (N_35353,N_33447,N_32146);
or U35354 (N_35354,N_32756,N_33980);
nor U35355 (N_35355,N_32479,N_30567);
xnor U35356 (N_35356,N_31399,N_31878);
or U35357 (N_35357,N_33333,N_31157);
nor U35358 (N_35358,N_31126,N_34126);
or U35359 (N_35359,N_32478,N_31985);
and U35360 (N_35360,N_32550,N_34904);
or U35361 (N_35361,N_34463,N_32643);
nor U35362 (N_35362,N_33378,N_34538);
nor U35363 (N_35363,N_33875,N_34763);
xor U35364 (N_35364,N_30413,N_31503);
or U35365 (N_35365,N_30547,N_31305);
nand U35366 (N_35366,N_34334,N_32219);
or U35367 (N_35367,N_32303,N_32249);
or U35368 (N_35368,N_31400,N_30521);
or U35369 (N_35369,N_32074,N_32049);
or U35370 (N_35370,N_31791,N_33932);
or U35371 (N_35371,N_33849,N_34069);
or U35372 (N_35372,N_31994,N_34390);
and U35373 (N_35373,N_32537,N_32162);
nand U35374 (N_35374,N_32380,N_31575);
or U35375 (N_35375,N_33648,N_31217);
nor U35376 (N_35376,N_31576,N_34084);
nand U35377 (N_35377,N_33578,N_30057);
and U35378 (N_35378,N_32071,N_32949);
and U35379 (N_35379,N_33906,N_32563);
and U35380 (N_35380,N_31230,N_30108);
nand U35381 (N_35381,N_33186,N_32523);
and U35382 (N_35382,N_33043,N_32188);
or U35383 (N_35383,N_33511,N_32511);
and U35384 (N_35384,N_33120,N_32189);
and U35385 (N_35385,N_31647,N_30167);
nor U35386 (N_35386,N_33633,N_30023);
nand U35387 (N_35387,N_32804,N_33368);
nand U35388 (N_35388,N_34725,N_32083);
or U35389 (N_35389,N_34790,N_32768);
xor U35390 (N_35390,N_31296,N_32586);
xnor U35391 (N_35391,N_32692,N_30012);
xnor U35392 (N_35392,N_30805,N_32662);
xor U35393 (N_35393,N_32081,N_34807);
nand U35394 (N_35394,N_32015,N_34337);
nor U35395 (N_35395,N_30297,N_33752);
xnor U35396 (N_35396,N_30149,N_31009);
xnor U35397 (N_35397,N_32483,N_31595);
xor U35398 (N_35398,N_32745,N_32426);
and U35399 (N_35399,N_34514,N_34393);
and U35400 (N_35400,N_34043,N_30006);
nand U35401 (N_35401,N_34040,N_34687);
and U35402 (N_35402,N_32153,N_34858);
or U35403 (N_35403,N_31172,N_33707);
nand U35404 (N_35404,N_30958,N_30139);
nand U35405 (N_35405,N_30904,N_33341);
and U35406 (N_35406,N_31191,N_32086);
or U35407 (N_35407,N_31345,N_34082);
nand U35408 (N_35408,N_32861,N_32468);
or U35409 (N_35409,N_31535,N_32048);
nand U35410 (N_35410,N_31622,N_31487);
or U35411 (N_35411,N_31633,N_33202);
nor U35412 (N_35412,N_34797,N_31995);
nand U35413 (N_35413,N_34720,N_34863);
or U35414 (N_35414,N_34607,N_30669);
xnor U35415 (N_35415,N_30615,N_34785);
and U35416 (N_35416,N_30428,N_31326);
nand U35417 (N_35417,N_34637,N_34199);
and U35418 (N_35418,N_33941,N_33937);
nand U35419 (N_35419,N_30193,N_33002);
xnor U35420 (N_35420,N_34382,N_30764);
nor U35421 (N_35421,N_30686,N_31260);
or U35422 (N_35422,N_34717,N_32032);
nor U35423 (N_35423,N_33719,N_32375);
or U35424 (N_35424,N_30972,N_31135);
or U35425 (N_35425,N_34468,N_34662);
nand U35426 (N_35426,N_34856,N_33812);
or U35427 (N_35427,N_30251,N_32183);
and U35428 (N_35428,N_31817,N_31324);
xor U35429 (N_35429,N_31561,N_32175);
or U35430 (N_35430,N_32555,N_33474);
and U35431 (N_35431,N_34640,N_34792);
nor U35432 (N_35432,N_34167,N_30968);
nand U35433 (N_35433,N_32909,N_30592);
xor U35434 (N_35434,N_31565,N_33340);
nor U35435 (N_35435,N_32459,N_33983);
and U35436 (N_35436,N_30208,N_30041);
xnor U35437 (N_35437,N_34566,N_30607);
nand U35438 (N_35438,N_34316,N_30574);
or U35439 (N_35439,N_34878,N_33958);
xor U35440 (N_35440,N_30868,N_30331);
and U35441 (N_35441,N_32946,N_32645);
and U35442 (N_35442,N_30401,N_31289);
or U35443 (N_35443,N_30142,N_33775);
or U35444 (N_35444,N_33419,N_30110);
or U35445 (N_35445,N_34285,N_31272);
nor U35446 (N_35446,N_34758,N_33944);
and U35447 (N_35447,N_32979,N_32758);
or U35448 (N_35448,N_33920,N_31318);
or U35449 (N_35449,N_32667,N_34307);
or U35450 (N_35450,N_33565,N_34546);
nor U35451 (N_35451,N_30235,N_34595);
or U35452 (N_35452,N_32322,N_31108);
xor U35453 (N_35453,N_32993,N_31864);
nor U35454 (N_35454,N_30707,N_33688);
nand U35455 (N_35455,N_31236,N_31455);
nor U35456 (N_35456,N_30674,N_30485);
nor U35457 (N_35457,N_31358,N_30800);
or U35458 (N_35458,N_33123,N_31807);
nand U35459 (N_35459,N_33096,N_32933);
nor U35460 (N_35460,N_33614,N_34736);
nand U35461 (N_35461,N_31927,N_33161);
nor U35462 (N_35462,N_34192,N_33725);
and U35463 (N_35463,N_32695,N_31222);
xor U35464 (N_35464,N_30770,N_31387);
nand U35465 (N_35465,N_34404,N_30834);
or U35466 (N_35466,N_33710,N_30813);
or U35467 (N_35467,N_33200,N_32950);
nor U35468 (N_35468,N_30802,N_34243);
and U35469 (N_35469,N_30104,N_33325);
and U35470 (N_35470,N_30743,N_34809);
nand U35471 (N_35471,N_30845,N_31520);
and U35472 (N_35472,N_34028,N_32433);
xnor U35473 (N_35473,N_32297,N_32529);
or U35474 (N_35474,N_30121,N_31115);
and U35475 (N_35475,N_33207,N_30148);
or U35476 (N_35476,N_33673,N_31295);
or U35477 (N_35477,N_33811,N_30582);
nand U35478 (N_35478,N_32829,N_33534);
and U35479 (N_35479,N_30541,N_30577);
nor U35480 (N_35480,N_32666,N_32379);
nand U35481 (N_35481,N_34688,N_34277);
xor U35482 (N_35482,N_34030,N_32954);
nor U35483 (N_35483,N_32827,N_33655);
nor U35484 (N_35484,N_31711,N_33454);
nor U35485 (N_35485,N_31228,N_34841);
nor U35486 (N_35486,N_30539,N_34465);
nor U35487 (N_35487,N_34054,N_33965);
and U35488 (N_35488,N_30927,N_33720);
or U35489 (N_35489,N_31966,N_31538);
nand U35490 (N_35490,N_33728,N_31431);
and U35491 (N_35491,N_30103,N_32233);
and U35492 (N_35492,N_33581,N_32159);
nand U35493 (N_35493,N_31499,N_30797);
xnor U35494 (N_35494,N_32655,N_31892);
nand U35495 (N_35495,N_32157,N_34472);
xor U35496 (N_35496,N_32597,N_31283);
and U35497 (N_35497,N_30703,N_30614);
nor U35498 (N_35498,N_34594,N_34062);
xor U35499 (N_35499,N_34845,N_31209);
nand U35500 (N_35500,N_31964,N_32392);
or U35501 (N_35501,N_32714,N_31862);
xor U35502 (N_35502,N_33636,N_33727);
xnor U35503 (N_35503,N_34170,N_31837);
nand U35504 (N_35504,N_30374,N_32200);
nor U35505 (N_35505,N_30411,N_31706);
nand U35506 (N_35506,N_34992,N_31643);
or U35507 (N_35507,N_33025,N_30284);
or U35508 (N_35508,N_32044,N_34229);
or U35509 (N_35509,N_31850,N_30848);
or U35510 (N_35510,N_33417,N_31630);
or U35511 (N_35511,N_34971,N_30693);
nor U35512 (N_35512,N_33751,N_30780);
nor U35513 (N_35513,N_31410,N_30599);
xor U35514 (N_35514,N_30403,N_30298);
or U35515 (N_35515,N_33376,N_33585);
and U35516 (N_35516,N_31835,N_31838);
xnor U35517 (N_35517,N_32431,N_30869);
nand U35518 (N_35518,N_30662,N_34670);
nand U35519 (N_35519,N_33577,N_34151);
nor U35520 (N_35520,N_32608,N_31910);
or U35521 (N_35521,N_34009,N_31975);
nor U35522 (N_35522,N_33360,N_30294);
nand U35523 (N_35523,N_33107,N_33424);
xor U35524 (N_35524,N_31225,N_34685);
nor U35525 (N_35525,N_33317,N_31424);
nor U35526 (N_35526,N_31241,N_31937);
xor U35527 (N_35527,N_32067,N_34800);
nor U35528 (N_35528,N_30250,N_30533);
xnor U35529 (N_35529,N_30116,N_34225);
nand U35530 (N_35530,N_31703,N_30606);
nor U35531 (N_35531,N_34756,N_33007);
nor U35532 (N_35532,N_33187,N_30376);
nand U35533 (N_35533,N_31282,N_31396);
and U35534 (N_35534,N_34755,N_34189);
xnor U35535 (N_35535,N_31978,N_30983);
xor U35536 (N_35536,N_34402,N_33800);
xnor U35537 (N_35537,N_33377,N_31379);
or U35538 (N_35538,N_30173,N_32711);
or U35539 (N_35539,N_34817,N_33687);
and U35540 (N_35540,N_34469,N_31382);
xor U35541 (N_35541,N_34590,N_30821);
nor U35542 (N_35542,N_30382,N_30286);
or U35543 (N_35543,N_31523,N_30957);
or U35544 (N_35544,N_30552,N_32669);
and U35545 (N_35545,N_34283,N_34777);
nand U35546 (N_35546,N_33478,N_30079);
xnor U35547 (N_35547,N_33519,N_33041);
nor U35548 (N_35548,N_33629,N_31188);
nor U35549 (N_35549,N_31265,N_31671);
and U35550 (N_35550,N_32430,N_30854);
nand U35551 (N_35551,N_31942,N_33686);
or U35552 (N_35552,N_32694,N_32115);
nand U35553 (N_35553,N_31039,N_30450);
and U35554 (N_35554,N_34516,N_32798);
xnor U35555 (N_35555,N_30131,N_33663);
xnor U35556 (N_35556,N_31980,N_34567);
or U35557 (N_35557,N_30724,N_32894);
nor U35558 (N_35558,N_34504,N_33231);
nor U35559 (N_35559,N_32627,N_31934);
nand U35560 (N_35560,N_30637,N_33984);
nand U35561 (N_35561,N_32510,N_33848);
xnor U35562 (N_35562,N_32603,N_33537);
or U35563 (N_35563,N_31234,N_30665);
or U35564 (N_35564,N_32671,N_30861);
nand U35565 (N_35565,N_34047,N_34875);
nand U35566 (N_35566,N_32874,N_30653);
nand U35567 (N_35567,N_31654,N_31339);
or U35568 (N_35568,N_32752,N_30252);
and U35569 (N_35569,N_30952,N_33690);
and U35570 (N_35570,N_34494,N_33109);
nand U35571 (N_35571,N_32163,N_34997);
nand U35572 (N_35572,N_30192,N_34416);
nor U35573 (N_35573,N_30771,N_34235);
nand U35574 (N_35574,N_31814,N_32204);
xnor U35575 (N_35575,N_32412,N_33220);
xnor U35576 (N_35576,N_31951,N_30332);
and U35577 (N_35577,N_32783,N_31642);
and U35578 (N_35578,N_30889,N_33490);
and U35579 (N_35579,N_32975,N_30923);
and U35580 (N_35580,N_33809,N_31516);
xor U35581 (N_35581,N_33644,N_33680);
nand U35582 (N_35582,N_33573,N_30452);
nor U35583 (N_35583,N_32496,N_34385);
and U35584 (N_35584,N_32543,N_33224);
nand U35585 (N_35585,N_34097,N_34448);
nand U35586 (N_35586,N_30836,N_30171);
xor U35587 (N_35587,N_33961,N_31276);
or U35588 (N_35588,N_30864,N_31635);
xor U35589 (N_35589,N_30901,N_33955);
and U35590 (N_35590,N_31845,N_31502);
and U35591 (N_35591,N_33763,N_34877);
xor U35592 (N_35592,N_30719,N_31253);
or U35593 (N_35593,N_34193,N_31356);
nor U35594 (N_35594,N_33842,N_30237);
xnor U35595 (N_35595,N_30329,N_34147);
xnor U35596 (N_35596,N_30863,N_30272);
nand U35597 (N_35597,N_32886,N_33726);
or U35598 (N_35598,N_33027,N_33136);
nor U35599 (N_35599,N_34798,N_34266);
nand U35600 (N_35600,N_30209,N_33917);
and U35601 (N_35601,N_34035,N_32678);
and U35602 (N_35602,N_33322,N_32998);
xnor U35603 (N_35603,N_33210,N_34141);
and U35604 (N_35604,N_31704,N_33786);
or U35605 (N_35605,N_33432,N_33355);
nand U35606 (N_35606,N_33538,N_30228);
nor U35607 (N_35607,N_30088,N_31320);
xor U35608 (N_35608,N_33523,N_34574);
or U35609 (N_35609,N_33267,N_34853);
xor U35610 (N_35610,N_34431,N_34087);
nand U35611 (N_35611,N_33426,N_32268);
or U35612 (N_35612,N_32325,N_32041);
or U35613 (N_35613,N_33595,N_34217);
nand U35614 (N_35614,N_32197,N_30449);
or U35615 (N_35615,N_34394,N_31314);
xor U35616 (N_35616,N_32251,N_32716);
nand U35617 (N_35617,N_34000,N_32437);
xor U35618 (N_35618,N_30946,N_33896);
and U35619 (N_35619,N_31383,N_32814);
and U35620 (N_35620,N_30342,N_30540);
nor U35621 (N_35621,N_34543,N_30078);
nor U35622 (N_35622,N_32924,N_32504);
or U35623 (N_35623,N_34526,N_34624);
or U35624 (N_35624,N_33524,N_33810);
xnor U35625 (N_35625,N_32624,N_33429);
nor U35626 (N_35626,N_30334,N_32145);
or U35627 (N_35627,N_30860,N_32274);
and U35628 (N_35628,N_32670,N_31069);
nand U35629 (N_35629,N_31397,N_32494);
and U35630 (N_35630,N_32366,N_30828);
xor U35631 (N_35631,N_31184,N_34014);
xnor U35632 (N_35632,N_30357,N_33182);
nand U35633 (N_35633,N_34200,N_34848);
xor U35634 (N_35634,N_33986,N_31112);
or U35635 (N_35635,N_30296,N_30440);
xnor U35636 (N_35636,N_34498,N_33013);
and U35637 (N_35637,N_33870,N_31187);
or U35638 (N_35638,N_31899,N_32438);
xnor U35639 (N_35639,N_34356,N_31923);
nor U35640 (N_35640,N_34881,N_34706);
and U35641 (N_35641,N_34220,N_30584);
xor U35642 (N_35642,N_33297,N_34579);
and U35643 (N_35643,N_30368,N_31125);
nor U35644 (N_35644,N_34535,N_30262);
or U35645 (N_35645,N_30825,N_33081);
nand U35646 (N_35646,N_30000,N_31805);
xor U35647 (N_35647,N_30361,N_32093);
and U35648 (N_35648,N_34822,N_34921);
nor U35649 (N_35649,N_34824,N_34842);
or U35650 (N_35650,N_31788,N_34521);
and U35651 (N_35651,N_32199,N_33087);
xnor U35652 (N_35652,N_34710,N_32945);
xor U35653 (N_35653,N_33883,N_32343);
nand U35654 (N_35654,N_30344,N_34341);
xor U35655 (N_35655,N_33179,N_33569);
or U35656 (N_35656,N_31763,N_32042);
xnor U35657 (N_35657,N_31461,N_34378);
xor U35658 (N_35658,N_33353,N_30621);
nand U35659 (N_35659,N_32245,N_34900);
nor U35660 (N_35660,N_33838,N_31466);
or U35661 (N_35661,N_34680,N_31693);
and U35662 (N_35662,N_32037,N_34654);
nand U35663 (N_35663,N_34555,N_34195);
nor U35664 (N_35664,N_34615,N_30995);
and U35665 (N_35665,N_33723,N_30354);
nor U35666 (N_35666,N_33326,N_32315);
and U35667 (N_35667,N_31033,N_34861);
and U35668 (N_35668,N_34573,N_32134);
and U35669 (N_35669,N_32718,N_32775);
or U35670 (N_35670,N_32980,N_30702);
or U35671 (N_35671,N_30846,N_34939);
nand U35672 (N_35672,N_33486,N_31577);
and U35673 (N_35673,N_33095,N_30808);
and U35674 (N_35674,N_34046,N_34304);
nor U35675 (N_35675,N_34006,N_31082);
or U35676 (N_35676,N_31821,N_31361);
nand U35677 (N_35677,N_32934,N_30604);
xor U35678 (N_35678,N_31210,N_30225);
nand U35679 (N_35679,N_32963,N_31560);
or U35680 (N_35680,N_34381,N_30691);
and U35681 (N_35681,N_33006,N_30723);
or U35682 (N_35682,N_30133,N_31855);
or U35683 (N_35683,N_31116,N_31099);
or U35684 (N_35684,N_32990,N_34805);
nor U35685 (N_35685,N_33162,N_34599);
nor U35686 (N_35686,N_31041,N_32749);
nor U35687 (N_35687,N_33222,N_33706);
or U35688 (N_35688,N_31325,N_30714);
nor U35689 (N_35689,N_30147,N_32012);
nor U35690 (N_35690,N_31739,N_31137);
nor U35691 (N_35691,N_32748,N_32276);
and U35692 (N_35692,N_34483,N_32321);
xnor U35693 (N_35693,N_33589,N_31486);
and U35694 (N_35694,N_33023,N_33431);
nand U35695 (N_35695,N_30658,N_30461);
or U35696 (N_35696,N_32088,N_34960);
nand U35697 (N_35697,N_30678,N_31915);
nand U35698 (N_35698,N_34981,N_32030);
and U35699 (N_35699,N_30488,N_34428);
xor U35700 (N_35700,N_32766,N_30335);
or U35701 (N_35701,N_32786,N_30305);
or U35702 (N_35702,N_31309,N_30162);
xnor U35703 (N_35703,N_31566,N_34156);
nor U35704 (N_35704,N_34617,N_30522);
or U35705 (N_35705,N_31973,N_31909);
or U35706 (N_35706,N_32072,N_33643);
nand U35707 (N_35707,N_31390,N_34411);
and U35708 (N_35708,N_33956,N_34236);
and U35709 (N_35709,N_33918,N_30934);
nand U35710 (N_35710,N_34986,N_33449);
nand U35711 (N_35711,N_30789,N_33548);
xor U35712 (N_35712,N_30360,N_30132);
nor U35713 (N_35713,N_34669,N_33201);
xnor U35714 (N_35714,N_30666,N_31246);
xor U35715 (N_35715,N_34460,N_32986);
or U35716 (N_35716,N_34572,N_30654);
nand U35717 (N_35717,N_33865,N_33452);
xor U35718 (N_35718,N_33184,N_33593);
and U35719 (N_35719,N_31347,N_33750);
nand U35720 (N_35720,N_34441,N_30090);
nand U35721 (N_35721,N_30679,N_30091);
or U35722 (N_35722,N_30060,N_34384);
xnor U35723 (N_35723,N_32432,N_33398);
or U35724 (N_35724,N_30550,N_31829);
nor U35725 (N_35725,N_34154,N_32367);
nand U35726 (N_35726,N_32022,N_32305);
or U35727 (N_35727,N_34258,N_30831);
or U35728 (N_35728,N_30512,N_34544);
nor U35729 (N_35729,N_33715,N_30215);
nor U35730 (N_35730,N_33859,N_30065);
xor U35731 (N_35731,N_31780,N_31232);
nor U35732 (N_35732,N_30328,N_32402);
nand U35733 (N_35733,N_32381,N_31783);
nand U35734 (N_35734,N_30906,N_31578);
nor U35735 (N_35735,N_32143,N_33351);
or U35736 (N_35736,N_30324,N_31772);
nand U35737 (N_35737,N_31355,N_31849);
nand U35738 (N_35738,N_32807,N_33926);
xnor U35739 (N_35739,N_32760,N_32326);
and U35740 (N_35740,N_32029,N_30682);
nor U35741 (N_35741,N_32195,N_32810);
and U35742 (N_35742,N_34984,N_32275);
and U35743 (N_35743,N_31353,N_30815);
nor U35744 (N_35744,N_30201,N_34295);
xnor U35745 (N_35745,N_33520,N_30292);
and U35746 (N_35746,N_34682,N_30082);
xor U35747 (N_35747,N_31364,N_32232);
or U35748 (N_35748,N_34517,N_31483);
or U35749 (N_35749,N_31498,N_33098);
nand U35750 (N_35750,N_33366,N_33494);
and U35751 (N_35751,N_31658,N_31334);
nor U35752 (N_35752,N_34532,N_32250);
or U35753 (N_35753,N_31036,N_34073);
nand U35754 (N_35754,N_30717,N_32617);
xor U35755 (N_35755,N_32584,N_33146);
nor U35756 (N_35756,N_34764,N_31771);
and U35757 (N_35757,N_34585,N_30166);
nand U35758 (N_35758,N_32733,N_33887);
or U35759 (N_35759,N_32908,N_30226);
nand U35760 (N_35760,N_31761,N_30024);
nand U35761 (N_35761,N_34296,N_34941);
nand U35762 (N_35762,N_30503,N_31441);
nand U35763 (N_35763,N_33959,N_30699);
nor U35764 (N_35764,N_32209,N_32571);
or U35765 (N_35765,N_34847,N_30076);
or U35766 (N_35766,N_30426,N_31426);
nand U35767 (N_35767,N_34360,N_31323);
nand U35768 (N_35768,N_32436,N_30501);
nand U35769 (N_35769,N_31465,N_31690);
nor U35770 (N_35770,N_33501,N_34086);
or U35771 (N_35771,N_33561,N_30453);
and U35772 (N_35772,N_34605,N_31668);
nor U35773 (N_35773,N_31081,N_31559);
and U35774 (N_35774,N_31078,N_34645);
xnor U35775 (N_35775,N_34423,N_33532);
and U35776 (N_35776,N_31542,N_30431);
xnor U35777 (N_35777,N_30516,N_34412);
and U35778 (N_35778,N_31146,N_34466);
or U35779 (N_35779,N_32317,N_31972);
or U35780 (N_35780,N_30211,N_31917);
and U35781 (N_35781,N_34353,N_33788);
xor U35782 (N_35782,N_32823,N_33627);
and U35783 (N_35783,N_32741,N_31480);
xnor U35784 (N_35784,N_33126,N_34410);
or U35785 (N_35785,N_33764,N_33826);
and U35786 (N_35786,N_34004,N_34161);
nand U35787 (N_35787,N_34525,N_30776);
or U35788 (N_35788,N_31149,N_33418);
nor U35789 (N_35789,N_33836,N_32360);
or U35790 (N_35790,N_30892,N_31641);
nor U35791 (N_35791,N_34547,N_32231);
and U35792 (N_35792,N_30620,N_34226);
or U35793 (N_35793,N_33443,N_31753);
and U35794 (N_35794,N_33394,N_33767);
nor U35795 (N_35795,N_33350,N_33625);
nand U35796 (N_35796,N_32725,N_34140);
xnor U35797 (N_35797,N_31485,N_30218);
nand U35798 (N_35798,N_34646,N_34368);
nor U35799 (N_35799,N_34182,N_34548);
nor U35800 (N_35800,N_31870,N_34883);
nand U35801 (N_35801,N_31030,N_31506);
nand U35802 (N_35802,N_31737,N_33789);
nand U35803 (N_35803,N_33890,N_30480);
xor U35804 (N_35804,N_32535,N_33453);
and U35805 (N_35805,N_32215,N_33059);
nand U35806 (N_35806,N_32912,N_30824);
xnor U35807 (N_35807,N_34584,N_30632);
nand U35808 (N_35808,N_33209,N_33653);
xnor U35809 (N_35809,N_33923,N_31287);
nor U35810 (N_35810,N_32845,N_30586);
and U35811 (N_35811,N_32105,N_34772);
or U35812 (N_35812,N_32607,N_31724);
nor U35813 (N_35813,N_34678,N_31330);
or U35814 (N_35814,N_33722,N_30753);
nor U35815 (N_35815,N_34128,N_31103);
or U35816 (N_35816,N_33557,N_32606);
xnor U35817 (N_35817,N_30617,N_30343);
nor U35818 (N_35818,N_33617,N_31893);
xnor U35819 (N_35819,N_30579,N_31645);
or U35820 (N_35820,N_30612,N_33156);
and U35821 (N_35821,N_32778,N_33793);
nor U35822 (N_35822,N_31017,N_32119);
or U35823 (N_35823,N_33434,N_34388);
and U35824 (N_35824,N_32485,N_31060);
xor U35825 (N_35825,N_32411,N_32887);
xor U35826 (N_35826,N_34512,N_32149);
nor U35827 (N_35827,N_30085,N_31087);
or U35828 (N_35828,N_31989,N_32242);
nor U35829 (N_35829,N_31254,N_30094);
xnor U35830 (N_35830,N_34601,N_32629);
nand U35831 (N_35831,N_33015,N_30535);
nand U35832 (N_35832,N_30515,N_30141);
and U35833 (N_35833,N_31843,N_33460);
or U35834 (N_35834,N_31800,N_34818);
or U35835 (N_35835,N_32885,N_32388);
nand U35836 (N_35836,N_32129,N_33635);
or U35837 (N_35837,N_34522,N_30973);
and U35838 (N_35838,N_32507,N_33597);
or U35839 (N_35839,N_32455,N_32239);
and U35840 (N_35840,N_31095,N_33083);
nor U35841 (N_35841,N_34524,N_33828);
nor U35842 (N_35842,N_32854,N_34834);
nor U35843 (N_35843,N_34172,N_31052);
and U35844 (N_35844,N_31795,N_30511);
and U35845 (N_35845,N_31414,N_33470);
xnor U35846 (N_35846,N_31607,N_30942);
and U35847 (N_35847,N_34237,N_33266);
xor U35848 (N_35848,N_33647,N_34718);
and U35849 (N_35849,N_32260,N_33696);
or U35850 (N_35850,N_32376,N_30959);
or U35851 (N_35851,N_31707,N_31712);
nand U35852 (N_35852,N_32445,N_31107);
xor U35853 (N_35853,N_30184,N_32279);
xor U35854 (N_35854,N_30049,N_31529);
and U35855 (N_35855,N_34895,N_34737);
nand U35856 (N_35856,N_33927,N_30954);
nor U35857 (N_35857,N_31891,N_30231);
xnor U35858 (N_35858,N_34520,N_32574);
xor U35859 (N_35859,N_30773,N_30603);
xor U35860 (N_35860,N_31370,N_34238);
or U35861 (N_35861,N_30447,N_34789);
or U35862 (N_35862,N_32965,N_34691);
xor U35863 (N_35863,N_30668,N_34899);
nand U35864 (N_35864,N_33094,N_34446);
nand U35865 (N_35865,N_32169,N_32542);
nand U35866 (N_35866,N_34614,N_33324);
nor U35867 (N_35867,N_32336,N_33545);
or U35868 (N_35868,N_33831,N_30327);
or U35869 (N_35869,N_30664,N_34036);
nor U35870 (N_35870,N_30660,N_34509);
nor U35871 (N_35871,N_32299,N_30156);
or U35872 (N_35872,N_31685,N_33229);
xnor U35873 (N_35873,N_32164,N_30976);
or U35874 (N_35874,N_32773,N_30545);
and U35875 (N_35875,N_30788,N_33912);
nor U35876 (N_35876,N_30560,N_31450);
and U35877 (N_35877,N_34928,N_31029);
xnor U35878 (N_35878,N_31093,N_31229);
or U35879 (N_35879,N_32973,N_33553);
xor U35880 (N_35880,N_30364,N_34215);
nand U35881 (N_35881,N_31479,N_34216);
or U35882 (N_35882,N_31787,N_30886);
nand U35883 (N_35883,N_34443,N_32942);
xor U35884 (N_35884,N_32620,N_30688);
nand U35885 (N_35885,N_31890,N_32833);
or U35886 (N_35886,N_34484,N_32806);
nor U35887 (N_35887,N_32000,N_32458);
or U35888 (N_35888,N_30210,N_32552);
nor U35889 (N_35889,N_33806,N_33198);
nor U35890 (N_35890,N_30713,N_34015);
xor U35891 (N_35891,N_34610,N_33549);
nand U35892 (N_35892,N_31495,N_32446);
or U35893 (N_35893,N_32619,N_31510);
nor U35894 (N_35894,N_31341,N_33294);
nand U35895 (N_35895,N_33881,N_32832);
xnor U35896 (N_35896,N_33603,N_33065);
or U35897 (N_35897,N_33466,N_34365);
xor U35898 (N_35898,N_30185,N_34641);
xor U35899 (N_35899,N_31308,N_32605);
xnor U35900 (N_35900,N_31969,N_34887);
xor U35901 (N_35901,N_30153,N_31804);
or U35902 (N_35902,N_32600,N_34133);
or U35903 (N_35903,N_34361,N_32601);
or U35904 (N_35904,N_31749,N_33544);
nand U35905 (N_35905,N_32880,N_32474);
xnor U35906 (N_35906,N_31378,N_32152);
nor U35907 (N_35907,N_31040,N_31471);
or U35908 (N_35908,N_32515,N_30003);
or U35909 (N_35909,N_32178,N_33296);
nor U35910 (N_35910,N_31429,N_34089);
nor U35911 (N_35911,N_30244,N_33933);
or U35912 (N_35912,N_32578,N_31176);
and U35913 (N_35913,N_32598,N_34305);
and U35914 (N_35914,N_33893,N_31610);
nand U35915 (N_35915,N_31544,N_34715);
nand U35916 (N_35916,N_33522,N_30421);
or U35917 (N_35917,N_32405,N_31153);
nand U35918 (N_35918,N_34152,N_32238);
xor U35919 (N_35919,N_31888,N_31022);
xor U35920 (N_35920,N_32442,N_34769);
or U35921 (N_35921,N_33957,N_34623);
or U35922 (N_35922,N_34998,N_33329);
and U35923 (N_35923,N_33191,N_34473);
and U35924 (N_35924,N_32547,N_32780);
xnor U35925 (N_35925,N_34289,N_32650);
nand U35926 (N_35926,N_32179,N_34784);
nor U35927 (N_35927,N_34529,N_33132);
or U35928 (N_35928,N_32813,N_30750);
nand U35929 (N_35929,N_30996,N_34134);
nand U35930 (N_35930,N_30455,N_33525);
or U35931 (N_35931,N_34372,N_34956);
xnor U35932 (N_35932,N_31709,N_30459);
nor U35933 (N_35933,N_33818,N_32877);
nor U35934 (N_35934,N_30349,N_30827);
nor U35935 (N_35935,N_34023,N_33405);
xnor U35936 (N_35936,N_30363,N_34977);
nor U35937 (N_35937,N_34095,N_31779);
and U35938 (N_35938,N_34600,N_30222);
nand U35939 (N_35939,N_33138,N_32161);
nor U35940 (N_35940,N_31887,N_32791);
nand U35941 (N_35941,N_30556,N_34144);
nand U35942 (N_35942,N_33320,N_31413);
nor U35943 (N_35943,N_34982,N_34796);
xor U35944 (N_35944,N_31306,N_30127);
nor U35945 (N_35945,N_34539,N_30380);
nor U35946 (N_35946,N_34891,N_34702);
xor U35947 (N_35947,N_33165,N_32094);
or U35948 (N_35948,N_31858,N_34059);
xor U35949 (N_35949,N_34705,N_32712);
and U35950 (N_35950,N_31242,N_34202);
and U35951 (N_35951,N_32365,N_31003);
and U35952 (N_35952,N_30026,N_32682);
or U35953 (N_35953,N_32220,N_33586);
nand U35954 (N_35954,N_34005,N_31477);
or U35955 (N_35955,N_32869,N_32622);
xor U35956 (N_35956,N_34648,N_34357);
nand U35957 (N_35957,N_33344,N_34475);
nand U35958 (N_35958,N_34434,N_33760);
nand U35959 (N_35959,N_33048,N_33124);
and U35960 (N_35960,N_31201,N_34482);
nor U35961 (N_35961,N_33012,N_31695);
and U35962 (N_35962,N_32591,N_31801);
and U35963 (N_35963,N_32394,N_33714);
xor U35964 (N_35964,N_30715,N_31067);
and U35965 (N_35965,N_32739,N_31869);
xor U35966 (N_35966,N_33943,N_32244);
nor U35967 (N_35967,N_34203,N_31597);
xnor U35968 (N_35968,N_34993,N_34424);
or U35969 (N_35969,N_30172,N_34180);
nand U35970 (N_35970,N_34766,N_33250);
or U35971 (N_35971,N_33777,N_33891);
and U35972 (N_35972,N_33411,N_31798);
nand U35973 (N_35973,N_31277,N_33060);
or U35974 (N_35974,N_33193,N_30027);
and U35975 (N_35975,N_33310,N_32095);
nand U35976 (N_35976,N_30855,N_32893);
or U35977 (N_35977,N_31818,N_34338);
and U35978 (N_35978,N_30196,N_31079);
nand U35979 (N_35979,N_33656,N_32019);
xor U35980 (N_35980,N_31286,N_31913);
nor U35981 (N_35981,N_30982,N_31943);
xor U35982 (N_35982,N_30623,N_30004);
and U35983 (N_35983,N_30883,N_33665);
and U35984 (N_35984,N_33543,N_34727);
nand U35985 (N_35985,N_30268,N_31011);
and U35986 (N_35986,N_31474,N_33649);
and U35987 (N_35987,N_34346,N_33101);
nand U35988 (N_35988,N_32782,N_33503);
xor U35989 (N_35989,N_32920,N_31898);
and U35990 (N_35990,N_30837,N_34291);
nand U35991 (N_35991,N_30438,N_30882);
nor U35992 (N_35992,N_31590,N_30093);
or U35993 (N_35993,N_30276,N_34485);
or U35994 (N_35994,N_33381,N_34570);
and U35995 (N_35995,N_31186,N_31539);
or U35996 (N_35996,N_32399,N_31109);
and U35997 (N_35997,N_34362,N_32590);
nor U35998 (N_35998,N_32300,N_33604);
and U35999 (N_35999,N_34506,N_31879);
nand U36000 (N_36000,N_33837,N_34301);
xor U36001 (N_36001,N_33817,N_33221);
nor U36002 (N_36002,N_32306,N_32539);
and U36003 (N_36003,N_34933,N_30847);
xnor U36004 (N_36004,N_30377,N_34273);
and U36005 (N_36005,N_34262,N_31526);
nor U36006 (N_36006,N_30709,N_31045);
xnor U36007 (N_36007,N_34198,N_33277);
or U36008 (N_36008,N_31357,N_31528);
and U36009 (N_36009,N_34609,N_32011);
or U36010 (N_36010,N_30267,N_30151);
nor U36011 (N_36011,N_30841,N_34839);
nor U36012 (N_36012,N_31790,N_33289);
nand U36013 (N_36013,N_32776,N_32961);
or U36014 (N_36014,N_32350,N_33862);
nor U36015 (N_36015,N_34527,N_33974);
and U36016 (N_36016,N_30865,N_33281);
nand U36017 (N_36017,N_32785,N_31743);
xor U36018 (N_36018,N_33374,N_34604);
and U36019 (N_36019,N_31983,N_32879);
nor U36020 (N_36020,N_32757,N_31785);
nand U36021 (N_36021,N_33576,N_33994);
nand U36022 (N_36022,N_32589,N_30940);
nand U36023 (N_36023,N_30590,N_32354);
and U36024 (N_36024,N_30233,N_32216);
and U36025 (N_36025,N_34788,N_31086);
xnor U36026 (N_36026,N_32170,N_34825);
nand U36027 (N_36027,N_33899,N_31659);
xor U36028 (N_36028,N_32594,N_32715);
or U36029 (N_36029,N_34496,N_34139);
and U36030 (N_36030,N_34391,N_32802);
nand U36031 (N_36031,N_31114,N_33801);
or U36032 (N_36032,N_33051,N_33492);
nand U36033 (N_36033,N_30224,N_34432);
and U36034 (N_36034,N_32288,N_34279);
and U36035 (N_36035,N_34674,N_33435);
nor U36036 (N_36036,N_31697,N_31440);
xnor U36037 (N_36037,N_34012,N_31959);
nor U36038 (N_36038,N_30955,N_32390);
xor U36039 (N_36039,N_32248,N_33276);
or U36040 (N_36040,N_34630,N_32057);
and U36041 (N_36041,N_32859,N_31632);
and U36042 (N_36042,N_30471,N_34892);
and U36043 (N_36043,N_34882,N_31700);
nor U36044 (N_36044,N_33497,N_33148);
and U36045 (N_36045,N_34924,N_34109);
or U36046 (N_36046,N_32139,N_32194);
nor U36047 (N_36047,N_30236,N_30056);
xor U36048 (N_36048,N_31860,N_30202);
xor U36049 (N_36049,N_34439,N_34415);
xnor U36050 (N_36050,N_33699,N_32837);
xor U36051 (N_36051,N_31901,N_32464);
nor U36052 (N_36052,N_30020,N_33713);
xor U36053 (N_36053,N_32502,N_32753);
or U36054 (N_36054,N_33596,N_31900);
or U36055 (N_36055,N_31548,N_34003);
and U36056 (N_36056,N_30096,N_33389);
or U36057 (N_36057,N_34723,N_34130);
nor U36058 (N_36058,N_32289,N_34757);
nand U36059 (N_36059,N_34739,N_31144);
nor U36060 (N_36060,N_31377,N_31002);
xor U36061 (N_36061,N_31911,N_31765);
xnor U36062 (N_36062,N_31662,N_30158);
xor U36063 (N_36063,N_31182,N_33099);
nand U36064 (N_36064,N_32928,N_31663);
xnor U36065 (N_36065,N_31416,N_34417);
nand U36066 (N_36066,N_31728,N_34056);
and U36067 (N_36067,N_33188,N_33967);
or U36068 (N_36068,N_34991,N_33425);
and U36069 (N_36069,N_32371,N_32848);
nor U36070 (N_36070,N_32907,N_30916);
xnor U36071 (N_36071,N_31740,N_33244);
and U36072 (N_36072,N_32988,N_34541);
or U36073 (N_36073,N_32937,N_34830);
nand U36074 (N_36074,N_34663,N_30646);
nor U36075 (N_36075,N_30330,N_32207);
nand U36076 (N_36076,N_33225,N_31925);
and U36077 (N_36077,N_34664,N_31902);
and U36078 (N_36078,N_34166,N_32626);
or U36079 (N_36079,N_34632,N_32107);
xor U36080 (N_36080,N_32010,N_34408);
nand U36081 (N_36081,N_32554,N_34105);
nand U36082 (N_36082,N_34696,N_30730);
or U36083 (N_36083,N_30546,N_32992);
and U36084 (N_36084,N_34775,N_30393);
or U36085 (N_36085,N_33963,N_34867);
nor U36086 (N_36086,N_33258,N_31601);
nand U36087 (N_36087,N_33141,N_30881);
nand U36088 (N_36088,N_30030,N_34563);
and U36089 (N_36089,N_31106,N_33314);
nor U36090 (N_36090,N_34700,N_30939);
or U36091 (N_36091,N_34503,N_31419);
or U36092 (N_36092,N_32205,N_30984);
or U36093 (N_36093,N_30396,N_34302);
nand U36094 (N_36094,N_30932,N_30102);
and U36095 (N_36095,N_31794,N_34131);
and U36096 (N_36096,N_32027,N_33346);
and U36097 (N_36097,N_30573,N_34729);
or U36098 (N_36098,N_34862,N_30746);
xor U36099 (N_36099,N_31439,N_32466);
nand U36100 (N_36100,N_30638,N_30087);
nor U36101 (N_36101,N_31042,N_32633);
and U36102 (N_36102,N_34342,N_30070);
xor U36103 (N_36103,N_31505,N_31274);
or U36104 (N_36104,N_31380,N_32765);
nor U36105 (N_36105,N_31512,N_31953);
nand U36106 (N_36106,N_31248,N_33678);
nand U36107 (N_36107,N_32014,N_30216);
nor U36108 (N_36108,N_31636,N_33703);
and U36109 (N_36109,N_30441,N_30255);
nor U36110 (N_36110,N_32944,N_31720);
nor U36111 (N_36111,N_33609,N_30953);
nand U36112 (N_36112,N_34944,N_32536);
nor U36113 (N_36113,N_34908,N_30731);
nand U36114 (N_36114,N_32811,N_32351);
xnor U36115 (N_36115,N_34284,N_30311);
nand U36116 (N_36116,N_33701,N_30880);
nor U36117 (N_36117,N_34153,N_33973);
or U36118 (N_36118,N_33213,N_30386);
or U36119 (N_36119,N_31627,N_30280);
and U36120 (N_36120,N_30609,N_30074);
nor U36121 (N_36121,N_30170,N_33547);
xnor U36122 (N_36122,N_34234,N_30729);
and U36123 (N_36123,N_34300,N_30517);
and U36124 (N_36124,N_32904,N_34957);
nor U36125 (N_36125,N_31047,N_34400);
nor U36126 (N_36126,N_34937,N_33650);
and U36127 (N_36127,N_34274,N_34429);
nand U36128 (N_36128,N_34693,N_32512);
or U36129 (N_36129,N_32658,N_32443);
nor U36130 (N_36130,N_32296,N_30310);
or U36131 (N_36131,N_30907,N_30493);
or U36132 (N_36132,N_34287,N_31611);
nand U36133 (N_36133,N_32269,N_34008);
or U36134 (N_36134,N_31725,N_33372);
nand U36135 (N_36135,N_34707,N_34099);
or U36136 (N_36136,N_33116,N_30817);
and U36137 (N_36137,N_30281,N_31008);
and U36138 (N_36138,N_30998,N_32024);
and U36139 (N_36139,N_30894,N_34031);
and U36140 (N_36140,N_34689,N_31977);
or U36141 (N_36141,N_30383,N_34973);
and U36142 (N_36142,N_32892,N_34803);
and U36143 (N_36143,N_33856,N_31713);
nor U36144 (N_36144,N_33981,N_32077);
nand U36145 (N_36145,N_31897,N_34681);
and U36146 (N_36146,N_33010,N_31759);
and U36147 (N_36147,N_32517,N_30025);
and U36148 (N_36148,N_32338,N_30395);
or U36149 (N_36149,N_30115,N_31681);
nor U36150 (N_36150,N_33171,N_33074);
or U36151 (N_36151,N_32636,N_30107);
and U36152 (N_36152,N_32497,N_34421);
or U36153 (N_36153,N_32729,N_30207);
nand U36154 (N_36154,N_30130,N_30464);
xnor U36155 (N_36155,N_30611,N_33869);
nor U36156 (N_36156,N_32040,N_34328);
nand U36157 (N_36157,N_34537,N_32025);
or U36158 (N_36158,N_30891,N_30526);
xnor U36159 (N_36159,N_30290,N_31637);
or U36160 (N_36160,N_30462,N_34048);
xnor U36161 (N_36161,N_30427,N_32847);
xor U36162 (N_36162,N_30299,N_31444);
nand U36163 (N_36163,N_33847,N_31957);
nand U36164 (N_36164,N_30439,N_33711);
nand U36165 (N_36165,N_30926,N_32976);
or U36166 (N_36166,N_34077,N_32246);
nand U36167 (N_36167,N_30613,N_31173);
and U36168 (N_36168,N_32710,N_34765);
xor U36169 (N_36169,N_34961,N_31974);
nand U36170 (N_36170,N_30016,N_31940);
and U36171 (N_36171,N_32688,N_32387);
and U36172 (N_36172,N_31993,N_30803);
or U36173 (N_36173,N_34314,N_32132);
nand U36174 (N_36174,N_31298,N_30204);
and U36175 (N_36175,N_30830,N_32841);
xnor U36176 (N_36176,N_30423,N_30350);
xor U36177 (N_36177,N_34732,N_31623);
and U36178 (N_36178,N_34345,N_31631);
or U36179 (N_36179,N_34823,N_31238);
or U36180 (N_36180,N_30075,N_30186);
nor U36181 (N_36181,N_30694,N_31001);
xor U36182 (N_36182,N_34335,N_32851);
or U36183 (N_36183,N_34233,N_32903);
nand U36184 (N_36184,N_30769,N_34844);
xor U36185 (N_36185,N_33876,N_34946);
xnor U36186 (N_36186,N_34241,N_30288);
or U36187 (N_36187,N_34183,N_30319);
or U36188 (N_36188,N_31288,N_30182);
nor U36189 (N_36189,N_31464,N_31988);
or U36190 (N_36190,N_31006,N_32258);
xnor U36191 (N_36191,N_33278,N_32492);
nor U36192 (N_36192,N_30062,N_31808);
or U36193 (N_36193,N_33410,N_30856);
xnor U36194 (N_36194,N_30458,N_30465);
or U36195 (N_36195,N_32836,N_30229);
and U36196 (N_36196,N_34611,N_31540);
and U36197 (N_36197,N_34985,N_33373);
nor U36198 (N_36198,N_33805,N_32664);
or U36199 (N_36199,N_31606,N_32463);
xnor U36200 (N_36200,N_33515,N_31683);
nand U36201 (N_36201,N_32236,N_32672);
nand U36202 (N_36202,N_30264,N_32021);
or U36203 (N_36203,N_32653,N_30572);
or U36204 (N_36204,N_32652,N_30655);
or U36205 (N_36205,N_34081,N_32345);
nand U36206 (N_36206,N_33861,N_34352);
or U36207 (N_36207,N_32576,N_33797);
or U36208 (N_36208,N_33335,N_32128);
xnor U36209 (N_36209,N_32460,N_33183);
and U36210 (N_36210,N_32038,N_30478);
and U36211 (N_36211,N_33552,N_30242);
or U36212 (N_36212,N_33384,N_33392);
nand U36213 (N_36213,N_33111,N_32913);
nand U36214 (N_36214,N_30492,N_32769);
nand U36215 (N_36215,N_34748,N_33331);
nor U36216 (N_36216,N_31684,N_33535);
nand U36217 (N_36217,N_32076,N_34879);
or U36218 (N_36218,N_30676,N_31628);
or U36219 (N_36219,N_31219,N_33167);
nand U36220 (N_36220,N_31612,N_33773);
or U36221 (N_36221,N_33273,N_33747);
xor U36222 (N_36222,N_34690,N_33499);
or U36223 (N_36223,N_33415,N_33472);
nand U36224 (N_36224,N_34426,N_32899);
and U36225 (N_36225,N_32696,N_30159);
xor U36226 (N_36226,N_32453,N_34556);
nor U36227 (N_36227,N_31133,N_34210);
xnor U36228 (N_36228,N_31148,N_33902);
xor U36229 (N_36229,N_30644,N_32651);
xnor U36230 (N_36230,N_31692,N_33858);
nor U36231 (N_36231,N_31048,N_32113);
and U36232 (N_36232,N_33840,N_31848);
nor U36233 (N_36233,N_33293,N_30576);
xnor U36234 (N_36234,N_33559,N_33992);
or U36235 (N_36235,N_33014,N_32370);
xor U36236 (N_36236,N_33485,N_32519);
and U36237 (N_36237,N_33461,N_34889);
xnor U36238 (N_36238,N_34228,N_31543);
nor U36239 (N_36239,N_34376,N_33285);
and U36240 (N_36240,N_30258,N_34651);
nand U36241 (N_36241,N_31436,N_30785);
nor U36242 (N_36242,N_33049,N_31136);
and U36243 (N_36243,N_33962,N_31852);
or U36244 (N_36244,N_34363,N_30456);
nor U36245 (N_36245,N_34749,N_34064);
xor U36246 (N_36246,N_33062,N_32101);
nor U36247 (N_36247,N_32720,N_30842);
or U36248 (N_36248,N_30144,N_32634);
nand U36249 (N_36249,N_34117,N_34492);
nor U36250 (N_36250,N_30627,N_34793);
nand U36251 (N_36251,N_31930,N_31489);
nand U36252 (N_36252,N_30663,N_30980);
or U36253 (N_36253,N_34349,N_34914);
xor U36254 (N_36254,N_31735,N_33830);
nand U36255 (N_36255,N_31259,N_30876);
xnor U36256 (N_36256,N_32198,N_34155);
nor U36257 (N_36257,N_31417,N_31368);
and U36258 (N_36258,N_34451,N_31281);
or U36259 (N_36259,N_30259,N_33787);
nor U36260 (N_36260,N_32566,N_34070);
or U36261 (N_36261,N_33571,N_33342);
or U36262 (N_36262,N_30799,N_32898);
and U36263 (N_36263,N_32822,N_32187);
nand U36264 (N_36264,N_34948,N_33462);
nor U36265 (N_36265,N_33457,N_33482);
xor U36266 (N_36266,N_33234,N_34045);
nand U36267 (N_36267,N_30850,N_31776);
and U36268 (N_36268,N_32985,N_32090);
xor U36269 (N_36269,N_34072,N_34150);
nand U36270 (N_36270,N_31223,N_33990);
xor U36271 (N_36271,N_32126,N_31190);
nor U36272 (N_36272,N_31245,N_32237);
or U36273 (N_36273,N_33832,N_30951);
and U36274 (N_36274,N_34510,N_32359);
xor U36275 (N_36275,N_30587,N_32817);
nand U36276 (N_36276,N_34958,N_33996);
xnor U36277 (N_36277,N_31160,N_34730);
nor U36278 (N_36278,N_32084,N_32895);
nor U36279 (N_36279,N_31603,N_34699);
and U36280 (N_36280,N_34831,N_30109);
and U36281 (N_36281,N_31183,N_33307);
xor U36282 (N_36282,N_30119,N_32862);
nor U36283 (N_36283,N_33737,N_32681);
nor U36284 (N_36284,N_33931,N_30902);
xnor U36285 (N_36285,N_34497,N_31918);
and U36286 (N_36286,N_31841,N_33886);
and U36287 (N_36287,N_34672,N_32800);
nand U36288 (N_36288,N_33253,N_33471);
or U36289 (N_36289,N_30469,N_33112);
nor U36290 (N_36290,N_32439,N_30125);
xnor U36291 (N_36291,N_30321,N_32556);
and U36292 (N_36292,N_34754,N_32424);
nand U36293 (N_36293,N_31586,N_33530);
xnor U36294 (N_36294,N_34930,N_31521);
nand U36295 (N_36295,N_34770,N_30787);
nor U36296 (N_36296,N_31063,N_32541);
nor U36297 (N_36297,N_32284,N_33483);
and U36298 (N_36298,N_33033,N_30183);
nand U36299 (N_36299,N_30217,N_33089);
or U36300 (N_36300,N_32968,N_31038);
or U36301 (N_36301,N_31430,N_32709);
nand U36302 (N_36302,N_34695,N_31375);
and U36303 (N_36303,N_33821,N_34406);
or U36304 (N_36304,N_31719,N_33045);
nand U36305 (N_36305,N_34491,N_34107);
and U36306 (N_36306,N_30581,N_34019);
or U36307 (N_36307,N_32465,N_33850);
nand U36308 (N_36308,N_30553,N_34661);
nor U36309 (N_36309,N_32393,N_32427);
nor U36310 (N_36310,N_30473,N_34259);
xnor U36311 (N_36311,N_34122,N_30840);
nor U36312 (N_36312,N_32641,N_31010);
or U36313 (N_36313,N_33206,N_30716);
nand U36314 (N_36314,N_31249,N_31731);
xnor U36315 (N_36315,N_30642,N_31158);
or U36316 (N_36316,N_30727,N_31459);
or U36317 (N_36317,N_32889,N_33495);
nand U36318 (N_36318,N_31752,N_32031);
nor U36319 (N_36319,N_34735,N_34033);
xor U36320 (N_36320,N_32123,N_32684);
nand U36321 (N_36321,N_33036,N_31562);
nand U36322 (N_36322,N_33439,N_30822);
nor U36323 (N_36323,N_31142,N_31208);
nand U36324 (N_36324,N_30801,N_34399);
nand U36325 (N_36325,N_31594,N_33412);
nand U36326 (N_36326,N_32007,N_34027);
xor U36327 (N_36327,N_31015,N_33484);
nor U36328 (N_36328,N_33061,N_30437);
or U36329 (N_36329,N_30875,N_31422);
nand U36330 (N_36330,N_34458,N_30790);
xnor U36331 (N_36331,N_32104,N_31203);
nand U36332 (N_36332,N_31088,N_34926);
or U36333 (N_36333,N_33219,N_30346);
nor U36334 (N_36334,N_33274,N_33078);
nor U36335 (N_36335,N_31582,N_31031);
nor U36336 (N_36336,N_34088,N_30657);
or U36337 (N_36337,N_33459,N_33364);
nand U36338 (N_36338,N_31279,N_31012);
and U36339 (N_36339,N_32222,N_30794);
xnor U36340 (N_36340,N_33166,N_31120);
xor U36341 (N_36341,N_31886,N_30925);
xnor U36342 (N_36342,N_33030,N_30240);
nand U36343 (N_36343,N_31652,N_30190);
and U36344 (N_36344,N_32830,N_30325);
nor U36345 (N_36345,N_34588,N_30295);
or U36346 (N_36346,N_30640,N_34179);
or U36347 (N_36347,N_30032,N_33303);
nor U36348 (N_36348,N_32362,N_34098);
nor U36349 (N_36349,N_32857,N_33732);
nand U36350 (N_36350,N_33021,N_30152);
nand U36351 (N_36351,N_33622,N_33942);
nand U36352 (N_36352,N_34495,N_32801);
or U36353 (N_36353,N_33243,N_31971);
nand U36354 (N_36354,N_31401,N_32616);
or U36355 (N_36355,N_33717,N_34138);
xor U36356 (N_36356,N_32567,N_33018);
and U36357 (N_36357,N_33507,N_34042);
nor U36358 (N_36358,N_33645,N_32434);
xor U36359 (N_36359,N_30928,N_33404);
nand U36360 (N_36360,N_30528,N_31667);
nor U36361 (N_36361,N_31155,N_33154);
or U36362 (N_36362,N_30339,N_30619);
and U36363 (N_36363,N_30810,N_31672);
nand U36364 (N_36364,N_31385,N_33080);
nand U36365 (N_36365,N_32298,N_31525);
or U36366 (N_36366,N_34919,N_31615);
nand U36367 (N_36367,N_31678,N_31941);
xor U36368 (N_36368,N_32384,N_31434);
nand U36369 (N_36369,N_33924,N_31299);
and U36370 (N_36370,N_30048,N_32277);
nor U36371 (N_36371,N_34906,N_31073);
or U36372 (N_36372,N_33236,N_32001);
xor U36373 (N_36373,N_34057,N_30333);
nand U36374 (N_36374,N_31409,N_34531);
and U36375 (N_36375,N_34470,N_32138);
xnor U36376 (N_36376,N_31134,N_32039);
nand U36377 (N_36377,N_30345,N_31754);
or U36378 (N_36378,N_30128,N_32562);
or U36379 (N_36379,N_32313,N_31343);
and U36380 (N_36380,N_32982,N_30338);
nor U36381 (N_36381,N_33620,N_30647);
nor U36382 (N_36382,N_32755,N_33618);
nand U36383 (N_36383,N_34208,N_32058);
and U36384 (N_36384,N_32052,N_34489);
or U36385 (N_36385,N_31608,N_32259);
and U36386 (N_36386,N_31833,N_33600);
xnor U36387 (N_36387,N_33868,N_30741);
and U36388 (N_36388,N_33143,N_31310);
nand U36389 (N_36389,N_33349,N_33097);
xor U36390 (N_36390,N_30497,N_30759);
or U36391 (N_36391,N_32940,N_32456);
or U36392 (N_36392,N_32960,N_31005);
nor U36393 (N_36393,N_33491,N_33125);
or U36394 (N_36394,N_32809,N_31640);
and U36395 (N_36395,N_32073,N_32377);
nor U36396 (N_36396,N_34116,N_32674);
and U36397 (N_36397,N_31322,N_34638);
xor U36398 (N_36398,N_33173,N_31866);
xor U36399 (N_36399,N_32059,N_32956);
or U36400 (N_36400,N_33496,N_34055);
xor U36401 (N_36401,N_33506,N_34132);
and U36402 (N_36402,N_31085,N_33054);
nor U36403 (N_36403,N_32821,N_30124);
nand U36404 (N_36404,N_34344,N_32312);
and U36405 (N_36405,N_33479,N_33379);
nand U36406 (N_36406,N_33951,N_31549);
nor U36407 (N_36407,N_30970,N_32254);
nand U36408 (N_36408,N_33248,N_33922);
xnor U36409 (N_36409,N_30721,N_34868);
or U36410 (N_36410,N_32281,N_34759);
xnor U36411 (N_36411,N_32792,N_34435);
nand U36412 (N_36412,N_33803,N_33892);
or U36413 (N_36413,N_31152,N_31618);
and U36414 (N_36414,N_30950,N_32192);
nand U36415 (N_36415,N_31264,N_34884);
or U36416 (N_36416,N_30991,N_31035);
nor U36417 (N_36417,N_34201,N_30733);
xnor U36418 (N_36418,N_33783,N_30685);
and U36419 (N_36419,N_33834,N_33759);
and U36420 (N_36420,N_33779,N_30530);
nand U36421 (N_36421,N_31649,N_33144);
nor U36422 (N_36422,N_34308,N_33739);
xor U36423 (N_36423,N_33964,N_30935);
xor U36424 (N_36424,N_32790,N_30002);
nor U36425 (N_36425,N_31698,N_31180);
xor U36426 (N_36426,N_30059,N_31258);
nor U36427 (N_36427,N_34942,N_33380);
xor U36428 (N_36428,N_33780,N_33437);
and U36429 (N_36429,N_34358,N_31113);
or U36430 (N_36430,N_31212,N_30651);
and U36431 (N_36431,N_34987,N_34827);
nand U36432 (N_36432,N_31130,N_33001);
or U36433 (N_36433,N_31213,N_30414);
and U36434 (N_36434,N_30680,N_34603);
nand U36435 (N_36435,N_34780,N_31263);
nor U36436 (N_36436,N_32061,N_32657);
and U36437 (N_36437,N_34747,N_34319);
xnor U36438 (N_36438,N_30796,N_30307);
xor U36439 (N_36439,N_32738,N_31484);
and U36440 (N_36440,N_31545,N_33385);
nor U36441 (N_36441,N_34731,N_33481);
and U36442 (N_36442,N_33846,N_30390);
and U36443 (N_36443,N_34320,N_32034);
nand U36444 (N_36444,N_32217,N_33756);
nor U36445 (N_36445,N_32096,N_34326);
xnor U36446 (N_36446,N_34318,N_34852);
or U36447 (N_36447,N_33077,N_30399);
nor U36448 (N_36448,N_30738,N_31756);
xnor U36449 (N_36449,N_31420,N_30247);
or U36450 (N_36450,N_31467,N_30446);
xnor U36451 (N_36451,N_30418,N_34734);
or U36452 (N_36452,N_32389,N_32610);
xor U36453 (N_36453,N_31748,N_33546);
or U36454 (N_36454,N_32337,N_33339);
and U36455 (N_36455,N_33287,N_34447);
nand U36456 (N_36456,N_30009,N_32932);
or U36457 (N_36457,N_31546,N_33934);
nor U36458 (N_36458,N_34851,N_30909);
nor U36459 (N_36459,N_30336,N_34181);
nand U36460 (N_36460,N_33262,N_32623);
nor U36461 (N_36461,N_30639,N_34826);
or U36462 (N_36462,N_34146,N_30490);
nor U36463 (N_36463,N_32346,N_33498);
or U36464 (N_36464,N_32349,N_33282);
nand U36465 (N_36465,N_32498,N_33729);
or U36466 (N_36466,N_32789,N_31381);
nor U36467 (N_36467,N_32561,N_32270);
and U36468 (N_36468,N_32915,N_34791);
nand U36469 (N_36469,N_32675,N_31657);
nand U36470 (N_36470,N_33762,N_34808);
and U36471 (N_36471,N_32522,N_30176);
or U36472 (N_36472,N_34545,N_32401);
or U36473 (N_36473,N_33500,N_33257);
or U36474 (N_36474,N_33634,N_34962);
nand U36475 (N_36475,N_30422,N_33681);
xnor U36476 (N_36476,N_34188,N_31194);
nor U36477 (N_36477,N_33323,N_34369);
xnor U36478 (N_36478,N_32560,N_34586);
and U36479 (N_36479,N_33566,N_31722);
xor U36480 (N_36480,N_31751,N_32521);
and U36481 (N_36481,N_33316,N_31702);
nand U36482 (N_36482,N_33716,N_30667);
xor U36483 (N_36483,N_33237,N_30055);
and U36484 (N_36484,N_33441,N_34951);
nand U36485 (N_36485,N_32087,N_30039);
and U36486 (N_36486,N_34980,N_34474);
and U36487 (N_36487,N_31056,N_30990);
or U36488 (N_36488,N_31871,N_31914);
nor U36489 (N_36489,N_34979,N_34684);
nand U36490 (N_36490,N_33133,N_34135);
xor U36491 (N_36491,N_33367,N_33147);
xnor U36492 (N_36492,N_30046,N_30058);
xor U36493 (N_36493,N_33640,N_30964);
and U36494 (N_36494,N_30194,N_34379);
nand U36495 (N_36495,N_32408,N_32112);
nor U36496 (N_36496,N_31616,N_34207);
nor U36497 (N_36497,N_30635,N_31237);
nor U36498 (N_36498,N_34371,N_30893);
and U36499 (N_36499,N_33804,N_31990);
or U36500 (N_36500,N_32644,N_31563);
or U36501 (N_36501,N_33409,N_33641);
or U36502 (N_36502,N_34952,N_32784);
nor U36503 (N_36503,N_30720,N_32770);
xor U36504 (N_36504,N_30408,N_31604);
nand U36505 (N_36505,N_31371,N_34430);
nor U36506 (N_36506,N_30687,N_30463);
and U36507 (N_36507,N_34963,N_31244);
nor U36508 (N_36508,N_34129,N_32875);
nor U36509 (N_36509,N_31360,N_32746);
and U36510 (N_36510,N_33968,N_30273);
nor U36511 (N_36511,N_31285,N_34565);
xor U36512 (N_36512,N_30213,N_31449);
and U36513 (N_36513,N_33909,N_34075);
nor U36514 (N_36514,N_34686,N_31206);
and U36515 (N_36515,N_34433,N_31453);
and U36516 (N_36516,N_32452,N_33671);
nand U36517 (N_36517,N_31317,N_32310);
or U36518 (N_36518,N_30406,N_31473);
nand U36519 (N_36519,N_31811,N_30695);
and U36520 (N_36520,N_31853,N_32391);
nand U36521 (N_36521,N_30466,N_31179);
nor U36522 (N_36522,N_30050,N_32028);
nand U36523 (N_36523,N_31307,N_30337);
or U36524 (N_36524,N_32005,N_34022);
nand U36525 (N_36525,N_32803,N_30482);
nor U36526 (N_36526,N_30467,N_33160);
nand U36527 (N_36527,N_32936,N_31162);
and U36528 (N_36528,N_31846,N_33085);
xor U36529 (N_36529,N_34231,N_30086);
nor U36530 (N_36530,N_31714,N_33403);
or U36531 (N_36531,N_33245,N_30518);
xor U36532 (N_36532,N_31151,N_32280);
nor U36533 (N_36533,N_31626,N_32581);
nand U36534 (N_36534,N_30683,N_32701);
or U36535 (N_36535,N_33879,N_34092);
or U36536 (N_36536,N_30555,N_34923);
or U36537 (N_36537,N_31768,N_30326);
nand U36538 (N_36538,N_31292,N_33674);
and U36539 (N_36539,N_30304,N_32097);
and U36540 (N_36540,N_31656,N_34761);
nand U36541 (N_36541,N_30443,N_31856);
or U36542 (N_36542,N_31268,N_31132);
or U36543 (N_36543,N_31638,N_30249);
and U36544 (N_36544,N_33359,N_33863);
xnor U36545 (N_36545,N_30429,N_33929);
or U36546 (N_36546,N_30498,N_32747);
nor U36547 (N_36547,N_33026,N_30454);
or U36548 (N_36548,N_31166,N_33682);
or U36549 (N_36549,N_33844,N_33989);
nor U36550 (N_36550,N_32654,N_32897);
nand U36551 (N_36551,N_33685,N_32261);
and U36552 (N_36552,N_33669,N_33330);
or U36553 (N_36553,N_34528,N_32168);
xor U36554 (N_36554,N_33463,N_32588);
nor U36555 (N_36555,N_32008,N_31170);
xnor U36556 (N_36556,N_31518,N_33386);
xnor U36557 (N_36557,N_31337,N_34873);
and U36558 (N_36558,N_31661,N_33516);
or U36559 (N_36559,N_33982,N_34025);
or U36560 (N_36560,N_33315,N_32642);
or U36561 (N_36561,N_33567,N_31374);
or U36562 (N_36562,N_33630,N_34804);
nand U36563 (N_36563,N_30405,N_34106);
or U36564 (N_36564,N_30113,N_33590);
nor U36565 (N_36565,N_31016,N_31408);
or U36566 (N_36566,N_32335,N_32374);
and U36567 (N_36567,N_31710,N_30956);
or U36568 (N_36568,N_32311,N_30795);
and U36569 (N_36569,N_32334,N_33391);
nor U36570 (N_36570,N_33233,N_31686);
nor U36571 (N_36571,N_32812,N_32834);
xor U36572 (N_36572,N_33291,N_30412);
and U36573 (N_36573,N_30067,N_30981);
and U36574 (N_36574,N_33157,N_34370);
and U36575 (N_36575,N_32687,N_32910);
xnor U36576 (N_36576,N_32410,N_31105);
or U36577 (N_36577,N_34751,N_31129);
and U36578 (N_36578,N_30031,N_31156);
nor U36579 (N_36579,N_34786,N_30191);
or U36580 (N_36580,N_31760,N_32930);
and U36581 (N_36581,N_33038,N_34303);
nand U36582 (N_36582,N_34581,N_31767);
nand U36583 (N_36583,N_34965,N_30722);
nor U36584 (N_36584,N_33791,N_32722);
nor U36585 (N_36585,N_33280,N_33003);
or U36586 (N_36586,N_32614,N_30737);
nor U36587 (N_36587,N_34549,N_30136);
nor U36588 (N_36588,N_32125,N_32068);
nand U36589 (N_36589,N_32385,N_33115);
xor U36590 (N_36590,N_30993,N_32085);
and U36591 (N_36591,N_31340,N_33900);
or U36592 (N_36592,N_31734,N_33845);
or U36593 (N_36593,N_30015,N_30146);
or U36594 (N_36594,N_30919,N_31200);
or U36595 (N_36595,N_34925,N_32583);
or U36596 (N_36596,N_34828,N_31131);
nand U36597 (N_36597,N_34343,N_30496);
nor U36598 (N_36598,N_32959,N_31979);
or U36599 (N_36599,N_30661,N_33336);
nor U36600 (N_36600,N_30322,N_32386);
or U36601 (N_36601,N_30690,N_34932);
xnor U36602 (N_36602,N_34034,N_33152);
xnor U36603 (N_36603,N_30037,N_31863);
nand U36604 (N_36604,N_31511,N_33011);
nor U36605 (N_36605,N_33311,N_33137);
nand U36606 (N_36606,N_32487,N_34859);
nor U36607 (N_36607,N_34621,N_31797);
nand U36608 (N_36608,N_31741,N_30160);
nor U36609 (N_36609,N_30312,N_33864);
or U36610 (N_36610,N_30899,N_34293);
nand U36611 (N_36611,N_31101,N_33815);
and U36612 (N_36612,N_31880,N_33623);
nand U36613 (N_36613,N_33261,N_32361);
nand U36614 (N_36614,N_33970,N_30266);
or U36615 (N_36615,N_30525,N_33371);
xor U36616 (N_36616,N_31352,N_32319);
nor U36617 (N_36617,N_30544,N_32462);
nor U36618 (N_36618,N_34165,N_34653);
nand U36619 (N_36619,N_30513,N_31810);
nor U36620 (N_36620,N_32332,N_33976);
or U36621 (N_36621,N_31290,N_34271);
xnor U36622 (N_36622,N_30756,N_33309);
nand U36623 (N_36623,N_33016,N_34519);
or U36624 (N_36624,N_31044,N_31463);
or U36625 (N_36625,N_30569,N_33272);
nor U36626 (N_36626,N_31929,N_34148);
or U36627 (N_36627,N_31926,N_34776);
xor U36628 (N_36628,N_30316,N_32301);
or U36629 (N_36629,N_31427,N_34288);
or U36630 (N_36630,N_32341,N_32996);
or U36631 (N_36631,N_34622,N_32831);
or U36632 (N_36632,N_30742,N_34377);
xnor U36633 (N_36633,N_32577,N_31344);
nand U36634 (N_36634,N_32706,N_33997);
and U36635 (N_36635,N_33978,N_32545);
xnor U36636 (N_36636,N_33275,N_33823);
xnor U36637 (N_36637,N_32509,N_33071);
or U36638 (N_36638,N_32177,N_34724);
and U36639 (N_36639,N_33464,N_33907);
xnor U36640 (N_36640,N_32717,N_33127);
or U36641 (N_36641,N_34855,N_34121);
and U36642 (N_36642,N_34350,N_31432);
nor U36643 (N_36643,N_32917,N_34888);
and U36644 (N_36644,N_32046,N_34922);
nand U36645 (N_36645,N_34281,N_32225);
nand U36646 (N_36646,N_34442,N_30248);
nand U36647 (N_36647,N_31192,N_33949);
nor U36648 (N_36648,N_30562,N_33615);
xnor U36649 (N_36649,N_33985,N_34246);
or U36650 (N_36650,N_34876,N_32471);
nor U36651 (N_36651,N_32409,N_31541);
or U36652 (N_36652,N_32240,N_32516);
xor U36653 (N_36653,N_30924,N_31536);
or U36654 (N_36654,N_32999,N_31517);
nand U36655 (N_36655,N_32793,N_30479);
nand U36656 (N_36656,N_31729,N_31660);
xnor U36657 (N_36657,N_30755,N_30922);
xor U36658 (N_36658,N_31117,N_30352);
and U36659 (N_36659,N_30154,N_32850);
xor U36660 (N_36660,N_34813,N_34559);
and U36661 (N_36661,N_31443,N_32291);
or U36662 (N_36662,N_32062,N_30870);
nand U36663 (N_36663,N_33448,N_30101);
or U36664 (N_36664,N_31428,N_30035);
nand U36665 (N_36665,N_31591,N_32273);
nor U36666 (N_36666,N_34375,N_31049);
or U36667 (N_36667,N_33218,N_30042);
nand U36668 (N_36668,N_31629,N_33375);
xor U36669 (N_36669,N_31261,N_34038);
nor U36670 (N_36670,N_32983,N_34066);
and U36671 (N_36671,N_33238,N_34256);
nand U36672 (N_36672,N_30816,N_33774);
xnor U36673 (N_36673,N_34523,N_30008);
xor U36674 (N_36674,N_30818,N_33423);
nor U36675 (N_36675,N_33660,N_30477);
or U36676 (N_36676,N_30243,N_31694);
and U36677 (N_36677,N_34490,N_30092);
nand U36678 (N_36678,N_34768,N_34943);
or U36679 (N_36679,N_31733,N_31773);
nand U36680 (N_36680,N_30890,N_30740);
nand U36681 (N_36681,N_31411,N_30385);
and U36682 (N_36682,N_30365,N_31831);
nor U36683 (N_36683,N_32407,N_34438);
and U36684 (N_36684,N_30969,N_32518);
nor U36685 (N_36685,N_30283,N_33772);
or U36686 (N_36686,N_31202,N_30859);
xor U36687 (N_36687,N_33613,N_30199);
and U36688 (N_36688,N_30778,N_34476);
or U36689 (N_36689,N_31061,N_34746);
nor U36690 (N_36690,N_31221,N_34901);
nand U36691 (N_36691,N_31291,N_32724);
and U36692 (N_36692,N_32406,N_33606);
and U36693 (N_36693,N_33004,N_33742);
nor U36694 (N_36694,N_34571,N_33521);
nand U36695 (N_36695,N_30862,N_34975);
and U36696 (N_36696,N_34508,N_34598);
and U36697 (N_36697,N_34814,N_33684);
or U36698 (N_36698,N_30585,N_32314);
nand U36699 (N_36699,N_31090,N_32148);
nor U36700 (N_36700,N_33121,N_34819);
nor U36701 (N_36701,N_33420,N_32166);
and U36702 (N_36702,N_33387,N_32461);
nor U36703 (N_36703,N_31812,N_31965);
nand U36704 (N_36704,N_31867,N_31625);
or U36705 (N_36705,N_33327,N_30670);
nor U36706 (N_36706,N_33456,N_31955);
nor U36707 (N_36707,N_33940,N_33866);
nor U36708 (N_36708,N_31100,N_33122);
nor U36709 (N_36709,N_31847,N_30774);
xor U36710 (N_36710,N_32223,N_34323);
xnor U36711 (N_36711,N_30505,N_30807);
and U36712 (N_36712,N_30570,N_34802);
xnor U36713 (N_36713,N_31059,N_32690);
xnor U36714 (N_36714,N_34918,N_32689);
and U36715 (N_36715,N_34374,N_34903);
nor U36716 (N_36716,N_31592,N_32927);
nor U36717 (N_36717,N_30083,N_31750);
xnor U36718 (N_36718,N_34596,N_32201);
and U36719 (N_36719,N_34569,N_30944);
or U36720 (N_36720,N_31256,N_33118);
xnor U36721 (N_36721,N_31111,N_34625);
and U36722 (N_36722,N_32404,N_32948);
and U36723 (N_36723,N_31376,N_34712);
nor U36724 (N_36724,N_31665,N_33741);
xor U36725 (N_36725,N_30838,N_31104);
and U36726 (N_36726,N_30100,N_33833);
and U36727 (N_36727,N_31908,N_31331);
and U36728 (N_36728,N_31679,N_30751);
xor U36729 (N_36729,N_31363,N_34104);
xor U36730 (N_36730,N_34263,N_33308);
nor U36731 (N_36731,N_31991,N_30011);
or U36732 (N_36732,N_34913,N_33839);
nor U36733 (N_36733,N_32508,N_33035);
or U36734 (N_36734,N_33178,N_31580);
and U36735 (N_36735,N_30072,N_32794);
nor U36736 (N_36736,N_33572,N_31581);
and U36737 (N_36737,N_32499,N_34620);
and U36738 (N_36738,N_30804,N_31981);
and U36739 (N_36739,N_34915,N_34967);
or U36740 (N_36740,N_30872,N_32506);
xnor U36741 (N_36741,N_30407,N_30618);
or U36742 (N_36742,N_32421,N_30726);
or U36743 (N_36743,N_33009,N_30948);
xor U36744 (N_36744,N_30309,N_30301);
nor U36745 (N_36745,N_32056,N_34071);
and U36746 (N_36746,N_32328,N_32767);
nor U36747 (N_36747,N_33288,N_33827);
nand U36748 (N_36748,N_34745,N_33180);
xor U36749 (N_36749,N_32530,N_33255);
and U36750 (N_36750,N_32190,N_30073);
or U36751 (N_36751,N_31032,N_32764);
nor U36752 (N_36752,N_31267,N_30293);
or U36753 (N_36753,N_30135,N_31836);
nor U36754 (N_36754,N_34553,N_30947);
and U36755 (N_36755,N_33822,N_31992);
xnor U36756 (N_36756,N_31827,N_33539);
or U36757 (N_36757,N_32186,N_33422);
nor U36758 (N_36758,N_31425,N_34694);
xnor U36759 (N_36759,N_33079,N_34185);
xnor U36760 (N_36760,N_31997,N_33008);
or U36761 (N_36761,N_33408,N_32357);
nand U36762 (N_36762,N_33915,N_31984);
nand U36763 (N_36763,N_32871,N_30188);
nor U36764 (N_36764,N_32513,N_31699);
and U36765 (N_36765,N_31004,N_31830);
xor U36766 (N_36766,N_31278,N_31556);
nand U36767 (N_36767,N_34007,N_33748);
nand U36768 (N_36768,N_34938,N_32100);
or U36769 (N_36769,N_33247,N_32649);
xor U36770 (N_36770,N_32415,N_31312);
xor U36771 (N_36771,N_33601,N_33877);
or U36772 (N_36772,N_32564,N_34647);
and U36773 (N_36773,N_34778,N_32130);
or U36774 (N_36774,N_30887,N_30677);
nor U36775 (N_36775,N_34969,N_33469);
nand U36776 (N_36776,N_31904,N_30992);
xor U36777 (N_36777,N_31820,N_31354);
nand U36778 (N_36778,N_32925,N_30200);
xor U36779 (N_36779,N_30044,N_31789);
nor U36780 (N_36780,N_34060,N_32287);
or U36781 (N_36781,N_31881,N_34178);
nor U36782 (N_36782,N_33271,N_31958);
or U36783 (N_36783,N_32867,N_34452);
and U36784 (N_36784,N_31999,N_32167);
and U36785 (N_36785,N_34211,N_33177);
xnor U36786 (N_36786,N_33766,N_33321);
and U36787 (N_36787,N_31097,N_34909);
nand U36788 (N_36788,N_32991,N_32185);
and U36789 (N_36789,N_32938,N_32418);
or U36790 (N_36790,N_33402,N_31359);
nor U36791 (N_36791,N_31519,N_34988);
or U36792 (N_36792,N_33819,N_33022);
xor U36793 (N_36793,N_32612,N_32661);
or U36794 (N_36794,N_31682,N_34564);
nor U36795 (N_36795,N_32013,N_30630);
xnor U36796 (N_36796,N_32484,N_32939);
nor U36797 (N_36797,N_30636,N_34989);
nor U36798 (N_36798,N_33860,N_31062);
xor U36799 (N_36799,N_34330,N_34501);
and U36800 (N_36800,N_33164,N_30900);
or U36801 (N_36801,N_31873,N_32816);
and U36802 (N_36802,N_30937,N_34500);
nor U36803 (N_36803,N_34692,N_34886);
nor U36804 (N_36804,N_31177,N_30728);
or U36805 (N_36805,N_31676,N_32202);
xor U36806 (N_36806,N_30835,N_33651);
nor U36807 (N_36807,N_31335,N_34558);
or U36808 (N_36808,N_30736,N_32952);
or U36809 (N_36809,N_34052,N_33493);
nand U36810 (N_36810,N_32978,N_30557);
or U36811 (N_36811,N_31558,N_31721);
and U36812 (N_36812,N_32218,N_32969);
and U36813 (N_36813,N_33347,N_33795);
xor U36814 (N_36814,N_34436,N_32796);
nor U36815 (N_36815,N_34955,N_33332);
nand U36816 (N_36816,N_32344,N_33369);
and U36817 (N_36817,N_33736,N_33657);
or U36818 (N_36818,N_30826,N_32528);
nor U36819 (N_36819,N_30302,N_31823);
or U36820 (N_36820,N_33897,N_31348);
or U36821 (N_36821,N_32308,N_34840);
or U36822 (N_36822,N_32203,N_32676);
xnor U36823 (N_36823,N_31572,N_30444);
or U36824 (N_36824,N_34602,N_30155);
nor U36825 (N_36825,N_32358,N_32323);
nor U36826 (N_36826,N_33223,N_32568);
xor U36827 (N_36827,N_32860,N_30829);
nor U36828 (N_36828,N_34656,N_30529);
xor U36829 (N_36829,N_33172,N_34870);
and U36830 (N_36830,N_33510,N_32327);
nand U36831 (N_36831,N_33873,N_31730);
and U36832 (N_36832,N_30111,N_33950);
nand U36833 (N_36833,N_34667,N_32699);
or U36834 (N_36834,N_30033,N_34722);
nand U36835 (N_36835,N_34425,N_32721);
xnor U36836 (N_36836,N_34340,N_32926);
and U36837 (N_36837,N_34593,N_31921);
or U36838 (N_36838,N_31313,N_33735);
or U36839 (N_36839,N_34026,N_33195);
or U36840 (N_36840,N_33249,N_33551);
nand U36841 (N_36841,N_32824,N_34812);
or U36842 (N_36842,N_32063,N_31894);
or U36843 (N_36843,N_30809,N_30602);
nand U36844 (N_36844,N_31470,N_33070);
nand U36845 (N_36845,N_34966,N_34204);
nor U36846 (N_36846,N_32719,N_31395);
or U36847 (N_36847,N_30768,N_30700);
nor U36848 (N_36848,N_32400,N_31275);
nand U36849 (N_36849,N_34479,N_34533);
nor U36850 (N_36850,N_34728,N_32971);
nor U36851 (N_36851,N_34158,N_34420);
or U36852 (N_36852,N_34359,N_30786);
nand U36853 (N_36853,N_30442,N_32089);
nand U36854 (N_36854,N_31655,N_31944);
and U36855 (N_36855,N_32141,N_30270);
and U36856 (N_36856,N_31415,N_32320);
xor U36857 (N_36857,N_30791,N_34742);
xor U36858 (N_36858,N_31723,N_33005);
and U36859 (N_36859,N_33465,N_34917);
and U36860 (N_36860,N_33232,N_30510);
or U36861 (N_36861,N_30227,N_34999);
nand U36862 (N_36862,N_34704,N_33765);
nor U36863 (N_36863,N_32615,N_30811);
xor U36864 (N_36864,N_33705,N_33259);
and U36865 (N_36865,N_30536,N_32224);
or U36866 (N_36866,N_34782,N_30593);
or U36867 (N_36867,N_34085,N_32873);
xnor U36868 (N_36868,N_32707,N_33925);
nor U36869 (N_36869,N_32481,N_33991);
or U36870 (N_36870,N_30832,N_30554);
nand U36871 (N_36871,N_30812,N_33155);
nand U36872 (N_36872,N_34996,N_30118);
or U36873 (N_36873,N_31599,N_33639);
and U36874 (N_36874,N_32429,N_34629);
nand U36875 (N_36875,N_32559,N_30436);
xor U36876 (N_36876,N_31501,N_33052);
xnor U36877 (N_36877,N_30285,N_32772);
nor U36878 (N_36878,N_31583,N_32538);
nand U36879 (N_36879,N_31701,N_33792);
or U36880 (N_36880,N_33969,N_33446);
xor U36881 (N_36881,N_31497,N_33270);
nand U36882 (N_36882,N_32330,N_33878);
nor U36883 (N_36883,N_33709,N_34927);
nand U36884 (N_36884,N_31255,N_32659);
and U36885 (N_36885,N_33608,N_31239);
nand U36886 (N_36886,N_31828,N_30896);
or U36887 (N_36887,N_33228,N_31302);
and U36888 (N_36888,N_30457,N_31982);
and U36889 (N_36889,N_33588,N_31270);
xnor U36890 (N_36890,N_34123,N_34912);
xnor U36891 (N_36891,N_32136,N_31648);
nor U36892 (N_36892,N_33945,N_30739);
and U36893 (N_36893,N_30777,N_32435);
nand U36894 (N_36894,N_32316,N_30416);
nand U36895 (N_36895,N_32703,N_34703);
xnor U36896 (N_36896,N_33730,N_32413);
and U36897 (N_36897,N_30117,N_33230);
nand U36898 (N_36898,N_30588,N_30610);
nand U36899 (N_36899,N_34931,N_34112);
or U36900 (N_36900,N_32700,N_34552);
nand U36901 (N_36901,N_32882,N_31026);
or U36902 (N_36902,N_30392,N_31799);
nand U36903 (N_36903,N_32454,N_32730);
nor U36904 (N_36904,N_32631,N_34920);
and U36905 (N_36905,N_30069,N_30417);
xor U36906 (N_36906,N_33745,N_31065);
or U36907 (N_36907,N_30494,N_34779);
nor U36908 (N_36908,N_31481,N_32763);
nor U36909 (N_36909,N_34644,N_34332);
nand U36910 (N_36910,N_33119,N_31952);
or U36911 (N_36911,N_30648,N_30965);
nor U36912 (N_36912,N_32635,N_30054);
and U36913 (N_36913,N_31018,N_33203);
nand U36914 (N_36914,N_32742,N_31758);
nand U36915 (N_36915,N_32896,N_33914);
nand U36916 (N_36916,N_31476,N_33352);
nand U36917 (N_36917,N_33704,N_34149);
or U36918 (N_36918,N_34176,N_31071);
and U36919 (N_36919,N_33852,N_32872);
or U36920 (N_36920,N_33664,N_31832);
nand U36921 (N_36921,N_32750,N_34815);
nor U36922 (N_36922,N_34849,N_30402);
and U36923 (N_36923,N_30706,N_33930);
nand U36924 (N_36924,N_34934,N_31777);
or U36925 (N_36925,N_34119,N_30275);
xor U36926 (N_36926,N_34650,N_33531);
nor U36927 (N_36927,N_30548,N_33235);
and U36928 (N_36928,N_32364,N_33046);
or U36929 (N_36929,N_33988,N_34418);
and U36930 (N_36930,N_30134,N_32450);
nor U36931 (N_36931,N_30099,N_32352);
nand U36932 (N_36932,N_32781,N_30910);
and U36933 (N_36933,N_34660,N_33607);
and U36934 (N_36934,N_31007,N_30165);
and U36935 (N_36935,N_30306,N_30433);
xor U36936 (N_36936,N_34254,N_32247);
and U36937 (N_36937,N_34953,N_32110);
xnor U36938 (N_36938,N_34701,N_32124);
or U36939 (N_36939,N_31613,N_32958);
nand U36940 (N_36940,N_31842,N_30749);
nand U36941 (N_36941,N_34311,N_34419);
and U36942 (N_36942,N_33550,N_31025);
nor U36943 (N_36943,N_31362,N_33702);
or U36944 (N_36944,N_32285,N_31257);
nand U36945 (N_36945,N_32396,N_30430);
nor U36946 (N_36946,N_33882,N_32580);
nand U36947 (N_36947,N_30180,N_30760);
or U36948 (N_36948,N_30246,N_34762);
xnor U36949 (N_36949,N_31231,N_32003);
and U36950 (N_36950,N_30931,N_33782);
xnor U36951 (N_36951,N_34351,N_32047);
or U36952 (N_36952,N_32191,N_33632);
nand U36953 (N_36953,N_34449,N_30999);
xor U36954 (N_36954,N_31653,N_32685);
nor U36955 (N_36955,N_31896,N_31895);
and U36956 (N_36956,N_34251,N_32398);
nor U36957 (N_36957,N_33174,N_32744);
xor U36958 (N_36958,N_30168,N_33204);
nand U36959 (N_36959,N_34437,N_31946);
or U36960 (N_36960,N_31224,N_33226);
nand U36961 (N_36961,N_30063,N_31280);
or U36962 (N_36962,N_31691,N_32214);
or U36963 (N_36963,N_34118,N_31865);
or U36964 (N_36964,N_33450,N_32265);
nand U36965 (N_36965,N_31311,N_34321);
and U36966 (N_36966,N_31742,N_30277);
or U36967 (N_36967,N_32656,N_32333);
nand U36968 (N_36968,N_30712,N_33816);
nand U36969 (N_36969,N_32241,N_32353);
and U36970 (N_36970,N_31718,N_30174);
or U36971 (N_36971,N_32091,N_34575);
and U36972 (N_36972,N_34787,N_32501);
nand U36973 (N_36973,N_31266,N_32919);
xnor U36974 (N_36974,N_31284,N_33283);
nand U36975 (N_36975,N_33872,N_34467);
nand U36976 (N_36976,N_30601,N_32665);
and U36977 (N_36977,N_32673,N_34869);
or U36978 (N_36978,N_31074,N_31365);
xnor U36979 (N_36979,N_34324,N_31423);
xor U36980 (N_36980,N_34224,N_33502);
nand U36981 (N_36981,N_32630,N_34657);
nand U36982 (N_36982,N_34866,N_32117);
nand U36983 (N_36983,N_30624,N_34636);
or U36984 (N_36984,N_32957,N_32221);
and U36985 (N_36985,N_34268,N_31178);
xnor U36986 (N_36986,N_33084,N_32863);
nor U36987 (N_36987,N_32210,N_30878);
xor U36988 (N_36988,N_30523,N_31034);
nor U36989 (N_36989,N_33798,N_34592);
xnor U36990 (N_36990,N_33853,N_30472);
nor U36991 (N_36991,N_30028,N_30483);
and U36992 (N_36992,N_33908,N_30143);
or U36993 (N_36993,N_34832,N_31054);
nand U36994 (N_36994,N_30710,N_33540);
nand U36995 (N_36995,N_30369,N_31327);
xor U36996 (N_36996,N_31949,N_34173);
and U36997 (N_36997,N_30971,N_30524);
or U36998 (N_36998,N_32422,N_32570);
nor U36999 (N_36999,N_34440,N_30766);
nor U37000 (N_37000,N_33901,N_31531);
nand U37001 (N_37001,N_34643,N_34110);
nor U37002 (N_37002,N_31596,N_33139);
and U37003 (N_37003,N_33508,N_30917);
and U37004 (N_37004,N_32705,N_34597);
xnor U37005 (N_37005,N_34414,N_33438);
and U37006 (N_37006,N_30318,N_34635);
nand U37007 (N_37007,N_31689,N_30120);
and U37008 (N_37008,N_31373,N_33370);
xnor U37009 (N_37009,N_34794,N_33776);
or U37010 (N_37010,N_30849,N_30271);
xor U37011 (N_37011,N_34315,N_33667);
or U37012 (N_37012,N_30629,N_34836);
or U37013 (N_37013,N_34905,N_34816);
and U37014 (N_37014,N_34221,N_34576);
nor U37015 (N_37015,N_31051,N_31803);
xnor U37016 (N_37016,N_32994,N_34810);
nand U37017 (N_37017,N_33100,N_33785);
nor U37018 (N_37018,N_33743,N_32150);
nor U37019 (N_37019,N_34536,N_30839);
or U37020 (N_37020,N_32534,N_32151);
or U37021 (N_37021,N_32467,N_33170);
nand U37022 (N_37022,N_30762,N_33708);
nand U37023 (N_37023,N_32064,N_30622);
nand U37024 (N_37024,N_32451,N_32355);
nand U37025 (N_37025,N_30014,N_34065);
xnor U37026 (N_37026,N_33295,N_33433);
and U37027 (N_37027,N_31140,N_33390);
or U37028 (N_37028,N_31600,N_33019);
or U37029 (N_37029,N_30748,N_32036);
or U37030 (N_37030,N_31882,N_34230);
nand U37031 (N_37031,N_33666,N_34163);
nor U37032 (N_37032,N_34113,N_32229);
or U37033 (N_37033,N_32235,N_31064);
xnor U37034 (N_37034,N_32732,N_31532);
or U37035 (N_37035,N_33069,N_31639);
and U37036 (N_37036,N_34171,N_33712);
or U37037 (N_37037,N_32099,N_31857);
xor U37038 (N_37038,N_31673,N_33905);
nor U37039 (N_37039,N_32066,N_33242);
or U37040 (N_37040,N_34248,N_32740);
xor U37041 (N_37041,N_34697,N_32558);
and U37042 (N_37042,N_34801,N_31435);
and U37043 (N_37043,N_34633,N_30047);
nand U37044 (N_37044,N_31482,N_33626);
nand U37045 (N_37045,N_30532,N_34478);
and U37046 (N_37046,N_31369,N_33334);
nor U37047 (N_37047,N_34910,N_33977);
and U37048 (N_37048,N_31247,N_32931);
or U37049 (N_37049,N_34331,N_34711);
or U37050 (N_37050,N_32989,N_30757);
and U37051 (N_37051,N_33106,N_30974);
xor U37052 (N_37052,N_33825,N_33913);
xor U37053 (N_37053,N_32009,N_33032);
xnor U37054 (N_37054,N_33064,N_32779);
nand U37055 (N_37055,N_31619,N_32761);
nand U37056 (N_37056,N_34995,N_33034);
xor U37057 (N_37057,N_34111,N_30732);
xnor U37058 (N_37058,N_33591,N_34854);
and U37059 (N_37059,N_30596,N_32686);
nand U37060 (N_37060,N_31504,N_30282);
nand U37061 (N_37061,N_33749,N_32176);
or U37062 (N_37062,N_34260,N_32525);
and U37063 (N_37063,N_33731,N_33697);
or U37064 (N_37064,N_31747,N_30782);
nand U37065 (N_37065,N_34639,N_33654);
or U37066 (N_37066,N_31053,N_32069);
nand U37067 (N_37067,N_31970,N_31680);
or U37068 (N_37068,N_33518,N_34582);
and U37069 (N_37069,N_32533,N_30181);
nor U37070 (N_37070,N_34740,N_31769);
nor U37071 (N_37071,N_31141,N_30966);
and U37072 (N_37072,N_30879,N_30867);
xnor U37073 (N_37073,N_34239,N_32395);
nand U37074 (N_37074,N_33884,N_31350);
nor U37075 (N_37075,N_31490,N_31128);
or U37076 (N_37076,N_31884,N_33382);
nand U37077 (N_37077,N_34401,N_33451);
nand U37078 (N_37078,N_31620,N_31813);
nand U37079 (N_37079,N_31515,N_30279);
xnor U37080 (N_37080,N_34355,N_34002);
nand U37081 (N_37081,N_30387,N_32734);
nor U37082 (N_37082,N_33694,N_32548);
and U37083 (N_37083,N_31346,N_32916);
xnor U37084 (N_37084,N_32647,N_33610);
nor U37085 (N_37085,N_34929,N_31077);
xor U37086 (N_37086,N_30157,N_33854);
nor U37087 (N_37087,N_30633,N_33698);
xnor U37088 (N_37088,N_32981,N_32680);
and U37089 (N_37089,N_33758,N_34264);
or U37090 (N_37090,N_34197,N_32881);
or U37091 (N_37091,N_31092,N_31854);
and U37092 (N_37092,N_34309,N_32106);
nand U37093 (N_37093,N_33799,N_32160);
nand U37094 (N_37094,N_32679,N_33436);
nand U37095 (N_37095,N_31567,N_33771);
nand U37096 (N_37096,N_32428,N_34568);
or U37097 (N_37097,N_32016,N_32213);
or U37098 (N_37098,N_32489,N_31456);
and U37099 (N_37099,N_31574,N_32425);
xor U37100 (N_37100,N_30375,N_34253);
or U37101 (N_37101,N_31555,N_33305);
and U37102 (N_37102,N_31046,N_30486);
nor U37103 (N_37103,N_33290,N_33151);
xor U37104 (N_37104,N_34017,N_31726);
and U37105 (N_37105,N_34214,N_34606);
nand U37106 (N_37106,N_31568,N_30415);
xnor U37107 (N_37107,N_31205,N_34222);
or U37108 (N_37108,N_31468,N_30145);
nand U37109 (N_37109,N_33214,N_34018);
nor U37110 (N_37110,N_31227,N_31840);
nand U37111 (N_37111,N_34885,N_34896);
nand U37112 (N_37112,N_31732,N_32663);
and U37113 (N_37113,N_30219,N_30269);
nand U37114 (N_37114,N_32704,N_34347);
and U37115 (N_37115,N_33754,N_30684);
and U37116 (N_37116,N_31163,N_30580);
and U37117 (N_37117,N_31677,N_30537);
nand U37118 (N_37118,N_34627,N_33570);
nand U37119 (N_37119,N_30798,N_31617);
nand U37120 (N_37120,N_34673,N_30013);
or U37121 (N_37121,N_33416,N_33790);
xnor U37122 (N_37122,N_30763,N_33128);
nor U37123 (N_37123,N_30534,N_31646);
xor U37124 (N_37124,N_31491,N_30994);
xor U37125 (N_37125,N_31602,N_30123);
or U37126 (N_37126,N_34871,N_31218);
and U37127 (N_37127,N_34339,N_32900);
nand U37128 (N_37128,N_33445,N_31746);
or U37129 (N_37129,N_31557,N_33240);
xor U37130 (N_37130,N_30689,N_34177);
and U37131 (N_37131,N_30765,N_32835);
and U37132 (N_37132,N_34049,N_31669);
xnor U37133 (N_37133,N_32828,N_34658);
or U37134 (N_37134,N_34067,N_31945);
or U37135 (N_37135,N_33718,N_33947);
nand U37136 (N_37136,N_31154,N_34714);
xnor U37137 (N_37137,N_33068,N_30122);
xor U37138 (N_37138,N_31418,N_31738);
xor U37139 (N_37139,N_32693,N_34562);
nand U37140 (N_37140,N_33575,N_32553);
nor U37141 (N_37141,N_30960,N_32271);
or U37142 (N_37142,N_31715,N_32318);
nand U37143 (N_37143,N_32754,N_31372);
nand U37144 (N_37144,N_33867,N_30656);
xor U37145 (N_37145,N_31118,N_33829);
nor U37146 (N_37146,N_34051,N_32488);
xnor U37147 (N_37147,N_33197,N_33268);
nor U37148 (N_37148,N_32356,N_32557);
nand U37149 (N_37149,N_33169,N_33611);
nor U37150 (N_37150,N_34405,N_31931);
or U37151 (N_37151,N_31349,N_31508);
nand U37152 (N_37152,N_34044,N_30114);
xnor U37153 (N_37153,N_30137,N_33489);
nor U37154 (N_37154,N_30595,N_32103);
xnor U37155 (N_37155,N_30701,N_31404);
xor U37156 (N_37156,N_33734,N_34983);
xor U37157 (N_37157,N_34292,N_33037);
and U37158 (N_37158,N_30223,N_34835);
nor U37159 (N_37159,N_31524,N_30608);
nor U37160 (N_37160,N_30874,N_31493);
xor U37161 (N_37161,N_32441,N_34587);
nor U37162 (N_37162,N_31806,N_30853);
xnor U37163 (N_37163,N_34872,N_34364);
nand U37164 (N_37164,N_33824,N_32646);
nand U37165 (N_37165,N_31696,N_30649);
or U37166 (N_37166,N_34145,N_34795);
nor U37167 (N_37167,N_31509,N_33768);
or U37168 (N_37168,N_34760,N_31488);
nand U37169 (N_37169,N_30625,N_31058);
nand U37170 (N_37170,N_34227,N_31472);
or U37171 (N_37171,N_32181,N_30021);
or U37172 (N_37172,N_31494,N_30943);
xor U37173 (N_37173,N_30089,N_30353);
xnor U37174 (N_37174,N_32133,N_30476);
nand U37175 (N_37175,N_34477,N_30735);
or U37176 (N_37176,N_34427,N_30558);
nand U37177 (N_37177,N_31438,N_31851);
or U37178 (N_37178,N_30549,N_31027);
and U37179 (N_37179,N_32842,N_34093);
and U37180 (N_37180,N_30671,N_30347);
nor U37181 (N_37181,N_31214,N_33781);
nand U37182 (N_37182,N_33889,N_30542);
xnor U37183 (N_37183,N_31235,N_32609);
xor U37184 (N_37184,N_34053,N_32902);
nor U37185 (N_37185,N_32286,N_33292);
or U37186 (N_37186,N_31755,N_30178);
or U37187 (N_37187,N_34668,N_30933);
or U37188 (N_37188,N_33903,N_30561);
and U37189 (N_37189,N_33093,N_30169);
and U37190 (N_37190,N_30038,N_34061);
and U37191 (N_37191,N_33057,N_31127);
or U37192 (N_37192,N_32256,N_34333);
nor U37193 (N_37193,N_32520,N_32102);
nand U37194 (N_37194,N_34665,N_32677);
nand U37195 (N_37195,N_30265,N_30460);
xor U37196 (N_37196,N_31000,N_34493);
and U37197 (N_37197,N_32759,N_30767);
and U37198 (N_37198,N_32043,N_30424);
or U37199 (N_37199,N_32818,N_33058);
and U37200 (N_37200,N_31171,N_34255);
or U37201 (N_37201,N_34626,N_32849);
nor U37202 (N_37202,N_33388,N_32120);
nor U37203 (N_37203,N_31165,N_31315);
nand U37204 (N_37204,N_31150,N_33208);
xnor U37205 (N_37205,N_32165,N_31189);
and U37206 (N_37206,N_31319,N_31705);
xnor U37207 (N_37207,N_34174,N_30578);
or U37208 (N_37208,N_34753,N_32075);
nor U37209 (N_37209,N_32477,N_30362);
and U37210 (N_37210,N_32226,N_34613);
or U37211 (N_37211,N_32449,N_32943);
xor U37212 (N_37212,N_34157,N_31883);
nand U37213 (N_37213,N_33163,N_34137);
nor U37214 (N_37214,N_31553,N_32751);
nor U37215 (N_37215,N_33954,N_32691);
nand U37216 (N_37216,N_31293,N_33638);
xnor U37217 (N_37217,N_30921,N_31986);
xor U37218 (N_37218,N_33302,N_30212);
xnor U37219 (N_37219,N_33440,N_33952);
and U37220 (N_37220,N_33150,N_33239);
or U37221 (N_37221,N_33953,N_30502);
or U37222 (N_37222,N_31584,N_33691);
or U37223 (N_37223,N_32174,N_31906);
xnor U37224 (N_37224,N_30698,N_30583);
xnor U37225 (N_37225,N_34652,N_34249);
nor U37226 (N_37226,N_30643,N_33251);
nand U37227 (N_37227,N_34037,N_32480);
and U37228 (N_37228,N_33383,N_34806);
or U37229 (N_37229,N_31240,N_32018);
xor U37230 (N_37230,N_30793,N_30920);
and U37231 (N_37231,N_30245,N_33721);
or U37232 (N_37232,N_30052,N_31174);
nand U37233 (N_37233,N_33562,N_34159);
xnor U37234 (N_37234,N_32613,N_30514);
nor U37235 (N_37235,N_32524,N_30001);
or U37236 (N_37236,N_32122,N_31384);
or U37237 (N_37237,N_31301,N_30645);
and U37238 (N_37238,N_31507,N_31262);
xnor U37239 (N_37239,N_32743,N_32051);
or U37240 (N_37240,N_31164,N_32180);
and U37241 (N_37241,N_30007,N_32368);
or U37242 (N_37242,N_31442,N_32457);
or U37243 (N_37243,N_30568,N_31961);
and U37244 (N_37244,N_30451,N_34294);
and U37245 (N_37245,N_30915,N_30641);
or U37246 (N_37246,N_34683,N_32572);
or U37247 (N_37247,N_30205,N_31216);
and U37248 (N_37248,N_33039,N_33076);
or U37249 (N_37249,N_30287,N_31876);
xor U37250 (N_37250,N_31919,N_31161);
nand U37251 (N_37251,N_31500,N_33796);
nor U37252 (N_37252,N_33073,N_34874);
xnor U37253 (N_37253,N_32278,N_31321);
nor U37254 (N_37254,N_34744,N_30997);
xor U37255 (N_37255,N_32476,N_30303);
or U37256 (N_37256,N_31122,N_31962);
nor U37257 (N_37257,N_32625,N_30040);
nor U37258 (N_37258,N_33874,N_30598);
nand U37259 (N_37259,N_31185,N_31716);
nand U37260 (N_37260,N_30885,N_31675);
nand U37261 (N_37261,N_33458,N_32777);
or U37262 (N_37262,N_31393,N_33189);
nor U37263 (N_37263,N_33689,N_33594);
nor U37264 (N_37264,N_34313,N_33755);
or U37265 (N_37265,N_33946,N_33757);
or U37266 (N_37266,N_33993,N_33476);
xnor U37267 (N_37267,N_34843,N_30912);
and U37268 (N_37268,N_31437,N_32727);
xor U37269 (N_37269,N_32055,N_33517);
and U37270 (N_37270,N_31885,N_34079);
and U37271 (N_37271,N_33199,N_32883);
nand U37272 (N_37272,N_31960,N_30563);
xnor U37273 (N_37273,N_31745,N_33975);
and U37274 (N_37274,N_33602,N_34016);
nand U37275 (N_37275,N_32382,N_30106);
nand U37276 (N_37276,N_32272,N_33807);
xor U37277 (N_37277,N_32230,N_33149);
nand U37278 (N_37278,N_30987,N_33652);
and U37279 (N_37279,N_34143,N_31211);
nor U37280 (N_37280,N_32531,N_32302);
xor U37281 (N_37281,N_34774,N_31609);
and U37282 (N_37282,N_30254,N_34245);
and U37283 (N_37283,N_32469,N_34487);
or U37284 (N_37284,N_33468,N_32788);
or U37285 (N_37285,N_33212,N_33642);
or U37286 (N_37286,N_34187,N_30905);
and U37287 (N_37287,N_32736,N_30397);
or U37288 (N_37288,N_32640,N_34194);
xnor U37289 (N_37289,N_34499,N_34833);
nor U37290 (N_37290,N_32079,N_34269);
or U37291 (N_37291,N_32054,N_30844);
or U37292 (N_37292,N_32787,N_34608);
or U37293 (N_37293,N_31938,N_30814);
and U37294 (N_37294,N_32668,N_30043);
nor U37295 (N_37295,N_32212,N_33612);
xnor U37296 (N_37296,N_34096,N_32551);
or U37297 (N_37297,N_33659,N_31023);
nor U37298 (N_37298,N_31954,N_30565);
nand U37299 (N_37299,N_33113,N_31935);
xnor U37300 (N_37300,N_32955,N_30754);
or U37301 (N_37301,N_33092,N_32774);
nand U37302 (N_37302,N_31666,N_32227);
and U37303 (N_37303,N_34964,N_30239);
or U37304 (N_37304,N_33692,N_30626);
or U37305 (N_37305,N_33592,N_30961);
or U37306 (N_37306,N_33345,N_33880);
nand U37307 (N_37307,N_30381,N_34671);
and U37308 (N_37308,N_34327,N_31530);
xor U37309 (N_37309,N_33194,N_34461);
or U37310 (N_37310,N_32815,N_34911);
nand U37311 (N_37311,N_30873,N_34213);
nor U37312 (N_37312,N_33299,N_30519);
nand U37313 (N_37313,N_34698,N_30066);
nor U37314 (N_37314,N_33679,N_33358);
and U37315 (N_37315,N_33928,N_33260);
nor U37316 (N_37316,N_34619,N_32182);
or U37317 (N_37317,N_33328,N_32891);
or U37318 (N_37318,N_34618,N_31889);
or U37319 (N_37319,N_30538,N_32726);
and U37320 (N_37320,N_33778,N_33108);
nand U37321 (N_37321,N_34752,N_33998);
nor U37322 (N_37322,N_32795,N_34480);
nand U37323 (N_37323,N_34090,N_31193);
or U37324 (N_37324,N_30819,N_31207);
nor U37325 (N_37325,N_34190,N_33215);
nor U37326 (N_37326,N_31674,N_30675);
or U37327 (N_37327,N_32611,N_34502);
xnor U37328 (N_37328,N_34218,N_31433);
and U37329 (N_37329,N_34530,N_33670);
nor U37330 (N_37330,N_32826,N_33090);
or U37331 (N_37331,N_34631,N_30551);
nand U37332 (N_37332,N_30898,N_32549);
nor U37333 (N_37333,N_34936,N_32292);
or U37334 (N_37334,N_34244,N_33662);
or U37335 (N_37335,N_30495,N_30391);
nand U37336 (N_37336,N_33740,N_30017);
or U37337 (N_37337,N_34649,N_30597);
or U37338 (N_37338,N_32065,N_34354);
nor U37339 (N_37339,N_30356,N_31587);
nor U37340 (N_37340,N_34829,N_34949);
and U37341 (N_37341,N_31624,N_31412);
nor U37342 (N_37342,N_33110,N_34186);
or U37343 (N_37343,N_32947,N_31844);
xnor U37344 (N_37344,N_34518,N_33356);
nor U37345 (N_37345,N_32735,N_33999);
nor U37346 (N_37346,N_33265,N_33580);
xor U37347 (N_37347,N_30566,N_34397);
xnor U37348 (N_37348,N_33176,N_32252);
nand U37349 (N_37349,N_32264,N_33911);
nor U37350 (N_37350,N_34743,N_33031);
or U37351 (N_37351,N_32257,N_33396);
nor U37352 (N_37352,N_32266,N_34708);
nand U37353 (N_37353,N_33428,N_31421);
nand U37354 (N_37354,N_33105,N_33979);
xor U37355 (N_37355,N_32923,N_34103);
and U37356 (N_37356,N_31096,N_34550);
xnor U37357 (N_37357,N_32648,N_32514);
xor U37358 (N_37358,N_30358,N_30253);
and U37359 (N_37359,N_31774,N_32473);
or U37360 (N_37360,N_30929,N_34513);
nor U37361 (N_37361,N_30161,N_30775);
nand U37362 (N_37362,N_31478,N_34507);
or U37363 (N_37363,N_30591,N_31475);
and U37364 (N_37364,N_30230,N_34124);
or U37365 (N_37365,N_32339,N_32582);
xor U37366 (N_37366,N_30034,N_33338);
or U37367 (N_37367,N_30341,N_31534);
nand U37368 (N_37368,N_30888,N_34799);
or U37369 (N_37369,N_34380,N_33319);
nand U37370 (N_37370,N_31300,N_31573);
or U37371 (N_37371,N_34219,N_32309);
nor U37372 (N_37372,N_31905,N_32846);
or U37373 (N_37373,N_32447,N_33504);
or U37374 (N_37374,N_31159,N_34726);
nand U37375 (N_37375,N_34894,N_34560);
nand U37376 (N_37376,N_32206,N_34457);
xor U37377 (N_37377,N_31019,N_33621);
nand U37378 (N_37378,N_31996,N_30370);
nand U37379 (N_37379,N_33185,N_31013);
xor U37380 (N_37380,N_30420,N_34577);
xnor U37381 (N_37381,N_32840,N_33399);
or U37382 (N_37382,N_31651,N_31351);
nand U37383 (N_37383,N_31462,N_33430);
nor U37384 (N_37384,N_30323,N_32962);
nand U37385 (N_37385,N_32154,N_32255);
nand U37386 (N_37386,N_31834,N_32283);
nand U37387 (N_37387,N_33028,N_30508);
xor U37388 (N_37388,N_30197,N_33936);
or U37389 (N_37389,N_31080,N_30384);
xnor U37390 (N_37390,N_32017,N_31124);
and U37391 (N_37391,N_31089,N_32683);
nor U37392 (N_37392,N_31175,N_31139);
nand U37393 (N_37393,N_33855,N_33313);
and U37394 (N_37394,N_30499,N_34175);
and U37395 (N_37395,N_32579,N_30564);
nor U37396 (N_37396,N_33312,N_31916);
nand U37397 (N_37397,N_31809,N_30851);
and U37398 (N_37398,N_30198,N_32723);
nand U37399 (N_37399,N_33624,N_30071);
nor U37400 (N_37400,N_32108,N_33599);
and U37401 (N_37401,N_30432,N_32290);
xnor U37402 (N_37402,N_33263,N_31394);
nand U37403 (N_37403,N_34041,N_31220);
xnor U37404 (N_37404,N_31956,N_32905);
or U37405 (N_37405,N_34733,N_33921);
xor U37406 (N_37406,N_30064,N_30126);
and U37407 (N_37407,N_31233,N_34094);
or U37408 (N_37408,N_31084,N_34413);
and U37409 (N_37409,N_30781,N_31250);
nor U37410 (N_37410,N_33541,N_32448);
or U37411 (N_37411,N_30913,N_34387);
nor U37412 (N_37412,N_33939,N_31269);
nor U37413 (N_37413,N_30394,N_33363);
or U37414 (N_37414,N_33158,N_32569);
or U37415 (N_37415,N_31014,N_32262);
nand U37416 (N_37416,N_33700,N_30903);
and U37417 (N_37417,N_34679,N_34713);
xor U37418 (N_37418,N_34282,N_30941);
nor U37419 (N_37419,N_30112,N_31252);
and U37420 (N_37420,N_31199,N_30945);
xor U37421 (N_37421,N_30745,N_30291);
or U37422 (N_37422,N_30005,N_32731);
nand U37423 (N_37423,N_30792,N_31303);
and U37424 (N_37424,N_30779,N_33401);
or U37425 (N_37425,N_33761,N_33794);
or U37426 (N_37426,N_34257,N_34616);
xor U37427 (N_37427,N_31569,N_31366);
nand U37428 (N_37428,N_34968,N_30470);
or U37429 (N_37429,N_30340,N_33286);
nor U37430 (N_37430,N_34212,N_33395);
nor U37431 (N_37431,N_31168,N_33102);
nand U37432 (N_37432,N_34058,N_31859);
or U37433 (N_37433,N_30975,N_33205);
or U37434 (N_37434,N_31110,N_33072);
nand U37435 (N_37435,N_34297,N_34278);
and U37436 (N_37436,N_34142,N_33587);
xor U37437 (N_37437,N_32070,N_31304);
xnor U37438 (N_37438,N_31138,N_34396);
nor U37439 (N_37439,N_33252,N_34078);
xnor U37440 (N_37440,N_30475,N_31197);
nand U37441 (N_37441,N_34108,N_30435);
and U37442 (N_37442,N_32135,N_33414);
xnor U37443 (N_37443,N_34232,N_34392);
and U37444 (N_37444,N_33631,N_34101);
and U37445 (N_37445,N_33217,N_33024);
or U37446 (N_37446,N_34540,N_33948);
or U37447 (N_37447,N_31169,N_33480);
xnor U37448 (N_37448,N_31924,N_33017);
nand U37449 (N_37449,N_34481,N_31551);
nand U37450 (N_37450,N_31083,N_31727);
or U37451 (N_37451,N_31145,N_30434);
nor U37452 (N_37452,N_33135,N_32033);
or U37453 (N_37453,N_30095,N_34945);
nor U37454 (N_37454,N_32575,N_30520);
nand U37455 (N_37455,N_34557,N_34395);
or U37456 (N_37456,N_31446,N_30509);
and U37457 (N_37457,N_34020,N_33348);
xor U37458 (N_37458,N_31533,N_34398);
nand U37459 (N_37459,N_31391,N_32172);
and U37460 (N_37460,N_32403,N_31447);
or U37461 (N_37461,N_30527,N_34655);
and U37462 (N_37462,N_33527,N_34032);
nand U37463 (N_37463,N_32602,N_33142);
nor U37464 (N_37464,N_30077,N_31839);
or U37465 (N_37465,N_31055,N_34972);
and U37466 (N_37466,N_30320,N_30366);
and U37467 (N_37467,N_32565,N_32348);
or U37468 (N_37468,N_32158,N_31717);
nand U37469 (N_37469,N_34454,N_30314);
xnor U37470 (N_37470,N_32006,N_33916);
or U37471 (N_37471,N_31294,N_32078);
nor U37472 (N_37472,N_32184,N_34011);
or U37473 (N_37473,N_30289,N_30504);
xor U37474 (N_37474,N_32020,N_31328);
nor U37475 (N_37475,N_32618,N_32109);
and U37476 (N_37476,N_32713,N_34994);
nand U37477 (N_37477,N_32970,N_34312);
nand U37478 (N_37478,N_34486,N_34050);
and U37479 (N_37479,N_32825,N_31861);
nor U37480 (N_37480,N_32987,N_31912);
and U37481 (N_37481,N_30150,N_30628);
xnor U37482 (N_37482,N_34741,N_30914);
or U37483 (N_37483,N_30373,N_34890);
xor U37484 (N_37484,N_32632,N_30871);
and U37485 (N_37485,N_30081,N_30138);
nor U37486 (N_37486,N_32621,N_34205);
and U37487 (N_37487,N_30962,N_32342);
and U37488 (N_37488,N_32964,N_34990);
or U37489 (N_37489,N_34115,N_33159);
xor U37490 (N_37490,N_34976,N_30543);
nor U37491 (N_37491,N_33400,N_31963);
nor U37492 (N_37492,N_33055,N_31102);
nand U37493 (N_37493,N_32053,N_34838);
nand U37494 (N_37494,N_34261,N_30097);
nand U37495 (N_37495,N_32295,N_31757);
xor U37496 (N_37496,N_34583,N_32573);
nand U37497 (N_37497,N_30404,N_33512);
nor U37498 (N_37498,N_31181,N_33820);
xnor U37499 (N_37499,N_33582,N_31457);
or U37500 (N_37500,N_32363,N_32292);
nand U37501 (N_37501,N_33597,N_34807);
nor U37502 (N_37502,N_33177,N_33388);
nor U37503 (N_37503,N_32145,N_34006);
nand U37504 (N_37504,N_33409,N_33151);
or U37505 (N_37505,N_30863,N_33680);
nand U37506 (N_37506,N_34192,N_34784);
or U37507 (N_37507,N_31835,N_31441);
or U37508 (N_37508,N_31043,N_30826);
xor U37509 (N_37509,N_30558,N_31831);
nand U37510 (N_37510,N_33187,N_30767);
nor U37511 (N_37511,N_33464,N_30518);
nand U37512 (N_37512,N_30330,N_32436);
nand U37513 (N_37513,N_31397,N_33393);
xnor U37514 (N_37514,N_34476,N_31103);
nor U37515 (N_37515,N_30143,N_31159);
or U37516 (N_37516,N_32284,N_30804);
or U37517 (N_37517,N_33414,N_33832);
nor U37518 (N_37518,N_33388,N_30405);
or U37519 (N_37519,N_32788,N_34745);
nand U37520 (N_37520,N_34544,N_30279);
xor U37521 (N_37521,N_31893,N_34952);
nand U37522 (N_37522,N_31652,N_33629);
nor U37523 (N_37523,N_33942,N_30124);
nor U37524 (N_37524,N_34927,N_31706);
nor U37525 (N_37525,N_32729,N_31860);
nor U37526 (N_37526,N_33450,N_31649);
nand U37527 (N_37527,N_34708,N_31207);
nor U37528 (N_37528,N_34621,N_31696);
and U37529 (N_37529,N_34864,N_33519);
or U37530 (N_37530,N_34767,N_32167);
nor U37531 (N_37531,N_30178,N_30474);
nand U37532 (N_37532,N_31626,N_30308);
and U37533 (N_37533,N_34300,N_32723);
or U37534 (N_37534,N_33877,N_33833);
nand U37535 (N_37535,N_30607,N_31245);
xor U37536 (N_37536,N_30374,N_31711);
nand U37537 (N_37537,N_33719,N_33362);
and U37538 (N_37538,N_30969,N_32099);
or U37539 (N_37539,N_31785,N_32037);
and U37540 (N_37540,N_33618,N_30363);
or U37541 (N_37541,N_32273,N_33937);
nor U37542 (N_37542,N_31263,N_32335);
nand U37543 (N_37543,N_31047,N_32868);
nand U37544 (N_37544,N_32590,N_31306);
xor U37545 (N_37545,N_33678,N_30618);
or U37546 (N_37546,N_34243,N_33950);
or U37547 (N_37547,N_34072,N_31653);
nand U37548 (N_37548,N_31042,N_32703);
xor U37549 (N_37549,N_32742,N_31842);
or U37550 (N_37550,N_31759,N_31673);
nor U37551 (N_37551,N_34768,N_32083);
nor U37552 (N_37552,N_32719,N_32961);
or U37553 (N_37553,N_33775,N_31552);
nor U37554 (N_37554,N_30325,N_32715);
nand U37555 (N_37555,N_31171,N_32848);
xnor U37556 (N_37556,N_34537,N_31043);
xnor U37557 (N_37557,N_33748,N_33394);
xnor U37558 (N_37558,N_30975,N_32702);
or U37559 (N_37559,N_30859,N_32290);
and U37560 (N_37560,N_33325,N_32100);
or U37561 (N_37561,N_30847,N_31760);
or U37562 (N_37562,N_30226,N_34162);
xnor U37563 (N_37563,N_30285,N_30815);
xnor U37564 (N_37564,N_32072,N_30649);
nor U37565 (N_37565,N_32352,N_33336);
nor U37566 (N_37566,N_31182,N_33802);
nand U37567 (N_37567,N_31631,N_31523);
nand U37568 (N_37568,N_33580,N_33366);
nor U37569 (N_37569,N_32575,N_31969);
nand U37570 (N_37570,N_33714,N_30459);
xor U37571 (N_37571,N_30330,N_30871);
nand U37572 (N_37572,N_33721,N_32439);
and U37573 (N_37573,N_34102,N_30358);
xnor U37574 (N_37574,N_33810,N_30012);
or U37575 (N_37575,N_32453,N_33764);
and U37576 (N_37576,N_30980,N_32307);
nor U37577 (N_37577,N_34721,N_34533);
or U37578 (N_37578,N_32201,N_30626);
nand U37579 (N_37579,N_31929,N_31175);
xor U37580 (N_37580,N_34638,N_30944);
xor U37581 (N_37581,N_33697,N_30542);
nand U37582 (N_37582,N_33788,N_31849);
or U37583 (N_37583,N_31111,N_33801);
xnor U37584 (N_37584,N_34575,N_31577);
and U37585 (N_37585,N_31713,N_32652);
and U37586 (N_37586,N_31721,N_31801);
nor U37587 (N_37587,N_30121,N_30096);
or U37588 (N_37588,N_33208,N_32882);
nand U37589 (N_37589,N_33313,N_30945);
or U37590 (N_37590,N_33127,N_33669);
nand U37591 (N_37591,N_30287,N_31937);
nand U37592 (N_37592,N_33805,N_33109);
nand U37593 (N_37593,N_34767,N_31570);
nand U37594 (N_37594,N_32459,N_33905);
nand U37595 (N_37595,N_30939,N_34235);
or U37596 (N_37596,N_31017,N_33300);
and U37597 (N_37597,N_30861,N_34935);
or U37598 (N_37598,N_31779,N_33324);
or U37599 (N_37599,N_34452,N_34811);
nor U37600 (N_37600,N_30504,N_31314);
nor U37601 (N_37601,N_33848,N_30218);
nor U37602 (N_37602,N_31554,N_31058);
nand U37603 (N_37603,N_30400,N_33303);
or U37604 (N_37604,N_32547,N_34446);
xor U37605 (N_37605,N_32058,N_34601);
and U37606 (N_37606,N_34980,N_31525);
xnor U37607 (N_37607,N_32410,N_33493);
nand U37608 (N_37608,N_33515,N_30138);
xnor U37609 (N_37609,N_30675,N_31466);
nor U37610 (N_37610,N_34061,N_32205);
or U37611 (N_37611,N_30364,N_34500);
and U37612 (N_37612,N_33591,N_30352);
or U37613 (N_37613,N_30680,N_30605);
and U37614 (N_37614,N_34610,N_30853);
nor U37615 (N_37615,N_33067,N_31193);
nor U37616 (N_37616,N_32792,N_30707);
nand U37617 (N_37617,N_34613,N_31364);
nand U37618 (N_37618,N_34438,N_32926);
nand U37619 (N_37619,N_30568,N_31183);
nand U37620 (N_37620,N_33796,N_32624);
or U37621 (N_37621,N_31013,N_31410);
nor U37622 (N_37622,N_33989,N_31710);
or U37623 (N_37623,N_31769,N_31937);
xnor U37624 (N_37624,N_32985,N_30788);
or U37625 (N_37625,N_33014,N_32580);
xor U37626 (N_37626,N_34639,N_30429);
xnor U37627 (N_37627,N_34282,N_31910);
or U37628 (N_37628,N_30997,N_31361);
or U37629 (N_37629,N_30734,N_30987);
or U37630 (N_37630,N_30226,N_30492);
xor U37631 (N_37631,N_32119,N_33652);
nor U37632 (N_37632,N_33920,N_30116);
xor U37633 (N_37633,N_30033,N_33416);
and U37634 (N_37634,N_31677,N_33503);
or U37635 (N_37635,N_31631,N_30546);
xnor U37636 (N_37636,N_34813,N_34307);
xnor U37637 (N_37637,N_30427,N_30754);
nand U37638 (N_37638,N_33124,N_33346);
and U37639 (N_37639,N_34769,N_31285);
nor U37640 (N_37640,N_30049,N_30683);
and U37641 (N_37641,N_31346,N_32765);
xor U37642 (N_37642,N_34941,N_34106);
or U37643 (N_37643,N_31525,N_33835);
and U37644 (N_37644,N_32180,N_30523);
and U37645 (N_37645,N_34567,N_31784);
or U37646 (N_37646,N_32292,N_31369);
nor U37647 (N_37647,N_32861,N_33129);
or U37648 (N_37648,N_33060,N_34132);
or U37649 (N_37649,N_30513,N_33779);
nand U37650 (N_37650,N_30583,N_31663);
or U37651 (N_37651,N_33236,N_33367);
or U37652 (N_37652,N_34865,N_32549);
xor U37653 (N_37653,N_32254,N_33341);
nand U37654 (N_37654,N_34698,N_33667);
nor U37655 (N_37655,N_31110,N_34184);
nor U37656 (N_37656,N_30805,N_32978);
or U37657 (N_37657,N_33977,N_31484);
xnor U37658 (N_37658,N_34351,N_34162);
or U37659 (N_37659,N_30442,N_33130);
or U37660 (N_37660,N_34525,N_33283);
xor U37661 (N_37661,N_30100,N_34778);
and U37662 (N_37662,N_33541,N_32859);
or U37663 (N_37663,N_33021,N_31514);
nor U37664 (N_37664,N_31701,N_30408);
or U37665 (N_37665,N_33005,N_30910);
xor U37666 (N_37666,N_33548,N_34467);
nand U37667 (N_37667,N_31432,N_31815);
xnor U37668 (N_37668,N_33550,N_31906);
nand U37669 (N_37669,N_32517,N_32777);
nand U37670 (N_37670,N_34342,N_30648);
xnor U37671 (N_37671,N_34098,N_34227);
xnor U37672 (N_37672,N_32691,N_31786);
nor U37673 (N_37673,N_31287,N_34949);
or U37674 (N_37674,N_33181,N_30400);
or U37675 (N_37675,N_32000,N_34803);
xor U37676 (N_37676,N_33015,N_31980);
nand U37677 (N_37677,N_32806,N_31621);
nor U37678 (N_37678,N_33856,N_30966);
nor U37679 (N_37679,N_31120,N_31011);
nor U37680 (N_37680,N_30010,N_34925);
nand U37681 (N_37681,N_31888,N_32304);
xor U37682 (N_37682,N_31563,N_32138);
nand U37683 (N_37683,N_32847,N_32019);
xor U37684 (N_37684,N_32688,N_34073);
and U37685 (N_37685,N_30111,N_34180);
nand U37686 (N_37686,N_34976,N_34447);
or U37687 (N_37687,N_34632,N_32109);
nor U37688 (N_37688,N_34302,N_32556);
nand U37689 (N_37689,N_30699,N_30182);
and U37690 (N_37690,N_31183,N_30233);
nor U37691 (N_37691,N_33538,N_34495);
or U37692 (N_37692,N_33022,N_30078);
nand U37693 (N_37693,N_31629,N_31229);
nand U37694 (N_37694,N_30438,N_33787);
or U37695 (N_37695,N_33965,N_32146);
xor U37696 (N_37696,N_31262,N_34391);
nand U37697 (N_37697,N_34579,N_31668);
xnor U37698 (N_37698,N_31182,N_34318);
xnor U37699 (N_37699,N_30493,N_30913);
xnor U37700 (N_37700,N_33359,N_32713);
nand U37701 (N_37701,N_31052,N_33152);
and U37702 (N_37702,N_32741,N_30667);
or U37703 (N_37703,N_32734,N_30253);
and U37704 (N_37704,N_31485,N_33075);
and U37705 (N_37705,N_31448,N_31560);
xnor U37706 (N_37706,N_33390,N_33743);
nor U37707 (N_37707,N_31347,N_31553);
xor U37708 (N_37708,N_33946,N_32671);
and U37709 (N_37709,N_33634,N_32861);
or U37710 (N_37710,N_34087,N_33271);
or U37711 (N_37711,N_31782,N_34345);
xor U37712 (N_37712,N_32258,N_33171);
and U37713 (N_37713,N_34689,N_32662);
or U37714 (N_37714,N_34570,N_33313);
xor U37715 (N_37715,N_32865,N_33031);
xnor U37716 (N_37716,N_31458,N_32787);
or U37717 (N_37717,N_32873,N_34394);
nor U37718 (N_37718,N_33724,N_33901);
and U37719 (N_37719,N_31283,N_33732);
or U37720 (N_37720,N_32635,N_30240);
and U37721 (N_37721,N_34699,N_32740);
or U37722 (N_37722,N_33930,N_33839);
xor U37723 (N_37723,N_31268,N_32365);
and U37724 (N_37724,N_33615,N_34898);
nand U37725 (N_37725,N_31150,N_33992);
or U37726 (N_37726,N_32027,N_32745);
nor U37727 (N_37727,N_30088,N_33687);
nor U37728 (N_37728,N_30511,N_32447);
nand U37729 (N_37729,N_32425,N_32823);
or U37730 (N_37730,N_33520,N_31262);
nand U37731 (N_37731,N_33489,N_34789);
and U37732 (N_37732,N_32456,N_31168);
nor U37733 (N_37733,N_34592,N_33102);
nand U37734 (N_37734,N_31372,N_30664);
xor U37735 (N_37735,N_30823,N_31616);
and U37736 (N_37736,N_33164,N_31080);
or U37737 (N_37737,N_32130,N_33050);
and U37738 (N_37738,N_34048,N_33545);
nand U37739 (N_37739,N_32577,N_33912);
and U37740 (N_37740,N_32568,N_31816);
nor U37741 (N_37741,N_30404,N_34286);
nor U37742 (N_37742,N_32280,N_33889);
or U37743 (N_37743,N_34790,N_32267);
nand U37744 (N_37744,N_30445,N_30897);
nand U37745 (N_37745,N_34038,N_30369);
nand U37746 (N_37746,N_34480,N_34550);
nand U37747 (N_37747,N_33991,N_34399);
nor U37748 (N_37748,N_31344,N_33206);
nor U37749 (N_37749,N_30761,N_30152);
xnor U37750 (N_37750,N_30490,N_33118);
xnor U37751 (N_37751,N_34793,N_33505);
and U37752 (N_37752,N_34740,N_33551);
and U37753 (N_37753,N_34998,N_33585);
or U37754 (N_37754,N_34743,N_33029);
or U37755 (N_37755,N_32737,N_31741);
nand U37756 (N_37756,N_30065,N_30662);
xnor U37757 (N_37757,N_30110,N_31947);
nand U37758 (N_37758,N_33567,N_32219);
nand U37759 (N_37759,N_31826,N_33535);
nand U37760 (N_37760,N_33537,N_32624);
nor U37761 (N_37761,N_33288,N_34042);
nand U37762 (N_37762,N_31852,N_33449);
and U37763 (N_37763,N_31587,N_31167);
nand U37764 (N_37764,N_33522,N_30398);
and U37765 (N_37765,N_33444,N_32834);
and U37766 (N_37766,N_31946,N_34618);
and U37767 (N_37767,N_30516,N_32192);
xnor U37768 (N_37768,N_34818,N_31378);
and U37769 (N_37769,N_34766,N_30783);
or U37770 (N_37770,N_33592,N_33218);
xor U37771 (N_37771,N_32034,N_33269);
and U37772 (N_37772,N_32590,N_30669);
nor U37773 (N_37773,N_32009,N_30400);
nand U37774 (N_37774,N_31329,N_31094);
nor U37775 (N_37775,N_30518,N_30212);
or U37776 (N_37776,N_31661,N_33880);
nand U37777 (N_37777,N_34615,N_32628);
or U37778 (N_37778,N_33733,N_33715);
xor U37779 (N_37779,N_30870,N_32647);
nor U37780 (N_37780,N_31072,N_34315);
nor U37781 (N_37781,N_34691,N_31637);
nand U37782 (N_37782,N_31864,N_32330);
or U37783 (N_37783,N_30837,N_30864);
nand U37784 (N_37784,N_33422,N_31129);
or U37785 (N_37785,N_34995,N_31146);
and U37786 (N_37786,N_31710,N_34898);
nor U37787 (N_37787,N_34445,N_32253);
or U37788 (N_37788,N_34883,N_33212);
or U37789 (N_37789,N_31164,N_31224);
nor U37790 (N_37790,N_30147,N_34545);
and U37791 (N_37791,N_34618,N_30828);
xnor U37792 (N_37792,N_33532,N_30443);
or U37793 (N_37793,N_32770,N_32153);
nand U37794 (N_37794,N_31888,N_30742);
or U37795 (N_37795,N_31808,N_31242);
or U37796 (N_37796,N_31369,N_31605);
and U37797 (N_37797,N_34853,N_32309);
nor U37798 (N_37798,N_32576,N_30000);
xnor U37799 (N_37799,N_30846,N_32369);
or U37800 (N_37800,N_34188,N_30726);
nor U37801 (N_37801,N_30191,N_30265);
nand U37802 (N_37802,N_32371,N_31244);
xnor U37803 (N_37803,N_33631,N_31863);
nor U37804 (N_37804,N_31711,N_34548);
nor U37805 (N_37805,N_30681,N_34200);
nor U37806 (N_37806,N_32351,N_30290);
or U37807 (N_37807,N_34389,N_30460);
and U37808 (N_37808,N_30403,N_30325);
and U37809 (N_37809,N_33471,N_30208);
nor U37810 (N_37810,N_31649,N_30307);
xnor U37811 (N_37811,N_33287,N_33088);
nor U37812 (N_37812,N_32579,N_31826);
nor U37813 (N_37813,N_34184,N_33266);
nand U37814 (N_37814,N_34803,N_32318);
xnor U37815 (N_37815,N_34063,N_33795);
and U37816 (N_37816,N_33945,N_34098);
nand U37817 (N_37817,N_33205,N_34302);
nor U37818 (N_37818,N_32943,N_32001);
nand U37819 (N_37819,N_34409,N_34488);
or U37820 (N_37820,N_30287,N_34208);
and U37821 (N_37821,N_30646,N_33859);
nand U37822 (N_37822,N_32470,N_30278);
nand U37823 (N_37823,N_31122,N_30630);
or U37824 (N_37824,N_34673,N_32156);
nor U37825 (N_37825,N_32555,N_34268);
and U37826 (N_37826,N_34937,N_31741);
or U37827 (N_37827,N_30032,N_30220);
or U37828 (N_37828,N_30125,N_32054);
and U37829 (N_37829,N_33063,N_31971);
xor U37830 (N_37830,N_31208,N_30006);
nor U37831 (N_37831,N_31932,N_31813);
or U37832 (N_37832,N_34116,N_34289);
or U37833 (N_37833,N_30138,N_32973);
nand U37834 (N_37834,N_34134,N_30946);
or U37835 (N_37835,N_34337,N_33189);
and U37836 (N_37836,N_32701,N_34901);
nand U37837 (N_37837,N_33799,N_31959);
nand U37838 (N_37838,N_32857,N_33169);
or U37839 (N_37839,N_34572,N_34297);
nand U37840 (N_37840,N_32271,N_32260);
xnor U37841 (N_37841,N_32246,N_30986);
or U37842 (N_37842,N_30289,N_33873);
or U37843 (N_37843,N_32426,N_34402);
and U37844 (N_37844,N_31026,N_30165);
nand U37845 (N_37845,N_31600,N_33534);
or U37846 (N_37846,N_32888,N_33668);
nand U37847 (N_37847,N_30249,N_32335);
xnor U37848 (N_37848,N_31555,N_34340);
and U37849 (N_37849,N_30237,N_30363);
xnor U37850 (N_37850,N_34988,N_33138);
nor U37851 (N_37851,N_33693,N_30905);
nand U37852 (N_37852,N_31086,N_31542);
or U37853 (N_37853,N_31303,N_31321);
and U37854 (N_37854,N_32750,N_33707);
or U37855 (N_37855,N_30998,N_32975);
nor U37856 (N_37856,N_31655,N_32932);
or U37857 (N_37857,N_30822,N_31000);
nand U37858 (N_37858,N_33595,N_31357);
and U37859 (N_37859,N_32353,N_30702);
or U37860 (N_37860,N_31878,N_33363);
and U37861 (N_37861,N_32305,N_31816);
nand U37862 (N_37862,N_30420,N_31905);
nor U37863 (N_37863,N_33966,N_33838);
or U37864 (N_37864,N_31009,N_32772);
or U37865 (N_37865,N_31372,N_33597);
xnor U37866 (N_37866,N_30421,N_33480);
xor U37867 (N_37867,N_30034,N_33071);
nand U37868 (N_37868,N_33679,N_34045);
or U37869 (N_37869,N_31658,N_30534);
xor U37870 (N_37870,N_32820,N_33310);
nor U37871 (N_37871,N_31759,N_32872);
and U37872 (N_37872,N_30460,N_31320);
nor U37873 (N_37873,N_34288,N_32849);
nor U37874 (N_37874,N_34270,N_34893);
and U37875 (N_37875,N_31886,N_33438);
nor U37876 (N_37876,N_32801,N_31400);
nor U37877 (N_37877,N_34931,N_32585);
nand U37878 (N_37878,N_34240,N_31349);
or U37879 (N_37879,N_34175,N_31503);
nand U37880 (N_37880,N_30923,N_31476);
xnor U37881 (N_37881,N_31644,N_30457);
nand U37882 (N_37882,N_31927,N_31235);
or U37883 (N_37883,N_31799,N_30271);
nor U37884 (N_37884,N_33393,N_30496);
and U37885 (N_37885,N_31417,N_32077);
xnor U37886 (N_37886,N_32723,N_33593);
xor U37887 (N_37887,N_31990,N_30243);
nor U37888 (N_37888,N_31629,N_30518);
and U37889 (N_37889,N_33753,N_34300);
or U37890 (N_37890,N_30773,N_34770);
and U37891 (N_37891,N_33669,N_30681);
and U37892 (N_37892,N_32959,N_32861);
nor U37893 (N_37893,N_31089,N_31631);
nand U37894 (N_37894,N_31060,N_34778);
xor U37895 (N_37895,N_34676,N_33850);
xor U37896 (N_37896,N_34843,N_32004);
nand U37897 (N_37897,N_33735,N_30475);
xnor U37898 (N_37898,N_30731,N_32943);
and U37899 (N_37899,N_31049,N_31446);
or U37900 (N_37900,N_32705,N_32394);
and U37901 (N_37901,N_33466,N_34478);
or U37902 (N_37902,N_32489,N_30825);
nor U37903 (N_37903,N_30358,N_30640);
xor U37904 (N_37904,N_33107,N_34806);
nand U37905 (N_37905,N_33247,N_34118);
nand U37906 (N_37906,N_33051,N_33466);
xor U37907 (N_37907,N_33362,N_32817);
xor U37908 (N_37908,N_34696,N_31474);
and U37909 (N_37909,N_31368,N_33334);
and U37910 (N_37910,N_34557,N_32508);
nand U37911 (N_37911,N_31149,N_32219);
xor U37912 (N_37912,N_31850,N_30015);
xor U37913 (N_37913,N_34187,N_31421);
xnor U37914 (N_37914,N_31574,N_30382);
xnor U37915 (N_37915,N_30168,N_34053);
and U37916 (N_37916,N_34615,N_32362);
xnor U37917 (N_37917,N_32620,N_30400);
nand U37918 (N_37918,N_32088,N_32802);
or U37919 (N_37919,N_30467,N_31700);
nand U37920 (N_37920,N_31466,N_32510);
nand U37921 (N_37921,N_32102,N_32317);
and U37922 (N_37922,N_34282,N_30270);
and U37923 (N_37923,N_32622,N_31901);
and U37924 (N_37924,N_31453,N_34032);
or U37925 (N_37925,N_33262,N_30146);
nand U37926 (N_37926,N_32417,N_34010);
nand U37927 (N_37927,N_30995,N_30705);
or U37928 (N_37928,N_32767,N_30852);
nor U37929 (N_37929,N_30273,N_33592);
and U37930 (N_37930,N_33905,N_33921);
or U37931 (N_37931,N_31551,N_33586);
nor U37932 (N_37932,N_33742,N_33962);
nor U37933 (N_37933,N_31034,N_34259);
xor U37934 (N_37934,N_30397,N_31364);
nand U37935 (N_37935,N_34695,N_30560);
nand U37936 (N_37936,N_31075,N_33652);
or U37937 (N_37937,N_32838,N_34657);
or U37938 (N_37938,N_30804,N_31603);
nand U37939 (N_37939,N_30020,N_30742);
nand U37940 (N_37940,N_33918,N_30595);
nand U37941 (N_37941,N_30250,N_30434);
nand U37942 (N_37942,N_33516,N_34181);
and U37943 (N_37943,N_30892,N_32702);
xnor U37944 (N_37944,N_31261,N_33711);
and U37945 (N_37945,N_33003,N_31399);
and U37946 (N_37946,N_31160,N_30450);
nor U37947 (N_37947,N_34137,N_32899);
and U37948 (N_37948,N_33756,N_33432);
or U37949 (N_37949,N_32791,N_30425);
and U37950 (N_37950,N_33267,N_34742);
xnor U37951 (N_37951,N_33504,N_32414);
or U37952 (N_37952,N_31462,N_30556);
nor U37953 (N_37953,N_32640,N_32292);
xnor U37954 (N_37954,N_34314,N_30535);
xor U37955 (N_37955,N_30078,N_32810);
or U37956 (N_37956,N_32903,N_32592);
and U37957 (N_37957,N_31938,N_34129);
nor U37958 (N_37958,N_33149,N_31211);
xor U37959 (N_37959,N_31825,N_30536);
or U37960 (N_37960,N_31710,N_31758);
nand U37961 (N_37961,N_31809,N_34271);
or U37962 (N_37962,N_31045,N_34422);
nor U37963 (N_37963,N_33467,N_34640);
or U37964 (N_37964,N_31152,N_33522);
or U37965 (N_37965,N_32926,N_32805);
nand U37966 (N_37966,N_30045,N_33315);
nand U37967 (N_37967,N_33585,N_33231);
xor U37968 (N_37968,N_32290,N_34710);
nand U37969 (N_37969,N_32818,N_34320);
and U37970 (N_37970,N_32870,N_34654);
or U37971 (N_37971,N_34422,N_31051);
and U37972 (N_37972,N_33450,N_30297);
nand U37973 (N_37973,N_30137,N_30375);
or U37974 (N_37974,N_32058,N_33695);
or U37975 (N_37975,N_32182,N_30289);
nand U37976 (N_37976,N_33504,N_32520);
nor U37977 (N_37977,N_30394,N_31885);
or U37978 (N_37978,N_30604,N_33989);
nor U37979 (N_37979,N_33291,N_34770);
xnor U37980 (N_37980,N_34521,N_32072);
xnor U37981 (N_37981,N_30703,N_30116);
xor U37982 (N_37982,N_34215,N_34049);
xnor U37983 (N_37983,N_32022,N_33838);
nor U37984 (N_37984,N_33846,N_34045);
and U37985 (N_37985,N_33002,N_34065);
xnor U37986 (N_37986,N_31638,N_32783);
and U37987 (N_37987,N_30444,N_33751);
nor U37988 (N_37988,N_31634,N_33306);
xnor U37989 (N_37989,N_31385,N_32736);
and U37990 (N_37990,N_34644,N_33386);
and U37991 (N_37991,N_33761,N_32934);
nand U37992 (N_37992,N_33327,N_33829);
nor U37993 (N_37993,N_33484,N_32039);
xnor U37994 (N_37994,N_34338,N_33458);
nor U37995 (N_37995,N_33633,N_32689);
or U37996 (N_37996,N_31941,N_31426);
and U37997 (N_37997,N_31543,N_34478);
nand U37998 (N_37998,N_34475,N_32946);
and U37999 (N_37999,N_31351,N_32784);
nor U38000 (N_38000,N_33759,N_32412);
xor U38001 (N_38001,N_31563,N_32100);
and U38002 (N_38002,N_32347,N_34276);
and U38003 (N_38003,N_32116,N_33131);
nor U38004 (N_38004,N_31861,N_32704);
nor U38005 (N_38005,N_30158,N_30467);
and U38006 (N_38006,N_33576,N_33004);
and U38007 (N_38007,N_31628,N_31508);
nand U38008 (N_38008,N_31010,N_34908);
or U38009 (N_38009,N_33249,N_33634);
or U38010 (N_38010,N_34160,N_31731);
or U38011 (N_38011,N_31733,N_34895);
or U38012 (N_38012,N_31696,N_30363);
xnor U38013 (N_38013,N_32553,N_30174);
or U38014 (N_38014,N_32294,N_33647);
or U38015 (N_38015,N_32490,N_31695);
nand U38016 (N_38016,N_31125,N_33284);
nand U38017 (N_38017,N_32000,N_34779);
nor U38018 (N_38018,N_30609,N_30837);
or U38019 (N_38019,N_31840,N_32339);
nand U38020 (N_38020,N_33527,N_33727);
xnor U38021 (N_38021,N_33214,N_31555);
and U38022 (N_38022,N_30518,N_34315);
xor U38023 (N_38023,N_32270,N_32872);
nand U38024 (N_38024,N_31187,N_34009);
xor U38025 (N_38025,N_34938,N_31612);
or U38026 (N_38026,N_32178,N_32772);
and U38027 (N_38027,N_34935,N_34892);
nand U38028 (N_38028,N_32936,N_32056);
or U38029 (N_38029,N_30505,N_34424);
nor U38030 (N_38030,N_32847,N_30998);
xor U38031 (N_38031,N_34485,N_34201);
nor U38032 (N_38032,N_31290,N_32721);
nor U38033 (N_38033,N_33406,N_30934);
nor U38034 (N_38034,N_31151,N_30097);
nand U38035 (N_38035,N_30188,N_31532);
xnor U38036 (N_38036,N_34051,N_30325);
nand U38037 (N_38037,N_32622,N_34235);
or U38038 (N_38038,N_31559,N_34637);
nand U38039 (N_38039,N_30097,N_30963);
or U38040 (N_38040,N_30237,N_30711);
or U38041 (N_38041,N_33370,N_32923);
nand U38042 (N_38042,N_31080,N_32143);
nand U38043 (N_38043,N_30752,N_33467);
nor U38044 (N_38044,N_30718,N_32591);
and U38045 (N_38045,N_31008,N_34772);
or U38046 (N_38046,N_34963,N_30856);
or U38047 (N_38047,N_33600,N_32929);
and U38048 (N_38048,N_34227,N_32122);
nor U38049 (N_38049,N_34618,N_31630);
nand U38050 (N_38050,N_30786,N_33868);
nand U38051 (N_38051,N_32844,N_33207);
or U38052 (N_38052,N_34599,N_30551);
nor U38053 (N_38053,N_33843,N_31835);
xnor U38054 (N_38054,N_30002,N_34670);
and U38055 (N_38055,N_33228,N_33361);
and U38056 (N_38056,N_34958,N_31871);
nor U38057 (N_38057,N_30863,N_31699);
and U38058 (N_38058,N_30502,N_32141);
nor U38059 (N_38059,N_31612,N_33674);
nor U38060 (N_38060,N_31936,N_30962);
nor U38061 (N_38061,N_34802,N_32313);
and U38062 (N_38062,N_31445,N_30580);
nor U38063 (N_38063,N_31187,N_33305);
xor U38064 (N_38064,N_31520,N_33007);
nand U38065 (N_38065,N_30879,N_33056);
xor U38066 (N_38066,N_31982,N_33018);
or U38067 (N_38067,N_32691,N_34603);
xnor U38068 (N_38068,N_30264,N_33171);
or U38069 (N_38069,N_30442,N_31400);
nor U38070 (N_38070,N_33295,N_34455);
nor U38071 (N_38071,N_31805,N_31083);
nand U38072 (N_38072,N_30806,N_34206);
nor U38073 (N_38073,N_33824,N_30956);
or U38074 (N_38074,N_33323,N_31312);
nand U38075 (N_38075,N_34084,N_34056);
nor U38076 (N_38076,N_33749,N_31528);
and U38077 (N_38077,N_32055,N_31758);
xnor U38078 (N_38078,N_34209,N_34171);
xnor U38079 (N_38079,N_33779,N_32866);
xnor U38080 (N_38080,N_32633,N_31428);
nand U38081 (N_38081,N_34778,N_30534);
and U38082 (N_38082,N_34592,N_33384);
nor U38083 (N_38083,N_31602,N_32861);
or U38084 (N_38084,N_31554,N_34188);
and U38085 (N_38085,N_33263,N_33143);
xnor U38086 (N_38086,N_33438,N_34537);
or U38087 (N_38087,N_30511,N_34033);
nand U38088 (N_38088,N_33109,N_32625);
nor U38089 (N_38089,N_32610,N_32895);
xnor U38090 (N_38090,N_32706,N_32658);
and U38091 (N_38091,N_34156,N_30378);
or U38092 (N_38092,N_34865,N_30226);
nand U38093 (N_38093,N_33725,N_31659);
and U38094 (N_38094,N_32365,N_31153);
nand U38095 (N_38095,N_30912,N_32365);
nor U38096 (N_38096,N_34462,N_34474);
and U38097 (N_38097,N_30610,N_30139);
or U38098 (N_38098,N_34858,N_30891);
or U38099 (N_38099,N_32504,N_32421);
and U38100 (N_38100,N_34306,N_34551);
nor U38101 (N_38101,N_33112,N_31028);
or U38102 (N_38102,N_34756,N_30590);
and U38103 (N_38103,N_34378,N_31615);
or U38104 (N_38104,N_32027,N_31228);
nor U38105 (N_38105,N_30697,N_32846);
and U38106 (N_38106,N_30844,N_31420);
or U38107 (N_38107,N_34092,N_31765);
or U38108 (N_38108,N_32108,N_34364);
or U38109 (N_38109,N_33034,N_33110);
or U38110 (N_38110,N_31287,N_31607);
or U38111 (N_38111,N_32882,N_33460);
and U38112 (N_38112,N_32195,N_31870);
nand U38113 (N_38113,N_30140,N_31147);
nand U38114 (N_38114,N_34848,N_30589);
nor U38115 (N_38115,N_30499,N_33745);
and U38116 (N_38116,N_32803,N_34970);
xor U38117 (N_38117,N_33148,N_33966);
nand U38118 (N_38118,N_32251,N_30755);
or U38119 (N_38119,N_31476,N_34832);
xnor U38120 (N_38120,N_32019,N_32932);
nor U38121 (N_38121,N_31375,N_31724);
or U38122 (N_38122,N_33065,N_30903);
xnor U38123 (N_38123,N_32921,N_34223);
and U38124 (N_38124,N_33379,N_33204);
xor U38125 (N_38125,N_32358,N_30113);
or U38126 (N_38126,N_34268,N_30808);
nor U38127 (N_38127,N_31305,N_31637);
or U38128 (N_38128,N_31976,N_32705);
or U38129 (N_38129,N_30726,N_33743);
or U38130 (N_38130,N_31377,N_30530);
xor U38131 (N_38131,N_30199,N_32736);
or U38132 (N_38132,N_32488,N_31878);
nor U38133 (N_38133,N_31806,N_32096);
xor U38134 (N_38134,N_30929,N_33749);
or U38135 (N_38135,N_31110,N_31401);
nand U38136 (N_38136,N_30813,N_30262);
or U38137 (N_38137,N_31088,N_31585);
and U38138 (N_38138,N_31125,N_30627);
or U38139 (N_38139,N_34234,N_31748);
and U38140 (N_38140,N_33446,N_32306);
nor U38141 (N_38141,N_30049,N_30437);
or U38142 (N_38142,N_33571,N_30417);
and U38143 (N_38143,N_30102,N_30854);
xnor U38144 (N_38144,N_33624,N_31136);
nand U38145 (N_38145,N_30526,N_31647);
and U38146 (N_38146,N_33847,N_31722);
and U38147 (N_38147,N_30574,N_30599);
and U38148 (N_38148,N_31688,N_34420);
and U38149 (N_38149,N_33916,N_30486);
nand U38150 (N_38150,N_31587,N_30231);
and U38151 (N_38151,N_32787,N_32773);
nor U38152 (N_38152,N_30033,N_31735);
xnor U38153 (N_38153,N_30971,N_31846);
nand U38154 (N_38154,N_30628,N_32203);
or U38155 (N_38155,N_33961,N_31013);
nand U38156 (N_38156,N_33425,N_34970);
xor U38157 (N_38157,N_31101,N_31523);
nand U38158 (N_38158,N_31498,N_32375);
nand U38159 (N_38159,N_32133,N_30739);
nand U38160 (N_38160,N_32743,N_34766);
and U38161 (N_38161,N_30644,N_32420);
nor U38162 (N_38162,N_32510,N_33844);
nand U38163 (N_38163,N_30998,N_30747);
nand U38164 (N_38164,N_31103,N_33341);
xor U38165 (N_38165,N_34459,N_33275);
nor U38166 (N_38166,N_34455,N_31259);
nor U38167 (N_38167,N_31897,N_34799);
and U38168 (N_38168,N_32411,N_32182);
or U38169 (N_38169,N_31834,N_34975);
nand U38170 (N_38170,N_32147,N_30554);
xor U38171 (N_38171,N_34947,N_34112);
nor U38172 (N_38172,N_30362,N_34859);
nor U38173 (N_38173,N_30323,N_32904);
nand U38174 (N_38174,N_31526,N_34541);
xnor U38175 (N_38175,N_30828,N_31683);
and U38176 (N_38176,N_30482,N_33347);
nand U38177 (N_38177,N_33765,N_33784);
xnor U38178 (N_38178,N_30101,N_32708);
or U38179 (N_38179,N_33806,N_33180);
xor U38180 (N_38180,N_30050,N_34750);
nand U38181 (N_38181,N_33745,N_31453);
or U38182 (N_38182,N_32335,N_34294);
and U38183 (N_38183,N_34511,N_30041);
nor U38184 (N_38184,N_32809,N_31869);
nand U38185 (N_38185,N_33919,N_32742);
and U38186 (N_38186,N_34045,N_32493);
or U38187 (N_38187,N_34893,N_32527);
nor U38188 (N_38188,N_30949,N_34168);
and U38189 (N_38189,N_34956,N_34032);
nand U38190 (N_38190,N_34745,N_34255);
nand U38191 (N_38191,N_34937,N_32616);
nand U38192 (N_38192,N_30223,N_33803);
nor U38193 (N_38193,N_30810,N_33757);
xor U38194 (N_38194,N_30230,N_34037);
nor U38195 (N_38195,N_33094,N_32847);
or U38196 (N_38196,N_32127,N_31284);
xor U38197 (N_38197,N_34619,N_33791);
nand U38198 (N_38198,N_33932,N_30917);
nor U38199 (N_38199,N_30500,N_30719);
xor U38200 (N_38200,N_34138,N_34196);
nand U38201 (N_38201,N_33912,N_32785);
xnor U38202 (N_38202,N_31345,N_33733);
or U38203 (N_38203,N_32760,N_34818);
xor U38204 (N_38204,N_32486,N_32112);
nor U38205 (N_38205,N_34882,N_32471);
xor U38206 (N_38206,N_32075,N_34775);
xor U38207 (N_38207,N_31514,N_31893);
xnor U38208 (N_38208,N_34713,N_30915);
xnor U38209 (N_38209,N_31248,N_34517);
nand U38210 (N_38210,N_32342,N_33485);
nor U38211 (N_38211,N_33759,N_32896);
nand U38212 (N_38212,N_30342,N_31077);
nor U38213 (N_38213,N_30296,N_33539);
xnor U38214 (N_38214,N_31865,N_34898);
nor U38215 (N_38215,N_34914,N_31105);
nand U38216 (N_38216,N_34568,N_33230);
nand U38217 (N_38217,N_32203,N_31251);
or U38218 (N_38218,N_30539,N_32019);
and U38219 (N_38219,N_34823,N_31446);
or U38220 (N_38220,N_33860,N_34037);
or U38221 (N_38221,N_32314,N_31153);
and U38222 (N_38222,N_30379,N_31064);
nor U38223 (N_38223,N_31981,N_32609);
xor U38224 (N_38224,N_31102,N_34912);
or U38225 (N_38225,N_34044,N_30962);
xor U38226 (N_38226,N_31748,N_33952);
xor U38227 (N_38227,N_33527,N_32320);
xnor U38228 (N_38228,N_31163,N_33344);
nor U38229 (N_38229,N_34770,N_30708);
and U38230 (N_38230,N_31659,N_31526);
nor U38231 (N_38231,N_31144,N_31585);
and U38232 (N_38232,N_33925,N_32688);
xnor U38233 (N_38233,N_30050,N_30083);
nand U38234 (N_38234,N_31892,N_31787);
and U38235 (N_38235,N_34854,N_34904);
and U38236 (N_38236,N_31241,N_31804);
xnor U38237 (N_38237,N_34628,N_32310);
and U38238 (N_38238,N_34457,N_33947);
or U38239 (N_38239,N_31058,N_33702);
and U38240 (N_38240,N_33749,N_32030);
nor U38241 (N_38241,N_32603,N_34071);
xnor U38242 (N_38242,N_32530,N_30701);
nor U38243 (N_38243,N_34443,N_30200);
nor U38244 (N_38244,N_34876,N_31366);
nand U38245 (N_38245,N_31382,N_31977);
or U38246 (N_38246,N_32972,N_31535);
nand U38247 (N_38247,N_31594,N_32926);
nand U38248 (N_38248,N_33260,N_34023);
nor U38249 (N_38249,N_33579,N_31813);
nor U38250 (N_38250,N_33014,N_31992);
or U38251 (N_38251,N_32209,N_33291);
nand U38252 (N_38252,N_31609,N_33733);
nor U38253 (N_38253,N_31303,N_32929);
and U38254 (N_38254,N_33064,N_34435);
or U38255 (N_38255,N_33555,N_31460);
and U38256 (N_38256,N_30190,N_33915);
and U38257 (N_38257,N_30671,N_32248);
or U38258 (N_38258,N_32947,N_31245);
nor U38259 (N_38259,N_34588,N_33144);
nor U38260 (N_38260,N_30660,N_33886);
xnor U38261 (N_38261,N_32083,N_33839);
nand U38262 (N_38262,N_32167,N_33979);
and U38263 (N_38263,N_30841,N_30566);
and U38264 (N_38264,N_33067,N_34533);
nor U38265 (N_38265,N_31467,N_33086);
and U38266 (N_38266,N_34057,N_31427);
nand U38267 (N_38267,N_30467,N_33608);
nor U38268 (N_38268,N_31101,N_30985);
or U38269 (N_38269,N_34320,N_30281);
nor U38270 (N_38270,N_31170,N_31576);
xor U38271 (N_38271,N_32527,N_34010);
or U38272 (N_38272,N_32325,N_33753);
or U38273 (N_38273,N_30608,N_31403);
xor U38274 (N_38274,N_33268,N_33328);
nor U38275 (N_38275,N_33105,N_33933);
or U38276 (N_38276,N_30362,N_30020);
xnor U38277 (N_38277,N_33811,N_33875);
or U38278 (N_38278,N_31950,N_32042);
and U38279 (N_38279,N_32614,N_32157);
and U38280 (N_38280,N_34165,N_31798);
xor U38281 (N_38281,N_33128,N_34077);
and U38282 (N_38282,N_30869,N_32840);
xnor U38283 (N_38283,N_33927,N_31012);
nor U38284 (N_38284,N_33662,N_31688);
nor U38285 (N_38285,N_32447,N_34026);
nand U38286 (N_38286,N_30421,N_32651);
nor U38287 (N_38287,N_32014,N_33375);
nor U38288 (N_38288,N_32560,N_31391);
nand U38289 (N_38289,N_33262,N_31767);
nand U38290 (N_38290,N_31979,N_34326);
xnor U38291 (N_38291,N_30495,N_30110);
and U38292 (N_38292,N_32214,N_33665);
or U38293 (N_38293,N_31480,N_33461);
or U38294 (N_38294,N_31450,N_31153);
nor U38295 (N_38295,N_31416,N_33357);
nand U38296 (N_38296,N_33496,N_31088);
nand U38297 (N_38297,N_33835,N_32851);
or U38298 (N_38298,N_30972,N_33766);
and U38299 (N_38299,N_31076,N_33811);
nand U38300 (N_38300,N_32234,N_34131);
nand U38301 (N_38301,N_34128,N_32149);
nor U38302 (N_38302,N_31768,N_30849);
nor U38303 (N_38303,N_32563,N_32942);
or U38304 (N_38304,N_32379,N_31506);
nand U38305 (N_38305,N_32721,N_33670);
or U38306 (N_38306,N_31546,N_34423);
xor U38307 (N_38307,N_32733,N_30353);
nand U38308 (N_38308,N_31346,N_34652);
or U38309 (N_38309,N_31926,N_30196);
nand U38310 (N_38310,N_32973,N_30017);
nand U38311 (N_38311,N_30577,N_32384);
nand U38312 (N_38312,N_32798,N_31380);
nor U38313 (N_38313,N_30179,N_33873);
nand U38314 (N_38314,N_30808,N_33808);
or U38315 (N_38315,N_30406,N_30965);
xnor U38316 (N_38316,N_34292,N_33969);
xor U38317 (N_38317,N_31027,N_31245);
nor U38318 (N_38318,N_33793,N_32042);
and U38319 (N_38319,N_34469,N_32348);
nand U38320 (N_38320,N_30219,N_33550);
xnor U38321 (N_38321,N_32179,N_33604);
nor U38322 (N_38322,N_34929,N_33071);
nor U38323 (N_38323,N_31138,N_33146);
and U38324 (N_38324,N_31510,N_31046);
xor U38325 (N_38325,N_34132,N_34704);
nand U38326 (N_38326,N_30773,N_32617);
xor U38327 (N_38327,N_31915,N_33229);
and U38328 (N_38328,N_32053,N_31663);
xnor U38329 (N_38329,N_31603,N_34708);
or U38330 (N_38330,N_32104,N_33350);
nor U38331 (N_38331,N_32295,N_32363);
nand U38332 (N_38332,N_34188,N_31237);
nand U38333 (N_38333,N_30562,N_31430);
xor U38334 (N_38334,N_31415,N_34295);
and U38335 (N_38335,N_32748,N_31199);
xnor U38336 (N_38336,N_31991,N_34495);
nand U38337 (N_38337,N_34125,N_30196);
nand U38338 (N_38338,N_30530,N_32877);
or U38339 (N_38339,N_30222,N_31193);
nor U38340 (N_38340,N_31903,N_31978);
and U38341 (N_38341,N_33479,N_30654);
and U38342 (N_38342,N_31966,N_34589);
or U38343 (N_38343,N_32319,N_33197);
xor U38344 (N_38344,N_30833,N_34882);
nand U38345 (N_38345,N_34132,N_31705);
or U38346 (N_38346,N_31426,N_32857);
xor U38347 (N_38347,N_32820,N_31048);
xor U38348 (N_38348,N_34131,N_32309);
nor U38349 (N_38349,N_31397,N_31424);
or U38350 (N_38350,N_34780,N_34424);
and U38351 (N_38351,N_33570,N_34516);
xor U38352 (N_38352,N_30915,N_32319);
nand U38353 (N_38353,N_33331,N_34428);
xnor U38354 (N_38354,N_34008,N_32218);
or U38355 (N_38355,N_31842,N_33635);
nand U38356 (N_38356,N_33538,N_31440);
nand U38357 (N_38357,N_31156,N_33887);
xor U38358 (N_38358,N_32244,N_33418);
nand U38359 (N_38359,N_33362,N_31464);
or U38360 (N_38360,N_33922,N_32981);
and U38361 (N_38361,N_31312,N_32684);
or U38362 (N_38362,N_34238,N_34185);
nor U38363 (N_38363,N_30392,N_30751);
nand U38364 (N_38364,N_33827,N_31693);
or U38365 (N_38365,N_34567,N_34884);
or U38366 (N_38366,N_31558,N_33479);
and U38367 (N_38367,N_30660,N_33029);
nor U38368 (N_38368,N_34360,N_34553);
and U38369 (N_38369,N_33030,N_34357);
or U38370 (N_38370,N_33166,N_32268);
or U38371 (N_38371,N_32910,N_33711);
or U38372 (N_38372,N_33140,N_32484);
nor U38373 (N_38373,N_31192,N_31449);
nand U38374 (N_38374,N_34607,N_30103);
xnor U38375 (N_38375,N_32084,N_33227);
xor U38376 (N_38376,N_30827,N_32705);
and U38377 (N_38377,N_34463,N_30005);
or U38378 (N_38378,N_33216,N_30357);
or U38379 (N_38379,N_30264,N_34703);
nor U38380 (N_38380,N_32530,N_32874);
xnor U38381 (N_38381,N_34261,N_31607);
nand U38382 (N_38382,N_32137,N_34751);
nor U38383 (N_38383,N_31284,N_33341);
nand U38384 (N_38384,N_33853,N_30199);
nor U38385 (N_38385,N_34064,N_31048);
xnor U38386 (N_38386,N_34372,N_33960);
nor U38387 (N_38387,N_32623,N_32113);
and U38388 (N_38388,N_32476,N_33214);
nand U38389 (N_38389,N_33926,N_33257);
xnor U38390 (N_38390,N_32480,N_32761);
and U38391 (N_38391,N_34276,N_31030);
and U38392 (N_38392,N_33531,N_31350);
xor U38393 (N_38393,N_33177,N_33144);
and U38394 (N_38394,N_30636,N_34336);
or U38395 (N_38395,N_30167,N_32570);
xnor U38396 (N_38396,N_32368,N_33203);
xnor U38397 (N_38397,N_32584,N_32757);
xnor U38398 (N_38398,N_31702,N_32342);
nor U38399 (N_38399,N_34166,N_32323);
nor U38400 (N_38400,N_32784,N_32209);
nand U38401 (N_38401,N_33503,N_30610);
nand U38402 (N_38402,N_32155,N_31284);
and U38403 (N_38403,N_32571,N_32844);
nand U38404 (N_38404,N_31342,N_33816);
nand U38405 (N_38405,N_34156,N_34418);
and U38406 (N_38406,N_31183,N_30534);
or U38407 (N_38407,N_30779,N_34017);
nor U38408 (N_38408,N_34978,N_33317);
xor U38409 (N_38409,N_32965,N_31371);
nor U38410 (N_38410,N_30868,N_33189);
or U38411 (N_38411,N_34305,N_33203);
and U38412 (N_38412,N_33486,N_32894);
nor U38413 (N_38413,N_31814,N_30082);
nor U38414 (N_38414,N_31864,N_30422);
or U38415 (N_38415,N_30752,N_33159);
and U38416 (N_38416,N_30652,N_34671);
nand U38417 (N_38417,N_34145,N_30557);
nor U38418 (N_38418,N_31754,N_34334);
nor U38419 (N_38419,N_32471,N_30140);
nand U38420 (N_38420,N_31620,N_34702);
or U38421 (N_38421,N_31795,N_33581);
and U38422 (N_38422,N_30815,N_34101);
xnor U38423 (N_38423,N_31644,N_33134);
and U38424 (N_38424,N_34010,N_33133);
nand U38425 (N_38425,N_33604,N_31727);
nor U38426 (N_38426,N_30108,N_34999);
or U38427 (N_38427,N_30728,N_32061);
nor U38428 (N_38428,N_33290,N_32235);
nand U38429 (N_38429,N_30622,N_30211);
and U38430 (N_38430,N_34878,N_32749);
or U38431 (N_38431,N_32212,N_33339);
nand U38432 (N_38432,N_34170,N_32955);
nand U38433 (N_38433,N_34509,N_30389);
or U38434 (N_38434,N_34531,N_34795);
nor U38435 (N_38435,N_30612,N_31764);
xnor U38436 (N_38436,N_31628,N_31680);
and U38437 (N_38437,N_34939,N_33063);
nand U38438 (N_38438,N_33720,N_32495);
and U38439 (N_38439,N_32679,N_31097);
or U38440 (N_38440,N_30528,N_33383);
and U38441 (N_38441,N_30130,N_33030);
xnor U38442 (N_38442,N_32942,N_34740);
xor U38443 (N_38443,N_31386,N_34955);
and U38444 (N_38444,N_34459,N_30192);
nor U38445 (N_38445,N_33029,N_33053);
xor U38446 (N_38446,N_30727,N_32804);
and U38447 (N_38447,N_30160,N_30503);
or U38448 (N_38448,N_33052,N_34598);
and U38449 (N_38449,N_30193,N_32332);
and U38450 (N_38450,N_30060,N_33805);
and U38451 (N_38451,N_30793,N_31120);
xor U38452 (N_38452,N_34874,N_33291);
or U38453 (N_38453,N_30336,N_30379);
or U38454 (N_38454,N_31060,N_33971);
nor U38455 (N_38455,N_31531,N_33847);
nand U38456 (N_38456,N_32732,N_33116);
and U38457 (N_38457,N_34319,N_32976);
and U38458 (N_38458,N_34866,N_31169);
xor U38459 (N_38459,N_31659,N_34365);
and U38460 (N_38460,N_33536,N_34526);
nand U38461 (N_38461,N_34916,N_31978);
or U38462 (N_38462,N_32763,N_31655);
nand U38463 (N_38463,N_34739,N_34938);
nand U38464 (N_38464,N_34262,N_32817);
and U38465 (N_38465,N_32490,N_30688);
or U38466 (N_38466,N_33596,N_34045);
nand U38467 (N_38467,N_34906,N_31695);
xnor U38468 (N_38468,N_34792,N_34811);
and U38469 (N_38469,N_30975,N_33746);
nor U38470 (N_38470,N_33724,N_34808);
nand U38471 (N_38471,N_33906,N_33061);
nand U38472 (N_38472,N_32002,N_31333);
and U38473 (N_38473,N_32568,N_30470);
nor U38474 (N_38474,N_34236,N_30289);
and U38475 (N_38475,N_34309,N_32608);
xor U38476 (N_38476,N_32587,N_30929);
and U38477 (N_38477,N_30492,N_31055);
xnor U38478 (N_38478,N_33735,N_33019);
nor U38479 (N_38479,N_32858,N_33231);
or U38480 (N_38480,N_33667,N_34791);
and U38481 (N_38481,N_34246,N_31528);
and U38482 (N_38482,N_33342,N_33029);
xor U38483 (N_38483,N_34810,N_31884);
xnor U38484 (N_38484,N_30237,N_31059);
xor U38485 (N_38485,N_34789,N_33531);
and U38486 (N_38486,N_32453,N_30520);
and U38487 (N_38487,N_30415,N_31911);
and U38488 (N_38488,N_31565,N_30061);
xor U38489 (N_38489,N_32079,N_30151);
or U38490 (N_38490,N_32424,N_31437);
or U38491 (N_38491,N_31416,N_33651);
and U38492 (N_38492,N_32391,N_32626);
and U38493 (N_38493,N_33217,N_31392);
nor U38494 (N_38494,N_30610,N_32144);
and U38495 (N_38495,N_30047,N_34705);
and U38496 (N_38496,N_31045,N_33299);
nand U38497 (N_38497,N_32994,N_30749);
nand U38498 (N_38498,N_33369,N_32952);
nor U38499 (N_38499,N_30152,N_30239);
and U38500 (N_38500,N_30939,N_33617);
nor U38501 (N_38501,N_30811,N_32785);
nor U38502 (N_38502,N_32863,N_30785);
nand U38503 (N_38503,N_33816,N_33781);
nor U38504 (N_38504,N_30834,N_33914);
and U38505 (N_38505,N_32260,N_30088);
xnor U38506 (N_38506,N_34016,N_31130);
and U38507 (N_38507,N_31721,N_33337);
or U38508 (N_38508,N_32569,N_30038);
nor U38509 (N_38509,N_30992,N_31621);
nand U38510 (N_38510,N_31805,N_34407);
and U38511 (N_38511,N_33091,N_33220);
xor U38512 (N_38512,N_32941,N_33909);
nor U38513 (N_38513,N_32436,N_34845);
nor U38514 (N_38514,N_33787,N_33124);
or U38515 (N_38515,N_30488,N_33678);
nand U38516 (N_38516,N_31766,N_32108);
xor U38517 (N_38517,N_30634,N_30005);
nor U38518 (N_38518,N_33229,N_31338);
nand U38519 (N_38519,N_30662,N_32981);
nand U38520 (N_38520,N_31502,N_31305);
and U38521 (N_38521,N_32803,N_32982);
nor U38522 (N_38522,N_31488,N_30859);
and U38523 (N_38523,N_31788,N_31689);
or U38524 (N_38524,N_32882,N_33500);
xor U38525 (N_38525,N_31184,N_32777);
nor U38526 (N_38526,N_33922,N_32893);
nand U38527 (N_38527,N_31242,N_31804);
or U38528 (N_38528,N_30010,N_33451);
nor U38529 (N_38529,N_32578,N_30422);
xnor U38530 (N_38530,N_31030,N_33103);
and U38531 (N_38531,N_33502,N_34594);
and U38532 (N_38532,N_34914,N_32345);
xnor U38533 (N_38533,N_31383,N_33255);
xnor U38534 (N_38534,N_34112,N_34540);
and U38535 (N_38535,N_31724,N_30134);
nand U38536 (N_38536,N_32503,N_33362);
xnor U38537 (N_38537,N_31241,N_32940);
nor U38538 (N_38538,N_33400,N_31052);
xnor U38539 (N_38539,N_31482,N_34210);
or U38540 (N_38540,N_31925,N_30361);
or U38541 (N_38541,N_30773,N_31292);
nand U38542 (N_38542,N_32786,N_30705);
nand U38543 (N_38543,N_30912,N_30801);
or U38544 (N_38544,N_30412,N_34325);
or U38545 (N_38545,N_30078,N_30440);
nand U38546 (N_38546,N_31659,N_30042);
nor U38547 (N_38547,N_32240,N_33051);
xnor U38548 (N_38548,N_33831,N_31266);
and U38549 (N_38549,N_32963,N_30882);
and U38550 (N_38550,N_31390,N_31551);
nor U38551 (N_38551,N_33502,N_32473);
or U38552 (N_38552,N_32057,N_32299);
or U38553 (N_38553,N_30577,N_31551);
nand U38554 (N_38554,N_30999,N_34974);
nor U38555 (N_38555,N_32173,N_30201);
nor U38556 (N_38556,N_31162,N_33540);
or U38557 (N_38557,N_33553,N_33709);
xor U38558 (N_38558,N_30819,N_30814);
and U38559 (N_38559,N_31191,N_31740);
nand U38560 (N_38560,N_34510,N_32623);
and U38561 (N_38561,N_34002,N_31465);
and U38562 (N_38562,N_30744,N_33946);
xnor U38563 (N_38563,N_32230,N_34457);
nand U38564 (N_38564,N_33238,N_30549);
and U38565 (N_38565,N_33833,N_30909);
or U38566 (N_38566,N_33610,N_34222);
nor U38567 (N_38567,N_32447,N_32625);
and U38568 (N_38568,N_34313,N_33309);
xnor U38569 (N_38569,N_31894,N_30280);
xnor U38570 (N_38570,N_33271,N_30093);
xnor U38571 (N_38571,N_34397,N_33467);
or U38572 (N_38572,N_34891,N_32987);
or U38573 (N_38573,N_34568,N_31334);
nor U38574 (N_38574,N_31463,N_32102);
xnor U38575 (N_38575,N_34527,N_31643);
xnor U38576 (N_38576,N_33444,N_32642);
or U38577 (N_38577,N_30295,N_31594);
nand U38578 (N_38578,N_33920,N_31894);
nor U38579 (N_38579,N_31281,N_31767);
and U38580 (N_38580,N_33998,N_30519);
nor U38581 (N_38581,N_34069,N_31414);
nand U38582 (N_38582,N_33156,N_32037);
nand U38583 (N_38583,N_30779,N_32764);
nor U38584 (N_38584,N_32948,N_31194);
xnor U38585 (N_38585,N_33254,N_32816);
or U38586 (N_38586,N_34132,N_32149);
nor U38587 (N_38587,N_31594,N_31406);
or U38588 (N_38588,N_31264,N_31891);
or U38589 (N_38589,N_33231,N_33183);
nor U38590 (N_38590,N_34723,N_33378);
nor U38591 (N_38591,N_33059,N_31054);
nand U38592 (N_38592,N_31089,N_33324);
nor U38593 (N_38593,N_32298,N_31188);
and U38594 (N_38594,N_30913,N_32676);
nand U38595 (N_38595,N_31695,N_33639);
nor U38596 (N_38596,N_34640,N_30353);
nand U38597 (N_38597,N_31933,N_33556);
xnor U38598 (N_38598,N_31498,N_34584);
or U38599 (N_38599,N_31318,N_31884);
and U38600 (N_38600,N_31853,N_33793);
xnor U38601 (N_38601,N_32885,N_34086);
or U38602 (N_38602,N_32193,N_31728);
xnor U38603 (N_38603,N_31434,N_32133);
and U38604 (N_38604,N_34659,N_31761);
or U38605 (N_38605,N_34050,N_32419);
nor U38606 (N_38606,N_32827,N_34502);
or U38607 (N_38607,N_33328,N_31399);
xor U38608 (N_38608,N_34860,N_32348);
xor U38609 (N_38609,N_32847,N_34704);
xnor U38610 (N_38610,N_32962,N_33473);
or U38611 (N_38611,N_33304,N_33262);
xnor U38612 (N_38612,N_33732,N_31594);
or U38613 (N_38613,N_33214,N_32409);
nor U38614 (N_38614,N_33096,N_34526);
and U38615 (N_38615,N_32784,N_31626);
or U38616 (N_38616,N_32838,N_30243);
xnor U38617 (N_38617,N_31759,N_32040);
or U38618 (N_38618,N_33563,N_34605);
and U38619 (N_38619,N_32271,N_30542);
xor U38620 (N_38620,N_31025,N_32055);
nor U38621 (N_38621,N_30294,N_32941);
nor U38622 (N_38622,N_32082,N_32690);
nor U38623 (N_38623,N_30719,N_31513);
or U38624 (N_38624,N_32004,N_30355);
or U38625 (N_38625,N_33937,N_32790);
and U38626 (N_38626,N_31899,N_30220);
nor U38627 (N_38627,N_33984,N_34102);
or U38628 (N_38628,N_33714,N_34836);
or U38629 (N_38629,N_33818,N_30338);
nor U38630 (N_38630,N_31788,N_31786);
and U38631 (N_38631,N_30254,N_33566);
xor U38632 (N_38632,N_31656,N_32331);
xnor U38633 (N_38633,N_31948,N_33235);
and U38634 (N_38634,N_31500,N_32280);
or U38635 (N_38635,N_32402,N_31624);
and U38636 (N_38636,N_34119,N_32161);
and U38637 (N_38637,N_30687,N_30579);
and U38638 (N_38638,N_31305,N_33339);
nand U38639 (N_38639,N_32016,N_30498);
nor U38640 (N_38640,N_33046,N_30661);
nor U38641 (N_38641,N_31227,N_33970);
xnor U38642 (N_38642,N_31368,N_34973);
nor U38643 (N_38643,N_31121,N_33676);
nor U38644 (N_38644,N_30934,N_34958);
and U38645 (N_38645,N_32367,N_33310);
xnor U38646 (N_38646,N_33100,N_33972);
nor U38647 (N_38647,N_32647,N_34727);
nand U38648 (N_38648,N_32807,N_31762);
nand U38649 (N_38649,N_34598,N_34698);
or U38650 (N_38650,N_33180,N_30120);
or U38651 (N_38651,N_30552,N_30439);
or U38652 (N_38652,N_30043,N_31027);
nor U38653 (N_38653,N_32762,N_31370);
nor U38654 (N_38654,N_34170,N_32010);
or U38655 (N_38655,N_34232,N_31479);
nor U38656 (N_38656,N_31790,N_32394);
nor U38657 (N_38657,N_30431,N_31667);
xor U38658 (N_38658,N_31764,N_31505);
and U38659 (N_38659,N_34942,N_34479);
nor U38660 (N_38660,N_32260,N_31339);
and U38661 (N_38661,N_34129,N_33357);
or U38662 (N_38662,N_33416,N_32973);
xor U38663 (N_38663,N_31106,N_30247);
nand U38664 (N_38664,N_33282,N_33661);
xnor U38665 (N_38665,N_32675,N_32706);
and U38666 (N_38666,N_34855,N_32484);
nor U38667 (N_38667,N_31994,N_32987);
xnor U38668 (N_38668,N_30933,N_30762);
nand U38669 (N_38669,N_30528,N_34839);
or U38670 (N_38670,N_33343,N_33729);
or U38671 (N_38671,N_33683,N_34647);
or U38672 (N_38672,N_31175,N_32187);
nor U38673 (N_38673,N_34395,N_30770);
or U38674 (N_38674,N_30503,N_34218);
xor U38675 (N_38675,N_33794,N_34795);
xnor U38676 (N_38676,N_32426,N_32282);
or U38677 (N_38677,N_34359,N_34106);
or U38678 (N_38678,N_34283,N_31157);
and U38679 (N_38679,N_33213,N_33491);
xnor U38680 (N_38680,N_32981,N_31203);
or U38681 (N_38681,N_31607,N_30129);
nor U38682 (N_38682,N_31804,N_30173);
xor U38683 (N_38683,N_30461,N_34114);
nor U38684 (N_38684,N_31231,N_30249);
and U38685 (N_38685,N_30412,N_34863);
or U38686 (N_38686,N_32445,N_32605);
and U38687 (N_38687,N_34739,N_34218);
nand U38688 (N_38688,N_33864,N_33086);
xnor U38689 (N_38689,N_30924,N_32101);
nor U38690 (N_38690,N_33998,N_30025);
or U38691 (N_38691,N_34191,N_32651);
nor U38692 (N_38692,N_33900,N_33117);
xnor U38693 (N_38693,N_33012,N_32503);
and U38694 (N_38694,N_33973,N_32897);
and U38695 (N_38695,N_32525,N_33303);
xor U38696 (N_38696,N_30302,N_34382);
or U38697 (N_38697,N_30098,N_34198);
nand U38698 (N_38698,N_30021,N_31062);
nand U38699 (N_38699,N_30019,N_30895);
nor U38700 (N_38700,N_31208,N_34068);
nor U38701 (N_38701,N_34572,N_31753);
xnor U38702 (N_38702,N_30651,N_33921);
or U38703 (N_38703,N_31738,N_30180);
or U38704 (N_38704,N_30101,N_33065);
xor U38705 (N_38705,N_34717,N_31341);
xor U38706 (N_38706,N_30524,N_31731);
nor U38707 (N_38707,N_34862,N_30301);
and U38708 (N_38708,N_33305,N_31475);
nand U38709 (N_38709,N_33095,N_34245);
nand U38710 (N_38710,N_32057,N_34709);
nand U38711 (N_38711,N_34010,N_34955);
and U38712 (N_38712,N_32863,N_30376);
xnor U38713 (N_38713,N_32387,N_30873);
and U38714 (N_38714,N_33122,N_30803);
xor U38715 (N_38715,N_32951,N_33855);
nor U38716 (N_38716,N_34180,N_30393);
nand U38717 (N_38717,N_33025,N_30772);
nand U38718 (N_38718,N_33715,N_33651);
and U38719 (N_38719,N_33156,N_33633);
or U38720 (N_38720,N_33645,N_32717);
or U38721 (N_38721,N_34124,N_32955);
or U38722 (N_38722,N_34974,N_31782);
and U38723 (N_38723,N_34080,N_33631);
or U38724 (N_38724,N_33496,N_33587);
or U38725 (N_38725,N_31379,N_31988);
nand U38726 (N_38726,N_34596,N_30169);
nand U38727 (N_38727,N_32770,N_31013);
nand U38728 (N_38728,N_32297,N_33242);
xnor U38729 (N_38729,N_30526,N_32331);
nor U38730 (N_38730,N_34419,N_31686);
xnor U38731 (N_38731,N_34642,N_32670);
or U38732 (N_38732,N_33073,N_33462);
or U38733 (N_38733,N_32834,N_30679);
or U38734 (N_38734,N_34266,N_30332);
and U38735 (N_38735,N_32150,N_32115);
nor U38736 (N_38736,N_34355,N_31975);
xnor U38737 (N_38737,N_33646,N_32694);
or U38738 (N_38738,N_33860,N_30423);
or U38739 (N_38739,N_32531,N_33390);
nor U38740 (N_38740,N_34640,N_33853);
or U38741 (N_38741,N_32873,N_34047);
and U38742 (N_38742,N_31886,N_30628);
nor U38743 (N_38743,N_34202,N_31372);
nand U38744 (N_38744,N_32273,N_34717);
or U38745 (N_38745,N_32858,N_34102);
xnor U38746 (N_38746,N_33334,N_32522);
or U38747 (N_38747,N_32438,N_33698);
and U38748 (N_38748,N_33292,N_33026);
and U38749 (N_38749,N_30442,N_30271);
nand U38750 (N_38750,N_30628,N_33844);
nor U38751 (N_38751,N_34884,N_33972);
xor U38752 (N_38752,N_32173,N_33217);
and U38753 (N_38753,N_34422,N_33356);
nor U38754 (N_38754,N_33543,N_33157);
nor U38755 (N_38755,N_33157,N_31435);
and U38756 (N_38756,N_32056,N_31928);
xor U38757 (N_38757,N_31990,N_33110);
or U38758 (N_38758,N_30949,N_34987);
nand U38759 (N_38759,N_31430,N_31804);
nand U38760 (N_38760,N_31709,N_31011);
or U38761 (N_38761,N_33635,N_32762);
nand U38762 (N_38762,N_34085,N_32383);
nor U38763 (N_38763,N_33499,N_30947);
nand U38764 (N_38764,N_33645,N_31036);
nor U38765 (N_38765,N_32039,N_32588);
and U38766 (N_38766,N_33557,N_34272);
or U38767 (N_38767,N_31713,N_30976);
or U38768 (N_38768,N_30212,N_32456);
xnor U38769 (N_38769,N_32994,N_34461);
or U38770 (N_38770,N_34334,N_33783);
nor U38771 (N_38771,N_32030,N_33170);
nor U38772 (N_38772,N_32697,N_31923);
nor U38773 (N_38773,N_31229,N_32319);
or U38774 (N_38774,N_32988,N_33972);
nand U38775 (N_38775,N_34399,N_33887);
and U38776 (N_38776,N_32032,N_33813);
and U38777 (N_38777,N_30037,N_32534);
and U38778 (N_38778,N_34451,N_33568);
nor U38779 (N_38779,N_33705,N_32249);
nor U38780 (N_38780,N_30617,N_31877);
and U38781 (N_38781,N_33621,N_31685);
and U38782 (N_38782,N_31103,N_34445);
and U38783 (N_38783,N_32903,N_32233);
nand U38784 (N_38784,N_30797,N_33360);
nor U38785 (N_38785,N_30614,N_34468);
xnor U38786 (N_38786,N_33309,N_30445);
nand U38787 (N_38787,N_31387,N_31325);
xor U38788 (N_38788,N_34461,N_31953);
or U38789 (N_38789,N_30887,N_32154);
nand U38790 (N_38790,N_32093,N_32009);
nand U38791 (N_38791,N_32712,N_32768);
xnor U38792 (N_38792,N_32430,N_31074);
xor U38793 (N_38793,N_33056,N_34308);
nand U38794 (N_38794,N_32675,N_32143);
or U38795 (N_38795,N_34830,N_30079);
xnor U38796 (N_38796,N_32170,N_33907);
nand U38797 (N_38797,N_30011,N_33051);
and U38798 (N_38798,N_32592,N_30477);
nand U38799 (N_38799,N_34479,N_32214);
nor U38800 (N_38800,N_33961,N_31531);
or U38801 (N_38801,N_32354,N_31795);
nor U38802 (N_38802,N_34685,N_32534);
nor U38803 (N_38803,N_32323,N_31049);
or U38804 (N_38804,N_34560,N_34459);
xnor U38805 (N_38805,N_33297,N_34530);
and U38806 (N_38806,N_34215,N_31798);
xor U38807 (N_38807,N_30519,N_32500);
xor U38808 (N_38808,N_30317,N_32722);
and U38809 (N_38809,N_34456,N_34233);
or U38810 (N_38810,N_33829,N_30507);
xor U38811 (N_38811,N_32584,N_34153);
and U38812 (N_38812,N_30254,N_33791);
and U38813 (N_38813,N_30575,N_33020);
or U38814 (N_38814,N_33532,N_31544);
nand U38815 (N_38815,N_33650,N_31174);
nor U38816 (N_38816,N_30522,N_31992);
nor U38817 (N_38817,N_34106,N_33068);
and U38818 (N_38818,N_32265,N_34015);
or U38819 (N_38819,N_32032,N_31375);
nand U38820 (N_38820,N_33120,N_32027);
and U38821 (N_38821,N_32230,N_32362);
nor U38822 (N_38822,N_33767,N_32898);
and U38823 (N_38823,N_30869,N_31464);
nand U38824 (N_38824,N_30367,N_34818);
nand U38825 (N_38825,N_33442,N_30660);
nor U38826 (N_38826,N_32908,N_31374);
xor U38827 (N_38827,N_31348,N_32889);
or U38828 (N_38828,N_33038,N_30922);
xnor U38829 (N_38829,N_34238,N_34846);
xor U38830 (N_38830,N_31934,N_33991);
xor U38831 (N_38831,N_33927,N_30417);
or U38832 (N_38832,N_34352,N_30755);
or U38833 (N_38833,N_31159,N_34538);
and U38834 (N_38834,N_34533,N_30415);
nor U38835 (N_38835,N_34522,N_30995);
nor U38836 (N_38836,N_31538,N_33635);
and U38837 (N_38837,N_30382,N_34619);
xor U38838 (N_38838,N_34787,N_33530);
xnor U38839 (N_38839,N_30286,N_32545);
nand U38840 (N_38840,N_34097,N_32198);
nand U38841 (N_38841,N_30142,N_30320);
nor U38842 (N_38842,N_31680,N_32129);
or U38843 (N_38843,N_34558,N_34725);
and U38844 (N_38844,N_30214,N_33875);
and U38845 (N_38845,N_31298,N_34582);
xnor U38846 (N_38846,N_34750,N_33363);
xnor U38847 (N_38847,N_31270,N_33322);
or U38848 (N_38848,N_31487,N_30496);
or U38849 (N_38849,N_31238,N_32356);
nor U38850 (N_38850,N_31344,N_30643);
nand U38851 (N_38851,N_32844,N_30589);
or U38852 (N_38852,N_30720,N_30602);
xnor U38853 (N_38853,N_33772,N_33187);
nand U38854 (N_38854,N_32398,N_34945);
nor U38855 (N_38855,N_33867,N_32833);
or U38856 (N_38856,N_33380,N_31869);
nor U38857 (N_38857,N_31673,N_31946);
nand U38858 (N_38858,N_30479,N_31934);
nand U38859 (N_38859,N_33510,N_31122);
or U38860 (N_38860,N_34552,N_31351);
nand U38861 (N_38861,N_31894,N_31830);
xnor U38862 (N_38862,N_31570,N_31301);
nand U38863 (N_38863,N_30238,N_34956);
or U38864 (N_38864,N_34986,N_33470);
nand U38865 (N_38865,N_33013,N_30069);
nor U38866 (N_38866,N_30916,N_31309);
nand U38867 (N_38867,N_33838,N_30313);
and U38868 (N_38868,N_33895,N_31278);
nor U38869 (N_38869,N_34090,N_33353);
and U38870 (N_38870,N_34138,N_33992);
and U38871 (N_38871,N_34236,N_30996);
or U38872 (N_38872,N_34739,N_32862);
nand U38873 (N_38873,N_32401,N_30478);
nand U38874 (N_38874,N_32341,N_33381);
and U38875 (N_38875,N_30037,N_33606);
and U38876 (N_38876,N_33527,N_34949);
nor U38877 (N_38877,N_30245,N_32817);
nor U38878 (N_38878,N_34786,N_32147);
nand U38879 (N_38879,N_31091,N_34985);
and U38880 (N_38880,N_32703,N_33158);
nor U38881 (N_38881,N_33727,N_34838);
nor U38882 (N_38882,N_33071,N_30254);
xnor U38883 (N_38883,N_34356,N_30521);
or U38884 (N_38884,N_34681,N_32194);
xnor U38885 (N_38885,N_31196,N_31393);
and U38886 (N_38886,N_33558,N_32679);
nand U38887 (N_38887,N_31456,N_31754);
nor U38888 (N_38888,N_30530,N_34259);
xnor U38889 (N_38889,N_32082,N_32689);
nor U38890 (N_38890,N_33723,N_34562);
or U38891 (N_38891,N_32985,N_30462);
xor U38892 (N_38892,N_32631,N_34596);
nor U38893 (N_38893,N_33409,N_33656);
nand U38894 (N_38894,N_30770,N_30364);
and U38895 (N_38895,N_31707,N_33590);
or U38896 (N_38896,N_33050,N_31012);
xnor U38897 (N_38897,N_30662,N_34613);
or U38898 (N_38898,N_34725,N_31212);
nand U38899 (N_38899,N_33765,N_33707);
nor U38900 (N_38900,N_30668,N_30586);
or U38901 (N_38901,N_34128,N_34111);
xnor U38902 (N_38902,N_30513,N_32971);
xor U38903 (N_38903,N_33415,N_31949);
and U38904 (N_38904,N_32814,N_31435);
and U38905 (N_38905,N_31634,N_32885);
nor U38906 (N_38906,N_34202,N_30152);
xnor U38907 (N_38907,N_31248,N_32826);
or U38908 (N_38908,N_30971,N_30429);
nand U38909 (N_38909,N_32784,N_30623);
nor U38910 (N_38910,N_33135,N_33134);
nand U38911 (N_38911,N_33662,N_32257);
or U38912 (N_38912,N_32602,N_30029);
or U38913 (N_38913,N_33705,N_32893);
or U38914 (N_38914,N_31705,N_30076);
xor U38915 (N_38915,N_33139,N_34170);
or U38916 (N_38916,N_31265,N_31870);
or U38917 (N_38917,N_34538,N_32372);
nor U38918 (N_38918,N_32828,N_31291);
xnor U38919 (N_38919,N_30419,N_32913);
nor U38920 (N_38920,N_32206,N_30492);
nor U38921 (N_38921,N_30925,N_32026);
and U38922 (N_38922,N_33423,N_31814);
and U38923 (N_38923,N_34150,N_30623);
nor U38924 (N_38924,N_30684,N_31334);
or U38925 (N_38925,N_33761,N_33175);
nor U38926 (N_38926,N_32336,N_31510);
nor U38927 (N_38927,N_33118,N_34435);
nand U38928 (N_38928,N_30851,N_32674);
nor U38929 (N_38929,N_33232,N_34114);
or U38930 (N_38930,N_30336,N_33982);
and U38931 (N_38931,N_34665,N_30790);
nor U38932 (N_38932,N_31698,N_33043);
and U38933 (N_38933,N_31328,N_33558);
nor U38934 (N_38934,N_33268,N_32420);
xor U38935 (N_38935,N_33826,N_32766);
and U38936 (N_38936,N_30785,N_33379);
xnor U38937 (N_38937,N_34290,N_33663);
xor U38938 (N_38938,N_34093,N_33982);
xor U38939 (N_38939,N_31245,N_30056);
or U38940 (N_38940,N_31977,N_31533);
or U38941 (N_38941,N_30542,N_32421);
or U38942 (N_38942,N_33314,N_31626);
and U38943 (N_38943,N_30747,N_32654);
and U38944 (N_38944,N_32817,N_33758);
nor U38945 (N_38945,N_34640,N_34626);
and U38946 (N_38946,N_31294,N_32964);
or U38947 (N_38947,N_34733,N_34313);
nand U38948 (N_38948,N_34798,N_32612);
or U38949 (N_38949,N_33748,N_30493);
and U38950 (N_38950,N_34536,N_33077);
nand U38951 (N_38951,N_30741,N_30222);
or U38952 (N_38952,N_33959,N_30072);
nor U38953 (N_38953,N_30819,N_30497);
or U38954 (N_38954,N_31931,N_33463);
nand U38955 (N_38955,N_31839,N_34415);
and U38956 (N_38956,N_34359,N_34620);
nor U38957 (N_38957,N_31970,N_33104);
or U38958 (N_38958,N_34548,N_33653);
or U38959 (N_38959,N_33962,N_31993);
nor U38960 (N_38960,N_34032,N_30627);
xnor U38961 (N_38961,N_31428,N_32596);
xnor U38962 (N_38962,N_33448,N_31649);
xor U38963 (N_38963,N_34781,N_31819);
nor U38964 (N_38964,N_32861,N_31634);
xor U38965 (N_38965,N_31846,N_34423);
nand U38966 (N_38966,N_32316,N_33713);
or U38967 (N_38967,N_30501,N_33624);
nand U38968 (N_38968,N_31398,N_31062);
or U38969 (N_38969,N_31628,N_30534);
and U38970 (N_38970,N_31181,N_31230);
xnor U38971 (N_38971,N_31395,N_31572);
and U38972 (N_38972,N_32731,N_34199);
and U38973 (N_38973,N_33416,N_30326);
and U38974 (N_38974,N_30748,N_34012);
and U38975 (N_38975,N_33875,N_31829);
xnor U38976 (N_38976,N_31057,N_30127);
nor U38977 (N_38977,N_30490,N_30908);
or U38978 (N_38978,N_32711,N_31227);
xor U38979 (N_38979,N_32921,N_33718);
nor U38980 (N_38980,N_34693,N_33049);
and U38981 (N_38981,N_32196,N_33892);
nand U38982 (N_38982,N_30403,N_33362);
nor U38983 (N_38983,N_34927,N_30387);
nand U38984 (N_38984,N_33041,N_32079);
and U38985 (N_38985,N_30067,N_32512);
and U38986 (N_38986,N_32768,N_30204);
nand U38987 (N_38987,N_32251,N_31388);
and U38988 (N_38988,N_34229,N_34692);
nand U38989 (N_38989,N_32185,N_32727);
xnor U38990 (N_38990,N_33592,N_34062);
nor U38991 (N_38991,N_33968,N_31721);
nand U38992 (N_38992,N_33463,N_31139);
or U38993 (N_38993,N_33203,N_32542);
or U38994 (N_38994,N_33793,N_32598);
xor U38995 (N_38995,N_33092,N_32591);
or U38996 (N_38996,N_30884,N_31409);
xnor U38997 (N_38997,N_30252,N_32750);
and U38998 (N_38998,N_33019,N_34702);
or U38999 (N_38999,N_30951,N_33230);
and U39000 (N_39000,N_34725,N_33219);
xnor U39001 (N_39001,N_31068,N_31349);
or U39002 (N_39002,N_31658,N_32406);
nor U39003 (N_39003,N_31944,N_31741);
and U39004 (N_39004,N_33683,N_31714);
or U39005 (N_39005,N_33231,N_34307);
or U39006 (N_39006,N_32660,N_31406);
nor U39007 (N_39007,N_31093,N_32210);
and U39008 (N_39008,N_34110,N_30819);
or U39009 (N_39009,N_34112,N_30243);
nand U39010 (N_39010,N_32675,N_33306);
nor U39011 (N_39011,N_31927,N_32728);
and U39012 (N_39012,N_34192,N_32744);
xor U39013 (N_39013,N_31895,N_32641);
nor U39014 (N_39014,N_31452,N_31786);
nand U39015 (N_39015,N_33359,N_30891);
nand U39016 (N_39016,N_33401,N_30985);
and U39017 (N_39017,N_32754,N_30013);
nand U39018 (N_39018,N_34362,N_33052);
nor U39019 (N_39019,N_31141,N_30815);
xnor U39020 (N_39020,N_32724,N_34174);
or U39021 (N_39021,N_32466,N_31263);
nand U39022 (N_39022,N_30897,N_32127);
or U39023 (N_39023,N_33833,N_31905);
and U39024 (N_39024,N_34731,N_30838);
nand U39025 (N_39025,N_32815,N_32049);
nand U39026 (N_39026,N_32251,N_31072);
nor U39027 (N_39027,N_32046,N_30858);
and U39028 (N_39028,N_30453,N_34359);
or U39029 (N_39029,N_33512,N_32305);
xor U39030 (N_39030,N_33031,N_33982);
and U39031 (N_39031,N_33743,N_30020);
and U39032 (N_39032,N_34868,N_30850);
nand U39033 (N_39033,N_34301,N_34012);
nand U39034 (N_39034,N_33597,N_32431);
or U39035 (N_39035,N_34162,N_34707);
xnor U39036 (N_39036,N_31159,N_32457);
nor U39037 (N_39037,N_34630,N_33289);
and U39038 (N_39038,N_34857,N_30816);
nor U39039 (N_39039,N_33532,N_33023);
and U39040 (N_39040,N_32953,N_34730);
nand U39041 (N_39041,N_32815,N_34578);
or U39042 (N_39042,N_31849,N_32191);
and U39043 (N_39043,N_30247,N_31320);
and U39044 (N_39044,N_30634,N_30462);
xnor U39045 (N_39045,N_31564,N_32056);
xor U39046 (N_39046,N_32625,N_34224);
or U39047 (N_39047,N_33335,N_34833);
xor U39048 (N_39048,N_30912,N_31223);
or U39049 (N_39049,N_32553,N_30059);
xnor U39050 (N_39050,N_30057,N_32494);
or U39051 (N_39051,N_30672,N_30994);
or U39052 (N_39052,N_33868,N_33066);
and U39053 (N_39053,N_31130,N_34386);
nand U39054 (N_39054,N_33479,N_34592);
nand U39055 (N_39055,N_31611,N_31966);
and U39056 (N_39056,N_33815,N_30445);
nand U39057 (N_39057,N_32592,N_34738);
and U39058 (N_39058,N_30938,N_30011);
nor U39059 (N_39059,N_34162,N_31938);
nor U39060 (N_39060,N_30652,N_34356);
nand U39061 (N_39061,N_30028,N_34865);
nand U39062 (N_39062,N_32559,N_34810);
or U39063 (N_39063,N_30546,N_32722);
or U39064 (N_39064,N_34668,N_31600);
and U39065 (N_39065,N_32837,N_33788);
or U39066 (N_39066,N_34005,N_33214);
nand U39067 (N_39067,N_34038,N_30221);
and U39068 (N_39068,N_31178,N_31885);
or U39069 (N_39069,N_33861,N_33709);
or U39070 (N_39070,N_34818,N_31587);
nor U39071 (N_39071,N_33899,N_34517);
and U39072 (N_39072,N_34552,N_33880);
xor U39073 (N_39073,N_31068,N_31563);
nor U39074 (N_39074,N_30684,N_32231);
nand U39075 (N_39075,N_33890,N_30794);
nor U39076 (N_39076,N_31430,N_31087);
and U39077 (N_39077,N_31952,N_31794);
nor U39078 (N_39078,N_34330,N_33647);
and U39079 (N_39079,N_34800,N_32284);
xor U39080 (N_39080,N_34592,N_30544);
nor U39081 (N_39081,N_34312,N_30921);
and U39082 (N_39082,N_31702,N_33584);
and U39083 (N_39083,N_32402,N_34662);
xor U39084 (N_39084,N_32733,N_33757);
or U39085 (N_39085,N_33223,N_34660);
nor U39086 (N_39086,N_31346,N_30325);
and U39087 (N_39087,N_30466,N_32125);
and U39088 (N_39088,N_33253,N_34389);
nor U39089 (N_39089,N_34421,N_32616);
or U39090 (N_39090,N_32303,N_30725);
nand U39091 (N_39091,N_30795,N_30504);
nand U39092 (N_39092,N_31947,N_31910);
and U39093 (N_39093,N_31026,N_34741);
nand U39094 (N_39094,N_30104,N_33955);
nor U39095 (N_39095,N_30451,N_30055);
and U39096 (N_39096,N_31325,N_31688);
or U39097 (N_39097,N_34313,N_34156);
and U39098 (N_39098,N_31544,N_34708);
or U39099 (N_39099,N_34342,N_34513);
or U39100 (N_39100,N_31477,N_32291);
nor U39101 (N_39101,N_30528,N_32177);
and U39102 (N_39102,N_32309,N_32127);
or U39103 (N_39103,N_32752,N_32461);
nor U39104 (N_39104,N_33006,N_32255);
nor U39105 (N_39105,N_30941,N_34226);
and U39106 (N_39106,N_33256,N_30983);
and U39107 (N_39107,N_30881,N_30182);
and U39108 (N_39108,N_32667,N_30226);
and U39109 (N_39109,N_34217,N_33485);
xor U39110 (N_39110,N_32597,N_33177);
and U39111 (N_39111,N_30788,N_31257);
nor U39112 (N_39112,N_32537,N_31246);
nor U39113 (N_39113,N_34296,N_30262);
nand U39114 (N_39114,N_33963,N_30455);
nor U39115 (N_39115,N_33358,N_34735);
and U39116 (N_39116,N_32311,N_31868);
and U39117 (N_39117,N_30287,N_31260);
xor U39118 (N_39118,N_31372,N_30633);
nor U39119 (N_39119,N_32422,N_33626);
or U39120 (N_39120,N_30303,N_31597);
xnor U39121 (N_39121,N_33881,N_34460);
nand U39122 (N_39122,N_33191,N_31772);
nand U39123 (N_39123,N_33727,N_34862);
nor U39124 (N_39124,N_30615,N_32325);
nor U39125 (N_39125,N_30309,N_32793);
or U39126 (N_39126,N_32839,N_33333);
nand U39127 (N_39127,N_34728,N_34260);
nor U39128 (N_39128,N_30648,N_30589);
nand U39129 (N_39129,N_32790,N_30735);
or U39130 (N_39130,N_33118,N_34313);
nor U39131 (N_39131,N_31661,N_32177);
or U39132 (N_39132,N_33302,N_34802);
nand U39133 (N_39133,N_30304,N_33029);
nand U39134 (N_39134,N_33453,N_32494);
xnor U39135 (N_39135,N_30224,N_33712);
or U39136 (N_39136,N_34666,N_33984);
nand U39137 (N_39137,N_32382,N_32059);
xnor U39138 (N_39138,N_31791,N_30566);
or U39139 (N_39139,N_30353,N_33253);
nor U39140 (N_39140,N_34790,N_32057);
or U39141 (N_39141,N_33416,N_32451);
and U39142 (N_39142,N_32513,N_32730);
nor U39143 (N_39143,N_34977,N_33560);
nor U39144 (N_39144,N_34113,N_33067);
nand U39145 (N_39145,N_34437,N_33275);
xnor U39146 (N_39146,N_32934,N_33552);
xor U39147 (N_39147,N_33095,N_30909);
or U39148 (N_39148,N_31741,N_32707);
xnor U39149 (N_39149,N_31421,N_33068);
nor U39150 (N_39150,N_32545,N_34153);
xnor U39151 (N_39151,N_30774,N_33390);
or U39152 (N_39152,N_31030,N_31393);
and U39153 (N_39153,N_30895,N_32796);
nand U39154 (N_39154,N_33942,N_34140);
xnor U39155 (N_39155,N_33549,N_30627);
nor U39156 (N_39156,N_30672,N_32882);
and U39157 (N_39157,N_32897,N_32485);
or U39158 (N_39158,N_31058,N_30299);
or U39159 (N_39159,N_30237,N_33009);
xor U39160 (N_39160,N_31396,N_34800);
nor U39161 (N_39161,N_31166,N_32574);
and U39162 (N_39162,N_34674,N_30710);
nor U39163 (N_39163,N_32876,N_30191);
or U39164 (N_39164,N_31828,N_31385);
xnor U39165 (N_39165,N_30679,N_32999);
xnor U39166 (N_39166,N_34236,N_30019);
nor U39167 (N_39167,N_33287,N_31505);
and U39168 (N_39168,N_30565,N_31625);
xnor U39169 (N_39169,N_32763,N_30576);
xor U39170 (N_39170,N_31593,N_31380);
xor U39171 (N_39171,N_33059,N_32945);
nand U39172 (N_39172,N_32039,N_33191);
nor U39173 (N_39173,N_31194,N_34170);
or U39174 (N_39174,N_34295,N_30749);
nand U39175 (N_39175,N_32880,N_33115);
and U39176 (N_39176,N_33446,N_31729);
xnor U39177 (N_39177,N_33412,N_33781);
and U39178 (N_39178,N_34835,N_32198);
or U39179 (N_39179,N_32036,N_32482);
nand U39180 (N_39180,N_31551,N_32406);
or U39181 (N_39181,N_32303,N_31545);
and U39182 (N_39182,N_34557,N_33267);
xnor U39183 (N_39183,N_33990,N_32933);
nor U39184 (N_39184,N_32672,N_32739);
nor U39185 (N_39185,N_30599,N_34592);
nand U39186 (N_39186,N_30197,N_34117);
or U39187 (N_39187,N_32335,N_31494);
nand U39188 (N_39188,N_32093,N_34277);
or U39189 (N_39189,N_32786,N_33897);
nand U39190 (N_39190,N_34338,N_31001);
nor U39191 (N_39191,N_34247,N_30033);
or U39192 (N_39192,N_33302,N_33136);
xor U39193 (N_39193,N_34542,N_30520);
nand U39194 (N_39194,N_33698,N_33176);
nand U39195 (N_39195,N_34459,N_33455);
and U39196 (N_39196,N_31677,N_31736);
xor U39197 (N_39197,N_33049,N_30437);
xnor U39198 (N_39198,N_32307,N_32241);
nor U39199 (N_39199,N_31839,N_34839);
or U39200 (N_39200,N_30557,N_30015);
nand U39201 (N_39201,N_30838,N_32635);
nand U39202 (N_39202,N_33551,N_33706);
and U39203 (N_39203,N_33163,N_30714);
xor U39204 (N_39204,N_33200,N_30531);
nor U39205 (N_39205,N_33270,N_32116);
nor U39206 (N_39206,N_32973,N_32833);
xor U39207 (N_39207,N_30979,N_33270);
or U39208 (N_39208,N_34089,N_31652);
or U39209 (N_39209,N_30999,N_31095);
nand U39210 (N_39210,N_30529,N_30266);
or U39211 (N_39211,N_33751,N_33295);
and U39212 (N_39212,N_33907,N_33381);
or U39213 (N_39213,N_33335,N_30116);
nand U39214 (N_39214,N_31710,N_32980);
nand U39215 (N_39215,N_33105,N_30360);
nor U39216 (N_39216,N_33990,N_32173);
and U39217 (N_39217,N_31291,N_33902);
and U39218 (N_39218,N_31109,N_33582);
and U39219 (N_39219,N_34777,N_30225);
and U39220 (N_39220,N_32460,N_31465);
nor U39221 (N_39221,N_33105,N_32664);
nor U39222 (N_39222,N_31250,N_31356);
and U39223 (N_39223,N_33000,N_34773);
or U39224 (N_39224,N_33375,N_31035);
or U39225 (N_39225,N_34209,N_30569);
or U39226 (N_39226,N_34911,N_33182);
xor U39227 (N_39227,N_34347,N_34944);
or U39228 (N_39228,N_33484,N_31994);
nand U39229 (N_39229,N_33103,N_31544);
xnor U39230 (N_39230,N_30861,N_30765);
xor U39231 (N_39231,N_30209,N_34907);
and U39232 (N_39232,N_33430,N_32125);
or U39233 (N_39233,N_33576,N_34980);
nand U39234 (N_39234,N_31287,N_30658);
nor U39235 (N_39235,N_30257,N_32053);
nor U39236 (N_39236,N_33404,N_30742);
nand U39237 (N_39237,N_34038,N_34926);
nand U39238 (N_39238,N_32263,N_32176);
xor U39239 (N_39239,N_30138,N_30998);
and U39240 (N_39240,N_34681,N_34240);
or U39241 (N_39241,N_33962,N_31307);
or U39242 (N_39242,N_31038,N_34600);
nand U39243 (N_39243,N_31275,N_30496);
and U39244 (N_39244,N_33057,N_30585);
or U39245 (N_39245,N_32833,N_30730);
and U39246 (N_39246,N_30813,N_30934);
nand U39247 (N_39247,N_30488,N_31191);
nor U39248 (N_39248,N_30252,N_31567);
xnor U39249 (N_39249,N_33098,N_31782);
nand U39250 (N_39250,N_31641,N_33792);
or U39251 (N_39251,N_32737,N_33899);
xnor U39252 (N_39252,N_33679,N_34290);
nand U39253 (N_39253,N_31801,N_34432);
and U39254 (N_39254,N_31957,N_31774);
and U39255 (N_39255,N_30569,N_31302);
xor U39256 (N_39256,N_30235,N_33312);
xor U39257 (N_39257,N_34994,N_33117);
xnor U39258 (N_39258,N_31809,N_33550);
nor U39259 (N_39259,N_34291,N_30070);
nand U39260 (N_39260,N_32897,N_31990);
and U39261 (N_39261,N_31690,N_34203);
nand U39262 (N_39262,N_33102,N_32551);
or U39263 (N_39263,N_31646,N_33027);
xor U39264 (N_39264,N_31568,N_33328);
nor U39265 (N_39265,N_32680,N_34332);
or U39266 (N_39266,N_34869,N_31245);
xor U39267 (N_39267,N_31073,N_32046);
or U39268 (N_39268,N_30426,N_34448);
nor U39269 (N_39269,N_31122,N_33842);
nand U39270 (N_39270,N_33121,N_30225);
nand U39271 (N_39271,N_31958,N_31764);
nand U39272 (N_39272,N_32236,N_33490);
xor U39273 (N_39273,N_32221,N_33780);
and U39274 (N_39274,N_34536,N_34133);
nor U39275 (N_39275,N_33219,N_31254);
or U39276 (N_39276,N_34667,N_32853);
xnor U39277 (N_39277,N_32885,N_34101);
and U39278 (N_39278,N_31552,N_32764);
and U39279 (N_39279,N_33325,N_34150);
xor U39280 (N_39280,N_30796,N_31750);
and U39281 (N_39281,N_30121,N_30390);
nor U39282 (N_39282,N_31061,N_32077);
and U39283 (N_39283,N_34313,N_34284);
and U39284 (N_39284,N_30556,N_30500);
xor U39285 (N_39285,N_31760,N_34450);
xor U39286 (N_39286,N_33840,N_34043);
nor U39287 (N_39287,N_34056,N_31424);
and U39288 (N_39288,N_34923,N_30644);
nand U39289 (N_39289,N_34809,N_33736);
nor U39290 (N_39290,N_33442,N_33622);
xnor U39291 (N_39291,N_30300,N_32058);
nor U39292 (N_39292,N_34997,N_31690);
and U39293 (N_39293,N_32414,N_34192);
nor U39294 (N_39294,N_30263,N_33562);
nand U39295 (N_39295,N_33515,N_32522);
nor U39296 (N_39296,N_31645,N_32986);
xor U39297 (N_39297,N_33452,N_32218);
or U39298 (N_39298,N_33078,N_30027);
xnor U39299 (N_39299,N_32203,N_31097);
xnor U39300 (N_39300,N_34919,N_33138);
nand U39301 (N_39301,N_30323,N_34369);
nand U39302 (N_39302,N_34421,N_33513);
or U39303 (N_39303,N_33753,N_34727);
nor U39304 (N_39304,N_34186,N_32413);
xnor U39305 (N_39305,N_32228,N_33143);
nand U39306 (N_39306,N_31253,N_31828);
and U39307 (N_39307,N_30457,N_32270);
or U39308 (N_39308,N_33743,N_30436);
or U39309 (N_39309,N_32266,N_31063);
or U39310 (N_39310,N_34152,N_32233);
nor U39311 (N_39311,N_32995,N_30265);
nand U39312 (N_39312,N_31824,N_32406);
nor U39313 (N_39313,N_31415,N_32256);
nor U39314 (N_39314,N_32946,N_30592);
or U39315 (N_39315,N_34796,N_32565);
nor U39316 (N_39316,N_32479,N_33649);
xnor U39317 (N_39317,N_33869,N_32808);
or U39318 (N_39318,N_34987,N_33188);
xnor U39319 (N_39319,N_32583,N_34766);
or U39320 (N_39320,N_30611,N_34927);
nand U39321 (N_39321,N_33874,N_31711);
or U39322 (N_39322,N_33462,N_33790);
xnor U39323 (N_39323,N_31763,N_33478);
or U39324 (N_39324,N_34340,N_32891);
or U39325 (N_39325,N_31648,N_31617);
xnor U39326 (N_39326,N_31036,N_30724);
nand U39327 (N_39327,N_32597,N_32478);
nor U39328 (N_39328,N_34581,N_32334);
xor U39329 (N_39329,N_31481,N_32495);
or U39330 (N_39330,N_31580,N_34196);
and U39331 (N_39331,N_32128,N_32987);
xor U39332 (N_39332,N_32635,N_32037);
nor U39333 (N_39333,N_31413,N_34371);
and U39334 (N_39334,N_30432,N_34620);
nor U39335 (N_39335,N_33683,N_34218);
nor U39336 (N_39336,N_32528,N_34156);
nor U39337 (N_39337,N_31295,N_34311);
nor U39338 (N_39338,N_30694,N_33192);
or U39339 (N_39339,N_30339,N_32724);
xor U39340 (N_39340,N_32840,N_30448);
xor U39341 (N_39341,N_32092,N_34299);
nand U39342 (N_39342,N_31099,N_30235);
or U39343 (N_39343,N_31595,N_32087);
nand U39344 (N_39344,N_31388,N_34318);
nand U39345 (N_39345,N_31259,N_32744);
and U39346 (N_39346,N_33494,N_32734);
or U39347 (N_39347,N_30667,N_31862);
xnor U39348 (N_39348,N_33637,N_34950);
nor U39349 (N_39349,N_33582,N_32036);
and U39350 (N_39350,N_30210,N_34839);
and U39351 (N_39351,N_34806,N_33370);
and U39352 (N_39352,N_31702,N_32739);
xnor U39353 (N_39353,N_30645,N_32534);
xnor U39354 (N_39354,N_31732,N_33709);
nor U39355 (N_39355,N_31486,N_33790);
xnor U39356 (N_39356,N_34846,N_33199);
nand U39357 (N_39357,N_31752,N_33414);
or U39358 (N_39358,N_30562,N_32605);
xor U39359 (N_39359,N_32092,N_32606);
or U39360 (N_39360,N_33435,N_31767);
or U39361 (N_39361,N_32782,N_30650);
nor U39362 (N_39362,N_32212,N_34802);
nor U39363 (N_39363,N_30609,N_33359);
or U39364 (N_39364,N_30229,N_32408);
nand U39365 (N_39365,N_33597,N_34280);
nand U39366 (N_39366,N_30535,N_30681);
xnor U39367 (N_39367,N_34281,N_34295);
xor U39368 (N_39368,N_32733,N_30568);
or U39369 (N_39369,N_32845,N_34986);
and U39370 (N_39370,N_34052,N_33835);
nor U39371 (N_39371,N_31613,N_33172);
xnor U39372 (N_39372,N_33133,N_33978);
or U39373 (N_39373,N_31056,N_31551);
nand U39374 (N_39374,N_31159,N_34050);
nor U39375 (N_39375,N_31590,N_32148);
nor U39376 (N_39376,N_31101,N_30127);
nand U39377 (N_39377,N_33372,N_30895);
xor U39378 (N_39378,N_30304,N_32670);
nor U39379 (N_39379,N_32930,N_30451);
nor U39380 (N_39380,N_30930,N_34026);
xnor U39381 (N_39381,N_30307,N_30057);
nor U39382 (N_39382,N_32000,N_30663);
and U39383 (N_39383,N_34174,N_31914);
xnor U39384 (N_39384,N_34454,N_33994);
or U39385 (N_39385,N_31829,N_31801);
and U39386 (N_39386,N_31963,N_30530);
xnor U39387 (N_39387,N_33305,N_30298);
xor U39388 (N_39388,N_31308,N_31358);
and U39389 (N_39389,N_31491,N_34671);
xnor U39390 (N_39390,N_31274,N_34270);
and U39391 (N_39391,N_30623,N_34008);
nor U39392 (N_39392,N_31392,N_32990);
or U39393 (N_39393,N_31745,N_33120);
nor U39394 (N_39394,N_31049,N_32576);
and U39395 (N_39395,N_32544,N_32611);
nand U39396 (N_39396,N_30897,N_34165);
or U39397 (N_39397,N_30416,N_33902);
nand U39398 (N_39398,N_31644,N_32843);
or U39399 (N_39399,N_34879,N_32451);
nand U39400 (N_39400,N_33961,N_32451);
xor U39401 (N_39401,N_32061,N_34658);
or U39402 (N_39402,N_33581,N_31474);
nand U39403 (N_39403,N_34894,N_31038);
xnor U39404 (N_39404,N_32070,N_30357);
nor U39405 (N_39405,N_33967,N_31528);
xnor U39406 (N_39406,N_31102,N_34747);
nor U39407 (N_39407,N_30614,N_32229);
or U39408 (N_39408,N_31344,N_33225);
and U39409 (N_39409,N_32032,N_30866);
and U39410 (N_39410,N_31874,N_31841);
nand U39411 (N_39411,N_30905,N_33918);
xnor U39412 (N_39412,N_33190,N_32866);
and U39413 (N_39413,N_30416,N_32555);
nand U39414 (N_39414,N_34892,N_30548);
nand U39415 (N_39415,N_32426,N_32457);
xnor U39416 (N_39416,N_32451,N_30986);
nand U39417 (N_39417,N_33664,N_31733);
xor U39418 (N_39418,N_33813,N_31595);
nand U39419 (N_39419,N_30366,N_34439);
nand U39420 (N_39420,N_32205,N_32276);
nand U39421 (N_39421,N_33317,N_33357);
nand U39422 (N_39422,N_32116,N_33354);
or U39423 (N_39423,N_33454,N_30766);
nand U39424 (N_39424,N_34221,N_30951);
nand U39425 (N_39425,N_32299,N_30185);
or U39426 (N_39426,N_31628,N_31127);
nand U39427 (N_39427,N_34226,N_30811);
xnor U39428 (N_39428,N_30901,N_33908);
xor U39429 (N_39429,N_32874,N_30138);
or U39430 (N_39430,N_33341,N_31441);
nand U39431 (N_39431,N_34240,N_31977);
nand U39432 (N_39432,N_30667,N_31670);
nand U39433 (N_39433,N_34370,N_30106);
nand U39434 (N_39434,N_32937,N_30975);
and U39435 (N_39435,N_32588,N_33300);
and U39436 (N_39436,N_33422,N_31120);
and U39437 (N_39437,N_34152,N_31698);
nand U39438 (N_39438,N_31265,N_30228);
nor U39439 (N_39439,N_30626,N_30936);
or U39440 (N_39440,N_33532,N_33514);
nor U39441 (N_39441,N_32187,N_32147);
or U39442 (N_39442,N_30358,N_32213);
and U39443 (N_39443,N_34381,N_33281);
or U39444 (N_39444,N_31661,N_34022);
and U39445 (N_39445,N_33745,N_30268);
or U39446 (N_39446,N_31728,N_32911);
and U39447 (N_39447,N_34593,N_34691);
nor U39448 (N_39448,N_34663,N_32896);
or U39449 (N_39449,N_34706,N_31815);
nor U39450 (N_39450,N_31023,N_31212);
xnor U39451 (N_39451,N_30055,N_31036);
xnor U39452 (N_39452,N_34657,N_32605);
nor U39453 (N_39453,N_31980,N_32295);
and U39454 (N_39454,N_32524,N_33614);
xor U39455 (N_39455,N_31052,N_33339);
or U39456 (N_39456,N_32430,N_34055);
nand U39457 (N_39457,N_34180,N_32152);
nand U39458 (N_39458,N_32276,N_32734);
nand U39459 (N_39459,N_34190,N_33056);
and U39460 (N_39460,N_34968,N_30250);
and U39461 (N_39461,N_34251,N_34804);
xnor U39462 (N_39462,N_32323,N_32432);
xor U39463 (N_39463,N_31423,N_33324);
nor U39464 (N_39464,N_32809,N_32401);
or U39465 (N_39465,N_34048,N_34860);
xor U39466 (N_39466,N_33210,N_34960);
xor U39467 (N_39467,N_33363,N_32354);
and U39468 (N_39468,N_31242,N_32718);
nor U39469 (N_39469,N_34886,N_33977);
nor U39470 (N_39470,N_33274,N_32667);
or U39471 (N_39471,N_31339,N_33499);
nand U39472 (N_39472,N_30679,N_31181);
xor U39473 (N_39473,N_30267,N_32056);
nand U39474 (N_39474,N_34069,N_30696);
and U39475 (N_39475,N_34801,N_30463);
nor U39476 (N_39476,N_33698,N_30277);
and U39477 (N_39477,N_31733,N_34793);
nand U39478 (N_39478,N_34083,N_32466);
nand U39479 (N_39479,N_34417,N_33497);
nor U39480 (N_39480,N_34075,N_30069);
xnor U39481 (N_39481,N_33872,N_33971);
xor U39482 (N_39482,N_33818,N_33245);
nand U39483 (N_39483,N_30722,N_34593);
and U39484 (N_39484,N_33809,N_34636);
xnor U39485 (N_39485,N_33747,N_32833);
nor U39486 (N_39486,N_33222,N_30081);
and U39487 (N_39487,N_32541,N_34791);
xnor U39488 (N_39488,N_34006,N_33140);
nand U39489 (N_39489,N_32266,N_32288);
or U39490 (N_39490,N_32417,N_30288);
and U39491 (N_39491,N_30047,N_32966);
and U39492 (N_39492,N_32315,N_30341);
or U39493 (N_39493,N_30284,N_32912);
nand U39494 (N_39494,N_30928,N_34921);
xnor U39495 (N_39495,N_34677,N_34913);
nor U39496 (N_39496,N_30624,N_32247);
nor U39497 (N_39497,N_33350,N_33775);
nor U39498 (N_39498,N_30464,N_30991);
or U39499 (N_39499,N_32770,N_31892);
xnor U39500 (N_39500,N_33071,N_32374);
and U39501 (N_39501,N_34897,N_34014);
nand U39502 (N_39502,N_30919,N_34219);
and U39503 (N_39503,N_34687,N_34458);
or U39504 (N_39504,N_31092,N_33001);
and U39505 (N_39505,N_32983,N_31898);
xnor U39506 (N_39506,N_30569,N_33182);
and U39507 (N_39507,N_31445,N_32927);
nor U39508 (N_39508,N_30897,N_31521);
and U39509 (N_39509,N_32270,N_34075);
xnor U39510 (N_39510,N_32132,N_32530);
xor U39511 (N_39511,N_32863,N_32885);
nor U39512 (N_39512,N_30958,N_32894);
xor U39513 (N_39513,N_34366,N_30742);
nor U39514 (N_39514,N_30543,N_34916);
xor U39515 (N_39515,N_30043,N_34117);
and U39516 (N_39516,N_34297,N_31878);
or U39517 (N_39517,N_31026,N_33076);
xnor U39518 (N_39518,N_33849,N_32314);
and U39519 (N_39519,N_32910,N_30338);
and U39520 (N_39520,N_31698,N_31720);
and U39521 (N_39521,N_33353,N_31543);
nor U39522 (N_39522,N_34147,N_30721);
and U39523 (N_39523,N_30415,N_34217);
and U39524 (N_39524,N_30433,N_30036);
xnor U39525 (N_39525,N_30370,N_33699);
and U39526 (N_39526,N_31545,N_30746);
and U39527 (N_39527,N_30497,N_30920);
and U39528 (N_39528,N_31473,N_33941);
and U39529 (N_39529,N_31433,N_34419);
xor U39530 (N_39530,N_33748,N_32170);
or U39531 (N_39531,N_31521,N_30735);
xnor U39532 (N_39532,N_32276,N_31953);
nand U39533 (N_39533,N_33538,N_34994);
or U39534 (N_39534,N_34081,N_33686);
xor U39535 (N_39535,N_33434,N_31062);
and U39536 (N_39536,N_33196,N_31055);
xor U39537 (N_39537,N_34946,N_32053);
nor U39538 (N_39538,N_32961,N_30182);
and U39539 (N_39539,N_33246,N_33004);
nand U39540 (N_39540,N_33540,N_32220);
xor U39541 (N_39541,N_32644,N_32168);
and U39542 (N_39542,N_31203,N_31982);
nor U39543 (N_39543,N_32220,N_34966);
nor U39544 (N_39544,N_30907,N_30519);
nor U39545 (N_39545,N_31760,N_33546);
xnor U39546 (N_39546,N_31298,N_32404);
xnor U39547 (N_39547,N_30645,N_32174);
and U39548 (N_39548,N_32027,N_32577);
and U39549 (N_39549,N_33763,N_30263);
and U39550 (N_39550,N_31456,N_30796);
xor U39551 (N_39551,N_31471,N_34580);
xor U39552 (N_39552,N_33513,N_34437);
nor U39553 (N_39553,N_34372,N_32477);
xor U39554 (N_39554,N_30965,N_31358);
nor U39555 (N_39555,N_30473,N_34954);
xor U39556 (N_39556,N_30467,N_30771);
and U39557 (N_39557,N_33508,N_33455);
nand U39558 (N_39558,N_34910,N_30921);
xnor U39559 (N_39559,N_33346,N_32380);
or U39560 (N_39560,N_33594,N_31474);
or U39561 (N_39561,N_32834,N_33079);
and U39562 (N_39562,N_32595,N_34147);
nor U39563 (N_39563,N_30264,N_31111);
xnor U39564 (N_39564,N_34763,N_30345);
xor U39565 (N_39565,N_33079,N_32036);
and U39566 (N_39566,N_32231,N_32086);
xnor U39567 (N_39567,N_32283,N_32153);
nor U39568 (N_39568,N_30713,N_33023);
and U39569 (N_39569,N_34332,N_32198);
xor U39570 (N_39570,N_30446,N_31064);
nor U39571 (N_39571,N_32056,N_30214);
or U39572 (N_39572,N_32434,N_32979);
nand U39573 (N_39573,N_34749,N_33506);
nand U39574 (N_39574,N_32563,N_32724);
or U39575 (N_39575,N_31777,N_34847);
or U39576 (N_39576,N_31754,N_33929);
nand U39577 (N_39577,N_32116,N_31662);
xnor U39578 (N_39578,N_32595,N_34422);
nand U39579 (N_39579,N_33022,N_34996);
and U39580 (N_39580,N_33551,N_32006);
or U39581 (N_39581,N_34645,N_34594);
and U39582 (N_39582,N_32764,N_31811);
nor U39583 (N_39583,N_30063,N_32292);
or U39584 (N_39584,N_32674,N_31503);
nor U39585 (N_39585,N_31036,N_33874);
nor U39586 (N_39586,N_30816,N_31959);
nor U39587 (N_39587,N_30333,N_30159);
nor U39588 (N_39588,N_31292,N_34597);
or U39589 (N_39589,N_31861,N_34214);
or U39590 (N_39590,N_31241,N_30292);
nor U39591 (N_39591,N_32558,N_32600);
xor U39592 (N_39592,N_33175,N_34409);
or U39593 (N_39593,N_30101,N_34760);
xnor U39594 (N_39594,N_30148,N_32607);
nor U39595 (N_39595,N_33865,N_33968);
xor U39596 (N_39596,N_31570,N_33835);
and U39597 (N_39597,N_31921,N_34189);
and U39598 (N_39598,N_33893,N_31117);
nor U39599 (N_39599,N_31492,N_33522);
or U39600 (N_39600,N_31256,N_34614);
nor U39601 (N_39601,N_33829,N_30105);
xor U39602 (N_39602,N_33623,N_33158);
and U39603 (N_39603,N_30067,N_33400);
and U39604 (N_39604,N_34439,N_34235);
or U39605 (N_39605,N_32144,N_30312);
or U39606 (N_39606,N_30734,N_30808);
and U39607 (N_39607,N_32703,N_31908);
or U39608 (N_39608,N_30627,N_31574);
xor U39609 (N_39609,N_34410,N_34265);
or U39610 (N_39610,N_30404,N_31700);
or U39611 (N_39611,N_30976,N_33067);
and U39612 (N_39612,N_31777,N_34225);
nand U39613 (N_39613,N_34291,N_33274);
or U39614 (N_39614,N_31839,N_33629);
nor U39615 (N_39615,N_30824,N_30403);
and U39616 (N_39616,N_33434,N_31815);
or U39617 (N_39617,N_33510,N_33001);
and U39618 (N_39618,N_31725,N_31157);
or U39619 (N_39619,N_33199,N_32549);
nand U39620 (N_39620,N_34139,N_31709);
xnor U39621 (N_39621,N_33679,N_30432);
xnor U39622 (N_39622,N_33874,N_32300);
xnor U39623 (N_39623,N_30342,N_31935);
and U39624 (N_39624,N_30888,N_33313);
and U39625 (N_39625,N_30931,N_30579);
and U39626 (N_39626,N_32177,N_34481);
or U39627 (N_39627,N_32519,N_34140);
nor U39628 (N_39628,N_32769,N_34161);
or U39629 (N_39629,N_33439,N_32959);
nor U39630 (N_39630,N_32387,N_31714);
and U39631 (N_39631,N_33879,N_33146);
or U39632 (N_39632,N_30238,N_33723);
nor U39633 (N_39633,N_30473,N_31439);
nor U39634 (N_39634,N_31058,N_34492);
or U39635 (N_39635,N_33942,N_34370);
and U39636 (N_39636,N_30639,N_32406);
and U39637 (N_39637,N_30210,N_31087);
nand U39638 (N_39638,N_31240,N_33748);
and U39639 (N_39639,N_32903,N_34952);
nor U39640 (N_39640,N_30887,N_30986);
and U39641 (N_39641,N_32297,N_34906);
nand U39642 (N_39642,N_32934,N_33385);
nand U39643 (N_39643,N_30194,N_33232);
nor U39644 (N_39644,N_31495,N_30121);
or U39645 (N_39645,N_30759,N_32144);
and U39646 (N_39646,N_30207,N_31958);
xnor U39647 (N_39647,N_33516,N_31789);
and U39648 (N_39648,N_31791,N_33675);
nor U39649 (N_39649,N_30089,N_33761);
nand U39650 (N_39650,N_31804,N_33972);
nor U39651 (N_39651,N_30840,N_32314);
or U39652 (N_39652,N_34977,N_30258);
or U39653 (N_39653,N_34699,N_30894);
nor U39654 (N_39654,N_30407,N_31781);
nand U39655 (N_39655,N_32408,N_31070);
and U39656 (N_39656,N_32750,N_32229);
nor U39657 (N_39657,N_31251,N_30821);
xnor U39658 (N_39658,N_30184,N_34713);
nand U39659 (N_39659,N_32351,N_34062);
and U39660 (N_39660,N_34226,N_32466);
nand U39661 (N_39661,N_34752,N_32973);
nand U39662 (N_39662,N_32259,N_34645);
xor U39663 (N_39663,N_34600,N_32028);
or U39664 (N_39664,N_34157,N_32341);
and U39665 (N_39665,N_30755,N_33853);
nor U39666 (N_39666,N_31019,N_31270);
or U39667 (N_39667,N_30654,N_30970);
xor U39668 (N_39668,N_34234,N_32959);
xor U39669 (N_39669,N_34665,N_32103);
or U39670 (N_39670,N_34079,N_30251);
or U39671 (N_39671,N_32877,N_32540);
and U39672 (N_39672,N_34789,N_31920);
nor U39673 (N_39673,N_30482,N_33750);
nor U39674 (N_39674,N_30153,N_31126);
nand U39675 (N_39675,N_34848,N_34182);
xnor U39676 (N_39676,N_32925,N_31832);
nand U39677 (N_39677,N_30891,N_31793);
xnor U39678 (N_39678,N_30376,N_32495);
or U39679 (N_39679,N_34558,N_31052);
nand U39680 (N_39680,N_32510,N_32169);
nor U39681 (N_39681,N_33968,N_34749);
xnor U39682 (N_39682,N_30716,N_31520);
and U39683 (N_39683,N_31917,N_34379);
nor U39684 (N_39684,N_33254,N_33767);
nor U39685 (N_39685,N_32399,N_32584);
or U39686 (N_39686,N_34300,N_33736);
xor U39687 (N_39687,N_33601,N_33188);
nor U39688 (N_39688,N_32140,N_31571);
nand U39689 (N_39689,N_33312,N_34183);
xor U39690 (N_39690,N_33237,N_34030);
and U39691 (N_39691,N_32110,N_34738);
xor U39692 (N_39692,N_34019,N_31325);
xor U39693 (N_39693,N_32310,N_30320);
nor U39694 (N_39694,N_33491,N_30248);
nor U39695 (N_39695,N_32880,N_33187);
nand U39696 (N_39696,N_33017,N_30380);
nand U39697 (N_39697,N_32390,N_34679);
xor U39698 (N_39698,N_30036,N_33209);
or U39699 (N_39699,N_33069,N_32105);
nand U39700 (N_39700,N_31413,N_32116);
nor U39701 (N_39701,N_30482,N_33130);
nor U39702 (N_39702,N_30780,N_31637);
or U39703 (N_39703,N_30454,N_32834);
or U39704 (N_39704,N_31437,N_34052);
nor U39705 (N_39705,N_34687,N_30223);
and U39706 (N_39706,N_34602,N_31378);
xnor U39707 (N_39707,N_32790,N_34614);
xnor U39708 (N_39708,N_31772,N_32762);
or U39709 (N_39709,N_31512,N_32205);
nand U39710 (N_39710,N_34770,N_32404);
xor U39711 (N_39711,N_33992,N_31858);
nand U39712 (N_39712,N_33158,N_30621);
or U39713 (N_39713,N_34404,N_30243);
nor U39714 (N_39714,N_30623,N_32311);
and U39715 (N_39715,N_33813,N_34119);
nor U39716 (N_39716,N_34147,N_32340);
nor U39717 (N_39717,N_30721,N_33474);
or U39718 (N_39718,N_31967,N_34966);
nand U39719 (N_39719,N_32829,N_33072);
and U39720 (N_39720,N_34822,N_32111);
and U39721 (N_39721,N_32728,N_34943);
nand U39722 (N_39722,N_33306,N_32751);
nand U39723 (N_39723,N_33543,N_33372);
xnor U39724 (N_39724,N_31127,N_30823);
nand U39725 (N_39725,N_33178,N_32745);
or U39726 (N_39726,N_33874,N_34183);
nand U39727 (N_39727,N_33118,N_30954);
nand U39728 (N_39728,N_31457,N_31339);
xor U39729 (N_39729,N_30265,N_34662);
xor U39730 (N_39730,N_34326,N_32136);
xor U39731 (N_39731,N_32844,N_30421);
nand U39732 (N_39732,N_30454,N_31517);
nand U39733 (N_39733,N_31032,N_30095);
nand U39734 (N_39734,N_30859,N_32884);
and U39735 (N_39735,N_33592,N_30413);
xor U39736 (N_39736,N_30503,N_30336);
and U39737 (N_39737,N_30179,N_30900);
nor U39738 (N_39738,N_30832,N_30122);
nand U39739 (N_39739,N_30332,N_32283);
and U39740 (N_39740,N_31879,N_32769);
or U39741 (N_39741,N_31327,N_33264);
nand U39742 (N_39742,N_30065,N_31305);
nand U39743 (N_39743,N_34898,N_32155);
nand U39744 (N_39744,N_32559,N_32972);
xor U39745 (N_39745,N_33040,N_31430);
nor U39746 (N_39746,N_33535,N_31784);
or U39747 (N_39747,N_31536,N_30825);
nand U39748 (N_39748,N_33275,N_34834);
xor U39749 (N_39749,N_30897,N_33795);
nor U39750 (N_39750,N_32275,N_30144);
and U39751 (N_39751,N_33319,N_34136);
nor U39752 (N_39752,N_34252,N_34066);
nor U39753 (N_39753,N_34731,N_31914);
nor U39754 (N_39754,N_31167,N_32488);
nor U39755 (N_39755,N_31198,N_33138);
and U39756 (N_39756,N_31473,N_31428);
xor U39757 (N_39757,N_32488,N_31864);
and U39758 (N_39758,N_34219,N_30540);
nand U39759 (N_39759,N_32460,N_34955);
nor U39760 (N_39760,N_33701,N_33072);
and U39761 (N_39761,N_33233,N_30840);
or U39762 (N_39762,N_30634,N_32292);
nand U39763 (N_39763,N_31208,N_34257);
nand U39764 (N_39764,N_33845,N_33337);
nand U39765 (N_39765,N_30179,N_30726);
nand U39766 (N_39766,N_32001,N_30562);
nor U39767 (N_39767,N_30371,N_33652);
and U39768 (N_39768,N_33838,N_33973);
nor U39769 (N_39769,N_34832,N_30792);
nand U39770 (N_39770,N_31918,N_34607);
nand U39771 (N_39771,N_33679,N_32286);
nand U39772 (N_39772,N_32869,N_31896);
xnor U39773 (N_39773,N_33885,N_31291);
nand U39774 (N_39774,N_30059,N_31463);
nor U39775 (N_39775,N_32974,N_32581);
and U39776 (N_39776,N_32390,N_31487);
nand U39777 (N_39777,N_31904,N_30289);
nor U39778 (N_39778,N_32785,N_32834);
and U39779 (N_39779,N_31364,N_32567);
nor U39780 (N_39780,N_34470,N_31017);
or U39781 (N_39781,N_34386,N_31712);
and U39782 (N_39782,N_33707,N_34744);
or U39783 (N_39783,N_30494,N_33145);
nor U39784 (N_39784,N_33282,N_31207);
nor U39785 (N_39785,N_33126,N_33933);
nor U39786 (N_39786,N_30664,N_34059);
nand U39787 (N_39787,N_30022,N_31716);
or U39788 (N_39788,N_32981,N_34898);
and U39789 (N_39789,N_34331,N_31668);
or U39790 (N_39790,N_31234,N_33984);
xnor U39791 (N_39791,N_34900,N_34834);
and U39792 (N_39792,N_33448,N_31719);
or U39793 (N_39793,N_31003,N_33390);
xor U39794 (N_39794,N_30133,N_30219);
and U39795 (N_39795,N_33839,N_31506);
and U39796 (N_39796,N_34680,N_32853);
nand U39797 (N_39797,N_30038,N_32392);
and U39798 (N_39798,N_33760,N_34313);
nand U39799 (N_39799,N_33024,N_33389);
and U39800 (N_39800,N_32536,N_32980);
or U39801 (N_39801,N_34109,N_34439);
and U39802 (N_39802,N_33990,N_30115);
or U39803 (N_39803,N_30167,N_30622);
or U39804 (N_39804,N_33243,N_31937);
nand U39805 (N_39805,N_34290,N_33040);
nand U39806 (N_39806,N_33222,N_30859);
xor U39807 (N_39807,N_31136,N_30892);
xnor U39808 (N_39808,N_31405,N_33729);
nor U39809 (N_39809,N_33840,N_34755);
nor U39810 (N_39810,N_32174,N_30048);
nand U39811 (N_39811,N_34113,N_34438);
nand U39812 (N_39812,N_30888,N_31927);
and U39813 (N_39813,N_31332,N_32076);
or U39814 (N_39814,N_33635,N_30688);
nor U39815 (N_39815,N_32829,N_31907);
nand U39816 (N_39816,N_34758,N_30296);
or U39817 (N_39817,N_33020,N_32104);
xor U39818 (N_39818,N_33325,N_32285);
xnor U39819 (N_39819,N_33034,N_33436);
xnor U39820 (N_39820,N_31383,N_31621);
xnor U39821 (N_39821,N_31048,N_32402);
and U39822 (N_39822,N_32263,N_32466);
xnor U39823 (N_39823,N_34645,N_33643);
xnor U39824 (N_39824,N_31899,N_34530);
xnor U39825 (N_39825,N_30032,N_34877);
or U39826 (N_39826,N_32674,N_30421);
or U39827 (N_39827,N_30548,N_33602);
nand U39828 (N_39828,N_32184,N_31127);
nor U39829 (N_39829,N_30545,N_32262);
nand U39830 (N_39830,N_31906,N_32822);
and U39831 (N_39831,N_34802,N_30525);
nor U39832 (N_39832,N_31634,N_34050);
or U39833 (N_39833,N_34036,N_33961);
and U39834 (N_39834,N_30559,N_30233);
and U39835 (N_39835,N_31346,N_32478);
xor U39836 (N_39836,N_33975,N_34822);
xor U39837 (N_39837,N_32115,N_30406);
xor U39838 (N_39838,N_32966,N_34353);
nand U39839 (N_39839,N_33524,N_30007);
or U39840 (N_39840,N_30766,N_30508);
xnor U39841 (N_39841,N_33221,N_32152);
xnor U39842 (N_39842,N_34862,N_32540);
or U39843 (N_39843,N_31140,N_33821);
and U39844 (N_39844,N_33523,N_34302);
and U39845 (N_39845,N_34652,N_34547);
nor U39846 (N_39846,N_30899,N_33380);
nand U39847 (N_39847,N_32533,N_30368);
nand U39848 (N_39848,N_31268,N_34972);
or U39849 (N_39849,N_33168,N_33224);
nor U39850 (N_39850,N_30021,N_31281);
nor U39851 (N_39851,N_31139,N_32078);
or U39852 (N_39852,N_31856,N_31565);
nand U39853 (N_39853,N_32857,N_32064);
or U39854 (N_39854,N_30651,N_33427);
xnor U39855 (N_39855,N_31119,N_32010);
or U39856 (N_39856,N_30259,N_32621);
xor U39857 (N_39857,N_32793,N_32198);
nor U39858 (N_39858,N_31639,N_31032);
nor U39859 (N_39859,N_33224,N_34479);
xnor U39860 (N_39860,N_34980,N_33779);
and U39861 (N_39861,N_31473,N_30815);
or U39862 (N_39862,N_32311,N_33549);
nand U39863 (N_39863,N_32785,N_32810);
or U39864 (N_39864,N_31792,N_30889);
and U39865 (N_39865,N_31483,N_33116);
and U39866 (N_39866,N_30956,N_34399);
nand U39867 (N_39867,N_30257,N_32003);
nand U39868 (N_39868,N_31554,N_32500);
and U39869 (N_39869,N_31473,N_32080);
and U39870 (N_39870,N_30541,N_33697);
and U39871 (N_39871,N_30710,N_30411);
nor U39872 (N_39872,N_31416,N_34726);
xnor U39873 (N_39873,N_31080,N_32829);
xor U39874 (N_39874,N_30426,N_31622);
or U39875 (N_39875,N_32867,N_31796);
nand U39876 (N_39876,N_34847,N_34791);
nand U39877 (N_39877,N_31051,N_33076);
or U39878 (N_39878,N_31253,N_31132);
nand U39879 (N_39879,N_32134,N_33164);
nor U39880 (N_39880,N_33569,N_31318);
nand U39881 (N_39881,N_32395,N_33859);
or U39882 (N_39882,N_34988,N_33802);
nand U39883 (N_39883,N_31210,N_34336);
nand U39884 (N_39884,N_31821,N_32357);
or U39885 (N_39885,N_30299,N_30180);
xor U39886 (N_39886,N_32136,N_34074);
or U39887 (N_39887,N_30013,N_30777);
or U39888 (N_39888,N_30943,N_31280);
or U39889 (N_39889,N_33016,N_30291);
and U39890 (N_39890,N_32685,N_30089);
or U39891 (N_39891,N_34698,N_32398);
xnor U39892 (N_39892,N_32262,N_33597);
nand U39893 (N_39893,N_34868,N_30354);
nand U39894 (N_39894,N_32316,N_31656);
and U39895 (N_39895,N_33606,N_30834);
or U39896 (N_39896,N_31291,N_34094);
or U39897 (N_39897,N_32647,N_33923);
xor U39898 (N_39898,N_31209,N_34922);
or U39899 (N_39899,N_34541,N_33679);
or U39900 (N_39900,N_32729,N_31882);
or U39901 (N_39901,N_30698,N_33919);
nand U39902 (N_39902,N_34301,N_32655);
nor U39903 (N_39903,N_34160,N_30236);
nor U39904 (N_39904,N_30446,N_32004);
nand U39905 (N_39905,N_30581,N_34243);
nor U39906 (N_39906,N_32630,N_31355);
or U39907 (N_39907,N_32348,N_33549);
xor U39908 (N_39908,N_33656,N_32219);
xnor U39909 (N_39909,N_34995,N_30284);
nand U39910 (N_39910,N_33988,N_30077);
nor U39911 (N_39911,N_34453,N_31173);
nand U39912 (N_39912,N_33207,N_30451);
nor U39913 (N_39913,N_33061,N_30017);
nand U39914 (N_39914,N_34467,N_31501);
xnor U39915 (N_39915,N_34719,N_33663);
xor U39916 (N_39916,N_31231,N_30745);
or U39917 (N_39917,N_32341,N_31775);
and U39918 (N_39918,N_32150,N_34050);
nor U39919 (N_39919,N_32617,N_32918);
and U39920 (N_39920,N_32933,N_32706);
nand U39921 (N_39921,N_30165,N_34963);
nor U39922 (N_39922,N_30502,N_33034);
nand U39923 (N_39923,N_30322,N_32731);
or U39924 (N_39924,N_32584,N_30852);
nand U39925 (N_39925,N_30527,N_30456);
xnor U39926 (N_39926,N_31615,N_32418);
nand U39927 (N_39927,N_32679,N_31530);
nor U39928 (N_39928,N_30234,N_32608);
nor U39929 (N_39929,N_30748,N_30460);
nand U39930 (N_39930,N_33094,N_32937);
nor U39931 (N_39931,N_30805,N_32695);
nor U39932 (N_39932,N_33344,N_32662);
xnor U39933 (N_39933,N_34279,N_32728);
and U39934 (N_39934,N_33807,N_34151);
xnor U39935 (N_39935,N_30876,N_30042);
nor U39936 (N_39936,N_31904,N_33645);
or U39937 (N_39937,N_34205,N_31677);
or U39938 (N_39938,N_33908,N_33826);
and U39939 (N_39939,N_32861,N_33985);
xor U39940 (N_39940,N_32150,N_30006);
or U39941 (N_39941,N_34782,N_31147);
and U39942 (N_39942,N_33159,N_32184);
and U39943 (N_39943,N_31215,N_33400);
and U39944 (N_39944,N_32700,N_31640);
nand U39945 (N_39945,N_34629,N_30461);
or U39946 (N_39946,N_31463,N_34411);
nand U39947 (N_39947,N_33762,N_31720);
xor U39948 (N_39948,N_32986,N_30949);
xor U39949 (N_39949,N_32667,N_30960);
and U39950 (N_39950,N_31780,N_31988);
and U39951 (N_39951,N_33967,N_32651);
nand U39952 (N_39952,N_33338,N_34690);
nand U39953 (N_39953,N_33487,N_32652);
nor U39954 (N_39954,N_34633,N_32613);
xor U39955 (N_39955,N_32661,N_33066);
and U39956 (N_39956,N_33739,N_30437);
xnor U39957 (N_39957,N_34208,N_33063);
or U39958 (N_39958,N_34427,N_33625);
xnor U39959 (N_39959,N_30740,N_34266);
and U39960 (N_39960,N_32439,N_31017);
nand U39961 (N_39961,N_34070,N_30145);
or U39962 (N_39962,N_32052,N_31948);
nor U39963 (N_39963,N_32539,N_33400);
xor U39964 (N_39964,N_34759,N_31634);
or U39965 (N_39965,N_33099,N_30588);
and U39966 (N_39966,N_32817,N_33402);
or U39967 (N_39967,N_31668,N_31195);
xnor U39968 (N_39968,N_33694,N_31853);
nand U39969 (N_39969,N_34731,N_30423);
and U39970 (N_39970,N_34220,N_32804);
nor U39971 (N_39971,N_30163,N_33452);
nand U39972 (N_39972,N_30156,N_34259);
xor U39973 (N_39973,N_33955,N_30245);
or U39974 (N_39974,N_30447,N_32755);
or U39975 (N_39975,N_32680,N_31211);
xor U39976 (N_39976,N_33814,N_30835);
nand U39977 (N_39977,N_32897,N_30219);
and U39978 (N_39978,N_33539,N_33951);
xor U39979 (N_39979,N_33656,N_30992);
xor U39980 (N_39980,N_33689,N_31309);
and U39981 (N_39981,N_33363,N_32562);
or U39982 (N_39982,N_32473,N_33513);
nor U39983 (N_39983,N_30753,N_30848);
nand U39984 (N_39984,N_33541,N_30013);
or U39985 (N_39985,N_31530,N_31409);
xor U39986 (N_39986,N_34852,N_32867);
nand U39987 (N_39987,N_33205,N_31710);
xor U39988 (N_39988,N_31806,N_31800);
xor U39989 (N_39989,N_30300,N_33722);
xnor U39990 (N_39990,N_32565,N_33326);
xor U39991 (N_39991,N_30792,N_34002);
nor U39992 (N_39992,N_31243,N_33129);
nand U39993 (N_39993,N_31133,N_31087);
or U39994 (N_39994,N_34687,N_33582);
xnor U39995 (N_39995,N_31414,N_31075);
nand U39996 (N_39996,N_32206,N_34208);
and U39997 (N_39997,N_34654,N_30887);
nor U39998 (N_39998,N_34536,N_34471);
and U39999 (N_39999,N_31505,N_34374);
nor U40000 (N_40000,N_39175,N_38743);
xor U40001 (N_40001,N_37299,N_36676);
nand U40002 (N_40002,N_35224,N_36139);
nand U40003 (N_40003,N_37691,N_38171);
nor U40004 (N_40004,N_35387,N_38236);
nand U40005 (N_40005,N_37255,N_36202);
and U40006 (N_40006,N_37371,N_36089);
nor U40007 (N_40007,N_39706,N_35554);
nand U40008 (N_40008,N_37151,N_38941);
xnor U40009 (N_40009,N_38953,N_38738);
xnor U40010 (N_40010,N_38485,N_37713);
and U40011 (N_40011,N_38603,N_39032);
and U40012 (N_40012,N_38257,N_36883);
xor U40013 (N_40013,N_38207,N_38042);
and U40014 (N_40014,N_37560,N_37445);
nor U40015 (N_40015,N_35966,N_37625);
xor U40016 (N_40016,N_37104,N_38669);
or U40017 (N_40017,N_37052,N_37665);
and U40018 (N_40018,N_39641,N_37499);
or U40019 (N_40019,N_37392,N_37931);
and U40020 (N_40020,N_38383,N_36802);
nand U40021 (N_40021,N_37131,N_37492);
or U40022 (N_40022,N_38612,N_35419);
nand U40023 (N_40023,N_37747,N_36307);
nor U40024 (N_40024,N_35599,N_37692);
xor U40025 (N_40025,N_39616,N_39995);
or U40026 (N_40026,N_37681,N_38378);
xor U40027 (N_40027,N_35201,N_36547);
or U40028 (N_40028,N_35027,N_37882);
xnor U40029 (N_40029,N_37021,N_39344);
and U40030 (N_40030,N_39850,N_39824);
or U40031 (N_40031,N_39454,N_39442);
xnor U40032 (N_40032,N_38949,N_37229);
nor U40033 (N_40033,N_35058,N_35729);
and U40034 (N_40034,N_35087,N_39337);
and U40035 (N_40035,N_37658,N_35824);
or U40036 (N_40036,N_39941,N_38896);
nor U40037 (N_40037,N_37087,N_39737);
or U40038 (N_40038,N_37136,N_39714);
nand U40039 (N_40039,N_36496,N_35032);
nand U40040 (N_40040,N_35162,N_35671);
nor U40041 (N_40041,N_38052,N_39860);
nor U40042 (N_40042,N_37077,N_36841);
nor U40043 (N_40043,N_36579,N_39167);
xor U40044 (N_40044,N_37535,N_35724);
or U40045 (N_40045,N_35461,N_35471);
or U40046 (N_40046,N_36261,N_35971);
or U40047 (N_40047,N_36673,N_38674);
xor U40048 (N_40048,N_38703,N_35026);
and U40049 (N_40049,N_35842,N_37615);
nor U40050 (N_40050,N_38475,N_37470);
nor U40051 (N_40051,N_35302,N_35636);
and U40052 (N_40052,N_38417,N_39245);
or U40053 (N_40053,N_39296,N_35832);
nand U40054 (N_40054,N_38777,N_35925);
or U40055 (N_40055,N_39434,N_37249);
and U40056 (N_40056,N_39488,N_35900);
nor U40057 (N_40057,N_39776,N_36978);
and U40058 (N_40058,N_36463,N_39393);
nand U40059 (N_40059,N_38157,N_37484);
or U40060 (N_40060,N_35979,N_37858);
nor U40061 (N_40061,N_36966,N_36095);
xor U40062 (N_40062,N_37836,N_35737);
xnor U40063 (N_40063,N_39387,N_35493);
nand U40064 (N_40064,N_36626,N_37770);
or U40065 (N_40065,N_39785,N_35287);
nor U40066 (N_40066,N_38254,N_39354);
or U40067 (N_40067,N_37483,N_36026);
or U40068 (N_40068,N_37965,N_38831);
or U40069 (N_40069,N_38027,N_39244);
nand U40070 (N_40070,N_37577,N_39186);
or U40071 (N_40071,N_37221,N_39038);
and U40072 (N_40072,N_35452,N_36554);
and U40073 (N_40073,N_35866,N_38387);
nand U40074 (N_40074,N_37324,N_35686);
xor U40075 (N_40075,N_36998,N_38039);
nor U40076 (N_40076,N_35303,N_38230);
and U40077 (N_40077,N_39106,N_39904);
nand U40078 (N_40078,N_37141,N_39794);
nand U40079 (N_40079,N_37944,N_37613);
xor U40080 (N_40080,N_38858,N_35080);
nand U40081 (N_40081,N_38182,N_36539);
nor U40082 (N_40082,N_36796,N_35407);
and U40083 (N_40083,N_39601,N_38734);
nand U40084 (N_40084,N_38906,N_36328);
xnor U40085 (N_40085,N_35383,N_38113);
xor U40086 (N_40086,N_36498,N_35219);
and U40087 (N_40087,N_38809,N_39916);
or U40088 (N_40088,N_39292,N_39265);
nand U40089 (N_40089,N_35542,N_37794);
xnor U40090 (N_40090,N_39473,N_39901);
or U40091 (N_40091,N_36321,N_38126);
and U40092 (N_40092,N_38249,N_36396);
nand U40093 (N_40093,N_37184,N_38062);
and U40094 (N_40094,N_35007,N_36381);
nor U40095 (N_40095,N_37070,N_39726);
nand U40096 (N_40096,N_37433,N_39382);
nand U40097 (N_40097,N_37870,N_35790);
xnor U40098 (N_40098,N_39788,N_38730);
and U40099 (N_40099,N_38801,N_36308);
nor U40100 (N_40100,N_36004,N_38694);
or U40101 (N_40101,N_37143,N_37404);
and U40102 (N_40102,N_36543,N_38471);
nand U40103 (N_40103,N_38465,N_35354);
nor U40104 (N_40104,N_35544,N_38707);
nor U40105 (N_40105,N_38793,N_37458);
nor U40106 (N_40106,N_36910,N_37901);
nand U40107 (N_40107,N_37972,N_37569);
xnor U40108 (N_40108,N_36657,N_37508);
nand U40109 (N_40109,N_38499,N_36532);
xor U40110 (N_40110,N_38851,N_38804);
nor U40111 (N_40111,N_37696,N_38141);
xor U40112 (N_40112,N_37773,N_36519);
nor U40113 (N_40113,N_35490,N_37271);
xor U40114 (N_40114,N_37817,N_37593);
or U40115 (N_40115,N_35752,N_38219);
and U40116 (N_40116,N_37695,N_35305);
xor U40117 (N_40117,N_39246,N_38129);
xor U40118 (N_40118,N_35972,N_39269);
xnor U40119 (N_40119,N_38544,N_35018);
nor U40120 (N_40120,N_36158,N_37015);
nand U40121 (N_40121,N_39126,N_39397);
nand U40122 (N_40122,N_36505,N_36552);
nor U40123 (N_40123,N_35973,N_36067);
nand U40124 (N_40124,N_39792,N_37262);
nor U40125 (N_40125,N_35516,N_35200);
and U40126 (N_40126,N_39999,N_37374);
or U40127 (N_40127,N_39515,N_39990);
and U40128 (N_40128,N_38296,N_38097);
nand U40129 (N_40129,N_39622,N_39055);
and U40130 (N_40130,N_37237,N_37095);
or U40131 (N_40131,N_39876,N_35336);
nand U40132 (N_40132,N_38842,N_37818);
nor U40133 (N_40133,N_35173,N_39567);
nand U40134 (N_40134,N_39880,N_39043);
xnor U40135 (N_40135,N_37285,N_37646);
xor U40136 (N_40136,N_38762,N_39896);
xor U40137 (N_40137,N_39070,N_39030);
and U40138 (N_40138,N_39683,N_36243);
nand U40139 (N_40139,N_39343,N_36355);
xor U40140 (N_40140,N_35564,N_36164);
or U40141 (N_40141,N_35584,N_39165);
and U40142 (N_40142,N_37573,N_39031);
nand U40143 (N_40143,N_35635,N_37551);
nor U40144 (N_40144,N_35556,N_35311);
xnor U40145 (N_40145,N_38456,N_39864);
and U40146 (N_40146,N_35702,N_38875);
xnor U40147 (N_40147,N_35100,N_37529);
xnor U40148 (N_40148,N_35112,N_35271);
xnor U40149 (N_40149,N_35454,N_39452);
xor U40150 (N_40150,N_37395,N_35951);
and U40151 (N_40151,N_38517,N_36290);
xor U40152 (N_40152,N_38711,N_35421);
nor U40153 (N_40153,N_36772,N_36990);
and U40154 (N_40154,N_36862,N_35946);
nand U40155 (N_40155,N_38224,N_36435);
and U40156 (N_40156,N_35353,N_35650);
and U40157 (N_40157,N_35897,N_39012);
or U40158 (N_40158,N_35758,N_35094);
nor U40159 (N_40159,N_37505,N_38772);
and U40160 (N_40160,N_37921,N_35869);
or U40161 (N_40161,N_37990,N_36981);
nor U40162 (N_40162,N_38285,N_39965);
and U40163 (N_40163,N_35196,N_36857);
nor U40164 (N_40164,N_35014,N_39029);
nand U40165 (N_40165,N_35432,N_38046);
nor U40166 (N_40166,N_35887,N_35507);
nand U40167 (N_40167,N_39383,N_36580);
nor U40168 (N_40168,N_37384,N_37074);
or U40169 (N_40169,N_37568,N_38754);
nor U40170 (N_40170,N_38019,N_39479);
or U40171 (N_40171,N_38839,N_38552);
nand U40172 (N_40172,N_36260,N_35155);
and U40173 (N_40173,N_39000,N_39644);
nor U40174 (N_40174,N_35130,N_35530);
xnor U40175 (N_40175,N_38739,N_36393);
xnor U40176 (N_40176,N_39893,N_39500);
and U40177 (N_40177,N_36369,N_37159);
or U40178 (N_40178,N_39624,N_39334);
xor U40179 (N_40179,N_35255,N_38859);
or U40180 (N_40180,N_35262,N_38946);
nor U40181 (N_40181,N_37339,N_38011);
and U40182 (N_40182,N_37664,N_35123);
or U40183 (N_40183,N_39604,N_38318);
and U40184 (N_40184,N_36336,N_39724);
or U40185 (N_40185,N_37047,N_36348);
and U40186 (N_40186,N_38108,N_38515);
nand U40187 (N_40187,N_35809,N_38290);
xnor U40188 (N_40188,N_39493,N_37419);
xor U40189 (N_40189,N_39404,N_36199);
and U40190 (N_40190,N_37083,N_39111);
and U40191 (N_40191,N_36378,N_35587);
and U40192 (N_40192,N_37631,N_35773);
nor U40193 (N_40193,N_37739,N_35601);
or U40194 (N_40194,N_35360,N_36662);
xor U40195 (N_40195,N_35669,N_37452);
or U40196 (N_40196,N_39594,N_39195);
and U40197 (N_40197,N_38758,N_35974);
xor U40198 (N_40198,N_38907,N_39221);
and U40199 (N_40199,N_38556,N_35010);
or U40200 (N_40200,N_36179,N_36891);
nand U40201 (N_40201,N_35395,N_36868);
or U40202 (N_40202,N_37154,N_36814);
or U40203 (N_40203,N_39820,N_39821);
xnor U40204 (N_40204,N_39749,N_39556);
nand U40205 (N_40205,N_37010,N_37148);
xnor U40206 (N_40206,N_36238,N_38960);
and U40207 (N_40207,N_36342,N_36610);
nand U40208 (N_40208,N_39056,N_35079);
and U40209 (N_40209,N_38643,N_39634);
or U40210 (N_40210,N_36134,N_37162);
nor U40211 (N_40211,N_35827,N_38461);
nand U40212 (N_40212,N_37734,N_37064);
or U40213 (N_40213,N_36959,N_37312);
and U40214 (N_40214,N_39710,N_38695);
nor U40215 (N_40215,N_39356,N_37116);
nor U40216 (N_40216,N_38699,N_38874);
and U40217 (N_40217,N_36402,N_39169);
xnor U40218 (N_40218,N_38176,N_37899);
and U40219 (N_40219,N_36939,N_39882);
nor U40220 (N_40220,N_35071,N_35846);
nor U40221 (N_40221,N_39329,N_35384);
nor U40222 (N_40222,N_39257,N_36175);
nor U40223 (N_40223,N_35644,N_39533);
nand U40224 (N_40224,N_36619,N_38657);
nor U40225 (N_40225,N_36473,N_39139);
or U40226 (N_40226,N_39808,N_35289);
and U40227 (N_40227,N_35132,N_38494);
and U40228 (N_40228,N_36176,N_39637);
or U40229 (N_40229,N_35486,N_35898);
or U40230 (N_40230,N_35975,N_35637);
or U40231 (N_40231,N_38281,N_36744);
nor U40232 (N_40232,N_36689,N_35046);
nand U40233 (N_40233,N_35822,N_36914);
nor U40234 (N_40234,N_38757,N_38597);
xor U40235 (N_40235,N_38186,N_38289);
nor U40236 (N_40236,N_37995,N_38197);
nand U40237 (N_40237,N_36390,N_38629);
xnor U40238 (N_40238,N_37690,N_38457);
nand U40239 (N_40239,N_39272,N_38449);
nor U40240 (N_40240,N_39077,N_38509);
nand U40241 (N_40241,N_35602,N_37466);
xor U40242 (N_40242,N_35894,N_38540);
and U40243 (N_40243,N_38355,N_35382);
nor U40244 (N_40244,N_39280,N_37081);
xnor U40245 (N_40245,N_39229,N_38838);
or U40246 (N_40246,N_39153,N_37630);
xnor U40247 (N_40247,N_35913,N_36082);
or U40248 (N_40248,N_35664,N_37055);
and U40249 (N_40249,N_36880,N_37843);
and U40250 (N_40250,N_38180,N_36251);
xor U40251 (N_40251,N_39017,N_38472);
nand U40252 (N_40252,N_39305,N_37698);
nand U40253 (N_40253,N_37133,N_37922);
or U40254 (N_40254,N_39587,N_35182);
and U40255 (N_40255,N_35772,N_38357);
and U40256 (N_40256,N_37938,N_38749);
xnor U40257 (N_40257,N_37795,N_38272);
and U40258 (N_40258,N_38969,N_39236);
or U40259 (N_40259,N_38425,N_37545);
nand U40260 (N_40260,N_37233,N_39028);
nand U40261 (N_40261,N_36596,N_38634);
or U40262 (N_40262,N_36613,N_39657);
or U40263 (N_40263,N_39781,N_38415);
nand U40264 (N_40264,N_39064,N_35133);
nand U40265 (N_40265,N_38265,N_35186);
xnor U40266 (N_40266,N_38366,N_35464);
nor U40267 (N_40267,N_38784,N_37934);
or U40268 (N_40268,N_38708,N_38879);
and U40269 (N_40269,N_35862,N_38479);
and U40270 (N_40270,N_36375,N_36096);
or U40271 (N_40271,N_37810,N_38395);
and U40272 (N_40272,N_37752,N_38534);
nand U40273 (N_40273,N_39342,N_36660);
or U40274 (N_40274,N_36138,N_39538);
xnor U40275 (N_40275,N_38825,N_36203);
nand U40276 (N_40276,N_37182,N_38309);
nor U40277 (N_40277,N_36540,N_36976);
and U40278 (N_40278,N_38312,N_36073);
and U40279 (N_40279,N_38174,N_37608);
and U40280 (N_40280,N_36852,N_36607);
and U40281 (N_40281,N_36156,N_36620);
and U40282 (N_40282,N_37600,N_36896);
nand U40283 (N_40283,N_35716,N_39478);
nor U40284 (N_40284,N_38218,N_37463);
or U40285 (N_40285,N_39203,N_35863);
or U40286 (N_40286,N_35300,N_35977);
nor U40287 (N_40287,N_38139,N_36823);
nor U40288 (N_40288,N_37910,N_37318);
and U40289 (N_40289,N_37506,N_38473);
xnor U40290 (N_40290,N_35796,N_36979);
and U40291 (N_40291,N_38592,N_36503);
or U40292 (N_40292,N_35472,N_35195);
and U40293 (N_40293,N_38950,N_36191);
and U40294 (N_40294,N_35704,N_39879);
and U40295 (N_40295,N_37661,N_35020);
and U40296 (N_40296,N_35778,N_38022);
xnor U40297 (N_40297,N_37949,N_36278);
xor U40298 (N_40298,N_36076,N_35498);
nand U40299 (N_40299,N_35188,N_39881);
nor U40300 (N_40300,N_37487,N_36001);
and U40301 (N_40301,N_39035,N_38028);
nand U40302 (N_40302,N_39540,N_37789);
nand U40303 (N_40303,N_37652,N_35470);
xnor U40304 (N_40304,N_35170,N_36597);
nand U40305 (N_40305,N_39079,N_37292);
and U40306 (N_40306,N_36833,N_35181);
xnor U40307 (N_40307,N_39095,N_39358);
or U40308 (N_40308,N_38870,N_35038);
or U40309 (N_40309,N_39608,N_35676);
xor U40310 (N_40310,N_39433,N_36143);
nand U40311 (N_40311,N_38342,N_35655);
and U40312 (N_40312,N_37926,N_35480);
nor U40313 (N_40313,N_36266,N_37044);
xor U40314 (N_40314,N_35418,N_38146);
nand U40315 (N_40315,N_37978,N_36403);
nor U40316 (N_40316,N_37641,N_35083);
or U40317 (N_40317,N_37422,N_36710);
xor U40318 (N_40318,N_39619,N_36545);
nand U40319 (N_40319,N_35138,N_38075);
or U40320 (N_40320,N_38454,N_35708);
or U40321 (N_40321,N_36112,N_35640);
xor U40322 (N_40322,N_38510,N_39279);
xor U40323 (N_40323,N_38590,N_39797);
and U40324 (N_40324,N_37620,N_36343);
nand U40325 (N_40325,N_35519,N_36709);
or U40326 (N_40326,N_35777,N_36454);
nor U40327 (N_40327,N_36031,N_35002);
and U40328 (N_40328,N_38700,N_37844);
xnor U40329 (N_40329,N_36037,N_35746);
and U40330 (N_40330,N_35060,N_37556);
or U40331 (N_40331,N_36758,N_38323);
or U40332 (N_40332,N_37796,N_39293);
nand U40333 (N_40333,N_36931,N_38687);
nand U40334 (N_40334,N_38910,N_35982);
and U40335 (N_40335,N_36904,N_36181);
nor U40336 (N_40336,N_38253,N_36229);
nand U40337 (N_40337,N_36424,N_38122);
or U40338 (N_40338,N_36086,N_36448);
nand U40339 (N_40339,N_39351,N_35738);
nor U40340 (N_40340,N_39579,N_38010);
nor U40341 (N_40341,N_38939,N_38353);
nand U40342 (N_40342,N_35926,N_38788);
and U40343 (N_40343,N_39859,N_39237);
or U40344 (N_40344,N_37937,N_35892);
xor U40345 (N_40345,N_36366,N_35786);
and U40346 (N_40346,N_39303,N_35412);
and U40347 (N_40347,N_39666,N_39123);
nand U40348 (N_40348,N_36510,N_36110);
or U40349 (N_40349,N_38764,N_35135);
xnor U40350 (N_40350,N_36080,N_37515);
nor U40351 (N_40351,N_38681,N_35627);
or U40352 (N_40352,N_35851,N_39371);
xnor U40353 (N_40353,N_35829,N_39044);
or U40354 (N_40354,N_35922,N_39900);
nor U40355 (N_40355,N_35312,N_36518);
nand U40356 (N_40356,N_36574,N_37357);
xor U40357 (N_40357,N_37375,N_39846);
nand U40358 (N_40358,N_36756,N_36337);
or U40359 (N_40359,N_35543,N_37627);
nor U40360 (N_40360,N_39671,N_35124);
or U40361 (N_40361,N_37190,N_36741);
and U40362 (N_40362,N_35625,N_35215);
xor U40363 (N_40363,N_38529,N_39348);
or U40364 (N_40364,N_37272,N_38343);
nor U40365 (N_40365,N_35469,N_37629);
xnor U40366 (N_40366,N_37587,N_38660);
or U40367 (N_40367,N_35485,N_35760);
nor U40368 (N_40368,N_39367,N_39467);
nor U40369 (N_40369,N_36386,N_39803);
nand U40370 (N_40370,N_37489,N_36791);
or U40371 (N_40371,N_39863,N_38761);
nand U40372 (N_40372,N_37401,N_36792);
or U40373 (N_40373,N_35216,N_36872);
xor U40374 (N_40374,N_39069,N_38892);
and U40375 (N_40375,N_37923,N_37779);
nand U40376 (N_40376,N_37171,N_36559);
nor U40377 (N_40377,N_36974,N_39232);
and U40378 (N_40378,N_39731,N_37056);
nor U40379 (N_40379,N_38106,N_36717);
xor U40380 (N_40380,N_36983,N_38142);
nand U40381 (N_40381,N_37442,N_36785);
nor U40382 (N_40382,N_36929,N_39325);
or U40383 (N_40383,N_37718,N_36021);
or U40384 (N_40384,N_37533,N_39906);
xnor U40385 (N_40385,N_38611,N_38880);
nor U40386 (N_40386,N_37114,N_37655);
xnor U40387 (N_40387,N_38393,N_38806);
nand U40388 (N_40388,N_37952,N_37050);
xnor U40389 (N_40389,N_38004,N_36887);
nor U40390 (N_40390,N_37111,N_38292);
nor U40391 (N_40391,N_36630,N_35097);
nand U40392 (N_40392,N_35441,N_38215);
nand U40393 (N_40393,N_36354,N_38388);
nand U40394 (N_40394,N_38966,N_37277);
nor U40395 (N_40395,N_38999,N_36712);
nand U40396 (N_40396,N_38242,N_35316);
nand U40397 (N_40397,N_35823,N_39968);
nor U40398 (N_40398,N_38688,N_38133);
or U40399 (N_40399,N_36609,N_38987);
xor U40400 (N_40400,N_35447,N_39048);
nor U40401 (N_40401,N_36578,N_36040);
or U40402 (N_40402,N_38557,N_39372);
or U40403 (N_40403,N_35742,N_35510);
or U40404 (N_40404,N_39867,N_37079);
nor U40405 (N_40405,N_36365,N_38427);
nand U40406 (N_40406,N_37389,N_39744);
and U40407 (N_40407,N_36136,N_37729);
nand U40408 (N_40408,N_35345,N_38134);
and U40409 (N_40409,N_39130,N_39670);
nor U40410 (N_40410,N_39027,N_35817);
xor U40411 (N_40411,N_37314,N_39886);
or U40412 (N_40412,N_35074,N_35500);
or U40413 (N_40413,N_38405,N_39625);
xnor U40414 (N_40414,N_38092,N_38581);
or U40415 (N_40415,N_35326,N_39872);
nor U40416 (N_40416,N_39685,N_38519);
or U40417 (N_40417,N_37820,N_38362);
xnor U40418 (N_40418,N_38310,N_36650);
and U40419 (N_40419,N_35552,N_37437);
nor U40420 (N_40420,N_37336,N_39914);
nand U40421 (N_40421,N_37859,N_35591);
nor U40422 (N_40422,N_39959,N_39003);
or U40423 (N_40423,N_38619,N_39779);
and U40424 (N_40424,N_35346,N_38955);
or U40425 (N_40425,N_38115,N_36687);
and U40426 (N_40426,N_39107,N_37837);
nand U40427 (N_40427,N_39837,N_35292);
nand U40428 (N_40428,N_36803,N_37181);
nor U40429 (N_40429,N_36070,N_35333);
nand U40430 (N_40430,N_37686,N_36252);
xor U40431 (N_40431,N_36331,N_37316);
nand U40432 (N_40432,N_35025,N_36735);
nor U40433 (N_40433,N_37707,N_39759);
nor U40434 (N_40434,N_35665,N_35781);
or U40435 (N_40435,N_38641,N_35684);
nand U40436 (N_40436,N_35914,N_36491);
and U40437 (N_40437,N_36416,N_36268);
nand U40438 (N_40438,N_37651,N_36999);
nor U40439 (N_40439,N_37955,N_38518);
xor U40440 (N_40440,N_35874,N_36779);
xnor U40441 (N_40441,N_36955,N_35288);
and U40442 (N_40442,N_38843,N_39613);
nand U40443 (N_40443,N_36264,N_37728);
nand U40444 (N_40444,N_37170,N_37367);
xor U40445 (N_40445,N_35902,N_38563);
nor U40446 (N_40446,N_37222,N_38948);
xor U40447 (N_40447,N_38931,N_36989);
xnor U40448 (N_40448,N_36697,N_37753);
nand U40449 (N_40449,N_38803,N_38390);
nand U40450 (N_40450,N_39969,N_35284);
xnor U40451 (N_40451,N_35482,N_38204);
xor U40452 (N_40452,N_38409,N_36392);
or U40453 (N_40453,N_37842,N_36973);
or U40454 (N_40454,N_39654,N_35313);
nand U40455 (N_40455,N_35899,N_37046);
xor U40456 (N_40456,N_37637,N_39739);
and U40457 (N_40457,N_39143,N_36899);
xnor U40458 (N_40458,N_36694,N_35298);
and U40459 (N_40459,N_36109,N_36279);
nand U40460 (N_40460,N_38338,N_37536);
nor U40461 (N_40461,N_36997,N_35129);
nor U40462 (N_40462,N_39199,N_35699);
nand U40463 (N_40463,N_39129,N_39703);
xnor U40464 (N_40464,N_36103,N_39173);
and U40465 (N_40465,N_39214,N_38496);
xor U40466 (N_40466,N_38691,N_35089);
or U40467 (N_40467,N_39956,N_36054);
nor U40468 (N_40468,N_37588,N_38579);
and U40469 (N_40469,N_37975,N_36430);
nor U40470 (N_40470,N_39388,N_36962);
nor U40471 (N_40471,N_35393,N_39224);
nor U40472 (N_40472,N_36917,N_38658);
or U40473 (N_40473,N_38091,N_38072);
or U40474 (N_40474,N_35828,N_39309);
nand U40475 (N_40475,N_39045,N_36077);
nor U40476 (N_40476,N_35411,N_38199);
nand U40477 (N_40477,N_37355,N_35558);
xnor U40478 (N_40478,N_38121,N_37228);
nand U40479 (N_40479,N_39525,N_36149);
nand U40480 (N_40480,N_39172,N_35947);
and U40481 (N_40481,N_38416,N_38169);
nand U40482 (N_40482,N_39004,N_35631);
nor U40483 (N_40483,N_38572,N_39696);
nor U40484 (N_40484,N_37542,N_35365);
xor U40485 (N_40485,N_36681,N_35950);
and U40486 (N_40486,N_35153,N_37302);
and U40487 (N_40487,N_35122,N_36882);
nor U40488 (N_40488,N_39420,N_36344);
and U40489 (N_40489,N_39469,N_37999);
or U40490 (N_40490,N_39593,N_35024);
nand U40491 (N_40491,N_36781,N_39066);
or U40492 (N_40492,N_37835,N_37390);
or U40493 (N_40493,N_39588,N_39888);
and U40494 (N_40494,N_38944,N_35810);
nor U40495 (N_40495,N_38869,N_37668);
or U40496 (N_40496,N_35279,N_37644);
nor U40497 (N_40497,N_36719,N_36595);
nor U40498 (N_40498,N_35244,N_37564);
and U40499 (N_40499,N_36668,N_35140);
nand U40500 (N_40500,N_35152,N_38368);
xor U40501 (N_40501,N_38912,N_38645);
nand U40502 (N_40502,N_36762,N_35662);
nand U40503 (N_40503,N_36520,N_38452);
and U40504 (N_40504,N_37400,N_39152);
and U40505 (N_40505,N_39840,N_38766);
or U40506 (N_40506,N_38566,N_35753);
xnor U40507 (N_40507,N_35672,N_39440);
xnor U40508 (N_40508,N_39966,N_35259);
nand U40509 (N_40509,N_39564,N_38017);
nand U40510 (N_40510,N_37449,N_37263);
and U40511 (N_40511,N_36043,N_37360);
or U40512 (N_40512,N_37240,N_38063);
xor U40513 (N_40513,N_37622,N_37227);
xnor U40514 (N_40514,N_36214,N_38434);
nand U40515 (N_40515,N_37998,N_36690);
xnor U40516 (N_40516,N_35595,N_37406);
and U40517 (N_40517,N_35763,N_37784);
nor U40518 (N_40518,N_35546,N_35301);
or U40519 (N_40519,N_35290,N_38630);
nor U40520 (N_40520,N_39887,N_37781);
and U40521 (N_40521,N_35506,N_39099);
or U40522 (N_40522,N_38817,N_36807);
nand U40523 (N_40523,N_35890,N_39252);
nand U40524 (N_40524,N_39891,N_38403);
or U40525 (N_40525,N_38511,N_39569);
xor U40526 (N_40526,N_38252,N_39205);
xor U40527 (N_40527,N_37887,N_35404);
nor U40528 (N_40528,N_39782,N_35831);
nor U40529 (N_40529,N_38714,N_37763);
or U40530 (N_40530,N_36345,N_38459);
xnor U40531 (N_40531,N_37900,N_38881);
and U40532 (N_40532,N_35849,N_36633);
xnor U40533 (N_40533,N_39428,N_37737);
or U40534 (N_40534,N_39162,N_38093);
nand U40535 (N_40535,N_39933,N_37428);
and U40536 (N_40536,N_36748,N_38025);
nor U40537 (N_40537,N_38702,N_35088);
and U40538 (N_40538,N_36172,N_36726);
or U40539 (N_40539,N_39057,N_38153);
nand U40540 (N_40540,N_39991,N_39184);
xnor U40541 (N_40541,N_39336,N_38038);
or U40542 (N_40542,N_36832,N_39427);
and U40543 (N_40543,N_37808,N_38627);
nor U40544 (N_40544,N_36783,N_39170);
or U40545 (N_40545,N_35037,N_39317);
nor U40546 (N_40546,N_36333,N_38591);
or U40547 (N_40547,N_36659,N_38000);
nand U40548 (N_40548,N_36192,N_37786);
or U40549 (N_40549,N_38363,N_35675);
nor U40550 (N_40550,N_38701,N_36154);
nand U40551 (N_40551,N_35852,N_39424);
and U40552 (N_40552,N_39958,N_35734);
nor U40553 (N_40553,N_36322,N_37596);
xnor U40554 (N_40554,N_38721,N_38808);
and U40555 (N_40555,N_38162,N_35990);
nor U40556 (N_40556,N_37501,N_38082);
and U40557 (N_40557,N_38018,N_39688);
nand U40558 (N_40558,N_39562,N_36384);
or U40559 (N_40559,N_38790,N_39176);
or U40560 (N_40560,N_36801,N_39519);
nand U40561 (N_40561,N_35160,N_36053);
nand U40562 (N_40562,N_39219,N_36319);
xnor U40563 (N_40563,N_35117,N_36774);
xor U40564 (N_40564,N_37675,N_36437);
and U40565 (N_40565,N_35513,N_35555);
nor U40566 (N_40566,N_36534,N_39104);
nand U40567 (N_40567,N_37523,N_36002);
or U40568 (N_40568,N_36851,N_35835);
xor U40569 (N_40569,N_39518,N_35323);
and U40570 (N_40570,N_36253,N_37412);
nand U40571 (N_40571,N_37597,N_35517);
and U40572 (N_40572,N_35011,N_36986);
or U40573 (N_40573,N_35363,N_37869);
xor U40574 (N_40574,N_36522,N_37498);
or U40575 (N_40575,N_39620,N_35803);
nor U40576 (N_40576,N_35009,N_36408);
and U40577 (N_40577,N_37238,N_39259);
nand U40578 (N_40578,N_39572,N_39676);
nand U40579 (N_40579,N_39947,N_39963);
or U40580 (N_40580,N_36315,N_37186);
or U40581 (N_40581,N_39929,N_35932);
nand U40582 (N_40582,N_36468,N_38088);
and U40583 (N_40583,N_35813,N_39482);
xor U40584 (N_40584,N_35369,N_36684);
nor U40585 (N_40585,N_36201,N_37599);
nor U40586 (N_40586,N_38668,N_38639);
or U40587 (N_40587,N_37623,N_37749);
nor U40588 (N_40588,N_38541,N_35717);
xnor U40589 (N_40589,N_36364,N_38277);
nor U40590 (N_40590,N_39128,N_35220);
nand U40591 (N_40591,N_36055,N_37555);
or U40592 (N_40592,N_35586,N_37929);
or U40593 (N_40593,N_35916,N_39502);
nor U40594 (N_40594,N_35771,N_37163);
nor U40595 (N_40595,N_38006,N_37574);
nand U40596 (N_40596,N_37543,N_35401);
or U40597 (N_40597,N_38671,N_38814);
xnor U40598 (N_40598,N_37063,N_35405);
or U40599 (N_40599,N_39728,N_37086);
nand U40600 (N_40600,N_35191,N_35068);
and U40601 (N_40601,N_39249,N_38005);
nor U40602 (N_40602,N_36221,N_35233);
nor U40603 (N_40603,N_37226,N_39302);
and U40604 (N_40604,N_39323,N_38787);
and U40605 (N_40605,N_39679,N_35611);
nand U40606 (N_40606,N_35962,N_35754);
xnor U40607 (N_40607,N_35864,N_39818);
xor U40608 (N_40608,N_35034,N_37744);
or U40609 (N_40609,N_35400,N_38905);
and U40610 (N_40610,N_38059,N_39379);
or U40611 (N_40611,N_35435,N_36631);
xnor U40612 (N_40612,N_36187,N_35527);
nand U40613 (N_40613,N_37746,N_37062);
or U40614 (N_40614,N_35172,N_35269);
and U40615 (N_40615,N_37269,N_38604);
nand U40616 (N_40616,N_35228,N_39815);
and U40617 (N_40617,N_36703,N_38505);
nor U40618 (N_40618,N_36793,N_37581);
nand U40619 (N_40619,N_36567,N_37275);
nor U40620 (N_40620,N_39185,N_35315);
xnor U40621 (N_40621,N_35197,N_36003);
or U40622 (N_40622,N_35652,N_37239);
and U40623 (N_40623,N_39885,N_35203);
xor U40624 (N_40624,N_37459,N_37478);
xor U40625 (N_40625,N_36444,N_36746);
and U40626 (N_40626,N_39196,N_37775);
xor U40627 (N_40627,N_38887,N_37471);
nor U40628 (N_40628,N_36871,N_35001);
nor U40629 (N_40629,N_37454,N_35232);
or U40630 (N_40630,N_38616,N_38663);
nor U40631 (N_40631,N_39415,N_37408);
nand U40632 (N_40632,N_38872,N_36525);
and U40633 (N_40633,N_38034,N_37082);
nor U40634 (N_40634,N_38271,N_37197);
xor U40635 (N_40635,N_35573,N_37425);
or U40636 (N_40636,N_39127,N_39970);
nor U40637 (N_40637,N_38287,N_39282);
or U40638 (N_40638,N_35528,N_35308);
xnor U40639 (N_40639,N_39610,N_37334);
xor U40640 (N_40640,N_38773,N_37212);
or U40641 (N_40641,N_38344,N_35993);
and U40642 (N_40642,N_39495,N_36141);
or U40643 (N_40643,N_35628,N_36132);
or U40644 (N_40644,N_36692,N_36301);
xor U40645 (N_40645,N_38098,N_37098);
and U40646 (N_40646,N_38512,N_37860);
nor U40647 (N_40647,N_38241,N_39228);
xnor U40648 (N_40648,N_37524,N_37361);
and U40649 (N_40649,N_36582,N_38374);
and U40650 (N_40650,N_35151,N_37252);
and U40651 (N_40651,N_37660,N_37298);
and U40652 (N_40652,N_39897,N_39444);
nand U40653 (N_40653,N_36737,N_39931);
or U40654 (N_40654,N_36995,N_36250);
or U40655 (N_40655,N_37467,N_35355);
nand U40656 (N_40656,N_39962,N_36713);
and U40657 (N_40657,N_39539,N_39135);
and U40658 (N_40658,N_37861,N_35910);
xnor U40659 (N_40659,N_36732,N_38873);
xnor U40660 (N_40660,N_39248,N_36600);
or U40661 (N_40661,N_35535,N_38064);
nand U40662 (N_40662,N_37963,N_36460);
nor U40663 (N_40663,N_37829,N_38545);
and U40664 (N_40664,N_35871,N_35670);
and U40665 (N_40665,N_38942,N_38369);
and U40666 (N_40666,N_36124,N_37880);
or U40667 (N_40667,N_37666,N_36296);
xnor U40668 (N_40668,N_35701,N_38262);
nor U40669 (N_40669,N_39211,N_38159);
or U40670 (N_40670,N_35938,N_38371);
nor U40671 (N_40671,N_38435,N_37798);
nand U40672 (N_40672,N_39376,N_36706);
nor U40673 (N_40673,N_39071,N_37871);
and U40674 (N_40674,N_39142,N_39485);
nand U40675 (N_40675,N_35350,N_38443);
nand U40676 (N_40676,N_38586,N_38615);
xor U40677 (N_40677,N_39357,N_39640);
nand U40678 (N_40678,N_39527,N_37078);
or U40679 (N_40679,N_38638,N_35649);
or U40680 (N_40680,N_35270,N_35901);
xor U40681 (N_40681,N_39513,N_35960);
or U40682 (N_40682,N_37806,N_37125);
and U40683 (N_40683,N_36930,N_36902);
or U40684 (N_40684,N_38516,N_38642);
xnor U40685 (N_40685,N_36407,N_36490);
nand U40686 (N_40686,N_39780,N_38255);
nor U40687 (N_40687,N_35171,N_36766);
xnor U40688 (N_40688,N_38882,N_37196);
and U40689 (N_40689,N_36818,N_37797);
nor U40690 (N_40690,N_38398,N_37916);
and U40691 (N_40691,N_37328,N_36024);
xnor U40692 (N_40692,N_37207,N_38086);
xnor U40693 (N_40693,N_38482,N_36449);
nor U40694 (N_40694,N_38151,N_35347);
xor U40695 (N_40695,N_36330,N_36679);
or U40696 (N_40696,N_37450,N_36213);
and U40697 (N_40697,N_38971,N_36151);
and U40698 (N_40698,N_39629,N_36541);
xor U40699 (N_40699,N_37838,N_39748);
xor U40700 (N_40700,N_35959,N_38123);
or U40701 (N_40701,N_36945,N_37805);
nor U40702 (N_40702,N_39116,N_38599);
nand U40703 (N_40703,N_35304,N_38903);
nor U40704 (N_40704,N_37917,N_36316);
xor U40705 (N_40705,N_39898,N_37853);
nor U40706 (N_40706,N_36953,N_35391);
nand U40707 (N_40707,N_35545,N_35429);
or U40708 (N_40708,N_36842,N_39270);
nand U40709 (N_40709,N_39800,N_36721);
nand U40710 (N_40710,N_37040,N_39465);
nor U40711 (N_40711,N_37007,N_35076);
nand U40712 (N_40712,N_38539,N_39766);
or U40713 (N_40713,N_37888,N_38746);
xnor U40714 (N_40714,N_37572,N_39051);
or U40715 (N_40715,N_38954,N_36122);
nand U40716 (N_40716,N_39516,N_37001);
xor U40717 (N_40717,N_35357,N_35961);
nand U40718 (N_40718,N_38661,N_39548);
xnor U40719 (N_40719,N_35057,N_36471);
xor U40720 (N_40720,N_35118,N_38648);
xnor U40721 (N_40721,N_35607,N_35836);
xor U40722 (N_40722,N_38431,N_35388);
nor U40723 (N_40723,N_35276,N_39431);
nor U40724 (N_40724,N_35580,N_38365);
or U40725 (N_40725,N_37935,N_39952);
xnor U40726 (N_40726,N_39338,N_38736);
or U40727 (N_40727,N_35168,N_35915);
or U40728 (N_40728,N_36924,N_38198);
xor U40729 (N_40729,N_37359,N_38300);
nor U40730 (N_40730,N_38439,N_37645);
or U40731 (N_40731,N_38484,N_38293);
nand U40732 (N_40732,N_39839,N_39487);
nand U40733 (N_40733,N_39691,N_38653);
nand U40734 (N_40734,N_35561,N_38811);
or U40735 (N_40735,N_37634,N_35307);
or U40736 (N_40736,N_35048,N_36798);
xor U40737 (N_40737,N_35450,N_39673);
or U40738 (N_40738,N_35502,N_39936);
nand U40739 (N_40739,N_36438,N_35750);
or U40740 (N_40740,N_39118,N_36215);
or U40741 (N_40741,N_36428,N_36729);
xnor U40742 (N_40742,N_35061,N_39403);
or U40743 (N_40743,N_37939,N_38911);
xnor U40744 (N_40744,N_38926,N_37697);
xor U40745 (N_40745,N_39732,N_36248);
or U40746 (N_40746,N_38846,N_35808);
nand U40747 (N_40747,N_35042,N_39817);
nor U40748 (N_40748,N_37563,N_36873);
or U40749 (N_40749,N_38883,N_37329);
and U40750 (N_40750,N_39994,N_38932);
nand U40751 (N_40751,N_39554,N_37873);
or U40752 (N_40752,N_36935,N_38014);
xnor U40753 (N_40753,N_39535,N_35731);
or U40754 (N_40754,N_39578,N_36432);
or U40755 (N_40755,N_35986,N_39979);
nand U40756 (N_40756,N_37030,N_39007);
or U40757 (N_40757,N_36612,N_38295);
nor U40758 (N_40758,N_38820,N_37828);
nor U40759 (N_40759,N_35062,N_38866);
xnor U40760 (N_40760,N_36380,N_38385);
and U40761 (N_40761,N_37293,N_36623);
and U40762 (N_40762,N_38074,N_39131);
nand U40763 (N_40763,N_38751,N_35820);
nand U40764 (N_40764,N_39986,N_36664);
or U40765 (N_40765,N_39178,N_35518);
and U40766 (N_40766,N_39586,N_36745);
and U40767 (N_40767,N_38468,N_38834);
nor U40768 (N_40768,N_37093,N_36527);
nand U40769 (N_40769,N_36184,N_38938);
or U40770 (N_40770,N_39677,N_39832);
nor U40771 (N_40771,N_37194,N_35756);
or U40772 (N_40772,N_36313,N_38455);
and U40773 (N_40773,N_36722,N_37430);
nor U40774 (N_40774,N_38677,N_37988);
or U40775 (N_40775,N_35840,N_39320);
xor U40776 (N_40776,N_36556,N_35968);
and U40777 (N_40777,N_38577,N_35257);
xor U40778 (N_40778,N_36224,N_37987);
nand U40779 (N_40779,N_35456,N_35185);
nand U40780 (N_40780,N_37033,N_36643);
or U40781 (N_40781,N_36038,N_37510);
nor U40782 (N_40782,N_39985,N_36087);
or U40783 (N_40783,N_35285,N_37997);
and U40784 (N_40784,N_37586,N_35217);
and U40785 (N_40785,N_36696,N_38543);
nor U40786 (N_40786,N_37800,N_35878);
nor U40787 (N_40787,N_38576,N_37742);
xor U40788 (N_40788,N_35251,N_39457);
or U40789 (N_40789,N_37821,N_35953);
nor U40790 (N_40790,N_37619,N_37013);
xor U40791 (N_40791,N_36538,N_39395);
and U40792 (N_40792,N_35620,N_37656);
xnor U40793 (N_40793,N_37059,N_36611);
nor U40794 (N_40794,N_39262,N_35804);
or U40795 (N_40795,N_37469,N_38261);
nand U40796 (N_40796,N_35695,N_39020);
nor U40797 (N_40797,N_35214,N_39076);
nand U40798 (N_40798,N_36346,N_38451);
and U40799 (N_40799,N_36361,N_36603);
xor U40800 (N_40800,N_38996,N_37254);
or U40801 (N_40801,N_35310,N_35022);
and U40802 (N_40802,N_35895,N_35722);
nor U40803 (N_40803,N_35949,N_39659);
and U40804 (N_40804,N_36410,N_37594);
and U40805 (N_40805,N_36764,N_35410);
xnor U40806 (N_40806,N_36933,N_36341);
nor U40807 (N_40807,N_39136,N_39783);
nand U40808 (N_40808,N_39526,N_38333);
nand U40809 (N_40809,N_36788,N_38913);
and U40810 (N_40810,N_36905,N_35463);
nand U40811 (N_40811,N_37168,N_37189);
nor U40812 (N_40812,N_36145,N_36434);
nor U40813 (N_40813,N_38481,N_36183);
nor U40814 (N_40814,N_38053,N_39543);
nor U40815 (N_40815,N_39549,N_39838);
nand U40816 (N_40816,N_37669,N_39772);
or U40817 (N_40817,N_39928,N_38350);
or U40818 (N_40818,N_36225,N_35161);
and U40819 (N_40819,N_36304,N_37122);
nor U40820 (N_40820,N_35988,N_35397);
or U40821 (N_40821,N_36325,N_35184);
nand U40822 (N_40822,N_36327,N_38084);
nor U40823 (N_40823,N_35096,N_36114);
or U40824 (N_40824,N_39822,N_39733);
nor U40825 (N_40825,N_39217,N_39346);
nor U40826 (N_40826,N_38165,N_36000);
nor U40827 (N_40827,N_37680,N_38968);
nor U40828 (N_40828,N_38536,N_38067);
nor U40829 (N_40829,N_37317,N_37160);
or U40830 (N_40830,N_39920,N_37223);
and U40831 (N_40831,N_35940,N_39103);
and U40832 (N_40832,N_38771,N_35525);
nand U40833 (N_40833,N_39767,N_37532);
or U40834 (N_40834,N_35816,N_36209);
or U40835 (N_40835,N_37772,N_36922);
nor U40836 (N_40836,N_35249,N_39132);
xnor U40837 (N_40837,N_35789,N_37205);
nand U40838 (N_40838,N_38904,N_38372);
and U40839 (N_40839,N_38555,N_39523);
xnor U40840 (N_40840,N_38217,N_39934);
nand U40841 (N_40841,N_36715,N_37409);
xor U40842 (N_40842,N_38348,N_35929);
xor U40843 (N_40843,N_38685,N_35077);
or U40844 (N_40844,N_38742,N_36399);
nand U40845 (N_40845,N_37693,N_38376);
or U40846 (N_40846,N_36749,N_37243);
or U40847 (N_40847,N_35505,N_38849);
nand U40848 (N_40848,N_35177,N_36035);
or U40849 (N_40849,N_37427,N_36671);
nor U40850 (N_40850,N_37120,N_38690);
and U40851 (N_40851,N_37591,N_38071);
nand U40852 (N_40852,N_39774,N_35449);
xnor U40853 (N_40853,N_39378,N_35327);
nand U40854 (N_40854,N_35614,N_36884);
and U40855 (N_40855,N_39147,N_36120);
and U40856 (N_40856,N_37852,N_35420);
xnor U40857 (N_40857,N_36566,N_39746);
nand U40858 (N_40858,N_39089,N_39836);
nor U40859 (N_40859,N_38538,N_35466);
xor U40860 (N_40860,N_35801,N_38178);
xnor U40861 (N_40861,N_39391,N_37167);
nand U40862 (N_40862,N_35691,N_37065);
xor U40863 (N_40863,N_36528,N_37793);
or U40864 (N_40864,N_37676,N_36569);
or U40865 (N_40865,N_37785,N_37348);
and U40866 (N_40866,N_38644,N_38320);
nand U40867 (N_40867,N_39894,N_37217);
nor U40868 (N_40868,N_38196,N_39163);
and U40869 (N_40869,N_35818,N_36812);
nand U40870 (N_40870,N_38193,N_35680);
nor U40871 (N_40871,N_38608,N_35157);
nor U40872 (N_40872,N_37420,N_35484);
and U40873 (N_40873,N_35212,N_35430);
and U40874 (N_40874,N_35710,N_35273);
or U40875 (N_40875,N_39187,N_37578);
nor U40876 (N_40876,N_37874,N_39417);
and U40877 (N_40877,N_37473,N_38023);
nor U40878 (N_40878,N_37178,N_37176);
nand U40879 (N_40879,N_35248,N_39067);
xnor U40880 (N_40880,N_35745,N_38394);
or U40881 (N_40881,N_35306,N_35385);
xnor U40882 (N_40882,N_35610,N_37671);
nor U40883 (N_40883,N_36615,N_35348);
or U40884 (N_40884,N_35479,N_36090);
nor U40885 (N_40885,N_37094,N_38990);
and U40886 (N_40886,N_39932,N_38917);
nor U40887 (N_40887,N_39108,N_36233);
and U40888 (N_40888,N_37106,N_39278);
xor U40889 (N_40889,N_35000,N_38447);
nand U40890 (N_40890,N_38266,N_37862);
nor U40891 (N_40891,N_35719,N_39695);
or U40892 (N_40892,N_37991,N_39660);
nor U40893 (N_40893,N_37363,N_35474);
and U40894 (N_40894,N_35293,N_39480);
xnor U40895 (N_40895,N_35945,N_38802);
and U40896 (N_40896,N_36349,N_39429);
xnor U40897 (N_40897,N_39496,N_35534);
xnor U40898 (N_40898,N_38797,N_36455);
nand U40899 (N_40899,N_36062,N_39456);
nor U40900 (N_40900,N_35783,N_35349);
xnor U40901 (N_40901,N_38807,N_39699);
or U40902 (N_40902,N_35263,N_37288);
nor U40903 (N_40903,N_35509,N_36677);
nand U40904 (N_40904,N_38340,N_37310);
nand U40905 (N_40905,N_36845,N_36100);
nand U40906 (N_40906,N_35029,N_36537);
and U40907 (N_40907,N_35991,N_35937);
nand U40908 (N_40908,N_39421,N_36377);
or U40909 (N_40909,N_35596,N_38593);
and U40910 (N_40910,N_35568,N_36502);
or U40911 (N_40911,N_36140,N_39981);
and U40912 (N_40912,N_37343,N_39735);
xnor U40913 (N_40913,N_36280,N_39407);
nand U40914 (N_40914,N_38716,N_35240);
nand U40915 (N_40915,N_38030,N_36442);
and U40916 (N_40916,N_37491,N_38578);
nand U40917 (N_40917,N_35314,N_38925);
and U40918 (N_40918,N_36093,N_39723);
and U40919 (N_40919,N_38497,N_39791);
and U40920 (N_40920,N_37758,N_36934);
xor U40921 (N_40921,N_35939,N_38232);
or U40922 (N_40922,N_37721,N_38399);
nand U40923 (N_40923,N_35660,N_37530);
nand U40924 (N_40924,N_37134,N_36177);
or U40925 (N_40925,N_38920,N_37018);
and U40926 (N_40926,N_38561,N_35524);
nand U40927 (N_40927,N_38209,N_38335);
nor U40928 (N_40928,N_38130,N_39568);
nand U40929 (N_40929,N_39288,N_36648);
xnor U40930 (N_40930,N_38020,N_35948);
nor U40931 (N_40931,N_39146,N_39945);
xor U40932 (N_40932,N_39258,N_39001);
or U40933 (N_40933,N_35639,N_37100);
xor U40934 (N_40934,N_37397,N_38136);
and U40935 (N_40935,N_38506,N_36769);
and U40936 (N_40936,N_36227,N_38601);
nand U40937 (N_40937,N_35043,N_37684);
nor U40938 (N_40938,N_36634,N_35780);
nor U40939 (N_40939,N_35164,N_36016);
nand U40940 (N_40940,N_36602,N_36754);
nand U40941 (N_40941,N_39805,N_35807);
nor U40942 (N_40942,N_35070,N_37598);
or U40943 (N_40943,N_38860,N_36018);
or U40944 (N_40944,N_37672,N_36890);
and U40945 (N_40945,N_39266,N_36773);
nand U40946 (N_40946,N_39092,N_37297);
nor U40947 (N_40947,N_39392,N_39542);
nand U40948 (N_40948,N_38172,N_36500);
and U40949 (N_40949,N_36276,N_38732);
nand U40950 (N_40950,N_36885,N_38109);
nor U40951 (N_40951,N_38240,N_39662);
or U40952 (N_40952,N_37416,N_39565);
nor U40953 (N_40953,N_37144,N_35896);
nand U40954 (N_40954,N_38205,N_37014);
nor U40955 (N_40955,N_38192,N_36827);
and U40956 (N_40956,N_39238,N_38741);
and U40957 (N_40957,N_37138,N_37762);
and U40958 (N_40958,N_37069,N_36670);
and U40959 (N_40959,N_37017,N_35918);
nand U40960 (N_40960,N_35206,N_38974);
nand U40961 (N_40961,N_35213,N_36064);
nor U40962 (N_40962,N_35150,N_39062);
nor U40963 (N_40963,N_36810,N_38201);
nand U40964 (N_40964,N_38675,N_36019);
xor U40965 (N_40965,N_37291,N_37258);
nor U40966 (N_40966,N_36599,N_35533);
and U40967 (N_40967,N_39655,N_38560);
or U40968 (N_40968,N_36244,N_37539);
nor U40969 (N_40969,N_38282,N_35199);
nand U40970 (N_40970,N_36817,N_36941);
nand U40971 (N_40971,N_36996,N_39693);
nand U40972 (N_40972,N_37809,N_37462);
xnor U40973 (N_40973,N_39580,N_39472);
nand U40974 (N_40974,N_35582,N_38582);
and U40975 (N_40975,N_37172,N_36317);
nor U40976 (N_40976,N_37043,N_36629);
nand U40977 (N_40977,N_37225,N_38723);
nor U40978 (N_40978,N_36092,N_38649);
xnor U40979 (N_40979,N_37628,N_38508);
nor U40980 (N_40980,N_36245,N_36632);
xor U40981 (N_40981,N_36309,N_36094);
nand U40982 (N_40982,N_39722,N_38476);
and U40983 (N_40983,N_37000,N_37626);
xor U40984 (N_40984,N_39024,N_36457);
and U40985 (N_40985,N_39939,N_35368);
or U40986 (N_40986,N_39284,N_37868);
nand U40987 (N_40987,N_36494,N_38624);
and U40988 (N_40988,N_37496,N_39909);
and U40989 (N_40989,N_37799,N_39982);
xor U40990 (N_40990,N_35843,N_35149);
and U40991 (N_40991,N_35770,N_37128);
nor U40992 (N_40992,N_35163,N_38503);
or U40993 (N_40993,N_36382,N_37831);
and U40994 (N_40994,N_35943,N_37146);
nand U40995 (N_40995,N_35893,N_35877);
nor U40996 (N_40996,N_39339,N_36830);
nand U40997 (N_40997,N_35682,N_38606);
xnor U40998 (N_40998,N_39015,N_39046);
and U40999 (N_40999,N_36198,N_39674);
xnor U41000 (N_41000,N_38893,N_35254);
nand U41001 (N_41001,N_35928,N_36461);
nand U41002 (N_41002,N_37989,N_38692);
or U41003 (N_41003,N_39289,N_37218);
nand U41004 (N_41004,N_37242,N_38623);
and U41005 (N_41005,N_36404,N_38760);
nor U41006 (N_41006,N_37204,N_37554);
nor U41007 (N_41007,N_36763,N_35075);
nor U41008 (N_41008,N_38554,N_35261);
and U41009 (N_41009,N_38725,N_37771);
nor U41010 (N_41010,N_37121,N_39917);
nand U41011 (N_41011,N_39755,N_36759);
xor U41012 (N_41012,N_39848,N_39450);
or U41013 (N_41013,N_39584,N_37219);
or U41014 (N_41014,N_37444,N_36376);
xnor U41015 (N_41015,N_36340,N_38867);
and U41016 (N_41016,N_36312,N_37231);
or U41017 (N_41017,N_38607,N_37147);
nand U41018 (N_41018,N_35028,N_37192);
or U41019 (N_41019,N_39607,N_36078);
nand U41020 (N_41020,N_35721,N_37438);
nor U41021 (N_41021,N_38567,N_38923);
and U41022 (N_41022,N_36853,N_36398);
and U41023 (N_41023,N_39085,N_39151);
nor U41024 (N_41024,N_36509,N_36289);
nand U41025 (N_41025,N_36374,N_38163);
and U41026 (N_41026,N_39830,N_36451);
nand U41027 (N_41027,N_39623,N_39823);
nor U41028 (N_41028,N_39852,N_35374);
nor U41029 (N_41029,N_36129,N_37886);
nand U41030 (N_41030,N_39406,N_35126);
or U41031 (N_41031,N_38956,N_36919);
xnor U41032 (N_41032,N_37827,N_37703);
xnor U41033 (N_41033,N_35854,N_38755);
xnor U41034 (N_41034,N_35084,N_36757);
xnor U41035 (N_41035,N_38313,N_39188);
or U41036 (N_41036,N_39633,N_37735);
or U41037 (N_41037,N_38190,N_37702);
and U41038 (N_41038,N_36714,N_38640);
xor U41039 (N_41039,N_38886,N_38048);
nor U41040 (N_41040,N_37475,N_39242);
xor U41041 (N_41041,N_37280,N_35183);
nand U41042 (N_41042,N_38429,N_38154);
nand U41043 (N_41043,N_37354,N_37722);
nand U41044 (N_41044,N_35139,N_35706);
nand U41045 (N_41045,N_37431,N_35406);
xnor U41046 (N_41046,N_37177,N_38596);
xor U41047 (N_41047,N_35208,N_38502);
nor U41048 (N_41048,N_38148,N_36881);
xnor U41049 (N_41049,N_37504,N_39112);
nand U41050 (N_41050,N_39254,N_38234);
xor U41051 (N_41051,N_39426,N_35376);
or U41052 (N_41052,N_37503,N_36863);
nor U41053 (N_41053,N_37962,N_35529);
nand U41054 (N_41054,N_35583,N_35653);
nor U41055 (N_41055,N_36107,N_36936);
and U41056 (N_41056,N_38238,N_38054);
xnor U41057 (N_41057,N_38036,N_39856);
nand U41058 (N_41058,N_35012,N_35996);
nor U41059 (N_41059,N_39047,N_39809);
or U41060 (N_41060,N_39026,N_35616);
xor U41061 (N_41061,N_37783,N_38617);
or U41062 (N_41062,N_35559,N_38750);
nor U41063 (N_41063,N_36819,N_35755);
nor U41064 (N_41064,N_36108,N_39855);
nor U41065 (N_41065,N_36504,N_37933);
or U41066 (N_41066,N_35379,N_35187);
or U41067 (N_41067,N_38278,N_35747);
and U41068 (N_41068,N_35439,N_36795);
and U41069 (N_41069,N_38037,N_37053);
and U41070 (N_41070,N_35229,N_37804);
and U41071 (N_41071,N_39350,N_37893);
and U41072 (N_41072,N_39875,N_39115);
nand U41073 (N_41073,N_37261,N_36324);
or U41074 (N_41074,N_38525,N_36169);
or U41075 (N_41075,N_37051,N_35047);
nand U41076 (N_41076,N_39512,N_36589);
and U41077 (N_41077,N_36686,N_37378);
or U41078 (N_41078,N_35459,N_36269);
nor U41079 (N_41079,N_35539,N_38495);
xnor U41080 (N_41080,N_39018,N_38728);
nor U41081 (N_41081,N_36993,N_39842);
nand U41082 (N_41082,N_39707,N_36014);
and U41083 (N_41083,N_36674,N_38135);
or U41084 (N_41084,N_37259,N_35615);
and U41085 (N_41085,N_39041,N_37481);
xnor U41086 (N_41086,N_35609,N_37802);
nor U41087 (N_41087,N_38364,N_36163);
xnor U41088 (N_41088,N_39425,N_38410);
nand U41089 (N_41089,N_36265,N_36865);
or U41090 (N_41090,N_38306,N_36071);
nand U41091 (N_41091,N_37399,N_36970);
nor U41092 (N_41092,N_39144,N_35531);
nand U41093 (N_41093,N_36780,N_39943);
and U41094 (N_41094,N_35204,N_35861);
nor U41095 (N_41095,N_35859,N_39443);
nor U41096 (N_41096,N_39019,N_37443);
nor U41097 (N_41097,N_35496,N_39052);
nand U41098 (N_41098,N_36693,N_38845);
xnor U41099 (N_41099,N_37407,N_38177);
nor U41100 (N_41100,N_38361,N_37417);
or U41101 (N_41101,N_37216,N_38523);
and U41102 (N_41102,N_38246,N_37076);
nand U41103 (N_41103,N_38175,N_35501);
nand U41104 (N_41104,N_38170,N_38450);
and U41105 (N_41105,N_36012,N_38856);
and U41106 (N_41106,N_35098,N_35361);
xnor U41107 (N_41107,N_35885,N_38977);
or U41108 (N_41108,N_39105,N_35833);
or U41109 (N_41109,N_38167,N_39948);
xor U41110 (N_41110,N_38765,N_39998);
nor U41111 (N_41111,N_39762,N_36414);
nor U41112 (N_41112,N_35508,N_38448);
nand U41113 (N_41113,N_39484,N_39294);
nand U41114 (N_41114,N_39438,N_39460);
nand U41115 (N_41115,N_35845,N_37954);
nand U41116 (N_41116,N_37777,N_38559);
xor U41117 (N_41117,N_37200,N_35330);
or U41118 (N_41118,N_39234,N_36666);
or U41119 (N_41119,N_37980,N_39923);
and U41120 (N_41120,N_36809,N_38991);
nand U41121 (N_41121,N_37156,N_36548);
and U41122 (N_41122,N_36123,N_35666);
nor U41123 (N_41123,N_37925,N_36022);
nand U41124 (N_41124,N_37319,N_38469);
nand U41125 (N_41125,N_36656,N_38101);
and U41126 (N_41126,N_38339,N_35797);
or U41127 (N_41127,N_35956,N_36050);
or U41128 (N_41128,N_35794,N_36583);
or U41129 (N_41129,N_39756,N_36332);
nand U41130 (N_41130,N_35218,N_39037);
nand U41131 (N_41131,N_39597,N_35723);
and U41132 (N_41132,N_39725,N_35134);
xnor U41133 (N_41133,N_39286,N_35390);
or U41134 (N_41134,N_38124,N_36678);
and U41135 (N_41135,N_35622,N_38813);
or U41136 (N_41136,N_36888,N_39890);
or U41137 (N_41137,N_36535,N_35253);
nand U41138 (N_41138,N_35839,N_38722);
and U41139 (N_41139,N_36299,N_38291);
nor U41140 (N_41140,N_38408,N_35222);
nor U41141 (N_41141,N_38975,N_36728);
and U41142 (N_41142,N_39878,N_37137);
xnor U41143 (N_41143,N_38040,N_39834);
nor U41144 (N_41144,N_35136,N_39093);
xor U41145 (N_41145,N_39441,N_39667);
and U41146 (N_41146,N_36222,N_39377);
or U41147 (N_41147,N_39312,N_39068);
xnor U41148 (N_41148,N_36226,N_38909);
xnor U41149 (N_41149,N_36858,N_38740);
nor U41150 (N_41150,N_37441,N_35984);
or U41151 (N_41151,N_38119,N_37943);
xnor U41152 (N_41152,N_38789,N_35492);
nand U41153 (N_41153,N_35581,N_36568);
or U41154 (N_41154,N_38031,N_39256);
xnor U41155 (N_41155,N_39612,N_36915);
xnor U41156 (N_41156,N_36452,N_39432);
nand U41157 (N_41157,N_36305,N_38462);
or U41158 (N_41158,N_39713,N_38780);
nor U41159 (N_41159,N_35433,N_35883);
or U41160 (N_41160,N_39150,N_36755);
nor U41161 (N_41161,N_35538,N_36052);
nand U41162 (N_41162,N_39075,N_37974);
nand U41163 (N_41163,N_37833,N_37413);
or U41164 (N_41164,N_37748,N_39918);
or U41165 (N_41165,N_38426,N_39757);
nor U41166 (N_41166,N_37115,N_39609);
nor U41167 (N_41167,N_36358,N_39180);
or U41168 (N_41168,N_37029,N_39806);
or U41169 (N_41169,N_37132,N_35970);
or U41170 (N_41170,N_35053,N_37382);
nand U41171 (N_41171,N_35954,N_38352);
xor U41172 (N_41172,N_36969,N_38090);
nand U41173 (N_41173,N_38747,N_38983);
and U41174 (N_41174,N_36440,N_39740);
and U41175 (N_41175,N_38706,N_39661);
xnor U41176 (N_41176,N_36529,N_39843);
nor U41177 (N_41177,N_36029,N_36775);
and U41178 (N_41178,N_37448,N_38709);
nand U41179 (N_41179,N_39574,N_37418);
and U41180 (N_41180,N_36831,N_37107);
or U41181 (N_41181,N_36507,N_39536);
nand U41182 (N_41182,N_36039,N_36048);
xor U41183 (N_41183,N_38021,N_35165);
nand U41184 (N_41184,N_35967,N_38621);
nand U41185 (N_41185,N_38144,N_38213);
and U41186 (N_41186,N_36824,N_35748);
or U41187 (N_41187,N_39529,N_36085);
nand U41188 (N_41188,N_37035,N_37307);
xnor U41189 (N_41189,N_35234,N_37436);
nand U41190 (N_41190,N_35236,N_38094);
xor U41191 (N_41191,N_35571,N_39040);
and U41192 (N_41192,N_36940,N_35904);
xnor U41193 (N_41193,N_39300,N_35757);
xnor U41194 (N_41194,N_36815,N_38164);
nor U41195 (N_41195,N_37103,N_36943);
nor U41196 (N_41196,N_39617,N_38958);
nand U41197 (N_41197,N_38225,N_38537);
and U41198 (N_41198,N_38962,N_36727);
nor U41199 (N_41199,N_37650,N_39719);
and U41200 (N_41200,N_38947,N_36958);
or U41201 (N_41201,N_36489,N_39649);
or U41202 (N_41202,N_36682,N_36608);
or U41203 (N_41203,N_37610,N_39133);
or U41204 (N_41204,N_39039,N_36370);
nor U41205 (N_41205,N_35965,N_36638);
nand U41206 (N_41206,N_37751,N_36592);
xnor U41207 (N_41207,N_35019,N_36799);
xnor U41208 (N_41208,N_39109,N_38189);
xor U41209 (N_41209,N_39384,N_36663);
or U41210 (N_41210,N_38487,N_37139);
or U41211 (N_41211,N_38636,N_36649);
and U41212 (N_41212,N_39149,N_36223);
nor U41213 (N_41213,N_37723,N_38463);
and U41214 (N_41214,N_36820,N_35371);
nor U41215 (N_41215,N_36778,N_38096);
nor U41216 (N_41216,N_36256,N_39097);
nor U41217 (N_41217,N_35180,N_37127);
and U41218 (N_41218,N_36300,N_35329);
nand U41219 (N_41219,N_38832,N_36283);
nand U41220 (N_41220,N_38898,N_35099);
nand U41221 (N_41221,N_39910,N_38901);
xnor U41222 (N_41222,N_37150,N_36571);
xor U41223 (N_41223,N_35499,N_36481);
and U41224 (N_41224,N_36517,N_38216);
xor U41225 (N_41225,N_35440,N_39650);
and U41226 (N_41226,N_36084,N_35462);
and U41227 (N_41227,N_39669,N_35434);
xor U41228 (N_41228,N_39489,N_39464);
or U41229 (N_41229,N_36614,N_37928);
or U41230 (N_41230,N_38493,N_38149);
and U41231 (N_41231,N_38620,N_35800);
nand U41232 (N_41232,N_39492,N_36486);
and U41233 (N_41233,N_36514,N_38445);
nand U41234 (N_41234,N_35109,N_36718);
nand U41235 (N_41235,N_39183,N_37550);
or U41236 (N_41236,N_35051,N_37678);
or U41237 (N_41237,N_36160,N_39812);
nor U41238 (N_41238,N_36549,N_35931);
xor U41239 (N_41239,N_38667,N_38035);
nor U41240 (N_41240,N_39734,N_37731);
nor U41241 (N_41241,N_35339,N_39632);
xnor U41242 (N_41242,N_37090,N_37527);
nand U41243 (N_41243,N_35557,N_39179);
xor U41244 (N_41244,N_36837,N_37265);
nor U41245 (N_41245,N_38520,N_37440);
xnor U41246 (N_41246,N_37927,N_38995);
nand U41247 (N_41247,N_36189,N_39304);
xor U41248 (N_41248,N_37346,N_35613);
nor U41249 (N_41249,N_39287,N_38251);
and U41250 (N_41250,N_38574,N_38637);
xnor U41251 (N_41251,N_35765,N_38354);
xor U41252 (N_41252,N_36733,N_36072);
or U41253 (N_41253,N_37589,N_35647);
and U41254 (N_41254,N_35567,N_38840);
or U41255 (N_41255,N_36695,N_36911);
xor U41256 (N_41256,N_36418,N_39462);
and U41257 (N_41257,N_37472,N_35193);
nor U41258 (N_41258,N_37959,N_38570);
nand U41259 (N_41259,N_39154,N_39975);
or U41260 (N_41260,N_36672,N_39760);
nor U41261 (N_41261,N_36133,N_36782);
xor U41262 (N_41262,N_35532,N_36952);
xor U41263 (N_41263,N_37642,N_39503);
or U41264 (N_41264,N_35733,N_35341);
and U41265 (N_41265,N_37918,N_35838);
and U41266 (N_41266,N_38442,N_38717);
and U41267 (N_41267,N_35989,N_36147);
nand U41268 (N_41268,N_36117,N_36180);
and U41269 (N_41269,N_37092,N_35282);
nor U41270 (N_41270,N_39884,N_38745);
or U41271 (N_41271,N_39697,N_36485);
and U41272 (N_41272,N_39422,N_36049);
xnor U41273 (N_41273,N_39600,N_37410);
xnor U41274 (N_41274,N_37356,N_38444);
and U41275 (N_41275,N_36044,N_37768);
or U41276 (N_41276,N_38065,N_36683);
xnor U41277 (N_41277,N_39447,N_39761);
nand U41278 (N_41278,N_39475,N_35725);
xor U41279 (N_41279,N_36961,N_36581);
and U41280 (N_41280,N_38440,N_37685);
or U41281 (N_41281,N_37049,N_35853);
nor U41282 (N_41282,N_39614,N_37725);
xnor U41283 (N_41283,N_38045,N_36889);
xor U41284 (N_41284,N_37099,N_37896);
nor U41285 (N_41285,N_39207,N_39577);
and U41286 (N_41286,N_35927,N_35617);
or U41287 (N_41287,N_39352,N_39702);
and U41288 (N_41288,N_39423,N_37279);
and U41289 (N_41289,N_36488,N_39532);
and U41290 (N_41290,N_35017,N_39686);
nand U41291 (N_41291,N_35590,N_37714);
nand U41292 (N_41292,N_39250,N_38844);
nand U41293 (N_41293,N_39102,N_38060);
xnor U41294 (N_41294,N_37006,N_38043);
and U41295 (N_41295,N_37727,N_39306);
nor U41296 (N_41296,N_39647,N_39555);
xnor U41297 (N_41297,N_36893,N_38729);
nand U41298 (N_41298,N_38753,N_38877);
nor U41299 (N_41299,N_35174,N_37022);
xnor U41300 (N_41300,N_37338,N_36894);
and U41301 (N_41301,N_38763,N_39507);
nor U41302 (N_41302,N_36558,N_35497);
or U41303 (N_41303,N_36005,N_35035);
or U41304 (N_41304,N_39125,N_38800);
and U41305 (N_41305,N_36051,N_38584);
and U41306 (N_41306,N_35769,N_37057);
xnor U41307 (N_41307,N_39260,N_35294);
xnor U41308 (N_41308,N_36483,N_37872);
or U41309 (N_41309,N_37611,N_37155);
xor U41310 (N_41310,N_39546,N_39140);
and U41311 (N_41311,N_39005,N_39277);
and U41312 (N_41312,N_35426,N_39090);
or U41313 (N_41313,N_35641,N_39769);
xor U41314 (N_41314,N_35826,N_35065);
nor U41315 (N_41315,N_36320,N_36848);
and U41316 (N_41316,N_39295,N_39198);
or U41317 (N_41317,N_37659,N_38847);
nor U41318 (N_41318,N_37867,N_37379);
or U41319 (N_41319,N_35681,N_39653);
xor U41320 (N_41320,N_36295,N_36994);
xor U41321 (N_41321,N_39796,N_38185);
or U41322 (N_41322,N_37235,N_35021);
nor U41323 (N_41323,N_35844,N_36353);
or U41324 (N_41324,N_39940,N_39159);
xnor U41325 (N_41325,N_37701,N_36472);
nand U41326 (N_41326,N_36314,N_38957);
nand U41327 (N_41327,N_35202,N_39996);
xnor U41328 (N_41328,N_39899,N_39889);
nor U41329 (N_41329,N_38351,N_39222);
nor U41330 (N_41330,N_37839,N_36878);
nand U41331 (N_41331,N_36023,N_37084);
and U41332 (N_41332,N_36524,N_37815);
nor U41333 (N_41333,N_39141,N_37792);
nand U41334 (N_41334,N_35522,N_39742);
nand U41335 (N_41335,N_35146,N_37439);
and U41336 (N_41336,N_36242,N_35727);
and U41337 (N_41337,N_35548,N_37061);
xor U41338 (N_41338,N_37461,N_39585);
and U41339 (N_41339,N_39072,N_39213);
or U41340 (N_41340,N_35812,N_36464);
nand U41341 (N_41341,N_36173,N_38080);
xor U41342 (N_41342,N_35547,N_37208);
and U41343 (N_41343,N_36113,N_38810);
nand U41344 (N_41344,N_37848,N_38267);
nand U41345 (N_41345,N_36789,N_36655);
or U41346 (N_41346,N_35154,N_35239);
and U41347 (N_41347,N_37526,N_39458);
nor U41348 (N_41348,N_37624,N_37026);
nand U41349 (N_41349,N_36383,N_35785);
xor U41350 (N_41350,N_35703,N_39380);
and U41351 (N_41351,N_39201,N_39913);
and U41352 (N_41352,N_36228,N_35779);
xor U41353 (N_41353,N_36825,N_36088);
nand U41354 (N_41354,N_38223,N_36544);
xor U41355 (N_41355,N_39110,N_37460);
nand U41356 (N_41356,N_38076,N_38194);
nor U41357 (N_41357,N_35848,N_35775);
nand U41358 (N_41358,N_38767,N_39160);
xnor U41359 (N_41359,N_37405,N_37951);
and U41360 (N_41360,N_35879,N_36926);
nand U41361 (N_41361,N_35997,N_39944);
nand U41362 (N_41362,N_35119,N_37108);
and U41363 (N_41363,N_38622,N_39233);
nand U41364 (N_41364,N_36008,N_39297);
and U41365 (N_41365,N_35740,N_38491);
nor U41366 (N_41366,N_35661,N_35402);
nand U41367 (N_41367,N_38827,N_38244);
nor U41368 (N_41368,N_38061,N_38531);
nor U41369 (N_41369,N_39060,N_37434);
or U41370 (N_41370,N_38928,N_37541);
nand U41371 (N_41371,N_36273,N_39715);
and U41372 (N_41372,N_39463,N_39971);
xor U41373 (N_41373,N_35275,N_36028);
xnor U41374 (N_41374,N_37774,N_39992);
xnor U41375 (N_41375,N_38208,N_38786);
nor U41376 (N_41376,N_37213,N_37304);
nand U41377 (N_41377,N_38498,N_36297);
nand U41378 (N_41378,N_37322,N_36367);
nand U41379 (N_41379,N_36379,N_37474);
nor U41380 (N_41380,N_39241,N_38527);
nor U41381 (N_41381,N_37032,N_36216);
or U41382 (N_41382,N_38982,N_36017);
xnor U41383 (N_41383,N_39182,N_35876);
nand U41384 (N_41384,N_38044,N_35632);
nor U41385 (N_41385,N_36843,N_39373);
and U41386 (N_41386,N_39819,N_35258);
nand U41387 (N_41387,N_35741,N_35373);
and U41388 (N_41388,N_35317,N_37704);
nand U41389 (N_41389,N_39793,N_38651);
and U41390 (N_41390,N_39581,N_36127);
nand U41391 (N_41391,N_36816,N_38779);
nor U41392 (N_41392,N_36702,N_37592);
nor U41393 (N_41393,N_37250,N_38103);
xor U41394 (N_41394,N_37278,N_39355);
and U41395 (N_41395,N_39771,N_39844);
nor U41396 (N_41396,N_37700,N_36210);
or U41397 (N_41397,N_39911,N_37429);
nor U41398 (N_41398,N_39611,N_37832);
or U41399 (N_41399,N_38127,N_37557);
xor U41400 (N_41400,N_35594,N_36813);
nor U41401 (N_41401,N_38029,N_39957);
nand U41402 (N_41402,N_37325,N_37755);
nand U41403 (N_41403,N_39314,N_37699);
or U41404 (N_41404,N_38704,N_35004);
nor U41405 (N_41405,N_38160,N_36476);
xnor U41406 (N_41406,N_37301,N_39396);
or U41407 (N_41407,N_37294,N_37245);
nand U41408 (N_41408,N_36422,N_36144);
nand U41409 (N_41409,N_37562,N_37919);
nor U41410 (N_41410,N_35889,N_36150);
nor U41411 (N_41411,N_36421,N_39754);
xor U41412 (N_41412,N_36119,N_39360);
nor U41413 (N_41413,N_39738,N_36326);
or U41414 (N_41414,N_36204,N_38418);
or U41415 (N_41415,N_38270,N_39138);
nor U41416 (N_41416,N_36985,N_38705);
nand U41417 (N_41417,N_37898,N_39631);
and U41418 (N_41418,N_35291,N_37973);
nand U41419 (N_41419,N_38214,N_36886);
or U41420 (N_41420,N_35066,N_38483);
or U41421 (N_41421,N_39307,N_35342);
nand U41422 (N_41422,N_38013,N_37477);
nand U41423 (N_41423,N_35030,N_39646);
xor U41424 (N_41424,N_35560,N_37276);
xnor U41425 (N_41425,N_35399,N_39937);
and U41426 (N_41426,N_38816,N_38229);
and U41427 (N_41427,N_36020,N_37790);
nand U41428 (N_41428,N_36640,N_37373);
nand U41429 (N_41429,N_37054,N_39073);
or U41430 (N_41430,N_39506,N_36285);
or U41431 (N_41431,N_35008,N_39606);
nor U41432 (N_41432,N_38396,N_37349);
xor U41433 (N_41433,N_35577,N_35205);
nand U41434 (N_41434,N_38885,N_38752);
and U41435 (N_41435,N_37788,N_39365);
and U41436 (N_41436,N_36513,N_38656);
xor U41437 (N_41437,N_35858,N_37451);
xnor U41438 (N_41438,N_38631,N_39255);
nor U41439 (N_41439,N_35964,N_39471);
or U41440 (N_41440,N_35992,N_37305);
and U41441 (N_41441,N_37866,N_35744);
nand U41442 (N_41442,N_39114,N_36446);
nor U41443 (N_41443,N_39750,N_39680);
nor U41444 (N_41444,N_39202,N_38542);
xnor U41445 (N_41445,N_39328,N_38050);
xnor U41446 (N_41446,N_36907,N_36065);
xnor U41447 (N_41447,N_37585,N_36984);
and U41448 (N_41448,N_35941,N_36646);
nor U41449 (N_41449,N_35598,N_37741);
nand U41450 (N_41450,N_38933,N_39570);
xnor U41451 (N_41451,N_37877,N_35942);
nand U41452 (N_41452,N_35933,N_39777);
nor U41453 (N_41453,N_36033,N_36137);
nand U41454 (N_41454,N_37089,N_38922);
or U41455 (N_41455,N_38822,N_38202);
or U41456 (N_41456,N_35052,N_38501);
and U41457 (N_41457,N_37012,N_35523);
nor U41458 (N_41458,N_36947,N_38386);
and U41459 (N_41459,N_35226,N_37720);
and U41460 (N_41460,N_35274,N_39412);
nor U41461 (N_41461,N_36310,N_39410);
nand U41462 (N_41462,N_36860,N_35629);
and U41463 (N_41463,N_39364,N_37091);
nand U41464 (N_41464,N_35194,N_35656);
xnor U41465 (N_41465,N_35735,N_37011);
and U41466 (N_41466,N_35422,N_35998);
nor U41467 (N_41467,N_36903,N_39340);
nand U41468 (N_41468,N_37214,N_38589);
or U41469 (N_41469,N_38986,N_39158);
and U41470 (N_41470,N_38614,N_37025);
and U41471 (N_41471,N_35955,N_35145);
or U41472 (N_41472,N_38110,N_39544);
nor U41473 (N_41473,N_37126,N_35396);
or U41474 (N_41474,N_39505,N_39752);
nand U41475 (N_41475,N_38818,N_36126);
and U41476 (N_41476,N_37230,N_39509);
nor U41477 (N_41477,N_36647,N_35179);
and U41478 (N_41478,N_39636,N_37123);
nor U41479 (N_41479,N_38432,N_37826);
or U41480 (N_41480,N_38967,N_39347);
and U41481 (N_41481,N_37060,N_36942);
nor U41482 (N_41482,N_35423,N_37290);
xnor U41483 (N_41483,N_36212,N_38521);
or U41484 (N_41484,N_35847,N_38565);
xor U41485 (N_41485,N_36627,N_37936);
nand U41486 (N_41486,N_38047,N_39455);
or U41487 (N_41487,N_36913,N_37516);
nor U41488 (N_41488,N_38547,N_39283);
and U41489 (N_41489,N_37969,N_39082);
nor U41490 (N_41490,N_37309,N_38012);
and U41491 (N_41491,N_37960,N_37447);
and U41492 (N_41492,N_37502,N_35585);
and U41493 (N_41493,N_36512,N_38147);
or U41494 (N_41494,N_36218,N_38927);
or U41495 (N_41495,N_37716,N_38138);
and U41496 (N_41496,N_39938,N_38698);
nand U41497 (N_41497,N_35178,N_39865);
and U41498 (N_41498,N_39590,N_36497);
nor U41499 (N_41499,N_36908,N_36923);
xor U41500 (N_41500,N_38423,N_37308);
nor U41501 (N_41501,N_36318,N_38294);
xor U41502 (N_41502,N_38551,N_37247);
nor U41503 (N_41503,N_35328,N_36356);
nor U41504 (N_41504,N_36220,N_36257);
or U41505 (N_41505,N_36030,N_37724);
nor U41506 (N_41506,N_37566,N_37740);
and U41507 (N_41507,N_38360,N_37039);
and U41508 (N_41508,N_38992,N_39866);
nand U41509 (N_41509,N_35237,N_36859);
and U41510 (N_41510,N_35667,N_38900);
nand U41511 (N_41511,N_35283,N_38055);
nand U41512 (N_41512,N_36736,N_35277);
xnor U41513 (N_41513,N_38349,N_35189);
or U41514 (N_41514,N_36246,N_36362);
xor U41515 (N_41515,N_39964,N_38381);
and U41516 (N_41516,N_39895,N_39770);
nand U41517 (N_41517,N_35209,N_39324);
nor U41518 (N_41518,N_36800,N_37377);
xnor U41519 (N_41519,N_35873,N_39319);
nor U41520 (N_41520,N_39006,N_35319);
or U41521 (N_41521,N_36963,N_37639);
nand U41522 (N_41522,N_35494,N_35888);
xor U41523 (N_41523,N_37241,N_37251);
and U41524 (N_41524,N_35256,N_37580);
nor U41525 (N_41525,N_37414,N_39498);
nand U41526 (N_41526,N_37854,N_35697);
nand U41527 (N_41527,N_39801,N_35281);
nor U41528 (N_41528,N_39504,N_39368);
nand U41529 (N_41529,N_37096,N_35881);
xnor U41530 (N_41530,N_36429,N_39736);
nor U41531 (N_41531,N_36667,N_36822);
xor U41532 (N_41532,N_39264,N_35541);
and U41533 (N_41533,N_38522,N_39530);
xor U41534 (N_41534,N_38112,N_37803);
nand U41535 (N_41535,N_38370,N_37575);
or U41536 (N_41536,N_36876,N_36135);
and U41537 (N_41537,N_38152,N_38116);
nand U41538 (N_41538,N_36458,N_38430);
nor U41539 (N_41539,N_39481,N_35668);
and U41540 (N_41540,N_37528,N_36708);
nand U41541 (N_41541,N_38332,N_35578);
nor U41542 (N_41542,N_36371,N_39022);
xor U41543 (N_41543,N_36099,N_38748);
nand U41544 (N_41544,N_35957,N_35920);
xnor U41545 (N_41545,N_38145,N_38056);
nor U41546 (N_41546,N_39230,N_37812);
and U41547 (N_41547,N_35242,N_39508);
nand U41548 (N_41548,N_37161,N_38981);
and U41549 (N_41549,N_39858,N_36784);
or U41550 (N_41550,N_39602,N_35963);
xor U41551 (N_41551,N_39274,N_35296);
nor U41552 (N_41552,N_35683,N_37712);
nor U41553 (N_41553,N_38654,N_36765);
or U41554 (N_41554,N_35128,N_37370);
nor U41555 (N_41555,N_36477,N_38002);
nor U41556 (N_41556,N_39087,N_36329);
or U41557 (N_41557,N_35102,N_37565);
nor U41558 (N_41558,N_38526,N_36351);
and U41559 (N_41559,N_37689,N_38673);
or U41560 (N_41560,N_37765,N_35605);
nor U41561 (N_41561,N_35855,N_38769);
nor U41562 (N_41562,N_35414,N_39078);
nor U41563 (N_41563,N_36188,N_35761);
nand U41564 (N_41564,N_35495,N_35821);
nor U41565 (N_41565,N_39517,N_37616);
or U41566 (N_41566,N_37706,N_37396);
nor U41567 (N_41567,N_37884,N_35651);
and U41568 (N_41568,N_39930,N_38268);
nor U41569 (N_41569,N_36015,N_36551);
or U41570 (N_41570,N_39598,N_36585);
xor U41571 (N_41571,N_38976,N_39868);
xor U41572 (N_41572,N_38486,N_35073);
nor U41573 (N_41573,N_37109,N_35266);
nand U41574 (N_41574,N_38916,N_35674);
xnor U41575 (N_41575,N_35857,N_35159);
nor U41576 (N_41576,N_36007,N_35648);
xnor U41577 (N_41577,N_38997,N_39156);
xnor U41578 (N_41578,N_38184,N_37465);
or U41579 (N_41579,N_38203,N_39816);
and U41580 (N_41580,N_39642,N_35764);
nand U41581 (N_41581,N_39566,N_37386);
xnor U41582 (N_41582,N_36751,N_37976);
nor U41583 (N_41583,N_37932,N_36879);
nor U41584 (N_41584,N_37042,N_35221);
nor U41585 (N_41585,N_36866,N_35870);
and U41586 (N_41586,N_39161,N_35325);
nor U41587 (N_41587,N_36194,N_35445);
nor U41588 (N_41588,N_35356,N_37966);
or U41589 (N_41589,N_39547,N_39275);
nor U41590 (N_41590,N_36628,N_39689);
nor U41591 (N_41591,N_36561,N_36950);
and U41592 (N_41592,N_36291,N_37558);
xor U41593 (N_41593,N_38696,N_35576);
nor U41594 (N_41594,N_37267,N_38422);
nand U41595 (N_41595,N_38273,N_35805);
and U41596 (N_41596,N_37248,N_35700);
nor U41597 (N_41597,N_35565,N_37767);
or U41598 (N_41598,N_39486,N_39081);
xor U41599 (N_41599,N_38664,N_35994);
and U41600 (N_41600,N_36701,N_37045);
or U41601 (N_41601,N_37961,N_37841);
and U41602 (N_41602,N_39639,N_36091);
and U41603 (N_41603,N_39137,N_37486);
xnor U41604 (N_41604,N_35999,N_38609);
nor U41605 (N_41605,N_39315,N_35381);
and U41606 (N_41606,N_39961,N_38467);
and U41607 (N_41607,N_36829,N_35646);
nand U41608 (N_41608,N_36861,N_38003);
or U41609 (N_41609,N_38618,N_36240);
xor U41610 (N_41610,N_35272,N_39227);
xnor U41611 (N_41611,N_37080,N_37009);
and U41612 (N_41612,N_37709,N_39583);
nor U41613 (N_41613,N_36423,N_38301);
and U41614 (N_41614,N_37892,N_36760);
and U41615 (N_41615,N_39253,N_36334);
xnor U41616 (N_41616,N_35016,N_37993);
nand U41617 (N_41617,N_39390,N_38679);
nor U41618 (N_41618,N_38118,N_37764);
nor U41619 (N_41619,N_37215,N_35919);
and U41620 (N_41620,N_37876,N_36101);
nor U41621 (N_41621,N_36593,N_39386);
nor U41622 (N_41622,N_38824,N_36193);
or U41623 (N_41623,N_37152,N_39416);
and U41624 (N_41624,N_37270,N_36621);
and U41625 (N_41625,N_37897,N_35113);
nand U41626 (N_41626,N_39413,N_36174);
xnor U41627 (N_41627,N_38275,N_37264);
or U41628 (N_41628,N_37067,N_35458);
nor U41629 (N_41629,N_35081,N_38336);
nand U41630 (N_41630,N_38239,N_38659);
nand U41631 (N_41631,N_36081,N_35225);
and U41632 (N_41632,N_36232,N_39960);
nor U41633 (N_41633,N_36653,N_35658);
nand U41634 (N_41634,N_39559,N_38382);
nor U41635 (N_41635,N_37364,N_37609);
nor U41636 (N_41636,N_39437,N_36968);
nand U41637 (N_41637,N_36944,N_39648);
nor U41638 (N_41638,N_39058,N_39626);
or U41639 (N_41639,N_37145,N_37825);
nand U41640 (N_41640,N_38314,N_36797);
nor U41641 (N_41641,N_38470,N_36698);
or U41642 (N_41642,N_37351,N_39950);
nand U41643 (N_41643,N_37632,N_39231);
nand U41644 (N_41644,N_37101,N_36954);
xnor U41645 (N_41645,N_38902,N_36237);
or U41646 (N_41646,N_37994,N_35107);
xor U41647 (N_41647,N_39361,N_37907);
nand U41648 (N_41648,N_37517,N_38453);
and U41649 (N_41649,N_37037,N_37518);
or U41650 (N_41650,N_36409,N_37345);
xor U41651 (N_41651,N_36617,N_37088);
xnor U41652 (N_41652,N_36395,N_35774);
nor U41653 (N_41653,N_39451,N_38421);
xnor U41654 (N_41654,N_36635,N_35425);
xor U41655 (N_41655,N_38908,N_39394);
nand U41656 (N_41656,N_39753,N_36011);
nor U41657 (N_41657,N_37649,N_37519);
nand U41658 (N_41658,N_39074,N_38235);
and U41659 (N_41659,N_39330,N_36846);
and U41660 (N_41660,N_39849,N_38549);
or U41661 (N_41661,N_37710,N_39016);
nand U41662 (N_41662,N_38571,N_38718);
nand U41663 (N_41663,N_36013,N_35514);
nand U41664 (N_41664,N_35477,N_36009);
nand U41665 (N_41665,N_35125,N_38774);
xnor U41666 (N_41666,N_36388,N_37889);
xor U41667 (N_41667,N_35453,N_39716);
and U41668 (N_41668,N_39008,N_39972);
and U41669 (N_41669,N_37391,N_39698);
xor U41670 (N_41670,N_39765,N_39088);
or U41671 (N_41671,N_35056,N_36259);
xor U41672 (N_41672,N_39171,N_36506);
nor U41673 (N_41673,N_39589,N_39193);
nand U41674 (N_41674,N_38317,N_36469);
xnor U41675 (N_41675,N_36128,N_36247);
nand U41676 (N_41676,N_39883,N_35912);
xor U41677 (N_41677,N_37169,N_35882);
and U41678 (N_41678,N_39276,N_37845);
and U41679 (N_41679,N_38680,N_35850);
nor U41680 (N_41680,N_36190,N_39335);
nor U41681 (N_41681,N_36771,N_35230);
nand U41682 (N_41682,N_36157,N_39263);
nor U41683 (N_41683,N_35526,N_36587);
nand U41684 (N_41684,N_36168,N_35712);
xor U41685 (N_41685,N_37673,N_39643);
nor U41686 (N_41686,N_39168,N_36641);
and U41687 (N_41687,N_38841,N_35872);
xor U41688 (N_41688,N_35465,N_39359);
nand U41689 (N_41689,N_36875,N_39775);
nand U41690 (N_41690,N_37303,N_37776);
nor U41691 (N_41691,N_36480,N_35147);
nand U41692 (N_41692,N_35334,N_36925);
or U41693 (N_41693,N_35362,N_35120);
nor U41694 (N_41694,N_37983,N_38297);
nand U41695 (N_41695,N_36453,N_39951);
xnor U41696 (N_41696,N_36121,N_38438);
or U41697 (N_41697,N_37494,N_35767);
or U41698 (N_41698,N_37638,N_37326);
or U41699 (N_41699,N_35265,N_38228);
xor U41700 (N_41700,N_36805,N_35806);
xnor U41701 (N_41701,N_38600,N_38795);
xor U41702 (N_41702,N_35238,N_37455);
xor U41703 (N_41703,N_35370,N_35366);
nor U41704 (N_41704,N_35476,N_39690);
nor U41705 (N_41705,N_35606,N_39385);
and U41706 (N_41706,N_39216,N_38460);
or U41707 (N_41707,N_39874,N_37497);
and U41708 (N_41708,N_36241,N_39537);
nand U41709 (N_41709,N_39786,N_37759);
or U41710 (N_41710,N_36462,N_38032);
nor U41711 (N_41711,N_37590,N_36870);
and U41712 (N_41712,N_37570,N_36083);
nor U41713 (N_41713,N_38358,N_36982);
or U41714 (N_41714,N_35759,N_36584);
nand U41715 (N_41715,N_35588,N_37253);
or U41716 (N_41716,N_39551,N_39663);
or U41717 (N_41717,N_36576,N_38009);
nand U41718 (N_41718,N_38424,N_35478);
xor U41719 (N_41719,N_39615,N_37941);
and U41720 (N_41720,N_35907,N_39730);
nor U41721 (N_41721,N_38891,N_37538);
nor U41722 (N_41722,N_39827,N_36937);
or U41723 (N_41723,N_36058,N_35192);
or U41724 (N_41724,N_38863,N_39476);
nor U41725 (N_41725,N_35015,N_35886);
and U41726 (N_41726,N_38489,N_39630);
xor U41727 (N_41727,N_37020,N_36211);
xnor U41728 (N_41728,N_37289,N_35115);
nand U41729 (N_41729,N_35488,N_36972);
xnor U41730 (N_41730,N_35657,N_37947);
xnor U41731 (N_41731,N_38437,N_38397);
nand U41732 (N_41732,N_38945,N_37068);
xnor U41733 (N_41733,N_37894,N_35106);
or U41734 (N_41734,N_38105,N_35475);
xor U41735 (N_41735,N_39718,N_39550);
nor U41736 (N_41736,N_39261,N_35642);
xnor U41737 (N_41737,N_37942,N_36010);
xor U41738 (N_41738,N_38951,N_37284);
or U41739 (N_41739,N_35103,N_38678);
nor U41740 (N_41740,N_36864,N_35343);
and U41741 (N_41741,N_38095,N_37811);
xnor U41742 (N_41742,N_38778,N_35377);
or U41743 (N_41743,N_39658,N_37579);
nor U41744 (N_41744,N_39399,N_37105);
xor U41745 (N_41745,N_38245,N_39727);
nand U41746 (N_41746,N_35455,N_39743);
xnor U41747 (N_41747,N_37640,N_39190);
nand U41748 (N_41748,N_37604,N_37164);
and U41749 (N_41749,N_36652,N_35732);
nor U41750 (N_41750,N_37891,N_39353);
or U41751 (N_41751,N_36906,N_39802);
nand U41752 (N_41752,N_36102,N_37957);
nor U41753 (N_41753,N_37614,N_39974);
nor U41754 (N_41754,N_37202,N_39010);
or U41755 (N_41755,N_36456,N_39790);
nand U41756 (N_41756,N_35340,N_36928);
xnor U41757 (N_41757,N_36263,N_38652);
and U41758 (N_41758,N_36642,N_36645);
nand U41759 (N_41759,N_36025,N_37195);
nor U41760 (N_41760,N_37846,N_39869);
or U41761 (N_41761,N_39461,N_39134);
xor U41762 (N_41762,N_35131,N_39374);
nor U41763 (N_41763,N_38466,N_36909);
and U41764 (N_41764,N_37511,N_35167);
xor U41765 (N_41765,N_38243,N_36292);
and U41766 (N_41766,N_37157,N_38279);
or U41767 (N_41767,N_39810,N_38719);
nand U41768 (N_41768,N_36467,N_38125);
and U41769 (N_41769,N_36281,N_36892);
and U41770 (N_41770,N_39402,N_35692);
nor U41771 (N_41771,N_37683,N_36975);
or U41772 (N_41772,N_35481,N_37822);
nand U41773 (N_41773,N_38380,N_36916);
xor U41774 (N_41774,N_39096,N_36508);
nor U41775 (N_41775,N_36598,N_38200);
and U41776 (N_41776,N_39925,N_35921);
nand U41777 (N_41777,N_37256,N_37236);
nand U41778 (N_41778,N_38836,N_37274);
nor U41779 (N_41779,N_35169,N_35364);
nand U41780 (N_41780,N_38233,N_38237);
xnor U41781 (N_41781,N_37890,N_35693);
or U41782 (N_41782,N_39061,N_39327);
and U41783 (N_41783,N_39120,N_36466);
nor U41784 (N_41784,N_37185,N_39672);
or U41785 (N_41785,N_37521,N_36895);
xor U41786 (N_41786,N_35045,N_38490);
nor U41787 (N_41787,N_39829,N_36898);
nor U41788 (N_41788,N_39826,N_38286);
xor U41789 (N_41789,N_36636,N_38324);
xnor U41790 (N_41790,N_38848,N_36804);
nor U41791 (N_41791,N_36912,N_39189);
or U41792 (N_41792,N_35280,N_36060);
or U41793 (N_41793,N_38041,N_38979);
nor U41794 (N_41794,N_36622,N_38326);
nor U41795 (N_41795,N_37595,N_38330);
and U41796 (N_41796,N_36752,N_38888);
or U41797 (N_41797,N_39795,N_36373);
nor U41798 (N_41798,N_38585,N_36965);
or U41799 (N_41799,N_39668,N_38710);
xor U41800 (N_41800,N_39873,N_35958);
nand U41801 (N_41801,N_35443,N_35597);
and U41802 (N_41802,N_38227,N_35264);
nor U41803 (N_41803,N_35575,N_35793);
nand U41804 (N_41804,N_39299,N_35643);
xor U41805 (N_41805,N_37085,N_36417);
and U41806 (N_41806,N_37191,N_37924);
xor U41807 (N_41807,N_35386,N_36161);
nor U41808 (N_41808,N_36063,N_35550);
or U41809 (N_41809,N_37118,N_37583);
nand U41810 (N_41810,N_36588,N_37028);
and U41811 (N_41811,N_38117,N_36484);
nand U41812 (N_41812,N_38857,N_35331);
or U41813 (N_41813,N_37296,N_37257);
nor U41814 (N_41814,N_39220,N_36546);
xnor U41815 (N_41815,N_35690,N_36413);
nor U41816 (N_41816,N_36564,N_35267);
and U41817 (N_41817,N_37982,N_38798);
or U41818 (N_41818,N_39768,N_35860);
or U41819 (N_41819,N_36704,N_37198);
nor U41820 (N_41820,N_36877,N_39908);
and U41821 (N_41821,N_37576,N_35562);
nand U41822 (N_41822,N_37482,N_37913);
or U41823 (N_41823,N_35156,N_39251);
xnor U41824 (N_41824,N_39773,N_36208);
nand U41825 (N_41825,N_37113,N_35487);
nor U41826 (N_41826,N_36550,N_39083);
nand U41827 (N_41827,N_35603,N_38595);
nor U41828 (N_41828,N_39223,N_37705);
nand U41829 (N_41829,N_39652,N_36594);
and U41830 (N_41830,N_39627,N_38524);
xnor U41831 (N_41831,N_38411,N_37682);
xnor U41832 (N_41832,N_37864,N_37260);
and U41833 (N_41833,N_38998,N_37670);
nor U41834 (N_41834,N_38078,N_36826);
and U41835 (N_41835,N_37787,N_36230);
or U41836 (N_41836,N_36479,N_39281);
nand U41837 (N_41837,N_37643,N_35612);
and U41838 (N_41838,N_38890,N_37342);
xor U41839 (N_41839,N_35802,N_38263);
xnor U41840 (N_41840,N_35324,N_38573);
or U41841 (N_41841,N_35408,N_39166);
nor U41842 (N_41842,N_38546,N_36590);
xnor U41843 (N_41843,N_38107,N_37209);
xor U41844 (N_41844,N_38532,N_35245);
nor U41845 (N_41845,N_37380,N_38670);
and U41846 (N_41846,N_38231,N_39942);
xnor U41847 (N_41847,N_39799,N_39080);
and U41848 (N_41848,N_36074,N_38850);
or U41849 (N_41849,N_35090,N_39215);
nor U41850 (N_41850,N_36790,N_38613);
nor U41851 (N_41851,N_38247,N_37875);
xnor U41852 (N_41852,N_35398,N_36412);
or U41853 (N_41853,N_39798,N_37824);
nor U41854 (N_41854,N_36835,N_36235);
nand U41855 (N_41855,N_35709,N_35924);
or U41856 (N_41856,N_35593,N_39405);
nand U41857 (N_41857,N_37730,N_38099);
and U41858 (N_41858,N_36688,N_39997);
xor U41859 (N_41859,N_36391,N_39098);
nor U41860 (N_41860,N_39366,N_35841);
xnor U41861 (N_41861,N_37840,N_36844);
xnor U41862 (N_41862,N_36130,N_36707);
nand U41863 (N_41863,N_37457,N_35659);
or U41864 (N_41864,N_35553,N_39804);
nand U41865 (N_41865,N_35031,N_36967);
or U41866 (N_41866,N_37715,N_37135);
xor U41867 (N_41867,N_35054,N_37332);
xor U41868 (N_41868,N_35403,N_37232);
nor U41869 (N_41869,N_36042,N_36482);
xor U41870 (N_41870,N_37340,N_37561);
or U41871 (N_41871,N_38783,N_35069);
nand U41872 (N_41872,N_36443,N_37865);
or U41873 (N_41873,N_35980,N_35837);
nor U41874 (N_41874,N_35815,N_39240);
and U41875 (N_41875,N_37582,N_37402);
nand U41876 (N_41876,N_39954,N_38248);
nand U41877 (N_41877,N_38821,N_39528);
nor U41878 (N_41878,N_36270,N_36311);
or U41879 (N_41879,N_38007,N_39717);
nor U41880 (N_41880,N_36478,N_37199);
nand U41881 (N_41881,N_38689,N_38480);
nand U41882 (N_41882,N_39470,N_36977);
or U41883 (N_41883,N_37863,N_38161);
nor U41884 (N_41884,N_37971,N_35437);
xnor U41885 (N_41885,N_39268,N_35442);
or U41886 (N_41886,N_39764,N_35619);
nand U41887 (N_41887,N_39758,N_35707);
xor U41888 (N_41888,N_38889,N_35318);
xor U41889 (N_41889,N_37287,N_37421);
nor U41890 (N_41890,N_35930,N_36420);
nor U41891 (N_41891,N_36400,N_36415);
or U41892 (N_41892,N_36236,N_39953);
nand U41893 (N_41893,N_37512,N_36750);
and U41894 (N_41894,N_38504,N_37281);
xnor U41895 (N_41895,N_35116,N_39225);
nand U41896 (N_41896,N_39448,N_38181);
nand U41897 (N_41897,N_39389,N_36115);
nand U41898 (N_41898,N_37005,N_35694);
nand U41899 (N_41899,N_37525,N_38474);
nor U41900 (N_41900,N_37058,N_35766);
nor U41901 (N_41901,N_35579,N_35121);
and U41902 (N_41902,N_36669,N_39531);
and U41903 (N_41903,N_37760,N_38871);
or U41904 (N_41904,N_39235,N_38964);
nand U41905 (N_41905,N_39596,N_35788);
or U41906 (N_41906,N_36980,N_35148);
nor U41907 (N_41907,N_36433,N_35040);
nand U41908 (N_41908,N_37480,N_36625);
xnor U41909 (N_41909,N_38073,N_37879);
nor U41910 (N_41910,N_38001,N_38833);
and U41911 (N_41911,N_36219,N_35776);
nand U41912 (N_41912,N_39497,N_38269);
xor U41913 (N_41913,N_39124,N_35198);
and U41914 (N_41914,N_39209,N_38733);
xnor U41915 (N_41915,N_39094,N_36560);
xnor U41916 (N_41916,N_38298,N_35952);
nand U41917 (N_41917,N_39847,N_38918);
nand U41918 (N_41918,N_39684,N_36155);
and U41919 (N_41919,N_38676,N_35736);
and U41920 (N_41920,N_36521,N_36992);
xnor U41921 (N_41921,N_39446,N_39983);
nor U41922 (N_41922,N_39927,N_38602);
xnor U41923 (N_41923,N_37016,N_39987);
xor U41924 (N_41924,N_35621,N_37149);
or U41925 (N_41925,N_36493,N_35158);
nor U41926 (N_41926,N_36523,N_38488);
and U41927 (N_41927,N_36445,N_36159);
nor U41928 (N_41928,N_35415,N_37423);
nand U41929 (N_41929,N_36957,N_37855);
nor U41930 (N_41930,N_37895,N_37347);
xnor U41931 (N_41931,N_37495,N_38346);
nand U41932 (N_41932,N_39926,N_38715);
nand U41933 (N_41933,N_35730,N_39326);
xor U41934 (N_41934,N_35696,N_35337);
and U41935 (N_41935,N_35416,N_37071);
nand U41936 (N_41936,N_38735,N_35572);
or U41937 (N_41937,N_37331,N_36665);
nor U41938 (N_41938,N_36431,N_36901);
nor U41939 (N_41939,N_39025,N_39298);
nand U41940 (N_41940,N_39468,N_36104);
nor U41941 (N_41941,N_38665,N_36419);
nand U41942 (N_41942,N_36591,N_39541);
xor U41943 (N_41943,N_35417,N_39813);
and U41944 (N_41944,N_36573,N_38548);
or U41945 (N_41945,N_39449,N_39694);
or U41946 (N_41946,N_39877,N_35995);
xnor U41947 (N_41947,N_39807,N_39381);
nand U41948 (N_41948,N_39977,N_39174);
or U41949 (N_41949,N_37344,N_39712);
or U41950 (N_41950,N_36767,N_39520);
and U41951 (N_41951,N_39845,N_35549);
nand U41952 (N_41952,N_37464,N_39605);
or U41953 (N_41953,N_39935,N_38775);
or U41954 (N_41954,N_36372,N_37036);
or U41955 (N_41955,N_39988,N_39332);
or U41956 (N_41956,N_38564,N_37878);
nor U41957 (N_41957,N_35875,N_38478);
nand U41958 (N_41958,N_36651,N_35521);
or U41959 (N_41959,N_36849,N_37979);
xor U41960 (N_41960,N_35041,N_36385);
nor U41961 (N_41961,N_37075,N_36350);
xnor U41962 (N_41962,N_35050,N_35241);
nand U41963 (N_41963,N_36287,N_35624);
nand U41964 (N_41964,N_36302,N_39177);
xnor U41965 (N_41965,N_37738,N_37612);
or U41966 (N_41966,N_35063,N_38568);
nor U41967 (N_41967,N_35227,N_35604);
and U41968 (N_41968,N_37124,N_36059);
or U41969 (N_41969,N_37950,N_39591);
xor U41970 (N_41970,N_39973,N_39592);
xor U41971 (N_41971,N_38256,N_36397);
nand U41972 (N_41972,N_39511,N_38934);
and U41973 (N_41973,N_35799,N_36644);
or U41974 (N_41974,N_35078,N_35210);
nand U41975 (N_41975,N_35768,N_39050);
nor U41976 (N_41976,N_35166,N_35297);
xnor U41977 (N_41977,N_37203,N_37601);
nand U41978 (N_41978,N_35321,N_38731);
nand U41979 (N_41979,N_35934,N_37187);
xnor U41980 (N_41980,N_38737,N_36405);
xor U41981 (N_41981,N_38724,N_36195);
nand U41982 (N_41982,N_35085,N_38535);
or U41983 (N_41983,N_39905,N_38407);
xor U41984 (N_41984,N_39682,N_39049);
and U41985 (N_41985,N_36178,N_37211);
and U41986 (N_41986,N_39922,N_39853);
or U41987 (N_41987,N_37507,N_38220);
xnor U41988 (N_41988,N_38051,N_35252);
or U41989 (N_41989,N_35243,N_35711);
and U41990 (N_41990,N_38791,N_38188);
nand U41991 (N_41991,N_39084,N_37341);
and U41992 (N_41992,N_38635,N_36027);
and U41993 (N_41993,N_36106,N_38412);
xnor U41994 (N_41994,N_35003,N_37220);
nor U41995 (N_41995,N_35728,N_35392);
xor U41996 (N_41996,N_39239,N_37769);
and U41997 (N_41997,N_35320,N_38024);
nor U41998 (N_41998,N_38768,N_39524);
or U41999 (N_41999,N_36239,N_35299);
xor U42000 (N_42000,N_37023,N_38959);
or U42001 (N_42001,N_36553,N_39628);
nand U42002 (N_42002,N_36357,N_35678);
and U42003 (N_42003,N_37130,N_35223);
nand U42004 (N_42004,N_36738,N_37323);
xnor U42005 (N_42005,N_37559,N_38389);
xor U42006 (N_42006,N_38259,N_36605);
and U42007 (N_42007,N_39014,N_38626);
xor U42008 (N_42008,N_39751,N_37509);
xnor U42009 (N_42009,N_35718,N_35906);
nand U42010 (N_42010,N_39009,N_37393);
or U42011 (N_42011,N_37295,N_35055);
and U42012 (N_42012,N_39409,N_38868);
nand U42013 (N_42013,N_38058,N_38280);
or U42014 (N_42014,N_37282,N_36639);
nor U42015 (N_42015,N_35923,N_36499);
xnor U42016 (N_42016,N_37004,N_38304);
xor U42017 (N_42017,N_35448,N_39291);
or U42018 (N_42018,N_39835,N_38131);
xnor U42019 (N_42019,N_35566,N_37383);
nand U42020 (N_42020,N_38655,N_37019);
xor U42021 (N_42021,N_37617,N_38016);
and U42022 (N_42022,N_37757,N_36821);
and U42023 (N_42023,N_37633,N_36731);
nand U42024 (N_42024,N_36389,N_37606);
nand U42025 (N_42025,N_39789,N_35044);
and U42026 (N_42026,N_36267,N_38156);
nor U42027 (N_42027,N_35332,N_36787);
xor U42028 (N_42028,N_39621,N_38963);
and U42029 (N_42029,N_38492,N_39741);
xnor U42030 (N_42030,N_38158,N_35468);
and U42031 (N_42031,N_37813,N_37778);
or U42032 (N_42032,N_37041,N_35141);
and U42033 (N_42033,N_38884,N_37903);
and U42034 (N_42034,N_36806,N_38143);
nand U42035 (N_42035,N_35460,N_39534);
nand U42036 (N_42036,N_38258,N_38173);
and U42037 (N_42037,N_39573,N_38598);
nor U42038 (N_42038,N_38980,N_39491);
and U42039 (N_42039,N_37791,N_37603);
nor U42040 (N_42040,N_38428,N_36705);
or U42041 (N_42041,N_37674,N_35413);
or U42042 (N_42042,N_35782,N_39226);
or U42043 (N_42043,N_39522,N_35714);
or U42044 (N_42044,N_37548,N_36960);
nand U42045 (N_42045,N_38876,N_39545);
and U42046 (N_42046,N_36450,N_36470);
or U42047 (N_42047,N_35856,N_37540);
and U42048 (N_42048,N_39345,N_35246);
nand U42049 (N_42049,N_36359,N_39483);
xor U42050 (N_42050,N_37908,N_39949);
nand U42051 (N_42051,N_38792,N_38436);
and U42052 (N_42052,N_39984,N_36637);
xor U42053 (N_42053,N_39993,N_35688);
nand U42054 (N_42054,N_39200,N_39678);
xnor U42055 (N_42055,N_36724,N_39208);
and U42056 (N_42056,N_36854,N_38812);
xnor U42057 (N_42057,N_38781,N_35689);
xor U42058 (N_42058,N_37353,N_38852);
and U42059 (N_42059,N_37394,N_38284);
and U42060 (N_42060,N_35127,N_39571);
nand U42061 (N_42061,N_39341,N_38720);
or U42062 (N_42062,N_37398,N_36284);
nand U42063 (N_42063,N_37687,N_38085);
nor U42064 (N_42064,N_39976,N_35438);
xor U42065 (N_42065,N_37300,N_36046);
xor U42066 (N_42066,N_38120,N_39635);
nor U42067 (N_42067,N_37352,N_35705);
or U42068 (N_42068,N_35638,N_36563);
and U42069 (N_42069,N_37210,N_37711);
or U42070 (N_42070,N_39053,N_36111);
and U42071 (N_42071,N_39267,N_35093);
nand U42072 (N_42072,N_38367,N_39708);
and U42073 (N_42073,N_36171,N_37717);
xor U42074 (N_42074,N_36987,N_38650);
nor U42075 (N_42075,N_35791,N_35424);
nor U42076 (N_42076,N_35909,N_38191);
nor U42077 (N_42077,N_37621,N_38759);
or U42078 (N_42078,N_36465,N_38855);
or U42079 (N_42079,N_39191,N_38662);
xor U42080 (N_42080,N_37985,N_37234);
xor U42081 (N_42081,N_37657,N_38973);
or U42082 (N_42082,N_38379,N_35072);
nand U42083 (N_42083,N_38805,N_37366);
nand U42084 (N_42084,N_38150,N_38137);
nor U42085 (N_42085,N_38799,N_35451);
and U42086 (N_42086,N_39192,N_38940);
nor U42087 (N_42087,N_37981,N_36839);
xnor U42088 (N_42088,N_39313,N_35654);
nor U42089 (N_42089,N_35473,N_37415);
xnor U42090 (N_42090,N_36927,N_35935);
nor U42091 (N_42091,N_36197,N_38605);
and U42092 (N_42092,N_39831,N_38325);
xor U42093 (N_42093,N_39197,N_38079);
or U42094 (N_42094,N_35589,N_38782);
nand U42095 (N_42095,N_38507,N_38693);
nand U42096 (N_42096,N_36618,N_36196);
and U42097 (N_42097,N_35378,N_38328);
and U42098 (N_42098,N_37940,N_37153);
or U42099 (N_42099,N_38195,N_39861);
xor U42100 (N_42100,N_36459,N_39912);
or U42101 (N_42101,N_37906,N_35359);
nand U42102 (N_42102,N_36165,N_36680);
nor U42103 (N_42103,N_35436,N_35713);
xor U42104 (N_42104,N_37350,N_38083);
and U42105 (N_42105,N_37648,N_35795);
nor U42106 (N_42106,N_38441,N_37385);
xor U42107 (N_42107,N_38930,N_38111);
xor U42108 (N_42108,N_39862,N_36352);
or U42109 (N_42109,N_39576,N_35268);
xnor U42110 (N_42110,N_37024,N_38283);
or U42111 (N_42111,N_37306,N_35908);
nor U42112 (N_42112,N_38864,N_37283);
nand U42113 (N_42113,N_38419,N_37745);
and U42114 (N_42114,N_36557,N_37034);
and U42115 (N_42115,N_38897,N_39675);
or U42116 (N_42116,N_36946,N_37173);
nand U42117 (N_42117,N_37102,N_37905);
or U42118 (N_42118,N_36838,N_35086);
nand U42119 (N_42119,N_36492,N_35491);
xor U42120 (N_42120,N_37268,N_39401);
nor U42121 (N_42121,N_35633,N_36401);
nand U42122 (N_42122,N_35884,N_36516);
nor U42123 (N_42123,N_38057,N_37881);
and U42124 (N_42124,N_37584,N_35868);
or U42125 (N_42125,N_37605,N_36836);
and U42126 (N_42126,N_39418,N_37726);
or U42127 (N_42127,N_36725,N_36116);
xnor U42128 (N_42128,N_38500,N_38327);
and U42129 (N_42129,N_36699,N_36776);
and U42130 (N_42130,N_35504,N_39042);
and U42131 (N_42131,N_36249,N_35483);
or U42132 (N_42132,N_39453,N_35457);
nand U42133 (N_42133,N_36360,N_36920);
and U42134 (N_42134,N_36427,N_39778);
and U42135 (N_42135,N_36900,N_36036);
nand U42136 (N_42136,N_36066,N_39857);
xnor U42137 (N_42137,N_37970,N_37635);
and U42138 (N_42138,N_36146,N_35551);
nand U42139 (N_42139,N_39408,N_39318);
nor U42140 (N_42140,N_36047,N_38477);
nand U42141 (N_42141,N_35082,N_35114);
and U42142 (N_42142,N_38686,N_36118);
xnor U42143 (N_42143,N_36734,N_36182);
nor U42144 (N_42144,N_36148,N_37911);
or U42145 (N_42145,N_37819,N_37520);
nor U42146 (N_42146,N_36170,N_35515);
xor U42147 (N_42147,N_36034,N_36700);
or U42148 (N_42148,N_36474,N_37662);
nor U42149 (N_42149,N_36056,N_35983);
nor U42150 (N_42150,N_38166,N_37500);
or U42151 (N_42151,N_38276,N_37335);
or U42152 (N_42152,N_38420,N_38861);
nor U42153 (N_42153,N_39870,N_38345);
nor U42154 (N_42154,N_39705,N_36964);
and U42155 (N_42155,N_35049,N_38391);
or U42156 (N_42156,N_35039,N_35787);
nor U42157 (N_42157,N_39558,N_38433);
xnor U42158 (N_42158,N_36565,N_38666);
nor U42159 (N_42159,N_35503,N_35446);
and U42160 (N_42160,N_37381,N_39362);
nand U42161 (N_42161,N_39687,N_38785);
nor U42162 (N_42162,N_38936,N_35987);
nand U42163 (N_42163,N_35715,N_37849);
or U42164 (N_42164,N_36570,N_39494);
or U42165 (N_42165,N_39121,N_38250);
nor U42166 (N_42166,N_37188,N_38569);
nor U42167 (N_42167,N_37549,N_35059);
nand U42168 (N_42168,N_38464,N_35698);
or U42169 (N_42169,N_36475,N_35563);
nand U42170 (N_42170,N_37365,N_37552);
or U42171 (N_42171,N_39955,N_37362);
and U42172 (N_42172,N_38319,N_38682);
nor U42173 (N_42173,N_37732,N_38315);
or U42174 (N_42174,N_38334,N_38533);
nor U42175 (N_42175,N_39369,N_35322);
xor U42176 (N_42176,N_37750,N_36768);
nand U42177 (N_42177,N_36411,N_35175);
xor U42178 (N_42178,N_35295,N_37647);
and U42179 (N_42179,N_38628,N_36794);
nor U42180 (N_42180,N_35626,N_37468);
nor U42181 (N_42181,N_39763,N_37856);
nand U42182 (N_42182,N_35944,N_35867);
and U42183 (N_42183,N_37201,N_39122);
or U42184 (N_42184,N_38587,N_36069);
and U42185 (N_42185,N_38970,N_36057);
xor U42186 (N_42186,N_38989,N_35092);
nand U42187 (N_42187,N_37166,N_36436);
or U42188 (N_42188,N_37547,N_35427);
or U42189 (N_42189,N_35743,N_37667);
and U42190 (N_42190,N_37048,N_39638);
xnor U42191 (N_42191,N_36167,N_38894);
and U42192 (N_42192,N_36723,N_37388);
and U42193 (N_42193,N_36932,N_36006);
xor U42194 (N_42194,N_36533,N_39681);
nand U42195 (N_42195,N_35444,N_38914);
or U42196 (N_42196,N_37072,N_35903);
nor U42197 (N_42197,N_38994,N_35537);
nand U42198 (N_42198,N_37984,N_35394);
or U42199 (N_42199,N_38756,N_36897);
nor U42200 (N_42200,N_37193,N_38341);
nand U42201 (N_42201,N_36770,N_36740);
nor U42202 (N_42202,N_35344,N_36949);
xor U42203 (N_42203,N_36658,N_35679);
or U42204 (N_42204,N_39701,N_37694);
xor U42205 (N_42205,N_36730,N_35190);
and U42206 (N_42206,N_38211,N_38830);
nand U42207 (N_42207,N_38819,N_36288);
xnor U42208 (N_42208,N_36616,N_36125);
or U42209 (N_42209,N_38972,N_39563);
or U42210 (N_42210,N_38308,N_37140);
nand U42211 (N_42211,N_39435,N_39333);
or U42212 (N_42212,N_37733,N_35389);
xnor U42213 (N_42213,N_36867,N_37027);
nor U42214 (N_42214,N_37031,N_39065);
nand U42215 (N_42215,N_39552,N_39204);
xnor U42216 (N_42216,N_39308,N_37708);
and U42217 (N_42217,N_35673,N_38288);
xnor U42218 (N_42218,N_39181,N_36339);
or U42219 (N_42219,N_38401,N_39787);
and U42220 (N_42220,N_39439,N_37224);
xor U42221 (N_42221,N_37337,N_38305);
and U42222 (N_42222,N_37719,N_38528);
or U42223 (N_42223,N_36271,N_36105);
nand U42224 (N_42224,N_38919,N_39430);
and U42225 (N_42225,N_35428,N_38087);
and U42226 (N_42226,N_39811,N_38414);
nor U42227 (N_42227,N_39510,N_37534);
nor U42228 (N_42228,N_36761,N_35064);
or U42229 (N_42229,N_39980,N_37073);
and U42230 (N_42230,N_37909,N_39036);
nor U42231 (N_42231,N_36739,N_39290);
nand U42232 (N_42232,N_35023,N_39902);
and U42233 (N_42233,N_39013,N_36394);
or U42234 (N_42234,N_38402,N_38646);
nand U42235 (N_42235,N_38337,N_38697);
and U42236 (N_42236,N_37904,N_38837);
nor U42237 (N_42237,N_38183,N_38400);
or U42238 (N_42238,N_39247,N_39729);
nand U42239 (N_42239,N_35830,N_37948);
nand U42240 (N_42240,N_39560,N_39331);
nand U42241 (N_42241,N_35260,N_39023);
and U42242 (N_42242,N_39721,N_39907);
nand U42243 (N_42243,N_39814,N_36166);
or U42244 (N_42244,N_36777,N_37320);
or U42245 (N_42245,N_35792,N_39011);
nand U42246 (N_42246,N_38583,N_39113);
nor U42247 (N_42247,N_38562,N_35751);
nor U42248 (N_42248,N_39651,N_37315);
or U42249 (N_42249,N_35235,N_39915);
xnor U42250 (N_42250,N_38530,N_38329);
nand U42251 (N_42251,N_38961,N_39664);
or U42252 (N_42252,N_37553,N_37531);
nand U42253 (N_42253,N_37945,N_35634);
xor U42254 (N_42254,N_36808,N_37967);
or U42255 (N_42255,N_38712,N_36293);
or U42256 (N_42256,N_35981,N_36032);
nor U42257 (N_42257,N_37369,N_38302);
or U42258 (N_42258,N_36921,N_39117);
and U42259 (N_42259,N_37782,N_35978);
xor U42260 (N_42260,N_35762,N_36098);
nand U42261 (N_42261,N_37372,N_35409);
nor U42262 (N_42262,N_38672,N_37920);
nor U42263 (N_42263,N_37761,N_39919);
nor U42264 (N_42264,N_38102,N_38633);
xnor U42265 (N_42265,N_35367,N_38575);
nor U42266 (N_42266,N_38347,N_39841);
and U42267 (N_42267,N_38155,N_36938);
xnor U42268 (N_42268,N_37206,N_35250);
xnor U42269 (N_42269,N_38580,N_37426);
nor U42270 (N_42270,N_35891,N_35570);
and U42271 (N_42271,N_38132,N_35352);
xnor U42272 (N_42272,N_37571,N_38413);
nand U42273 (N_42273,N_36786,N_35685);
nor U42274 (N_42274,N_39466,N_37679);
nor U42275 (N_42275,N_36231,N_38632);
nand U42276 (N_42276,N_38921,N_35985);
xnor U42277 (N_42277,N_36363,N_39903);
xor U42278 (N_42278,N_39311,N_36675);
nand U42279 (N_42279,N_36661,N_36272);
xor U42280 (N_42280,N_38823,N_38070);
nor U42281 (N_42281,N_39414,N_35819);
nand U42282 (N_42282,N_38081,N_37544);
and U42283 (N_42283,N_37514,N_39148);
or U42284 (N_42284,N_39833,N_38458);
and U42285 (N_42285,N_38978,N_37485);
and U42286 (N_42286,N_39054,N_35013);
nor U42287 (N_42287,N_39553,N_38264);
and U42288 (N_42288,N_37636,N_37756);
xnor U42289 (N_42289,N_35574,N_37002);
nor U42290 (N_42290,N_35720,N_36850);
and U42291 (N_42291,N_36586,N_37183);
or U42292 (N_42292,N_39477,N_37119);
or U42293 (N_42293,N_36834,N_35917);
nand U42294 (N_42294,N_35431,N_38683);
and U42295 (N_42295,N_35540,N_37567);
and U42296 (N_42296,N_38713,N_36338);
xor U42297 (N_42297,N_37946,N_39828);
or U42298 (N_42298,N_38965,N_39745);
and U42299 (N_42299,N_37174,N_36991);
or U42300 (N_42300,N_36956,N_36041);
nand U42301 (N_42301,N_37110,N_39363);
nand U42302 (N_42302,N_38985,N_38993);
nand U42303 (N_42303,N_37411,N_36572);
or U42304 (N_42304,N_36716,N_37851);
and U42305 (N_42305,N_38550,N_36303);
and U42306 (N_42306,N_36531,N_35905);
and U42307 (N_42307,N_39119,N_38377);
nor U42308 (N_42308,N_37830,N_39582);
or U42309 (N_42309,N_35101,N_35592);
xnor U42310 (N_42310,N_36079,N_36200);
or U42311 (N_42311,N_39273,N_35309);
nor U42312 (N_42312,N_39157,N_35278);
or U42313 (N_42313,N_37008,N_37996);
xnor U42314 (N_42314,N_35067,N_38943);
xor U42315 (N_42315,N_37286,N_37958);
or U42316 (N_42316,N_36515,N_36205);
and U42317 (N_42317,N_35372,N_36045);
xnor U42318 (N_42318,N_38299,N_35749);
xnor U42319 (N_42319,N_37607,N_38727);
nor U42320 (N_42320,N_36606,N_37885);
nor U42321 (N_42321,N_35969,N_36234);
or U42322 (N_42322,N_36323,N_37142);
and U42323 (N_42323,N_37688,N_35005);
and U42324 (N_42324,N_39091,N_37964);
nor U42325 (N_42325,N_37883,N_39445);
and U42326 (N_42326,N_37432,N_35489);
and U42327 (N_42327,N_38100,N_35110);
and U42328 (N_42328,N_35677,N_37602);
nand U42329 (N_42329,N_35536,N_35569);
or U42330 (N_42330,N_38815,N_35104);
and U42331 (N_42331,N_37165,N_39243);
and U42332 (N_42332,N_39034,N_38077);
or U42333 (N_42333,N_36542,N_39499);
xnor U42334 (N_42334,N_39218,N_39599);
xor U42335 (N_42335,N_37368,N_35520);
or U42336 (N_42336,N_37066,N_35911);
nand U42337 (N_42337,N_36874,N_37387);
nor U42338 (N_42338,N_39059,N_36555);
or U42339 (N_42339,N_37992,N_36720);
or U42340 (N_42340,N_36368,N_38513);
and U42341 (N_42341,N_39924,N_35608);
or U42342 (N_42342,N_38588,N_38049);
nand U42343 (N_42343,N_35630,N_39206);
or U42344 (N_42344,N_37246,N_35095);
nor U42345 (N_42345,N_38311,N_37446);
and U42346 (N_42346,N_36335,N_38826);
xnor U42347 (N_42347,N_36347,N_37968);
nor U42348 (N_42348,N_39164,N_36511);
xor U42349 (N_42349,N_38307,N_37823);
or U42350 (N_42350,N_38796,N_38726);
or U42351 (N_42351,N_39704,N_38069);
or U42352 (N_42352,N_39398,N_36258);
and U42353 (N_42353,N_38937,N_37618);
xor U42354 (N_42354,N_36097,N_36441);
xor U42355 (N_42355,N_37097,N_38446);
nand U42356 (N_42356,N_35512,N_38303);
nand U42357 (N_42357,N_38952,N_39501);
xor U42358 (N_42358,N_38862,N_35784);
or U42359 (N_42359,N_36061,N_36206);
nor U42360 (N_42360,N_38066,N_38260);
and U42361 (N_42361,N_37158,N_37175);
or U42362 (N_42362,N_39285,N_39557);
nor U42363 (N_42363,N_36855,N_35144);
nand U42364 (N_42364,N_38865,N_36294);
xnor U42365 (N_42365,N_39709,N_35811);
and U42366 (N_42366,N_35142,N_36275);
nand U42367 (N_42367,N_37313,N_39033);
nor U42368 (N_42368,N_36536,N_38222);
nor U42369 (N_42369,N_39419,N_36742);
nor U42370 (N_42370,N_35091,N_39212);
or U42371 (N_42371,N_36425,N_37129);
nor U42372 (N_42372,N_39490,N_39692);
or U42373 (N_42373,N_36918,N_36562);
nor U42374 (N_42374,N_37424,N_35687);
and U42375 (N_42375,N_35511,N_36487);
or U42376 (N_42376,N_39720,N_35108);
and U42377 (N_42377,N_39145,N_38594);
and U42378 (N_42378,N_35231,N_39322);
nand U42379 (N_42379,N_38210,N_38068);
and U42380 (N_42380,N_38406,N_36068);
nand U42381 (N_42381,N_35286,N_38988);
or U42382 (N_42382,N_36624,N_37766);
nand U42383 (N_42383,N_36131,N_36075);
and U42384 (N_42384,N_37546,N_38514);
or U42385 (N_42385,N_36577,N_35006);
or U42386 (N_42386,N_39784,N_39851);
and U42387 (N_42387,N_39700,N_38015);
nor U42388 (N_42388,N_36988,N_37986);
or U42389 (N_42389,N_39871,N_36685);
xnor U42390 (N_42390,N_38331,N_39101);
xor U42391 (N_42391,N_38878,N_38835);
or U42392 (N_42392,N_36282,N_37179);
and U42393 (N_42393,N_39194,N_36152);
or U42394 (N_42394,N_38179,N_38828);
or U42395 (N_42395,N_38935,N_36254);
and U42396 (N_42396,N_35143,N_35600);
and U42397 (N_42397,N_37358,N_39618);
xor U42398 (N_42398,N_37654,N_38929);
nor U42399 (N_42399,N_38104,N_39349);
xor U42400 (N_42400,N_37311,N_38321);
xnor U42401 (N_42401,N_36869,N_39595);
nor U42402 (N_42402,N_37814,N_35111);
and U42403 (N_42403,N_36743,N_38895);
nand U42404 (N_42404,N_38610,N_35351);
or U42405 (N_42405,N_39436,N_37914);
or U42406 (N_42406,N_35105,N_39645);
xnor U42407 (N_42407,N_36306,N_36711);
nand U42408 (N_42408,N_39370,N_36262);
nand U42409 (N_42409,N_37376,N_37850);
xor U42410 (N_42410,N_39021,N_35798);
nor U42411 (N_42411,N_38854,N_38008);
xor U42412 (N_42412,N_37663,N_37476);
xnor U42413 (N_42413,N_37327,N_39854);
xor U42414 (N_42414,N_38359,N_38221);
nor U42415 (N_42415,N_38553,N_36426);
nand U42416 (N_42416,N_39521,N_39063);
or U42417 (N_42417,N_37244,N_37953);
nand U42418 (N_42418,N_37003,N_35825);
and U42419 (N_42419,N_39603,N_36948);
nor U42420 (N_42420,N_38089,N_36387);
nor U42421 (N_42421,N_37912,N_37273);
xnor U42422 (N_42422,N_35880,N_35176);
nor U42423 (N_42423,N_35976,N_38128);
or U42424 (N_42424,N_37513,N_39561);
nand U42425 (N_42425,N_38899,N_36691);
xor U42426 (N_42426,N_38187,N_36277);
nand U42427 (N_42427,N_36840,N_36207);
xnor U42428 (N_42428,N_36447,N_38625);
or U42429 (N_42429,N_36856,N_37743);
or U42430 (N_42430,N_36501,N_35739);
xnor U42431 (N_42431,N_38647,N_37977);
nor U42432 (N_42432,N_38375,N_38274);
xor U42433 (N_42433,N_38384,N_38114);
or U42434 (N_42434,N_39210,N_36186);
or U42435 (N_42435,N_38316,N_39665);
or U42436 (N_42436,N_39989,N_39921);
nand U42437 (N_42437,N_37807,N_39474);
or U42438 (N_42438,N_35623,N_36828);
nand U42439 (N_42439,N_36654,N_36601);
xnor U42440 (N_42440,N_37453,N_37321);
xnor U42441 (N_42441,N_39747,N_38226);
xor U42442 (N_42442,N_38853,N_36575);
and U42443 (N_42443,N_39411,N_39301);
xor U42444 (N_42444,N_35338,N_37490);
and U42445 (N_42445,N_35645,N_36971);
or U42446 (N_42446,N_36847,N_36753);
nor U42447 (N_42447,N_37403,N_35335);
nor U42448 (N_42448,N_37816,N_39321);
and U42449 (N_42449,N_35936,N_38744);
and U42450 (N_42450,N_35033,N_39155);
nand U42451 (N_42451,N_38356,N_36530);
nand U42452 (N_42452,N_36526,N_36185);
nor U42453 (N_42453,N_35865,N_39967);
nor U42454 (N_42454,N_37736,N_37488);
or U42455 (N_42455,N_37902,N_39002);
nand U42456 (N_42456,N_39978,N_39459);
and U42457 (N_42457,N_36406,N_36811);
xnor U42458 (N_42458,N_37834,N_36951);
xnor U42459 (N_42459,N_35663,N_39711);
xnor U42460 (N_42460,N_37956,N_36495);
nor U42461 (N_42461,N_35358,N_35467);
nor U42462 (N_42462,N_38404,N_38168);
or U42463 (N_42463,N_37456,N_36255);
xor U42464 (N_42464,N_39946,N_37266);
and U42465 (N_42465,N_37754,N_38373);
or U42466 (N_42466,N_39310,N_38794);
xnor U42467 (N_42467,N_39575,N_37117);
nor U42468 (N_42468,N_37493,N_38915);
or U42469 (N_42469,N_35137,N_37537);
and U42470 (N_42470,N_35207,N_39514);
or U42471 (N_42471,N_38684,N_37780);
nand U42472 (N_42472,N_37847,N_35247);
nor U42473 (N_42473,N_36274,N_35834);
nand U42474 (N_42474,N_35036,N_35375);
or U42475 (N_42475,N_39825,N_38770);
nor U42476 (N_42476,N_38140,N_38392);
or U42477 (N_42477,N_37653,N_39400);
or U42478 (N_42478,N_36142,N_35814);
and U42479 (N_42479,N_37330,N_38212);
or U42480 (N_42480,N_37479,N_35726);
and U42481 (N_42481,N_38924,N_38206);
xnor U42482 (N_42482,N_38776,N_35380);
nor U42483 (N_42483,N_35618,N_39100);
and U42484 (N_42484,N_36217,N_36604);
nor U42485 (N_42485,N_36162,N_35211);
xnor U42486 (N_42486,N_36747,N_36153);
nor U42487 (N_42487,N_37801,N_39656);
nand U42488 (N_42488,N_37180,N_37038);
or U42489 (N_42489,N_39086,N_39271);
or U42490 (N_42490,N_39375,N_37522);
or U42491 (N_42491,N_36298,N_38984);
or U42492 (N_42492,N_37857,N_37112);
nand U42493 (N_42493,N_38033,N_38829);
or U42494 (N_42494,N_39892,N_37435);
or U42495 (N_42495,N_37930,N_38026);
or U42496 (N_42496,N_36439,N_37915);
nand U42497 (N_42497,N_37677,N_37333);
nor U42498 (N_42498,N_36286,N_39316);
nand U42499 (N_42499,N_38322,N_38558);
or U42500 (N_42500,N_37421,N_35752);
xnor U42501 (N_42501,N_36730,N_37967);
nor U42502 (N_42502,N_37806,N_39798);
nor U42503 (N_42503,N_37710,N_37330);
xnor U42504 (N_42504,N_36509,N_37289);
nand U42505 (N_42505,N_39770,N_38572);
and U42506 (N_42506,N_36344,N_36771);
nor U42507 (N_42507,N_38043,N_39447);
xor U42508 (N_42508,N_39106,N_37624);
or U42509 (N_42509,N_39699,N_38470);
xnor U42510 (N_42510,N_38482,N_39737);
nor U42511 (N_42511,N_36983,N_39577);
or U42512 (N_42512,N_39621,N_39142);
nor U42513 (N_42513,N_35398,N_38554);
nand U42514 (N_42514,N_38506,N_36767);
nor U42515 (N_42515,N_39929,N_35154);
or U42516 (N_42516,N_35456,N_39027);
and U42517 (N_42517,N_39825,N_37106);
xnor U42518 (N_42518,N_35335,N_37084);
or U42519 (N_42519,N_36604,N_36961);
or U42520 (N_42520,N_37865,N_37324);
or U42521 (N_42521,N_35913,N_37481);
and U42522 (N_42522,N_36502,N_38121);
xor U42523 (N_42523,N_36246,N_39743);
nand U42524 (N_42524,N_36251,N_38114);
or U42525 (N_42525,N_38731,N_36191);
and U42526 (N_42526,N_35894,N_36139);
or U42527 (N_42527,N_37342,N_39795);
nand U42528 (N_42528,N_36057,N_37785);
nand U42529 (N_42529,N_39783,N_38095);
xor U42530 (N_42530,N_38228,N_36379);
xor U42531 (N_42531,N_35915,N_38039);
and U42532 (N_42532,N_38278,N_36017);
or U42533 (N_42533,N_37409,N_35267);
xnor U42534 (N_42534,N_37215,N_35248);
nor U42535 (N_42535,N_35710,N_37794);
xor U42536 (N_42536,N_35876,N_39419);
or U42537 (N_42537,N_39755,N_39741);
nor U42538 (N_42538,N_36872,N_37541);
or U42539 (N_42539,N_39616,N_38567);
xor U42540 (N_42540,N_36042,N_39359);
xnor U42541 (N_42541,N_35696,N_36580);
and U42542 (N_42542,N_38700,N_35639);
and U42543 (N_42543,N_37082,N_39138);
nor U42544 (N_42544,N_36880,N_37410);
and U42545 (N_42545,N_37353,N_38654);
nand U42546 (N_42546,N_39479,N_36657);
or U42547 (N_42547,N_35887,N_36374);
nor U42548 (N_42548,N_38534,N_35058);
and U42549 (N_42549,N_37400,N_35513);
and U42550 (N_42550,N_35967,N_39130);
xnor U42551 (N_42551,N_39514,N_35634);
and U42552 (N_42552,N_37165,N_37777);
and U42553 (N_42553,N_36211,N_37298);
or U42554 (N_42554,N_35656,N_36882);
or U42555 (N_42555,N_37621,N_35129);
and U42556 (N_42556,N_37623,N_39801);
xor U42557 (N_42557,N_38678,N_38884);
nor U42558 (N_42558,N_35688,N_39435);
or U42559 (N_42559,N_35325,N_35905);
nor U42560 (N_42560,N_38308,N_37326);
or U42561 (N_42561,N_36443,N_37375);
nand U42562 (N_42562,N_39296,N_37763);
and U42563 (N_42563,N_35628,N_35639);
xnor U42564 (N_42564,N_35282,N_36917);
nor U42565 (N_42565,N_37872,N_39561);
or U42566 (N_42566,N_38158,N_37640);
xor U42567 (N_42567,N_36612,N_35614);
xnor U42568 (N_42568,N_37125,N_36816);
nor U42569 (N_42569,N_38766,N_36670);
nand U42570 (N_42570,N_38906,N_39022);
and U42571 (N_42571,N_37271,N_36735);
nand U42572 (N_42572,N_36868,N_37260);
nor U42573 (N_42573,N_39440,N_36134);
and U42574 (N_42574,N_35996,N_39232);
xor U42575 (N_42575,N_38050,N_37111);
xor U42576 (N_42576,N_38618,N_39341);
xnor U42577 (N_42577,N_38234,N_38736);
nand U42578 (N_42578,N_39478,N_37247);
or U42579 (N_42579,N_39001,N_35925);
nor U42580 (N_42580,N_38556,N_38699);
or U42581 (N_42581,N_35411,N_39735);
and U42582 (N_42582,N_38616,N_37856);
xor U42583 (N_42583,N_37654,N_36803);
or U42584 (N_42584,N_37604,N_35205);
or U42585 (N_42585,N_37515,N_37400);
nand U42586 (N_42586,N_36407,N_35858);
or U42587 (N_42587,N_35276,N_35584);
nand U42588 (N_42588,N_35382,N_36500);
xor U42589 (N_42589,N_36291,N_38173);
xnor U42590 (N_42590,N_35681,N_35727);
nand U42591 (N_42591,N_38294,N_38153);
nor U42592 (N_42592,N_39837,N_39523);
or U42593 (N_42593,N_35975,N_39210);
nor U42594 (N_42594,N_39801,N_35883);
nand U42595 (N_42595,N_38027,N_36677);
nor U42596 (N_42596,N_37891,N_35340);
nand U42597 (N_42597,N_36452,N_37532);
xor U42598 (N_42598,N_39224,N_35086);
xor U42599 (N_42599,N_35913,N_35867);
nand U42600 (N_42600,N_36167,N_36773);
and U42601 (N_42601,N_38624,N_39534);
or U42602 (N_42602,N_36006,N_39189);
or U42603 (N_42603,N_35967,N_38971);
and U42604 (N_42604,N_39829,N_38941);
or U42605 (N_42605,N_39927,N_36163);
nand U42606 (N_42606,N_36960,N_38992);
nand U42607 (N_42607,N_39950,N_37969);
nor U42608 (N_42608,N_35795,N_39354);
nor U42609 (N_42609,N_37548,N_38812);
or U42610 (N_42610,N_37316,N_39494);
nand U42611 (N_42611,N_36605,N_35402);
nor U42612 (N_42612,N_39463,N_37736);
or U42613 (N_42613,N_35425,N_38848);
or U42614 (N_42614,N_35996,N_35622);
xor U42615 (N_42615,N_39373,N_37050);
xor U42616 (N_42616,N_39696,N_38216);
xnor U42617 (N_42617,N_35807,N_37008);
xor U42618 (N_42618,N_38017,N_36082);
or U42619 (N_42619,N_37098,N_35595);
nand U42620 (N_42620,N_39020,N_37118);
xnor U42621 (N_42621,N_37434,N_37220);
or U42622 (N_42622,N_39716,N_37679);
nand U42623 (N_42623,N_37606,N_39918);
nand U42624 (N_42624,N_35186,N_38074);
xor U42625 (N_42625,N_37097,N_38605);
xnor U42626 (N_42626,N_37820,N_36664);
and U42627 (N_42627,N_37502,N_39881);
nor U42628 (N_42628,N_39145,N_39686);
nand U42629 (N_42629,N_36385,N_38248);
and U42630 (N_42630,N_38033,N_35544);
nand U42631 (N_42631,N_36082,N_37255);
or U42632 (N_42632,N_36700,N_37681);
nor U42633 (N_42633,N_38152,N_36279);
xor U42634 (N_42634,N_39360,N_38851);
nand U42635 (N_42635,N_35980,N_39429);
nor U42636 (N_42636,N_37237,N_37707);
nand U42637 (N_42637,N_37357,N_35540);
nor U42638 (N_42638,N_35870,N_36096);
xnor U42639 (N_42639,N_35237,N_38957);
and U42640 (N_42640,N_37960,N_36774);
and U42641 (N_42641,N_35215,N_39910);
nor U42642 (N_42642,N_35654,N_35821);
and U42643 (N_42643,N_39197,N_37514);
and U42644 (N_42644,N_39283,N_37478);
xnor U42645 (N_42645,N_35013,N_39369);
and U42646 (N_42646,N_38331,N_35139);
nor U42647 (N_42647,N_36094,N_38991);
or U42648 (N_42648,N_35941,N_37499);
nand U42649 (N_42649,N_37059,N_37753);
and U42650 (N_42650,N_39938,N_39888);
and U42651 (N_42651,N_39797,N_37364);
xor U42652 (N_42652,N_37841,N_38276);
and U42653 (N_42653,N_39541,N_35429);
and U42654 (N_42654,N_37147,N_37994);
nand U42655 (N_42655,N_39663,N_37668);
nand U42656 (N_42656,N_35053,N_39909);
nor U42657 (N_42657,N_36087,N_38653);
or U42658 (N_42658,N_36234,N_36938);
xor U42659 (N_42659,N_39969,N_39530);
nor U42660 (N_42660,N_38973,N_38492);
nand U42661 (N_42661,N_38601,N_38532);
nand U42662 (N_42662,N_38226,N_36958);
xnor U42663 (N_42663,N_38662,N_38816);
or U42664 (N_42664,N_36437,N_36858);
nand U42665 (N_42665,N_36858,N_39241);
nand U42666 (N_42666,N_36425,N_38587);
xnor U42667 (N_42667,N_37914,N_38371);
or U42668 (N_42668,N_39097,N_35833);
xor U42669 (N_42669,N_36523,N_38682);
and U42670 (N_42670,N_37550,N_36463);
nor U42671 (N_42671,N_38921,N_37078);
xor U42672 (N_42672,N_37576,N_36417);
and U42673 (N_42673,N_36286,N_37798);
and U42674 (N_42674,N_37801,N_39323);
nand U42675 (N_42675,N_37284,N_38498);
and U42676 (N_42676,N_35934,N_37220);
nand U42677 (N_42677,N_37984,N_36551);
and U42678 (N_42678,N_37215,N_38196);
and U42679 (N_42679,N_38941,N_37279);
and U42680 (N_42680,N_39524,N_37819);
or U42681 (N_42681,N_37427,N_37388);
nand U42682 (N_42682,N_38645,N_35642);
xor U42683 (N_42683,N_37995,N_38584);
nand U42684 (N_42684,N_36726,N_39967);
and U42685 (N_42685,N_35587,N_37964);
xnor U42686 (N_42686,N_36578,N_35940);
nand U42687 (N_42687,N_36717,N_35837);
xor U42688 (N_42688,N_38109,N_39687);
nand U42689 (N_42689,N_38651,N_36073);
xor U42690 (N_42690,N_37482,N_36582);
xnor U42691 (N_42691,N_37814,N_36016);
or U42692 (N_42692,N_39622,N_36155);
or U42693 (N_42693,N_35635,N_35262);
nor U42694 (N_42694,N_38627,N_36481);
nor U42695 (N_42695,N_38619,N_38909);
nor U42696 (N_42696,N_39782,N_36894);
and U42697 (N_42697,N_37752,N_35496);
nor U42698 (N_42698,N_38295,N_38536);
xnor U42699 (N_42699,N_39452,N_39460);
or U42700 (N_42700,N_36624,N_35445);
and U42701 (N_42701,N_37145,N_39566);
nor U42702 (N_42702,N_37246,N_35946);
xnor U42703 (N_42703,N_39332,N_37654);
and U42704 (N_42704,N_38282,N_36021);
nor U42705 (N_42705,N_39068,N_37740);
or U42706 (N_42706,N_36626,N_35492);
xnor U42707 (N_42707,N_35822,N_39307);
or U42708 (N_42708,N_37877,N_35191);
and U42709 (N_42709,N_38667,N_35625);
or U42710 (N_42710,N_38650,N_38143);
nand U42711 (N_42711,N_35134,N_35064);
nand U42712 (N_42712,N_39150,N_35836);
and U42713 (N_42713,N_39402,N_35940);
nand U42714 (N_42714,N_38345,N_39485);
or U42715 (N_42715,N_38223,N_38872);
nand U42716 (N_42716,N_36838,N_38327);
nor U42717 (N_42717,N_38110,N_37336);
nand U42718 (N_42718,N_36694,N_39185);
nor U42719 (N_42719,N_36090,N_37999);
nor U42720 (N_42720,N_38526,N_35299);
nor U42721 (N_42721,N_37455,N_36433);
or U42722 (N_42722,N_38122,N_35310);
and U42723 (N_42723,N_39230,N_36040);
nor U42724 (N_42724,N_38395,N_37985);
and U42725 (N_42725,N_37198,N_37529);
nor U42726 (N_42726,N_37251,N_35140);
nor U42727 (N_42727,N_36597,N_35485);
and U42728 (N_42728,N_39481,N_37545);
and U42729 (N_42729,N_38449,N_37344);
nand U42730 (N_42730,N_36861,N_38073);
or U42731 (N_42731,N_37987,N_38451);
or U42732 (N_42732,N_36751,N_36235);
nor U42733 (N_42733,N_39346,N_37898);
nand U42734 (N_42734,N_39663,N_37433);
and U42735 (N_42735,N_37229,N_37969);
nand U42736 (N_42736,N_35850,N_37104);
xnor U42737 (N_42737,N_37592,N_36244);
xor U42738 (N_42738,N_38402,N_35640);
nor U42739 (N_42739,N_35798,N_35474);
nor U42740 (N_42740,N_37665,N_37858);
or U42741 (N_42741,N_36368,N_39478);
nor U42742 (N_42742,N_37584,N_38849);
xnor U42743 (N_42743,N_39862,N_37185);
and U42744 (N_42744,N_39153,N_39491);
or U42745 (N_42745,N_35384,N_36281);
and U42746 (N_42746,N_38726,N_39466);
and U42747 (N_42747,N_37132,N_36809);
nor U42748 (N_42748,N_38584,N_36405);
nand U42749 (N_42749,N_35287,N_37467);
nor U42750 (N_42750,N_39219,N_35242);
xnor U42751 (N_42751,N_38827,N_35522);
xor U42752 (N_42752,N_35007,N_35348);
and U42753 (N_42753,N_35977,N_38933);
xor U42754 (N_42754,N_35881,N_35109);
or U42755 (N_42755,N_37760,N_39207);
nand U42756 (N_42756,N_39584,N_38769);
xnor U42757 (N_42757,N_35286,N_35319);
nand U42758 (N_42758,N_36785,N_38297);
xnor U42759 (N_42759,N_35541,N_37138);
xor U42760 (N_42760,N_39329,N_36032);
nor U42761 (N_42761,N_36576,N_37545);
and U42762 (N_42762,N_37337,N_39899);
nand U42763 (N_42763,N_36903,N_35929);
nand U42764 (N_42764,N_38879,N_36266);
xnor U42765 (N_42765,N_37373,N_38832);
nand U42766 (N_42766,N_37318,N_36119);
nand U42767 (N_42767,N_36802,N_36403);
or U42768 (N_42768,N_35984,N_36692);
and U42769 (N_42769,N_36143,N_38236);
or U42770 (N_42770,N_38868,N_35995);
nand U42771 (N_42771,N_37778,N_38512);
nor U42772 (N_42772,N_39849,N_38913);
xor U42773 (N_42773,N_36853,N_36048);
and U42774 (N_42774,N_35384,N_36254);
xnor U42775 (N_42775,N_35028,N_37812);
nand U42776 (N_42776,N_35918,N_35691);
nor U42777 (N_42777,N_39428,N_39188);
and U42778 (N_42778,N_39833,N_39450);
or U42779 (N_42779,N_37931,N_36349);
nor U42780 (N_42780,N_35773,N_36983);
nor U42781 (N_42781,N_38035,N_36100);
nand U42782 (N_42782,N_36356,N_35634);
nand U42783 (N_42783,N_35930,N_38674);
nand U42784 (N_42784,N_36274,N_37329);
nor U42785 (N_42785,N_37094,N_36771);
and U42786 (N_42786,N_39813,N_37550);
nor U42787 (N_42787,N_35380,N_37293);
nor U42788 (N_42788,N_38781,N_37830);
nor U42789 (N_42789,N_37926,N_38112);
xor U42790 (N_42790,N_38307,N_37191);
xnor U42791 (N_42791,N_39931,N_36779);
nand U42792 (N_42792,N_37409,N_37792);
nand U42793 (N_42793,N_38601,N_35832);
and U42794 (N_42794,N_37032,N_37985);
xor U42795 (N_42795,N_39267,N_38824);
or U42796 (N_42796,N_35320,N_38151);
or U42797 (N_42797,N_38006,N_38534);
and U42798 (N_42798,N_36600,N_37709);
and U42799 (N_42799,N_36712,N_39637);
and U42800 (N_42800,N_36285,N_37226);
and U42801 (N_42801,N_39814,N_35511);
nor U42802 (N_42802,N_35916,N_37854);
xor U42803 (N_42803,N_36947,N_36609);
nor U42804 (N_42804,N_38153,N_39572);
or U42805 (N_42805,N_37162,N_37880);
or U42806 (N_42806,N_36710,N_39212);
xor U42807 (N_42807,N_35682,N_39562);
or U42808 (N_42808,N_37678,N_38231);
or U42809 (N_42809,N_35445,N_36499);
nand U42810 (N_42810,N_37942,N_37672);
nand U42811 (N_42811,N_37047,N_36114);
nand U42812 (N_42812,N_35660,N_36485);
xnor U42813 (N_42813,N_37552,N_37525);
nor U42814 (N_42814,N_37395,N_38670);
or U42815 (N_42815,N_39460,N_35539);
nor U42816 (N_42816,N_39559,N_37197);
xnor U42817 (N_42817,N_39255,N_38919);
or U42818 (N_42818,N_37394,N_39720);
nand U42819 (N_42819,N_35885,N_38036);
xor U42820 (N_42820,N_37186,N_39171);
xor U42821 (N_42821,N_38348,N_35324);
nand U42822 (N_42822,N_38485,N_37322);
or U42823 (N_42823,N_36547,N_37402);
nor U42824 (N_42824,N_36096,N_35519);
nand U42825 (N_42825,N_38062,N_37074);
nor U42826 (N_42826,N_36025,N_39166);
nor U42827 (N_42827,N_36253,N_37059);
nor U42828 (N_42828,N_37551,N_35310);
and U42829 (N_42829,N_39506,N_36266);
or U42830 (N_42830,N_36871,N_35074);
nor U42831 (N_42831,N_38260,N_38099);
or U42832 (N_42832,N_35886,N_36995);
xnor U42833 (N_42833,N_39941,N_38783);
nand U42834 (N_42834,N_35843,N_39478);
xor U42835 (N_42835,N_37905,N_39407);
nor U42836 (N_42836,N_38417,N_38187);
nor U42837 (N_42837,N_38778,N_37321);
nor U42838 (N_42838,N_38522,N_37077);
or U42839 (N_42839,N_38374,N_39083);
or U42840 (N_42840,N_37018,N_37488);
nor U42841 (N_42841,N_38855,N_35716);
and U42842 (N_42842,N_37177,N_37938);
or U42843 (N_42843,N_36910,N_36445);
and U42844 (N_42844,N_39629,N_35276);
or U42845 (N_42845,N_35525,N_39371);
nor U42846 (N_42846,N_35709,N_36412);
and U42847 (N_42847,N_39461,N_39320);
or U42848 (N_42848,N_39122,N_37548);
xnor U42849 (N_42849,N_39367,N_37046);
nand U42850 (N_42850,N_38198,N_35457);
and U42851 (N_42851,N_37749,N_38784);
nand U42852 (N_42852,N_36856,N_38323);
xnor U42853 (N_42853,N_38163,N_39401);
nand U42854 (N_42854,N_38491,N_36595);
xor U42855 (N_42855,N_36382,N_37174);
nand U42856 (N_42856,N_36193,N_38097);
or U42857 (N_42857,N_36934,N_37360);
nor U42858 (N_42858,N_36772,N_35769);
and U42859 (N_42859,N_36581,N_37755);
xor U42860 (N_42860,N_35393,N_35855);
or U42861 (N_42861,N_37683,N_39180);
and U42862 (N_42862,N_35949,N_35035);
and U42863 (N_42863,N_35719,N_39446);
xor U42864 (N_42864,N_37751,N_38892);
and U42865 (N_42865,N_39527,N_37248);
xnor U42866 (N_42866,N_38940,N_36415);
nand U42867 (N_42867,N_38010,N_36627);
nor U42868 (N_42868,N_38349,N_37100);
xor U42869 (N_42869,N_35410,N_38418);
xor U42870 (N_42870,N_39500,N_38480);
nand U42871 (N_42871,N_37275,N_37196);
xor U42872 (N_42872,N_39543,N_36255);
xor U42873 (N_42873,N_35581,N_38771);
or U42874 (N_42874,N_36519,N_36602);
and U42875 (N_42875,N_37372,N_35715);
nand U42876 (N_42876,N_39501,N_38554);
nand U42877 (N_42877,N_39718,N_39324);
or U42878 (N_42878,N_38723,N_37711);
nand U42879 (N_42879,N_37564,N_35994);
or U42880 (N_42880,N_37387,N_39065);
xor U42881 (N_42881,N_38661,N_38253);
xor U42882 (N_42882,N_35313,N_38794);
and U42883 (N_42883,N_39723,N_38074);
or U42884 (N_42884,N_35865,N_38620);
and U42885 (N_42885,N_37947,N_35415);
xnor U42886 (N_42886,N_35728,N_36130);
or U42887 (N_42887,N_36809,N_38210);
nor U42888 (N_42888,N_37026,N_37721);
nor U42889 (N_42889,N_36519,N_39943);
xor U42890 (N_42890,N_37737,N_36048);
or U42891 (N_42891,N_38803,N_35122);
xnor U42892 (N_42892,N_39969,N_37244);
and U42893 (N_42893,N_35669,N_36574);
nand U42894 (N_42894,N_36886,N_39697);
or U42895 (N_42895,N_38620,N_35950);
xor U42896 (N_42896,N_37906,N_38713);
or U42897 (N_42897,N_37413,N_37309);
xor U42898 (N_42898,N_39954,N_36947);
and U42899 (N_42899,N_38555,N_35138);
or U42900 (N_42900,N_36115,N_39782);
nor U42901 (N_42901,N_38378,N_39709);
nor U42902 (N_42902,N_36475,N_36899);
xor U42903 (N_42903,N_36268,N_38822);
or U42904 (N_42904,N_36308,N_36297);
nand U42905 (N_42905,N_37691,N_38447);
xor U42906 (N_42906,N_35944,N_39046);
and U42907 (N_42907,N_37182,N_38725);
nor U42908 (N_42908,N_35436,N_38107);
and U42909 (N_42909,N_38010,N_39572);
nand U42910 (N_42910,N_37035,N_38561);
xnor U42911 (N_42911,N_37256,N_36046);
nand U42912 (N_42912,N_38518,N_37288);
or U42913 (N_42913,N_36425,N_37842);
nor U42914 (N_42914,N_37493,N_36792);
nand U42915 (N_42915,N_38562,N_36872);
xnor U42916 (N_42916,N_36043,N_35669);
xor U42917 (N_42917,N_36241,N_39224);
and U42918 (N_42918,N_37832,N_35279);
xnor U42919 (N_42919,N_37077,N_35824);
xor U42920 (N_42920,N_35906,N_39998);
xnor U42921 (N_42921,N_38511,N_39232);
or U42922 (N_42922,N_37600,N_35974);
nor U42923 (N_42923,N_39108,N_37363);
nor U42924 (N_42924,N_35674,N_35330);
nor U42925 (N_42925,N_36785,N_36232);
or U42926 (N_42926,N_35230,N_39658);
xor U42927 (N_42927,N_37066,N_37512);
nand U42928 (N_42928,N_36367,N_36809);
xor U42929 (N_42929,N_37424,N_35364);
and U42930 (N_42930,N_39398,N_38768);
xnor U42931 (N_42931,N_36438,N_38897);
and U42932 (N_42932,N_37252,N_38879);
and U42933 (N_42933,N_36974,N_35039);
nand U42934 (N_42934,N_37250,N_38127);
xor U42935 (N_42935,N_39563,N_36398);
xnor U42936 (N_42936,N_38349,N_35820);
nor U42937 (N_42937,N_37233,N_38039);
xor U42938 (N_42938,N_36060,N_38178);
and U42939 (N_42939,N_37220,N_39614);
xnor U42940 (N_42940,N_37827,N_35371);
or U42941 (N_42941,N_37845,N_35340);
xnor U42942 (N_42942,N_39615,N_38312);
xor U42943 (N_42943,N_36904,N_39362);
nor U42944 (N_42944,N_37724,N_35115);
and U42945 (N_42945,N_38620,N_39019);
nor U42946 (N_42946,N_39132,N_37749);
nor U42947 (N_42947,N_37990,N_35499);
xnor U42948 (N_42948,N_37351,N_39265);
nand U42949 (N_42949,N_39731,N_35325);
nand U42950 (N_42950,N_37441,N_35023);
or U42951 (N_42951,N_39976,N_39140);
and U42952 (N_42952,N_39460,N_37395);
nor U42953 (N_42953,N_37197,N_38144);
xnor U42954 (N_42954,N_35681,N_38562);
nand U42955 (N_42955,N_35606,N_38622);
and U42956 (N_42956,N_35383,N_38300);
nor U42957 (N_42957,N_39917,N_37190);
xor U42958 (N_42958,N_36472,N_39979);
xor U42959 (N_42959,N_38880,N_36612);
and U42960 (N_42960,N_35888,N_37972);
nor U42961 (N_42961,N_38887,N_39473);
nor U42962 (N_42962,N_38371,N_37252);
or U42963 (N_42963,N_37864,N_36016);
and U42964 (N_42964,N_38008,N_39684);
nor U42965 (N_42965,N_36869,N_39193);
or U42966 (N_42966,N_37099,N_39180);
xor U42967 (N_42967,N_36954,N_38639);
and U42968 (N_42968,N_35469,N_38920);
or U42969 (N_42969,N_38549,N_35373);
nand U42970 (N_42970,N_39341,N_39796);
nor U42971 (N_42971,N_39128,N_35629);
nand U42972 (N_42972,N_37808,N_38440);
or U42973 (N_42973,N_39508,N_35950);
nor U42974 (N_42974,N_39948,N_37157);
or U42975 (N_42975,N_37225,N_35599);
nor U42976 (N_42976,N_35341,N_36504);
or U42977 (N_42977,N_39097,N_39806);
and U42978 (N_42978,N_35701,N_38681);
nor U42979 (N_42979,N_36139,N_38192);
and U42980 (N_42980,N_39642,N_37168);
and U42981 (N_42981,N_35088,N_38232);
or U42982 (N_42982,N_35291,N_39475);
xnor U42983 (N_42983,N_39022,N_37838);
nor U42984 (N_42984,N_35453,N_37053);
nor U42985 (N_42985,N_38214,N_39523);
xnor U42986 (N_42986,N_38584,N_37822);
nand U42987 (N_42987,N_39458,N_36656);
nor U42988 (N_42988,N_38530,N_35061);
or U42989 (N_42989,N_37327,N_38799);
nor U42990 (N_42990,N_37989,N_35532);
or U42991 (N_42991,N_36018,N_35528);
nor U42992 (N_42992,N_36273,N_38567);
xnor U42993 (N_42993,N_37093,N_35734);
xor U42994 (N_42994,N_36829,N_39951);
nand U42995 (N_42995,N_38444,N_38828);
nor U42996 (N_42996,N_35171,N_39949);
nor U42997 (N_42997,N_36814,N_39419);
or U42998 (N_42998,N_37836,N_35764);
or U42999 (N_42999,N_37655,N_35579);
or U43000 (N_43000,N_38830,N_37224);
and U43001 (N_43001,N_38103,N_35650);
and U43002 (N_43002,N_39001,N_36048);
xor U43003 (N_43003,N_35252,N_35915);
xnor U43004 (N_43004,N_35522,N_39368);
or U43005 (N_43005,N_39753,N_35548);
and U43006 (N_43006,N_38134,N_38328);
nor U43007 (N_43007,N_38947,N_39180);
and U43008 (N_43008,N_38056,N_38434);
or U43009 (N_43009,N_35579,N_35499);
nand U43010 (N_43010,N_35705,N_36135);
and U43011 (N_43011,N_39790,N_36762);
nor U43012 (N_43012,N_35159,N_35621);
nand U43013 (N_43013,N_37649,N_36330);
nor U43014 (N_43014,N_37937,N_36408);
nor U43015 (N_43015,N_36625,N_37065);
nor U43016 (N_43016,N_35091,N_37991);
and U43017 (N_43017,N_35358,N_35424);
or U43018 (N_43018,N_37238,N_36484);
nor U43019 (N_43019,N_37285,N_35690);
nand U43020 (N_43020,N_39716,N_36416);
nor U43021 (N_43021,N_35903,N_36529);
nand U43022 (N_43022,N_38635,N_36413);
or U43023 (N_43023,N_39754,N_37320);
nor U43024 (N_43024,N_39443,N_36689);
nor U43025 (N_43025,N_35135,N_38214);
nor U43026 (N_43026,N_37706,N_39004);
and U43027 (N_43027,N_36626,N_38956);
nor U43028 (N_43028,N_35376,N_38019);
nand U43029 (N_43029,N_39295,N_37934);
nor U43030 (N_43030,N_38767,N_37701);
nor U43031 (N_43031,N_38424,N_35036);
nand U43032 (N_43032,N_39310,N_35077);
nand U43033 (N_43033,N_37706,N_39277);
or U43034 (N_43034,N_37284,N_35058);
nand U43035 (N_43035,N_35223,N_39164);
xor U43036 (N_43036,N_37898,N_36173);
or U43037 (N_43037,N_39564,N_36207);
and U43038 (N_43038,N_37181,N_38890);
and U43039 (N_43039,N_39451,N_35679);
nand U43040 (N_43040,N_39128,N_36466);
and U43041 (N_43041,N_37613,N_38399);
or U43042 (N_43042,N_35106,N_38216);
nand U43043 (N_43043,N_39653,N_35368);
xnor U43044 (N_43044,N_38793,N_38161);
xnor U43045 (N_43045,N_38254,N_38975);
nor U43046 (N_43046,N_35538,N_38067);
nor U43047 (N_43047,N_35968,N_39350);
nand U43048 (N_43048,N_37078,N_37781);
nand U43049 (N_43049,N_37067,N_36182);
and U43050 (N_43050,N_38911,N_37795);
nand U43051 (N_43051,N_38498,N_38840);
or U43052 (N_43052,N_38436,N_38655);
xor U43053 (N_43053,N_36270,N_38169);
nand U43054 (N_43054,N_39959,N_37638);
nor U43055 (N_43055,N_37528,N_36451);
and U43056 (N_43056,N_39200,N_35005);
nand U43057 (N_43057,N_39111,N_37328);
and U43058 (N_43058,N_35956,N_36760);
nor U43059 (N_43059,N_35557,N_39043);
or U43060 (N_43060,N_35496,N_38918);
and U43061 (N_43061,N_39606,N_39430);
or U43062 (N_43062,N_37325,N_35640);
nor U43063 (N_43063,N_37037,N_38920);
xnor U43064 (N_43064,N_35244,N_38314);
nor U43065 (N_43065,N_39184,N_38931);
xor U43066 (N_43066,N_38328,N_39128);
and U43067 (N_43067,N_37665,N_38281);
nand U43068 (N_43068,N_35475,N_39363);
nor U43069 (N_43069,N_38599,N_37207);
xnor U43070 (N_43070,N_36437,N_36080);
or U43071 (N_43071,N_35818,N_39634);
xnor U43072 (N_43072,N_35281,N_35323);
and U43073 (N_43073,N_35412,N_39050);
xnor U43074 (N_43074,N_38538,N_35099);
xor U43075 (N_43075,N_35980,N_35740);
nor U43076 (N_43076,N_36511,N_38049);
nor U43077 (N_43077,N_36321,N_35745);
nand U43078 (N_43078,N_38315,N_35202);
nor U43079 (N_43079,N_37495,N_38375);
or U43080 (N_43080,N_39633,N_36714);
and U43081 (N_43081,N_38587,N_38132);
xor U43082 (N_43082,N_36822,N_39612);
xor U43083 (N_43083,N_36062,N_36544);
nor U43084 (N_43084,N_39224,N_36740);
or U43085 (N_43085,N_38359,N_37001);
or U43086 (N_43086,N_38208,N_39634);
or U43087 (N_43087,N_37544,N_37495);
xor U43088 (N_43088,N_37390,N_35919);
nor U43089 (N_43089,N_36266,N_35202);
or U43090 (N_43090,N_37634,N_36878);
nor U43091 (N_43091,N_38994,N_37152);
nand U43092 (N_43092,N_37939,N_36222);
xor U43093 (N_43093,N_36322,N_35390);
nand U43094 (N_43094,N_38653,N_38721);
xor U43095 (N_43095,N_35869,N_38735);
nor U43096 (N_43096,N_37650,N_38573);
nand U43097 (N_43097,N_38890,N_35274);
nor U43098 (N_43098,N_35286,N_38064);
nor U43099 (N_43099,N_38358,N_37155);
and U43100 (N_43100,N_35706,N_38698);
nor U43101 (N_43101,N_39157,N_39079);
nor U43102 (N_43102,N_38704,N_37185);
or U43103 (N_43103,N_39574,N_35993);
or U43104 (N_43104,N_38924,N_39813);
and U43105 (N_43105,N_37386,N_35533);
nor U43106 (N_43106,N_36784,N_37480);
xnor U43107 (N_43107,N_35596,N_38451);
nor U43108 (N_43108,N_36719,N_37043);
xnor U43109 (N_43109,N_39066,N_37070);
nor U43110 (N_43110,N_37177,N_35806);
nor U43111 (N_43111,N_39765,N_38259);
nor U43112 (N_43112,N_38316,N_35705);
nand U43113 (N_43113,N_36322,N_38411);
nand U43114 (N_43114,N_36592,N_38746);
or U43115 (N_43115,N_38622,N_35760);
or U43116 (N_43116,N_37401,N_38538);
or U43117 (N_43117,N_38944,N_35695);
xnor U43118 (N_43118,N_38148,N_39794);
nor U43119 (N_43119,N_39069,N_36479);
nor U43120 (N_43120,N_36483,N_37353);
and U43121 (N_43121,N_37411,N_39225);
nor U43122 (N_43122,N_35717,N_39094);
or U43123 (N_43123,N_37901,N_39026);
and U43124 (N_43124,N_38207,N_36367);
and U43125 (N_43125,N_37469,N_39377);
or U43126 (N_43126,N_36789,N_36324);
nand U43127 (N_43127,N_37812,N_38832);
xor U43128 (N_43128,N_37579,N_35763);
nor U43129 (N_43129,N_35738,N_36874);
xnor U43130 (N_43130,N_38140,N_39352);
or U43131 (N_43131,N_36589,N_39715);
nand U43132 (N_43132,N_39204,N_38961);
nand U43133 (N_43133,N_37274,N_37741);
nand U43134 (N_43134,N_37725,N_36386);
nor U43135 (N_43135,N_39525,N_38123);
xor U43136 (N_43136,N_38119,N_39854);
or U43137 (N_43137,N_38556,N_37800);
nor U43138 (N_43138,N_36741,N_35577);
or U43139 (N_43139,N_35974,N_39773);
xnor U43140 (N_43140,N_35973,N_39530);
nand U43141 (N_43141,N_37704,N_39921);
or U43142 (N_43142,N_38744,N_37162);
xnor U43143 (N_43143,N_36325,N_39297);
or U43144 (N_43144,N_35564,N_35838);
nand U43145 (N_43145,N_36762,N_36440);
nor U43146 (N_43146,N_38845,N_36387);
xnor U43147 (N_43147,N_35189,N_35464);
or U43148 (N_43148,N_36000,N_38120);
xnor U43149 (N_43149,N_36994,N_36190);
or U43150 (N_43150,N_36182,N_37971);
and U43151 (N_43151,N_36386,N_36627);
nor U43152 (N_43152,N_37854,N_36671);
xor U43153 (N_43153,N_37277,N_38092);
xor U43154 (N_43154,N_37477,N_37612);
nor U43155 (N_43155,N_35441,N_35361);
and U43156 (N_43156,N_39393,N_37240);
and U43157 (N_43157,N_36738,N_39062);
and U43158 (N_43158,N_38260,N_37013);
or U43159 (N_43159,N_35902,N_38557);
nand U43160 (N_43160,N_36212,N_36889);
nor U43161 (N_43161,N_36162,N_39955);
or U43162 (N_43162,N_38215,N_39807);
xnor U43163 (N_43163,N_36271,N_39639);
xnor U43164 (N_43164,N_37072,N_36249);
or U43165 (N_43165,N_37402,N_36707);
and U43166 (N_43166,N_38731,N_36647);
and U43167 (N_43167,N_37984,N_35850);
and U43168 (N_43168,N_36998,N_38501);
or U43169 (N_43169,N_39366,N_37349);
or U43170 (N_43170,N_36743,N_38801);
nand U43171 (N_43171,N_38077,N_38588);
nand U43172 (N_43172,N_39921,N_36363);
nor U43173 (N_43173,N_37363,N_35843);
or U43174 (N_43174,N_35539,N_37796);
xnor U43175 (N_43175,N_35499,N_39711);
nand U43176 (N_43176,N_36227,N_35167);
nor U43177 (N_43177,N_38827,N_36793);
and U43178 (N_43178,N_36747,N_39343);
xor U43179 (N_43179,N_38410,N_35642);
nor U43180 (N_43180,N_37493,N_36178);
nand U43181 (N_43181,N_36885,N_36584);
and U43182 (N_43182,N_39529,N_35636);
xor U43183 (N_43183,N_38076,N_36753);
and U43184 (N_43184,N_38394,N_39066);
and U43185 (N_43185,N_36106,N_38991);
or U43186 (N_43186,N_37879,N_39777);
nor U43187 (N_43187,N_37679,N_36373);
nor U43188 (N_43188,N_38577,N_35209);
or U43189 (N_43189,N_35125,N_35858);
or U43190 (N_43190,N_38420,N_39664);
nand U43191 (N_43191,N_38679,N_39729);
nand U43192 (N_43192,N_35342,N_38082);
nor U43193 (N_43193,N_39006,N_36674);
and U43194 (N_43194,N_36882,N_38637);
xor U43195 (N_43195,N_39438,N_39854);
xnor U43196 (N_43196,N_38405,N_35194);
and U43197 (N_43197,N_36675,N_37463);
nor U43198 (N_43198,N_37948,N_39805);
or U43199 (N_43199,N_39097,N_39159);
and U43200 (N_43200,N_35062,N_36626);
nor U43201 (N_43201,N_37578,N_37016);
or U43202 (N_43202,N_36543,N_38006);
nor U43203 (N_43203,N_35459,N_38126);
xor U43204 (N_43204,N_37051,N_35490);
and U43205 (N_43205,N_35546,N_37106);
nor U43206 (N_43206,N_36416,N_37628);
and U43207 (N_43207,N_37682,N_37916);
xnor U43208 (N_43208,N_35829,N_38015);
xor U43209 (N_43209,N_37064,N_35367);
and U43210 (N_43210,N_36413,N_36534);
nor U43211 (N_43211,N_38036,N_35553);
nor U43212 (N_43212,N_37903,N_37431);
xnor U43213 (N_43213,N_36649,N_36214);
nand U43214 (N_43214,N_37340,N_38946);
or U43215 (N_43215,N_39374,N_36801);
nand U43216 (N_43216,N_39260,N_37937);
xnor U43217 (N_43217,N_35502,N_36081);
nor U43218 (N_43218,N_39970,N_35292);
and U43219 (N_43219,N_37860,N_38144);
xnor U43220 (N_43220,N_37077,N_35053);
xnor U43221 (N_43221,N_39516,N_38245);
xor U43222 (N_43222,N_36951,N_38036);
or U43223 (N_43223,N_38742,N_38853);
or U43224 (N_43224,N_39453,N_38660);
nand U43225 (N_43225,N_35196,N_38600);
xor U43226 (N_43226,N_35322,N_37631);
and U43227 (N_43227,N_39861,N_36395);
and U43228 (N_43228,N_38603,N_39985);
or U43229 (N_43229,N_36991,N_39052);
nor U43230 (N_43230,N_36306,N_39253);
and U43231 (N_43231,N_39410,N_37997);
xor U43232 (N_43232,N_37345,N_38326);
or U43233 (N_43233,N_36906,N_38625);
and U43234 (N_43234,N_38180,N_39271);
nor U43235 (N_43235,N_38177,N_35908);
and U43236 (N_43236,N_37970,N_37758);
or U43237 (N_43237,N_38024,N_37800);
xnor U43238 (N_43238,N_35517,N_36160);
or U43239 (N_43239,N_37818,N_38276);
and U43240 (N_43240,N_39663,N_39253);
or U43241 (N_43241,N_37834,N_39977);
or U43242 (N_43242,N_36140,N_37243);
nor U43243 (N_43243,N_39819,N_35281);
nand U43244 (N_43244,N_36291,N_35915);
nand U43245 (N_43245,N_39850,N_38864);
xnor U43246 (N_43246,N_38960,N_36373);
xor U43247 (N_43247,N_39168,N_36926);
xnor U43248 (N_43248,N_38068,N_39874);
or U43249 (N_43249,N_36924,N_36213);
nor U43250 (N_43250,N_38670,N_35010);
nor U43251 (N_43251,N_35761,N_39602);
nor U43252 (N_43252,N_39614,N_36397);
xor U43253 (N_43253,N_37002,N_38434);
and U43254 (N_43254,N_38127,N_36957);
nor U43255 (N_43255,N_35887,N_35102);
nand U43256 (N_43256,N_37916,N_36545);
xor U43257 (N_43257,N_39108,N_38759);
or U43258 (N_43258,N_38168,N_37547);
or U43259 (N_43259,N_37726,N_39317);
nand U43260 (N_43260,N_36798,N_38653);
xnor U43261 (N_43261,N_39432,N_36725);
and U43262 (N_43262,N_35055,N_39442);
or U43263 (N_43263,N_39120,N_36205);
and U43264 (N_43264,N_36094,N_38622);
and U43265 (N_43265,N_35793,N_35992);
nor U43266 (N_43266,N_36219,N_39861);
and U43267 (N_43267,N_38916,N_38845);
xnor U43268 (N_43268,N_35215,N_36745);
xnor U43269 (N_43269,N_37983,N_37730);
or U43270 (N_43270,N_39882,N_36753);
nor U43271 (N_43271,N_36205,N_38053);
xnor U43272 (N_43272,N_39847,N_36798);
xor U43273 (N_43273,N_35915,N_39218);
nor U43274 (N_43274,N_39714,N_39577);
or U43275 (N_43275,N_37739,N_35062);
or U43276 (N_43276,N_36177,N_39069);
xnor U43277 (N_43277,N_38475,N_39372);
xor U43278 (N_43278,N_36537,N_39776);
or U43279 (N_43279,N_36863,N_36494);
xor U43280 (N_43280,N_36362,N_38513);
nor U43281 (N_43281,N_35889,N_35806);
xor U43282 (N_43282,N_37833,N_36641);
nor U43283 (N_43283,N_36687,N_38391);
and U43284 (N_43284,N_35673,N_37637);
and U43285 (N_43285,N_37411,N_36763);
or U43286 (N_43286,N_39114,N_37613);
xor U43287 (N_43287,N_38488,N_38793);
nor U43288 (N_43288,N_39241,N_38344);
or U43289 (N_43289,N_36662,N_38451);
nand U43290 (N_43290,N_37787,N_37339);
and U43291 (N_43291,N_38841,N_36969);
xnor U43292 (N_43292,N_37312,N_37550);
or U43293 (N_43293,N_35946,N_37204);
nand U43294 (N_43294,N_38441,N_35115);
or U43295 (N_43295,N_35013,N_39756);
or U43296 (N_43296,N_36788,N_36174);
nand U43297 (N_43297,N_35955,N_38209);
nor U43298 (N_43298,N_39871,N_35076);
nand U43299 (N_43299,N_37597,N_39842);
nand U43300 (N_43300,N_36838,N_37748);
or U43301 (N_43301,N_38829,N_38447);
nand U43302 (N_43302,N_35277,N_35641);
xor U43303 (N_43303,N_35720,N_39580);
nand U43304 (N_43304,N_36755,N_35330);
or U43305 (N_43305,N_36568,N_38686);
and U43306 (N_43306,N_37471,N_39892);
xnor U43307 (N_43307,N_39189,N_36514);
xor U43308 (N_43308,N_35998,N_35830);
nand U43309 (N_43309,N_37559,N_36134);
or U43310 (N_43310,N_37666,N_39269);
or U43311 (N_43311,N_39414,N_37213);
or U43312 (N_43312,N_38652,N_38162);
or U43313 (N_43313,N_38097,N_39435);
nor U43314 (N_43314,N_35306,N_37588);
xor U43315 (N_43315,N_39245,N_39016);
nor U43316 (N_43316,N_37870,N_39893);
nor U43317 (N_43317,N_36216,N_39919);
and U43318 (N_43318,N_37495,N_38519);
nand U43319 (N_43319,N_37443,N_35567);
and U43320 (N_43320,N_37801,N_35922);
and U43321 (N_43321,N_39948,N_36256);
nor U43322 (N_43322,N_38452,N_37861);
or U43323 (N_43323,N_39549,N_39783);
or U43324 (N_43324,N_36546,N_38176);
and U43325 (N_43325,N_36808,N_38217);
or U43326 (N_43326,N_37134,N_35741);
nor U43327 (N_43327,N_37924,N_38698);
nand U43328 (N_43328,N_36885,N_39458);
and U43329 (N_43329,N_35530,N_36436);
or U43330 (N_43330,N_39005,N_35673);
xor U43331 (N_43331,N_35941,N_35563);
nor U43332 (N_43332,N_36500,N_38499);
or U43333 (N_43333,N_37606,N_38368);
nand U43334 (N_43334,N_38819,N_38323);
xor U43335 (N_43335,N_35060,N_38160);
xnor U43336 (N_43336,N_39050,N_38386);
nand U43337 (N_43337,N_35077,N_36982);
nand U43338 (N_43338,N_35075,N_36940);
or U43339 (N_43339,N_35617,N_35815);
or U43340 (N_43340,N_35800,N_36303);
or U43341 (N_43341,N_38543,N_37056);
nor U43342 (N_43342,N_38531,N_37993);
and U43343 (N_43343,N_35938,N_39547);
xor U43344 (N_43344,N_37914,N_39928);
or U43345 (N_43345,N_35063,N_36332);
nor U43346 (N_43346,N_38007,N_36856);
xnor U43347 (N_43347,N_38242,N_36798);
and U43348 (N_43348,N_38226,N_39850);
or U43349 (N_43349,N_38693,N_39479);
or U43350 (N_43350,N_37392,N_38025);
or U43351 (N_43351,N_38946,N_36630);
or U43352 (N_43352,N_39394,N_37920);
nand U43353 (N_43353,N_39619,N_37705);
nand U43354 (N_43354,N_39005,N_38472);
nand U43355 (N_43355,N_36222,N_39270);
or U43356 (N_43356,N_37795,N_39331);
nor U43357 (N_43357,N_36617,N_36725);
or U43358 (N_43358,N_35063,N_38781);
or U43359 (N_43359,N_39251,N_37844);
nand U43360 (N_43360,N_35725,N_39203);
nor U43361 (N_43361,N_39604,N_35511);
nand U43362 (N_43362,N_39332,N_39556);
nor U43363 (N_43363,N_37763,N_39049);
nor U43364 (N_43364,N_38281,N_37172);
nor U43365 (N_43365,N_35199,N_39397);
nor U43366 (N_43366,N_38295,N_38429);
nor U43367 (N_43367,N_39727,N_38247);
or U43368 (N_43368,N_37085,N_36249);
or U43369 (N_43369,N_39193,N_38522);
nand U43370 (N_43370,N_36317,N_36903);
or U43371 (N_43371,N_37926,N_35421);
nor U43372 (N_43372,N_37561,N_39738);
xnor U43373 (N_43373,N_37725,N_37524);
nor U43374 (N_43374,N_35764,N_37470);
nor U43375 (N_43375,N_37436,N_36179);
and U43376 (N_43376,N_37952,N_37962);
xor U43377 (N_43377,N_39345,N_36646);
or U43378 (N_43378,N_36645,N_36474);
nand U43379 (N_43379,N_39860,N_38017);
and U43380 (N_43380,N_35029,N_36960);
nand U43381 (N_43381,N_35170,N_35520);
nor U43382 (N_43382,N_37481,N_35170);
or U43383 (N_43383,N_38329,N_36869);
nor U43384 (N_43384,N_37216,N_35428);
nor U43385 (N_43385,N_35767,N_35892);
nor U43386 (N_43386,N_39829,N_37970);
nor U43387 (N_43387,N_36899,N_35294);
or U43388 (N_43388,N_35852,N_35702);
and U43389 (N_43389,N_37806,N_37691);
or U43390 (N_43390,N_38418,N_39716);
and U43391 (N_43391,N_38003,N_35987);
xnor U43392 (N_43392,N_39135,N_36864);
or U43393 (N_43393,N_37898,N_38898);
nor U43394 (N_43394,N_35355,N_37358);
or U43395 (N_43395,N_39818,N_35808);
xor U43396 (N_43396,N_39783,N_37146);
xor U43397 (N_43397,N_36781,N_35024);
or U43398 (N_43398,N_39843,N_37647);
nor U43399 (N_43399,N_39867,N_37789);
nor U43400 (N_43400,N_35402,N_39665);
nor U43401 (N_43401,N_35088,N_39575);
or U43402 (N_43402,N_39440,N_37930);
xor U43403 (N_43403,N_39028,N_37824);
and U43404 (N_43404,N_37259,N_39226);
nor U43405 (N_43405,N_37439,N_39168);
or U43406 (N_43406,N_39254,N_37015);
xnor U43407 (N_43407,N_36309,N_39050);
xor U43408 (N_43408,N_39966,N_37073);
or U43409 (N_43409,N_39446,N_37542);
and U43410 (N_43410,N_37777,N_35751);
xnor U43411 (N_43411,N_37415,N_35875);
or U43412 (N_43412,N_36974,N_35507);
and U43413 (N_43413,N_35119,N_38804);
or U43414 (N_43414,N_35104,N_37922);
nor U43415 (N_43415,N_35326,N_39555);
xnor U43416 (N_43416,N_35539,N_39282);
nor U43417 (N_43417,N_35650,N_39215);
nand U43418 (N_43418,N_35101,N_39494);
xor U43419 (N_43419,N_37701,N_36580);
and U43420 (N_43420,N_36308,N_36304);
and U43421 (N_43421,N_37156,N_38879);
nand U43422 (N_43422,N_35158,N_36768);
or U43423 (N_43423,N_35428,N_36195);
nor U43424 (N_43424,N_39057,N_38949);
xnor U43425 (N_43425,N_38589,N_36838);
nor U43426 (N_43426,N_36494,N_38805);
nand U43427 (N_43427,N_35716,N_39134);
nand U43428 (N_43428,N_36782,N_38969);
or U43429 (N_43429,N_35036,N_39044);
xor U43430 (N_43430,N_39677,N_36022);
nor U43431 (N_43431,N_36878,N_39107);
and U43432 (N_43432,N_38544,N_37262);
nand U43433 (N_43433,N_37826,N_36612);
nor U43434 (N_43434,N_35359,N_37181);
nor U43435 (N_43435,N_39079,N_39054);
nor U43436 (N_43436,N_36756,N_35427);
and U43437 (N_43437,N_37439,N_39269);
and U43438 (N_43438,N_35885,N_35062);
xor U43439 (N_43439,N_37983,N_39858);
or U43440 (N_43440,N_36338,N_37453);
nand U43441 (N_43441,N_39071,N_37144);
nand U43442 (N_43442,N_35490,N_35065);
nand U43443 (N_43443,N_36175,N_35243);
nor U43444 (N_43444,N_36056,N_37522);
xor U43445 (N_43445,N_35044,N_36621);
and U43446 (N_43446,N_38702,N_38357);
or U43447 (N_43447,N_37379,N_35530);
nand U43448 (N_43448,N_35054,N_37772);
nand U43449 (N_43449,N_37036,N_37990);
xor U43450 (N_43450,N_35929,N_39227);
and U43451 (N_43451,N_38456,N_39676);
xor U43452 (N_43452,N_38160,N_37792);
or U43453 (N_43453,N_35744,N_39944);
nor U43454 (N_43454,N_37915,N_36603);
nor U43455 (N_43455,N_36833,N_35633);
nand U43456 (N_43456,N_36231,N_39404);
nor U43457 (N_43457,N_36929,N_35490);
xnor U43458 (N_43458,N_38230,N_36651);
and U43459 (N_43459,N_37855,N_36238);
and U43460 (N_43460,N_37309,N_37518);
or U43461 (N_43461,N_35482,N_37728);
nor U43462 (N_43462,N_36077,N_38880);
xor U43463 (N_43463,N_35104,N_37817);
nor U43464 (N_43464,N_36841,N_36341);
or U43465 (N_43465,N_35406,N_39398);
and U43466 (N_43466,N_37372,N_37523);
xor U43467 (N_43467,N_37774,N_36350);
nor U43468 (N_43468,N_36342,N_38319);
and U43469 (N_43469,N_36428,N_39809);
or U43470 (N_43470,N_38322,N_39756);
and U43471 (N_43471,N_38113,N_35884);
or U43472 (N_43472,N_38288,N_36410);
and U43473 (N_43473,N_35429,N_35084);
and U43474 (N_43474,N_37167,N_38486);
and U43475 (N_43475,N_36121,N_36163);
and U43476 (N_43476,N_37513,N_35640);
or U43477 (N_43477,N_36137,N_38787);
xor U43478 (N_43478,N_36415,N_37344);
or U43479 (N_43479,N_38197,N_38345);
nand U43480 (N_43480,N_37221,N_39489);
nand U43481 (N_43481,N_35237,N_35572);
nor U43482 (N_43482,N_35854,N_37117);
nor U43483 (N_43483,N_36975,N_36440);
xor U43484 (N_43484,N_36403,N_39677);
or U43485 (N_43485,N_35511,N_38544);
nor U43486 (N_43486,N_37986,N_36820);
nand U43487 (N_43487,N_35097,N_39130);
nor U43488 (N_43488,N_39951,N_35379);
nand U43489 (N_43489,N_37324,N_36864);
and U43490 (N_43490,N_37525,N_35135);
and U43491 (N_43491,N_37243,N_37604);
and U43492 (N_43492,N_39014,N_35016);
or U43493 (N_43493,N_39653,N_36217);
nand U43494 (N_43494,N_39585,N_38581);
nand U43495 (N_43495,N_35813,N_39652);
or U43496 (N_43496,N_38910,N_36669);
and U43497 (N_43497,N_39512,N_35791);
or U43498 (N_43498,N_39307,N_38400);
nor U43499 (N_43499,N_39168,N_37506);
nand U43500 (N_43500,N_36687,N_36818);
nand U43501 (N_43501,N_39497,N_37020);
or U43502 (N_43502,N_38659,N_35975);
nand U43503 (N_43503,N_39998,N_37562);
nor U43504 (N_43504,N_36053,N_38679);
or U43505 (N_43505,N_37528,N_36933);
nor U43506 (N_43506,N_36266,N_35441);
and U43507 (N_43507,N_39375,N_39252);
or U43508 (N_43508,N_39092,N_37587);
xor U43509 (N_43509,N_35386,N_36830);
and U43510 (N_43510,N_37467,N_38419);
nor U43511 (N_43511,N_37347,N_36715);
xnor U43512 (N_43512,N_37285,N_39582);
xor U43513 (N_43513,N_36905,N_37049);
nor U43514 (N_43514,N_35252,N_35969);
or U43515 (N_43515,N_37640,N_39763);
nor U43516 (N_43516,N_39569,N_37389);
nand U43517 (N_43517,N_38197,N_37744);
nand U43518 (N_43518,N_35839,N_36068);
and U43519 (N_43519,N_38928,N_37134);
xor U43520 (N_43520,N_39054,N_39194);
xor U43521 (N_43521,N_38155,N_38044);
nor U43522 (N_43522,N_38786,N_38283);
or U43523 (N_43523,N_36821,N_39769);
or U43524 (N_43524,N_39463,N_35960);
and U43525 (N_43525,N_39897,N_35779);
nand U43526 (N_43526,N_38392,N_36598);
nor U43527 (N_43527,N_36081,N_38653);
nand U43528 (N_43528,N_35224,N_35771);
nand U43529 (N_43529,N_39941,N_38813);
xor U43530 (N_43530,N_39105,N_39602);
or U43531 (N_43531,N_39399,N_38083);
nor U43532 (N_43532,N_36744,N_35408);
nor U43533 (N_43533,N_38044,N_36949);
xnor U43534 (N_43534,N_37211,N_36115);
nand U43535 (N_43535,N_35172,N_39588);
or U43536 (N_43536,N_37701,N_39703);
nor U43537 (N_43537,N_39203,N_39334);
or U43538 (N_43538,N_35695,N_36216);
nor U43539 (N_43539,N_37862,N_39124);
nor U43540 (N_43540,N_38176,N_38251);
or U43541 (N_43541,N_35262,N_37359);
nor U43542 (N_43542,N_38149,N_37579);
and U43543 (N_43543,N_38808,N_39331);
or U43544 (N_43544,N_37891,N_39442);
nand U43545 (N_43545,N_36502,N_38552);
xor U43546 (N_43546,N_39053,N_39451);
nor U43547 (N_43547,N_38206,N_39865);
nor U43548 (N_43548,N_38436,N_36595);
or U43549 (N_43549,N_35897,N_39399);
nor U43550 (N_43550,N_36358,N_37766);
nand U43551 (N_43551,N_39561,N_36339);
xnor U43552 (N_43552,N_35576,N_35740);
and U43553 (N_43553,N_38525,N_37058);
and U43554 (N_43554,N_37524,N_37939);
and U43555 (N_43555,N_35321,N_37541);
or U43556 (N_43556,N_38421,N_38494);
and U43557 (N_43557,N_39300,N_35185);
nand U43558 (N_43558,N_35279,N_39524);
nand U43559 (N_43559,N_39006,N_37961);
or U43560 (N_43560,N_37866,N_38616);
xor U43561 (N_43561,N_37229,N_38948);
xnor U43562 (N_43562,N_35607,N_39630);
xor U43563 (N_43563,N_35825,N_36339);
nand U43564 (N_43564,N_35737,N_35800);
nand U43565 (N_43565,N_38718,N_37776);
or U43566 (N_43566,N_38702,N_35274);
xnor U43567 (N_43567,N_36254,N_38639);
nand U43568 (N_43568,N_35471,N_36698);
and U43569 (N_43569,N_35203,N_35032);
nor U43570 (N_43570,N_36595,N_37507);
and U43571 (N_43571,N_37523,N_37804);
nand U43572 (N_43572,N_36317,N_39242);
nor U43573 (N_43573,N_36234,N_39826);
nand U43574 (N_43574,N_39096,N_39766);
xnor U43575 (N_43575,N_39905,N_38628);
or U43576 (N_43576,N_38104,N_35914);
nand U43577 (N_43577,N_35957,N_36764);
or U43578 (N_43578,N_37835,N_35329);
xnor U43579 (N_43579,N_35636,N_39493);
or U43580 (N_43580,N_37483,N_39452);
xnor U43581 (N_43581,N_38151,N_39173);
nor U43582 (N_43582,N_35932,N_39694);
or U43583 (N_43583,N_36165,N_35682);
nand U43584 (N_43584,N_38710,N_37372);
or U43585 (N_43585,N_39568,N_38161);
nand U43586 (N_43586,N_38701,N_36091);
nor U43587 (N_43587,N_36353,N_35926);
and U43588 (N_43588,N_39565,N_37519);
nand U43589 (N_43589,N_35717,N_39151);
nor U43590 (N_43590,N_35852,N_37530);
nor U43591 (N_43591,N_35557,N_37070);
xnor U43592 (N_43592,N_37107,N_39665);
nor U43593 (N_43593,N_35516,N_35840);
or U43594 (N_43594,N_38816,N_38800);
or U43595 (N_43595,N_38319,N_36831);
nand U43596 (N_43596,N_36982,N_39422);
nand U43597 (N_43597,N_36207,N_38231);
xnor U43598 (N_43598,N_39567,N_37685);
xor U43599 (N_43599,N_37232,N_38881);
xor U43600 (N_43600,N_35274,N_39334);
and U43601 (N_43601,N_39865,N_39041);
nand U43602 (N_43602,N_38551,N_35453);
nor U43603 (N_43603,N_38718,N_39617);
nand U43604 (N_43604,N_39550,N_37299);
or U43605 (N_43605,N_37314,N_38666);
nand U43606 (N_43606,N_38251,N_38543);
and U43607 (N_43607,N_38418,N_39425);
xnor U43608 (N_43608,N_35218,N_38718);
nor U43609 (N_43609,N_37124,N_38298);
nand U43610 (N_43610,N_37338,N_37292);
or U43611 (N_43611,N_38730,N_38742);
nor U43612 (N_43612,N_36990,N_37352);
or U43613 (N_43613,N_39827,N_37055);
xnor U43614 (N_43614,N_38500,N_35140);
xor U43615 (N_43615,N_37518,N_39062);
and U43616 (N_43616,N_35901,N_37349);
nor U43617 (N_43617,N_39008,N_37128);
and U43618 (N_43618,N_35967,N_37543);
xor U43619 (N_43619,N_37689,N_36246);
nor U43620 (N_43620,N_39613,N_37949);
nand U43621 (N_43621,N_35540,N_39569);
nand U43622 (N_43622,N_38192,N_36135);
or U43623 (N_43623,N_36458,N_36428);
xnor U43624 (N_43624,N_35581,N_38053);
xor U43625 (N_43625,N_35376,N_35624);
nor U43626 (N_43626,N_36333,N_35454);
xor U43627 (N_43627,N_37700,N_39230);
and U43628 (N_43628,N_36740,N_36939);
or U43629 (N_43629,N_35326,N_35866);
and U43630 (N_43630,N_37498,N_35002);
and U43631 (N_43631,N_37125,N_36992);
nand U43632 (N_43632,N_38986,N_36454);
and U43633 (N_43633,N_36453,N_39716);
nor U43634 (N_43634,N_36291,N_37748);
xor U43635 (N_43635,N_37691,N_36947);
nor U43636 (N_43636,N_35333,N_39684);
or U43637 (N_43637,N_37044,N_37741);
nand U43638 (N_43638,N_39613,N_36380);
and U43639 (N_43639,N_39081,N_39251);
and U43640 (N_43640,N_39756,N_36968);
nand U43641 (N_43641,N_37647,N_39921);
and U43642 (N_43642,N_39337,N_38925);
and U43643 (N_43643,N_39261,N_35806);
and U43644 (N_43644,N_37433,N_39290);
nand U43645 (N_43645,N_39188,N_38311);
xnor U43646 (N_43646,N_36129,N_37484);
nand U43647 (N_43647,N_35638,N_38710);
nor U43648 (N_43648,N_38413,N_37942);
or U43649 (N_43649,N_35750,N_35008);
and U43650 (N_43650,N_39063,N_39624);
and U43651 (N_43651,N_38548,N_39102);
and U43652 (N_43652,N_37905,N_37703);
or U43653 (N_43653,N_38664,N_37070);
and U43654 (N_43654,N_37867,N_38256);
or U43655 (N_43655,N_38945,N_38889);
xnor U43656 (N_43656,N_35563,N_35125);
or U43657 (N_43657,N_36792,N_36894);
nand U43658 (N_43658,N_38502,N_38229);
nor U43659 (N_43659,N_35846,N_39539);
nand U43660 (N_43660,N_38748,N_36065);
nor U43661 (N_43661,N_39693,N_36003);
nand U43662 (N_43662,N_39995,N_36225);
nor U43663 (N_43663,N_36435,N_38832);
nor U43664 (N_43664,N_37506,N_36231);
and U43665 (N_43665,N_36888,N_35779);
xnor U43666 (N_43666,N_36891,N_38724);
xor U43667 (N_43667,N_38340,N_35702);
nand U43668 (N_43668,N_36875,N_38923);
nand U43669 (N_43669,N_39516,N_38215);
or U43670 (N_43670,N_35843,N_39923);
nand U43671 (N_43671,N_38476,N_39757);
nor U43672 (N_43672,N_37305,N_37283);
and U43673 (N_43673,N_39072,N_39672);
nand U43674 (N_43674,N_35885,N_35147);
and U43675 (N_43675,N_37397,N_36111);
nor U43676 (N_43676,N_38251,N_35169);
xnor U43677 (N_43677,N_38303,N_39105);
xnor U43678 (N_43678,N_36494,N_39046);
xnor U43679 (N_43679,N_36082,N_35386);
nor U43680 (N_43680,N_35862,N_38873);
nand U43681 (N_43681,N_36775,N_38950);
xor U43682 (N_43682,N_37680,N_36031);
and U43683 (N_43683,N_37460,N_35253);
or U43684 (N_43684,N_36138,N_36865);
and U43685 (N_43685,N_36380,N_36082);
and U43686 (N_43686,N_38007,N_38496);
and U43687 (N_43687,N_37007,N_38829);
nor U43688 (N_43688,N_38644,N_35249);
nor U43689 (N_43689,N_36160,N_35230);
and U43690 (N_43690,N_36079,N_37031);
or U43691 (N_43691,N_35337,N_36960);
xnor U43692 (N_43692,N_38112,N_38286);
nand U43693 (N_43693,N_35439,N_38653);
xnor U43694 (N_43694,N_38081,N_38560);
nor U43695 (N_43695,N_36232,N_37528);
or U43696 (N_43696,N_39242,N_36034);
or U43697 (N_43697,N_38889,N_36526);
or U43698 (N_43698,N_39422,N_35917);
nor U43699 (N_43699,N_37216,N_38671);
or U43700 (N_43700,N_38852,N_39512);
nor U43701 (N_43701,N_37709,N_36929);
xnor U43702 (N_43702,N_38716,N_39526);
nand U43703 (N_43703,N_38349,N_39698);
and U43704 (N_43704,N_37445,N_39327);
or U43705 (N_43705,N_39112,N_37279);
or U43706 (N_43706,N_37673,N_39289);
nor U43707 (N_43707,N_36336,N_37409);
xor U43708 (N_43708,N_36862,N_39291);
or U43709 (N_43709,N_35104,N_39637);
nand U43710 (N_43710,N_39610,N_37424);
or U43711 (N_43711,N_36017,N_37529);
or U43712 (N_43712,N_35762,N_39788);
or U43713 (N_43713,N_36287,N_36227);
or U43714 (N_43714,N_37834,N_39502);
nor U43715 (N_43715,N_38992,N_35079);
xor U43716 (N_43716,N_39745,N_35800);
or U43717 (N_43717,N_37467,N_37257);
or U43718 (N_43718,N_35185,N_36330);
xnor U43719 (N_43719,N_36590,N_39500);
nand U43720 (N_43720,N_39468,N_39996);
nand U43721 (N_43721,N_36443,N_38562);
nand U43722 (N_43722,N_38675,N_36882);
nand U43723 (N_43723,N_36730,N_39055);
and U43724 (N_43724,N_38015,N_38459);
or U43725 (N_43725,N_38670,N_38910);
and U43726 (N_43726,N_35783,N_37305);
or U43727 (N_43727,N_39715,N_39518);
xor U43728 (N_43728,N_35381,N_39172);
nor U43729 (N_43729,N_38587,N_39398);
nand U43730 (N_43730,N_38651,N_38669);
xnor U43731 (N_43731,N_37328,N_37111);
nand U43732 (N_43732,N_35748,N_37668);
xnor U43733 (N_43733,N_38378,N_38392);
or U43734 (N_43734,N_36579,N_35714);
xor U43735 (N_43735,N_35946,N_38508);
or U43736 (N_43736,N_35375,N_35255);
and U43737 (N_43737,N_35823,N_39297);
nor U43738 (N_43738,N_36016,N_36937);
nand U43739 (N_43739,N_39357,N_37423);
xor U43740 (N_43740,N_37197,N_38576);
nor U43741 (N_43741,N_37202,N_35233);
xor U43742 (N_43742,N_39869,N_36020);
nor U43743 (N_43743,N_38093,N_39938);
xor U43744 (N_43744,N_37031,N_37843);
nand U43745 (N_43745,N_37701,N_38138);
nand U43746 (N_43746,N_37478,N_38771);
or U43747 (N_43747,N_36507,N_37843);
or U43748 (N_43748,N_39080,N_37185);
and U43749 (N_43749,N_38820,N_35691);
xor U43750 (N_43750,N_38594,N_36184);
and U43751 (N_43751,N_38710,N_36338);
or U43752 (N_43752,N_37704,N_35505);
or U43753 (N_43753,N_37478,N_36193);
and U43754 (N_43754,N_36771,N_36166);
xnor U43755 (N_43755,N_35317,N_39060);
xor U43756 (N_43756,N_39032,N_39348);
nor U43757 (N_43757,N_39401,N_38781);
nor U43758 (N_43758,N_36822,N_38887);
and U43759 (N_43759,N_38933,N_36923);
and U43760 (N_43760,N_39436,N_35013);
and U43761 (N_43761,N_39761,N_38267);
xnor U43762 (N_43762,N_37458,N_38006);
and U43763 (N_43763,N_39324,N_36201);
xor U43764 (N_43764,N_37986,N_38359);
or U43765 (N_43765,N_39969,N_38018);
xnor U43766 (N_43766,N_39362,N_37664);
and U43767 (N_43767,N_35812,N_38360);
nand U43768 (N_43768,N_37263,N_36886);
xor U43769 (N_43769,N_38014,N_38281);
xnor U43770 (N_43770,N_37970,N_35076);
nor U43771 (N_43771,N_39130,N_38228);
xnor U43772 (N_43772,N_35474,N_35423);
nor U43773 (N_43773,N_37761,N_38046);
nor U43774 (N_43774,N_39089,N_36076);
or U43775 (N_43775,N_37383,N_39314);
nor U43776 (N_43776,N_39322,N_37446);
or U43777 (N_43777,N_37649,N_37111);
nor U43778 (N_43778,N_39320,N_36706);
nand U43779 (N_43779,N_37579,N_35252);
and U43780 (N_43780,N_36025,N_36535);
and U43781 (N_43781,N_36009,N_38288);
and U43782 (N_43782,N_38116,N_38338);
xnor U43783 (N_43783,N_35011,N_35397);
nor U43784 (N_43784,N_38747,N_39489);
xor U43785 (N_43785,N_37361,N_38574);
and U43786 (N_43786,N_38839,N_36888);
nand U43787 (N_43787,N_36908,N_38927);
or U43788 (N_43788,N_38365,N_37103);
xnor U43789 (N_43789,N_36070,N_35326);
or U43790 (N_43790,N_36694,N_38873);
xnor U43791 (N_43791,N_35470,N_38996);
nand U43792 (N_43792,N_37756,N_39029);
or U43793 (N_43793,N_35533,N_35572);
nand U43794 (N_43794,N_39051,N_36907);
nand U43795 (N_43795,N_39336,N_37377);
xnor U43796 (N_43796,N_35184,N_35273);
nand U43797 (N_43797,N_38742,N_39068);
xor U43798 (N_43798,N_37248,N_35073);
xnor U43799 (N_43799,N_35727,N_38380);
nand U43800 (N_43800,N_39899,N_39166);
nand U43801 (N_43801,N_39082,N_38009);
nor U43802 (N_43802,N_37347,N_39042);
nand U43803 (N_43803,N_37100,N_35637);
or U43804 (N_43804,N_36453,N_35119);
or U43805 (N_43805,N_39055,N_38381);
and U43806 (N_43806,N_39001,N_35578);
or U43807 (N_43807,N_37887,N_37861);
or U43808 (N_43808,N_36175,N_36787);
nor U43809 (N_43809,N_35643,N_37832);
or U43810 (N_43810,N_35905,N_39729);
nand U43811 (N_43811,N_38263,N_35955);
nor U43812 (N_43812,N_36343,N_39402);
or U43813 (N_43813,N_37417,N_36641);
and U43814 (N_43814,N_38038,N_36917);
or U43815 (N_43815,N_37450,N_36457);
or U43816 (N_43816,N_39121,N_39423);
nor U43817 (N_43817,N_37880,N_36747);
nand U43818 (N_43818,N_35096,N_35848);
or U43819 (N_43819,N_38442,N_39421);
or U43820 (N_43820,N_35869,N_39953);
nand U43821 (N_43821,N_35409,N_36373);
nand U43822 (N_43822,N_36564,N_36079);
nor U43823 (N_43823,N_39177,N_39448);
nor U43824 (N_43824,N_37929,N_39412);
xor U43825 (N_43825,N_38359,N_36115);
xnor U43826 (N_43826,N_36628,N_37489);
or U43827 (N_43827,N_35699,N_38032);
xor U43828 (N_43828,N_38284,N_37906);
nor U43829 (N_43829,N_35456,N_37711);
xor U43830 (N_43830,N_36086,N_38292);
and U43831 (N_43831,N_36876,N_35749);
and U43832 (N_43832,N_36520,N_39968);
or U43833 (N_43833,N_35425,N_37756);
and U43834 (N_43834,N_35476,N_38751);
nand U43835 (N_43835,N_37511,N_35614);
and U43836 (N_43836,N_39706,N_37961);
and U43837 (N_43837,N_35254,N_36662);
or U43838 (N_43838,N_36714,N_36048);
or U43839 (N_43839,N_39425,N_35075);
or U43840 (N_43840,N_35271,N_37539);
nand U43841 (N_43841,N_38803,N_38535);
xnor U43842 (N_43842,N_39821,N_37577);
nand U43843 (N_43843,N_35030,N_36704);
nor U43844 (N_43844,N_37094,N_36846);
or U43845 (N_43845,N_37924,N_37374);
nand U43846 (N_43846,N_37791,N_35940);
nand U43847 (N_43847,N_35956,N_36759);
nor U43848 (N_43848,N_37202,N_39409);
nor U43849 (N_43849,N_35941,N_39177);
xor U43850 (N_43850,N_37897,N_39767);
nor U43851 (N_43851,N_37243,N_38652);
and U43852 (N_43852,N_39375,N_38068);
nand U43853 (N_43853,N_38898,N_35370);
nand U43854 (N_43854,N_36770,N_39415);
xnor U43855 (N_43855,N_36316,N_38491);
nand U43856 (N_43856,N_35946,N_39813);
xor U43857 (N_43857,N_36738,N_35758);
or U43858 (N_43858,N_35992,N_35796);
or U43859 (N_43859,N_38387,N_37571);
xor U43860 (N_43860,N_35572,N_37288);
and U43861 (N_43861,N_37067,N_39587);
nand U43862 (N_43862,N_39608,N_38743);
and U43863 (N_43863,N_36326,N_39943);
nand U43864 (N_43864,N_36174,N_35481);
nor U43865 (N_43865,N_38098,N_38537);
or U43866 (N_43866,N_35402,N_36058);
and U43867 (N_43867,N_36856,N_38665);
nand U43868 (N_43868,N_37589,N_39063);
nand U43869 (N_43869,N_35126,N_37598);
nand U43870 (N_43870,N_37038,N_39767);
nand U43871 (N_43871,N_36959,N_38228);
xnor U43872 (N_43872,N_39043,N_36728);
nor U43873 (N_43873,N_36700,N_38186);
xnor U43874 (N_43874,N_35576,N_37816);
xnor U43875 (N_43875,N_38297,N_38662);
xnor U43876 (N_43876,N_36769,N_36980);
xor U43877 (N_43877,N_36671,N_38629);
nand U43878 (N_43878,N_39558,N_39146);
or U43879 (N_43879,N_38107,N_37190);
and U43880 (N_43880,N_37420,N_35450);
or U43881 (N_43881,N_37053,N_37261);
nand U43882 (N_43882,N_36713,N_39845);
xnor U43883 (N_43883,N_37103,N_37059);
nand U43884 (N_43884,N_38030,N_37605);
or U43885 (N_43885,N_36085,N_35362);
nand U43886 (N_43886,N_35577,N_38398);
xnor U43887 (N_43887,N_35476,N_37657);
or U43888 (N_43888,N_35757,N_35802);
or U43889 (N_43889,N_35806,N_37588);
and U43890 (N_43890,N_38558,N_36819);
nor U43891 (N_43891,N_39184,N_39619);
xnor U43892 (N_43892,N_39222,N_39826);
or U43893 (N_43893,N_36807,N_38123);
nor U43894 (N_43894,N_39540,N_36181);
nand U43895 (N_43895,N_35846,N_36253);
xnor U43896 (N_43896,N_38059,N_39032);
and U43897 (N_43897,N_36764,N_37031);
nand U43898 (N_43898,N_37183,N_35901);
and U43899 (N_43899,N_35124,N_35194);
or U43900 (N_43900,N_38569,N_37341);
or U43901 (N_43901,N_37571,N_38351);
xnor U43902 (N_43902,N_36209,N_36330);
and U43903 (N_43903,N_38029,N_38470);
or U43904 (N_43904,N_38120,N_35563);
and U43905 (N_43905,N_38967,N_36768);
or U43906 (N_43906,N_38877,N_38244);
and U43907 (N_43907,N_38564,N_36182);
and U43908 (N_43908,N_38394,N_37263);
and U43909 (N_43909,N_36536,N_36103);
nand U43910 (N_43910,N_39820,N_38225);
nor U43911 (N_43911,N_36598,N_36189);
nand U43912 (N_43912,N_38184,N_39199);
nor U43913 (N_43913,N_37706,N_36162);
or U43914 (N_43914,N_37512,N_39035);
nand U43915 (N_43915,N_39767,N_38739);
xnor U43916 (N_43916,N_35330,N_38917);
and U43917 (N_43917,N_36310,N_39308);
nand U43918 (N_43918,N_36139,N_39492);
and U43919 (N_43919,N_39967,N_35767);
xor U43920 (N_43920,N_37842,N_39712);
nor U43921 (N_43921,N_35383,N_36581);
xnor U43922 (N_43922,N_36258,N_39258);
and U43923 (N_43923,N_35387,N_38325);
nand U43924 (N_43924,N_35629,N_39352);
and U43925 (N_43925,N_36428,N_37774);
nand U43926 (N_43926,N_39289,N_35673);
nand U43927 (N_43927,N_35951,N_39556);
xor U43928 (N_43928,N_35310,N_37921);
and U43929 (N_43929,N_38730,N_39846);
nor U43930 (N_43930,N_37176,N_36902);
and U43931 (N_43931,N_39609,N_39912);
or U43932 (N_43932,N_39828,N_37742);
and U43933 (N_43933,N_38094,N_35929);
nor U43934 (N_43934,N_39399,N_39016);
or U43935 (N_43935,N_38995,N_37299);
and U43936 (N_43936,N_36949,N_37045);
or U43937 (N_43937,N_39926,N_38755);
nand U43938 (N_43938,N_39220,N_37451);
nor U43939 (N_43939,N_39362,N_39095);
nor U43940 (N_43940,N_37168,N_37934);
nand U43941 (N_43941,N_37436,N_36299);
or U43942 (N_43942,N_36542,N_36688);
or U43943 (N_43943,N_35644,N_36212);
xnor U43944 (N_43944,N_38631,N_38440);
and U43945 (N_43945,N_39269,N_39987);
or U43946 (N_43946,N_35133,N_39744);
xnor U43947 (N_43947,N_37589,N_39919);
or U43948 (N_43948,N_37934,N_37042);
and U43949 (N_43949,N_38717,N_35762);
nor U43950 (N_43950,N_39580,N_37201);
nor U43951 (N_43951,N_39345,N_39373);
nand U43952 (N_43952,N_35321,N_37602);
and U43953 (N_43953,N_36618,N_37506);
or U43954 (N_43954,N_39097,N_37301);
or U43955 (N_43955,N_35850,N_36389);
nand U43956 (N_43956,N_35721,N_36776);
nor U43957 (N_43957,N_35787,N_39035);
xor U43958 (N_43958,N_36404,N_39112);
xnor U43959 (N_43959,N_35694,N_35330);
and U43960 (N_43960,N_35184,N_38375);
xor U43961 (N_43961,N_37901,N_39570);
or U43962 (N_43962,N_39778,N_39654);
nand U43963 (N_43963,N_38584,N_36120);
xor U43964 (N_43964,N_39913,N_35846);
nor U43965 (N_43965,N_39724,N_36108);
nand U43966 (N_43966,N_38655,N_36146);
and U43967 (N_43967,N_37737,N_38236);
nor U43968 (N_43968,N_39129,N_38114);
nand U43969 (N_43969,N_39113,N_35989);
or U43970 (N_43970,N_39670,N_39212);
and U43971 (N_43971,N_38128,N_38684);
nand U43972 (N_43972,N_38902,N_36328);
nor U43973 (N_43973,N_36690,N_38181);
and U43974 (N_43974,N_38483,N_39542);
xor U43975 (N_43975,N_35105,N_37326);
xor U43976 (N_43976,N_37953,N_35332);
and U43977 (N_43977,N_39481,N_35584);
or U43978 (N_43978,N_38595,N_39483);
or U43979 (N_43979,N_36664,N_36082);
nor U43980 (N_43980,N_38446,N_39309);
or U43981 (N_43981,N_37142,N_36585);
xor U43982 (N_43982,N_39317,N_36971);
nor U43983 (N_43983,N_39129,N_35254);
or U43984 (N_43984,N_35371,N_37208);
and U43985 (N_43985,N_35823,N_39401);
and U43986 (N_43986,N_35374,N_36547);
and U43987 (N_43987,N_39166,N_36980);
nor U43988 (N_43988,N_37679,N_37786);
or U43989 (N_43989,N_35230,N_38225);
xor U43990 (N_43990,N_36655,N_38819);
nand U43991 (N_43991,N_38702,N_39414);
and U43992 (N_43992,N_39625,N_35602);
and U43993 (N_43993,N_35396,N_39496);
nand U43994 (N_43994,N_35963,N_35135);
nor U43995 (N_43995,N_37126,N_38233);
nor U43996 (N_43996,N_38814,N_36681);
and U43997 (N_43997,N_38502,N_38239);
nor U43998 (N_43998,N_36339,N_38392);
xnor U43999 (N_43999,N_39998,N_39625);
nand U44000 (N_44000,N_36819,N_35792);
nor U44001 (N_44001,N_37487,N_36581);
nor U44002 (N_44002,N_38654,N_35075);
nand U44003 (N_44003,N_35872,N_37793);
nor U44004 (N_44004,N_38392,N_35835);
or U44005 (N_44005,N_38424,N_36597);
and U44006 (N_44006,N_37684,N_35819);
xor U44007 (N_44007,N_36142,N_38649);
nand U44008 (N_44008,N_37908,N_35537);
xnor U44009 (N_44009,N_38104,N_38440);
or U44010 (N_44010,N_39561,N_37110);
xor U44011 (N_44011,N_39958,N_38841);
and U44012 (N_44012,N_39375,N_37317);
or U44013 (N_44013,N_35705,N_38471);
or U44014 (N_44014,N_36288,N_39156);
nor U44015 (N_44015,N_37631,N_38229);
xor U44016 (N_44016,N_36090,N_38845);
or U44017 (N_44017,N_38107,N_37074);
xor U44018 (N_44018,N_36055,N_38005);
nand U44019 (N_44019,N_38225,N_36152);
nand U44020 (N_44020,N_36696,N_38639);
nand U44021 (N_44021,N_38252,N_37566);
xnor U44022 (N_44022,N_35310,N_35800);
and U44023 (N_44023,N_38217,N_39953);
nand U44024 (N_44024,N_39594,N_38846);
xor U44025 (N_44025,N_39268,N_36239);
xor U44026 (N_44026,N_36644,N_36684);
and U44027 (N_44027,N_38296,N_36449);
and U44028 (N_44028,N_36914,N_37317);
or U44029 (N_44029,N_36461,N_38509);
or U44030 (N_44030,N_38746,N_38030);
and U44031 (N_44031,N_35404,N_35288);
xnor U44032 (N_44032,N_39107,N_35499);
nor U44033 (N_44033,N_37456,N_35970);
nand U44034 (N_44034,N_38361,N_35292);
nand U44035 (N_44035,N_39491,N_38890);
nand U44036 (N_44036,N_35555,N_35381);
xnor U44037 (N_44037,N_38914,N_38464);
nand U44038 (N_44038,N_35978,N_38389);
nand U44039 (N_44039,N_35186,N_35504);
and U44040 (N_44040,N_37105,N_39032);
nand U44041 (N_44041,N_37519,N_39879);
and U44042 (N_44042,N_35125,N_36655);
or U44043 (N_44043,N_35957,N_36857);
nand U44044 (N_44044,N_38496,N_36579);
nor U44045 (N_44045,N_35927,N_38575);
nand U44046 (N_44046,N_36171,N_36865);
nor U44047 (N_44047,N_36651,N_35916);
xnor U44048 (N_44048,N_36509,N_36627);
or U44049 (N_44049,N_35225,N_36654);
and U44050 (N_44050,N_38188,N_39776);
xor U44051 (N_44051,N_35190,N_35222);
and U44052 (N_44052,N_39702,N_39536);
or U44053 (N_44053,N_36566,N_37096);
and U44054 (N_44054,N_38159,N_37571);
nor U44055 (N_44055,N_36225,N_39528);
and U44056 (N_44056,N_39826,N_38991);
nor U44057 (N_44057,N_39889,N_36490);
xnor U44058 (N_44058,N_37055,N_38904);
nor U44059 (N_44059,N_39161,N_38616);
or U44060 (N_44060,N_39609,N_36494);
nor U44061 (N_44061,N_38504,N_37822);
xor U44062 (N_44062,N_39634,N_37279);
nor U44063 (N_44063,N_39160,N_39398);
or U44064 (N_44064,N_38573,N_38447);
nand U44065 (N_44065,N_38133,N_36029);
nand U44066 (N_44066,N_35957,N_36234);
or U44067 (N_44067,N_37644,N_39232);
xor U44068 (N_44068,N_36082,N_39364);
nor U44069 (N_44069,N_35681,N_37149);
or U44070 (N_44070,N_37737,N_39167);
or U44071 (N_44071,N_38266,N_39711);
nor U44072 (N_44072,N_37900,N_38622);
and U44073 (N_44073,N_39556,N_37867);
nor U44074 (N_44074,N_37840,N_36569);
and U44075 (N_44075,N_39009,N_38124);
nand U44076 (N_44076,N_39998,N_37948);
nand U44077 (N_44077,N_38311,N_37710);
xor U44078 (N_44078,N_39952,N_38810);
nor U44079 (N_44079,N_39101,N_39566);
nor U44080 (N_44080,N_39582,N_35816);
xnor U44081 (N_44081,N_37852,N_39807);
nand U44082 (N_44082,N_38165,N_39120);
nand U44083 (N_44083,N_37028,N_37195);
xor U44084 (N_44084,N_38198,N_36621);
nor U44085 (N_44085,N_38618,N_37893);
xnor U44086 (N_44086,N_35050,N_38092);
nor U44087 (N_44087,N_39337,N_37025);
nor U44088 (N_44088,N_38955,N_37834);
nand U44089 (N_44089,N_36557,N_36696);
and U44090 (N_44090,N_35813,N_35894);
xnor U44091 (N_44091,N_37154,N_37885);
and U44092 (N_44092,N_39796,N_38927);
nand U44093 (N_44093,N_39009,N_37176);
nand U44094 (N_44094,N_36965,N_38254);
nor U44095 (N_44095,N_38717,N_35549);
and U44096 (N_44096,N_38982,N_35691);
nand U44097 (N_44097,N_35785,N_39385);
and U44098 (N_44098,N_37499,N_36746);
nand U44099 (N_44099,N_38621,N_38829);
or U44100 (N_44100,N_36110,N_37842);
xnor U44101 (N_44101,N_35975,N_36573);
nand U44102 (N_44102,N_39721,N_37366);
nor U44103 (N_44103,N_37518,N_35262);
nor U44104 (N_44104,N_39184,N_38998);
nand U44105 (N_44105,N_36450,N_36006);
or U44106 (N_44106,N_39755,N_35064);
nor U44107 (N_44107,N_39334,N_37751);
and U44108 (N_44108,N_36507,N_38955);
or U44109 (N_44109,N_39355,N_38164);
or U44110 (N_44110,N_38740,N_37800);
nor U44111 (N_44111,N_38111,N_37515);
nor U44112 (N_44112,N_37300,N_35298);
xor U44113 (N_44113,N_39918,N_38555);
xnor U44114 (N_44114,N_39897,N_36831);
or U44115 (N_44115,N_35745,N_36148);
nor U44116 (N_44116,N_38006,N_37716);
xor U44117 (N_44117,N_36028,N_38443);
or U44118 (N_44118,N_39954,N_36297);
nor U44119 (N_44119,N_37156,N_38738);
nor U44120 (N_44120,N_36200,N_36799);
or U44121 (N_44121,N_36486,N_36883);
or U44122 (N_44122,N_36533,N_37573);
nand U44123 (N_44123,N_36896,N_36237);
and U44124 (N_44124,N_37828,N_38133);
nor U44125 (N_44125,N_37804,N_35521);
or U44126 (N_44126,N_37560,N_37964);
nand U44127 (N_44127,N_35253,N_35458);
xor U44128 (N_44128,N_37298,N_35333);
and U44129 (N_44129,N_39794,N_36699);
and U44130 (N_44130,N_36758,N_37803);
and U44131 (N_44131,N_35677,N_39721);
or U44132 (N_44132,N_36689,N_35619);
or U44133 (N_44133,N_36714,N_37604);
or U44134 (N_44134,N_38155,N_39044);
xor U44135 (N_44135,N_38977,N_38880);
nor U44136 (N_44136,N_36848,N_38506);
and U44137 (N_44137,N_35910,N_39819);
and U44138 (N_44138,N_38358,N_35930);
nand U44139 (N_44139,N_35446,N_38286);
xnor U44140 (N_44140,N_37042,N_39312);
or U44141 (N_44141,N_37303,N_36882);
xor U44142 (N_44142,N_39423,N_39633);
xor U44143 (N_44143,N_36424,N_37052);
and U44144 (N_44144,N_37542,N_38347);
or U44145 (N_44145,N_37887,N_36799);
and U44146 (N_44146,N_39582,N_37521);
nand U44147 (N_44147,N_36843,N_38742);
xnor U44148 (N_44148,N_39037,N_37247);
nor U44149 (N_44149,N_39942,N_36554);
and U44150 (N_44150,N_38393,N_36540);
xor U44151 (N_44151,N_36190,N_35581);
nand U44152 (N_44152,N_37256,N_36292);
or U44153 (N_44153,N_35471,N_39857);
and U44154 (N_44154,N_38993,N_36714);
and U44155 (N_44155,N_38242,N_38459);
xor U44156 (N_44156,N_39744,N_35194);
and U44157 (N_44157,N_35350,N_37954);
nor U44158 (N_44158,N_39006,N_38404);
and U44159 (N_44159,N_39641,N_39528);
and U44160 (N_44160,N_38444,N_35771);
nand U44161 (N_44161,N_36543,N_37858);
or U44162 (N_44162,N_36593,N_36377);
or U44163 (N_44163,N_37214,N_38899);
nor U44164 (N_44164,N_38199,N_35675);
nand U44165 (N_44165,N_35119,N_38925);
or U44166 (N_44166,N_35379,N_37481);
or U44167 (N_44167,N_36799,N_39936);
or U44168 (N_44168,N_36942,N_37015);
and U44169 (N_44169,N_35558,N_36602);
nand U44170 (N_44170,N_35597,N_38876);
xor U44171 (N_44171,N_38301,N_36552);
nor U44172 (N_44172,N_38148,N_35140);
or U44173 (N_44173,N_38695,N_39657);
nor U44174 (N_44174,N_36084,N_36173);
and U44175 (N_44175,N_37734,N_38552);
xor U44176 (N_44176,N_38872,N_36154);
nor U44177 (N_44177,N_35136,N_39539);
and U44178 (N_44178,N_35540,N_38476);
nor U44179 (N_44179,N_38954,N_39527);
xnor U44180 (N_44180,N_37112,N_39026);
and U44181 (N_44181,N_39463,N_39930);
or U44182 (N_44182,N_38908,N_35340);
or U44183 (N_44183,N_38363,N_37643);
nor U44184 (N_44184,N_38301,N_36415);
xor U44185 (N_44185,N_39874,N_38203);
xnor U44186 (N_44186,N_35560,N_36825);
and U44187 (N_44187,N_37864,N_38007);
or U44188 (N_44188,N_37907,N_36469);
and U44189 (N_44189,N_36923,N_37048);
xnor U44190 (N_44190,N_36915,N_38008);
and U44191 (N_44191,N_39347,N_37702);
xnor U44192 (N_44192,N_38057,N_35698);
and U44193 (N_44193,N_38033,N_38267);
nor U44194 (N_44194,N_38443,N_39404);
nand U44195 (N_44195,N_39586,N_37293);
and U44196 (N_44196,N_36184,N_38142);
and U44197 (N_44197,N_35902,N_38617);
and U44198 (N_44198,N_36555,N_37516);
or U44199 (N_44199,N_37096,N_37463);
xnor U44200 (N_44200,N_36105,N_35431);
nand U44201 (N_44201,N_35921,N_35819);
xnor U44202 (N_44202,N_35831,N_39352);
nor U44203 (N_44203,N_38564,N_36826);
nor U44204 (N_44204,N_37960,N_36797);
and U44205 (N_44205,N_37182,N_38094);
nor U44206 (N_44206,N_36356,N_38745);
and U44207 (N_44207,N_35389,N_35354);
and U44208 (N_44208,N_39999,N_35846);
or U44209 (N_44209,N_35116,N_38324);
and U44210 (N_44210,N_37874,N_35107);
and U44211 (N_44211,N_36392,N_36113);
nor U44212 (N_44212,N_38750,N_39790);
nor U44213 (N_44213,N_36911,N_36427);
or U44214 (N_44214,N_38334,N_37303);
and U44215 (N_44215,N_38831,N_36290);
nand U44216 (N_44216,N_38603,N_38307);
or U44217 (N_44217,N_35900,N_37476);
xor U44218 (N_44218,N_38120,N_36794);
nand U44219 (N_44219,N_37653,N_36369);
and U44220 (N_44220,N_38352,N_35235);
nor U44221 (N_44221,N_35154,N_39719);
xnor U44222 (N_44222,N_39698,N_37893);
nand U44223 (N_44223,N_37886,N_36251);
xnor U44224 (N_44224,N_39354,N_38990);
xnor U44225 (N_44225,N_35699,N_38951);
and U44226 (N_44226,N_39806,N_37969);
or U44227 (N_44227,N_38089,N_37479);
xnor U44228 (N_44228,N_36349,N_39661);
nand U44229 (N_44229,N_38568,N_39247);
nand U44230 (N_44230,N_36639,N_38510);
nor U44231 (N_44231,N_37171,N_37361);
xnor U44232 (N_44232,N_39053,N_37396);
nand U44233 (N_44233,N_37325,N_36474);
nand U44234 (N_44234,N_35696,N_36410);
and U44235 (N_44235,N_38787,N_39776);
or U44236 (N_44236,N_35974,N_35380);
nand U44237 (N_44237,N_39826,N_35994);
or U44238 (N_44238,N_38872,N_37570);
or U44239 (N_44239,N_37656,N_38549);
and U44240 (N_44240,N_39372,N_38079);
and U44241 (N_44241,N_36040,N_36468);
or U44242 (N_44242,N_36380,N_35308);
and U44243 (N_44243,N_37052,N_35201);
and U44244 (N_44244,N_37938,N_39176);
or U44245 (N_44245,N_37770,N_39546);
xor U44246 (N_44246,N_35432,N_36008);
nor U44247 (N_44247,N_36803,N_39424);
and U44248 (N_44248,N_37220,N_39313);
nand U44249 (N_44249,N_35131,N_36431);
and U44250 (N_44250,N_35869,N_37367);
xnor U44251 (N_44251,N_38738,N_35935);
nand U44252 (N_44252,N_39824,N_35370);
or U44253 (N_44253,N_39973,N_36837);
nand U44254 (N_44254,N_38376,N_38642);
nand U44255 (N_44255,N_37049,N_39225);
nand U44256 (N_44256,N_36015,N_37677);
xor U44257 (N_44257,N_37321,N_38703);
nor U44258 (N_44258,N_38589,N_38163);
nor U44259 (N_44259,N_35154,N_36890);
nand U44260 (N_44260,N_35354,N_36847);
nor U44261 (N_44261,N_39949,N_38953);
and U44262 (N_44262,N_36815,N_36995);
and U44263 (N_44263,N_37939,N_38601);
xnor U44264 (N_44264,N_39705,N_36781);
and U44265 (N_44265,N_37235,N_39822);
and U44266 (N_44266,N_38916,N_39887);
and U44267 (N_44267,N_39032,N_35806);
nor U44268 (N_44268,N_35905,N_38236);
xnor U44269 (N_44269,N_36399,N_37231);
or U44270 (N_44270,N_36968,N_38998);
nand U44271 (N_44271,N_35767,N_35028);
and U44272 (N_44272,N_36714,N_36164);
xnor U44273 (N_44273,N_38983,N_35852);
and U44274 (N_44274,N_38613,N_35165);
nor U44275 (N_44275,N_35381,N_36554);
nand U44276 (N_44276,N_37316,N_38439);
nand U44277 (N_44277,N_37865,N_36917);
or U44278 (N_44278,N_36561,N_38785);
and U44279 (N_44279,N_39851,N_36159);
or U44280 (N_44280,N_38641,N_38888);
nor U44281 (N_44281,N_36769,N_36265);
nor U44282 (N_44282,N_38481,N_37160);
and U44283 (N_44283,N_38286,N_38102);
nor U44284 (N_44284,N_35692,N_35230);
and U44285 (N_44285,N_38393,N_37925);
xor U44286 (N_44286,N_35190,N_36857);
nand U44287 (N_44287,N_36865,N_35174);
nand U44288 (N_44288,N_37174,N_38923);
and U44289 (N_44289,N_36257,N_38897);
xnor U44290 (N_44290,N_39012,N_35919);
nor U44291 (N_44291,N_35180,N_37713);
nand U44292 (N_44292,N_38815,N_39272);
nor U44293 (N_44293,N_39325,N_36197);
nand U44294 (N_44294,N_38012,N_39748);
nor U44295 (N_44295,N_39742,N_37068);
nor U44296 (N_44296,N_38777,N_39969);
or U44297 (N_44297,N_38166,N_37796);
xnor U44298 (N_44298,N_39095,N_35227);
and U44299 (N_44299,N_35389,N_35880);
nand U44300 (N_44300,N_36314,N_36715);
and U44301 (N_44301,N_36477,N_38388);
xor U44302 (N_44302,N_39905,N_38973);
and U44303 (N_44303,N_38238,N_36902);
nor U44304 (N_44304,N_39497,N_35074);
nor U44305 (N_44305,N_37999,N_39633);
and U44306 (N_44306,N_36765,N_35221);
xor U44307 (N_44307,N_35372,N_35221);
nand U44308 (N_44308,N_37988,N_39623);
xnor U44309 (N_44309,N_37439,N_37771);
nand U44310 (N_44310,N_37586,N_38842);
nand U44311 (N_44311,N_39648,N_39345);
xor U44312 (N_44312,N_36489,N_38805);
and U44313 (N_44313,N_39598,N_38036);
nor U44314 (N_44314,N_35732,N_39188);
and U44315 (N_44315,N_35616,N_37112);
nor U44316 (N_44316,N_35939,N_38166);
and U44317 (N_44317,N_39861,N_37014);
xor U44318 (N_44318,N_37652,N_38288);
xor U44319 (N_44319,N_35074,N_38282);
nand U44320 (N_44320,N_36304,N_37456);
and U44321 (N_44321,N_37026,N_38066);
xnor U44322 (N_44322,N_36819,N_36045);
and U44323 (N_44323,N_35819,N_39687);
or U44324 (N_44324,N_36623,N_38059);
nor U44325 (N_44325,N_35597,N_37463);
or U44326 (N_44326,N_39744,N_38351);
xnor U44327 (N_44327,N_36167,N_37563);
or U44328 (N_44328,N_38624,N_37032);
nor U44329 (N_44329,N_36776,N_39034);
nand U44330 (N_44330,N_36173,N_36652);
nor U44331 (N_44331,N_39354,N_38305);
xnor U44332 (N_44332,N_38334,N_39703);
xor U44333 (N_44333,N_37942,N_37486);
and U44334 (N_44334,N_38574,N_38268);
and U44335 (N_44335,N_37275,N_37926);
or U44336 (N_44336,N_37893,N_38944);
and U44337 (N_44337,N_37442,N_37563);
or U44338 (N_44338,N_38804,N_35500);
xnor U44339 (N_44339,N_39527,N_37440);
xnor U44340 (N_44340,N_38971,N_37860);
nor U44341 (N_44341,N_38951,N_37119);
nand U44342 (N_44342,N_37876,N_37254);
nand U44343 (N_44343,N_38371,N_38383);
nor U44344 (N_44344,N_38391,N_35452);
xor U44345 (N_44345,N_37586,N_35518);
nor U44346 (N_44346,N_37266,N_35117);
nand U44347 (N_44347,N_39724,N_37159);
or U44348 (N_44348,N_37820,N_36102);
and U44349 (N_44349,N_39016,N_37126);
nor U44350 (N_44350,N_35637,N_36483);
or U44351 (N_44351,N_38046,N_35743);
nand U44352 (N_44352,N_39277,N_35966);
xnor U44353 (N_44353,N_38610,N_37564);
xnor U44354 (N_44354,N_38875,N_37357);
nand U44355 (N_44355,N_38536,N_35053);
nor U44356 (N_44356,N_39059,N_36870);
and U44357 (N_44357,N_38999,N_35907);
and U44358 (N_44358,N_38087,N_39140);
and U44359 (N_44359,N_35809,N_38026);
or U44360 (N_44360,N_38717,N_37409);
or U44361 (N_44361,N_37476,N_35280);
nand U44362 (N_44362,N_35006,N_35013);
and U44363 (N_44363,N_38583,N_36478);
nand U44364 (N_44364,N_36371,N_36238);
nor U44365 (N_44365,N_38901,N_36275);
and U44366 (N_44366,N_35761,N_37428);
or U44367 (N_44367,N_35333,N_39235);
nand U44368 (N_44368,N_38674,N_39525);
and U44369 (N_44369,N_36914,N_36067);
nor U44370 (N_44370,N_37035,N_39358);
nor U44371 (N_44371,N_36668,N_36206);
nor U44372 (N_44372,N_38893,N_39597);
xor U44373 (N_44373,N_39800,N_37407);
nor U44374 (N_44374,N_36666,N_36042);
or U44375 (N_44375,N_37891,N_36795);
or U44376 (N_44376,N_35067,N_36393);
nor U44377 (N_44377,N_37915,N_39548);
xnor U44378 (N_44378,N_37882,N_37570);
xnor U44379 (N_44379,N_39286,N_36587);
nand U44380 (N_44380,N_35317,N_36891);
xor U44381 (N_44381,N_38055,N_35740);
or U44382 (N_44382,N_39469,N_38668);
nor U44383 (N_44383,N_35879,N_35417);
nand U44384 (N_44384,N_36564,N_39890);
nor U44385 (N_44385,N_35579,N_38749);
or U44386 (N_44386,N_36179,N_38516);
nand U44387 (N_44387,N_39898,N_35700);
nand U44388 (N_44388,N_38275,N_39735);
and U44389 (N_44389,N_39022,N_39773);
nand U44390 (N_44390,N_37977,N_36923);
xor U44391 (N_44391,N_39894,N_38406);
or U44392 (N_44392,N_37292,N_36165);
nand U44393 (N_44393,N_36719,N_39995);
xnor U44394 (N_44394,N_36817,N_36667);
and U44395 (N_44395,N_38381,N_37627);
xor U44396 (N_44396,N_39021,N_36902);
nand U44397 (N_44397,N_35504,N_37933);
or U44398 (N_44398,N_35622,N_38086);
nand U44399 (N_44399,N_37102,N_36376);
or U44400 (N_44400,N_39005,N_36086);
nor U44401 (N_44401,N_39679,N_39650);
xnor U44402 (N_44402,N_36355,N_37558);
xor U44403 (N_44403,N_38336,N_39778);
and U44404 (N_44404,N_37734,N_37702);
or U44405 (N_44405,N_35333,N_39105);
nor U44406 (N_44406,N_38143,N_39208);
xnor U44407 (N_44407,N_35496,N_37249);
and U44408 (N_44408,N_35608,N_36424);
xnor U44409 (N_44409,N_36695,N_37659);
nor U44410 (N_44410,N_36305,N_39353);
xor U44411 (N_44411,N_35663,N_35606);
or U44412 (N_44412,N_36231,N_35378);
nand U44413 (N_44413,N_36989,N_36013);
nor U44414 (N_44414,N_37175,N_39079);
or U44415 (N_44415,N_37664,N_39523);
and U44416 (N_44416,N_38795,N_35419);
nor U44417 (N_44417,N_36039,N_37978);
nor U44418 (N_44418,N_35322,N_37345);
and U44419 (N_44419,N_36781,N_38705);
xnor U44420 (N_44420,N_36410,N_37338);
and U44421 (N_44421,N_39585,N_38911);
nand U44422 (N_44422,N_38390,N_38856);
nor U44423 (N_44423,N_36206,N_38952);
xor U44424 (N_44424,N_37810,N_36100);
nand U44425 (N_44425,N_36879,N_36780);
xor U44426 (N_44426,N_35298,N_37551);
nand U44427 (N_44427,N_38603,N_36659);
and U44428 (N_44428,N_36345,N_38606);
and U44429 (N_44429,N_36612,N_36457);
xnor U44430 (N_44430,N_38308,N_39276);
xnor U44431 (N_44431,N_39947,N_39250);
and U44432 (N_44432,N_35625,N_37924);
xor U44433 (N_44433,N_35354,N_35152);
nand U44434 (N_44434,N_37333,N_35790);
nand U44435 (N_44435,N_36333,N_36994);
xnor U44436 (N_44436,N_36118,N_37027);
xnor U44437 (N_44437,N_35185,N_36782);
or U44438 (N_44438,N_39873,N_38993);
or U44439 (N_44439,N_37069,N_38310);
nor U44440 (N_44440,N_37620,N_39510);
nand U44441 (N_44441,N_35038,N_36367);
and U44442 (N_44442,N_36606,N_36414);
xor U44443 (N_44443,N_35217,N_38648);
or U44444 (N_44444,N_37523,N_37710);
xor U44445 (N_44445,N_36763,N_37533);
and U44446 (N_44446,N_37109,N_35470);
or U44447 (N_44447,N_37651,N_37858);
nor U44448 (N_44448,N_38572,N_38174);
or U44449 (N_44449,N_35507,N_38615);
nor U44450 (N_44450,N_36879,N_36068);
nor U44451 (N_44451,N_37634,N_38672);
or U44452 (N_44452,N_36452,N_39026);
or U44453 (N_44453,N_37768,N_36170);
and U44454 (N_44454,N_38901,N_37336);
or U44455 (N_44455,N_35542,N_38424);
and U44456 (N_44456,N_38908,N_37614);
and U44457 (N_44457,N_36739,N_39790);
nor U44458 (N_44458,N_37334,N_38763);
nand U44459 (N_44459,N_37625,N_37295);
nand U44460 (N_44460,N_36358,N_39713);
xor U44461 (N_44461,N_39598,N_35251);
nand U44462 (N_44462,N_39245,N_35851);
nand U44463 (N_44463,N_36025,N_35651);
nor U44464 (N_44464,N_37509,N_37131);
nor U44465 (N_44465,N_37632,N_35700);
nor U44466 (N_44466,N_38693,N_36409);
nor U44467 (N_44467,N_36167,N_35132);
nand U44468 (N_44468,N_37666,N_35316);
or U44469 (N_44469,N_35353,N_37763);
xor U44470 (N_44470,N_38966,N_36079);
nor U44471 (N_44471,N_38212,N_36694);
nor U44472 (N_44472,N_38663,N_36993);
and U44473 (N_44473,N_37309,N_37332);
xor U44474 (N_44474,N_37096,N_35811);
and U44475 (N_44475,N_37066,N_38946);
nand U44476 (N_44476,N_35376,N_38900);
nand U44477 (N_44477,N_35256,N_36558);
xor U44478 (N_44478,N_36219,N_38383);
or U44479 (N_44479,N_37685,N_36173);
nor U44480 (N_44480,N_39462,N_35613);
nor U44481 (N_44481,N_37871,N_38517);
nor U44482 (N_44482,N_36686,N_36142);
nor U44483 (N_44483,N_35546,N_35052);
nand U44484 (N_44484,N_35783,N_35301);
or U44485 (N_44485,N_38395,N_36501);
nand U44486 (N_44486,N_35009,N_38789);
nor U44487 (N_44487,N_36311,N_37442);
xnor U44488 (N_44488,N_35354,N_35396);
nand U44489 (N_44489,N_36314,N_36703);
and U44490 (N_44490,N_38073,N_35817);
nor U44491 (N_44491,N_35538,N_37804);
nor U44492 (N_44492,N_38697,N_36588);
nor U44493 (N_44493,N_37023,N_39724);
and U44494 (N_44494,N_39580,N_37715);
and U44495 (N_44495,N_39997,N_37615);
or U44496 (N_44496,N_36603,N_39810);
and U44497 (N_44497,N_37666,N_38875);
nand U44498 (N_44498,N_35237,N_37439);
nand U44499 (N_44499,N_35787,N_36148);
and U44500 (N_44500,N_39269,N_35916);
or U44501 (N_44501,N_36915,N_37949);
nor U44502 (N_44502,N_39878,N_36735);
nor U44503 (N_44503,N_35575,N_38858);
nand U44504 (N_44504,N_39364,N_38166);
and U44505 (N_44505,N_36097,N_37341);
nand U44506 (N_44506,N_39273,N_35292);
xor U44507 (N_44507,N_36049,N_35090);
xor U44508 (N_44508,N_35898,N_36722);
nor U44509 (N_44509,N_38503,N_38714);
or U44510 (N_44510,N_39380,N_39858);
nor U44511 (N_44511,N_37544,N_38016);
and U44512 (N_44512,N_37734,N_38255);
nor U44513 (N_44513,N_36576,N_36228);
nor U44514 (N_44514,N_38188,N_38042);
and U44515 (N_44515,N_38906,N_39330);
xor U44516 (N_44516,N_35668,N_39745);
nor U44517 (N_44517,N_39446,N_37409);
nand U44518 (N_44518,N_35736,N_36431);
xnor U44519 (N_44519,N_38972,N_35419);
nand U44520 (N_44520,N_36874,N_39983);
nand U44521 (N_44521,N_39595,N_36504);
nand U44522 (N_44522,N_38837,N_37825);
nand U44523 (N_44523,N_37082,N_37582);
nand U44524 (N_44524,N_36466,N_37230);
or U44525 (N_44525,N_39675,N_36986);
nor U44526 (N_44526,N_39548,N_37854);
and U44527 (N_44527,N_36947,N_36530);
nand U44528 (N_44528,N_36335,N_37157);
nor U44529 (N_44529,N_35359,N_36554);
xnor U44530 (N_44530,N_35326,N_37373);
nand U44531 (N_44531,N_36557,N_39373);
nor U44532 (N_44532,N_37339,N_35497);
and U44533 (N_44533,N_37189,N_37488);
and U44534 (N_44534,N_38946,N_36526);
and U44535 (N_44535,N_36746,N_36050);
nand U44536 (N_44536,N_39110,N_36086);
nor U44537 (N_44537,N_36998,N_36547);
nand U44538 (N_44538,N_38036,N_36990);
or U44539 (N_44539,N_37387,N_39309);
and U44540 (N_44540,N_37961,N_37184);
and U44541 (N_44541,N_38531,N_35965);
and U44542 (N_44542,N_39310,N_38151);
nand U44543 (N_44543,N_38317,N_38148);
xnor U44544 (N_44544,N_37073,N_39257);
xnor U44545 (N_44545,N_36884,N_36763);
nor U44546 (N_44546,N_37288,N_36098);
xnor U44547 (N_44547,N_38473,N_37275);
or U44548 (N_44548,N_39778,N_36506);
nand U44549 (N_44549,N_38140,N_39760);
nand U44550 (N_44550,N_38719,N_39664);
nor U44551 (N_44551,N_37394,N_38720);
and U44552 (N_44552,N_38880,N_37194);
nor U44553 (N_44553,N_35697,N_37229);
nor U44554 (N_44554,N_36437,N_37038);
and U44555 (N_44555,N_38947,N_35607);
xnor U44556 (N_44556,N_39852,N_36181);
or U44557 (N_44557,N_39556,N_38660);
or U44558 (N_44558,N_38174,N_39571);
xnor U44559 (N_44559,N_37167,N_38879);
xnor U44560 (N_44560,N_39650,N_35296);
nand U44561 (N_44561,N_35727,N_39602);
and U44562 (N_44562,N_37874,N_38780);
nand U44563 (N_44563,N_37108,N_38995);
nor U44564 (N_44564,N_36536,N_37975);
or U44565 (N_44565,N_37488,N_35562);
nor U44566 (N_44566,N_35652,N_37467);
and U44567 (N_44567,N_39788,N_37170);
and U44568 (N_44568,N_38108,N_38034);
nand U44569 (N_44569,N_39462,N_36938);
nand U44570 (N_44570,N_36753,N_35339);
and U44571 (N_44571,N_35724,N_39710);
xnor U44572 (N_44572,N_37527,N_35555);
or U44573 (N_44573,N_36328,N_38798);
xor U44574 (N_44574,N_39810,N_38116);
nand U44575 (N_44575,N_35748,N_35379);
xor U44576 (N_44576,N_36131,N_39761);
xor U44577 (N_44577,N_39126,N_38163);
and U44578 (N_44578,N_35308,N_38211);
or U44579 (N_44579,N_36036,N_38187);
nand U44580 (N_44580,N_39803,N_35353);
xnor U44581 (N_44581,N_35467,N_37922);
or U44582 (N_44582,N_37112,N_36898);
nor U44583 (N_44583,N_36255,N_37181);
or U44584 (N_44584,N_37774,N_37691);
xor U44585 (N_44585,N_35644,N_38898);
nor U44586 (N_44586,N_39547,N_39049);
nor U44587 (N_44587,N_37846,N_37030);
and U44588 (N_44588,N_36372,N_39079);
or U44589 (N_44589,N_38890,N_36205);
nand U44590 (N_44590,N_36169,N_35980);
nand U44591 (N_44591,N_39251,N_37645);
xnor U44592 (N_44592,N_35312,N_39791);
or U44593 (N_44593,N_35170,N_36818);
or U44594 (N_44594,N_37537,N_36755);
nand U44595 (N_44595,N_39403,N_38884);
xor U44596 (N_44596,N_37299,N_36973);
nand U44597 (N_44597,N_36342,N_39324);
nand U44598 (N_44598,N_35737,N_36544);
and U44599 (N_44599,N_39371,N_39357);
nor U44600 (N_44600,N_39144,N_35213);
nand U44601 (N_44601,N_39615,N_35368);
nand U44602 (N_44602,N_39814,N_35558);
or U44603 (N_44603,N_35672,N_38514);
xnor U44604 (N_44604,N_39326,N_37183);
nand U44605 (N_44605,N_39732,N_38702);
xnor U44606 (N_44606,N_35925,N_36776);
or U44607 (N_44607,N_35543,N_36043);
nand U44608 (N_44608,N_36043,N_38590);
xor U44609 (N_44609,N_36524,N_37325);
nor U44610 (N_44610,N_38710,N_38126);
xor U44611 (N_44611,N_36868,N_37637);
nor U44612 (N_44612,N_37625,N_35909);
nor U44613 (N_44613,N_39628,N_36692);
nand U44614 (N_44614,N_38068,N_35017);
or U44615 (N_44615,N_39613,N_39604);
nor U44616 (N_44616,N_37411,N_38198);
and U44617 (N_44617,N_36815,N_37282);
xnor U44618 (N_44618,N_37381,N_35596);
and U44619 (N_44619,N_38464,N_39653);
and U44620 (N_44620,N_39977,N_36472);
nand U44621 (N_44621,N_35493,N_35029);
or U44622 (N_44622,N_39334,N_38707);
and U44623 (N_44623,N_36152,N_36526);
or U44624 (N_44624,N_36166,N_36485);
and U44625 (N_44625,N_39620,N_39924);
or U44626 (N_44626,N_37364,N_39347);
xnor U44627 (N_44627,N_39679,N_36704);
or U44628 (N_44628,N_35038,N_36317);
and U44629 (N_44629,N_38543,N_39434);
nor U44630 (N_44630,N_36027,N_35939);
and U44631 (N_44631,N_35412,N_37039);
or U44632 (N_44632,N_39721,N_39834);
nor U44633 (N_44633,N_37789,N_35332);
nand U44634 (N_44634,N_38599,N_36251);
or U44635 (N_44635,N_39516,N_39967);
nand U44636 (N_44636,N_39359,N_37478);
nand U44637 (N_44637,N_35773,N_38422);
nor U44638 (N_44638,N_39041,N_38124);
or U44639 (N_44639,N_37456,N_36865);
or U44640 (N_44640,N_37017,N_38886);
xnor U44641 (N_44641,N_38324,N_38344);
or U44642 (N_44642,N_37867,N_37649);
nand U44643 (N_44643,N_39204,N_36880);
or U44644 (N_44644,N_35435,N_39007);
or U44645 (N_44645,N_35373,N_38779);
nor U44646 (N_44646,N_35426,N_37452);
nor U44647 (N_44647,N_36213,N_39781);
nor U44648 (N_44648,N_38044,N_39191);
nor U44649 (N_44649,N_36631,N_38759);
and U44650 (N_44650,N_35176,N_38560);
and U44651 (N_44651,N_37950,N_36122);
nand U44652 (N_44652,N_38719,N_36069);
and U44653 (N_44653,N_39460,N_39061);
or U44654 (N_44654,N_37459,N_38762);
and U44655 (N_44655,N_35675,N_38559);
and U44656 (N_44656,N_39856,N_38966);
nor U44657 (N_44657,N_38814,N_38264);
or U44658 (N_44658,N_38927,N_36269);
xor U44659 (N_44659,N_36153,N_37528);
nor U44660 (N_44660,N_39809,N_39275);
nand U44661 (N_44661,N_35153,N_35119);
or U44662 (N_44662,N_39501,N_37159);
and U44663 (N_44663,N_36560,N_39058);
xnor U44664 (N_44664,N_36722,N_36931);
nor U44665 (N_44665,N_39478,N_35509);
or U44666 (N_44666,N_37106,N_36375);
nand U44667 (N_44667,N_37297,N_35937);
xnor U44668 (N_44668,N_37146,N_37592);
or U44669 (N_44669,N_36646,N_36303);
and U44670 (N_44670,N_37645,N_38314);
xor U44671 (N_44671,N_38843,N_38845);
nor U44672 (N_44672,N_38952,N_35221);
xnor U44673 (N_44673,N_36787,N_37554);
and U44674 (N_44674,N_39902,N_37351);
and U44675 (N_44675,N_39454,N_35088);
nor U44676 (N_44676,N_35507,N_38749);
xor U44677 (N_44677,N_38175,N_35278);
nand U44678 (N_44678,N_39511,N_38906);
nor U44679 (N_44679,N_39826,N_36764);
xnor U44680 (N_44680,N_35492,N_39350);
xnor U44681 (N_44681,N_39117,N_38498);
nand U44682 (N_44682,N_36561,N_36655);
nor U44683 (N_44683,N_37325,N_35115);
nor U44684 (N_44684,N_39399,N_35279);
nand U44685 (N_44685,N_35303,N_36052);
nor U44686 (N_44686,N_37100,N_36786);
xnor U44687 (N_44687,N_35571,N_38452);
xnor U44688 (N_44688,N_37856,N_37748);
nand U44689 (N_44689,N_36001,N_37261);
nand U44690 (N_44690,N_37419,N_37616);
xnor U44691 (N_44691,N_37932,N_38344);
xor U44692 (N_44692,N_36665,N_38447);
nor U44693 (N_44693,N_37089,N_35002);
nand U44694 (N_44694,N_37896,N_39985);
nor U44695 (N_44695,N_39076,N_35519);
or U44696 (N_44696,N_36361,N_37310);
nor U44697 (N_44697,N_38232,N_39794);
nor U44698 (N_44698,N_38863,N_36096);
or U44699 (N_44699,N_38411,N_39149);
or U44700 (N_44700,N_35064,N_38325);
xor U44701 (N_44701,N_37056,N_35922);
nor U44702 (N_44702,N_39675,N_35177);
nor U44703 (N_44703,N_37972,N_35000);
xor U44704 (N_44704,N_37155,N_36580);
nor U44705 (N_44705,N_37270,N_36155);
nor U44706 (N_44706,N_38892,N_37154);
xor U44707 (N_44707,N_39432,N_37645);
nor U44708 (N_44708,N_38983,N_38776);
or U44709 (N_44709,N_39142,N_38206);
xor U44710 (N_44710,N_38134,N_37002);
nor U44711 (N_44711,N_36042,N_35368);
nand U44712 (N_44712,N_37913,N_37283);
or U44713 (N_44713,N_37922,N_37002);
and U44714 (N_44714,N_37485,N_39066);
and U44715 (N_44715,N_35652,N_35465);
xor U44716 (N_44716,N_35398,N_38090);
nand U44717 (N_44717,N_35386,N_39309);
nand U44718 (N_44718,N_36692,N_36417);
nor U44719 (N_44719,N_36001,N_39152);
and U44720 (N_44720,N_38870,N_36917);
and U44721 (N_44721,N_36913,N_38529);
nor U44722 (N_44722,N_35200,N_36866);
xor U44723 (N_44723,N_35453,N_37417);
nor U44724 (N_44724,N_39240,N_38570);
xnor U44725 (N_44725,N_37113,N_38193);
xnor U44726 (N_44726,N_38962,N_35583);
xor U44727 (N_44727,N_35661,N_39370);
or U44728 (N_44728,N_35084,N_39000);
or U44729 (N_44729,N_37560,N_39940);
or U44730 (N_44730,N_38664,N_36134);
or U44731 (N_44731,N_39966,N_37651);
nand U44732 (N_44732,N_38142,N_37973);
nor U44733 (N_44733,N_38850,N_38439);
nor U44734 (N_44734,N_36009,N_38507);
and U44735 (N_44735,N_38384,N_36425);
or U44736 (N_44736,N_38452,N_38330);
xnor U44737 (N_44737,N_37374,N_36128);
nand U44738 (N_44738,N_37973,N_36839);
xnor U44739 (N_44739,N_37335,N_36980);
and U44740 (N_44740,N_36146,N_39854);
and U44741 (N_44741,N_37084,N_35546);
nand U44742 (N_44742,N_37917,N_39435);
nand U44743 (N_44743,N_37529,N_39918);
or U44744 (N_44744,N_39401,N_36895);
xnor U44745 (N_44745,N_39766,N_36733);
xnor U44746 (N_44746,N_39580,N_35272);
or U44747 (N_44747,N_37097,N_37256);
nor U44748 (N_44748,N_37700,N_37471);
nor U44749 (N_44749,N_38877,N_38384);
xnor U44750 (N_44750,N_35887,N_37464);
and U44751 (N_44751,N_35587,N_36612);
xor U44752 (N_44752,N_39335,N_37109);
xnor U44753 (N_44753,N_36649,N_39938);
and U44754 (N_44754,N_39727,N_39729);
and U44755 (N_44755,N_39655,N_38497);
or U44756 (N_44756,N_35790,N_38340);
nand U44757 (N_44757,N_39681,N_39321);
nor U44758 (N_44758,N_35591,N_36747);
or U44759 (N_44759,N_36012,N_37318);
or U44760 (N_44760,N_36728,N_38991);
or U44761 (N_44761,N_36375,N_37777);
nor U44762 (N_44762,N_39879,N_37077);
or U44763 (N_44763,N_38059,N_36315);
nor U44764 (N_44764,N_38198,N_38690);
nand U44765 (N_44765,N_38905,N_37040);
nor U44766 (N_44766,N_35857,N_38593);
xor U44767 (N_44767,N_39210,N_39275);
or U44768 (N_44768,N_38087,N_39552);
nor U44769 (N_44769,N_36231,N_36263);
and U44770 (N_44770,N_37491,N_36397);
xor U44771 (N_44771,N_38136,N_38110);
and U44772 (N_44772,N_39935,N_37033);
nor U44773 (N_44773,N_35054,N_35950);
xor U44774 (N_44774,N_36234,N_39582);
xnor U44775 (N_44775,N_36218,N_37807);
nand U44776 (N_44776,N_35761,N_39461);
nand U44777 (N_44777,N_37509,N_37944);
nor U44778 (N_44778,N_37736,N_37881);
xor U44779 (N_44779,N_35304,N_39378);
nand U44780 (N_44780,N_35878,N_39890);
xor U44781 (N_44781,N_36726,N_36716);
and U44782 (N_44782,N_35053,N_39960);
xnor U44783 (N_44783,N_39261,N_37101);
nand U44784 (N_44784,N_35979,N_35717);
and U44785 (N_44785,N_36413,N_35285);
or U44786 (N_44786,N_36067,N_39302);
nand U44787 (N_44787,N_38242,N_39859);
nor U44788 (N_44788,N_38590,N_37001);
nand U44789 (N_44789,N_36925,N_35548);
or U44790 (N_44790,N_36613,N_37329);
or U44791 (N_44791,N_35971,N_36679);
nand U44792 (N_44792,N_38937,N_39090);
or U44793 (N_44793,N_35486,N_36503);
nor U44794 (N_44794,N_39404,N_38774);
nand U44795 (N_44795,N_39762,N_37645);
nor U44796 (N_44796,N_35496,N_37800);
nand U44797 (N_44797,N_39920,N_39632);
and U44798 (N_44798,N_36577,N_39619);
xor U44799 (N_44799,N_36541,N_35869);
or U44800 (N_44800,N_35073,N_39909);
nor U44801 (N_44801,N_36761,N_39734);
and U44802 (N_44802,N_35398,N_35239);
nor U44803 (N_44803,N_36343,N_38312);
or U44804 (N_44804,N_35335,N_37684);
nand U44805 (N_44805,N_35533,N_37174);
or U44806 (N_44806,N_36640,N_39505);
and U44807 (N_44807,N_35644,N_39039);
xor U44808 (N_44808,N_38115,N_39946);
and U44809 (N_44809,N_36767,N_36110);
nor U44810 (N_44810,N_39849,N_39167);
xor U44811 (N_44811,N_35581,N_37634);
nand U44812 (N_44812,N_37454,N_39594);
nand U44813 (N_44813,N_36134,N_35412);
and U44814 (N_44814,N_35610,N_37257);
or U44815 (N_44815,N_37461,N_35895);
or U44816 (N_44816,N_37178,N_35297);
nand U44817 (N_44817,N_39973,N_35613);
and U44818 (N_44818,N_35017,N_36030);
and U44819 (N_44819,N_37611,N_36722);
nor U44820 (N_44820,N_38716,N_38454);
nand U44821 (N_44821,N_39342,N_37499);
nand U44822 (N_44822,N_39711,N_36472);
xor U44823 (N_44823,N_37963,N_39572);
xor U44824 (N_44824,N_36487,N_35026);
nor U44825 (N_44825,N_39706,N_37307);
nand U44826 (N_44826,N_35974,N_37564);
xnor U44827 (N_44827,N_36020,N_36838);
or U44828 (N_44828,N_37239,N_36058);
or U44829 (N_44829,N_37321,N_38262);
nand U44830 (N_44830,N_37075,N_39681);
xnor U44831 (N_44831,N_37869,N_39863);
nor U44832 (N_44832,N_35158,N_36815);
or U44833 (N_44833,N_36280,N_37733);
xnor U44834 (N_44834,N_39022,N_35859);
and U44835 (N_44835,N_38432,N_36646);
or U44836 (N_44836,N_39770,N_35144);
nor U44837 (N_44837,N_36812,N_37432);
nor U44838 (N_44838,N_37702,N_36232);
nand U44839 (N_44839,N_37092,N_35182);
nor U44840 (N_44840,N_39283,N_35689);
or U44841 (N_44841,N_38902,N_35478);
xnor U44842 (N_44842,N_36725,N_35943);
or U44843 (N_44843,N_37195,N_36599);
and U44844 (N_44844,N_39961,N_38176);
and U44845 (N_44845,N_38434,N_36210);
nand U44846 (N_44846,N_36819,N_37707);
xor U44847 (N_44847,N_36636,N_37255);
or U44848 (N_44848,N_39744,N_38679);
and U44849 (N_44849,N_36586,N_36581);
or U44850 (N_44850,N_36683,N_38938);
or U44851 (N_44851,N_39209,N_39363);
nor U44852 (N_44852,N_35699,N_35640);
nand U44853 (N_44853,N_35822,N_39345);
xor U44854 (N_44854,N_35054,N_39752);
and U44855 (N_44855,N_39023,N_36434);
nand U44856 (N_44856,N_36145,N_38834);
nand U44857 (N_44857,N_36917,N_38685);
and U44858 (N_44858,N_38582,N_36226);
nand U44859 (N_44859,N_39466,N_38424);
xor U44860 (N_44860,N_39257,N_35412);
and U44861 (N_44861,N_39069,N_39446);
nor U44862 (N_44862,N_36597,N_35206);
and U44863 (N_44863,N_35679,N_38529);
and U44864 (N_44864,N_38934,N_36083);
and U44865 (N_44865,N_36355,N_35168);
nand U44866 (N_44866,N_36508,N_37482);
and U44867 (N_44867,N_39154,N_38189);
and U44868 (N_44868,N_36938,N_39760);
nor U44869 (N_44869,N_35197,N_36359);
and U44870 (N_44870,N_39934,N_37021);
or U44871 (N_44871,N_37389,N_35076);
nand U44872 (N_44872,N_37046,N_36984);
nor U44873 (N_44873,N_38214,N_35605);
or U44874 (N_44874,N_39313,N_39235);
nand U44875 (N_44875,N_36043,N_39580);
xor U44876 (N_44876,N_38998,N_36575);
or U44877 (N_44877,N_39487,N_35125);
xnor U44878 (N_44878,N_38435,N_35628);
or U44879 (N_44879,N_39707,N_35531);
or U44880 (N_44880,N_35231,N_38242);
nor U44881 (N_44881,N_36519,N_38301);
nor U44882 (N_44882,N_36499,N_38505);
nor U44883 (N_44883,N_36632,N_39738);
nor U44884 (N_44884,N_37578,N_35622);
or U44885 (N_44885,N_35617,N_39428);
nor U44886 (N_44886,N_38223,N_35390);
nand U44887 (N_44887,N_39901,N_37033);
and U44888 (N_44888,N_38135,N_38323);
nor U44889 (N_44889,N_39123,N_36990);
nand U44890 (N_44890,N_35975,N_39209);
and U44891 (N_44891,N_38277,N_37181);
or U44892 (N_44892,N_36956,N_39919);
or U44893 (N_44893,N_37053,N_36875);
nand U44894 (N_44894,N_36172,N_37337);
xor U44895 (N_44895,N_36408,N_35875);
and U44896 (N_44896,N_36919,N_37746);
nand U44897 (N_44897,N_35597,N_35747);
or U44898 (N_44898,N_35953,N_36917);
xor U44899 (N_44899,N_38777,N_38570);
nand U44900 (N_44900,N_38271,N_37410);
xnor U44901 (N_44901,N_36628,N_37090);
xor U44902 (N_44902,N_38514,N_38432);
or U44903 (N_44903,N_39531,N_37648);
xor U44904 (N_44904,N_36081,N_38530);
nor U44905 (N_44905,N_37442,N_36805);
nand U44906 (N_44906,N_35959,N_35170);
nand U44907 (N_44907,N_35939,N_37350);
nand U44908 (N_44908,N_35596,N_37583);
nand U44909 (N_44909,N_37533,N_35854);
or U44910 (N_44910,N_36424,N_38284);
nor U44911 (N_44911,N_38221,N_38032);
nor U44912 (N_44912,N_36266,N_35903);
nand U44913 (N_44913,N_38463,N_36207);
nand U44914 (N_44914,N_37214,N_39325);
xnor U44915 (N_44915,N_35794,N_36552);
nor U44916 (N_44916,N_37563,N_36678);
nor U44917 (N_44917,N_37005,N_35791);
nand U44918 (N_44918,N_39887,N_37929);
xnor U44919 (N_44919,N_35353,N_37456);
xnor U44920 (N_44920,N_37424,N_38928);
and U44921 (N_44921,N_37375,N_37576);
xor U44922 (N_44922,N_39715,N_35418);
xnor U44923 (N_44923,N_35423,N_35685);
xor U44924 (N_44924,N_36671,N_39094);
and U44925 (N_44925,N_39221,N_36548);
or U44926 (N_44926,N_35168,N_36285);
or U44927 (N_44927,N_37594,N_36748);
nand U44928 (N_44928,N_36897,N_39096);
xor U44929 (N_44929,N_36058,N_39809);
nor U44930 (N_44930,N_36052,N_38340);
and U44931 (N_44931,N_35765,N_38544);
nor U44932 (N_44932,N_38929,N_35181);
or U44933 (N_44933,N_38304,N_38761);
nor U44934 (N_44934,N_37207,N_37178);
xnor U44935 (N_44935,N_39793,N_39194);
nand U44936 (N_44936,N_38701,N_36085);
xor U44937 (N_44937,N_39144,N_38445);
xnor U44938 (N_44938,N_38908,N_35325);
nor U44939 (N_44939,N_35395,N_37099);
nand U44940 (N_44940,N_37695,N_35246);
and U44941 (N_44941,N_36923,N_36652);
xnor U44942 (N_44942,N_39449,N_38697);
xor U44943 (N_44943,N_36012,N_38613);
nand U44944 (N_44944,N_39370,N_39184);
nor U44945 (N_44945,N_38687,N_37912);
and U44946 (N_44946,N_36508,N_38184);
nor U44947 (N_44947,N_35823,N_37494);
or U44948 (N_44948,N_36677,N_38967);
xor U44949 (N_44949,N_38151,N_38475);
nor U44950 (N_44950,N_35592,N_35452);
xnor U44951 (N_44951,N_39871,N_36080);
or U44952 (N_44952,N_36787,N_35517);
nor U44953 (N_44953,N_36569,N_38944);
nand U44954 (N_44954,N_37120,N_38082);
xor U44955 (N_44955,N_35155,N_35454);
nor U44956 (N_44956,N_35500,N_36023);
nand U44957 (N_44957,N_37428,N_39605);
nor U44958 (N_44958,N_38205,N_36044);
nor U44959 (N_44959,N_36295,N_39432);
nor U44960 (N_44960,N_35849,N_39037);
nand U44961 (N_44961,N_38241,N_37443);
or U44962 (N_44962,N_36127,N_39164);
nor U44963 (N_44963,N_35797,N_36217);
or U44964 (N_44964,N_37908,N_35103);
and U44965 (N_44965,N_37208,N_37980);
nand U44966 (N_44966,N_37753,N_38090);
xor U44967 (N_44967,N_37573,N_36945);
xor U44968 (N_44968,N_39488,N_39943);
nor U44969 (N_44969,N_38357,N_35758);
or U44970 (N_44970,N_37198,N_36007);
xor U44971 (N_44971,N_39421,N_38769);
and U44972 (N_44972,N_39776,N_35279);
xor U44973 (N_44973,N_39776,N_35065);
or U44974 (N_44974,N_38084,N_36745);
nand U44975 (N_44975,N_38434,N_35723);
nor U44976 (N_44976,N_38519,N_35405);
and U44977 (N_44977,N_37085,N_35818);
nand U44978 (N_44978,N_37503,N_38217);
nor U44979 (N_44979,N_39106,N_38358);
xnor U44980 (N_44980,N_35524,N_38127);
or U44981 (N_44981,N_37201,N_36666);
nor U44982 (N_44982,N_35557,N_37033);
nor U44983 (N_44983,N_39217,N_37177);
and U44984 (N_44984,N_35796,N_35795);
nand U44985 (N_44985,N_36195,N_36673);
and U44986 (N_44986,N_35619,N_39714);
xor U44987 (N_44987,N_35498,N_38191);
nand U44988 (N_44988,N_39546,N_37568);
xnor U44989 (N_44989,N_37894,N_38298);
nor U44990 (N_44990,N_39549,N_35695);
nor U44991 (N_44991,N_37503,N_39033);
and U44992 (N_44992,N_38970,N_37861);
or U44993 (N_44993,N_37487,N_38310);
nor U44994 (N_44994,N_35093,N_38225);
nand U44995 (N_44995,N_35884,N_35604);
xor U44996 (N_44996,N_38249,N_38381);
xnor U44997 (N_44997,N_39984,N_37848);
and U44998 (N_44998,N_39882,N_36388);
nor U44999 (N_44999,N_37241,N_38231);
nand U45000 (N_45000,N_41525,N_43990);
nand U45001 (N_45001,N_41482,N_44097);
nor U45002 (N_45002,N_42618,N_43662);
nand U45003 (N_45003,N_42743,N_44481);
and U45004 (N_45004,N_44425,N_43544);
xor U45005 (N_45005,N_41669,N_42348);
and U45006 (N_45006,N_43713,N_43198);
nand U45007 (N_45007,N_44270,N_44666);
nand U45008 (N_45008,N_44434,N_40665);
xnor U45009 (N_45009,N_40875,N_40310);
xor U45010 (N_45010,N_40801,N_42909);
nand U45011 (N_45011,N_40193,N_44935);
nand U45012 (N_45012,N_44546,N_42509);
xnor U45013 (N_45013,N_44934,N_43059);
nand U45014 (N_45014,N_44414,N_40189);
or U45015 (N_45015,N_43040,N_42475);
xor U45016 (N_45016,N_40485,N_43307);
nand U45017 (N_45017,N_40768,N_43365);
xnor U45018 (N_45018,N_44537,N_42110);
nor U45019 (N_45019,N_42032,N_44592);
or U45020 (N_45020,N_44337,N_43354);
xor U45021 (N_45021,N_40754,N_42931);
and U45022 (N_45022,N_44076,N_44526);
or U45023 (N_45023,N_40976,N_43344);
nand U45024 (N_45024,N_41441,N_41010);
nand U45025 (N_45025,N_44602,N_40314);
xnor U45026 (N_45026,N_43087,N_44564);
or U45027 (N_45027,N_41803,N_43734);
nand U45028 (N_45028,N_40234,N_44792);
nor U45029 (N_45029,N_44961,N_40970);
or U45030 (N_45030,N_41367,N_41090);
or U45031 (N_45031,N_41458,N_41487);
nor U45032 (N_45032,N_42470,N_41602);
nor U45033 (N_45033,N_40795,N_44018);
xnor U45034 (N_45034,N_41480,N_42222);
or U45035 (N_45035,N_44755,N_42825);
xnor U45036 (N_45036,N_40915,N_41930);
and U45037 (N_45037,N_43751,N_40027);
and U45038 (N_45038,N_41667,N_44279);
or U45039 (N_45039,N_41318,N_44585);
or U45040 (N_45040,N_41808,N_43954);
nor U45041 (N_45041,N_42734,N_44743);
or U45042 (N_45042,N_42327,N_40625);
xnor U45043 (N_45043,N_44290,N_44143);
xnor U45044 (N_45044,N_42691,N_41864);
xnor U45045 (N_45045,N_42882,N_42566);
nand U45046 (N_45046,N_41361,N_40644);
nand U45047 (N_45047,N_41842,N_44895);
or U45048 (N_45048,N_43572,N_42506);
nor U45049 (N_45049,N_44883,N_40999);
xnor U45050 (N_45050,N_41511,N_44039);
and U45051 (N_45051,N_43542,N_44408);
and U45052 (N_45052,N_43188,N_40538);
and U45053 (N_45053,N_44104,N_43810);
or U45054 (N_45054,N_41611,N_40524);
nor U45055 (N_45055,N_43639,N_41261);
nand U45056 (N_45056,N_42605,N_41568);
and U45057 (N_45057,N_40652,N_40537);
and U45058 (N_45058,N_41969,N_40765);
nand U45059 (N_45059,N_43591,N_43192);
nor U45060 (N_45060,N_44350,N_41530);
or U45061 (N_45061,N_43057,N_42558);
or U45062 (N_45062,N_40143,N_40706);
xor U45063 (N_45063,N_41027,N_42805);
and U45064 (N_45064,N_44791,N_42568);
or U45065 (N_45065,N_40584,N_40482);
nand U45066 (N_45066,N_44102,N_41160);
nand U45067 (N_45067,N_41211,N_42384);
nand U45068 (N_45068,N_42742,N_41134);
nor U45069 (N_45069,N_43285,N_44413);
or U45070 (N_45070,N_42156,N_43458);
xnor U45071 (N_45071,N_42923,N_43688);
or U45072 (N_45072,N_40006,N_44927);
and U45073 (N_45073,N_42541,N_44074);
or U45074 (N_45074,N_40924,N_41861);
and U45075 (N_45075,N_41491,N_40009);
and U45076 (N_45076,N_40983,N_42940);
or U45077 (N_45077,N_40592,N_40435);
or U45078 (N_45078,N_44432,N_41989);
xor U45079 (N_45079,N_43903,N_41396);
nor U45080 (N_45080,N_41682,N_41642);
and U45081 (N_45081,N_41300,N_43674);
and U45082 (N_45082,N_43958,N_41745);
xor U45083 (N_45083,N_42154,N_40626);
nor U45084 (N_45084,N_42946,N_40406);
nand U45085 (N_45085,N_43024,N_41323);
xor U45086 (N_45086,N_41932,N_41869);
and U45087 (N_45087,N_44750,N_41496);
nand U45088 (N_45088,N_42696,N_41684);
or U45089 (N_45089,N_44989,N_43876);
and U45090 (N_45090,N_43573,N_42853);
xnor U45091 (N_45091,N_44171,N_40546);
nor U45092 (N_45092,N_44304,N_43977);
xnor U45093 (N_45093,N_40569,N_44158);
xnor U45094 (N_45094,N_40530,N_44181);
nor U45095 (N_45095,N_42177,N_41689);
or U45096 (N_45096,N_41192,N_43604);
and U45097 (N_45097,N_44735,N_43871);
and U45098 (N_45098,N_42326,N_41529);
xor U45099 (N_45099,N_41003,N_40883);
xor U45100 (N_45100,N_42397,N_41537);
nand U45101 (N_45101,N_43250,N_40588);
or U45102 (N_45102,N_42792,N_44229);
nand U45103 (N_45103,N_42037,N_41133);
xor U45104 (N_45104,N_44393,N_40283);
and U45105 (N_45105,N_40824,N_40511);
xor U45106 (N_45106,N_43756,N_41651);
nor U45107 (N_45107,N_42720,N_44625);
and U45108 (N_45108,N_42108,N_43816);
xor U45109 (N_45109,N_41325,N_40750);
nand U45110 (N_45110,N_44411,N_44294);
and U45111 (N_45111,N_40220,N_41687);
nand U45112 (N_45112,N_43656,N_44710);
and U45113 (N_45113,N_43174,N_43461);
xor U45114 (N_45114,N_43730,N_40050);
nor U45115 (N_45115,N_41424,N_41650);
and U45116 (N_45116,N_42984,N_40807);
nand U45117 (N_45117,N_43923,N_40829);
nand U45118 (N_45118,N_44347,N_43375);
xnor U45119 (N_45119,N_44015,N_44921);
nor U45120 (N_45120,N_40746,N_43237);
or U45121 (N_45121,N_43817,N_41970);
xor U45122 (N_45122,N_41117,N_40835);
nor U45123 (N_45123,N_44151,N_41404);
nand U45124 (N_45124,N_41303,N_40262);
xnor U45125 (N_45125,N_40430,N_42235);
or U45126 (N_45126,N_40440,N_41370);
nor U45127 (N_45127,N_44048,N_42416);
xnor U45128 (N_45128,N_43044,N_41958);
nor U45129 (N_45129,N_43380,N_41654);
and U45130 (N_45130,N_41384,N_40491);
nor U45131 (N_45131,N_40529,N_40198);
and U45132 (N_45132,N_40912,N_41196);
and U45133 (N_45133,N_44964,N_41783);
xor U45134 (N_45134,N_43624,N_41671);
xor U45135 (N_45135,N_42545,N_43254);
xnor U45136 (N_45136,N_43212,N_41101);
and U45137 (N_45137,N_40167,N_44569);
xnor U45138 (N_45138,N_41715,N_44781);
xnor U45139 (N_45139,N_40036,N_42058);
xnor U45140 (N_45140,N_41900,N_42547);
nor U45141 (N_45141,N_42074,N_40145);
xor U45142 (N_45142,N_43006,N_41005);
and U45143 (N_45143,N_40926,N_42823);
nor U45144 (N_45144,N_43852,N_42829);
nor U45145 (N_45145,N_44253,N_43909);
or U45146 (N_45146,N_40270,N_42574);
nor U45147 (N_45147,N_42069,N_44706);
nor U45148 (N_45148,N_43336,N_41157);
nor U45149 (N_45149,N_42970,N_44506);
nor U45150 (N_45150,N_42758,N_41412);
nor U45151 (N_45151,N_44700,N_42830);
or U45152 (N_45152,N_41341,N_42698);
and U45153 (N_45153,N_40183,N_41416);
xnor U45154 (N_45154,N_43549,N_41193);
xor U45155 (N_45155,N_43041,N_44619);
nand U45156 (N_45156,N_42524,N_41891);
or U45157 (N_45157,N_43889,N_42878);
and U45158 (N_45158,N_42025,N_41702);
and U45159 (N_45159,N_42081,N_44802);
nor U45160 (N_45160,N_43866,N_40423);
and U45161 (N_45161,N_40077,N_40506);
nand U45162 (N_45162,N_42113,N_41378);
xor U45163 (N_45163,N_41645,N_40536);
nand U45164 (N_45164,N_42866,N_44522);
or U45165 (N_45165,N_40097,N_43182);
nor U45166 (N_45166,N_40995,N_42392);
and U45167 (N_45167,N_43640,N_43914);
xnor U45168 (N_45168,N_43614,N_41169);
and U45169 (N_45169,N_43769,N_43615);
nand U45170 (N_45170,N_41678,N_42738);
nand U45171 (N_45171,N_41968,N_40636);
nand U45172 (N_45172,N_43488,N_40574);
and U45173 (N_45173,N_40522,N_42057);
nand U45174 (N_45174,N_40560,N_42442);
xor U45175 (N_45175,N_40195,N_43781);
xor U45176 (N_45176,N_44795,N_42939);
nand U45177 (N_45177,N_44343,N_40273);
nor U45178 (N_45178,N_43976,N_44361);
xnor U45179 (N_45179,N_42906,N_40732);
nor U45180 (N_45180,N_43595,N_40377);
nor U45181 (N_45181,N_44949,N_43811);
or U45182 (N_45182,N_43278,N_43943);
nor U45183 (N_45183,N_44046,N_44129);
nor U45184 (N_45184,N_44331,N_42471);
and U45185 (N_45185,N_40532,N_44184);
nor U45186 (N_45186,N_42644,N_44991);
xor U45187 (N_45187,N_43989,N_44212);
nand U45188 (N_45188,N_42672,N_41841);
or U45189 (N_45189,N_41171,N_40129);
nand U45190 (N_45190,N_42255,N_41987);
nor U45191 (N_45191,N_43991,N_41610);
xnor U45192 (N_45192,N_44175,N_42234);
xnor U45193 (N_45193,N_41447,N_43825);
nor U45194 (N_45194,N_42662,N_41121);
or U45195 (N_45195,N_40771,N_43176);
and U45196 (N_45196,N_42847,N_42903);
and U45197 (N_45197,N_43735,N_43398);
or U45198 (N_45198,N_40638,N_41187);
xor U45199 (N_45199,N_44507,N_43102);
nor U45200 (N_45200,N_41538,N_42907);
and U45201 (N_45201,N_42010,N_44876);
or U45202 (N_45202,N_44003,N_44038);
or U45203 (N_45203,N_41259,N_44589);
nor U45204 (N_45204,N_42701,N_40397);
xor U45205 (N_45205,N_44868,N_43204);
nand U45206 (N_45206,N_43761,N_43140);
nand U45207 (N_45207,N_43642,N_41631);
nor U45208 (N_45208,N_41024,N_42223);
or U45209 (N_45209,N_41852,N_40150);
or U45210 (N_45210,N_41348,N_44887);
and U45211 (N_45211,N_43519,N_42400);
xor U45212 (N_45212,N_41552,N_43100);
or U45213 (N_45213,N_43629,N_43266);
nor U45214 (N_45214,N_42135,N_42925);
xor U45215 (N_45215,N_42964,N_42789);
nor U45216 (N_45216,N_43167,N_40842);
and U45217 (N_45217,N_41223,N_40816);
or U45218 (N_45218,N_40047,N_41419);
nor U45219 (N_45219,N_41203,N_41063);
or U45220 (N_45220,N_41004,N_42368);
or U45221 (N_45221,N_43836,N_44892);
and U45222 (N_45222,N_44012,N_44006);
or U45223 (N_45223,N_43352,N_40596);
and U45224 (N_45224,N_44977,N_43585);
nand U45225 (N_45225,N_42752,N_42050);
nor U45226 (N_45226,N_42928,N_42033);
and U45227 (N_45227,N_42601,N_42669);
nand U45228 (N_45228,N_43547,N_44079);
nor U45229 (N_45229,N_41204,N_43228);
xnor U45230 (N_45230,N_41536,N_44731);
nor U45231 (N_45231,N_42841,N_41020);
and U45232 (N_45232,N_40320,N_42873);
nand U45233 (N_45233,N_44732,N_44264);
or U45234 (N_45234,N_44647,N_43881);
nand U45235 (N_45235,N_42085,N_44156);
nand U45236 (N_45236,N_42862,N_41104);
nor U45237 (N_45237,N_44226,N_41657);
or U45238 (N_45238,N_44520,N_43835);
nand U45239 (N_45239,N_40725,N_41385);
xnor U45240 (N_45240,N_40024,N_40632);
nor U45241 (N_45241,N_41840,N_43789);
xor U45242 (N_45242,N_42374,N_42371);
nor U45243 (N_45243,N_43370,N_44951);
and U45244 (N_45244,N_41873,N_44775);
and U45245 (N_45245,N_43478,N_44099);
nor U45246 (N_45246,N_43259,N_41199);
and U45247 (N_45247,N_40082,N_43736);
or U45248 (N_45248,N_43834,N_41307);
xor U45249 (N_45249,N_43243,N_42351);
xnor U45250 (N_45250,N_42459,N_40822);
nand U45251 (N_45251,N_43828,N_41890);
nor U45252 (N_45252,N_44349,N_41519);
and U45253 (N_45253,N_43805,N_43199);
or U45254 (N_45254,N_40434,N_41084);
nand U45255 (N_45255,N_44453,N_44418);
or U45256 (N_45256,N_40663,N_42477);
or U45257 (N_45257,N_44634,N_40263);
nor U45258 (N_45258,N_40882,N_41036);
xnor U45259 (N_45259,N_42540,N_40940);
or U45260 (N_45260,N_40726,N_43104);
nor U45261 (N_45261,N_44769,N_40946);
nor U45262 (N_45262,N_44445,N_41079);
nand U45263 (N_45263,N_42994,N_44239);
nand U45264 (N_45264,N_40080,N_41432);
and U45265 (N_45265,N_40634,N_43062);
and U45266 (N_45266,N_44225,N_40897);
nand U45267 (N_45267,N_43251,N_42163);
nor U45268 (N_45268,N_43854,N_40555);
and U45269 (N_45269,N_42158,N_44227);
nand U45270 (N_45270,N_41787,N_40087);
or U45271 (N_45271,N_41763,N_41945);
xor U45272 (N_45272,N_42622,N_40982);
xnor U45273 (N_45273,N_41793,N_40114);
xor U45274 (N_45274,N_43879,N_44306);
nor U45275 (N_45275,N_40952,N_42063);
nand U45276 (N_45276,N_43080,N_43890);
and U45277 (N_45277,N_40595,N_40023);
or U45278 (N_45278,N_43492,N_42275);
or U45279 (N_45279,N_40798,N_44093);
and U45280 (N_45280,N_44482,N_41995);
nor U45281 (N_45281,N_40950,N_40229);
nor U45282 (N_45282,N_43043,N_40691);
nor U45283 (N_45283,N_44494,N_41697);
nor U45284 (N_45284,N_40639,N_43306);
xnor U45285 (N_45285,N_40606,N_44947);
and U45286 (N_45286,N_43514,N_43787);
xnor U45287 (N_45287,N_43779,N_42487);
and U45288 (N_45288,N_42003,N_42145);
or U45289 (N_45289,N_40155,N_40741);
xor U45290 (N_45290,N_42686,N_44815);
and U45291 (N_45291,N_43754,N_42491);
nor U45292 (N_45292,N_44152,N_40124);
and U45293 (N_45293,N_40113,N_41640);
nor U45294 (N_45294,N_43130,N_40216);
or U45295 (N_45295,N_43540,N_42856);
or U45296 (N_45296,N_42211,N_44773);
or U45297 (N_45297,N_44441,N_41755);
nand U45298 (N_45298,N_43555,N_44861);
xnor U45299 (N_45299,N_40572,N_41163);
nor U45300 (N_45300,N_43063,N_42339);
xor U45301 (N_45301,N_42100,N_44704);
xnor U45302 (N_45302,N_41469,N_43728);
xnor U45303 (N_45303,N_41288,N_42298);
and U45304 (N_45304,N_44095,N_42592);
nor U45305 (N_45305,N_40866,N_42246);
nor U45306 (N_45306,N_40432,N_42630);
and U45307 (N_45307,N_41878,N_42412);
and U45308 (N_45308,N_42771,N_43103);
and U45309 (N_45309,N_44050,N_44386);
nand U45310 (N_45310,N_40031,N_44941);
nor U45311 (N_45311,N_44409,N_42353);
or U45312 (N_45312,N_42563,N_43466);
xnor U45313 (N_45313,N_42122,N_42242);
and U45314 (N_45314,N_42510,N_40965);
xnor U45315 (N_45315,N_43833,N_42681);
xor U45316 (N_45316,N_42450,N_40547);
nand U45317 (N_45317,N_41912,N_44889);
nand U45318 (N_45318,N_41733,N_44673);
nand U45319 (N_45319,N_40608,N_41732);
nand U45320 (N_45320,N_40543,N_43635);
or U45321 (N_45321,N_43911,N_42064);
xor U45322 (N_45322,N_44854,N_42851);
and U45323 (N_45323,N_41350,N_43297);
and U45324 (N_45324,N_43382,N_44450);
nor U45325 (N_45325,N_41159,N_44501);
nand U45326 (N_45326,N_43993,N_44240);
nand U45327 (N_45327,N_42983,N_44500);
nor U45328 (N_45328,N_41575,N_41479);
xnor U45329 (N_45329,N_40980,N_42913);
nor U45330 (N_45330,N_40601,N_43785);
xor U45331 (N_45331,N_44163,N_43858);
or U45332 (N_45332,N_42167,N_42581);
nor U45333 (N_45333,N_43244,N_42286);
and U45334 (N_45334,N_44913,N_41809);
xnor U45335 (N_45335,N_43027,N_43669);
xor U45336 (N_45336,N_40154,N_40045);
and U45337 (N_45337,N_41607,N_40773);
nor U45338 (N_45338,N_43312,N_41100);
nor U45339 (N_45339,N_40000,N_42075);
xnor U45340 (N_45340,N_40762,N_42590);
nand U45341 (N_45341,N_42208,N_42249);
nor U45342 (N_45342,N_44816,N_41009);
nor U45343 (N_45343,N_42214,N_41670);
nand U45344 (N_45344,N_41465,N_43113);
nand U45345 (N_45345,N_41413,N_41843);
nand U45346 (N_45346,N_43288,N_40730);
or U45347 (N_45347,N_40677,N_44203);
nand U45348 (N_45348,N_41521,N_43839);
and U45349 (N_45349,N_44812,N_44684);
and U45350 (N_45350,N_44907,N_43275);
or U45351 (N_45351,N_44374,N_40056);
and U45352 (N_45352,N_44696,N_41835);
xnor U45353 (N_45353,N_40831,N_40052);
xnor U45354 (N_45354,N_41927,N_42857);
and U45355 (N_45355,N_44479,N_43632);
xor U45356 (N_45356,N_43843,N_44954);
and U45357 (N_45357,N_42201,N_43981);
and U45358 (N_45358,N_43508,N_44528);
nand U45359 (N_45359,N_44348,N_43536);
nand U45360 (N_45360,N_44842,N_42889);
xnor U45361 (N_45361,N_44255,N_42318);
xnor U45362 (N_45362,N_44274,N_44745);
xor U45363 (N_45363,N_43141,N_41097);
xnor U45364 (N_45364,N_44643,N_41831);
xor U45365 (N_45365,N_41218,N_40810);
xnor U45366 (N_45366,N_42048,N_43047);
nor U45367 (N_45367,N_43533,N_44182);
and U45368 (N_45368,N_41254,N_43011);
or U45369 (N_45369,N_44410,N_40736);
nand U45370 (N_45370,N_41032,N_43242);
nor U45371 (N_45371,N_44194,N_42272);
nand U45372 (N_45372,N_42276,N_40863);
nand U45373 (N_45373,N_43133,N_43528);
and U45374 (N_45374,N_41474,N_44114);
or U45375 (N_45375,N_41500,N_40439);
or U45376 (N_45376,N_42842,N_42804);
nor U45377 (N_45377,N_40680,N_43737);
nor U45378 (N_45378,N_43837,N_42452);
and U45379 (N_45379,N_42807,N_41504);
or U45380 (N_45380,N_43289,N_42800);
and U45381 (N_45381,N_43733,N_42653);
and U45382 (N_45382,N_42306,N_42355);
and U45383 (N_45383,N_42591,N_42257);
and U45384 (N_45384,N_43806,N_42426);
xnor U45385 (N_45385,N_42930,N_44944);
and U45386 (N_45386,N_40141,N_40269);
or U45387 (N_45387,N_43869,N_41235);
nor U45388 (N_45388,N_41944,N_43822);
and U45389 (N_45389,N_42582,N_40481);
or U45390 (N_45390,N_44258,N_40748);
or U45391 (N_45391,N_43601,N_43083);
or U45392 (N_45392,N_40947,N_44424);
or U45393 (N_45393,N_44514,N_42949);
nand U45394 (N_45394,N_42405,N_44578);
or U45395 (N_45395,N_40731,N_44397);
or U45396 (N_45396,N_44025,N_43137);
xor U45397 (N_45397,N_40046,N_41053);
xor U45398 (N_45398,N_42224,N_40176);
or U45399 (N_45399,N_40015,N_42526);
nand U45400 (N_45400,N_43791,N_42036);
nand U45401 (N_45401,N_41872,N_43746);
nor U45402 (N_45402,N_44800,N_42365);
nor U45403 (N_45403,N_41372,N_43218);
or U45404 (N_45404,N_40668,N_43792);
and U45405 (N_45405,N_43868,N_41178);
nand U45406 (N_45406,N_41085,N_43767);
nand U45407 (N_45407,N_41105,N_41527);
and U45408 (N_45408,N_40065,N_40782);
nand U45409 (N_45409,N_41179,N_44694);
or U45410 (N_45410,N_43227,N_43527);
or U45411 (N_45411,N_44828,N_41015);
and U45412 (N_45412,N_42718,N_42107);
nand U45413 (N_45413,N_42958,N_41811);
nand U45414 (N_45414,N_44049,N_41414);
or U45415 (N_45415,N_44936,N_42457);
or U45416 (N_45416,N_44000,N_40276);
xnor U45417 (N_45417,N_40819,N_43502);
or U45418 (N_45418,N_43064,N_43223);
nor U45419 (N_45419,N_43195,N_40694);
and U45420 (N_45420,N_42456,N_40914);
nand U45421 (N_45421,N_41124,N_44945);
nand U45422 (N_45422,N_44068,N_40319);
nor U45423 (N_45423,N_42231,N_43768);
or U45424 (N_45424,N_42640,N_43951);
xnor U45425 (N_45425,N_42240,N_43972);
and U45426 (N_45426,N_43975,N_43487);
xor U45427 (N_45427,N_43968,N_44466);
or U45428 (N_45428,N_43337,N_41782);
nand U45429 (N_45429,N_44768,N_43494);
nand U45430 (N_45430,N_41749,N_40450);
and U45431 (N_45431,N_44319,N_42082);
nor U45432 (N_45432,N_40989,N_40655);
xnor U45433 (N_45433,N_43532,N_41127);
or U45434 (N_45434,N_40772,N_40007);
or U45435 (N_45435,N_42359,N_40421);
and U45436 (N_45436,N_43727,N_40647);
nor U45437 (N_45437,N_42944,N_43631);
or U45438 (N_45438,N_40932,N_43840);
or U45439 (N_45439,N_40437,N_41909);
xnor U45440 (N_45440,N_40629,N_44044);
or U45441 (N_45441,N_41923,N_42362);
nand U45442 (N_45442,N_40681,N_43477);
xor U45443 (N_45443,N_41244,N_43281);
or U45444 (N_45444,N_44621,N_41423);
nor U45445 (N_45445,N_43170,N_41400);
xor U45446 (N_45446,N_41227,N_40303);
and U45447 (N_45447,N_41125,N_40117);
xnor U45448 (N_45448,N_42200,N_43691);
nand U45449 (N_45449,N_42103,N_44254);
xnor U45450 (N_45450,N_43098,N_44549);
xnor U45451 (N_45451,N_43623,N_42389);
nor U45452 (N_45452,N_42833,N_44760);
or U45453 (N_45453,N_44185,N_41531);
nor U45454 (N_45454,N_41477,N_41436);
or U45455 (N_45455,N_40541,N_42514);
nand U45456 (N_45456,N_41734,N_41076);
or U45457 (N_45457,N_40488,N_42097);
nand U45458 (N_45458,N_42756,N_42285);
or U45459 (N_45459,N_44273,N_42824);
or U45460 (N_45460,N_41248,N_41088);
nor U45461 (N_45461,N_43740,N_44765);
and U45462 (N_45462,N_42594,N_41761);
or U45463 (N_45463,N_44882,N_44461);
nor U45464 (N_45464,N_41446,N_40177);
and U45465 (N_45465,N_40159,N_42625);
nand U45466 (N_45466,N_40548,N_41172);
xor U45467 (N_45467,N_43016,N_44512);
or U45468 (N_45468,N_42380,N_41660);
nor U45469 (N_45469,N_40783,N_41991);
and U45470 (N_45470,N_42973,N_41295);
and U45471 (N_45471,N_43543,N_40757);
nor U45472 (N_45472,N_43596,N_42479);
xnor U45473 (N_45473,N_43898,N_41791);
or U45474 (N_45474,N_40436,N_43798);
and U45475 (N_45475,N_42993,N_43763);
or U45476 (N_45476,N_44328,N_42711);
and U45477 (N_45477,N_42736,N_42445);
nor U45478 (N_45478,N_42198,N_44772);
and U45479 (N_45479,N_43467,N_40242);
nand U45480 (N_45480,N_42464,N_42331);
nand U45481 (N_45481,N_40431,N_40418);
nand U45482 (N_45482,N_42521,N_41753);
or U45483 (N_45483,N_40540,N_41397);
xnor U45484 (N_45484,N_42496,N_43731);
nor U45485 (N_45485,N_40252,N_40770);
or U45486 (N_45486,N_43033,N_41886);
nand U45487 (N_45487,N_44309,N_41920);
and U45488 (N_45488,N_40194,N_42264);
nand U45489 (N_45489,N_44297,N_42783);
nor U45490 (N_45490,N_44733,N_43035);
or U45491 (N_45491,N_41850,N_41550);
or U45492 (N_45492,N_43169,N_44631);
xor U45493 (N_45493,N_44122,N_40131);
nand U45494 (N_45494,N_44825,N_41593);
nand U45495 (N_45495,N_41365,N_44837);
and U45496 (N_45496,N_41152,N_44368);
nor U45497 (N_45497,N_40751,N_40362);
nor U45498 (N_45498,N_43607,N_44004);
nor U45499 (N_45499,N_43374,N_40071);
xnor U45500 (N_45500,N_41621,N_41353);
and U45501 (N_45501,N_42030,N_40018);
or U45502 (N_45502,N_44749,N_43205);
and U45503 (N_45503,N_43877,N_43755);
xnor U45504 (N_45504,N_44953,N_42562);
and U45505 (N_45505,N_44804,N_41741);
nor U45506 (N_45506,N_41016,N_43672);
xor U45507 (N_45507,N_44135,N_43219);
or U45508 (N_45508,N_43110,N_41558);
xor U45509 (N_45509,N_42084,N_40166);
nor U45510 (N_45510,N_40956,N_42101);
nor U45511 (N_45511,N_40521,N_40121);
nand U45512 (N_45512,N_44665,N_44189);
and U45513 (N_45513,N_43933,N_42128);
nor U45514 (N_45514,N_44089,N_44125);
nor U45515 (N_45515,N_43155,N_43610);
xor U45516 (N_45516,N_43132,N_43495);
nor U45517 (N_45517,N_40806,N_42334);
xnor U45518 (N_45518,N_40413,N_42375);
or U45519 (N_45519,N_44510,N_41764);
or U45520 (N_45520,N_41613,N_41770);
nand U45521 (N_45521,N_40717,N_40675);
nand U45522 (N_45522,N_41271,N_44010);
nor U45523 (N_45523,N_42806,N_40739);
or U45524 (N_45524,N_43511,N_44077);
nand U45525 (N_45525,N_44860,N_41089);
nor U45526 (N_45526,N_41876,N_44789);
and U45527 (N_45527,N_43960,N_40937);
or U45528 (N_45528,N_42624,N_44636);
nor U45529 (N_45529,N_41478,N_42072);
and U45530 (N_45530,N_41164,N_41108);
and U45531 (N_45531,N_41953,N_41586);
xor U45532 (N_45532,N_41700,N_41266);
nor U45533 (N_45533,N_42409,N_41420);
nor U45534 (N_45534,N_42497,N_42022);
and U45535 (N_45535,N_40173,N_42440);
or U45536 (N_45536,N_43938,N_42687);
nand U45537 (N_45537,N_40698,N_40692);
nor U45538 (N_45538,N_44915,N_43394);
or U45539 (N_45539,N_40582,N_42441);
nor U45540 (N_45540,N_42684,N_41454);
xor U45541 (N_45541,N_41959,N_44833);
nor U45542 (N_45542,N_40387,N_42432);
and U45543 (N_45543,N_44154,N_41492);
nor U45544 (N_45544,N_40539,N_42259);
nor U45545 (N_45545,N_43409,N_43522);
nand U45546 (N_45546,N_40471,N_44641);
nand U45547 (N_45547,N_43929,N_43927);
nand U45548 (N_45548,N_43556,N_41618);
nor U45549 (N_45549,N_43657,N_40920);
nand U45550 (N_45550,N_43826,N_40908);
nor U45551 (N_45551,N_43979,N_44439);
or U45552 (N_45552,N_41138,N_43444);
nand U45553 (N_45553,N_44055,N_43308);
nand U45554 (N_45554,N_40869,N_44906);
nand U45555 (N_45555,N_40854,N_40962);
nor U45556 (N_45556,N_41747,N_44417);
nand U45557 (N_45557,N_43621,N_43025);
nand U45558 (N_45558,N_42619,N_42190);
and U45559 (N_45559,N_41467,N_42765);
nand U45560 (N_45560,N_44435,N_40057);
nor U45561 (N_45561,N_41941,N_41302);
and U45562 (N_45562,N_44443,N_41331);
and U45563 (N_45563,N_44712,N_43628);
or U45564 (N_45564,N_40375,N_42617);
and U45565 (N_45565,N_41317,N_42350);
or U45566 (N_45566,N_41514,N_43844);
and U45567 (N_45567,N_44529,N_41245);
nor U45568 (N_45568,N_43918,N_41986);
or U45569 (N_45569,N_40711,N_44511);
or U45570 (N_45570,N_41595,N_42733);
nand U45571 (N_45571,N_40987,N_41055);
nor U45572 (N_45572,N_41498,N_41691);
and U45573 (N_45573,N_40508,N_43460);
nor U45574 (N_45574,N_40179,N_41115);
xnor U45575 (N_45575,N_42905,N_42537);
and U45576 (N_45576,N_42843,N_43129);
nor U45577 (N_45577,N_42029,N_44862);
nor U45578 (N_45578,N_43368,N_41065);
xor U45579 (N_45579,N_43588,N_43135);
nand U45580 (N_45580,N_44384,N_43996);
nand U45581 (N_45581,N_42040,N_40498);
and U45582 (N_45582,N_44451,N_44365);
xor U45583 (N_45583,N_41542,N_42182);
nand U45584 (N_45584,N_40526,N_42448);
nor U45585 (N_45585,N_40654,N_42166);
nor U45586 (N_45586,N_40852,N_40949);
and U45587 (N_45587,N_44560,N_41949);
nand U45588 (N_45588,N_41429,N_41128);
or U45589 (N_45589,N_43340,N_44841);
or U45590 (N_45590,N_42729,N_40528);
and U45591 (N_45591,N_44686,N_40593);
xor U45592 (N_45592,N_44007,N_42160);
and U45593 (N_45593,N_40653,N_44670);
xor U45594 (N_45594,N_44793,N_41778);
or U45595 (N_45595,N_41584,N_40724);
or U45596 (N_45596,N_40580,N_42626);
and U45597 (N_45597,N_44611,N_44681);
and U45598 (N_45598,N_41810,N_40978);
xnor U45599 (N_45599,N_41546,N_40805);
and U45600 (N_45600,N_40038,N_41379);
nand U45601 (N_45601,N_40709,N_43490);
nand U45602 (N_45602,N_44295,N_44983);
nor U45603 (N_45603,N_42294,N_43974);
and U45604 (N_45604,N_41951,N_40487);
or U45605 (N_45605,N_41590,N_43910);
and U45606 (N_45606,N_44072,N_43338);
or U45607 (N_45607,N_42076,N_41495);
nand U45608 (N_45608,N_42087,N_43964);
nand U45609 (N_45609,N_41450,N_43097);
and U45610 (N_45610,N_43703,N_44237);
or U45611 (N_45611,N_42481,N_43764);
xnor U45612 (N_45612,N_41094,N_41281);
xnor U45613 (N_45613,N_41154,N_44215);
and U45614 (N_45614,N_41442,N_40549);
nand U45615 (N_45615,N_43774,N_42955);
nor U45616 (N_45616,N_42615,N_41408);
nand U45617 (N_45617,N_44886,N_43611);
nand U45618 (N_45618,N_44267,N_41449);
and U45619 (N_45619,N_44758,N_40585);
and U45620 (N_45620,N_44918,N_44094);
xor U45621 (N_45621,N_44790,N_42062);
or U45622 (N_45622,N_44766,N_41870);
and U45623 (N_45623,N_40998,N_44870);
nand U45624 (N_45624,N_42014,N_41013);
xor U45625 (N_45625,N_43395,N_43012);
nand U45626 (N_45626,N_41475,N_44810);
nand U45627 (N_45627,N_40058,N_41683);
nand U45628 (N_45628,N_43807,N_41289);
nor U45629 (N_45629,N_44101,N_43664);
xnor U45630 (N_45630,N_41865,N_42106);
nor U45631 (N_45631,N_43284,N_43094);
nand U45632 (N_45632,N_42606,N_40520);
nand U45633 (N_45633,N_40994,N_43217);
nand U45634 (N_45634,N_41484,N_41405);
and U45635 (N_45635,N_42213,N_41879);
and U45636 (N_45636,N_41309,N_44455);
and U45637 (N_45637,N_41176,N_42123);
or U45638 (N_45638,N_44940,N_41626);
nand U45639 (N_45639,N_41236,N_42340);
xnor U45640 (N_45640,N_40469,N_44740);
or U45641 (N_45641,N_43883,N_43548);
and U45642 (N_45642,N_42611,N_41377);
nor U45643 (N_45643,N_43046,N_43641);
nor U45644 (N_45644,N_40918,N_42358);
and U45645 (N_45645,N_42056,N_42697);
nor U45646 (N_45646,N_44370,N_44463);
nor U45647 (N_45647,N_42891,N_43566);
nor U45648 (N_45648,N_41703,N_42879);
nand U45649 (N_45649,N_40656,N_42760);
nand U45650 (N_45650,N_40374,N_41068);
and U45651 (N_45651,N_41962,N_42472);
nor U45652 (N_45652,N_44955,N_40451);
and U45653 (N_45653,N_41011,N_42155);
nand U45654 (N_45654,N_41389,N_44394);
xnor U45655 (N_45655,N_40637,N_42894);
nand U45656 (N_45656,N_42612,N_44624);
nor U45657 (N_45657,N_42768,N_41622);
and U45658 (N_45658,N_42324,N_44137);
and U45659 (N_45659,N_41116,N_41371);
or U45660 (N_45660,N_44027,N_43017);
nand U45661 (N_45661,N_41262,N_40891);
or U45662 (N_45662,N_44470,N_41239);
nand U45663 (N_45663,N_43687,N_40109);
or U45664 (N_45664,N_41383,N_42478);
or U45665 (N_45665,N_44865,N_44959);
and U45666 (N_45666,N_43955,N_40602);
nand U45667 (N_45667,N_43333,N_43111);
or U45668 (N_45668,N_43450,N_41785);
or U45669 (N_45669,N_41643,N_44912);
nor U45670 (N_45670,N_41756,N_40325);
nand U45671 (N_45671,N_44614,N_44469);
and U45672 (N_45672,N_40938,N_44969);
xnor U45673 (N_45673,N_42726,N_42425);
nor U45674 (N_45674,N_43179,N_44813);
or U45675 (N_45675,N_44498,N_44493);
or U45676 (N_45676,N_43973,N_40222);
or U45677 (N_45677,N_43481,N_40324);
nor U45678 (N_45678,N_44748,N_43020);
or U45679 (N_45679,N_41427,N_44248);
and U45680 (N_45680,N_41533,N_43997);
or U45681 (N_45681,N_44301,N_40158);
and U45682 (N_45682,N_44899,N_42937);
nor U45683 (N_45683,N_44960,N_42370);
nand U45684 (N_45684,N_41114,N_40017);
nand U45685 (N_45685,N_42778,N_42372);
nor U45686 (N_45686,N_41743,N_43850);
nand U45687 (N_45687,N_44399,N_44838);
and U45688 (N_45688,N_42390,N_44782);
xor U45689 (N_45689,N_44799,N_40620);
xor U45690 (N_45690,N_40353,N_42401);
nor U45691 (N_45691,N_40004,N_42092);
nor U45692 (N_45692,N_43626,N_40490);
and U45693 (N_45693,N_43247,N_43729);
xor U45694 (N_45694,N_43031,N_41056);
and U45695 (N_45695,N_40054,N_41091);
nor U45696 (N_45696,N_42858,N_44967);
nor U45697 (N_45697,N_44778,N_42042);
and U45698 (N_45698,N_44342,N_43940);
nor U45699 (N_45699,N_41821,N_40477);
nor U45700 (N_45700,N_43745,N_41535);
nor U45701 (N_45701,N_41571,N_42336);
nor U45702 (N_45702,N_42838,N_40321);
nand U45703 (N_45703,N_40255,N_44353);
and U45704 (N_45704,N_42694,N_40333);
and U45705 (N_45705,N_44797,N_40975);
nand U45706 (N_45706,N_44542,N_42347);
nor U45707 (N_45707,N_43520,N_43268);
or U45708 (N_45708,N_42124,N_40422);
nor U45709 (N_45709,N_43049,N_43917);
nand U45710 (N_45710,N_42817,N_41033);
xnor U45711 (N_45711,N_40881,N_41624);
xnor U45712 (N_45712,N_43439,N_40414);
nor U45713 (N_45713,N_40368,N_41506);
xnor U45714 (N_45714,N_43421,N_42196);
or U45715 (N_45715,N_43002,N_44186);
xnor U45716 (N_45716,N_41041,N_44903);
nand U45717 (N_45717,N_41522,N_44034);
nor U45718 (N_45718,N_43014,N_43575);
nor U45719 (N_45719,N_44310,N_40766);
xor U45720 (N_45720,N_40876,N_44335);
or U45721 (N_45721,N_42349,N_41907);
nand U45722 (N_45722,N_43515,N_40329);
nand U45723 (N_45723,N_43440,N_43554);
or U45724 (N_45724,N_41625,N_44321);
or U45725 (N_45725,N_42835,N_40561);
xnor U45726 (N_45726,N_43241,N_40389);
nor U45727 (N_45727,N_44579,N_44901);
nand U45728 (N_45728,N_41877,N_42572);
nand U45729 (N_45729,N_42245,N_43697);
nor U45730 (N_45730,N_40266,N_42408);
nand U45731 (N_45731,N_44806,N_42034);
or U45732 (N_45732,N_42710,N_43448);
nor U45733 (N_45733,N_44963,N_43353);
xnor U45734 (N_45734,N_43963,N_42776);
xnor U45735 (N_45735,N_44807,N_41398);
or U45736 (N_45736,N_43117,N_44360);
nand U45737 (N_45737,N_43861,N_41139);
or U45738 (N_45738,N_43056,N_40633);
and U45739 (N_45739,N_43928,N_40136);
xor U45740 (N_45740,N_44820,N_44164);
xor U45741 (N_45741,N_43841,N_43862);
or U45742 (N_45742,N_44558,N_41773);
xor U45743 (N_45743,N_44638,N_43603);
and U45744 (N_45744,N_41981,N_44130);
nor U45745 (N_45745,N_41663,N_41561);
nand U45746 (N_45746,N_41815,N_44090);
and U45747 (N_45747,N_43298,N_43474);
nand U45748 (N_45748,N_40925,N_42268);
nor U45749 (N_45749,N_43813,N_41052);
xor U45750 (N_45750,N_40786,N_42536);
or U45751 (N_45751,N_42660,N_40185);
nor U45752 (N_45752,N_44709,N_42585);
and U45753 (N_45753,N_44047,N_41705);
nor U45754 (N_45754,N_41744,N_43470);
or U45755 (N_45755,N_42614,N_40293);
nand U45756 (N_45756,N_42164,N_41950);
nand U45757 (N_45757,N_42966,N_40817);
or U45758 (N_45758,N_40612,N_41410);
xor U45759 (N_45759,N_42577,N_40500);
and U45760 (N_45760,N_42038,N_42692);
nand U45761 (N_45761,N_40452,N_40370);
or U45762 (N_45762,N_43676,N_41863);
xnor U45763 (N_45763,N_43456,N_41078);
or U45764 (N_45764,N_44826,N_41532);
nor U45765 (N_45765,N_43086,N_43932);
nor U45766 (N_45766,N_43946,N_42283);
xor U45767 (N_45767,N_40986,N_44873);
or U45768 (N_45768,N_44262,N_44483);
or U45769 (N_45769,N_40091,N_40820);
or U45770 (N_45770,N_40338,N_40642);
and U45771 (N_45771,N_42171,N_44617);
nand U45772 (N_45772,N_42185,N_44604);
nand U45773 (N_45773,N_42466,N_42205);
nand U45774 (N_45774,N_41232,N_43778);
and U45775 (N_45775,N_41976,N_41294);
or U45776 (N_45776,N_41982,N_44875);
nor U45777 (N_45777,N_43386,N_40108);
or U45778 (N_45778,N_40426,N_44167);
nand U45779 (N_45779,N_41264,N_44881);
nand U45780 (N_45780,N_41382,N_42543);
nor U45781 (N_45781,N_42600,N_42498);
nand U45782 (N_45782,N_40070,N_42621);
or U45783 (N_45783,N_43738,N_44562);
xnor U45784 (N_45784,N_40197,N_43377);
and U45785 (N_45785,N_42436,N_40061);
and U45786 (N_45786,N_43644,N_43213);
and U45787 (N_45787,N_41364,N_40285);
or U45788 (N_45788,N_42377,N_40679);
and U45789 (N_45789,N_40896,N_41023);
or U45790 (N_45790,N_44702,N_40209);
nand U45791 (N_45791,N_42885,N_42273);
nor U45792 (N_45792,N_44277,N_44211);
and U45793 (N_45793,N_40749,N_43136);
nor U45794 (N_45794,N_42430,N_43633);
or U45795 (N_45795,N_43373,N_41931);
or U45796 (N_45796,N_43023,N_42675);
and U45797 (N_45797,N_42043,N_42381);
nor U45798 (N_45798,N_40366,N_41113);
or U45799 (N_45799,N_40256,N_41213);
nor U45800 (N_45800,N_42274,N_42844);
xnor U45801 (N_45801,N_43079,N_41308);
nand U45802 (N_45802,N_42821,N_43559);
or U45803 (N_45803,N_43078,N_41366);
nor U45804 (N_45804,N_40497,N_42530);
nand U45805 (N_45805,N_43463,N_40718);
and U45806 (N_45806,N_40225,N_42304);
nand U45807 (N_45807,N_43121,N_40433);
nor U45808 (N_45808,N_41174,N_44020);
nor U45809 (N_45809,N_42328,N_40743);
nor U45810 (N_45810,N_40853,N_42314);
nor U45811 (N_45811,N_44674,N_40954);
xnor U45812 (N_45812,N_44460,N_42419);
nor U45813 (N_45813,N_42573,N_41612);
nand U45814 (N_45814,N_43292,N_41844);
nand U45815 (N_45815,N_44863,N_43699);
and U45816 (N_45816,N_40716,N_42777);
nand U45817 (N_45817,N_40196,N_41656);
nand U45818 (N_45818,N_41795,N_41483);
nand U45819 (N_45819,N_43517,N_43563);
or U45820 (N_45820,N_44180,N_41581);
nor U45821 (N_45821,N_40249,N_44259);
xnor U45822 (N_45822,N_43673,N_40212);
and U45823 (N_45823,N_40404,N_43874);
nand U45824 (N_45824,N_40086,N_44465);
xor U45825 (N_45825,N_41576,N_43311);
nand U45826 (N_45826,N_43897,N_40044);
or U45827 (N_45827,N_40729,N_40605);
nor U45828 (N_45828,N_44639,N_40715);
nand U45829 (N_45829,N_43510,N_44380);
nor U45830 (N_45830,N_44161,N_42361);
xor U45831 (N_45831,N_41230,N_44884);
or U45832 (N_45832,N_41471,N_42564);
xnor U45833 (N_45833,N_41272,N_41122);
nor U45834 (N_45834,N_43401,N_42394);
or U45835 (N_45835,N_44324,N_43842);
and U45836 (N_45836,N_41964,N_43108);
nand U45837 (N_45837,N_44420,N_40769);
and U45838 (N_45838,N_43509,N_44610);
nor U45839 (N_45839,N_42987,N_43969);
and U45840 (N_45840,N_40858,N_41727);
nor U45841 (N_45841,N_43647,N_43287);
and U45842 (N_45842,N_40100,N_43704);
or U45843 (N_45843,N_40011,N_41035);
and U45844 (N_45844,N_40631,N_41661);
xnor U45845 (N_45845,N_43649,N_44123);
or U45846 (N_45846,N_42398,N_41249);
xor U45847 (N_45847,N_42785,N_42338);
or U45848 (N_45848,N_44318,N_43873);
nor U45849 (N_45849,N_40240,N_43919);
xnor U45850 (N_45850,N_43355,N_41751);
and U45851 (N_45851,N_41726,N_41918);
xor U45852 (N_45852,N_44162,N_42935);
or U45853 (N_45853,N_40657,N_42080);
nand U45854 (N_45854,N_41352,N_42289);
or U45855 (N_45855,N_42632,N_42981);
nand U45856 (N_45856,N_41083,N_40384);
nand U45857 (N_45857,N_44218,N_40870);
nor U45858 (N_45858,N_43710,N_40509);
nand U45859 (N_45859,N_40877,N_43902);
xnor U45860 (N_45860,N_42525,N_41208);
and U45861 (N_45861,N_41180,N_41854);
xnor U45862 (N_45862,N_41888,N_41131);
nor U45863 (N_45863,N_44852,N_43303);
nand U45864 (N_45864,N_41140,N_42252);
nor U45865 (N_45865,N_41069,N_40651);
or U45866 (N_45866,N_41418,N_42433);
or U45867 (N_45867,N_42315,N_43061);
or U45868 (N_45868,N_41025,N_42623);
nor U45869 (N_45869,N_41766,N_44855);
nor U45870 (N_45870,N_42386,N_44919);
xnor U45871 (N_45871,N_40175,N_41057);
xor U45872 (N_45872,N_40328,N_43894);
and U45873 (N_45873,N_41714,N_43683);
and U45874 (N_45874,N_41319,N_41954);
or U45875 (N_45875,N_42130,N_40126);
xnor U45876 (N_45876,N_43209,N_44155);
or U45877 (N_45877,N_44176,N_42871);
nand U45878 (N_45878,N_41857,N_44794);
xnor U45879 (N_45879,N_42175,N_40096);
nand U45880 (N_45880,N_44376,N_43711);
or U45881 (N_45881,N_43360,N_41925);
nor U45882 (N_45882,N_44478,N_40025);
or U45883 (N_45883,N_41098,N_44682);
or U45884 (N_45884,N_40157,N_44630);
nor U45885 (N_45885,N_42149,N_44334);
and U45886 (N_45886,N_44195,N_44238);
xnor U45887 (N_45887,N_43124,N_42636);
nor U45888 (N_45888,N_40019,N_40146);
or U45889 (N_45889,N_41583,N_41327);
or U45890 (N_45890,N_43005,N_40132);
or U45891 (N_45891,N_40153,N_41615);
nor U45892 (N_45892,N_43950,N_42111);
xnor U45893 (N_45893,N_43295,N_40862);
nor U45894 (N_45894,N_42959,N_44464);
or U45895 (N_45895,N_41395,N_42233);
xor U45896 (N_45896,N_40372,N_43082);
nand U45897 (N_45897,N_44808,N_43855);
nor U45898 (N_45898,N_42447,N_43498);
or U45899 (N_45899,N_43957,N_43378);
xor U45900 (N_45900,N_44285,N_40466);
or U45901 (N_45901,N_41387,N_44851);
xnor U45902 (N_45902,N_44725,N_40503);
or U45903 (N_45903,N_42897,N_43742);
and U45904 (N_45904,N_40827,N_41439);
and U45905 (N_45905,N_43586,N_42287);
nor U45906 (N_45906,N_44685,N_41186);
and U45907 (N_45907,N_42991,N_44109);
xnor U45908 (N_45908,N_41286,N_44351);
nor U45909 (N_45909,N_42609,N_41096);
xor U45910 (N_45910,N_44149,N_41620);
or U45911 (N_45911,N_40966,N_44146);
nand U45912 (N_45912,N_40236,N_43332);
nand U45913 (N_45913,N_42810,N_42647);
nand U45914 (N_45914,N_42967,N_43202);
or U45915 (N_45915,N_41881,N_43489);
nor U45916 (N_45916,N_44739,N_41594);
nor U45917 (N_45917,N_43587,N_42652);
nand U45918 (N_45918,N_41461,N_43551);
nand U45919 (N_45919,N_41111,N_44291);
nand U45920 (N_45920,N_40735,N_42512);
nand U45921 (N_45921,N_44723,N_42628);
xnor U45922 (N_45922,N_43441,N_42699);
nor U45923 (N_45923,N_41112,N_44722);
xor U45924 (N_45924,N_41819,N_43516);
or U45925 (N_45925,N_44014,N_43349);
nor U45926 (N_45926,N_44216,N_44021);
nand U45927 (N_45927,N_42679,N_40696);
xnor U45928 (N_45928,N_40111,N_41508);
or U45929 (N_45929,N_42417,N_44317);
nand U45930 (N_45930,N_43567,N_44691);
nand U45931 (N_45931,N_40340,N_41276);
xor U45932 (N_45932,N_42924,N_42820);
nand U45933 (N_45933,N_42356,N_43724);
nand U45934 (N_45934,N_44958,N_44737);
or U45935 (N_45935,N_40834,N_41043);
and U45936 (N_45936,N_43208,N_40210);
xor U45937 (N_45937,N_44382,N_41588);
xnor U45938 (N_45938,N_41095,N_43252);
nand U45939 (N_45939,N_40168,N_40461);
nor U45940 (N_45940,N_43884,N_44533);
nor U45941 (N_45941,N_40566,N_41636);
nand U45942 (N_45942,N_44107,N_40534);
nor U45943 (N_45943,N_41731,N_42845);
or U45944 (N_45944,N_40722,N_42876);
nand U45945 (N_45945,N_43425,N_42295);
xor U45946 (N_45946,N_44312,N_44503);
nor U45947 (N_45947,N_43685,N_40453);
or U45948 (N_45948,N_42446,N_40910);
or U45949 (N_45949,N_40583,N_40279);
or U45950 (N_45950,N_44689,N_41786);
xor U45951 (N_45951,N_42199,N_42120);
and U45952 (N_45952,N_43007,N_43707);
nor U45953 (N_45953,N_40643,N_42798);
nand U45954 (N_45954,N_43886,N_43073);
or U45955 (N_45955,N_42008,N_41356);
and U45956 (N_45956,N_44657,N_43507);
xor U45957 (N_45957,N_42290,N_41072);
nand U45958 (N_45958,N_42277,N_43863);
nand U45959 (N_45959,N_42238,N_40873);
or U45960 (N_45960,N_40504,N_41915);
nor U45961 (N_45961,N_42766,N_42757);
nor U45962 (N_45962,N_42028,N_42676);
or U45963 (N_45963,N_40049,N_44849);
xnor U45964 (N_45964,N_41771,N_42658);
nor U45965 (N_45965,N_44037,N_40151);
or U45966 (N_45966,N_44819,N_44879);
or U45967 (N_45967,N_41375,N_40617);
nand U45968 (N_45968,N_42168,N_42429);
nor U45969 (N_45969,N_40420,N_41392);
or U45970 (N_45970,N_43838,N_43695);
or U45971 (N_45971,N_43022,N_41758);
or U45972 (N_45972,N_42176,N_40944);
or U45973 (N_45973,N_43194,N_43175);
nor U45974 (N_45974,N_44429,N_43985);
xor U45975 (N_45975,N_43535,N_43766);
or U45976 (N_45976,N_44284,N_40137);
nor U45977 (N_45977,N_40211,N_44664);
nand U45978 (N_45978,N_41999,N_44777);
and U45979 (N_45979,N_41790,N_41401);
or U45980 (N_45980,N_40846,N_43096);
nor U45981 (N_45981,N_42938,N_41673);
or U45982 (N_45982,N_44774,N_43036);
xor U45983 (N_45983,N_40021,N_42578);
and U45984 (N_45984,N_41996,N_44581);
or U45985 (N_45985,N_42629,N_43994);
xor U45986 (N_45986,N_43501,N_42717);
nand U45987 (N_45987,N_40713,N_44219);
nand U45988 (N_45988,N_43908,N_41928);
or U45989 (N_45989,N_40190,N_42714);
and U45990 (N_45990,N_41933,N_44214);
xor U45991 (N_45991,N_43831,N_44448);
nand U45992 (N_45992,N_41913,N_42313);
or U45993 (N_45993,N_41490,N_44144);
and U45994 (N_45994,N_42202,N_41614);
xnor U45995 (N_45995,N_42716,N_42613);
nand U45996 (N_45996,N_40719,N_44821);
nand U45997 (N_45997,N_40922,N_42688);
nor U45998 (N_45998,N_44454,N_41963);
or U45999 (N_45999,N_43053,N_43154);
nand U46000 (N_46000,N_44992,N_43700);
and U46001 (N_46001,N_42918,N_40797);
nor U46002 (N_46002,N_41979,N_42502);
and U46003 (N_46003,N_44190,N_43952);
xnor U46004 (N_46004,N_41883,N_43084);
nand U46005 (N_46005,N_43339,N_43803);
nand U46006 (N_46006,N_42948,N_42517);
nand U46007 (N_46007,N_44687,N_44518);
nand U46008 (N_46008,N_41237,N_42953);
nor U46009 (N_46009,N_44026,N_44188);
or U46010 (N_46010,N_40218,N_44261);
or U46011 (N_46011,N_42309,N_44720);
or U46012 (N_46012,N_43185,N_42588);
nor U46013 (N_46013,N_40744,N_44869);
nor U46014 (N_46014,N_43891,N_40659);
and U46015 (N_46015,N_40610,N_41324);
or U46016 (N_46016,N_40104,N_40300);
and U46017 (N_46017,N_40089,N_42713);
xor U46018 (N_46018,N_43065,N_40233);
xnor U46019 (N_46019,N_41468,N_44583);
xor U46020 (N_46020,N_41523,N_44588);
xor U46021 (N_46021,N_42985,N_40405);
xor U46022 (N_46022,N_44866,N_42709);
and U46023 (N_46023,N_43678,N_41765);
or U46024 (N_46024,N_41344,N_41167);
or U46025 (N_46025,N_42232,N_44582);
xnor U46026 (N_46026,N_42301,N_41834);
xor U46027 (N_46027,N_42007,N_44024);
nor U46028 (N_46028,N_41882,N_41388);
or U46029 (N_46029,N_40627,N_44620);
and U46030 (N_46030,N_40465,N_41333);
or U46031 (N_46031,N_41895,N_41214);
nor U46032 (N_46032,N_41274,N_42753);
or U46033 (N_46033,N_41644,N_40034);
xor U46034 (N_46034,N_40514,N_42483);
or U46035 (N_46035,N_43783,N_43385);
and U46036 (N_46036,N_40419,N_44252);
xnor U46037 (N_46037,N_43230,N_43088);
xor U46038 (N_46038,N_42439,N_44978);
or U46039 (N_46039,N_43147,N_40513);
or U46040 (N_46040,N_41173,N_43634);
nand U46041 (N_46041,N_41146,N_43570);
xnor U46042 (N_46042,N_44160,N_42322);
nor U46043 (N_46043,N_44986,N_43257);
and U46044 (N_46044,N_43913,N_43126);
nand U46045 (N_46045,N_42702,N_40960);
nor U46046 (N_46046,N_42096,N_42670);
nor U46047 (N_46047,N_44544,N_41346);
nor U46048 (N_46048,N_43274,N_44705);
xnor U46049 (N_46049,N_40401,N_43316);
xor U46050 (N_46050,N_41580,N_44220);
xor U46051 (N_46051,N_44667,N_40934);
and U46052 (N_46052,N_43430,N_44660);
or U46053 (N_46053,N_41415,N_44244);
nor U46054 (N_46054,N_44437,N_41887);
nor U46055 (N_46055,N_41363,N_40721);
xor U46056 (N_46056,N_41399,N_44054);
and U46057 (N_46057,N_40048,N_42936);
xnor U46058 (N_46058,N_44419,N_43356);
nand U46059 (N_46059,N_42508,N_40268);
xnor U46060 (N_46060,N_44521,N_40930);
xor U46061 (N_46061,N_41241,N_40836);
xnor U46062 (N_46062,N_41426,N_40902);
xnor U46063 (N_46063,N_44332,N_42719);
xnor U46064 (N_46064,N_40764,N_41585);
nand U46065 (N_46065,N_40554,N_42974);
nor U46066 (N_46066,N_43953,N_44433);
and U46067 (N_46067,N_41037,N_42013);
nand U46068 (N_46068,N_43496,N_42006);
nand U46069 (N_46069,N_41489,N_40067);
nor U46070 (N_46070,N_43361,N_43272);
nand U46071 (N_46071,N_44957,N_43907);
nor U46072 (N_46072,N_42677,N_40010);
nor U46073 (N_46073,N_44729,N_44043);
nand U46074 (N_46074,N_42671,N_43847);
xor U46075 (N_46075,N_41200,N_41699);
xnor U46076 (N_46076,N_42423,N_43435);
xor U46077 (N_46077,N_41359,N_44289);
xnor U46078 (N_46078,N_42519,N_40814);
nand U46079 (N_46079,N_41940,N_42551);
xnor U46080 (N_46080,N_42451,N_42039);
or U46081 (N_46081,N_43705,N_41911);
nor U46082 (N_46082,N_43650,N_44056);
or U46083 (N_46083,N_42604,N_42253);
nor U46084 (N_46084,N_42216,N_41772);
or U46085 (N_46085,N_43593,N_41695);
or U46086 (N_46086,N_40138,N_44535);
and U46087 (N_46087,N_44245,N_40449);
nor U46088 (N_46088,N_44456,N_44036);
and U46089 (N_46089,N_40265,N_44985);
and U46090 (N_46090,N_44475,N_44928);
and U46091 (N_46091,N_40839,N_40826);
nor U46092 (N_46092,N_43153,N_43592);
or U46093 (N_46093,N_40030,N_43702);
or U46094 (N_46094,N_41080,N_41805);
or U46095 (N_46095,N_41802,N_42834);
and U46096 (N_46096,N_43348,N_43240);
nand U46097 (N_46097,N_44708,N_44741);
and U46098 (N_46098,N_42015,N_41407);
or U46099 (N_46099,N_44213,N_44557);
nor U46100 (N_46100,N_43653,N_42865);
or U46101 (N_46101,N_42217,N_43857);
nor U46102 (N_46102,N_41868,N_41548);
nand U46103 (N_46103,N_41460,N_43645);
and U46104 (N_46104,N_41796,N_40648);
and U46105 (N_46105,N_44035,N_44966);
xnor U46106 (N_46106,N_44359,N_42421);
or U46107 (N_46107,N_43905,N_43823);
nor U46108 (N_46108,N_40945,N_44933);
nor U46109 (N_46109,N_41845,N_40475);
nor U46110 (N_46110,N_40299,N_43347);
xor U46111 (N_46111,N_40341,N_41578);
and U46112 (N_46112,N_43546,N_41658);
and U46113 (N_46113,N_41647,N_41443);
nand U46114 (N_46114,N_40336,N_42258);
xnor U46115 (N_46115,N_43335,N_44840);
xor U46116 (N_46116,N_42271,N_42910);
nand U46117 (N_46117,N_40202,N_42250);
nand U46118 (N_46118,N_41216,N_42476);
or U46119 (N_46119,N_43663,N_42266);
or U46120 (N_46120,N_42663,N_42212);
nor U46121 (N_46121,N_40818,N_44595);
nand U46122 (N_46122,N_44524,N_41369);
nand U46123 (N_46123,N_43388,N_44551);
or U46124 (N_46124,N_44354,N_41028);
and U46125 (N_46125,N_43829,N_43034);
and U46126 (N_46126,N_40342,N_40075);
xor U46127 (N_46127,N_41902,N_44543);
xnor U46128 (N_46128,N_42895,N_42443);
nor U46129 (N_46129,N_44206,N_43172);
and U46130 (N_46130,N_42500,N_43032);
and U46131 (N_46131,N_41956,N_44746);
nor U46132 (N_46132,N_42755,N_40258);
xor U46133 (N_46133,N_41297,N_40685);
nand U46134 (N_46134,N_41884,N_40243);
or U46135 (N_46135,N_43849,N_41494);
or U46136 (N_46136,N_43666,N_42209);
xor U46137 (N_46137,N_42575,N_44931);
nand U46138 (N_46138,N_40289,N_40727);
nor U46139 (N_46139,N_43569,N_43602);
or U46140 (N_46140,N_44041,N_42861);
nand U46141 (N_46141,N_40281,N_44509);
and U46142 (N_46142,N_40868,N_40382);
and U46143 (N_46143,N_42403,N_40237);
nor U46144 (N_46144,N_43719,N_40615);
xor U46145 (N_46145,N_43538,N_41328);
nor U46146 (N_46146,N_40428,N_42772);
or U46147 (N_46147,N_40105,N_43226);
nor U46148 (N_46148,N_41801,N_41740);
and U46149 (N_46149,N_43341,N_41735);
or U46150 (N_46150,N_43794,N_44207);
nor U46151 (N_46151,N_40078,N_43895);
nor U46152 (N_46152,N_43146,N_44085);
xor U46153 (N_46153,N_44340,N_44690);
nor U46154 (N_46154,N_44121,N_41730);
and U46155 (N_46155,N_41434,N_42320);
nand U46156 (N_46156,N_43162,N_44292);
and U46157 (N_46157,N_42538,N_44431);
xor U46158 (N_46158,N_40161,N_41222);
xnor U46159 (N_46159,N_43229,N_44644);
nor U46160 (N_46160,N_41198,N_43777);
or U46161 (N_46161,N_44022,N_42321);
and U46162 (N_46162,N_41233,N_44168);
nand U46163 (N_46163,N_43416,N_44100);
nor U46164 (N_46164,N_41330,N_43149);
nor U46165 (N_46165,N_41485,N_41600);
xor U46166 (N_46166,N_40380,N_41182);
xnor U46167 (N_46167,N_40085,N_42325);
xnor U46168 (N_46168,N_44232,N_44426);
or U46169 (N_46169,N_44398,N_40412);
nor U46170 (N_46170,N_44609,N_41440);
xor U46171 (N_46171,N_41825,N_44990);
nor U46172 (N_46172,N_43859,N_40609);
and U46173 (N_46173,N_43246,N_42904);
nor U46174 (N_46174,N_40712,N_44699);
nor U46175 (N_46175,N_40516,N_43762);
nand U46176 (N_46176,N_43931,N_44982);
xor U46177 (N_46177,N_40684,N_42059);
nand U46178 (N_46178,N_42173,N_44530);
nand U46179 (N_46179,N_42269,N_43090);
and U46180 (N_46180,N_43122,N_44192);
or U46181 (N_46181,N_42979,N_43576);
xnor U46182 (N_46182,N_41189,N_42555);
nand U46183 (N_46183,N_42988,N_43403);
xor U46184 (N_46184,N_41718,N_41143);
or U46185 (N_46185,N_43315,N_40351);
nand U46186 (N_46186,N_43521,N_44116);
nand U46187 (N_46187,N_44067,N_43116);
nor U46188 (N_46188,N_40611,N_43402);
xor U46189 (N_46189,N_42415,N_42383);
and U46190 (N_46190,N_41569,N_41889);
nand U46191 (N_46191,N_43075,N_43371);
or U46192 (N_46192,N_41760,N_41019);
xnor U46193 (N_46193,N_40674,N_40755);
nand U46194 (N_46194,N_41713,N_44302);
xnor U46195 (N_46195,N_43772,N_44596);
nor U46196 (N_46196,N_43970,N_41042);
xor U46197 (N_46197,N_43582,N_42639);
and U46198 (N_46198,N_41081,N_42635);
nor U46199 (N_46199,N_42189,N_41917);
or U46200 (N_46200,N_42599,N_42256);
xnor U46201 (N_46201,N_42620,N_42654);
nand U46202 (N_46202,N_40261,N_40170);
nand U46203 (N_46203,N_44440,N_40326);
xor U46204 (N_46204,N_43625,N_40600);
or U46205 (N_46205,N_40192,N_44904);
xnor U46206 (N_46206,N_44196,N_44711);
and U46207 (N_46207,N_40660,N_43471);
or U46208 (N_46208,N_40367,N_41769);
xor U46209 (N_46209,N_43714,N_44764);
xnor U46210 (N_46210,N_40417,N_40900);
and U46211 (N_46211,N_41150,N_40053);
or U46212 (N_46212,N_44233,N_42706);
or U46213 (N_46213,N_40345,N_42586);
nand U46214 (N_46214,N_44975,N_40913);
and U46215 (N_46215,N_44580,N_44824);
and U46216 (N_46216,N_41488,N_43541);
and U46217 (N_46217,N_44798,N_44221);
or U46218 (N_46218,N_43359,N_40110);
nand U46219 (N_46219,N_43485,N_43750);
or U46220 (N_46220,N_41711,N_43427);
nand U46221 (N_46221,N_42427,N_42197);
xnor U46222 (N_46222,N_41141,N_41291);
nand U46223 (N_46223,N_43961,N_41102);
xnor U46224 (N_46224,N_41547,N_40165);
xnor U46225 (N_46225,N_43887,N_44984);
or U46226 (N_46226,N_41267,N_40664);
and U46227 (N_46227,N_43177,N_41012);
nor U46228 (N_46228,N_43899,N_41634);
and U46229 (N_46229,N_43070,N_42666);
nand U46230 (N_46230,N_43579,N_40295);
or U46231 (N_46231,N_41534,N_43404);
nand U46232 (N_46232,N_40090,N_41935);
nor U46233 (N_46233,N_41574,N_44338);
nand U46234 (N_46234,N_41243,N_42019);
nand U46235 (N_46235,N_41524,N_41685);
xnor U46236 (N_46236,N_40106,N_44563);
xor U46237 (N_46237,N_40953,N_43173);
nor U46238 (N_46238,N_44724,N_40221);
and U46239 (N_46239,N_43000,N_44505);
and U46240 (N_46240,N_42667,N_44362);
xnor U46241 (N_46241,N_42796,N_40012);
or U46242 (N_46242,N_41543,N_42887);
nor U46243 (N_46243,N_41021,N_40304);
nor U46244 (N_46244,N_41942,N_41207);
or U46245 (N_46245,N_41599,N_43978);
xnor U46246 (N_46246,N_40040,N_43343);
xor U46247 (N_46247,N_44716,N_40358);
nand U46248 (N_46248,N_42703,N_44659);
or U46249 (N_46249,N_40144,N_42992);
xnor U46250 (N_46250,N_42933,N_44117);
nand U46251 (N_46251,N_42192,N_40361);
and U46252 (N_46252,N_43752,N_44556);
nand U46253 (N_46253,N_41794,N_43216);
xor U46254 (N_46254,N_42191,N_40282);
or U46255 (N_46255,N_41250,N_41871);
nor U46256 (N_46256,N_44761,N_40803);
or U46257 (N_46257,N_43397,N_43580);
xnor U46258 (N_46258,N_41051,N_40098);
and U46259 (N_46259,N_40562,N_42300);
nor U46260 (N_46260,N_41690,N_43399);
and U46261 (N_46261,N_41444,N_40041);
xnor U46262 (N_46262,N_43915,N_42559);
nor U46263 (N_46263,N_44344,N_41556);
or U46264 (N_46264,N_41292,N_44692);
xor U46265 (N_46265,N_42989,N_44909);
nand U46266 (N_46266,N_42546,N_44950);
nor U46267 (N_46267,N_40224,N_42826);
or U46268 (N_46268,N_41000,N_40148);
nand U46269 (N_46269,N_42422,N_44126);
nand U46270 (N_46270,N_42352,N_40525);
or U46271 (N_46271,N_44488,N_40317);
nor U46272 (N_46272,N_43984,N_43944);
xor U46273 (N_46273,N_42399,N_43475);
and U46274 (N_46274,N_42715,N_40936);
or U46275 (N_46275,N_42583,N_41393);
nand U46276 (N_46276,N_40492,N_43814);
nor U46277 (N_46277,N_41464,N_44999);
nand U46278 (N_46278,N_44293,N_41906);
and U46279 (N_46279,N_41721,N_41217);
nor U46280 (N_46280,N_40169,N_42094);
or U46281 (N_46281,N_42863,N_40005);
nor U46282 (N_46282,N_42126,N_43937);
nor U46283 (N_46283,N_43659,N_42060);
and U46284 (N_46284,N_40544,N_41551);
and U46285 (N_46285,N_40575,N_44375);
and U46286 (N_46286,N_43827,N_43015);
and U46287 (N_46287,N_41255,N_40125);
and U46288 (N_46288,N_41676,N_43619);
and U46289 (N_46289,N_44323,N_40758);
nand U46290 (N_46290,N_40951,N_40519);
xnor U46291 (N_46291,N_42929,N_40784);
or U46292 (N_46292,N_41807,N_40931);
nor U46293 (N_46293,N_41851,N_42520);
or U46294 (N_46294,N_41298,N_43220);
nor U46295 (N_46295,N_43305,N_41830);
or U46296 (N_46296,N_41296,N_42005);
or U46297 (N_46297,N_42972,N_41431);
nand U46298 (N_46298,N_42117,N_42941);
xnor U46299 (N_46299,N_44814,N_40535);
and U46300 (N_46300,N_44201,N_41848);
and U46301 (N_46301,N_40542,N_40028);
and U46302 (N_46302,N_40667,N_44333);
xnor U46303 (N_46303,N_43934,N_42184);
nor U46304 (N_46304,N_44139,N_42363);
and U46305 (N_46305,N_40072,N_43718);
or U46306 (N_46306,N_41185,N_40343);
xnor U46307 (N_46307,N_43134,N_43464);
nand U46308 (N_46308,N_40903,N_42947);
nor U46309 (N_46309,N_42641,N_44011);
nand U46310 (N_46310,N_44662,N_42814);
and U46311 (N_46311,N_40039,N_44943);
and U46312 (N_46312,N_43925,N_42683);
nand U46313 (N_46313,N_41007,N_43334);
or U46314 (N_46314,N_44256,N_40840);
xnor U46315 (N_46315,N_41336,N_40832);
nor U46316 (N_46316,N_44477,N_43565);
or U46317 (N_46317,N_43042,N_43712);
nand U46318 (N_46318,N_44531,N_41838);
or U46319 (N_46319,N_40076,N_42595);
nand U46320 (N_46320,N_41435,N_42695);
xnor U46321 (N_46321,N_43995,N_40043);
nand U46322 (N_46322,N_40738,N_44019);
nand U46323 (N_46323,N_41045,N_40352);
or U46324 (N_46324,N_44061,N_43462);
and U46325 (N_46325,N_41505,N_40695);
xor U46326 (N_46326,N_44257,N_40622);
nand U46327 (N_46327,N_44243,N_42086);
or U46328 (N_46328,N_40927,N_42453);
or U46329 (N_46329,N_41662,N_43181);
nor U46330 (N_46330,N_44962,N_44668);
and U46331 (N_46331,N_40760,N_42542);
and U46332 (N_46332,N_44565,N_43447);
nor U46333 (N_46333,N_40073,N_44864);
nor U46334 (N_46334,N_40199,N_44430);
xor U46335 (N_46335,N_41337,N_42098);
nor U46336 (N_46336,N_41638,N_44898);
xor U46337 (N_46337,N_44893,N_44770);
nand U46338 (N_46338,N_40219,N_43872);
and U46339 (N_46339,N_40029,N_43263);
nor U46340 (N_46340,N_40968,N_44199);
and U46341 (N_46341,N_43214,N_40899);
nor U46342 (N_46342,N_41946,N_41191);
or U46343 (N_46343,N_44584,N_42109);
and U46344 (N_46344,N_44930,N_42465);
xnor U46345 (N_46345,N_42225,N_44835);
xor U46346 (N_46346,N_40128,N_44462);
nor U46347 (N_46347,N_44345,N_42179);
or U46348 (N_46348,N_42046,N_44187);
nor U46349 (N_46349,N_43280,N_43962);
nor U46350 (N_46350,N_42261,N_44391);
or U46351 (N_46351,N_40483,N_43417);
and U46352 (N_46352,N_43491,N_43443);
and U46353 (N_46353,N_41767,N_44276);
or U46354 (N_46354,N_42550,N_44385);
nand U46355 (N_46355,N_40446,N_44679);
or U46356 (N_46356,N_44205,N_44495);
nor U46357 (N_46357,N_43419,N_44390);
nand U46358 (N_46358,N_42090,N_44106);
or U46359 (N_46359,N_43583,N_44707);
nor U46360 (N_46360,N_42721,N_43423);
nor U46361 (N_46361,N_41774,N_42157);
nor U46362 (N_46362,N_41839,N_40093);
nand U46363 (N_46363,N_40244,N_44033);
nand U46364 (N_46364,N_44173,N_41694);
and U46365 (N_46365,N_42759,N_44946);
xnor U46366 (N_46366,N_41462,N_44998);
xnor U46367 (N_46367,N_41209,N_43561);
xor U46368 (N_46368,N_40275,N_44066);
nand U46369 (N_46369,N_44677,N_41073);
nor U46370 (N_46370,N_41284,N_42957);
nor U46371 (N_46371,N_41880,N_40101);
xnor U46372 (N_46372,N_41287,N_42608);
and U46373 (N_46373,N_44446,N_40699);
or U46374 (N_46374,N_44008,N_44676);
and U46375 (N_46375,N_40977,N_40394);
or U46376 (N_46376,N_42215,N_40981);
and U46377 (N_46377,N_42420,N_44751);
or U46378 (N_46378,N_41269,N_42685);
nor U46379 (N_46379,N_41194,N_41153);
nand U46380 (N_46380,N_43318,N_40332);
or U46381 (N_46381,N_42754,N_44995);
nor U46382 (N_46382,N_40672,N_40889);
or U46383 (N_46383,N_40473,N_42237);
nand U46384 (N_46384,N_44124,N_41677);
or U46385 (N_46385,N_41156,N_44305);
or U46386 (N_46386,N_43351,N_43534);
or U46387 (N_46387,N_44783,N_42828);
nand U46388 (N_46388,N_43648,N_41066);
xnor U46389 (N_46389,N_42723,N_44327);
and U46390 (N_46390,N_42975,N_44651);
xnor U46391 (N_46391,N_44771,N_40178);
or U46392 (N_46392,N_42875,N_42357);
and U46393 (N_46393,N_43253,N_42291);
xnor U46394 (N_46394,N_40885,N_44646);
nand U46395 (N_46395,N_41894,N_40823);
or U46396 (N_46396,N_42877,N_40650);
or U46397 (N_46397,N_43759,N_40884);
nand U46398 (N_46398,N_40756,N_41729);
nor U46399 (N_46399,N_40571,N_42589);
or U46400 (N_46400,N_40775,N_44567);
or U46401 (N_46401,N_42902,N_44972);
and U46402 (N_46402,N_41301,N_44843);
or U46403 (N_46403,N_40499,N_41978);
nand U46404 (N_46404,N_44336,N_42218);
and U46405 (N_46405,N_40103,N_43245);
nor U46406 (N_46406,N_40967,N_40369);
and U46407 (N_46407,N_43802,N_40472);
or U46408 (N_46408,N_43163,N_41598);
nand U46409 (N_46409,N_40139,N_44779);
and U46410 (N_46410,N_41316,N_42461);
and U46411 (N_46411,N_44260,N_44858);
nand U46412 (N_46412,N_43472,N_42343);
xnor U46413 (N_46413,N_42784,N_43191);
xor U46414 (N_46414,N_44272,N_42872);
and U46415 (N_46415,N_41526,N_40172);
or U46416 (N_46416,N_40559,N_40174);
nor U46417 (N_46417,N_44224,N_41860);
nor U46418 (N_46418,N_42342,N_42170);
or U46419 (N_46419,N_40855,N_40395);
or U46420 (N_46420,N_42018,N_42523);
nand U46421 (N_46421,N_40895,N_44829);
or U46422 (N_46422,N_40051,N_43434);
or U46423 (N_46423,N_44540,N_43598);
or U46424 (N_46424,N_43389,N_42016);
xnor U46425 (N_46425,N_44603,N_40898);
and U46426 (N_46426,N_42934,N_44486);
xor U46427 (N_46427,N_43609,N_41693);
and U46428 (N_46428,N_44948,N_40893);
xor U46429 (N_46429,N_40874,N_44894);
xnor U46430 (N_46430,N_41746,N_40223);
nor U46431 (N_46431,N_42646,N_42668);
nand U46432 (N_46432,N_40294,N_41257);
or U46433 (N_46433,N_43820,N_43066);
nand U46434 (N_46434,N_43935,N_40690);
and U46435 (N_46435,N_43207,N_41071);
nand U46436 (N_46436,N_42311,N_42645);
nand U46437 (N_46437,N_41827,N_40002);
and U46438 (N_46438,N_40331,N_44575);
xnor U46439 (N_46439,N_44718,N_42705);
nor U46440 (N_46440,N_41967,N_44920);
and U46441 (N_46441,N_41696,N_41481);
nor U46442 (N_46442,N_42596,N_44830);
xnor U46443 (N_46443,N_43026,N_44131);
and U46444 (N_46444,N_40723,N_44728);
xnor U46445 (N_46445,N_40505,N_42382);
nand U46446 (N_46446,N_40697,N_44063);
nand U46447 (N_46447,N_40928,N_40669);
xnor U46448 (N_46448,N_43622,N_44447);
nor U46449 (N_46449,N_42587,N_40238);
and U46450 (N_46450,N_41339,N_44355);
nor U46451 (N_46451,N_44346,N_42642);
nand U46452 (N_46452,N_44591,N_42655);
nor U46453 (N_46453,N_41567,N_40800);
nor U46454 (N_46454,N_43983,N_43545);
and U46455 (N_46455,N_43383,N_42597);
nand U46456 (N_46456,N_41853,N_42133);
nand U46457 (N_46457,N_43776,N_43715);
nor U46458 (N_46458,N_43030,N_40767);
nand U46459 (N_46459,N_43893,N_40360);
or U46460 (N_46460,N_43716,N_42418);
and U46461 (N_46461,N_40359,N_42284);
xnor U46462 (N_46462,N_40939,N_40042);
nor U46463 (N_46463,N_43429,N_43726);
xnor U46464 (N_46464,N_41728,N_40296);
and U46465 (N_46465,N_41867,N_40594);
or U46466 (N_46466,N_42172,N_42567);
xor U46467 (N_46467,N_42961,N_42730);
xnor U46468 (N_46468,N_44287,N_44142);
nand U46469 (N_46469,N_42649,N_41335);
and U46470 (N_46470,N_42344,N_41655);
nand U46471 (N_46471,N_42886,N_41381);
or U46472 (N_46472,N_42187,N_43658);
or U46473 (N_46473,N_42548,N_43708);
and U46474 (N_46474,N_44598,N_40905);
nor U46475 (N_46475,N_43482,N_43967);
nand U46476 (N_46476,N_40055,N_42186);
nor U46477 (N_46477,N_42206,N_41280);
xnor U46478 (N_46478,N_40553,N_41587);
or U46479 (N_46479,N_40689,N_44785);
or U46480 (N_46480,N_44358,N_41510);
nor U46481 (N_46481,N_41161,N_44547);
nand U46482 (N_46482,N_43959,N_42576);
or U46483 (N_46483,N_44652,N_40411);
xnor U46484 (N_46484,N_43279,N_43069);
nand U46485 (N_46485,N_43652,N_43796);
nor U46486 (N_46486,N_44402,N_41077);
xor U46487 (N_46487,N_40201,N_44719);
xor U46488 (N_46488,N_41438,N_42797);
and U46489 (N_46489,N_40095,N_43309);
xnor U46490 (N_46490,N_44805,N_44157);
xnor U46491 (N_46491,N_42438,N_41540);
xor U46492 (N_46492,N_42735,N_42118);
and U46493 (N_46493,N_40590,N_43686);
nor U46494 (N_46494,N_41637,N_42490);
xnor U46495 (N_46495,N_42779,N_41998);
or U46496 (N_46496,N_40830,N_40251);
nand U46497 (N_46497,N_44846,N_41338);
nand U46498 (N_46498,N_44499,N_44200);
and U46499 (N_46499,N_41736,N_41517);
nor U46500 (N_46500,N_42178,N_44278);
or U46501 (N_46501,N_44970,N_44316);
and U46502 (N_46502,N_44635,N_43885);
nand U46503 (N_46503,N_40478,N_41646);
nand U46504 (N_46504,N_43486,N_44427);
or U46505 (N_46505,N_44059,N_42104);
nor U46506 (N_46506,N_44599,N_40813);
xor U46507 (N_46507,N_44088,N_41897);
or U46508 (N_46508,N_40988,N_41265);
or U46509 (N_46509,N_43597,N_42724);
nor U46510 (N_46510,N_41305,N_43577);
xnor U46511 (N_46511,N_43260,N_40714);
nor U46512 (N_46512,N_41768,N_41118);
or U46513 (N_46513,N_41349,N_40292);
nand U46514 (N_46514,N_44096,N_42378);
nand U46515 (N_46515,N_44320,N_44586);
and U46516 (N_46516,N_44654,N_41202);
or U46517 (N_46517,N_40408,N_43732);
xnor U46518 (N_46518,N_43660,N_41820);
xnor U46519 (N_46519,N_40720,N_40467);
xor U46520 (N_46520,N_44282,N_40230);
xnor U46521 (N_46521,N_44680,N_43438);
and U46522 (N_46522,N_40603,N_43321);
nor U46523 (N_46523,N_41789,N_44401);
xor U46524 (N_46524,N_41107,N_42329);
nor U46525 (N_46525,N_43068,N_44759);
nor U46526 (N_46526,N_43291,N_44669);
nor U46527 (N_46527,N_42244,N_43151);
nand U46528 (N_46528,N_43693,N_40014);
and U46529 (N_46529,N_41263,N_42332);
nor U46530 (N_46530,N_43342,N_41067);
nor U46531 (N_46531,N_44444,N_44084);
and U46532 (N_46532,N_42219,N_43013);
nand U46533 (N_46533,N_41503,N_41148);
nor U46534 (N_46534,N_43865,N_44923);
nand U46535 (N_46535,N_42385,N_41062);
or U46536 (N_46536,N_44553,N_44979);
xor U46537 (N_46537,N_43882,N_44523);
or U46538 (N_46538,N_43560,N_42920);
or U46539 (N_46539,N_41553,N_42335);
nand U46540 (N_46540,N_40861,N_40567);
or U46541 (N_46541,N_41675,N_41824);
and U46542 (N_46542,N_42414,N_40923);
nand U46543 (N_46543,N_44573,N_43630);
nor U46544 (N_46544,N_41993,N_42908);
xor U46545 (N_46545,N_40363,N_41183);
nand U46546 (N_46546,N_43426,N_40871);
or U46547 (N_46547,N_40063,N_40843);
and U46548 (N_46548,N_42544,N_43613);
or U46549 (N_46549,N_42682,N_41376);
or U46550 (N_46550,N_41499,N_40587);
nand U46551 (N_46551,N_42262,N_42065);
and U46552 (N_46552,N_40231,N_44629);
nor U46553 (N_46553,N_43325,N_42428);
nor U46554 (N_46554,N_42511,N_42148);
or U46555 (N_46555,N_41509,N_42299);
and U46556 (N_46556,N_40570,N_40079);
nor U46557 (N_46557,N_40415,N_41742);
nand U46558 (N_46558,N_40311,N_42962);
xnor U46559 (N_46559,N_41855,N_44416);
nand U46560 (N_46560,N_42474,N_40838);
or U46561 (N_46561,N_44098,N_42795);
or U46562 (N_46562,N_40182,N_44817);
or U46563 (N_46563,N_44105,N_40272);
and U46564 (N_46564,N_40035,N_40470);
nor U46565 (N_46565,N_43608,N_42207);
or U46566 (N_46566,N_43028,N_44103);
or U46567 (N_46567,N_41983,N_44896);
nand U46568 (N_46568,N_42061,N_40957);
nor U46569 (N_46569,N_43187,N_43600);
xnor U46570 (N_46570,N_41374,N_42770);
xor U46571 (N_46571,N_44092,N_44449);
nand U46572 (N_46572,N_43304,N_42137);
or U46573 (N_46573,N_40305,N_42278);
and U46574 (N_46574,N_41597,N_41149);
nor U46575 (N_46575,N_42610,N_43249);
nand U46576 (N_46576,N_44064,N_43832);
nor U46577 (N_46577,N_40847,N_44423);
nand U46578 (N_46578,N_42969,N_42898);
nor U46579 (N_46579,N_40686,N_40578);
nor U46580 (N_46580,N_41228,N_40848);
xor U46581 (N_46581,N_42849,N_43159);
nand U46582 (N_46582,N_41919,N_44313);
and U46583 (N_46583,N_43095,N_44236);
nor U46584 (N_46584,N_41064,N_44490);
xnor U46585 (N_46585,N_40890,N_41896);
nor U46586 (N_46586,N_44752,N_43168);
and U46587 (N_46587,N_41748,N_40271);
nand U46588 (N_46588,N_40330,N_41788);
nor U46589 (N_46589,N_40545,N_40274);
nor U46590 (N_46590,N_41784,N_41893);
and U46591 (N_46591,N_42638,N_40640);
and U46592 (N_46592,N_42864,N_44590);
nor U46593 (N_46593,N_42116,N_43085);
nand U46594 (N_46594,N_41541,N_42580);
xor U46595 (N_46595,N_40979,N_44288);
nand U46596 (N_46596,N_44571,N_40973);
or U46597 (N_46597,N_42549,N_43812);
and U46598 (N_46598,N_40457,N_44976);
nor U46599 (N_46599,N_41278,N_40455);
and U46600 (N_46600,N_43270,N_41092);
and U46601 (N_46601,N_43696,N_44476);
nor U46602 (N_46602,N_41544,N_41591);
nand U46603 (N_46603,N_40410,N_44110);
nand U46604 (N_46604,N_42330,N_41109);
nor U46605 (N_46605,N_42637,N_43393);
nand U46606 (N_46606,N_40306,N_42774);
or U46607 (N_46607,N_40507,N_40164);
or U46608 (N_46608,N_43483,N_41501);
xor U46609 (N_46609,N_41652,N_44713);
and U46610 (N_46610,N_40123,N_44127);
xor U46611 (N_46611,N_43469,N_42088);
xor U46612 (N_46612,N_41238,N_40140);
xnor U46613 (N_46613,N_44996,N_42884);
nor U46614 (N_46614,N_43099,N_41126);
xor U46615 (N_46615,N_41659,N_43457);
xnor U46616 (N_46616,N_44023,N_44519);
nor U46617 (N_46617,N_42741,N_41031);
xor U46618 (N_46618,N_41229,N_44383);
and U46619 (N_46619,N_40257,N_40468);
or U46620 (N_46620,N_42602,N_42556);
or U46621 (N_46621,N_41242,N_41823);
or U46622 (N_46622,N_43684,N_42673);
nor U46623 (N_46623,N_44576,N_44671);
xnor U46624 (N_46624,N_40120,N_42319);
nand U46625 (N_46625,N_41679,N_43262);
and U46626 (N_46626,N_40837,N_44952);
nand U46627 (N_46627,N_40191,N_41804);
xor U46628 (N_46628,N_43590,N_43921);
nand U46629 (N_46629,N_40886,N_41630);
nand U46630 (N_46630,N_43142,N_40607);
xnor U46631 (N_46631,N_41937,N_41985);
nor U46632 (N_46632,N_43526,N_41921);
or U46633 (N_46633,N_44683,N_43468);
and U46634 (N_46634,N_43196,N_43878);
nor U46635 (N_46635,N_44527,N_44566);
xnor U46636 (N_46636,N_44784,N_42144);
xnor U46637 (N_46637,N_40576,N_43143);
nor U46638 (N_46638,N_41798,N_41780);
nor U46639 (N_46639,N_40438,N_42727);
or U46640 (N_46640,N_44373,N_41409);
xnor U46641 (N_46641,N_44539,N_41437);
nand U46642 (N_46642,N_40013,N_44251);
xor U46643 (N_46643,N_40811,N_43357);
or U46644 (N_46644,N_43029,N_41486);
and U46645 (N_46645,N_41936,N_43081);
nand U46646 (N_46646,N_42722,N_44701);
nor U46647 (N_46647,N_40392,N_41849);
and U46648 (N_46648,N_43484,N_43682);
xor U46649 (N_46649,N_40969,N_42899);
nor U46650 (N_46650,N_40347,N_43156);
xor U46651 (N_46651,N_44053,N_40581);
or U46652 (N_46652,N_41992,N_41390);
or U46653 (N_46653,N_41357,N_44714);
nand U46654 (N_46654,N_44263,N_40635);
xor U46655 (N_46655,N_42011,N_40849);
nor U46656 (N_46656,N_42971,N_42815);
and U46657 (N_46657,N_40628,N_43739);
nor U46658 (N_46658,N_44974,N_43605);
xor U46659 (N_46659,N_41421,N_41528);
xnor U46660 (N_46660,N_40494,N_44890);
nor U46661 (N_46661,N_44070,N_42407);
nor U46662 (N_46662,N_44897,N_43052);
nand U46663 (N_46663,N_41320,N_44377);
or U46664 (N_46664,N_43112,N_41188);
nor U46665 (N_46665,N_41050,N_42813);
nand U46666 (N_46666,N_44653,N_41251);
xor U46667 (N_46667,N_43193,N_41380);
and U46668 (N_46668,N_42499,N_43231);
nand U46669 (N_46669,N_42341,N_41762);
nor U46670 (N_46670,N_44108,N_43618);
nor U46671 (N_46671,N_44128,N_42832);
or U46672 (N_46672,N_41943,N_40996);
nand U46673 (N_46673,N_43350,N_42174);
xor U46674 (N_46674,N_41957,N_41816);
or U46675 (N_46675,N_44612,N_44271);
nand U46676 (N_46676,N_43848,N_41706);
xnor U46677 (N_46677,N_41417,N_41738);
and U46678 (N_46678,N_40613,N_40687);
and U46679 (N_46679,N_44057,N_41445);
nand U46680 (N_46680,N_42044,N_42803);
nand U46681 (N_46681,N_41672,N_40563);
xnor U46682 (N_46682,N_42083,N_40026);
nor U46683 (N_46683,N_41648,N_41075);
xnor U46684 (N_46684,N_43406,N_40993);
or U46685 (N_46685,N_40162,N_43864);
or U46686 (N_46686,N_42749,N_43637);
and U46687 (N_46687,N_44717,N_43821);
or U46688 (N_46688,N_40752,N_40865);
nand U46689 (N_46689,N_43384,N_44939);
xnor U46690 (N_46690,N_43301,N_44115);
nand U46691 (N_46691,N_41832,N_42978);
xor U46692 (N_46692,N_42995,N_43255);
or U46693 (N_46693,N_42532,N_44570);
nand U46694 (N_46694,N_42467,N_43988);
or U46695 (N_46695,N_42527,N_41926);
nand U46696 (N_46696,N_44228,N_43449);
nor U46697 (N_46697,N_41875,N_43680);
nand U46698 (N_46698,N_43345,N_42424);
nor U46699 (N_46699,N_42704,N_41026);
nor U46700 (N_46700,N_43019,N_42593);
and U46701 (N_46701,N_42152,N_44118);
or U46702 (N_46702,N_41219,N_44322);
or U46703 (N_46703,N_41922,N_40407);
nor U46704 (N_46704,N_42827,N_42454);
nand U46705 (N_46705,N_40348,N_43689);
xor U46706 (N_46706,N_42230,N_42119);
xor U46707 (N_46707,N_44525,N_44938);
or U46708 (N_46708,N_41960,N_42954);
and U46709 (N_46709,N_43221,N_42846);
xor U46710 (N_46710,N_42002,N_43076);
or U46711 (N_46711,N_41934,N_42648);
nor U46712 (N_46712,N_44296,N_44616);
and U46713 (N_46713,N_41649,N_40804);
and U46714 (N_46714,N_41617,N_41456);
or U46715 (N_46715,N_44031,N_43446);
nor U46716 (N_46716,N_43055,N_42360);
or U46717 (N_46717,N_40447,N_41060);
or U46718 (N_46718,N_42288,N_44695);
nor U46719 (N_46719,N_40964,N_41184);
and U46720 (N_46720,N_43322,N_42911);
and U46721 (N_46721,N_44082,N_41136);
and U46722 (N_46722,N_44917,N_42888);
nand U46723 (N_46723,N_40564,N_42468);
or U46724 (N_46724,N_43058,N_42047);
xnor U46725 (N_46725,N_42919,N_40250);
xor U46726 (N_46726,N_42455,N_43654);
nand U46727 (N_46727,N_43553,N_42449);
or U46728 (N_46728,N_43667,N_41258);
and U46729 (N_46729,N_40791,N_41030);
and U46730 (N_46730,N_41952,N_43797);
nor U46731 (N_46731,N_43171,N_40493);
or U46732 (N_46732,N_44832,N_44534);
and U46733 (N_46733,N_41293,N_43051);
or U46734 (N_46734,N_44081,N_44246);
or U46735 (N_46735,N_42850,N_40156);
nand U46736 (N_46736,N_41463,N_42883);
nor U46737 (N_46737,N_41231,N_41939);
nand U46738 (N_46738,N_43529,N_44922);
xor U46739 (N_46739,N_40794,N_43999);
and U46740 (N_46740,N_43722,N_44541);
nand U46741 (N_46741,N_43283,N_44605);
or U46742 (N_46742,N_42747,N_40589);
or U46743 (N_46743,N_42528,N_42584);
or U46744 (N_46744,N_44367,N_43391);
nor U46745 (N_46745,N_41433,N_43293);
nand U46746 (N_46746,N_40502,N_40409);
nand U46747 (N_46747,N_42210,N_43107);
and U46748 (N_46748,N_40935,N_44017);
xnor U46749 (N_46749,N_42125,N_42963);
nor U46750 (N_46750,N_41448,N_41476);
xnor U46751 (N_46751,N_40879,N_41847);
xnor U46752 (N_46752,N_43286,N_40016);
and U46753 (N_46753,N_40531,N_43433);
or U46754 (N_46754,N_44908,N_44468);
and U46755 (N_46755,N_43093,N_42965);
xnor U46756 (N_46756,N_40851,N_42413);
nand U46757 (N_46757,N_44177,N_41220);
xnor U46758 (N_46758,N_44513,N_41966);
and U46759 (N_46759,N_41701,N_41047);
and U46760 (N_46760,N_40812,N_42147);
and U46761 (N_46761,N_41905,N_42860);
nor U46762 (N_46762,N_43599,N_40441);
nand U46763 (N_46763,N_44378,N_42848);
nand U46764 (N_46764,N_42914,N_43770);
xor U46765 (N_46765,N_41633,N_41322);
and U46766 (N_46766,N_44120,N_42303);
and U46767 (N_46767,N_40400,N_41119);
nor U46768 (N_46768,N_42012,N_41175);
and U46769 (N_46769,N_42728,N_40323);
xnor U46770 (N_46770,N_40184,N_40020);
nor U46771 (N_46771,N_43366,N_41616);
and U46772 (N_46772,N_40682,N_44561);
nor U46773 (N_46773,N_43328,N_44988);
nand U46774 (N_46774,N_42707,N_41800);
and U46775 (N_46775,N_44645,N_42270);
xor U46776 (N_46776,N_40187,N_42533);
nor U46777 (N_46777,N_42518,N_44299);
and U46778 (N_46778,N_40334,N_41972);
xnor U46779 (N_46779,N_43184,N_41430);
or U46780 (N_46780,N_42793,N_42066);
nand U46781 (N_46781,N_42229,N_40037);
nor U46782 (N_46782,N_43926,N_42077);
and U46783 (N_46783,N_43299,N_41812);
and U46784 (N_46784,N_43118,N_43574);
nor U46785 (N_46785,N_43497,N_43379);
and U46786 (N_46786,N_43018,N_44268);
xnor U46787 (N_46787,N_42790,N_40984);
and U46788 (N_46788,N_44859,N_40399);
or U46789 (N_46789,N_43161,N_41273);
nor U46790 (N_46790,N_42808,N_40152);
and U46791 (N_46791,N_41306,N_40700);
and U46792 (N_46792,N_42055,N_43636);
or U46793 (N_46793,N_42522,N_44210);
and U46794 (N_46794,N_43420,N_44753);
and U46795 (N_46795,N_41910,N_43920);
xor U46796 (N_46796,N_41792,N_42153);
and U46797 (N_46797,N_42296,N_44726);
xor U46798 (N_46798,N_44926,N_42631);
and U46799 (N_46799,N_43818,N_41632);
and U46800 (N_46800,N_40833,N_43523);
nor U46801 (N_46801,N_42854,N_40133);
nor U46802 (N_46802,N_43670,N_43236);
nand U46803 (N_46803,N_41162,N_42769);
and U46804 (N_46804,N_40708,N_41470);
nand U46805 (N_46805,N_44703,N_40398);
xor U46806 (N_46806,N_43232,N_40246);
xnor U46807 (N_46807,N_44508,N_41168);
xor U46808 (N_46808,N_44311,N_43775);
xor U46809 (N_46809,N_41502,N_41129);
nand U46810 (N_46810,N_42926,N_44459);
or U46811 (N_46811,N_42183,N_42915);
nand U46812 (N_46812,N_44314,N_43982);
xnor U46813 (N_46813,N_42226,N_42280);
nor U46814 (N_46814,N_43500,N_44159);
nor U46815 (N_46815,N_44877,N_43681);
or U46816 (N_46816,N_40264,N_43210);
nor U46817 (N_46817,N_41862,N_40486);
nor U46818 (N_46818,N_43452,N_41725);
or U46819 (N_46819,N_41994,N_41070);
and U46820 (N_46820,N_40102,N_41029);
nand U46821 (N_46821,N_42869,N_41002);
xnor U46822 (N_46822,N_40309,N_41628);
and U46823 (N_46823,N_42302,N_40339);
nor U46824 (N_46824,N_40740,N_40774);
xor U46825 (N_46825,N_43396,N_41779);
and U46826 (N_46826,N_42852,N_42818);
or U46827 (N_46827,N_40841,N_43499);
nor U46828 (N_46828,N_42333,N_44648);
nand U46829 (N_46829,N_42411,N_44742);
nor U46830 (N_46830,N_44661,N_41158);
or U46831 (N_46831,N_43277,N_44853);
and U46832 (N_46832,N_40135,N_40789);
or U46833 (N_46833,N_41515,N_43144);
xor U46834 (N_46834,N_40552,N_40365);
nand U46835 (N_46835,N_43454,N_41406);
xor U46836 (N_46836,N_40445,N_40710);
nor U46837 (N_46837,N_43387,N_44994);
or U46838 (N_46838,N_42788,N_42305);
or U46839 (N_46839,N_40702,N_42786);
and U46840 (N_46840,N_40008,N_42188);
xnor U46841 (N_46841,N_44230,N_42571);
or U46842 (N_46842,N_40181,N_42565);
nor U46843 (N_46843,N_44388,N_42001);
xnor U46844 (N_46844,N_40828,N_40163);
nor U46845 (N_46845,N_40084,N_43627);
xor U46846 (N_46846,N_40278,N_42391);
and U46847 (N_46847,N_43760,N_44178);
xor U46848 (N_46848,N_44480,N_42712);
xnor U46849 (N_46849,N_43413,N_44415);
or U46850 (N_46850,N_43367,N_42376);
or U46851 (N_46851,N_44597,N_40127);
or U46852 (N_46852,N_43790,N_41609);
nand U46853 (N_46853,N_42159,N_41201);
nand U46854 (N_46854,N_41665,N_43302);
nand U46855 (N_46855,N_40248,N_42310);
xnor U46856 (N_46856,N_42236,N_40239);
nand U46857 (N_46857,N_42435,N_40186);
nand U46858 (N_46858,N_44045,N_44787);
and U46859 (N_46859,N_40092,N_43901);
xnor U46860 (N_46860,N_44971,N_41914);
nand U46861 (N_46861,N_43753,N_40200);
nand U46862 (N_46862,N_41997,N_40992);
and U46863 (N_46863,N_43888,N_42221);
xnor U46864 (N_46864,N_40462,N_43411);
nand U46865 (N_46865,N_43867,N_43743);
nor U46866 (N_46866,N_43265,N_44834);
and U46867 (N_46867,N_44788,N_40371);
nor U46868 (N_46868,N_41898,N_42345);
xnor U46869 (N_46869,N_42136,N_42952);
xnor U46870 (N_46870,N_43956,N_40208);
nand U46871 (N_46871,N_44356,N_40022);
nand U46872 (N_46872,N_42661,N_40456);
nor U46873 (N_46873,N_43089,N_40290);
and U46874 (N_46874,N_41582,N_43001);
nand U46875 (N_46875,N_40429,N_40614);
or U46876 (N_46876,N_41822,N_44352);
nor U46877 (N_46877,N_43310,N_43224);
nor U46878 (N_46878,N_41757,N_40213);
xnor U46879 (N_46879,N_43410,N_41358);
nand U46880 (N_46880,N_42775,N_41560);
xnor U46881 (N_46881,N_40107,N_44727);
nor U46882 (N_46882,N_41386,N_42035);
nand U46883 (N_46883,N_43152,N_42811);
xor U46884 (N_46884,N_41206,N_40880);
xor U46885 (N_46885,N_40060,N_43037);
nand U46886 (N_46886,N_40459,N_44169);
nand U46887 (N_46887,N_40227,N_43127);
and U46888 (N_46888,N_41566,N_42960);
xor U46889 (N_46889,N_43808,N_43319);
or U46890 (N_46890,N_40747,N_41859);
or U46891 (N_46891,N_42434,N_44554);
nor U46892 (N_46892,N_40059,N_43106);
or U46893 (N_46893,N_43800,N_44471);
nor U46894 (N_46894,N_41518,N_40666);
nand U46895 (N_46895,N_44001,N_44836);
nor U46896 (N_46896,N_41212,N_44911);
nor U46897 (N_46897,N_44069,N_41570);
or U46898 (N_46898,N_43924,N_41061);
xnor U46899 (N_46899,N_43021,N_41874);
and U46900 (N_46900,N_40515,N_43101);
xnor U46901 (N_46901,N_42997,N_40518);
xnor U46902 (N_46902,N_41623,N_41955);
xnor U46903 (N_46903,N_41692,N_44613);
and U46904 (N_46904,N_42656,N_43782);
xnor U46905 (N_46905,N_42396,N_42977);
xor U46906 (N_46906,N_43986,N_40383);
nor U46907 (N_46907,N_41123,N_40188);
xnor U46908 (N_46908,N_42951,N_42689);
and U46909 (N_46909,N_44658,N_40512);
nand U46910 (N_46910,N_42402,N_41722);
xor U46911 (N_46911,N_41668,N_42725);
xor U46912 (N_46912,N_44300,N_43780);
or U46913 (N_46913,N_43256,N_42129);
xor U46914 (N_46914,N_44241,N_43186);
nand U46915 (N_46915,N_42513,N_43248);
xor U46916 (N_46916,N_42529,N_42819);
or U46917 (N_46917,N_40403,N_41428);
nor U46918 (N_46918,N_42678,N_42870);
or U46919 (N_46919,N_41974,N_44762);
xor U46920 (N_46920,N_43594,N_41681);
nand U46921 (N_46921,N_42346,N_40955);
xnor U46922 (N_46922,N_43123,N_41402);
nor U46923 (N_46923,N_44615,N_43987);
nor U46924 (N_46924,N_43139,N_40315);
nand U46925 (N_46925,N_43201,N_43400);
nor U46926 (N_46926,N_41737,N_41562);
and U46927 (N_46927,N_42690,N_40245);
or U46928 (N_46928,N_44809,N_44028);
xnor U46929 (N_46929,N_41343,N_43493);
nand U46930 (N_46930,N_43148,N_40809);
and U46931 (N_46931,N_44071,N_42737);
or U46932 (N_46932,N_43290,N_41087);
nor U46933 (N_46933,N_43651,N_40298);
nand U46934 (N_46934,N_41559,N_40350);
nand U46935 (N_46935,N_43415,N_43358);
nand U46936 (N_46936,N_41130,N_40396);
nand U46937 (N_46937,N_41452,N_43276);
nor U46938 (N_46938,N_42998,N_44474);
or U46939 (N_46939,N_42162,N_41181);
or U46940 (N_46940,N_42840,N_42494);
nand U46941 (N_46941,N_40917,N_42890);
nand U46942 (N_46942,N_43892,N_43296);
and U46943 (N_46943,N_42912,N_43455);
or U46944 (N_46944,N_44298,N_42150);
xnor U46945 (N_46945,N_40088,N_40933);
or U46946 (N_46946,N_43709,N_40489);
or U46947 (N_46947,N_42354,N_42091);
nor U46948 (N_46948,N_44392,N_41313);
and U46949 (N_46949,N_44801,N_44675);
or U46950 (N_46950,N_44065,N_42151);
nor U46951 (N_46951,N_43568,N_44141);
or U46952 (N_46952,N_42773,N_41017);
nand U46953 (N_46953,N_41151,N_44608);
or U46954 (N_46954,N_43668,N_44878);
or U46955 (N_46955,N_43178,N_41516);
nor U46956 (N_46956,N_42227,N_40301);
xnor U46957 (N_46957,N_43824,N_42570);
and U46958 (N_46958,N_43949,N_43010);
xor U46959 (N_46959,N_42143,N_43786);
nor U46960 (N_46960,N_40792,N_44372);
and U46961 (N_46961,N_42579,N_42463);
or U46962 (N_46962,N_44552,N_43091);
and U46963 (N_46963,N_40496,N_44396);
and U46964 (N_46964,N_42482,N_42495);
or U46965 (N_46965,N_40815,N_41058);
nor U46966 (N_46966,N_41828,N_44839);
or U46967 (N_46967,N_40349,N_40904);
or U46968 (N_46968,N_42437,N_41836);
nor U46969 (N_46969,N_42802,N_43407);
nor U46970 (N_46970,N_43518,N_41604);
or U46971 (N_46971,N_40916,N_40872);
nor U46972 (N_46972,N_42444,N_40402);
nor U46973 (N_46973,N_40523,N_41221);
nor U46974 (N_46974,N_42095,N_44678);
nand U46975 (N_46975,N_44436,N_43643);
nor U46976 (N_46976,N_42659,N_43138);
nor U46977 (N_46977,N_44754,N_43428);
and U46978 (N_46978,N_41022,N_43552);
or U46979 (N_46979,N_44555,N_43799);
nor U46980 (N_46980,N_40259,N_44942);
or U46981 (N_46981,N_44822,N_41916);
nand U46982 (N_46982,N_44823,N_44428);
nand U46983 (N_46983,N_41754,N_42026);
xnor U46984 (N_46984,N_40779,N_44381);
xor U46985 (N_46985,N_44040,N_41014);
or U46986 (N_46986,N_44269,N_41373);
or U46987 (N_46987,N_40291,N_43418);
nor U46988 (N_46988,N_42469,N_43801);
nand U46989 (N_46989,N_44132,N_40844);
nand U46990 (N_46990,N_43109,N_44811);
and U46991 (N_46991,N_40327,N_43119);
or U46992 (N_46992,N_42868,N_40776);
or U46993 (N_46993,N_43720,N_41554);
xor U46994 (N_46994,N_40510,N_44087);
or U46995 (N_46995,N_40228,N_44632);
nor U46996 (N_46996,N_40793,N_43513);
or U46997 (N_46997,N_40344,N_40671);
xor U46998 (N_46998,N_41716,N_42127);
or U46999 (N_46999,N_41717,N_42816);
nand U47000 (N_47000,N_40214,N_40649);
xnor U47001 (N_47001,N_42307,N_40790);
nand U47002 (N_47002,N_42071,N_43505);
nor U47003 (N_47003,N_44009,N_41247);
nor U47004 (N_47004,N_42867,N_40501);
or U47005 (N_47005,N_41929,N_40630);
nand U47006 (N_47006,N_42194,N_40337);
or U47007 (N_47007,N_41990,N_42916);
or U47008 (N_47008,N_42700,N_40857);
and U47009 (N_47009,N_40068,N_42809);
or U47010 (N_47010,N_40906,N_42369);
nor U47011 (N_47011,N_42945,N_41627);
xor U47012 (N_47012,N_44730,N_43939);
xnor U47013 (N_47013,N_44738,N_40943);
xor U47014 (N_47014,N_40416,N_44140);
and U47015 (N_47015,N_42708,N_44172);
xor U47016 (N_47016,N_43414,N_40785);
nand U47017 (N_47017,N_42248,N_43323);
and U47018 (N_47018,N_42410,N_44845);
nor U47019 (N_47019,N_41603,N_44086);
and U47020 (N_47020,N_44655,N_41304);
nand U47021 (N_47021,N_40990,N_41001);
and U47022 (N_47022,N_41641,N_41224);
or U47023 (N_47023,N_43203,N_42799);
and U47024 (N_47024,N_44153,N_42260);
nand U47025 (N_47025,N_42503,N_44150);
nor U47026 (N_47026,N_42220,N_41797);
nand U47027 (N_47027,N_44497,N_41197);
and U47028 (N_47028,N_41048,N_44234);
and U47029 (N_47029,N_40364,N_40427);
and U47030 (N_47030,N_42516,N_40062);
nand U47031 (N_47031,N_41345,N_41829);
and U47032 (N_47032,N_41712,N_40753);
xor U47033 (N_47033,N_42070,N_44850);
nand U47034 (N_47034,N_44005,N_44856);
and U47035 (N_47035,N_44138,N_44231);
and U47036 (N_47036,N_44400,N_40604);
nor U47037 (N_47037,N_42263,N_41472);
or U47038 (N_47038,N_43936,N_41315);
or U47039 (N_47039,N_43150,N_41355);
nor U47040 (N_47040,N_42317,N_42780);
nor U47041 (N_47041,N_43324,N_40565);
xnor U47042 (N_47042,N_43376,N_40808);
or U47043 (N_47043,N_42900,N_42105);
xnor U47044 (N_47044,N_44202,N_43706);
nor U47045 (N_47045,N_40479,N_41018);
nor U47046 (N_47046,N_44757,N_44968);
nand U47047 (N_47047,N_41866,N_41709);
nor U47048 (N_47048,N_44548,N_43408);
nand U47049 (N_47049,N_41984,N_40693);
nor U47050 (N_47050,N_40204,N_44997);
or U47051 (N_47051,N_42751,N_40066);
xor U47052 (N_47052,N_42746,N_42239);
xor U47053 (N_47053,N_42099,N_40888);
nand U47054 (N_47054,N_41282,N_41564);
and U47055 (N_47055,N_44637,N_43431);
xor U47056 (N_47056,N_41311,N_41110);
and U47057 (N_47057,N_42922,N_40001);
or U47058 (N_47058,N_43317,N_41215);
xnor U47059 (N_47059,N_42067,N_43331);
or U47060 (N_47060,N_40232,N_42767);
nand U47061 (N_47061,N_42265,N_44559);
or U47062 (N_47062,N_41145,N_43050);
nor U47063 (N_47063,N_41739,N_42633);
or U47064 (N_47064,N_43432,N_43965);
xor U47065 (N_47065,N_43942,N_43578);
nor U47066 (N_47066,N_42921,N_44136);
or U47067 (N_47067,N_41059,N_43424);
xor U47068 (N_47068,N_42180,N_41253);
or U47069 (N_47069,N_40577,N_42267);
or U47070 (N_47070,N_42836,N_44847);
or U47071 (N_47071,N_40069,N_41977);
and U47072 (N_47072,N_40355,N_44516);
nand U47073 (N_47073,N_44786,N_42787);
nor U47074 (N_47074,N_42243,N_42763);
xnor U47075 (N_47075,N_43200,N_40381);
nand U47076 (N_47076,N_40495,N_42535);
and U47077 (N_47077,N_40598,N_42115);
and U47078 (N_47078,N_40556,N_40864);
xnor U47079 (N_47079,N_43571,N_41132);
and U47080 (N_47080,N_40856,N_41106);
nand U47081 (N_47081,N_43904,N_44744);
xor U47082 (N_47082,N_42561,N_40579);
and U47083 (N_47083,N_41283,N_42505);
xnor U47084 (N_47084,N_43930,N_40247);
and U47085 (N_47085,N_43166,N_40911);
and U47086 (N_47086,N_42387,N_43692);
or U47087 (N_47087,N_43665,N_40302);
nand U47088 (N_47088,N_42507,N_43896);
xnor U47089 (N_47089,N_40373,N_41290);
or U47090 (N_47090,N_44339,N_42079);
nor U47091 (N_47091,N_41704,N_44618);
nand U47092 (N_47092,N_43039,N_44421);
and U47093 (N_47093,N_43646,N_44517);
nand U47094 (N_47094,N_41155,N_43267);
nor U47095 (N_47095,N_43160,N_44848);
and U47096 (N_47096,N_41539,N_43346);
xnor U47097 (N_47097,N_42297,N_44395);
nand U47098 (N_47098,N_44242,N_41965);
and U47099 (N_47099,N_43525,N_42293);
nand U47100 (N_47100,N_40517,N_40284);
nor U47101 (N_47101,N_40484,N_40624);
and U47102 (N_47102,N_40974,N_40253);
and U47103 (N_47103,N_44485,N_40799);
nor U47104 (N_47104,N_44032,N_41904);
xnor U47105 (N_47105,N_40662,N_41971);
nand U47106 (N_47106,N_41285,N_43694);
xnor U47107 (N_47107,N_41565,N_44389);
or U47108 (N_47108,N_42161,N_44283);
nor U47109 (N_47109,N_40670,N_42366);
and U47110 (N_47110,N_41817,N_40678);
xnor U47111 (N_47111,N_42254,N_40616);
nor U47112 (N_47112,N_43870,N_40379);
nand U47113 (N_47113,N_44929,N_42504);
xor U47114 (N_47114,N_40909,N_42431);
and U47115 (N_47115,N_43269,N_41899);
nand U47116 (N_47116,N_44062,N_42492);
or U47117 (N_47117,N_42942,N_43473);
and U47118 (N_47118,N_42282,N_43537);
xor U47119 (N_47119,N_41234,N_41351);
xnor U47120 (N_47120,N_44329,N_44357);
and U47121 (N_47121,N_40568,N_43077);
nor U47122 (N_47122,N_40676,N_44341);
nor U47123 (N_47123,N_43773,N_42480);
or U47124 (N_47124,N_43612,N_42782);
nor U47125 (N_47125,N_44871,N_42489);
xnor U47126 (N_47126,N_40728,N_44827);
nor U47127 (N_47127,N_41166,N_42943);
and U47128 (N_47128,N_41321,N_40142);
xor U47129 (N_47129,N_44672,N_44404);
nand U47130 (N_47130,N_44656,N_42999);
nor U47131 (N_47131,N_40094,N_43616);
xnor U47132 (N_47132,N_44736,N_42458);
xnor U47133 (N_47133,N_40991,N_41170);
or U47134 (N_47134,N_42693,N_40821);
nor U47135 (N_47135,N_43748,N_40442);
xor U47136 (N_47136,N_43675,N_42831);
or U47137 (N_47137,N_40788,N_43211);
nand U47138 (N_47138,N_41277,N_41635);
nand U47139 (N_47139,N_44183,N_42791);
and U47140 (N_47140,N_40963,N_41947);
or U47141 (N_47141,N_42027,N_41252);
xor U47142 (N_47142,N_42917,N_42138);
xor U47143 (N_47143,N_42073,N_43846);
nand U47144 (N_47144,N_40701,N_42627);
nor U47145 (N_47145,N_44594,N_40985);
and U47146 (N_47146,N_41948,N_43793);
nor U47147 (N_47147,N_44148,N_43405);
or U47148 (N_47148,N_41425,N_40171);
xor U47149 (N_47149,N_43422,N_44073);
nor U47150 (N_47150,N_40845,N_44166);
nand U47151 (N_47151,N_44688,N_42956);
nand U47152 (N_47152,N_42114,N_43105);
and U47153 (N_47153,N_41466,N_42552);
xnor U47154 (N_47154,N_43581,N_42893);
nor U47155 (N_47155,N_41572,N_44818);
nand U47156 (N_47156,N_40646,N_42053);
nand U47157 (N_47157,N_41135,N_40658);
nand U47158 (N_47158,N_43273,N_41457);
or U47159 (N_47159,N_40203,N_41555);
or U47160 (N_47160,N_43531,N_43655);
nor U47161 (N_47161,N_44467,N_44536);
xor U47162 (N_47162,N_43550,N_43476);
and U47163 (N_47163,N_41451,N_42041);
and U47164 (N_47164,N_44042,N_44491);
nand U47165 (N_47165,N_42488,N_43845);
and U47166 (N_47166,N_44052,N_40860);
nand U47167 (N_47167,N_41074,N_40742);
nand U47168 (N_47168,N_41512,N_44235);
xnor U47169 (N_47169,N_40318,N_43804);
xnor U47170 (N_47170,N_43264,N_43606);
xnor U47171 (N_47171,N_43045,N_42404);
and U47172 (N_47172,N_41279,N_41310);
xnor U47173 (N_47173,N_41557,N_44363);
and U47174 (N_47174,N_41806,N_42021);
and U47175 (N_47175,N_43906,N_44734);
or U47176 (N_47176,N_41698,N_40391);
and U47177 (N_47177,N_43912,N_40458);
xor U47178 (N_47178,N_40480,N_41723);
and U47179 (N_47179,N_42251,N_44422);
or U47180 (N_47180,N_44987,N_41329);
and U47181 (N_47181,N_40448,N_44280);
xor U47182 (N_47182,N_42473,N_41601);
and U47183 (N_47183,N_44403,N_44145);
xor U47184 (N_47184,N_41629,N_43459);
nor U47185 (N_47185,N_43941,N_41776);
xnor U47186 (N_47186,N_41885,N_40761);
nor U47187 (N_47187,N_40661,N_42139);
nand U47188 (N_47188,N_41314,N_44133);
or U47189 (N_47189,N_43363,N_43294);
xor U47190 (N_47190,N_41165,N_42739);
xnor U47191 (N_47191,N_41362,N_41403);
and U47192 (N_47192,N_40206,N_40557);
nor U47193 (N_47193,N_40707,N_41777);
and U47194 (N_47194,N_41818,N_41334);
or U47195 (N_47195,N_43564,N_43314);
nand U47196 (N_47196,N_44640,N_40254);
nand U47197 (N_47197,N_43131,N_42515);
or U47198 (N_47198,N_42373,N_43180);
or U47199 (N_47199,N_44029,N_41453);
nand U47200 (N_47200,N_40217,N_40235);
nand U47201 (N_47201,N_41596,N_41312);
and U47202 (N_47202,N_40972,N_40424);
nand U47203 (N_47203,N_43225,N_43749);
nand U47204 (N_47204,N_42812,N_41545);
or U47205 (N_47205,N_42054,N_43128);
nor U47206 (N_47206,N_42195,N_42976);
xnor U47207 (N_47207,N_44767,N_41724);
nand U47208 (N_47208,N_42140,N_43190);
and U47209 (N_47209,N_42744,N_40316);
or U47210 (N_47210,N_42968,N_40997);
nand U47211 (N_47211,N_42657,N_41046);
nand U47212 (N_47212,N_44281,N_42560);
xor U47213 (N_47213,N_42680,N_44303);
nor U47214 (N_47214,N_44888,N_43271);
nor U47215 (N_47215,N_42531,N_44058);
xnor U47216 (N_47216,N_42598,N_41813);
xor U47217 (N_47217,N_44545,N_44387);
nor U47218 (N_47218,N_43830,N_41210);
xor U47219 (N_47219,N_40386,N_42181);
xor U47220 (N_47220,N_41275,N_42781);
nor U47221 (N_47221,N_43795,N_40354);
and U47222 (N_47222,N_40288,N_44956);
and U47223 (N_47223,N_40393,N_42004);
nand U47224 (N_47224,N_44693,N_40781);
nand U47225 (N_47225,N_40802,N_43072);
xor U47226 (N_47226,N_44532,N_40683);
nor U47227 (N_47227,N_43003,N_42134);
nor U47228 (N_47228,N_44796,N_43980);
and U47229 (N_47229,N_42901,N_41680);
nand U47230 (N_47230,N_43004,N_43922);
and U47231 (N_47231,N_41147,N_42279);
or U47232 (N_47232,N_42102,N_43437);
nand U47233 (N_47233,N_43479,N_43589);
xnor U47234 (N_47234,N_41988,N_41459);
nor U47235 (N_47235,N_42762,N_43765);
or U47236 (N_47236,N_40907,N_44932);
xor U47237 (N_47237,N_41360,N_43539);
nand U47238 (N_47238,N_40287,N_44973);
and U47239 (N_47239,N_40463,N_43235);
xnor U47240 (N_47240,N_41473,N_40959);
or U47241 (N_47241,N_44217,N_40032);
nor U47242 (N_47242,N_44698,N_41038);
nand U47243 (N_47243,N_42501,N_43992);
or U47244 (N_47244,N_40443,N_41975);
nand U47245 (N_47245,N_40297,N_44174);
xnor U47246 (N_47246,N_41326,N_43445);
and U47247 (N_47247,N_40388,N_41666);
or U47248 (N_47248,N_43717,N_43503);
xnor U47249 (N_47249,N_44633,N_44780);
nand U47250 (N_47250,N_43504,N_41781);
or U47251 (N_47251,N_43197,N_40550);
xnor U47252 (N_47252,N_43524,N_44568);
or U47253 (N_47253,N_43788,N_40734);
nand U47254 (N_47254,N_44574,N_42121);
and U47255 (N_47255,N_44776,N_40759);
nor U47256 (N_47256,N_44980,N_41008);
nor U47257 (N_47257,N_40591,N_44900);
xnor U47258 (N_47258,N_44484,N_43971);
xnor U47259 (N_47259,N_43060,N_40733);
nand U47260 (N_47260,N_42193,N_42950);
nor U47261 (N_47261,N_44266,N_40385);
xnor U47262 (N_47262,N_44885,N_41099);
nor U47263 (N_47263,N_42896,N_42553);
nor U47264 (N_47264,N_43819,N_40134);
nor U47265 (N_47265,N_44222,N_42045);
xor U47266 (N_47266,N_44091,N_41961);
xor U47267 (N_47267,N_41938,N_40160);
nand U47268 (N_47268,N_42204,N_42650);
and U47269 (N_47269,N_44275,N_42607);
and U47270 (N_47270,N_44204,N_44627);
and U47271 (N_47271,N_41497,N_40533);
and U47272 (N_47272,N_44013,N_42794);
nor U47273 (N_47273,N_40286,N_44330);
xnor U47274 (N_47274,N_40207,N_44628);
xnor U47275 (N_47275,N_43330,N_43617);
nor U47276 (N_47276,N_40703,N_41177);
nand U47277 (N_47277,N_41846,N_43741);
and U47278 (N_47278,N_42980,N_40322);
nand U47279 (N_47279,N_41347,N_44981);
nand U47280 (N_47280,N_42982,N_41799);
or U47281 (N_47281,N_44965,N_42839);
nor U47282 (N_47282,N_44438,N_44747);
xnor U47283 (N_47283,N_42316,N_43115);
nand U47284 (N_47284,N_40673,N_40558);
nor U47285 (N_47285,N_40378,N_44925);
or U47286 (N_47286,N_40894,N_43947);
or U47287 (N_47287,N_40887,N_43392);
or U47288 (N_47288,N_41082,N_41619);
xor U47289 (N_47289,N_40787,N_41826);
or U47290 (N_47290,N_40083,N_42616);
and U47291 (N_47291,N_40112,N_42203);
nor U47292 (N_47292,N_44442,N_42323);
xor U47293 (N_47293,N_40425,N_40597);
or U47294 (N_47294,N_43851,N_44650);
and U47295 (N_47295,N_44113,N_44250);
or U47296 (N_47296,N_44325,N_41708);
nor U47297 (N_47297,N_41750,N_43158);
nand U47298 (N_47298,N_43557,N_44924);
nor U47299 (N_47299,N_43679,N_41814);
xnor U47300 (N_47300,N_41720,N_44606);
nand U47301 (N_47301,N_40280,N_40573);
nor U47302 (N_47302,N_43562,N_44315);
nand U47303 (N_47303,N_42337,N_42484);
and U47304 (N_47304,N_43165,N_41664);
and U47305 (N_47305,N_44607,N_44914);
and U47306 (N_47306,N_42880,N_40599);
nor U47307 (N_47307,N_43506,N_41039);
xor U47308 (N_47308,N_44405,N_44060);
nor U47309 (N_47309,N_42643,N_40003);
and U47310 (N_47310,N_42000,N_43998);
nand U47311 (N_47311,N_40704,N_43558);
and U47312 (N_47312,N_42068,N_43690);
nor U47313 (N_47313,N_44663,N_42379);
and U47314 (N_47314,N_41973,N_43327);
and U47315 (N_47315,N_40474,N_44147);
nand U47316 (N_47316,N_40147,N_44193);
nor U47317 (N_47317,N_43183,N_43234);
xnor U47318 (N_47318,N_44601,N_41034);
nand U47319 (N_47319,N_43916,N_40130);
nor U47320 (N_47320,N_42292,N_41639);
or U47321 (N_47321,N_40464,N_42822);
or U47322 (N_47322,N_41411,N_42078);
nor U47323 (N_47323,N_40460,N_42986);
nor U47324 (N_47324,N_44209,N_41775);
and U47325 (N_47325,N_41093,N_44030);
nand U47326 (N_47326,N_41493,N_40929);
or U47327 (N_47327,N_40357,N_43071);
nand U47328 (N_47328,N_42020,N_43698);
or U47329 (N_47329,N_43054,N_42996);
xnor U47330 (N_47330,N_44502,N_41137);
nand U47331 (N_47331,N_41719,N_40115);
xnor U47332 (N_47332,N_40033,N_44649);
nand U47333 (N_47333,N_40241,N_43048);
or U47334 (N_47334,N_42165,N_40878);
or U47335 (N_47335,N_42395,N_43412);
nand U47336 (N_47336,N_43620,N_41225);
nand U47337 (N_47337,N_43238,N_40074);
nand U47338 (N_47338,N_41342,N_41579);
xnor U47339 (N_47339,N_44457,N_42634);
and U47340 (N_47340,N_41195,N_44623);
and U47341 (N_47341,N_44600,N_44831);
and U47342 (N_47342,N_44326,N_43239);
and U47343 (N_47343,N_44587,N_44051);
nand U47344 (N_47344,N_44265,N_43436);
and U47345 (N_47345,N_44492,N_42031);
nor U47346 (N_47346,N_43677,N_42051);
nor U47347 (N_47347,N_43074,N_41044);
xor U47348 (N_47348,N_42049,N_40527);
xnor U47349 (N_47349,N_42462,N_41707);
nor U47350 (N_47350,N_40778,N_44867);
or U47351 (N_47351,N_42485,N_44577);
nand U47352 (N_47352,N_41299,N_41688);
xnor U47353 (N_47353,N_40737,N_42024);
xnor U47354 (N_47354,N_40892,N_44993);
xnor U47355 (N_47355,N_41563,N_40641);
and U47356 (N_47356,N_43853,N_40867);
and U47357 (N_47357,N_43966,N_42486);
or U47358 (N_47358,N_43114,N_44223);
nand U47359 (N_47359,N_40476,N_40118);
or U47360 (N_47360,N_40116,N_44197);
nand U47361 (N_47361,N_40376,N_42874);
or U47362 (N_47362,N_42534,N_43381);
nor U47363 (N_47363,N_41901,N_41240);
or U47364 (N_47364,N_42748,N_43584);
or U47365 (N_47365,N_44489,N_41142);
nand U47366 (N_47366,N_42892,N_42367);
nand U47367 (N_47367,N_42281,N_42732);
and U47368 (N_47368,N_41354,N_41856);
nand U47369 (N_47369,N_40081,N_44721);
and U47370 (N_47370,N_41759,N_44844);
nand U47371 (N_47371,N_44515,N_41086);
or U47372 (N_47372,N_43362,N_44369);
and U47373 (N_47373,N_43480,N_42932);
nor U47374 (N_47374,N_41833,N_44249);
or U47375 (N_47375,N_43067,N_41606);
xor U47376 (N_47376,N_43530,N_42881);
xnor U47377 (N_47377,N_44857,N_44080);
and U47378 (N_47378,N_41577,N_42052);
or U47379 (N_47379,N_41549,N_42745);
and U47380 (N_47380,N_41837,N_40205);
and U47381 (N_47381,N_43120,N_43661);
nand U47382 (N_47382,N_43948,N_43206);
nand U47383 (N_47383,N_41903,N_44487);
xnor U47384 (N_47384,N_42731,N_43329);
xnor U47385 (N_47385,N_40859,N_42603);
xnor U47386 (N_47386,N_43758,N_43008);
xor U47387 (N_47387,N_44880,N_43771);
nor U47388 (N_47388,N_43744,N_40312);
nand U47389 (N_47389,N_42569,N_41332);
nor U47390 (N_47390,N_40745,N_42406);
and U47391 (N_47391,N_40149,N_43900);
nor U47392 (N_47392,N_40099,N_44910);
xnor U47393 (N_47393,N_41270,N_44002);
or U47394 (N_47394,N_41686,N_42112);
xor U47395 (N_47395,N_40619,N_43364);
and U47396 (N_47396,N_40919,N_43313);
nor U47397 (N_47397,N_43222,N_41120);
nand U47398 (N_47398,N_41391,N_44504);
and U47399 (N_47399,N_44208,N_41054);
xnor U47400 (N_47400,N_44165,N_44538);
nand U47401 (N_47401,N_41368,N_40180);
nor U47402 (N_47402,N_40825,N_42664);
or U47403 (N_47403,N_40688,N_43856);
or U47404 (N_47404,N_44572,N_43945);
or U47405 (N_47405,N_43721,N_43442);
or U47406 (N_47406,N_43671,N_43747);
nor U47407 (N_47407,N_41040,N_40119);
xor U47408 (N_47408,N_44112,N_43701);
nor U47409 (N_47409,N_41573,N_42493);
xor U47410 (N_47410,N_42651,N_44902);
nand U47411 (N_47411,N_43372,N_41455);
xnor U47412 (N_47412,N_44872,N_41205);
xnor U47413 (N_47413,N_40313,N_44550);
nor U47414 (N_47414,N_42855,N_41340);
xor U47415 (N_47415,N_43320,N_42146);
and U47416 (N_47416,N_43189,N_42247);
or U47417 (N_47417,N_42141,N_41980);
or U47418 (N_47418,N_40705,N_44458);
nor U47419 (N_47419,N_44198,N_43875);
xnor U47420 (N_47420,N_42393,N_44406);
or U47421 (N_47421,N_44307,N_43261);
nand U47422 (N_47422,N_43638,N_42017);
or U47423 (N_47423,N_44379,N_43809);
nor U47424 (N_47424,N_43757,N_40267);
or U47425 (N_47425,N_43009,N_43725);
xnor U47426 (N_47426,N_42927,N_40454);
nand U47427 (N_47427,N_41246,N_41520);
nor U47428 (N_47428,N_42801,N_40621);
nand U47429 (N_47429,N_41260,N_43784);
nor U47430 (N_47430,N_44937,N_40346);
and U47431 (N_47431,N_43038,N_40901);
or U47432 (N_47432,N_42132,N_43453);
nor U47433 (N_47433,N_40850,N_41103);
and U47434 (N_47434,N_40777,N_44473);
nor U47435 (N_47435,N_40277,N_40958);
and U47436 (N_47436,N_42460,N_41268);
and U47437 (N_47437,N_42539,N_42740);
nand U47438 (N_47438,N_44472,N_42093);
and U47439 (N_47439,N_43300,N_43233);
nor U47440 (N_47440,N_40551,N_44874);
xnor U47441 (N_47441,N_44371,N_40335);
xnor U47442 (N_47442,N_42665,N_41608);
nand U47443 (N_47443,N_42009,N_44891);
xnor U47444 (N_47444,N_41605,N_40064);
nand U47445 (N_47445,N_44756,N_42557);
nand U47446 (N_47446,N_42131,N_43258);
or U47447 (N_47447,N_40780,N_41226);
xnor U47448 (N_47448,N_41190,N_41006);
nand U47449 (N_47449,N_41592,N_44452);
nand U47450 (N_47450,N_42142,N_40122);
nor U47451 (N_47451,N_40356,N_42312);
xor U47452 (N_47452,N_42764,N_40971);
nand U47453 (N_47453,N_44286,N_44111);
nand U47454 (N_47454,N_44916,N_44626);
and U47455 (N_47455,N_42228,N_43164);
or U47456 (N_47456,N_44366,N_41710);
and U47457 (N_47457,N_40645,N_44016);
or U47458 (N_47458,N_43465,N_44364);
xnor U47459 (N_47459,N_44642,N_44905);
or U47460 (N_47460,N_42990,N_40796);
nand U47461 (N_47461,N_42837,N_44308);
xnor U47462 (N_47462,N_40215,N_42388);
xnor U47463 (N_47463,N_44179,N_41513);
and U47464 (N_47464,N_42554,N_40618);
and U47465 (N_47465,N_43390,N_41256);
and U47466 (N_47466,N_42089,N_43215);
and U47467 (N_47467,N_44763,N_40942);
nor U47468 (N_47468,N_41858,N_44078);
and U47469 (N_47469,N_43815,N_40308);
xor U47470 (N_47470,N_44083,N_42750);
and U47471 (N_47471,N_41589,N_43451);
nand U47472 (N_47472,N_43157,N_44803);
nand U47473 (N_47473,N_41752,N_44191);
nor U47474 (N_47474,N_40948,N_41892);
nor U47475 (N_47475,N_44496,N_44170);
or U47476 (N_47476,N_43092,N_40921);
or U47477 (N_47477,N_40586,N_40763);
and U47478 (N_47478,N_41653,N_44697);
nand U47479 (N_47479,N_43723,N_42364);
nand U47480 (N_47480,N_41144,N_44407);
nor U47481 (N_47481,N_44622,N_40226);
xor U47482 (N_47482,N_42674,N_44412);
nand U47483 (N_47483,N_44715,N_43860);
or U47484 (N_47484,N_44134,N_43369);
nor U47485 (N_47485,N_43326,N_41908);
or U47486 (N_47486,N_43880,N_41507);
or U47487 (N_47487,N_40444,N_42859);
nand U47488 (N_47488,N_40623,N_44119);
xor U47489 (N_47489,N_42241,N_42308);
nor U47490 (N_47490,N_40390,N_43282);
nor U47491 (N_47491,N_41674,N_44247);
and U47492 (N_47492,N_42761,N_44593);
or U47493 (N_47493,N_44075,N_40941);
nor U47494 (N_47494,N_40307,N_41049);
nand U47495 (N_47495,N_41422,N_43145);
xnor U47496 (N_47496,N_43125,N_40260);
or U47497 (N_47497,N_41394,N_40961);
and U47498 (N_47498,N_42023,N_41924);
and U47499 (N_47499,N_43512,N_42169);
xnor U47500 (N_47500,N_44552,N_40487);
and U47501 (N_47501,N_43676,N_41415);
and U47502 (N_47502,N_40382,N_41093);
or U47503 (N_47503,N_43600,N_42263);
or U47504 (N_47504,N_43640,N_44391);
or U47505 (N_47505,N_44287,N_41447);
or U47506 (N_47506,N_44879,N_40104);
nand U47507 (N_47507,N_44646,N_41802);
nand U47508 (N_47508,N_41879,N_42096);
or U47509 (N_47509,N_44890,N_41785);
or U47510 (N_47510,N_42210,N_41924);
xor U47511 (N_47511,N_44957,N_40467);
and U47512 (N_47512,N_44263,N_44649);
and U47513 (N_47513,N_42106,N_44457);
xnor U47514 (N_47514,N_40115,N_44294);
nor U47515 (N_47515,N_43419,N_44284);
or U47516 (N_47516,N_40024,N_43338);
or U47517 (N_47517,N_42363,N_42263);
xnor U47518 (N_47518,N_43696,N_43360);
nand U47519 (N_47519,N_41063,N_44078);
nand U47520 (N_47520,N_44085,N_44922);
nor U47521 (N_47521,N_41884,N_43709);
and U47522 (N_47522,N_40781,N_41162);
nand U47523 (N_47523,N_40722,N_40834);
or U47524 (N_47524,N_41420,N_42981);
and U47525 (N_47525,N_41540,N_44813);
nand U47526 (N_47526,N_44770,N_42989);
nand U47527 (N_47527,N_40408,N_43753);
nor U47528 (N_47528,N_44357,N_42163);
nor U47529 (N_47529,N_44565,N_41881);
xor U47530 (N_47530,N_40327,N_44775);
or U47531 (N_47531,N_41488,N_43964);
and U47532 (N_47532,N_44808,N_44489);
nor U47533 (N_47533,N_41583,N_41165);
nand U47534 (N_47534,N_43341,N_42729);
nor U47535 (N_47535,N_44802,N_44701);
nand U47536 (N_47536,N_44345,N_43254);
nor U47537 (N_47537,N_40611,N_44906);
xor U47538 (N_47538,N_43879,N_43896);
nand U47539 (N_47539,N_43570,N_41691);
xor U47540 (N_47540,N_44378,N_43026);
nor U47541 (N_47541,N_41010,N_42432);
xor U47542 (N_47542,N_42887,N_40145);
nor U47543 (N_47543,N_44836,N_44881);
and U47544 (N_47544,N_41683,N_41026);
and U47545 (N_47545,N_41689,N_42865);
nand U47546 (N_47546,N_40545,N_43689);
and U47547 (N_47547,N_40645,N_41313);
nor U47548 (N_47548,N_42296,N_44953);
nor U47549 (N_47549,N_40645,N_43584);
xnor U47550 (N_47550,N_41858,N_43671);
xor U47551 (N_47551,N_41395,N_42569);
or U47552 (N_47552,N_43890,N_43506);
and U47553 (N_47553,N_41577,N_42082);
and U47554 (N_47554,N_43517,N_43918);
and U47555 (N_47555,N_44698,N_41093);
nor U47556 (N_47556,N_44058,N_40886);
xnor U47557 (N_47557,N_42918,N_44203);
nor U47558 (N_47558,N_41397,N_44634);
and U47559 (N_47559,N_43871,N_40971);
xnor U47560 (N_47560,N_40763,N_44764);
nand U47561 (N_47561,N_42546,N_40229);
or U47562 (N_47562,N_40997,N_42253);
xor U47563 (N_47563,N_43021,N_42620);
nor U47564 (N_47564,N_40953,N_44244);
or U47565 (N_47565,N_44794,N_40213);
or U47566 (N_47566,N_44092,N_42728);
nand U47567 (N_47567,N_41334,N_43909);
xnor U47568 (N_47568,N_44179,N_44509);
xnor U47569 (N_47569,N_44340,N_42291);
or U47570 (N_47570,N_43152,N_44703);
nor U47571 (N_47571,N_40799,N_43049);
nand U47572 (N_47572,N_43639,N_40939);
nand U47573 (N_47573,N_44781,N_44168);
nor U47574 (N_47574,N_44398,N_40261);
or U47575 (N_47575,N_40521,N_43434);
nor U47576 (N_47576,N_41644,N_40155);
nand U47577 (N_47577,N_43041,N_44079);
nor U47578 (N_47578,N_43173,N_42287);
and U47579 (N_47579,N_40642,N_44953);
nor U47580 (N_47580,N_40255,N_41699);
or U47581 (N_47581,N_41640,N_44355);
or U47582 (N_47582,N_40714,N_40217);
xor U47583 (N_47583,N_41232,N_43869);
xor U47584 (N_47584,N_41487,N_40155);
or U47585 (N_47585,N_43301,N_42268);
nor U47586 (N_47586,N_42174,N_43486);
nor U47587 (N_47587,N_43015,N_44509);
nand U47588 (N_47588,N_41410,N_40147);
nor U47589 (N_47589,N_43378,N_40938);
nor U47590 (N_47590,N_44427,N_42662);
nor U47591 (N_47591,N_40035,N_44015);
or U47592 (N_47592,N_43995,N_41063);
and U47593 (N_47593,N_42203,N_42435);
nor U47594 (N_47594,N_44558,N_43103);
and U47595 (N_47595,N_42930,N_43181);
or U47596 (N_47596,N_44054,N_41001);
nor U47597 (N_47597,N_41990,N_44894);
xnor U47598 (N_47598,N_41922,N_44029);
nor U47599 (N_47599,N_42557,N_41666);
nor U47600 (N_47600,N_41533,N_42823);
xor U47601 (N_47601,N_43033,N_40085);
and U47602 (N_47602,N_41841,N_44889);
or U47603 (N_47603,N_40175,N_40838);
nor U47604 (N_47604,N_42155,N_41140);
nand U47605 (N_47605,N_44698,N_43034);
xor U47606 (N_47606,N_43416,N_44700);
and U47607 (N_47607,N_43631,N_44273);
nor U47608 (N_47608,N_40416,N_41856);
xor U47609 (N_47609,N_40366,N_41175);
and U47610 (N_47610,N_40984,N_43888);
xor U47611 (N_47611,N_40286,N_42977);
or U47612 (N_47612,N_43316,N_41430);
xor U47613 (N_47613,N_42354,N_42613);
nor U47614 (N_47614,N_43013,N_40867);
xnor U47615 (N_47615,N_40220,N_42171);
or U47616 (N_47616,N_40374,N_40546);
xor U47617 (N_47617,N_40662,N_41427);
nor U47618 (N_47618,N_42001,N_42349);
and U47619 (N_47619,N_40886,N_44737);
xor U47620 (N_47620,N_41774,N_42832);
nand U47621 (N_47621,N_41492,N_44253);
and U47622 (N_47622,N_42196,N_41924);
nand U47623 (N_47623,N_43031,N_43558);
xor U47624 (N_47624,N_40914,N_44772);
nor U47625 (N_47625,N_40864,N_40887);
and U47626 (N_47626,N_40189,N_40335);
nand U47627 (N_47627,N_42078,N_44580);
xnor U47628 (N_47628,N_43228,N_40002);
or U47629 (N_47629,N_40129,N_41158);
nand U47630 (N_47630,N_42764,N_40844);
or U47631 (N_47631,N_42691,N_42384);
nand U47632 (N_47632,N_41910,N_41889);
nor U47633 (N_47633,N_41382,N_43899);
nor U47634 (N_47634,N_43963,N_41643);
nand U47635 (N_47635,N_40443,N_42773);
and U47636 (N_47636,N_42722,N_40526);
xor U47637 (N_47637,N_43007,N_40964);
nand U47638 (N_47638,N_43389,N_40337);
and U47639 (N_47639,N_40952,N_41395);
and U47640 (N_47640,N_42611,N_41422);
or U47641 (N_47641,N_41226,N_42221);
xor U47642 (N_47642,N_41316,N_41340);
and U47643 (N_47643,N_44957,N_40818);
nand U47644 (N_47644,N_43786,N_43016);
nor U47645 (N_47645,N_41144,N_40090);
nor U47646 (N_47646,N_40616,N_41749);
xnor U47647 (N_47647,N_44926,N_40283);
nand U47648 (N_47648,N_42166,N_43479);
and U47649 (N_47649,N_40798,N_40391);
xor U47650 (N_47650,N_43616,N_40319);
or U47651 (N_47651,N_40872,N_43163);
or U47652 (N_47652,N_40669,N_43359);
nor U47653 (N_47653,N_42341,N_42985);
and U47654 (N_47654,N_42311,N_42027);
or U47655 (N_47655,N_43856,N_40089);
and U47656 (N_47656,N_43336,N_40830);
or U47657 (N_47657,N_44939,N_43210);
nor U47658 (N_47658,N_44149,N_42497);
xor U47659 (N_47659,N_43637,N_40227);
xor U47660 (N_47660,N_44494,N_44547);
xnor U47661 (N_47661,N_42675,N_44310);
or U47662 (N_47662,N_44473,N_41590);
and U47663 (N_47663,N_42566,N_42001);
or U47664 (N_47664,N_43424,N_40189);
nand U47665 (N_47665,N_40838,N_40630);
nor U47666 (N_47666,N_40071,N_40596);
nor U47667 (N_47667,N_43654,N_42601);
nor U47668 (N_47668,N_40457,N_41976);
nor U47669 (N_47669,N_42704,N_40473);
nand U47670 (N_47670,N_41084,N_40930);
xnor U47671 (N_47671,N_44444,N_41583);
and U47672 (N_47672,N_43784,N_41268);
and U47673 (N_47673,N_43362,N_44975);
or U47674 (N_47674,N_44771,N_40518);
nor U47675 (N_47675,N_43496,N_44980);
xor U47676 (N_47676,N_42004,N_40100);
xnor U47677 (N_47677,N_42364,N_41433);
nand U47678 (N_47678,N_42767,N_40321);
and U47679 (N_47679,N_44600,N_42322);
and U47680 (N_47680,N_43849,N_44245);
or U47681 (N_47681,N_42178,N_41850);
or U47682 (N_47682,N_42051,N_41064);
nor U47683 (N_47683,N_43900,N_40340);
nor U47684 (N_47684,N_42860,N_44571);
or U47685 (N_47685,N_40772,N_41371);
nor U47686 (N_47686,N_44099,N_42283);
nand U47687 (N_47687,N_40843,N_41049);
nand U47688 (N_47688,N_41967,N_42891);
and U47689 (N_47689,N_44459,N_44621);
nor U47690 (N_47690,N_43743,N_43624);
or U47691 (N_47691,N_43034,N_42683);
and U47692 (N_47692,N_43112,N_41141);
xnor U47693 (N_47693,N_42812,N_41094);
and U47694 (N_47694,N_41622,N_43514);
nand U47695 (N_47695,N_41778,N_40073);
or U47696 (N_47696,N_44406,N_42856);
and U47697 (N_47697,N_44554,N_41356);
nor U47698 (N_47698,N_43013,N_42178);
nand U47699 (N_47699,N_41452,N_44097);
nor U47700 (N_47700,N_43978,N_41659);
xor U47701 (N_47701,N_42277,N_43363);
nor U47702 (N_47702,N_41426,N_42990);
xnor U47703 (N_47703,N_41246,N_44759);
xnor U47704 (N_47704,N_43861,N_43554);
nor U47705 (N_47705,N_42814,N_41751);
or U47706 (N_47706,N_40151,N_44618);
and U47707 (N_47707,N_41973,N_41022);
nor U47708 (N_47708,N_41843,N_42409);
nor U47709 (N_47709,N_44440,N_41001);
or U47710 (N_47710,N_40597,N_41292);
xnor U47711 (N_47711,N_40210,N_42580);
and U47712 (N_47712,N_43127,N_43601);
or U47713 (N_47713,N_40101,N_44212);
nand U47714 (N_47714,N_42042,N_41107);
nor U47715 (N_47715,N_43717,N_41947);
nand U47716 (N_47716,N_44480,N_44211);
xor U47717 (N_47717,N_43543,N_42689);
and U47718 (N_47718,N_42593,N_42297);
and U47719 (N_47719,N_42278,N_42630);
xnor U47720 (N_47720,N_41632,N_40340);
xor U47721 (N_47721,N_44978,N_41654);
xnor U47722 (N_47722,N_41144,N_40697);
and U47723 (N_47723,N_41331,N_43942);
nor U47724 (N_47724,N_42788,N_40007);
and U47725 (N_47725,N_40563,N_40648);
nand U47726 (N_47726,N_41170,N_43324);
nor U47727 (N_47727,N_44047,N_40574);
xnor U47728 (N_47728,N_41493,N_40934);
or U47729 (N_47729,N_43378,N_44604);
xor U47730 (N_47730,N_42599,N_44188);
and U47731 (N_47731,N_44052,N_40603);
nor U47732 (N_47732,N_44239,N_40290);
xnor U47733 (N_47733,N_42245,N_42959);
nand U47734 (N_47734,N_43806,N_41531);
and U47735 (N_47735,N_40521,N_42194);
or U47736 (N_47736,N_41466,N_42484);
nand U47737 (N_47737,N_40377,N_43531);
xor U47738 (N_47738,N_43414,N_42716);
xnor U47739 (N_47739,N_44291,N_41229);
xor U47740 (N_47740,N_40997,N_41688);
or U47741 (N_47741,N_41370,N_43575);
xor U47742 (N_47742,N_41437,N_43118);
or U47743 (N_47743,N_42926,N_40980);
and U47744 (N_47744,N_41746,N_43488);
nand U47745 (N_47745,N_44084,N_41131);
nor U47746 (N_47746,N_43981,N_40242);
xor U47747 (N_47747,N_44221,N_44954);
nand U47748 (N_47748,N_44442,N_44264);
nand U47749 (N_47749,N_42645,N_42910);
nor U47750 (N_47750,N_42560,N_43463);
xnor U47751 (N_47751,N_44206,N_42685);
and U47752 (N_47752,N_42720,N_43733);
nor U47753 (N_47753,N_44830,N_43157);
nor U47754 (N_47754,N_42498,N_41480);
xnor U47755 (N_47755,N_43472,N_41985);
nor U47756 (N_47756,N_41695,N_40089);
or U47757 (N_47757,N_40731,N_44935);
and U47758 (N_47758,N_40707,N_42409);
and U47759 (N_47759,N_43220,N_44706);
nor U47760 (N_47760,N_42165,N_40768);
and U47761 (N_47761,N_41941,N_42917);
and U47762 (N_47762,N_43654,N_41800);
xor U47763 (N_47763,N_42480,N_41965);
or U47764 (N_47764,N_44541,N_43236);
nor U47765 (N_47765,N_41791,N_43143);
nand U47766 (N_47766,N_44882,N_43820);
nand U47767 (N_47767,N_42581,N_43094);
xor U47768 (N_47768,N_41863,N_44311);
nand U47769 (N_47769,N_43117,N_44128);
and U47770 (N_47770,N_42397,N_41216);
and U47771 (N_47771,N_44732,N_43404);
xnor U47772 (N_47772,N_40956,N_40456);
nor U47773 (N_47773,N_42556,N_43223);
and U47774 (N_47774,N_42101,N_44192);
and U47775 (N_47775,N_44821,N_44060);
or U47776 (N_47776,N_42541,N_40899);
nand U47777 (N_47777,N_44480,N_42972);
nand U47778 (N_47778,N_41098,N_40818);
nand U47779 (N_47779,N_42948,N_44257);
nand U47780 (N_47780,N_42382,N_44995);
nand U47781 (N_47781,N_43534,N_43217);
xnor U47782 (N_47782,N_43832,N_41432);
xor U47783 (N_47783,N_41291,N_44266);
xor U47784 (N_47784,N_40282,N_42749);
or U47785 (N_47785,N_43687,N_43328);
xor U47786 (N_47786,N_42175,N_43578);
xor U47787 (N_47787,N_41056,N_40956);
xnor U47788 (N_47788,N_41852,N_40457);
or U47789 (N_47789,N_42829,N_44078);
xor U47790 (N_47790,N_43899,N_43534);
xor U47791 (N_47791,N_43652,N_42153);
xnor U47792 (N_47792,N_41142,N_40192);
nand U47793 (N_47793,N_44984,N_40287);
or U47794 (N_47794,N_44259,N_40866);
nor U47795 (N_47795,N_41530,N_44628);
nand U47796 (N_47796,N_42377,N_44508);
nor U47797 (N_47797,N_41625,N_44896);
or U47798 (N_47798,N_40722,N_41881);
or U47799 (N_47799,N_43124,N_41498);
and U47800 (N_47800,N_43399,N_40382);
and U47801 (N_47801,N_43556,N_42598);
and U47802 (N_47802,N_42044,N_42402);
nand U47803 (N_47803,N_44080,N_41824);
nand U47804 (N_47804,N_42340,N_40785);
nor U47805 (N_47805,N_40375,N_43577);
nor U47806 (N_47806,N_40588,N_40211);
nor U47807 (N_47807,N_42650,N_41208);
nor U47808 (N_47808,N_41804,N_41006);
and U47809 (N_47809,N_42698,N_43412);
xor U47810 (N_47810,N_41958,N_43387);
nor U47811 (N_47811,N_40207,N_42888);
or U47812 (N_47812,N_43609,N_44596);
and U47813 (N_47813,N_44000,N_43416);
nand U47814 (N_47814,N_44622,N_44375);
nor U47815 (N_47815,N_44449,N_43121);
xnor U47816 (N_47816,N_41913,N_40912);
or U47817 (N_47817,N_41073,N_43685);
xnor U47818 (N_47818,N_41638,N_41525);
and U47819 (N_47819,N_41430,N_43519);
xor U47820 (N_47820,N_44048,N_41039);
or U47821 (N_47821,N_40840,N_42506);
or U47822 (N_47822,N_41612,N_41570);
and U47823 (N_47823,N_40789,N_42918);
xor U47824 (N_47824,N_44031,N_44819);
xnor U47825 (N_47825,N_41678,N_43608);
and U47826 (N_47826,N_42894,N_44844);
nand U47827 (N_47827,N_44962,N_44610);
or U47828 (N_47828,N_41396,N_41755);
and U47829 (N_47829,N_41225,N_40969);
nor U47830 (N_47830,N_41302,N_43113);
and U47831 (N_47831,N_40937,N_40917);
nor U47832 (N_47832,N_40760,N_42619);
nand U47833 (N_47833,N_41900,N_40841);
or U47834 (N_47834,N_43263,N_41885);
and U47835 (N_47835,N_40860,N_40738);
nor U47836 (N_47836,N_41954,N_43125);
nor U47837 (N_47837,N_42535,N_44249);
nor U47838 (N_47838,N_44463,N_43611);
xnor U47839 (N_47839,N_44179,N_40520);
and U47840 (N_47840,N_43234,N_44914);
and U47841 (N_47841,N_41771,N_42950);
nand U47842 (N_47842,N_42747,N_40311);
nor U47843 (N_47843,N_42543,N_40585);
nor U47844 (N_47844,N_43321,N_42062);
xor U47845 (N_47845,N_40723,N_41739);
nor U47846 (N_47846,N_44310,N_41357);
nor U47847 (N_47847,N_44908,N_43144);
nor U47848 (N_47848,N_43577,N_44448);
nor U47849 (N_47849,N_43971,N_43703);
or U47850 (N_47850,N_44206,N_42987);
nor U47851 (N_47851,N_40730,N_43021);
and U47852 (N_47852,N_41264,N_43810);
xnor U47853 (N_47853,N_43263,N_41468);
xnor U47854 (N_47854,N_41439,N_43731);
xor U47855 (N_47855,N_43314,N_42164);
nor U47856 (N_47856,N_41299,N_40333);
or U47857 (N_47857,N_43231,N_43396);
nand U47858 (N_47858,N_40425,N_44502);
and U47859 (N_47859,N_42106,N_42008);
nor U47860 (N_47860,N_43498,N_43719);
nand U47861 (N_47861,N_42809,N_44408);
nand U47862 (N_47862,N_41422,N_42417);
or U47863 (N_47863,N_40589,N_42577);
xor U47864 (N_47864,N_42283,N_44860);
nor U47865 (N_47865,N_44164,N_42249);
xnor U47866 (N_47866,N_42946,N_42123);
nand U47867 (N_47867,N_43604,N_44821);
xor U47868 (N_47868,N_40701,N_41212);
and U47869 (N_47869,N_41745,N_43840);
nand U47870 (N_47870,N_40539,N_40397);
nor U47871 (N_47871,N_43277,N_44011);
nor U47872 (N_47872,N_43871,N_40106);
or U47873 (N_47873,N_41787,N_42927);
and U47874 (N_47874,N_44448,N_42903);
nand U47875 (N_47875,N_42911,N_40060);
nand U47876 (N_47876,N_43618,N_41945);
or U47877 (N_47877,N_43745,N_43008);
nor U47878 (N_47878,N_44878,N_44240);
nor U47879 (N_47879,N_44928,N_43016);
or U47880 (N_47880,N_43179,N_41438);
and U47881 (N_47881,N_42310,N_44354);
nor U47882 (N_47882,N_41325,N_44175);
xnor U47883 (N_47883,N_42760,N_40050);
nor U47884 (N_47884,N_40910,N_40438);
or U47885 (N_47885,N_40044,N_41854);
and U47886 (N_47886,N_42591,N_42222);
or U47887 (N_47887,N_43277,N_43039);
or U47888 (N_47888,N_43469,N_44753);
and U47889 (N_47889,N_42272,N_41776);
nor U47890 (N_47890,N_44401,N_42858);
nor U47891 (N_47891,N_44027,N_43883);
nand U47892 (N_47892,N_41841,N_40456);
xor U47893 (N_47893,N_40801,N_41443);
nand U47894 (N_47894,N_44000,N_42290);
and U47895 (N_47895,N_44079,N_42468);
or U47896 (N_47896,N_43041,N_42523);
or U47897 (N_47897,N_40483,N_42287);
or U47898 (N_47898,N_40204,N_43154);
nor U47899 (N_47899,N_43174,N_43653);
nand U47900 (N_47900,N_44658,N_40182);
nor U47901 (N_47901,N_41794,N_43848);
and U47902 (N_47902,N_43364,N_41716);
and U47903 (N_47903,N_41544,N_40551);
nor U47904 (N_47904,N_44712,N_40275);
and U47905 (N_47905,N_42245,N_40079);
nand U47906 (N_47906,N_40373,N_42273);
or U47907 (N_47907,N_43856,N_41210);
nand U47908 (N_47908,N_42500,N_44113);
nor U47909 (N_47909,N_40468,N_40133);
nand U47910 (N_47910,N_43314,N_41750);
and U47911 (N_47911,N_40745,N_43627);
nor U47912 (N_47912,N_41292,N_40898);
nand U47913 (N_47913,N_43152,N_42657);
and U47914 (N_47914,N_40248,N_44466);
nor U47915 (N_47915,N_40416,N_44436);
nor U47916 (N_47916,N_42699,N_42253);
or U47917 (N_47917,N_41238,N_43046);
xnor U47918 (N_47918,N_43684,N_40467);
nand U47919 (N_47919,N_43922,N_42592);
xor U47920 (N_47920,N_40391,N_40473);
and U47921 (N_47921,N_41705,N_40517);
nor U47922 (N_47922,N_41391,N_44319);
xor U47923 (N_47923,N_43343,N_44113);
xor U47924 (N_47924,N_40983,N_42237);
or U47925 (N_47925,N_41018,N_43650);
nor U47926 (N_47926,N_40288,N_44121);
xor U47927 (N_47927,N_44359,N_41621);
and U47928 (N_47928,N_42433,N_44608);
or U47929 (N_47929,N_41479,N_40275);
or U47930 (N_47930,N_40355,N_41900);
or U47931 (N_47931,N_42486,N_41709);
and U47932 (N_47932,N_41582,N_43764);
xor U47933 (N_47933,N_44718,N_43894);
nor U47934 (N_47934,N_40993,N_40792);
nor U47935 (N_47935,N_42850,N_42327);
and U47936 (N_47936,N_42936,N_41325);
nand U47937 (N_47937,N_44653,N_42600);
nor U47938 (N_47938,N_44143,N_43362);
and U47939 (N_47939,N_42358,N_41661);
or U47940 (N_47940,N_43469,N_40139);
or U47941 (N_47941,N_41406,N_41819);
and U47942 (N_47942,N_43174,N_44690);
and U47943 (N_47943,N_41355,N_44574);
xor U47944 (N_47944,N_44247,N_41631);
and U47945 (N_47945,N_41988,N_42333);
xor U47946 (N_47946,N_40491,N_41902);
nand U47947 (N_47947,N_44301,N_44501);
xnor U47948 (N_47948,N_44252,N_44930);
and U47949 (N_47949,N_43155,N_41734);
nor U47950 (N_47950,N_40538,N_44005);
nor U47951 (N_47951,N_44964,N_44245);
nor U47952 (N_47952,N_42056,N_44281);
xor U47953 (N_47953,N_41047,N_41952);
nand U47954 (N_47954,N_40110,N_41863);
nor U47955 (N_47955,N_42751,N_44354);
xnor U47956 (N_47956,N_40044,N_42340);
or U47957 (N_47957,N_41811,N_42618);
nand U47958 (N_47958,N_44815,N_44711);
or U47959 (N_47959,N_43831,N_44341);
nand U47960 (N_47960,N_43182,N_42360);
and U47961 (N_47961,N_41024,N_40033);
nand U47962 (N_47962,N_42857,N_43763);
and U47963 (N_47963,N_40329,N_43067);
or U47964 (N_47964,N_42201,N_43793);
or U47965 (N_47965,N_40596,N_44205);
xor U47966 (N_47966,N_41466,N_40023);
or U47967 (N_47967,N_44856,N_44590);
nor U47968 (N_47968,N_43264,N_41216);
xnor U47969 (N_47969,N_43277,N_43174);
nand U47970 (N_47970,N_41924,N_43656);
and U47971 (N_47971,N_42119,N_40343);
xor U47972 (N_47972,N_40143,N_42530);
and U47973 (N_47973,N_43633,N_41019);
xor U47974 (N_47974,N_44342,N_43927);
nand U47975 (N_47975,N_42627,N_43915);
nand U47976 (N_47976,N_41275,N_41968);
or U47977 (N_47977,N_43074,N_42450);
nand U47978 (N_47978,N_43746,N_42510);
and U47979 (N_47979,N_40965,N_40517);
xor U47980 (N_47980,N_41893,N_41026);
xnor U47981 (N_47981,N_44796,N_43775);
nor U47982 (N_47982,N_41036,N_43878);
xnor U47983 (N_47983,N_43963,N_44090);
and U47984 (N_47984,N_41015,N_41679);
or U47985 (N_47985,N_42778,N_43145);
nor U47986 (N_47986,N_42505,N_41885);
nand U47987 (N_47987,N_41743,N_42426);
and U47988 (N_47988,N_41685,N_43834);
nand U47989 (N_47989,N_43928,N_44326);
nand U47990 (N_47990,N_44546,N_43463);
and U47991 (N_47991,N_42534,N_40571);
nand U47992 (N_47992,N_42522,N_40554);
and U47993 (N_47993,N_44985,N_44169);
or U47994 (N_47994,N_40190,N_44918);
or U47995 (N_47995,N_44222,N_40477);
or U47996 (N_47996,N_40896,N_42574);
nand U47997 (N_47997,N_43228,N_42177);
nand U47998 (N_47998,N_41262,N_42189);
and U47999 (N_47999,N_40915,N_44016);
xor U48000 (N_48000,N_43693,N_43438);
nor U48001 (N_48001,N_40626,N_44169);
nor U48002 (N_48002,N_42202,N_42034);
xnor U48003 (N_48003,N_40425,N_42974);
xor U48004 (N_48004,N_41166,N_40637);
nand U48005 (N_48005,N_40947,N_43573);
nand U48006 (N_48006,N_41144,N_40896);
xor U48007 (N_48007,N_42664,N_40429);
nor U48008 (N_48008,N_44293,N_44964);
xor U48009 (N_48009,N_44056,N_43272);
nor U48010 (N_48010,N_43378,N_41420);
nand U48011 (N_48011,N_41291,N_41089);
xnor U48012 (N_48012,N_40723,N_41935);
nand U48013 (N_48013,N_42110,N_40375);
or U48014 (N_48014,N_43109,N_44306);
or U48015 (N_48015,N_44268,N_41289);
xnor U48016 (N_48016,N_40705,N_42573);
xor U48017 (N_48017,N_42377,N_43189);
and U48018 (N_48018,N_41320,N_42994);
nor U48019 (N_48019,N_42718,N_44342);
nor U48020 (N_48020,N_43204,N_40844);
or U48021 (N_48021,N_42358,N_44077);
or U48022 (N_48022,N_40880,N_43687);
or U48023 (N_48023,N_41710,N_43196);
nor U48024 (N_48024,N_42765,N_43484);
or U48025 (N_48025,N_42680,N_40898);
or U48026 (N_48026,N_44836,N_43568);
nand U48027 (N_48027,N_44866,N_44137);
or U48028 (N_48028,N_43163,N_43363);
nor U48029 (N_48029,N_40742,N_42462);
xor U48030 (N_48030,N_42111,N_40793);
xnor U48031 (N_48031,N_44170,N_42814);
or U48032 (N_48032,N_41152,N_42116);
nand U48033 (N_48033,N_44363,N_44615);
xnor U48034 (N_48034,N_44155,N_42522);
and U48035 (N_48035,N_43664,N_42396);
nand U48036 (N_48036,N_43234,N_42874);
nand U48037 (N_48037,N_40275,N_41180);
or U48038 (N_48038,N_42325,N_41503);
and U48039 (N_48039,N_42579,N_41111);
xor U48040 (N_48040,N_44173,N_41164);
nand U48041 (N_48041,N_41206,N_41510);
nor U48042 (N_48042,N_40022,N_40070);
nor U48043 (N_48043,N_44269,N_42558);
nand U48044 (N_48044,N_44793,N_40509);
nand U48045 (N_48045,N_41353,N_43752);
xnor U48046 (N_48046,N_40776,N_43891);
or U48047 (N_48047,N_44802,N_41684);
or U48048 (N_48048,N_41214,N_40327);
or U48049 (N_48049,N_44019,N_40459);
nand U48050 (N_48050,N_40808,N_44903);
or U48051 (N_48051,N_44052,N_43330);
xor U48052 (N_48052,N_42114,N_40125);
nor U48053 (N_48053,N_42442,N_40050);
xor U48054 (N_48054,N_43053,N_41846);
or U48055 (N_48055,N_43632,N_42898);
or U48056 (N_48056,N_41421,N_44282);
and U48057 (N_48057,N_41671,N_41384);
or U48058 (N_48058,N_43506,N_43316);
or U48059 (N_48059,N_44764,N_40207);
or U48060 (N_48060,N_43488,N_40674);
xnor U48061 (N_48061,N_42737,N_40568);
xnor U48062 (N_48062,N_40951,N_44799);
nor U48063 (N_48063,N_43188,N_42467);
xor U48064 (N_48064,N_43323,N_40168);
nand U48065 (N_48065,N_40927,N_41498);
xor U48066 (N_48066,N_41552,N_41550);
nand U48067 (N_48067,N_40602,N_40042);
nor U48068 (N_48068,N_42924,N_41897);
and U48069 (N_48069,N_41626,N_41908);
and U48070 (N_48070,N_40251,N_41775);
or U48071 (N_48071,N_43659,N_43768);
and U48072 (N_48072,N_43272,N_40620);
nor U48073 (N_48073,N_43742,N_41459);
or U48074 (N_48074,N_41711,N_40469);
nor U48075 (N_48075,N_40003,N_40854);
nand U48076 (N_48076,N_44240,N_42756);
and U48077 (N_48077,N_44286,N_44214);
or U48078 (N_48078,N_41729,N_40506);
nor U48079 (N_48079,N_43869,N_42750);
or U48080 (N_48080,N_44198,N_41228);
nor U48081 (N_48081,N_41447,N_42585);
nand U48082 (N_48082,N_42079,N_40566);
xnor U48083 (N_48083,N_42546,N_42621);
and U48084 (N_48084,N_40437,N_42349);
nor U48085 (N_48085,N_41847,N_41476);
xor U48086 (N_48086,N_42747,N_41176);
nand U48087 (N_48087,N_40590,N_41146);
xor U48088 (N_48088,N_44210,N_43116);
and U48089 (N_48089,N_41880,N_41008);
nor U48090 (N_48090,N_41310,N_43264);
nor U48091 (N_48091,N_42467,N_42574);
or U48092 (N_48092,N_41915,N_41340);
and U48093 (N_48093,N_41747,N_40958);
and U48094 (N_48094,N_44262,N_40651);
and U48095 (N_48095,N_43011,N_41593);
nand U48096 (N_48096,N_41181,N_43384);
nand U48097 (N_48097,N_43465,N_43858);
nand U48098 (N_48098,N_40301,N_40243);
nor U48099 (N_48099,N_41313,N_41290);
xor U48100 (N_48100,N_43654,N_41243);
and U48101 (N_48101,N_41101,N_41980);
or U48102 (N_48102,N_41862,N_41080);
nor U48103 (N_48103,N_41333,N_42042);
or U48104 (N_48104,N_40585,N_42710);
or U48105 (N_48105,N_41901,N_44763);
or U48106 (N_48106,N_44347,N_42452);
nor U48107 (N_48107,N_42979,N_44110);
or U48108 (N_48108,N_40770,N_44912);
nand U48109 (N_48109,N_41566,N_42670);
or U48110 (N_48110,N_40605,N_40684);
nor U48111 (N_48111,N_43417,N_41627);
or U48112 (N_48112,N_42134,N_42345);
nand U48113 (N_48113,N_43933,N_44358);
and U48114 (N_48114,N_40986,N_42754);
nor U48115 (N_48115,N_41243,N_43168);
nand U48116 (N_48116,N_40263,N_42940);
nor U48117 (N_48117,N_42131,N_42352);
or U48118 (N_48118,N_40199,N_41864);
xor U48119 (N_48119,N_42790,N_41941);
nand U48120 (N_48120,N_42923,N_43669);
nand U48121 (N_48121,N_41789,N_44573);
or U48122 (N_48122,N_40416,N_44905);
and U48123 (N_48123,N_43475,N_44091);
or U48124 (N_48124,N_41129,N_42262);
nand U48125 (N_48125,N_42151,N_40722);
nor U48126 (N_48126,N_44855,N_41361);
nand U48127 (N_48127,N_40390,N_42172);
xor U48128 (N_48128,N_42927,N_43134);
and U48129 (N_48129,N_43926,N_41455);
xnor U48130 (N_48130,N_40642,N_40209);
xnor U48131 (N_48131,N_44617,N_43786);
nand U48132 (N_48132,N_43216,N_42686);
nand U48133 (N_48133,N_41229,N_41436);
xnor U48134 (N_48134,N_42376,N_44952);
nand U48135 (N_48135,N_41865,N_42294);
or U48136 (N_48136,N_42445,N_41668);
nand U48137 (N_48137,N_41506,N_41289);
nor U48138 (N_48138,N_44937,N_40217);
nand U48139 (N_48139,N_40665,N_44595);
nor U48140 (N_48140,N_43746,N_41202);
or U48141 (N_48141,N_41848,N_40896);
nand U48142 (N_48142,N_40626,N_41164);
nor U48143 (N_48143,N_42796,N_40973);
nor U48144 (N_48144,N_41889,N_43222);
nand U48145 (N_48145,N_42916,N_44476);
xor U48146 (N_48146,N_41055,N_42387);
or U48147 (N_48147,N_44911,N_44784);
nor U48148 (N_48148,N_43871,N_43188);
xor U48149 (N_48149,N_40771,N_43964);
xnor U48150 (N_48150,N_43328,N_43910);
or U48151 (N_48151,N_44450,N_42949);
or U48152 (N_48152,N_43606,N_44810);
nand U48153 (N_48153,N_44888,N_44203);
or U48154 (N_48154,N_42178,N_43813);
xnor U48155 (N_48155,N_41653,N_41576);
nand U48156 (N_48156,N_42444,N_40378);
xor U48157 (N_48157,N_42301,N_42844);
xnor U48158 (N_48158,N_42233,N_41801);
and U48159 (N_48159,N_43013,N_43185);
nor U48160 (N_48160,N_43941,N_44888);
nor U48161 (N_48161,N_44275,N_44121);
xnor U48162 (N_48162,N_43627,N_42598);
xnor U48163 (N_48163,N_43781,N_41669);
xnor U48164 (N_48164,N_42526,N_44860);
xor U48165 (N_48165,N_42882,N_40697);
nor U48166 (N_48166,N_40561,N_42627);
xor U48167 (N_48167,N_41515,N_44553);
nand U48168 (N_48168,N_41726,N_41300);
and U48169 (N_48169,N_44437,N_44483);
and U48170 (N_48170,N_41772,N_42739);
or U48171 (N_48171,N_41150,N_40552);
nor U48172 (N_48172,N_42816,N_41864);
xnor U48173 (N_48173,N_40025,N_44113);
or U48174 (N_48174,N_42922,N_44026);
nor U48175 (N_48175,N_44732,N_40424);
or U48176 (N_48176,N_43255,N_42874);
or U48177 (N_48177,N_41717,N_43885);
xnor U48178 (N_48178,N_44682,N_44923);
nor U48179 (N_48179,N_42734,N_42867);
or U48180 (N_48180,N_43172,N_41249);
nor U48181 (N_48181,N_41203,N_44738);
nor U48182 (N_48182,N_44630,N_43889);
or U48183 (N_48183,N_40355,N_40023);
or U48184 (N_48184,N_44612,N_42591);
xnor U48185 (N_48185,N_43202,N_43372);
nor U48186 (N_48186,N_44886,N_40234);
or U48187 (N_48187,N_42595,N_44851);
or U48188 (N_48188,N_43036,N_41209);
nor U48189 (N_48189,N_40517,N_41308);
nor U48190 (N_48190,N_43005,N_42772);
and U48191 (N_48191,N_41380,N_40270);
nor U48192 (N_48192,N_43537,N_42384);
nand U48193 (N_48193,N_43698,N_42965);
or U48194 (N_48194,N_41121,N_44040);
nand U48195 (N_48195,N_44859,N_40598);
xnor U48196 (N_48196,N_44073,N_43471);
xnor U48197 (N_48197,N_41933,N_44369);
or U48198 (N_48198,N_42818,N_40620);
nand U48199 (N_48199,N_43789,N_43022);
nor U48200 (N_48200,N_44520,N_44430);
and U48201 (N_48201,N_43838,N_41232);
or U48202 (N_48202,N_43197,N_43437);
and U48203 (N_48203,N_41151,N_40698);
and U48204 (N_48204,N_43868,N_43633);
nor U48205 (N_48205,N_40820,N_42703);
nor U48206 (N_48206,N_40234,N_42462);
or U48207 (N_48207,N_43016,N_40159);
nand U48208 (N_48208,N_43807,N_43992);
nor U48209 (N_48209,N_43316,N_40971);
xnor U48210 (N_48210,N_41752,N_43840);
and U48211 (N_48211,N_44703,N_43613);
and U48212 (N_48212,N_42709,N_44825);
or U48213 (N_48213,N_43564,N_41540);
nor U48214 (N_48214,N_42204,N_42939);
xor U48215 (N_48215,N_44345,N_41657);
xor U48216 (N_48216,N_40022,N_41945);
or U48217 (N_48217,N_42658,N_41444);
nor U48218 (N_48218,N_44635,N_40316);
nor U48219 (N_48219,N_43521,N_43385);
nand U48220 (N_48220,N_40452,N_43264);
nand U48221 (N_48221,N_41002,N_40726);
xnor U48222 (N_48222,N_43865,N_44975);
xor U48223 (N_48223,N_43197,N_41665);
nor U48224 (N_48224,N_41958,N_44234);
or U48225 (N_48225,N_40050,N_44806);
nor U48226 (N_48226,N_44755,N_44112);
xor U48227 (N_48227,N_42911,N_40269);
or U48228 (N_48228,N_43865,N_44257);
or U48229 (N_48229,N_43604,N_42814);
or U48230 (N_48230,N_44476,N_40120);
nor U48231 (N_48231,N_44710,N_44962);
xnor U48232 (N_48232,N_41454,N_43879);
or U48233 (N_48233,N_43133,N_42640);
nand U48234 (N_48234,N_44983,N_43426);
nor U48235 (N_48235,N_40990,N_41725);
xor U48236 (N_48236,N_40080,N_41361);
nor U48237 (N_48237,N_44676,N_43626);
and U48238 (N_48238,N_44481,N_42380);
nor U48239 (N_48239,N_42928,N_44130);
and U48240 (N_48240,N_42401,N_41490);
nor U48241 (N_48241,N_42332,N_42862);
and U48242 (N_48242,N_42718,N_42389);
and U48243 (N_48243,N_42308,N_40577);
and U48244 (N_48244,N_44372,N_41082);
nor U48245 (N_48245,N_40138,N_44598);
and U48246 (N_48246,N_41225,N_43920);
and U48247 (N_48247,N_44228,N_43927);
and U48248 (N_48248,N_41968,N_43379);
nand U48249 (N_48249,N_44290,N_41640);
nor U48250 (N_48250,N_43491,N_40428);
or U48251 (N_48251,N_42692,N_42891);
or U48252 (N_48252,N_44370,N_41053);
or U48253 (N_48253,N_40928,N_43000);
nor U48254 (N_48254,N_44735,N_41237);
and U48255 (N_48255,N_42918,N_44674);
nand U48256 (N_48256,N_44683,N_40561);
nand U48257 (N_48257,N_43391,N_42915);
xor U48258 (N_48258,N_43073,N_44911);
xor U48259 (N_48259,N_43274,N_40892);
and U48260 (N_48260,N_40799,N_42134);
xor U48261 (N_48261,N_43401,N_42132);
xnor U48262 (N_48262,N_41528,N_42557);
nand U48263 (N_48263,N_40364,N_44371);
and U48264 (N_48264,N_42973,N_43581);
or U48265 (N_48265,N_43858,N_40065);
nor U48266 (N_48266,N_42963,N_42611);
nand U48267 (N_48267,N_40483,N_40574);
or U48268 (N_48268,N_44063,N_42460);
nor U48269 (N_48269,N_40913,N_40103);
nor U48270 (N_48270,N_41609,N_40830);
or U48271 (N_48271,N_43792,N_41373);
nand U48272 (N_48272,N_42649,N_40873);
nor U48273 (N_48273,N_42412,N_40359);
xor U48274 (N_48274,N_41138,N_44091);
nand U48275 (N_48275,N_40152,N_44794);
nand U48276 (N_48276,N_40177,N_41727);
xor U48277 (N_48277,N_41428,N_44263);
xor U48278 (N_48278,N_43435,N_43026);
or U48279 (N_48279,N_40289,N_41284);
or U48280 (N_48280,N_43086,N_44198);
xor U48281 (N_48281,N_43569,N_43419);
nor U48282 (N_48282,N_42271,N_41200);
or U48283 (N_48283,N_41298,N_42986);
nand U48284 (N_48284,N_42375,N_41136);
or U48285 (N_48285,N_40098,N_43980);
nor U48286 (N_48286,N_40621,N_41130);
nand U48287 (N_48287,N_41323,N_42773);
xor U48288 (N_48288,N_40691,N_42052);
xor U48289 (N_48289,N_42560,N_44048);
nand U48290 (N_48290,N_44175,N_40789);
and U48291 (N_48291,N_42296,N_42102);
nand U48292 (N_48292,N_41317,N_40061);
or U48293 (N_48293,N_44124,N_43746);
and U48294 (N_48294,N_44638,N_41011);
nand U48295 (N_48295,N_41750,N_44818);
and U48296 (N_48296,N_44195,N_44223);
nor U48297 (N_48297,N_42332,N_44528);
and U48298 (N_48298,N_44442,N_42326);
or U48299 (N_48299,N_42084,N_43151);
xor U48300 (N_48300,N_44698,N_43164);
xnor U48301 (N_48301,N_41378,N_40530);
nor U48302 (N_48302,N_42760,N_44570);
xnor U48303 (N_48303,N_42102,N_43599);
or U48304 (N_48304,N_43721,N_40370);
or U48305 (N_48305,N_42394,N_42437);
or U48306 (N_48306,N_43021,N_41067);
or U48307 (N_48307,N_40038,N_44367);
xor U48308 (N_48308,N_43241,N_41420);
and U48309 (N_48309,N_41742,N_41018);
xnor U48310 (N_48310,N_43376,N_44129);
and U48311 (N_48311,N_42649,N_42194);
xor U48312 (N_48312,N_43737,N_42725);
or U48313 (N_48313,N_41094,N_40401);
nand U48314 (N_48314,N_42287,N_44094);
or U48315 (N_48315,N_40955,N_42103);
nand U48316 (N_48316,N_43226,N_43784);
nand U48317 (N_48317,N_42841,N_43318);
nand U48318 (N_48318,N_44667,N_41226);
and U48319 (N_48319,N_40053,N_42402);
nand U48320 (N_48320,N_42819,N_43715);
nand U48321 (N_48321,N_44593,N_40960);
nand U48322 (N_48322,N_44423,N_43553);
nand U48323 (N_48323,N_41788,N_43025);
xnor U48324 (N_48324,N_40283,N_42406);
nor U48325 (N_48325,N_44739,N_43019);
nand U48326 (N_48326,N_41884,N_40807);
nand U48327 (N_48327,N_42786,N_40752);
or U48328 (N_48328,N_42021,N_42252);
nor U48329 (N_48329,N_43238,N_43703);
and U48330 (N_48330,N_42922,N_43191);
nor U48331 (N_48331,N_41119,N_40813);
or U48332 (N_48332,N_42171,N_43789);
xnor U48333 (N_48333,N_43344,N_42486);
or U48334 (N_48334,N_41296,N_40961);
or U48335 (N_48335,N_41684,N_42184);
nand U48336 (N_48336,N_44715,N_40055);
and U48337 (N_48337,N_44125,N_42320);
or U48338 (N_48338,N_44409,N_40659);
nor U48339 (N_48339,N_44639,N_44679);
and U48340 (N_48340,N_44874,N_40227);
and U48341 (N_48341,N_42992,N_40606);
xnor U48342 (N_48342,N_43050,N_41478);
nor U48343 (N_48343,N_44518,N_43912);
or U48344 (N_48344,N_41710,N_42696);
or U48345 (N_48345,N_43465,N_40848);
and U48346 (N_48346,N_44930,N_42773);
and U48347 (N_48347,N_43091,N_42622);
nor U48348 (N_48348,N_43490,N_41676);
nor U48349 (N_48349,N_44997,N_44698);
or U48350 (N_48350,N_44973,N_43658);
nand U48351 (N_48351,N_44291,N_40458);
or U48352 (N_48352,N_41205,N_42812);
or U48353 (N_48353,N_42939,N_42130);
nand U48354 (N_48354,N_41148,N_42936);
or U48355 (N_48355,N_41562,N_41522);
and U48356 (N_48356,N_43186,N_42671);
nand U48357 (N_48357,N_40105,N_44871);
or U48358 (N_48358,N_42192,N_44001);
nor U48359 (N_48359,N_42209,N_41819);
and U48360 (N_48360,N_43924,N_43950);
and U48361 (N_48361,N_44264,N_42449);
or U48362 (N_48362,N_42857,N_41398);
nor U48363 (N_48363,N_40636,N_40126);
nand U48364 (N_48364,N_42820,N_40097);
xor U48365 (N_48365,N_44426,N_44694);
nor U48366 (N_48366,N_43020,N_41762);
nand U48367 (N_48367,N_44613,N_42756);
xnor U48368 (N_48368,N_44882,N_43410);
or U48369 (N_48369,N_40440,N_42694);
nor U48370 (N_48370,N_43451,N_44297);
or U48371 (N_48371,N_44737,N_43047);
or U48372 (N_48372,N_41118,N_40074);
nor U48373 (N_48373,N_44795,N_42377);
nor U48374 (N_48374,N_43353,N_44830);
nor U48375 (N_48375,N_44153,N_43611);
or U48376 (N_48376,N_43718,N_40990);
xnor U48377 (N_48377,N_44357,N_41309);
nor U48378 (N_48378,N_40654,N_44467);
xor U48379 (N_48379,N_41196,N_43480);
and U48380 (N_48380,N_40122,N_41921);
or U48381 (N_48381,N_44451,N_43092);
nand U48382 (N_48382,N_41817,N_41692);
and U48383 (N_48383,N_41946,N_43606);
or U48384 (N_48384,N_44324,N_43667);
xor U48385 (N_48385,N_43446,N_41655);
nand U48386 (N_48386,N_41563,N_40308);
nor U48387 (N_48387,N_40435,N_41211);
nor U48388 (N_48388,N_44290,N_42937);
xor U48389 (N_48389,N_43270,N_41633);
nor U48390 (N_48390,N_43602,N_44689);
or U48391 (N_48391,N_43142,N_40399);
nor U48392 (N_48392,N_42246,N_42411);
xnor U48393 (N_48393,N_40132,N_43879);
or U48394 (N_48394,N_41632,N_43010);
or U48395 (N_48395,N_42724,N_41934);
nand U48396 (N_48396,N_43287,N_42678);
or U48397 (N_48397,N_43812,N_40927);
nor U48398 (N_48398,N_40389,N_43511);
xnor U48399 (N_48399,N_41561,N_43228);
nand U48400 (N_48400,N_44720,N_40690);
or U48401 (N_48401,N_43697,N_41163);
xnor U48402 (N_48402,N_44743,N_40379);
xor U48403 (N_48403,N_44946,N_43185);
and U48404 (N_48404,N_41016,N_40210);
nand U48405 (N_48405,N_41171,N_44912);
and U48406 (N_48406,N_44351,N_43903);
nand U48407 (N_48407,N_40136,N_40141);
nand U48408 (N_48408,N_42371,N_43459);
and U48409 (N_48409,N_43864,N_44246);
nand U48410 (N_48410,N_41182,N_42768);
xor U48411 (N_48411,N_43342,N_43223);
nor U48412 (N_48412,N_40782,N_41012);
and U48413 (N_48413,N_40081,N_40306);
and U48414 (N_48414,N_44370,N_44733);
xor U48415 (N_48415,N_40413,N_43678);
nor U48416 (N_48416,N_43104,N_41122);
nand U48417 (N_48417,N_43528,N_41445);
nand U48418 (N_48418,N_41790,N_43090);
xor U48419 (N_48419,N_40264,N_43218);
nor U48420 (N_48420,N_40213,N_43418);
nand U48421 (N_48421,N_43259,N_44528);
nor U48422 (N_48422,N_40685,N_42388);
xor U48423 (N_48423,N_44204,N_41560);
nor U48424 (N_48424,N_41265,N_40945);
and U48425 (N_48425,N_40191,N_41504);
nand U48426 (N_48426,N_42221,N_41794);
or U48427 (N_48427,N_42454,N_40957);
and U48428 (N_48428,N_42219,N_41167);
nand U48429 (N_48429,N_44683,N_44006);
nand U48430 (N_48430,N_41403,N_44955);
or U48431 (N_48431,N_44431,N_44549);
or U48432 (N_48432,N_40814,N_42434);
xnor U48433 (N_48433,N_43647,N_40516);
and U48434 (N_48434,N_41419,N_42422);
and U48435 (N_48435,N_42024,N_41331);
and U48436 (N_48436,N_41398,N_44614);
xor U48437 (N_48437,N_44266,N_42830);
or U48438 (N_48438,N_44446,N_41430);
and U48439 (N_48439,N_43021,N_40499);
nor U48440 (N_48440,N_41738,N_44861);
nand U48441 (N_48441,N_41684,N_40812);
nand U48442 (N_48442,N_44297,N_44607);
nor U48443 (N_48443,N_44870,N_40214);
nor U48444 (N_48444,N_40393,N_40307);
nand U48445 (N_48445,N_42577,N_44815);
nor U48446 (N_48446,N_44181,N_43100);
nand U48447 (N_48447,N_41187,N_43285);
or U48448 (N_48448,N_41172,N_44481);
or U48449 (N_48449,N_42544,N_40202);
and U48450 (N_48450,N_43866,N_42155);
xnor U48451 (N_48451,N_42806,N_40397);
nand U48452 (N_48452,N_44697,N_42328);
or U48453 (N_48453,N_42946,N_42707);
and U48454 (N_48454,N_43910,N_40752);
or U48455 (N_48455,N_42990,N_42910);
and U48456 (N_48456,N_41766,N_44803);
or U48457 (N_48457,N_41621,N_41559);
nor U48458 (N_48458,N_41568,N_44357);
xor U48459 (N_48459,N_43590,N_43048);
nor U48460 (N_48460,N_42251,N_44237);
xor U48461 (N_48461,N_42145,N_40996);
nor U48462 (N_48462,N_43291,N_40742);
nor U48463 (N_48463,N_44066,N_42590);
nor U48464 (N_48464,N_43017,N_44572);
nor U48465 (N_48465,N_40232,N_44203);
nor U48466 (N_48466,N_40280,N_40758);
nor U48467 (N_48467,N_42438,N_41682);
xor U48468 (N_48468,N_44440,N_40944);
and U48469 (N_48469,N_40883,N_41833);
xnor U48470 (N_48470,N_44602,N_42419);
xor U48471 (N_48471,N_40405,N_44003);
nor U48472 (N_48472,N_43709,N_44564);
xnor U48473 (N_48473,N_41580,N_44632);
or U48474 (N_48474,N_44662,N_42098);
xnor U48475 (N_48475,N_40775,N_44070);
nor U48476 (N_48476,N_44679,N_40608);
nor U48477 (N_48477,N_44322,N_43257);
nor U48478 (N_48478,N_41203,N_44015);
or U48479 (N_48479,N_44426,N_40288);
or U48480 (N_48480,N_43565,N_44022);
nor U48481 (N_48481,N_43927,N_43010);
and U48482 (N_48482,N_43562,N_44951);
and U48483 (N_48483,N_42171,N_42183);
nand U48484 (N_48484,N_41928,N_44962);
nor U48485 (N_48485,N_44840,N_44931);
and U48486 (N_48486,N_42421,N_40601);
nand U48487 (N_48487,N_43779,N_42873);
nand U48488 (N_48488,N_42059,N_40020);
nand U48489 (N_48489,N_42604,N_41670);
nand U48490 (N_48490,N_43600,N_43444);
or U48491 (N_48491,N_43310,N_42308);
and U48492 (N_48492,N_40411,N_42987);
xnor U48493 (N_48493,N_43804,N_41606);
and U48494 (N_48494,N_42608,N_43414);
nor U48495 (N_48495,N_40032,N_41472);
nor U48496 (N_48496,N_43332,N_44735);
xor U48497 (N_48497,N_41716,N_42959);
or U48498 (N_48498,N_40026,N_40220);
xor U48499 (N_48499,N_42240,N_42128);
and U48500 (N_48500,N_44575,N_42356);
and U48501 (N_48501,N_43708,N_44079);
xnor U48502 (N_48502,N_42000,N_40266);
nand U48503 (N_48503,N_40783,N_43761);
and U48504 (N_48504,N_40175,N_41735);
and U48505 (N_48505,N_41150,N_44865);
or U48506 (N_48506,N_42695,N_44366);
and U48507 (N_48507,N_40309,N_40468);
nand U48508 (N_48508,N_42009,N_42592);
and U48509 (N_48509,N_40544,N_41845);
xnor U48510 (N_48510,N_44573,N_41121);
nor U48511 (N_48511,N_42556,N_41803);
xor U48512 (N_48512,N_44956,N_44979);
xnor U48513 (N_48513,N_40613,N_44342);
xor U48514 (N_48514,N_44438,N_41824);
or U48515 (N_48515,N_42676,N_42931);
nor U48516 (N_48516,N_41999,N_40910);
nand U48517 (N_48517,N_44048,N_40475);
and U48518 (N_48518,N_41550,N_41774);
nand U48519 (N_48519,N_41196,N_41739);
xnor U48520 (N_48520,N_43198,N_42040);
xnor U48521 (N_48521,N_44172,N_41858);
nand U48522 (N_48522,N_44490,N_44977);
nor U48523 (N_48523,N_42792,N_44863);
and U48524 (N_48524,N_41450,N_42794);
xor U48525 (N_48525,N_41144,N_40869);
xor U48526 (N_48526,N_42594,N_42149);
or U48527 (N_48527,N_43160,N_40040);
xor U48528 (N_48528,N_43664,N_43506);
nand U48529 (N_48529,N_43437,N_42552);
xnor U48530 (N_48530,N_40848,N_40813);
nand U48531 (N_48531,N_41323,N_43867);
xor U48532 (N_48532,N_42225,N_41129);
xor U48533 (N_48533,N_41141,N_40603);
and U48534 (N_48534,N_40976,N_44752);
nor U48535 (N_48535,N_42468,N_42927);
nand U48536 (N_48536,N_42447,N_42891);
and U48537 (N_48537,N_40969,N_43907);
and U48538 (N_48538,N_40213,N_41204);
nor U48539 (N_48539,N_44863,N_44379);
nand U48540 (N_48540,N_40922,N_43491);
or U48541 (N_48541,N_44618,N_42410);
xnor U48542 (N_48542,N_44169,N_41067);
and U48543 (N_48543,N_40005,N_42808);
or U48544 (N_48544,N_43589,N_42116);
xnor U48545 (N_48545,N_41754,N_44597);
or U48546 (N_48546,N_42842,N_43304);
and U48547 (N_48547,N_41840,N_43624);
or U48548 (N_48548,N_44539,N_44498);
xor U48549 (N_48549,N_44285,N_43552);
xnor U48550 (N_48550,N_41678,N_41730);
xnor U48551 (N_48551,N_44946,N_42715);
xor U48552 (N_48552,N_43161,N_43619);
xnor U48553 (N_48553,N_41017,N_44539);
or U48554 (N_48554,N_40024,N_40660);
and U48555 (N_48555,N_40480,N_44147);
and U48556 (N_48556,N_44389,N_40135);
and U48557 (N_48557,N_41414,N_42685);
or U48558 (N_48558,N_41395,N_42948);
nor U48559 (N_48559,N_41245,N_40917);
nor U48560 (N_48560,N_41155,N_44549);
nand U48561 (N_48561,N_40522,N_43557);
nor U48562 (N_48562,N_44902,N_41267);
or U48563 (N_48563,N_40024,N_42063);
nor U48564 (N_48564,N_41504,N_40321);
xnor U48565 (N_48565,N_40166,N_43887);
nor U48566 (N_48566,N_40202,N_44445);
nor U48567 (N_48567,N_40018,N_41726);
xnor U48568 (N_48568,N_43978,N_40881);
and U48569 (N_48569,N_42711,N_43029);
nand U48570 (N_48570,N_41235,N_41533);
and U48571 (N_48571,N_44371,N_40073);
nand U48572 (N_48572,N_41422,N_40230);
and U48573 (N_48573,N_41401,N_44800);
nor U48574 (N_48574,N_44830,N_44923);
xor U48575 (N_48575,N_40009,N_42333);
xnor U48576 (N_48576,N_42761,N_41529);
nor U48577 (N_48577,N_40341,N_42015);
xor U48578 (N_48578,N_44119,N_40501);
nor U48579 (N_48579,N_42013,N_42954);
nor U48580 (N_48580,N_44436,N_42629);
and U48581 (N_48581,N_41471,N_41386);
nor U48582 (N_48582,N_42076,N_42095);
or U48583 (N_48583,N_41828,N_41145);
or U48584 (N_48584,N_41859,N_43546);
and U48585 (N_48585,N_40940,N_42275);
and U48586 (N_48586,N_43342,N_40443);
nor U48587 (N_48587,N_42835,N_41924);
xor U48588 (N_48588,N_43757,N_43216);
xnor U48589 (N_48589,N_41385,N_40720);
nor U48590 (N_48590,N_44129,N_41839);
nor U48591 (N_48591,N_43779,N_41009);
or U48592 (N_48592,N_44512,N_44331);
or U48593 (N_48593,N_42660,N_44586);
nor U48594 (N_48594,N_41655,N_40711);
xor U48595 (N_48595,N_42916,N_43276);
or U48596 (N_48596,N_41938,N_41752);
or U48597 (N_48597,N_40654,N_40857);
nor U48598 (N_48598,N_44781,N_41320);
or U48599 (N_48599,N_43687,N_43817);
xor U48600 (N_48600,N_40991,N_44547);
nor U48601 (N_48601,N_44393,N_42595);
nand U48602 (N_48602,N_44532,N_41200);
nor U48603 (N_48603,N_40908,N_43557);
and U48604 (N_48604,N_44564,N_42329);
and U48605 (N_48605,N_40164,N_42659);
or U48606 (N_48606,N_44921,N_43777);
nor U48607 (N_48607,N_40023,N_44489);
and U48608 (N_48608,N_40865,N_43114);
or U48609 (N_48609,N_40783,N_42272);
and U48610 (N_48610,N_40754,N_42166);
nor U48611 (N_48611,N_41694,N_44070);
or U48612 (N_48612,N_40853,N_43565);
and U48613 (N_48613,N_41602,N_41091);
xor U48614 (N_48614,N_41987,N_44830);
nand U48615 (N_48615,N_44476,N_43924);
nor U48616 (N_48616,N_41448,N_41010);
nand U48617 (N_48617,N_41009,N_41798);
or U48618 (N_48618,N_42001,N_40076);
nand U48619 (N_48619,N_44640,N_40040);
xor U48620 (N_48620,N_44434,N_42785);
nor U48621 (N_48621,N_44399,N_44016);
nand U48622 (N_48622,N_44875,N_41692);
xor U48623 (N_48623,N_40676,N_43494);
xnor U48624 (N_48624,N_44191,N_41094);
or U48625 (N_48625,N_44864,N_43951);
xor U48626 (N_48626,N_43305,N_41117);
nand U48627 (N_48627,N_40133,N_40176);
xnor U48628 (N_48628,N_42409,N_44072);
and U48629 (N_48629,N_41616,N_40563);
or U48630 (N_48630,N_40845,N_41792);
and U48631 (N_48631,N_41826,N_44841);
xnor U48632 (N_48632,N_40397,N_42241);
or U48633 (N_48633,N_43312,N_43698);
nor U48634 (N_48634,N_44629,N_43601);
and U48635 (N_48635,N_42351,N_41575);
xor U48636 (N_48636,N_44174,N_44626);
xnor U48637 (N_48637,N_42790,N_42353);
nand U48638 (N_48638,N_40176,N_44643);
nor U48639 (N_48639,N_44654,N_40917);
nor U48640 (N_48640,N_43220,N_41329);
or U48641 (N_48641,N_41502,N_44451);
xnor U48642 (N_48642,N_44026,N_42090);
nand U48643 (N_48643,N_43901,N_44854);
nor U48644 (N_48644,N_42321,N_41223);
or U48645 (N_48645,N_40174,N_44280);
nor U48646 (N_48646,N_40530,N_43485);
and U48647 (N_48647,N_40512,N_42343);
or U48648 (N_48648,N_44636,N_42681);
nor U48649 (N_48649,N_44478,N_41202);
and U48650 (N_48650,N_41727,N_43500);
nand U48651 (N_48651,N_43076,N_41572);
nor U48652 (N_48652,N_44493,N_42432);
and U48653 (N_48653,N_41797,N_40049);
nor U48654 (N_48654,N_42142,N_42126);
or U48655 (N_48655,N_43738,N_44301);
nor U48656 (N_48656,N_44352,N_43793);
or U48657 (N_48657,N_41112,N_42089);
nor U48658 (N_48658,N_40596,N_41340);
and U48659 (N_48659,N_43541,N_41093);
or U48660 (N_48660,N_44049,N_42359);
nand U48661 (N_48661,N_41291,N_44407);
nor U48662 (N_48662,N_41960,N_43345);
or U48663 (N_48663,N_40997,N_43190);
nor U48664 (N_48664,N_41345,N_43735);
nor U48665 (N_48665,N_43286,N_42887);
xor U48666 (N_48666,N_43092,N_41020);
nand U48667 (N_48667,N_40303,N_40801);
nor U48668 (N_48668,N_40345,N_44962);
xnor U48669 (N_48669,N_41018,N_43552);
nand U48670 (N_48670,N_44935,N_40679);
xnor U48671 (N_48671,N_43916,N_44353);
xnor U48672 (N_48672,N_43815,N_41044);
xnor U48673 (N_48673,N_41593,N_43748);
nor U48674 (N_48674,N_41316,N_41141);
xor U48675 (N_48675,N_43307,N_42550);
nor U48676 (N_48676,N_40132,N_43287);
xnor U48677 (N_48677,N_40164,N_41482);
or U48678 (N_48678,N_41574,N_42799);
nor U48679 (N_48679,N_41006,N_44384);
or U48680 (N_48680,N_42558,N_40452);
nand U48681 (N_48681,N_43921,N_44351);
xnor U48682 (N_48682,N_44073,N_40707);
and U48683 (N_48683,N_43312,N_43552);
and U48684 (N_48684,N_43590,N_43271);
xor U48685 (N_48685,N_40642,N_40357);
xnor U48686 (N_48686,N_41583,N_40915);
or U48687 (N_48687,N_42340,N_43832);
nand U48688 (N_48688,N_44886,N_40274);
and U48689 (N_48689,N_41225,N_41428);
and U48690 (N_48690,N_42017,N_41686);
and U48691 (N_48691,N_43543,N_40308);
nor U48692 (N_48692,N_44085,N_44852);
and U48693 (N_48693,N_43589,N_43690);
nor U48694 (N_48694,N_40498,N_40453);
nor U48695 (N_48695,N_40422,N_43153);
and U48696 (N_48696,N_43288,N_42755);
nand U48697 (N_48697,N_40274,N_41005);
nor U48698 (N_48698,N_44120,N_43794);
or U48699 (N_48699,N_43056,N_44039);
xor U48700 (N_48700,N_40990,N_41349);
and U48701 (N_48701,N_44078,N_42602);
nand U48702 (N_48702,N_43427,N_40045);
nor U48703 (N_48703,N_41012,N_44942);
and U48704 (N_48704,N_44686,N_42290);
nand U48705 (N_48705,N_43451,N_40236);
and U48706 (N_48706,N_43844,N_41336);
and U48707 (N_48707,N_43361,N_40935);
xor U48708 (N_48708,N_42096,N_40885);
or U48709 (N_48709,N_40900,N_42934);
nor U48710 (N_48710,N_41921,N_40877);
xnor U48711 (N_48711,N_40061,N_41304);
and U48712 (N_48712,N_41461,N_44099);
and U48713 (N_48713,N_43225,N_40537);
or U48714 (N_48714,N_41227,N_40018);
xnor U48715 (N_48715,N_44798,N_41670);
nor U48716 (N_48716,N_40917,N_43727);
nor U48717 (N_48717,N_42909,N_42779);
and U48718 (N_48718,N_43925,N_41484);
or U48719 (N_48719,N_40945,N_40644);
and U48720 (N_48720,N_40594,N_40716);
or U48721 (N_48721,N_43062,N_40758);
or U48722 (N_48722,N_41091,N_44311);
and U48723 (N_48723,N_42842,N_44113);
nor U48724 (N_48724,N_44695,N_44511);
or U48725 (N_48725,N_40439,N_44879);
nand U48726 (N_48726,N_42964,N_41294);
or U48727 (N_48727,N_42851,N_42202);
or U48728 (N_48728,N_42823,N_40261);
and U48729 (N_48729,N_43681,N_44280);
and U48730 (N_48730,N_42168,N_40657);
xnor U48731 (N_48731,N_44213,N_42597);
nand U48732 (N_48732,N_40157,N_42250);
nor U48733 (N_48733,N_43051,N_40332);
nor U48734 (N_48734,N_43873,N_43912);
or U48735 (N_48735,N_42356,N_44335);
and U48736 (N_48736,N_44270,N_43504);
or U48737 (N_48737,N_43791,N_43720);
nor U48738 (N_48738,N_41090,N_42142);
nor U48739 (N_48739,N_40212,N_44658);
and U48740 (N_48740,N_44307,N_44019);
nand U48741 (N_48741,N_42443,N_40815);
or U48742 (N_48742,N_43882,N_44592);
or U48743 (N_48743,N_42374,N_43065);
nand U48744 (N_48744,N_42305,N_40140);
nor U48745 (N_48745,N_44526,N_40554);
or U48746 (N_48746,N_44915,N_41143);
xnor U48747 (N_48747,N_42119,N_42354);
nand U48748 (N_48748,N_41858,N_43001);
nand U48749 (N_48749,N_44228,N_42059);
and U48750 (N_48750,N_43781,N_42492);
xor U48751 (N_48751,N_40085,N_41873);
nand U48752 (N_48752,N_41716,N_44192);
nor U48753 (N_48753,N_43030,N_42963);
nand U48754 (N_48754,N_40987,N_40392);
nor U48755 (N_48755,N_44235,N_40944);
xnor U48756 (N_48756,N_44210,N_40141);
and U48757 (N_48757,N_40748,N_44083);
or U48758 (N_48758,N_43728,N_41762);
nor U48759 (N_48759,N_41828,N_41972);
and U48760 (N_48760,N_40260,N_42615);
and U48761 (N_48761,N_41666,N_41162);
nor U48762 (N_48762,N_42765,N_43066);
or U48763 (N_48763,N_42321,N_40742);
nand U48764 (N_48764,N_40640,N_44661);
nand U48765 (N_48765,N_41633,N_40211);
xnor U48766 (N_48766,N_43460,N_42737);
nor U48767 (N_48767,N_43242,N_44896);
and U48768 (N_48768,N_42499,N_42279);
nand U48769 (N_48769,N_41462,N_40790);
and U48770 (N_48770,N_41101,N_42663);
nand U48771 (N_48771,N_40736,N_44375);
and U48772 (N_48772,N_40945,N_41730);
xor U48773 (N_48773,N_43109,N_43323);
nor U48774 (N_48774,N_43670,N_40749);
nand U48775 (N_48775,N_42569,N_41294);
or U48776 (N_48776,N_41384,N_44495);
or U48777 (N_48777,N_40316,N_43750);
or U48778 (N_48778,N_41911,N_42361);
nand U48779 (N_48779,N_40759,N_44440);
xnor U48780 (N_48780,N_41441,N_43329);
nor U48781 (N_48781,N_41225,N_44264);
nor U48782 (N_48782,N_40350,N_43584);
or U48783 (N_48783,N_43630,N_41586);
or U48784 (N_48784,N_43702,N_40368);
xor U48785 (N_48785,N_41830,N_44589);
and U48786 (N_48786,N_43102,N_43582);
nor U48787 (N_48787,N_44048,N_44282);
xnor U48788 (N_48788,N_42885,N_40558);
and U48789 (N_48789,N_40349,N_44243);
nand U48790 (N_48790,N_40537,N_43827);
or U48791 (N_48791,N_42943,N_44802);
nor U48792 (N_48792,N_41740,N_44128);
nand U48793 (N_48793,N_41020,N_42436);
xor U48794 (N_48794,N_43198,N_40846);
nor U48795 (N_48795,N_43194,N_43105);
xnor U48796 (N_48796,N_41544,N_42568);
xnor U48797 (N_48797,N_42539,N_43560);
nand U48798 (N_48798,N_41825,N_40508);
xor U48799 (N_48799,N_42406,N_42908);
or U48800 (N_48800,N_41071,N_40387);
or U48801 (N_48801,N_44171,N_42222);
and U48802 (N_48802,N_40606,N_44109);
nor U48803 (N_48803,N_42912,N_42820);
nand U48804 (N_48804,N_41676,N_44441);
or U48805 (N_48805,N_42824,N_40523);
xor U48806 (N_48806,N_43890,N_43664);
nor U48807 (N_48807,N_42065,N_41040);
nor U48808 (N_48808,N_41624,N_44207);
xnor U48809 (N_48809,N_42118,N_43851);
nand U48810 (N_48810,N_43929,N_40177);
nor U48811 (N_48811,N_43908,N_42474);
nor U48812 (N_48812,N_42950,N_40708);
nor U48813 (N_48813,N_41752,N_41152);
nand U48814 (N_48814,N_42352,N_44038);
or U48815 (N_48815,N_41899,N_44947);
or U48816 (N_48816,N_42808,N_40229);
or U48817 (N_48817,N_42835,N_41962);
nand U48818 (N_48818,N_40196,N_40004);
xnor U48819 (N_48819,N_44788,N_43085);
nor U48820 (N_48820,N_44832,N_41486);
xnor U48821 (N_48821,N_41691,N_44282);
nand U48822 (N_48822,N_43985,N_44572);
or U48823 (N_48823,N_40325,N_40144);
and U48824 (N_48824,N_44591,N_42719);
nand U48825 (N_48825,N_40912,N_42331);
xnor U48826 (N_48826,N_40841,N_41951);
nor U48827 (N_48827,N_41541,N_44602);
nor U48828 (N_48828,N_43527,N_44358);
nand U48829 (N_48829,N_43632,N_44163);
xnor U48830 (N_48830,N_40960,N_43041);
nor U48831 (N_48831,N_44301,N_40835);
nor U48832 (N_48832,N_44087,N_41564);
nor U48833 (N_48833,N_43189,N_43562);
or U48834 (N_48834,N_44123,N_44750);
nand U48835 (N_48835,N_42251,N_43977);
nor U48836 (N_48836,N_44031,N_40666);
nor U48837 (N_48837,N_43232,N_41229);
nand U48838 (N_48838,N_41348,N_42798);
or U48839 (N_48839,N_43198,N_44563);
xnor U48840 (N_48840,N_40544,N_42940);
nand U48841 (N_48841,N_42302,N_41117);
nor U48842 (N_48842,N_42782,N_44609);
xnor U48843 (N_48843,N_42039,N_44633);
xnor U48844 (N_48844,N_42548,N_44416);
nor U48845 (N_48845,N_43166,N_43834);
xor U48846 (N_48846,N_41294,N_41939);
and U48847 (N_48847,N_40435,N_41471);
nand U48848 (N_48848,N_43199,N_40812);
and U48849 (N_48849,N_43631,N_43253);
xor U48850 (N_48850,N_40875,N_42968);
nand U48851 (N_48851,N_40058,N_41714);
or U48852 (N_48852,N_42409,N_44992);
nand U48853 (N_48853,N_44628,N_44154);
and U48854 (N_48854,N_42874,N_42429);
nor U48855 (N_48855,N_44217,N_40579);
or U48856 (N_48856,N_42884,N_43736);
nor U48857 (N_48857,N_41668,N_41835);
nor U48858 (N_48858,N_43812,N_43989);
and U48859 (N_48859,N_41658,N_44023);
nor U48860 (N_48860,N_43528,N_44315);
and U48861 (N_48861,N_41408,N_42502);
or U48862 (N_48862,N_42439,N_40289);
xor U48863 (N_48863,N_41270,N_44834);
or U48864 (N_48864,N_41413,N_42180);
or U48865 (N_48865,N_41053,N_43268);
xnor U48866 (N_48866,N_43280,N_44452);
xor U48867 (N_48867,N_41467,N_44204);
nor U48868 (N_48868,N_41221,N_40612);
xnor U48869 (N_48869,N_43611,N_42983);
or U48870 (N_48870,N_41309,N_43093);
or U48871 (N_48871,N_41151,N_41572);
or U48872 (N_48872,N_41414,N_40315);
xor U48873 (N_48873,N_42215,N_42005);
xnor U48874 (N_48874,N_42048,N_40249);
nand U48875 (N_48875,N_44299,N_40127);
or U48876 (N_48876,N_42136,N_42871);
xor U48877 (N_48877,N_40112,N_44463);
or U48878 (N_48878,N_41880,N_41396);
xnor U48879 (N_48879,N_41298,N_43617);
or U48880 (N_48880,N_43860,N_41779);
xnor U48881 (N_48881,N_44834,N_43086);
and U48882 (N_48882,N_43980,N_42004);
xnor U48883 (N_48883,N_40177,N_40145);
and U48884 (N_48884,N_44910,N_40978);
nor U48885 (N_48885,N_43773,N_40046);
xnor U48886 (N_48886,N_43415,N_43627);
xnor U48887 (N_48887,N_44788,N_40498);
xor U48888 (N_48888,N_42494,N_44749);
and U48889 (N_48889,N_40429,N_43964);
and U48890 (N_48890,N_44233,N_43632);
nor U48891 (N_48891,N_44795,N_43460);
nand U48892 (N_48892,N_40678,N_43466);
and U48893 (N_48893,N_40336,N_41356);
nand U48894 (N_48894,N_44898,N_43670);
nand U48895 (N_48895,N_44981,N_44765);
nor U48896 (N_48896,N_44644,N_42667);
and U48897 (N_48897,N_40660,N_41345);
xnor U48898 (N_48898,N_43030,N_41919);
nand U48899 (N_48899,N_40746,N_41282);
xor U48900 (N_48900,N_41684,N_43072);
nand U48901 (N_48901,N_42436,N_44553);
or U48902 (N_48902,N_44499,N_43005);
or U48903 (N_48903,N_44051,N_41585);
xor U48904 (N_48904,N_40333,N_41816);
or U48905 (N_48905,N_44843,N_40295);
and U48906 (N_48906,N_40007,N_43903);
or U48907 (N_48907,N_40967,N_44682);
xnor U48908 (N_48908,N_42043,N_42169);
or U48909 (N_48909,N_43044,N_40591);
and U48910 (N_48910,N_42852,N_43456);
nand U48911 (N_48911,N_41213,N_43069);
xor U48912 (N_48912,N_43959,N_42497);
nor U48913 (N_48913,N_43480,N_44000);
nand U48914 (N_48914,N_44230,N_44345);
or U48915 (N_48915,N_40307,N_44539);
nor U48916 (N_48916,N_40560,N_40857);
and U48917 (N_48917,N_42094,N_44362);
and U48918 (N_48918,N_41515,N_40153);
nand U48919 (N_48919,N_44858,N_42834);
xnor U48920 (N_48920,N_44640,N_41370);
and U48921 (N_48921,N_43044,N_43394);
nor U48922 (N_48922,N_42401,N_41844);
and U48923 (N_48923,N_41302,N_44735);
nor U48924 (N_48924,N_42640,N_41178);
or U48925 (N_48925,N_43514,N_42542);
xnor U48926 (N_48926,N_43752,N_43775);
nor U48927 (N_48927,N_43840,N_41860);
nand U48928 (N_48928,N_44974,N_41478);
nor U48929 (N_48929,N_43613,N_43082);
xor U48930 (N_48930,N_40168,N_43579);
nand U48931 (N_48931,N_44125,N_41911);
and U48932 (N_48932,N_42243,N_40771);
xnor U48933 (N_48933,N_42864,N_43185);
and U48934 (N_48934,N_43068,N_40322);
and U48935 (N_48935,N_41949,N_40161);
nand U48936 (N_48936,N_42183,N_41339);
and U48937 (N_48937,N_40938,N_42713);
or U48938 (N_48938,N_44488,N_43668);
nand U48939 (N_48939,N_44162,N_40741);
and U48940 (N_48940,N_43523,N_44140);
and U48941 (N_48941,N_42832,N_40929);
nor U48942 (N_48942,N_41984,N_42593);
nand U48943 (N_48943,N_40980,N_44407);
or U48944 (N_48944,N_44273,N_40121);
xnor U48945 (N_48945,N_44578,N_43792);
or U48946 (N_48946,N_43982,N_42323);
or U48947 (N_48947,N_42644,N_40825);
xnor U48948 (N_48948,N_41165,N_40769);
nor U48949 (N_48949,N_41757,N_42512);
nor U48950 (N_48950,N_43137,N_43953);
nor U48951 (N_48951,N_43062,N_41307);
nor U48952 (N_48952,N_40516,N_40725);
or U48953 (N_48953,N_43698,N_42841);
xnor U48954 (N_48954,N_41703,N_41021);
or U48955 (N_48955,N_41818,N_42476);
or U48956 (N_48956,N_40405,N_44590);
or U48957 (N_48957,N_40025,N_42725);
or U48958 (N_48958,N_41743,N_43121);
nand U48959 (N_48959,N_41374,N_44108);
xnor U48960 (N_48960,N_44449,N_42708);
nand U48961 (N_48961,N_44298,N_43038);
nor U48962 (N_48962,N_40256,N_41889);
nand U48963 (N_48963,N_42313,N_43518);
and U48964 (N_48964,N_42207,N_44310);
and U48965 (N_48965,N_41747,N_43888);
nor U48966 (N_48966,N_42659,N_44779);
nor U48967 (N_48967,N_40622,N_42419);
and U48968 (N_48968,N_43740,N_41951);
xor U48969 (N_48969,N_43449,N_43199);
xor U48970 (N_48970,N_43980,N_42864);
and U48971 (N_48971,N_43415,N_44486);
and U48972 (N_48972,N_44389,N_42314);
nand U48973 (N_48973,N_40753,N_44373);
xor U48974 (N_48974,N_40229,N_42715);
nand U48975 (N_48975,N_40391,N_44685);
nor U48976 (N_48976,N_42952,N_40559);
xnor U48977 (N_48977,N_40078,N_43816);
and U48978 (N_48978,N_44707,N_43319);
nor U48979 (N_48979,N_44360,N_40247);
nor U48980 (N_48980,N_41916,N_41220);
and U48981 (N_48981,N_44627,N_40473);
and U48982 (N_48982,N_43332,N_44630);
nand U48983 (N_48983,N_42757,N_44336);
nand U48984 (N_48984,N_44628,N_44732);
or U48985 (N_48985,N_41767,N_43418);
or U48986 (N_48986,N_42983,N_40330);
and U48987 (N_48987,N_44537,N_41032);
and U48988 (N_48988,N_42898,N_42092);
nand U48989 (N_48989,N_41873,N_40591);
or U48990 (N_48990,N_43427,N_41335);
nor U48991 (N_48991,N_43637,N_41815);
or U48992 (N_48992,N_40181,N_40486);
nor U48993 (N_48993,N_40396,N_43409);
or U48994 (N_48994,N_40239,N_44223);
and U48995 (N_48995,N_40897,N_40197);
nor U48996 (N_48996,N_44631,N_43057);
nand U48997 (N_48997,N_42805,N_41618);
nor U48998 (N_48998,N_41018,N_43794);
and U48999 (N_48999,N_41155,N_42962);
and U49000 (N_49000,N_41209,N_40636);
or U49001 (N_49001,N_41078,N_41368);
xnor U49002 (N_49002,N_40627,N_44662);
and U49003 (N_49003,N_44921,N_44437);
nor U49004 (N_49004,N_41106,N_40632);
nor U49005 (N_49005,N_41238,N_44295);
xnor U49006 (N_49006,N_42014,N_44599);
and U49007 (N_49007,N_40451,N_43222);
nor U49008 (N_49008,N_43157,N_42398);
nor U49009 (N_49009,N_41854,N_43676);
nand U49010 (N_49010,N_40959,N_44490);
nand U49011 (N_49011,N_41722,N_41340);
xor U49012 (N_49012,N_44165,N_42741);
nor U49013 (N_49013,N_40963,N_40799);
or U49014 (N_49014,N_42692,N_40776);
nand U49015 (N_49015,N_40830,N_44137);
nand U49016 (N_49016,N_43292,N_42056);
xor U49017 (N_49017,N_40663,N_42215);
and U49018 (N_49018,N_42230,N_40984);
or U49019 (N_49019,N_43696,N_41974);
xor U49020 (N_49020,N_42768,N_40547);
nand U49021 (N_49021,N_41265,N_42289);
nand U49022 (N_49022,N_43630,N_43098);
or U49023 (N_49023,N_41937,N_43774);
nor U49024 (N_49024,N_43559,N_41731);
nand U49025 (N_49025,N_40518,N_44811);
nor U49026 (N_49026,N_41712,N_44067);
xor U49027 (N_49027,N_40264,N_42631);
and U49028 (N_49028,N_41060,N_41588);
nand U49029 (N_49029,N_43778,N_40148);
nand U49030 (N_49030,N_44191,N_40255);
or U49031 (N_49031,N_44025,N_41347);
nand U49032 (N_49032,N_44405,N_44813);
and U49033 (N_49033,N_43251,N_40469);
nor U49034 (N_49034,N_40798,N_42489);
nor U49035 (N_49035,N_41519,N_41040);
nand U49036 (N_49036,N_40826,N_42279);
and U49037 (N_49037,N_40828,N_44319);
or U49038 (N_49038,N_41221,N_40943);
xnor U49039 (N_49039,N_40573,N_40562);
nor U49040 (N_49040,N_42560,N_43718);
xor U49041 (N_49041,N_42718,N_44070);
xor U49042 (N_49042,N_40593,N_43950);
and U49043 (N_49043,N_44831,N_44733);
nand U49044 (N_49044,N_42597,N_41131);
nor U49045 (N_49045,N_42302,N_43703);
xnor U49046 (N_49046,N_41091,N_42774);
nand U49047 (N_49047,N_42163,N_40224);
and U49048 (N_49048,N_40100,N_41449);
and U49049 (N_49049,N_44497,N_43930);
xnor U49050 (N_49050,N_44121,N_43386);
and U49051 (N_49051,N_41649,N_43729);
and U49052 (N_49052,N_44695,N_41284);
xor U49053 (N_49053,N_41806,N_44359);
and U49054 (N_49054,N_42790,N_42123);
nand U49055 (N_49055,N_44909,N_41695);
and U49056 (N_49056,N_43597,N_43137);
nand U49057 (N_49057,N_44423,N_43323);
nand U49058 (N_49058,N_43828,N_41171);
and U49059 (N_49059,N_41214,N_41578);
nor U49060 (N_49060,N_41018,N_41466);
and U49061 (N_49061,N_43471,N_43363);
and U49062 (N_49062,N_40111,N_41914);
xor U49063 (N_49063,N_42323,N_41571);
nand U49064 (N_49064,N_43328,N_40854);
nor U49065 (N_49065,N_42133,N_40506);
xor U49066 (N_49066,N_41624,N_40887);
and U49067 (N_49067,N_42835,N_44763);
nand U49068 (N_49068,N_41705,N_43776);
nor U49069 (N_49069,N_41763,N_40877);
or U49070 (N_49070,N_41098,N_40595);
nor U49071 (N_49071,N_41524,N_42556);
and U49072 (N_49072,N_40822,N_42783);
xor U49073 (N_49073,N_41889,N_44463);
xnor U49074 (N_49074,N_41780,N_43390);
or U49075 (N_49075,N_41522,N_40665);
xor U49076 (N_49076,N_41045,N_41623);
and U49077 (N_49077,N_44983,N_41957);
xnor U49078 (N_49078,N_44670,N_41343);
xnor U49079 (N_49079,N_40447,N_42763);
or U49080 (N_49080,N_42305,N_40332);
nor U49081 (N_49081,N_44804,N_41898);
nand U49082 (N_49082,N_43071,N_40927);
nand U49083 (N_49083,N_40029,N_43913);
nor U49084 (N_49084,N_43867,N_43068);
nor U49085 (N_49085,N_42390,N_40562);
xor U49086 (N_49086,N_42936,N_42085);
or U49087 (N_49087,N_41059,N_42554);
or U49088 (N_49088,N_44676,N_42899);
nor U49089 (N_49089,N_40841,N_42286);
and U49090 (N_49090,N_42020,N_42680);
nand U49091 (N_49091,N_43761,N_44885);
and U49092 (N_49092,N_41090,N_42360);
nand U49093 (N_49093,N_44239,N_40005);
and U49094 (N_49094,N_44574,N_42259);
nand U49095 (N_49095,N_40904,N_41458);
nand U49096 (N_49096,N_42658,N_40027);
xnor U49097 (N_49097,N_44442,N_41092);
or U49098 (N_49098,N_40588,N_43316);
nand U49099 (N_49099,N_44163,N_42779);
xnor U49100 (N_49100,N_42867,N_43366);
or U49101 (N_49101,N_41909,N_40691);
nand U49102 (N_49102,N_42285,N_44267);
nor U49103 (N_49103,N_40641,N_41776);
and U49104 (N_49104,N_40308,N_42098);
xnor U49105 (N_49105,N_41739,N_43265);
and U49106 (N_49106,N_42770,N_42303);
nand U49107 (N_49107,N_43778,N_41980);
and U49108 (N_49108,N_42483,N_42660);
or U49109 (N_49109,N_42507,N_40711);
and U49110 (N_49110,N_41824,N_42003);
nor U49111 (N_49111,N_44916,N_40220);
xnor U49112 (N_49112,N_43025,N_41680);
nor U49113 (N_49113,N_41218,N_44885);
nand U49114 (N_49114,N_40796,N_43786);
or U49115 (N_49115,N_44668,N_43080);
or U49116 (N_49116,N_40167,N_42316);
xnor U49117 (N_49117,N_40354,N_44012);
nor U49118 (N_49118,N_44684,N_42342);
nand U49119 (N_49119,N_43657,N_40941);
or U49120 (N_49120,N_43272,N_43386);
xor U49121 (N_49121,N_44198,N_44490);
and U49122 (N_49122,N_44502,N_41911);
or U49123 (N_49123,N_43517,N_41456);
nor U49124 (N_49124,N_43911,N_40517);
nor U49125 (N_49125,N_40245,N_41153);
nand U49126 (N_49126,N_41969,N_40814);
nand U49127 (N_49127,N_40045,N_41209);
xnor U49128 (N_49128,N_40160,N_42776);
nand U49129 (N_49129,N_40673,N_40776);
nand U49130 (N_49130,N_42764,N_44999);
and U49131 (N_49131,N_42689,N_44531);
nor U49132 (N_49132,N_41222,N_40120);
xnor U49133 (N_49133,N_41999,N_42079);
nand U49134 (N_49134,N_41114,N_42410);
nor U49135 (N_49135,N_44115,N_41124);
xor U49136 (N_49136,N_44741,N_44099);
and U49137 (N_49137,N_41540,N_42629);
xnor U49138 (N_49138,N_42586,N_43315);
xnor U49139 (N_49139,N_42331,N_41948);
and U49140 (N_49140,N_41264,N_40364);
or U49141 (N_49141,N_42395,N_43580);
and U49142 (N_49142,N_41011,N_40326);
or U49143 (N_49143,N_42693,N_41065);
xnor U49144 (N_49144,N_41276,N_41035);
or U49145 (N_49145,N_44328,N_43310);
xnor U49146 (N_49146,N_41766,N_43033);
nand U49147 (N_49147,N_42109,N_43710);
or U49148 (N_49148,N_43999,N_43690);
nand U49149 (N_49149,N_44952,N_42036);
nand U49150 (N_49150,N_42809,N_44412);
nor U49151 (N_49151,N_40498,N_44979);
and U49152 (N_49152,N_43122,N_44238);
nor U49153 (N_49153,N_43391,N_41599);
and U49154 (N_49154,N_41714,N_43337);
xnor U49155 (N_49155,N_40525,N_41538);
or U49156 (N_49156,N_43085,N_43748);
nand U49157 (N_49157,N_42212,N_44762);
or U49158 (N_49158,N_43817,N_40199);
nor U49159 (N_49159,N_44005,N_41929);
nand U49160 (N_49160,N_41150,N_41970);
nand U49161 (N_49161,N_41847,N_40059);
nor U49162 (N_49162,N_42810,N_42409);
or U49163 (N_49163,N_42272,N_41405);
nand U49164 (N_49164,N_42301,N_43920);
and U49165 (N_49165,N_44224,N_42162);
nor U49166 (N_49166,N_40580,N_42993);
nor U49167 (N_49167,N_40712,N_43130);
and U49168 (N_49168,N_43506,N_41917);
nand U49169 (N_49169,N_43846,N_44887);
nor U49170 (N_49170,N_40703,N_43728);
and U49171 (N_49171,N_41920,N_43312);
xnor U49172 (N_49172,N_44378,N_42103);
xor U49173 (N_49173,N_43395,N_41154);
nand U49174 (N_49174,N_44858,N_44706);
nor U49175 (N_49175,N_44561,N_40258);
nand U49176 (N_49176,N_41537,N_41513);
nand U49177 (N_49177,N_44232,N_40906);
and U49178 (N_49178,N_41375,N_40155);
nor U49179 (N_49179,N_42405,N_44941);
or U49180 (N_49180,N_44695,N_44697);
nand U49181 (N_49181,N_43931,N_42889);
and U49182 (N_49182,N_44279,N_43458);
nor U49183 (N_49183,N_40351,N_42566);
and U49184 (N_49184,N_43934,N_44177);
xor U49185 (N_49185,N_43198,N_43519);
and U49186 (N_49186,N_40187,N_44876);
and U49187 (N_49187,N_42771,N_42314);
xor U49188 (N_49188,N_43630,N_40817);
and U49189 (N_49189,N_44204,N_44632);
or U49190 (N_49190,N_40291,N_40928);
nand U49191 (N_49191,N_42290,N_42413);
nand U49192 (N_49192,N_42082,N_42792);
and U49193 (N_49193,N_40558,N_40762);
and U49194 (N_49194,N_43087,N_41497);
or U49195 (N_49195,N_44449,N_43283);
or U49196 (N_49196,N_41001,N_44745);
or U49197 (N_49197,N_43843,N_40470);
and U49198 (N_49198,N_41542,N_44764);
xnor U49199 (N_49199,N_40417,N_40287);
nor U49200 (N_49200,N_44302,N_44214);
nor U49201 (N_49201,N_44230,N_40862);
or U49202 (N_49202,N_43959,N_43451);
and U49203 (N_49203,N_41149,N_41362);
nor U49204 (N_49204,N_43625,N_42834);
xnor U49205 (N_49205,N_42291,N_42145);
or U49206 (N_49206,N_40312,N_42068);
nand U49207 (N_49207,N_40434,N_43687);
and U49208 (N_49208,N_44825,N_41426);
or U49209 (N_49209,N_42935,N_43192);
xnor U49210 (N_49210,N_41226,N_44919);
nand U49211 (N_49211,N_42438,N_40290);
nor U49212 (N_49212,N_42061,N_43218);
xnor U49213 (N_49213,N_41179,N_44936);
nand U49214 (N_49214,N_43528,N_44130);
and U49215 (N_49215,N_42052,N_44430);
nand U49216 (N_49216,N_42910,N_44034);
or U49217 (N_49217,N_43692,N_43616);
or U49218 (N_49218,N_40447,N_41178);
nand U49219 (N_49219,N_42890,N_44990);
nand U49220 (N_49220,N_41056,N_42202);
xor U49221 (N_49221,N_41163,N_41202);
nor U49222 (N_49222,N_42431,N_42804);
nor U49223 (N_49223,N_41428,N_40379);
or U49224 (N_49224,N_41652,N_43320);
nor U49225 (N_49225,N_44193,N_42343);
or U49226 (N_49226,N_42212,N_43208);
or U49227 (N_49227,N_44834,N_44053);
and U49228 (N_49228,N_43545,N_41412);
and U49229 (N_49229,N_40613,N_44626);
xor U49230 (N_49230,N_42040,N_42462);
and U49231 (N_49231,N_43250,N_40405);
and U49232 (N_49232,N_42579,N_43607);
xnor U49233 (N_49233,N_44884,N_42117);
nand U49234 (N_49234,N_44316,N_42685);
and U49235 (N_49235,N_41363,N_43964);
or U49236 (N_49236,N_42175,N_43645);
xor U49237 (N_49237,N_43829,N_43732);
and U49238 (N_49238,N_43222,N_44697);
or U49239 (N_49239,N_43310,N_42816);
nand U49240 (N_49240,N_44415,N_40682);
xnor U49241 (N_49241,N_41203,N_44859);
xnor U49242 (N_49242,N_44293,N_44358);
nor U49243 (N_49243,N_42270,N_41225);
and U49244 (N_49244,N_41755,N_43578);
xor U49245 (N_49245,N_41095,N_42284);
nor U49246 (N_49246,N_44459,N_42819);
nand U49247 (N_49247,N_42776,N_40408);
and U49248 (N_49248,N_40768,N_42997);
or U49249 (N_49249,N_40830,N_40918);
and U49250 (N_49250,N_41629,N_44269);
nor U49251 (N_49251,N_42461,N_44871);
nor U49252 (N_49252,N_42415,N_40255);
and U49253 (N_49253,N_42143,N_43851);
nor U49254 (N_49254,N_44847,N_41947);
and U49255 (N_49255,N_42282,N_42426);
xnor U49256 (N_49256,N_41622,N_41354);
nand U49257 (N_49257,N_40251,N_44058);
xnor U49258 (N_49258,N_42344,N_41290);
nand U49259 (N_49259,N_40518,N_41805);
nand U49260 (N_49260,N_40895,N_44550);
xnor U49261 (N_49261,N_42279,N_43554);
and U49262 (N_49262,N_44196,N_40552);
nand U49263 (N_49263,N_43591,N_41448);
nor U49264 (N_49264,N_44588,N_43230);
nand U49265 (N_49265,N_42886,N_41539);
or U49266 (N_49266,N_40648,N_41092);
xnor U49267 (N_49267,N_42325,N_40869);
nor U49268 (N_49268,N_40702,N_41747);
nand U49269 (N_49269,N_41007,N_44765);
xor U49270 (N_49270,N_40618,N_43278);
xor U49271 (N_49271,N_43769,N_43717);
xor U49272 (N_49272,N_41517,N_41001);
nor U49273 (N_49273,N_44973,N_42122);
and U49274 (N_49274,N_43269,N_40146);
or U49275 (N_49275,N_40838,N_42161);
nor U49276 (N_49276,N_40420,N_40296);
and U49277 (N_49277,N_44038,N_41808);
xnor U49278 (N_49278,N_41514,N_43246);
nor U49279 (N_49279,N_43859,N_40991);
or U49280 (N_49280,N_42505,N_43521);
xor U49281 (N_49281,N_41887,N_40697);
and U49282 (N_49282,N_40096,N_44508);
and U49283 (N_49283,N_44689,N_41113);
xor U49284 (N_49284,N_40578,N_41223);
and U49285 (N_49285,N_42288,N_42020);
nand U49286 (N_49286,N_40988,N_40269);
or U49287 (N_49287,N_42548,N_44549);
nand U49288 (N_49288,N_44021,N_44295);
or U49289 (N_49289,N_41355,N_42109);
xnor U49290 (N_49290,N_41667,N_42818);
or U49291 (N_49291,N_43089,N_41659);
or U49292 (N_49292,N_42265,N_42452);
or U49293 (N_49293,N_42714,N_44626);
xnor U49294 (N_49294,N_41287,N_42498);
xor U49295 (N_49295,N_42912,N_41001);
or U49296 (N_49296,N_44563,N_42560);
nand U49297 (N_49297,N_41689,N_42104);
nand U49298 (N_49298,N_44024,N_44841);
xnor U49299 (N_49299,N_42500,N_42213);
or U49300 (N_49300,N_41644,N_43639);
nand U49301 (N_49301,N_40611,N_43701);
or U49302 (N_49302,N_41161,N_40093);
nor U49303 (N_49303,N_44845,N_44973);
or U49304 (N_49304,N_40293,N_42034);
and U49305 (N_49305,N_44538,N_40670);
xnor U49306 (N_49306,N_43206,N_44817);
nand U49307 (N_49307,N_42577,N_43131);
or U49308 (N_49308,N_44801,N_43914);
xnor U49309 (N_49309,N_43974,N_43621);
or U49310 (N_49310,N_40836,N_40729);
nor U49311 (N_49311,N_44566,N_40786);
and U49312 (N_49312,N_44805,N_40562);
xor U49313 (N_49313,N_43445,N_44286);
or U49314 (N_49314,N_42653,N_42703);
and U49315 (N_49315,N_42152,N_40876);
nand U49316 (N_49316,N_40818,N_41337);
xor U49317 (N_49317,N_44530,N_44654);
or U49318 (N_49318,N_43500,N_40718);
and U49319 (N_49319,N_44750,N_42482);
xor U49320 (N_49320,N_43080,N_44607);
xnor U49321 (N_49321,N_42559,N_43510);
nor U49322 (N_49322,N_41453,N_43646);
nand U49323 (N_49323,N_44266,N_42320);
or U49324 (N_49324,N_41453,N_40213);
nand U49325 (N_49325,N_42345,N_44787);
nor U49326 (N_49326,N_42423,N_40825);
or U49327 (N_49327,N_44401,N_41436);
nor U49328 (N_49328,N_44746,N_44494);
or U49329 (N_49329,N_43295,N_43731);
nand U49330 (N_49330,N_43062,N_44265);
nand U49331 (N_49331,N_42218,N_40669);
and U49332 (N_49332,N_44355,N_44247);
or U49333 (N_49333,N_44749,N_42352);
nand U49334 (N_49334,N_43863,N_40956);
xnor U49335 (N_49335,N_40963,N_41485);
and U49336 (N_49336,N_44811,N_42117);
nand U49337 (N_49337,N_44628,N_43330);
xor U49338 (N_49338,N_43654,N_42011);
and U49339 (N_49339,N_43657,N_42220);
nand U49340 (N_49340,N_40628,N_41704);
and U49341 (N_49341,N_44455,N_44220);
xor U49342 (N_49342,N_42803,N_40811);
or U49343 (N_49343,N_42970,N_43408);
nand U49344 (N_49344,N_43307,N_44794);
nor U49345 (N_49345,N_40913,N_40331);
xnor U49346 (N_49346,N_42645,N_41119);
and U49347 (N_49347,N_43282,N_43169);
and U49348 (N_49348,N_40784,N_40013);
nand U49349 (N_49349,N_44809,N_44323);
nor U49350 (N_49350,N_42072,N_42319);
nand U49351 (N_49351,N_43003,N_43797);
nand U49352 (N_49352,N_42123,N_40079);
nand U49353 (N_49353,N_40008,N_44458);
nor U49354 (N_49354,N_42523,N_43536);
and U49355 (N_49355,N_41688,N_43228);
xnor U49356 (N_49356,N_40837,N_43767);
or U49357 (N_49357,N_41333,N_40509);
and U49358 (N_49358,N_40954,N_41735);
and U49359 (N_49359,N_44823,N_44462);
nand U49360 (N_49360,N_40034,N_41009);
nor U49361 (N_49361,N_44792,N_40661);
nor U49362 (N_49362,N_44179,N_42680);
and U49363 (N_49363,N_41046,N_43065);
nand U49364 (N_49364,N_42014,N_40704);
nand U49365 (N_49365,N_43497,N_41432);
nand U49366 (N_49366,N_44555,N_42833);
nor U49367 (N_49367,N_43727,N_41849);
and U49368 (N_49368,N_42106,N_42621);
xor U49369 (N_49369,N_43644,N_40046);
xnor U49370 (N_49370,N_42427,N_41239);
nand U49371 (N_49371,N_42710,N_40619);
nor U49372 (N_49372,N_42259,N_40636);
xor U49373 (N_49373,N_43230,N_42836);
or U49374 (N_49374,N_43568,N_42487);
nor U49375 (N_49375,N_43433,N_41866);
or U49376 (N_49376,N_43281,N_42127);
nor U49377 (N_49377,N_42209,N_41034);
nand U49378 (N_49378,N_44961,N_44628);
and U49379 (N_49379,N_41985,N_41502);
nand U49380 (N_49380,N_43928,N_41425);
xnor U49381 (N_49381,N_41126,N_43827);
nand U49382 (N_49382,N_41609,N_42009);
nor U49383 (N_49383,N_41431,N_42445);
nand U49384 (N_49384,N_42942,N_40444);
or U49385 (N_49385,N_43453,N_42124);
nor U49386 (N_49386,N_42604,N_43130);
and U49387 (N_49387,N_43876,N_41104);
and U49388 (N_49388,N_44491,N_44429);
nor U49389 (N_49389,N_42993,N_40195);
and U49390 (N_49390,N_43110,N_43019);
xnor U49391 (N_49391,N_41079,N_43885);
xnor U49392 (N_49392,N_43625,N_41586);
and U49393 (N_49393,N_41464,N_40507);
nor U49394 (N_49394,N_40355,N_43909);
nand U49395 (N_49395,N_44857,N_43058);
or U49396 (N_49396,N_40171,N_41504);
nor U49397 (N_49397,N_41639,N_40259);
and U49398 (N_49398,N_41945,N_40245);
nand U49399 (N_49399,N_40478,N_40125);
nor U49400 (N_49400,N_40449,N_40822);
and U49401 (N_49401,N_43370,N_41116);
or U49402 (N_49402,N_40059,N_40842);
xor U49403 (N_49403,N_43442,N_41808);
nor U49404 (N_49404,N_41297,N_43293);
or U49405 (N_49405,N_43238,N_44125);
and U49406 (N_49406,N_42480,N_41001);
nor U49407 (N_49407,N_43464,N_41838);
and U49408 (N_49408,N_40957,N_44652);
xnor U49409 (N_49409,N_41528,N_42599);
or U49410 (N_49410,N_41037,N_40501);
nand U49411 (N_49411,N_43160,N_40747);
nor U49412 (N_49412,N_42191,N_40874);
nand U49413 (N_49413,N_40828,N_43493);
nand U49414 (N_49414,N_44869,N_43618);
and U49415 (N_49415,N_43022,N_42414);
and U49416 (N_49416,N_44493,N_43283);
or U49417 (N_49417,N_41697,N_41271);
and U49418 (N_49418,N_43964,N_41283);
nand U49419 (N_49419,N_42948,N_44729);
nor U49420 (N_49420,N_42753,N_44506);
nor U49421 (N_49421,N_42755,N_41442);
or U49422 (N_49422,N_41806,N_41662);
and U49423 (N_49423,N_40535,N_44159);
xnor U49424 (N_49424,N_44822,N_43720);
nand U49425 (N_49425,N_42441,N_41259);
xor U49426 (N_49426,N_41354,N_44886);
nor U49427 (N_49427,N_42558,N_42430);
or U49428 (N_49428,N_43168,N_40015);
nand U49429 (N_49429,N_43344,N_41391);
xor U49430 (N_49430,N_40984,N_43135);
or U49431 (N_49431,N_42446,N_41477);
xnor U49432 (N_49432,N_44942,N_41479);
or U49433 (N_49433,N_42604,N_42747);
xnor U49434 (N_49434,N_41865,N_44289);
nor U49435 (N_49435,N_44567,N_44496);
xnor U49436 (N_49436,N_44915,N_40081);
nor U49437 (N_49437,N_41782,N_44587);
xor U49438 (N_49438,N_41312,N_44207);
xor U49439 (N_49439,N_44783,N_42735);
nor U49440 (N_49440,N_41793,N_42736);
or U49441 (N_49441,N_43683,N_42409);
and U49442 (N_49442,N_44997,N_41667);
nand U49443 (N_49443,N_40355,N_42905);
nand U49444 (N_49444,N_44453,N_44596);
xor U49445 (N_49445,N_44936,N_42429);
or U49446 (N_49446,N_40636,N_41331);
nand U49447 (N_49447,N_44052,N_40940);
nand U49448 (N_49448,N_41254,N_43812);
or U49449 (N_49449,N_41249,N_42460);
xnor U49450 (N_49450,N_44788,N_40723);
nor U49451 (N_49451,N_42320,N_42116);
nand U49452 (N_49452,N_43594,N_44567);
nor U49453 (N_49453,N_42477,N_41270);
or U49454 (N_49454,N_42543,N_41039);
nor U49455 (N_49455,N_44966,N_43798);
nor U49456 (N_49456,N_43362,N_44092);
xor U49457 (N_49457,N_40590,N_40436);
and U49458 (N_49458,N_44134,N_40186);
and U49459 (N_49459,N_40529,N_41652);
and U49460 (N_49460,N_41055,N_42758);
nand U49461 (N_49461,N_43118,N_44508);
xnor U49462 (N_49462,N_42060,N_40019);
nand U49463 (N_49463,N_43769,N_43959);
or U49464 (N_49464,N_44181,N_43820);
nand U49465 (N_49465,N_40199,N_42807);
nand U49466 (N_49466,N_42037,N_44066);
nand U49467 (N_49467,N_43648,N_42380);
or U49468 (N_49468,N_43505,N_41829);
or U49469 (N_49469,N_43344,N_43400);
nor U49470 (N_49470,N_40645,N_44478);
nand U49471 (N_49471,N_43180,N_40345);
or U49472 (N_49472,N_43346,N_41329);
nor U49473 (N_49473,N_40950,N_40038);
or U49474 (N_49474,N_41855,N_42579);
xnor U49475 (N_49475,N_41150,N_40913);
nor U49476 (N_49476,N_43525,N_44435);
and U49477 (N_49477,N_42686,N_41374);
or U49478 (N_49478,N_41200,N_42487);
nand U49479 (N_49479,N_42640,N_44967);
or U49480 (N_49480,N_40212,N_41721);
nand U49481 (N_49481,N_41197,N_40126);
xor U49482 (N_49482,N_41567,N_42198);
xor U49483 (N_49483,N_42873,N_42372);
or U49484 (N_49484,N_42926,N_42527);
nor U49485 (N_49485,N_40406,N_41343);
nor U49486 (N_49486,N_42492,N_43042);
nand U49487 (N_49487,N_40897,N_40918);
or U49488 (N_49488,N_43300,N_44797);
nand U49489 (N_49489,N_44023,N_43177);
xnor U49490 (N_49490,N_44320,N_44265);
and U49491 (N_49491,N_42142,N_43732);
nand U49492 (N_49492,N_41563,N_42308);
xor U49493 (N_49493,N_43788,N_44314);
nand U49494 (N_49494,N_44600,N_42943);
and U49495 (N_49495,N_43568,N_43094);
xnor U49496 (N_49496,N_41539,N_40318);
nor U49497 (N_49497,N_40896,N_41234);
nor U49498 (N_49498,N_41297,N_40168);
nand U49499 (N_49499,N_43127,N_41929);
xnor U49500 (N_49500,N_41448,N_44319);
and U49501 (N_49501,N_40311,N_44091);
nand U49502 (N_49502,N_41967,N_42021);
and U49503 (N_49503,N_43713,N_40558);
nand U49504 (N_49504,N_44587,N_41864);
and U49505 (N_49505,N_40535,N_43865);
and U49506 (N_49506,N_41262,N_42309);
and U49507 (N_49507,N_42129,N_41437);
and U49508 (N_49508,N_42014,N_42824);
nor U49509 (N_49509,N_41105,N_41746);
nor U49510 (N_49510,N_43656,N_42423);
or U49511 (N_49511,N_40578,N_43081);
nor U49512 (N_49512,N_42699,N_44980);
or U49513 (N_49513,N_44569,N_44051);
xor U49514 (N_49514,N_42727,N_42492);
and U49515 (N_49515,N_42919,N_42870);
nor U49516 (N_49516,N_41974,N_40124);
xor U49517 (N_49517,N_44360,N_44420);
and U49518 (N_49518,N_43367,N_44101);
xor U49519 (N_49519,N_41205,N_44790);
nand U49520 (N_49520,N_42677,N_43306);
xor U49521 (N_49521,N_44841,N_40333);
xor U49522 (N_49522,N_42501,N_41848);
nand U49523 (N_49523,N_44341,N_40912);
and U49524 (N_49524,N_42159,N_41653);
nor U49525 (N_49525,N_43236,N_41081);
and U49526 (N_49526,N_40498,N_40187);
nand U49527 (N_49527,N_40650,N_41457);
or U49528 (N_49528,N_42368,N_43413);
nor U49529 (N_49529,N_42201,N_43710);
nand U49530 (N_49530,N_43815,N_44335);
nand U49531 (N_49531,N_40195,N_41790);
xor U49532 (N_49532,N_41956,N_41386);
and U49533 (N_49533,N_43505,N_41144);
xor U49534 (N_49534,N_40768,N_44488);
or U49535 (N_49535,N_41246,N_44935);
xor U49536 (N_49536,N_42389,N_43609);
nor U49537 (N_49537,N_42062,N_42518);
xnor U49538 (N_49538,N_40599,N_40904);
xor U49539 (N_49539,N_42328,N_42487);
xnor U49540 (N_49540,N_44687,N_40410);
xor U49541 (N_49541,N_41953,N_43521);
nor U49542 (N_49542,N_43762,N_43446);
or U49543 (N_49543,N_44109,N_41265);
nor U49544 (N_49544,N_43723,N_41079);
and U49545 (N_49545,N_44687,N_43659);
or U49546 (N_49546,N_43882,N_44331);
nor U49547 (N_49547,N_44611,N_43297);
and U49548 (N_49548,N_42087,N_43889);
nor U49549 (N_49549,N_44089,N_44940);
nand U49550 (N_49550,N_40516,N_44751);
xor U49551 (N_49551,N_40721,N_41391);
or U49552 (N_49552,N_43241,N_40988);
xnor U49553 (N_49553,N_42106,N_43344);
nor U49554 (N_49554,N_44868,N_43725);
nand U49555 (N_49555,N_40677,N_44817);
nand U49556 (N_49556,N_42529,N_40401);
nand U49557 (N_49557,N_41206,N_42333);
or U49558 (N_49558,N_44105,N_43062);
and U49559 (N_49559,N_43713,N_42398);
xor U49560 (N_49560,N_42549,N_43043);
xor U49561 (N_49561,N_40882,N_42575);
xor U49562 (N_49562,N_40744,N_40680);
and U49563 (N_49563,N_40245,N_40104);
and U49564 (N_49564,N_41917,N_40538);
nor U49565 (N_49565,N_44114,N_42327);
nor U49566 (N_49566,N_41865,N_43146);
and U49567 (N_49567,N_43733,N_42324);
nand U49568 (N_49568,N_44398,N_43423);
or U49569 (N_49569,N_40589,N_42520);
nand U49570 (N_49570,N_44874,N_41589);
xnor U49571 (N_49571,N_42737,N_41548);
or U49572 (N_49572,N_40000,N_42294);
and U49573 (N_49573,N_42028,N_43924);
xnor U49574 (N_49574,N_41267,N_40466);
and U49575 (N_49575,N_43410,N_44888);
xor U49576 (N_49576,N_43741,N_41023);
or U49577 (N_49577,N_40580,N_42627);
nor U49578 (N_49578,N_43474,N_44696);
or U49579 (N_49579,N_41957,N_43708);
and U49580 (N_49580,N_42027,N_42387);
or U49581 (N_49581,N_40135,N_42046);
xor U49582 (N_49582,N_40376,N_44184);
nand U49583 (N_49583,N_41274,N_43531);
nor U49584 (N_49584,N_42219,N_42532);
nor U49585 (N_49585,N_40272,N_43353);
xnor U49586 (N_49586,N_43500,N_43653);
or U49587 (N_49587,N_43896,N_41083);
nor U49588 (N_49588,N_43290,N_43709);
nor U49589 (N_49589,N_42895,N_44071);
nor U49590 (N_49590,N_44537,N_43343);
xnor U49591 (N_49591,N_44398,N_40430);
nand U49592 (N_49592,N_44813,N_41008);
nand U49593 (N_49593,N_44125,N_40016);
nor U49594 (N_49594,N_42800,N_43281);
nor U49595 (N_49595,N_42844,N_44557);
nand U49596 (N_49596,N_41660,N_43644);
xnor U49597 (N_49597,N_42400,N_43562);
or U49598 (N_49598,N_43221,N_42661);
nor U49599 (N_49599,N_40734,N_43374);
or U49600 (N_49600,N_44321,N_41836);
or U49601 (N_49601,N_42746,N_40449);
and U49602 (N_49602,N_42121,N_41174);
xor U49603 (N_49603,N_40709,N_40033);
and U49604 (N_49604,N_40385,N_43368);
nor U49605 (N_49605,N_41683,N_42434);
xnor U49606 (N_49606,N_42154,N_44847);
and U49607 (N_49607,N_42726,N_43334);
and U49608 (N_49608,N_42437,N_41085);
nand U49609 (N_49609,N_42297,N_40543);
nand U49610 (N_49610,N_40133,N_42313);
xor U49611 (N_49611,N_41809,N_40058);
or U49612 (N_49612,N_42235,N_43671);
nor U49613 (N_49613,N_42519,N_44751);
xor U49614 (N_49614,N_42869,N_43202);
nand U49615 (N_49615,N_44209,N_41723);
and U49616 (N_49616,N_43916,N_44059);
nor U49617 (N_49617,N_43275,N_44405);
and U49618 (N_49618,N_41686,N_41588);
or U49619 (N_49619,N_42313,N_42871);
or U49620 (N_49620,N_43398,N_42948);
and U49621 (N_49621,N_44516,N_44956);
or U49622 (N_49622,N_42411,N_44052);
and U49623 (N_49623,N_41466,N_42917);
nor U49624 (N_49624,N_42980,N_41084);
nand U49625 (N_49625,N_43495,N_41815);
and U49626 (N_49626,N_40040,N_44012);
nand U49627 (N_49627,N_41015,N_41190);
nand U49628 (N_49628,N_43066,N_41092);
or U49629 (N_49629,N_44044,N_43145);
xnor U49630 (N_49630,N_40300,N_44192);
or U49631 (N_49631,N_40955,N_42536);
and U49632 (N_49632,N_40980,N_42152);
or U49633 (N_49633,N_41935,N_40201);
nand U49634 (N_49634,N_41338,N_41305);
xor U49635 (N_49635,N_43327,N_42922);
xnor U49636 (N_49636,N_43432,N_42374);
and U49637 (N_49637,N_42043,N_43038);
nand U49638 (N_49638,N_43738,N_40320);
and U49639 (N_49639,N_43355,N_40689);
nor U49640 (N_49640,N_43113,N_40482);
nor U49641 (N_49641,N_40539,N_40796);
nor U49642 (N_49642,N_43582,N_40876);
nand U49643 (N_49643,N_44960,N_42429);
nand U49644 (N_49644,N_44810,N_43458);
xnor U49645 (N_49645,N_40287,N_44126);
xor U49646 (N_49646,N_42133,N_44921);
xnor U49647 (N_49647,N_41866,N_42347);
nand U49648 (N_49648,N_40179,N_40380);
nor U49649 (N_49649,N_42147,N_44108);
xor U49650 (N_49650,N_43985,N_42931);
nand U49651 (N_49651,N_40246,N_40410);
xnor U49652 (N_49652,N_42106,N_44320);
nand U49653 (N_49653,N_42362,N_44375);
nand U49654 (N_49654,N_42835,N_44996);
nand U49655 (N_49655,N_41093,N_41393);
xnor U49656 (N_49656,N_43831,N_44052);
and U49657 (N_49657,N_42938,N_40758);
and U49658 (N_49658,N_41494,N_41428);
nor U49659 (N_49659,N_43326,N_41320);
nor U49660 (N_49660,N_42368,N_43897);
or U49661 (N_49661,N_41449,N_43484);
nand U49662 (N_49662,N_44619,N_41834);
xnor U49663 (N_49663,N_42394,N_41157);
nand U49664 (N_49664,N_43533,N_42063);
or U49665 (N_49665,N_44856,N_44162);
and U49666 (N_49666,N_44505,N_44975);
and U49667 (N_49667,N_43136,N_43227);
and U49668 (N_49668,N_42223,N_42991);
nor U49669 (N_49669,N_44850,N_44957);
xnor U49670 (N_49670,N_41165,N_41709);
xnor U49671 (N_49671,N_43940,N_44109);
nor U49672 (N_49672,N_44715,N_44087);
nand U49673 (N_49673,N_43410,N_44514);
and U49674 (N_49674,N_41531,N_41735);
or U49675 (N_49675,N_42218,N_40200);
or U49676 (N_49676,N_41539,N_42347);
nand U49677 (N_49677,N_42525,N_42335);
or U49678 (N_49678,N_42890,N_42203);
nor U49679 (N_49679,N_41350,N_43514);
nor U49680 (N_49680,N_40016,N_42927);
nand U49681 (N_49681,N_43924,N_44707);
nand U49682 (N_49682,N_40194,N_43165);
xnor U49683 (N_49683,N_44920,N_44526);
or U49684 (N_49684,N_40598,N_40088);
or U49685 (N_49685,N_40303,N_44250);
nand U49686 (N_49686,N_40036,N_43951);
or U49687 (N_49687,N_42239,N_42939);
xor U49688 (N_49688,N_44154,N_44047);
and U49689 (N_49689,N_44529,N_44552);
xor U49690 (N_49690,N_41497,N_43778);
xor U49691 (N_49691,N_41626,N_44216);
and U49692 (N_49692,N_44152,N_40304);
nor U49693 (N_49693,N_41030,N_43645);
nor U49694 (N_49694,N_42988,N_42931);
or U49695 (N_49695,N_44003,N_41144);
nand U49696 (N_49696,N_42596,N_43346);
nand U49697 (N_49697,N_43104,N_44765);
or U49698 (N_49698,N_40471,N_40022);
nor U49699 (N_49699,N_44091,N_40049);
nor U49700 (N_49700,N_44647,N_40902);
and U49701 (N_49701,N_41251,N_43022);
nor U49702 (N_49702,N_44525,N_40652);
and U49703 (N_49703,N_44110,N_40406);
nor U49704 (N_49704,N_44268,N_40612);
or U49705 (N_49705,N_44364,N_44372);
nand U49706 (N_49706,N_41478,N_43238);
or U49707 (N_49707,N_41689,N_42334);
or U49708 (N_49708,N_44403,N_44078);
nor U49709 (N_49709,N_40737,N_40920);
nor U49710 (N_49710,N_43115,N_43876);
nand U49711 (N_49711,N_44633,N_42947);
xor U49712 (N_49712,N_42017,N_43614);
nand U49713 (N_49713,N_44044,N_41758);
and U49714 (N_49714,N_40020,N_42235);
and U49715 (N_49715,N_44284,N_42043);
nand U49716 (N_49716,N_40505,N_43835);
or U49717 (N_49717,N_44528,N_44806);
and U49718 (N_49718,N_40426,N_43112);
or U49719 (N_49719,N_43086,N_42176);
nand U49720 (N_49720,N_41956,N_42012);
nor U49721 (N_49721,N_44259,N_40630);
nand U49722 (N_49722,N_42845,N_40756);
nand U49723 (N_49723,N_40763,N_42835);
and U49724 (N_49724,N_40580,N_41247);
and U49725 (N_49725,N_41621,N_43446);
xnor U49726 (N_49726,N_44956,N_41989);
or U49727 (N_49727,N_44691,N_43979);
and U49728 (N_49728,N_43056,N_43262);
and U49729 (N_49729,N_43291,N_44828);
or U49730 (N_49730,N_43295,N_41942);
or U49731 (N_49731,N_40334,N_43079);
nor U49732 (N_49732,N_44632,N_41349);
and U49733 (N_49733,N_42802,N_44585);
nand U49734 (N_49734,N_40714,N_41863);
or U49735 (N_49735,N_43849,N_41784);
nand U49736 (N_49736,N_42646,N_40908);
nand U49737 (N_49737,N_40411,N_40691);
or U49738 (N_49738,N_43764,N_44245);
nand U49739 (N_49739,N_43943,N_41274);
nor U49740 (N_49740,N_44518,N_40452);
xor U49741 (N_49741,N_43326,N_44584);
nor U49742 (N_49742,N_41240,N_41329);
or U49743 (N_49743,N_42534,N_41691);
nand U49744 (N_49744,N_44754,N_43479);
and U49745 (N_49745,N_44565,N_41298);
xnor U49746 (N_49746,N_43393,N_41447);
nor U49747 (N_49747,N_43735,N_43116);
xor U49748 (N_49748,N_41436,N_40762);
or U49749 (N_49749,N_42300,N_44485);
or U49750 (N_49750,N_40616,N_41914);
nand U49751 (N_49751,N_41455,N_44934);
and U49752 (N_49752,N_44003,N_43479);
xor U49753 (N_49753,N_42845,N_42697);
and U49754 (N_49754,N_42416,N_40820);
or U49755 (N_49755,N_40075,N_43824);
and U49756 (N_49756,N_43532,N_43231);
and U49757 (N_49757,N_40994,N_41608);
nand U49758 (N_49758,N_40944,N_43610);
nand U49759 (N_49759,N_41153,N_44973);
nand U49760 (N_49760,N_44504,N_40584);
and U49761 (N_49761,N_43982,N_44703);
or U49762 (N_49762,N_43873,N_42684);
nor U49763 (N_49763,N_41468,N_43258);
or U49764 (N_49764,N_43063,N_44411);
xor U49765 (N_49765,N_41886,N_42374);
nor U49766 (N_49766,N_40382,N_42325);
or U49767 (N_49767,N_40851,N_41916);
xor U49768 (N_49768,N_41328,N_42606);
and U49769 (N_49769,N_41753,N_42050);
xor U49770 (N_49770,N_44825,N_42472);
nor U49771 (N_49771,N_40023,N_41604);
and U49772 (N_49772,N_41792,N_40100);
xor U49773 (N_49773,N_40947,N_40194);
and U49774 (N_49774,N_43171,N_44572);
xnor U49775 (N_49775,N_42310,N_42739);
and U49776 (N_49776,N_44790,N_41771);
nor U49777 (N_49777,N_44092,N_44358);
nand U49778 (N_49778,N_41071,N_43184);
or U49779 (N_49779,N_44037,N_42797);
or U49780 (N_49780,N_41949,N_43553);
or U49781 (N_49781,N_44578,N_43319);
nand U49782 (N_49782,N_40824,N_40484);
nor U49783 (N_49783,N_43089,N_40947);
xnor U49784 (N_49784,N_40257,N_40143);
and U49785 (N_49785,N_44303,N_42251);
and U49786 (N_49786,N_42113,N_44952);
nand U49787 (N_49787,N_40668,N_40260);
nor U49788 (N_49788,N_41664,N_43521);
nor U49789 (N_49789,N_41067,N_40206);
nand U49790 (N_49790,N_41214,N_40441);
nand U49791 (N_49791,N_44930,N_42707);
and U49792 (N_49792,N_42691,N_42128);
nor U49793 (N_49793,N_44351,N_42006);
or U49794 (N_49794,N_44447,N_44559);
or U49795 (N_49795,N_42848,N_41008);
and U49796 (N_49796,N_40169,N_40263);
nand U49797 (N_49797,N_43583,N_43104);
or U49798 (N_49798,N_41764,N_40826);
and U49799 (N_49799,N_41575,N_42237);
nand U49800 (N_49800,N_40933,N_42893);
and U49801 (N_49801,N_43427,N_40737);
nor U49802 (N_49802,N_41683,N_44883);
or U49803 (N_49803,N_40174,N_41693);
xor U49804 (N_49804,N_40826,N_42169);
xor U49805 (N_49805,N_41246,N_42329);
and U49806 (N_49806,N_42613,N_40671);
and U49807 (N_49807,N_41283,N_40021);
nand U49808 (N_49808,N_43542,N_44198);
xor U49809 (N_49809,N_43133,N_42552);
xnor U49810 (N_49810,N_41762,N_42956);
and U49811 (N_49811,N_40896,N_44605);
nor U49812 (N_49812,N_43847,N_41737);
nand U49813 (N_49813,N_42152,N_43985);
or U49814 (N_49814,N_44706,N_43097);
and U49815 (N_49815,N_43944,N_42807);
nand U49816 (N_49816,N_40890,N_40016);
nor U49817 (N_49817,N_42141,N_42877);
nor U49818 (N_49818,N_44405,N_41340);
xor U49819 (N_49819,N_44803,N_41594);
and U49820 (N_49820,N_44222,N_43491);
nor U49821 (N_49821,N_42006,N_42355);
nor U49822 (N_49822,N_43471,N_42330);
or U49823 (N_49823,N_44698,N_42672);
nand U49824 (N_49824,N_40275,N_44307);
nor U49825 (N_49825,N_40976,N_44535);
or U49826 (N_49826,N_43442,N_41751);
nand U49827 (N_49827,N_43990,N_44285);
or U49828 (N_49828,N_43603,N_42283);
xnor U49829 (N_49829,N_44397,N_44260);
or U49830 (N_49830,N_40969,N_40349);
nand U49831 (N_49831,N_44618,N_43522);
nand U49832 (N_49832,N_41236,N_42443);
nor U49833 (N_49833,N_44695,N_43436);
nor U49834 (N_49834,N_41483,N_40696);
and U49835 (N_49835,N_43032,N_44111);
nand U49836 (N_49836,N_43947,N_44384);
xor U49837 (N_49837,N_43453,N_44131);
xnor U49838 (N_49838,N_43410,N_44255);
nor U49839 (N_49839,N_43061,N_42067);
or U49840 (N_49840,N_44583,N_43242);
xor U49841 (N_49841,N_41276,N_44729);
or U49842 (N_49842,N_44788,N_40183);
nand U49843 (N_49843,N_43646,N_44004);
and U49844 (N_49844,N_40013,N_40864);
and U49845 (N_49845,N_41859,N_40422);
xor U49846 (N_49846,N_41889,N_43913);
nor U49847 (N_49847,N_43617,N_43022);
and U49848 (N_49848,N_40367,N_40954);
and U49849 (N_49849,N_43990,N_42654);
nor U49850 (N_49850,N_44165,N_41714);
or U49851 (N_49851,N_43592,N_43978);
nor U49852 (N_49852,N_41693,N_44434);
and U49853 (N_49853,N_41837,N_44784);
nor U49854 (N_49854,N_44745,N_43139);
nor U49855 (N_49855,N_43279,N_44264);
nor U49856 (N_49856,N_44173,N_44702);
xor U49857 (N_49857,N_40848,N_41462);
nor U49858 (N_49858,N_41139,N_42497);
and U49859 (N_49859,N_41171,N_42102);
xnor U49860 (N_49860,N_44864,N_42968);
and U49861 (N_49861,N_42894,N_44580);
nor U49862 (N_49862,N_40864,N_40052);
or U49863 (N_49863,N_43338,N_43556);
nor U49864 (N_49864,N_43873,N_41791);
or U49865 (N_49865,N_41481,N_44939);
nand U49866 (N_49866,N_42582,N_43300);
nand U49867 (N_49867,N_41671,N_44863);
xnor U49868 (N_49868,N_40327,N_43944);
or U49869 (N_49869,N_41101,N_42651);
and U49870 (N_49870,N_43565,N_44105);
nor U49871 (N_49871,N_40757,N_42274);
and U49872 (N_49872,N_40897,N_44552);
and U49873 (N_49873,N_40455,N_43604);
or U49874 (N_49874,N_43176,N_42221);
xor U49875 (N_49875,N_41285,N_40092);
and U49876 (N_49876,N_41863,N_43055);
and U49877 (N_49877,N_41585,N_42355);
or U49878 (N_49878,N_41781,N_43934);
nor U49879 (N_49879,N_41347,N_43095);
or U49880 (N_49880,N_40080,N_40871);
and U49881 (N_49881,N_40202,N_40684);
nand U49882 (N_49882,N_40208,N_42461);
and U49883 (N_49883,N_43382,N_41683);
xnor U49884 (N_49884,N_41888,N_44468);
or U49885 (N_49885,N_40929,N_44299);
and U49886 (N_49886,N_40747,N_41659);
xnor U49887 (N_49887,N_42210,N_42601);
or U49888 (N_49888,N_44676,N_43726);
and U49889 (N_49889,N_44339,N_40796);
nand U49890 (N_49890,N_44198,N_43728);
nand U49891 (N_49891,N_43460,N_40915);
nand U49892 (N_49892,N_41615,N_43415);
nor U49893 (N_49893,N_41165,N_42530);
and U49894 (N_49894,N_42660,N_44041);
and U49895 (N_49895,N_42911,N_42805);
xnor U49896 (N_49896,N_43012,N_40710);
or U49897 (N_49897,N_42815,N_42659);
and U49898 (N_49898,N_41557,N_43668);
or U49899 (N_49899,N_44321,N_41169);
xor U49900 (N_49900,N_43785,N_41061);
and U49901 (N_49901,N_43656,N_43176);
xnor U49902 (N_49902,N_41832,N_41279);
xnor U49903 (N_49903,N_44998,N_42187);
nor U49904 (N_49904,N_41069,N_41505);
nor U49905 (N_49905,N_42259,N_43837);
xnor U49906 (N_49906,N_44487,N_42217);
and U49907 (N_49907,N_42192,N_40830);
and U49908 (N_49908,N_44262,N_42675);
nand U49909 (N_49909,N_42092,N_40681);
nand U49910 (N_49910,N_41766,N_40853);
xor U49911 (N_49911,N_40674,N_40814);
nor U49912 (N_49912,N_41425,N_44087);
and U49913 (N_49913,N_43544,N_43104);
and U49914 (N_49914,N_44285,N_40185);
xnor U49915 (N_49915,N_44045,N_43176);
and U49916 (N_49916,N_42191,N_41593);
or U49917 (N_49917,N_42465,N_41573);
xor U49918 (N_49918,N_43606,N_40718);
and U49919 (N_49919,N_42735,N_44711);
or U49920 (N_49920,N_41776,N_41862);
nor U49921 (N_49921,N_40820,N_44401);
or U49922 (N_49922,N_41972,N_44294);
xnor U49923 (N_49923,N_41846,N_42030);
or U49924 (N_49924,N_43366,N_41475);
and U49925 (N_49925,N_40979,N_44367);
nor U49926 (N_49926,N_40138,N_42416);
nor U49927 (N_49927,N_43398,N_40634);
and U49928 (N_49928,N_43727,N_41684);
nand U49929 (N_49929,N_43352,N_44249);
nor U49930 (N_49930,N_42579,N_44094);
nand U49931 (N_49931,N_42786,N_43693);
xor U49932 (N_49932,N_43783,N_40985);
or U49933 (N_49933,N_44261,N_41677);
nor U49934 (N_49934,N_40452,N_44477);
nor U49935 (N_49935,N_43503,N_41484);
nor U49936 (N_49936,N_40237,N_40831);
nor U49937 (N_49937,N_43598,N_40834);
nor U49938 (N_49938,N_42673,N_44733);
xnor U49939 (N_49939,N_43512,N_41182);
xnor U49940 (N_49940,N_41606,N_43214);
and U49941 (N_49941,N_41939,N_40186);
nand U49942 (N_49942,N_40706,N_43706);
or U49943 (N_49943,N_41739,N_41460);
or U49944 (N_49944,N_42567,N_40649);
nor U49945 (N_49945,N_41612,N_43626);
nor U49946 (N_49946,N_40454,N_40259);
nor U49947 (N_49947,N_43437,N_42611);
and U49948 (N_49948,N_43842,N_44129);
nor U49949 (N_49949,N_41355,N_41989);
nor U49950 (N_49950,N_42673,N_40222);
nor U49951 (N_49951,N_43054,N_41988);
nand U49952 (N_49952,N_44944,N_44156);
or U49953 (N_49953,N_43468,N_44386);
or U49954 (N_49954,N_41418,N_40831);
xor U49955 (N_49955,N_40119,N_42471);
or U49956 (N_49956,N_43117,N_42819);
or U49957 (N_49957,N_42325,N_40844);
and U49958 (N_49958,N_44598,N_41682);
nand U49959 (N_49959,N_40664,N_44091);
nand U49960 (N_49960,N_42693,N_44413);
or U49961 (N_49961,N_40561,N_42854);
nor U49962 (N_49962,N_41050,N_41499);
nor U49963 (N_49963,N_40895,N_43807);
nand U49964 (N_49964,N_43720,N_40580);
nor U49965 (N_49965,N_40786,N_44258);
nand U49966 (N_49966,N_44521,N_40941);
xnor U49967 (N_49967,N_40193,N_41261);
and U49968 (N_49968,N_43591,N_41595);
and U49969 (N_49969,N_42614,N_43755);
nor U49970 (N_49970,N_44828,N_44958);
nor U49971 (N_49971,N_44643,N_42030);
nor U49972 (N_49972,N_40912,N_42004);
or U49973 (N_49973,N_44126,N_41729);
or U49974 (N_49974,N_41296,N_41462);
and U49975 (N_49975,N_40979,N_40790);
nand U49976 (N_49976,N_41255,N_43168);
and U49977 (N_49977,N_42058,N_41263);
and U49978 (N_49978,N_40227,N_44721);
or U49979 (N_49979,N_44342,N_41009);
or U49980 (N_49980,N_41700,N_44889);
nor U49981 (N_49981,N_44587,N_42329);
nand U49982 (N_49982,N_42503,N_42533);
or U49983 (N_49983,N_43805,N_44753);
and U49984 (N_49984,N_43552,N_43871);
and U49985 (N_49985,N_43179,N_43708);
nor U49986 (N_49986,N_40017,N_41828);
nor U49987 (N_49987,N_41700,N_44737);
xnor U49988 (N_49988,N_43409,N_44640);
nor U49989 (N_49989,N_42408,N_40677);
nand U49990 (N_49990,N_42587,N_44173);
and U49991 (N_49991,N_41438,N_41645);
and U49992 (N_49992,N_43198,N_44161);
nor U49993 (N_49993,N_44981,N_43591);
nand U49994 (N_49994,N_42469,N_40640);
nand U49995 (N_49995,N_42133,N_41356);
xor U49996 (N_49996,N_40594,N_43523);
or U49997 (N_49997,N_43253,N_40245);
and U49998 (N_49998,N_40096,N_44670);
nand U49999 (N_49999,N_43025,N_44864);
nand UO_0 (O_0,N_47022,N_48449);
xnor UO_1 (O_1,N_49941,N_49574);
and UO_2 (O_2,N_47927,N_45341);
and UO_3 (O_3,N_47143,N_46920);
nand UO_4 (O_4,N_49079,N_45885);
and UO_5 (O_5,N_48947,N_47170);
nor UO_6 (O_6,N_45588,N_48456);
and UO_7 (O_7,N_46647,N_49255);
and UO_8 (O_8,N_48338,N_49405);
xnor UO_9 (O_9,N_49608,N_49025);
and UO_10 (O_10,N_45016,N_45519);
nand UO_11 (O_11,N_47919,N_45658);
nand UO_12 (O_12,N_49174,N_45955);
or UO_13 (O_13,N_48157,N_45175);
xor UO_14 (O_14,N_49814,N_45534);
xnor UO_15 (O_15,N_45582,N_46852);
xor UO_16 (O_16,N_45418,N_46485);
nor UO_17 (O_17,N_45265,N_48336);
nor UO_18 (O_18,N_45893,N_49873);
nor UO_19 (O_19,N_48598,N_45493);
nor UO_20 (O_20,N_48906,N_49224);
or UO_21 (O_21,N_46011,N_45567);
nand UO_22 (O_22,N_48039,N_47419);
nand UO_23 (O_23,N_45252,N_47522);
nand UO_24 (O_24,N_48396,N_46827);
xor UO_25 (O_25,N_47724,N_45335);
nor UO_26 (O_26,N_49508,N_49301);
and UO_27 (O_27,N_46550,N_47381);
and UO_28 (O_28,N_45507,N_49982);
nand UO_29 (O_29,N_46951,N_48724);
xnor UO_30 (O_30,N_49577,N_48193);
and UO_31 (O_31,N_46947,N_46790);
and UO_32 (O_32,N_46090,N_47227);
nand UO_33 (O_33,N_47979,N_49695);
nor UO_34 (O_34,N_45954,N_47035);
or UO_35 (O_35,N_46955,N_49893);
nand UO_36 (O_36,N_48965,N_47192);
and UO_37 (O_37,N_47161,N_47693);
nor UO_38 (O_38,N_46361,N_46423);
and UO_39 (O_39,N_46813,N_46718);
or UO_40 (O_40,N_49402,N_49753);
xnor UO_41 (O_41,N_49961,N_46892);
nor UO_42 (O_42,N_49864,N_45553);
nand UO_43 (O_43,N_46482,N_48446);
xor UO_44 (O_44,N_49113,N_49259);
nand UO_45 (O_45,N_48458,N_47416);
xnor UO_46 (O_46,N_46948,N_47972);
xor UO_47 (O_47,N_45200,N_46703);
or UO_48 (O_48,N_47296,N_48326);
xor UO_49 (O_49,N_49926,N_49112);
and UO_50 (O_50,N_48876,N_49850);
xnor UO_51 (O_51,N_46379,N_47073);
and UO_52 (O_52,N_45443,N_48240);
or UO_53 (O_53,N_47696,N_49005);
nand UO_54 (O_54,N_45469,N_49016);
xnor UO_55 (O_55,N_45634,N_45540);
and UO_56 (O_56,N_48806,N_48636);
nor UO_57 (O_57,N_46979,N_45239);
nand UO_58 (O_58,N_49952,N_45967);
xnor UO_59 (O_59,N_46987,N_49258);
nand UO_60 (O_60,N_47313,N_46152);
nand UO_61 (O_61,N_49871,N_47141);
and UO_62 (O_62,N_47831,N_47189);
xor UO_63 (O_63,N_49249,N_49722);
nor UO_64 (O_64,N_48923,N_45213);
nor UO_65 (O_65,N_46704,N_48090);
and UO_66 (O_66,N_46507,N_45691);
nor UO_67 (O_67,N_48773,N_47753);
nand UO_68 (O_68,N_45746,N_47262);
nor UO_69 (O_69,N_45836,N_49392);
nand UO_70 (O_70,N_47656,N_46083);
nand UO_71 (O_71,N_49180,N_49665);
and UO_72 (O_72,N_49832,N_45502);
nor UO_73 (O_73,N_49037,N_46949);
xnor UO_74 (O_74,N_46742,N_46172);
and UO_75 (O_75,N_47437,N_45703);
nand UO_76 (O_76,N_46405,N_45161);
nor UO_77 (O_77,N_48627,N_45512);
or UO_78 (O_78,N_46092,N_48436);
nand UO_79 (O_79,N_47238,N_47671);
and UO_80 (O_80,N_46097,N_48596);
or UO_81 (O_81,N_48179,N_49707);
and UO_82 (O_82,N_48382,N_46942);
or UO_83 (O_83,N_45310,N_49983);
and UO_84 (O_84,N_48614,N_46546);
and UO_85 (O_85,N_48303,N_46102);
nand UO_86 (O_86,N_46241,N_46262);
or UO_87 (O_87,N_46660,N_45420);
or UO_88 (O_88,N_47020,N_45759);
or UO_89 (O_89,N_46671,N_49976);
or UO_90 (O_90,N_47925,N_47074);
and UO_91 (O_91,N_48873,N_46478);
nand UO_92 (O_92,N_45145,N_46940);
xor UO_93 (O_93,N_47249,N_46815);
xor UO_94 (O_94,N_48025,N_48891);
nor UO_95 (O_95,N_46196,N_45218);
nand UO_96 (O_96,N_47835,N_45078);
xor UO_97 (O_97,N_48710,N_45586);
or UO_98 (O_98,N_46394,N_48853);
nand UO_99 (O_99,N_45521,N_48212);
and UO_100 (O_100,N_49472,N_46508);
nand UO_101 (O_101,N_48500,N_46571);
xnor UO_102 (O_102,N_48694,N_46359);
nor UO_103 (O_103,N_48073,N_47991);
and UO_104 (O_104,N_46716,N_48572);
nor UO_105 (O_105,N_46329,N_45255);
nand UO_106 (O_106,N_45049,N_45854);
nor UO_107 (O_107,N_46182,N_48444);
and UO_108 (O_108,N_45777,N_49383);
nor UO_109 (O_109,N_46975,N_46213);
and UO_110 (O_110,N_46766,N_48824);
xnor UO_111 (O_111,N_48316,N_48644);
and UO_112 (O_112,N_48922,N_45160);
nor UO_113 (O_113,N_45392,N_47644);
nor UO_114 (O_114,N_45610,N_46270);
nand UO_115 (O_115,N_47006,N_47038);
or UO_116 (O_116,N_46653,N_49422);
or UO_117 (O_117,N_49043,N_47534);
nor UO_118 (O_118,N_47001,N_46166);
or UO_119 (O_119,N_46226,N_47108);
and UO_120 (O_120,N_46014,N_46500);
and UO_121 (O_121,N_47078,N_47316);
nand UO_122 (O_122,N_45504,N_49784);
and UO_123 (O_123,N_46958,N_46617);
nor UO_124 (O_124,N_47795,N_47590);
and UO_125 (O_125,N_48419,N_47362);
nand UO_126 (O_126,N_49008,N_45071);
or UO_127 (O_127,N_45859,N_48526);
nand UO_128 (O_128,N_46125,N_46689);
and UO_129 (O_129,N_45959,N_47700);
nand UO_130 (O_130,N_49721,N_46695);
nor UO_131 (O_131,N_49783,N_47737);
or UO_132 (O_132,N_48994,N_48606);
xnor UO_133 (O_133,N_45452,N_47819);
and UO_134 (O_134,N_48224,N_46927);
nor UO_135 (O_135,N_46242,N_48631);
and UO_136 (O_136,N_45989,N_47286);
and UO_137 (O_137,N_45794,N_47946);
and UO_138 (O_138,N_48677,N_47789);
nor UO_139 (O_139,N_49662,N_45375);
xnor UO_140 (O_140,N_48898,N_46491);
or UO_141 (O_141,N_49892,N_46877);
or UO_142 (O_142,N_47360,N_46786);
xnor UO_143 (O_143,N_46407,N_48159);
or UO_144 (O_144,N_49275,N_45915);
or UO_145 (O_145,N_49126,N_48187);
and UO_146 (O_146,N_49208,N_48675);
or UO_147 (O_147,N_47175,N_47486);
xnor UO_148 (O_148,N_48542,N_47081);
nand UO_149 (O_149,N_46227,N_47276);
xnor UO_150 (O_150,N_45370,N_49423);
xnor UO_151 (O_151,N_49364,N_47312);
nand UO_152 (O_152,N_48975,N_49884);
nor UO_153 (O_153,N_45414,N_46572);
nand UO_154 (O_154,N_46749,N_47428);
xor UO_155 (O_155,N_46103,N_46380);
and UO_156 (O_156,N_47767,N_48155);
xnor UO_157 (O_157,N_46128,N_47202);
xnor UO_158 (O_158,N_46882,N_45640);
nor UO_159 (O_159,N_48678,N_49420);
nand UO_160 (O_160,N_48190,N_48993);
nand UO_161 (O_161,N_48652,N_49847);
nor UO_162 (O_162,N_49800,N_46952);
xor UO_163 (O_163,N_49481,N_47910);
or UO_164 (O_164,N_48253,N_45972);
nand UO_165 (O_165,N_48924,N_47197);
nand UO_166 (O_166,N_49311,N_47114);
and UO_167 (O_167,N_49750,N_48028);
and UO_168 (O_168,N_46957,N_47063);
xor UO_169 (O_169,N_49936,N_49973);
nand UO_170 (O_170,N_46510,N_49903);
or UO_171 (O_171,N_47587,N_48474);
or UO_172 (O_172,N_48378,N_47032);
and UO_173 (O_173,N_47666,N_47096);
and UO_174 (O_174,N_46116,N_47931);
or UO_175 (O_175,N_48388,N_49457);
and UO_176 (O_176,N_45075,N_49082);
and UO_177 (O_177,N_47068,N_46086);
xnor UO_178 (O_178,N_46669,N_45681);
nor UO_179 (O_179,N_47278,N_48881);
or UO_180 (O_180,N_46576,N_46526);
xor UO_181 (O_181,N_48620,N_49188);
or UO_182 (O_182,N_48697,N_46169);
nor UO_183 (O_183,N_47889,N_45224);
and UO_184 (O_184,N_46739,N_45251);
nand UO_185 (O_185,N_47990,N_48805);
or UO_186 (O_186,N_49621,N_46818);
and UO_187 (O_187,N_45987,N_45867);
xor UO_188 (O_188,N_48086,N_48418);
or UO_189 (O_189,N_46186,N_48580);
and UO_190 (O_190,N_46401,N_46791);
nor UO_191 (O_191,N_46627,N_48012);
xor UO_192 (O_192,N_48768,N_49114);
nand UO_193 (O_193,N_48935,N_45608);
or UO_194 (O_194,N_45063,N_47564);
nand UO_195 (O_195,N_47824,N_45424);
or UO_196 (O_196,N_49388,N_49632);
and UO_197 (O_197,N_48814,N_48549);
xnor UO_198 (O_198,N_46613,N_46972);
nand UO_199 (O_199,N_45587,N_49195);
xnor UO_200 (O_200,N_49416,N_49116);
and UO_201 (O_201,N_46495,N_49849);
nand UO_202 (O_202,N_49386,N_46980);
nor UO_203 (O_203,N_49379,N_48988);
nand UO_204 (O_204,N_49561,N_46006);
or UO_205 (O_205,N_47691,N_49261);
nand UO_206 (O_206,N_46537,N_47011);
and UO_207 (O_207,N_49914,N_47764);
nand UO_208 (O_208,N_47475,N_46604);
nor UO_209 (O_209,N_45481,N_47476);
and UO_210 (O_210,N_46875,N_47040);
nor UO_211 (O_211,N_49857,N_46734);
or UO_212 (O_212,N_49504,N_45296);
nand UO_213 (O_213,N_48173,N_46301);
nand UO_214 (O_214,N_48750,N_46905);
xor UO_215 (O_215,N_49466,N_48461);
xor UO_216 (O_216,N_48793,N_46878);
nand UO_217 (O_217,N_48639,N_45739);
and UO_218 (O_218,N_49763,N_45377);
or UO_219 (O_219,N_45283,N_46857);
nor UO_220 (O_220,N_49128,N_49776);
and UO_221 (O_221,N_48566,N_47023);
and UO_222 (O_222,N_49162,N_47290);
and UO_223 (O_223,N_46352,N_47086);
xor UO_224 (O_224,N_48995,N_47817);
xor UO_225 (O_225,N_49532,N_46904);
and UO_226 (O_226,N_46838,N_49524);
and UO_227 (O_227,N_48297,N_45520);
or UO_228 (O_228,N_48331,N_46767);
nor UO_229 (O_229,N_48719,N_49173);
and UO_230 (O_230,N_47525,N_46305);
and UO_231 (O_231,N_46364,N_49506);
or UO_232 (O_232,N_49501,N_46035);
nor UO_233 (O_233,N_46474,N_47460);
nand UO_234 (O_234,N_47779,N_45128);
or UO_235 (O_235,N_46117,N_47709);
nor UO_236 (O_236,N_46966,N_45118);
nand UO_237 (O_237,N_47222,N_46907);
nand UO_238 (O_238,N_46265,N_48539);
and UO_239 (O_239,N_46012,N_48105);
nor UO_240 (O_240,N_49478,N_48040);
xnor UO_241 (O_241,N_48348,N_45108);
and UO_242 (O_242,N_49748,N_47256);
nor UO_243 (O_243,N_47966,N_49705);
or UO_244 (O_244,N_47399,N_46712);
and UO_245 (O_245,N_45004,N_49339);
nand UO_246 (O_246,N_48963,N_47639);
nand UO_247 (O_247,N_49980,N_46637);
or UO_248 (O_248,N_46831,N_45548);
and UO_249 (O_249,N_46466,N_48912);
xnor UO_250 (O_250,N_47037,N_47593);
and UO_251 (O_251,N_49634,N_49734);
nor UO_252 (O_252,N_46315,N_47388);
nand UO_253 (O_253,N_47548,N_48797);
and UO_254 (O_254,N_46538,N_49684);
nand UO_255 (O_255,N_46559,N_47341);
nor UO_256 (O_256,N_46009,N_46177);
and UO_257 (O_257,N_46887,N_49266);
xor UO_258 (O_258,N_49670,N_45349);
xor UO_259 (O_259,N_48521,N_47883);
nand UO_260 (O_260,N_47214,N_45646);
nand UO_261 (O_261,N_45358,N_49288);
nor UO_262 (O_262,N_46414,N_49842);
nand UO_263 (O_263,N_47766,N_47251);
nand UO_264 (O_264,N_48263,N_49635);
nand UO_265 (O_265,N_46017,N_48133);
nor UO_266 (O_266,N_46280,N_47849);
xnor UO_267 (O_267,N_47224,N_46098);
nand UO_268 (O_268,N_48037,N_46354);
nor UO_269 (O_269,N_46341,N_45483);
or UO_270 (O_270,N_48299,N_46038);
and UO_271 (O_271,N_48200,N_48358);
nor UO_272 (O_272,N_46385,N_48546);
nor UO_273 (O_273,N_49744,N_45602);
nand UO_274 (O_274,N_47894,N_47259);
and UO_275 (O_275,N_49889,N_45581);
or UO_276 (O_276,N_48967,N_45393);
or UO_277 (O_277,N_46434,N_48269);
nor UO_278 (O_278,N_49579,N_47390);
nor UO_279 (O_279,N_45735,N_46454);
xnor UO_280 (O_280,N_46614,N_45242);
xnor UO_281 (O_281,N_45912,N_47859);
xnor UO_282 (O_282,N_49046,N_47716);
nor UO_283 (O_283,N_47368,N_45903);
nor UO_284 (O_284,N_47075,N_45917);
xnor UO_285 (O_285,N_47225,N_48953);
and UO_286 (O_286,N_46939,N_45665);
and UO_287 (O_287,N_48001,N_46594);
nor UO_288 (O_288,N_47595,N_45355);
nor UO_289 (O_289,N_49841,N_45147);
and UO_290 (O_290,N_47461,N_48060);
and UO_291 (O_291,N_46593,N_47828);
or UO_292 (O_292,N_46457,N_47790);
nand UO_293 (O_293,N_46238,N_48648);
and UO_294 (O_294,N_45883,N_49446);
nand UO_295 (O_295,N_45829,N_46727);
nor UO_296 (O_296,N_49764,N_45121);
or UO_297 (O_297,N_47483,N_49024);
xor UO_298 (O_298,N_49026,N_45659);
xor UO_299 (O_299,N_45523,N_48587);
nor UO_300 (O_300,N_47999,N_49071);
nand UO_301 (O_301,N_49681,N_45998);
nor UO_302 (O_302,N_46597,N_49434);
nand UO_303 (O_303,N_45828,N_47855);
nor UO_304 (O_304,N_49310,N_48799);
nand UO_305 (O_305,N_48296,N_45130);
nand UO_306 (O_306,N_46105,N_45485);
nor UO_307 (O_307,N_45573,N_48616);
or UO_308 (O_308,N_48279,N_47447);
and UO_309 (O_309,N_45473,N_45804);
and UO_310 (O_310,N_45497,N_47097);
xnor UO_311 (O_311,N_45457,N_45631);
nor UO_312 (O_312,N_48385,N_49384);
nor UO_313 (O_313,N_45053,N_45231);
nand UO_314 (O_314,N_46570,N_47794);
nand UO_315 (O_315,N_48513,N_48264);
nand UO_316 (O_316,N_49555,N_49751);
nor UO_317 (O_317,N_46568,N_47029);
nor UO_318 (O_318,N_45192,N_49916);
nor UO_319 (O_319,N_48051,N_46475);
nand UO_320 (O_320,N_48381,N_49771);
xnor UO_321 (O_321,N_47203,N_49158);
nor UO_322 (O_322,N_45280,N_45228);
nand UO_323 (O_323,N_49804,N_45708);
nand UO_324 (O_324,N_48803,N_46312);
and UO_325 (O_325,N_45813,N_48150);
xor UO_326 (O_326,N_48579,N_48445);
nor UO_327 (O_327,N_45527,N_46112);
or UO_328 (O_328,N_45333,N_48515);
nand UO_329 (O_329,N_49161,N_46525);
nand UO_330 (O_330,N_45660,N_47206);
nor UO_331 (O_331,N_48680,N_49051);
xnor UO_332 (O_332,N_47705,N_49318);
xnor UO_333 (O_333,N_47961,N_45788);
or UO_334 (O_334,N_48091,N_48158);
nor UO_335 (O_335,N_46591,N_47007);
or UO_336 (O_336,N_46504,N_48266);
or UO_337 (O_337,N_47338,N_45918);
and UO_338 (O_338,N_45749,N_48076);
xor UO_339 (O_339,N_46677,N_49290);
nor UO_340 (O_340,N_46517,N_48682);
nor UO_341 (O_341,N_45680,N_47746);
nand UO_342 (O_342,N_49510,N_46416);
nand UO_343 (O_343,N_49595,N_46626);
or UO_344 (O_344,N_48543,N_46258);
or UO_345 (O_345,N_49152,N_46473);
and UO_346 (O_346,N_46839,N_45058);
nor UO_347 (O_347,N_47048,N_46427);
nand UO_348 (O_348,N_48071,N_47757);
or UO_349 (O_349,N_48392,N_48576);
and UO_350 (O_350,N_47721,N_47787);
nand UO_351 (O_351,N_47454,N_45402);
nor UO_352 (O_352,N_46319,N_47344);
or UO_353 (O_353,N_46409,N_49337);
nand UO_354 (O_354,N_48477,N_48490);
and UO_355 (O_355,N_49709,N_48555);
or UO_356 (O_356,N_49436,N_45704);
nor UO_357 (O_357,N_49792,N_46350);
or UO_358 (O_358,N_48172,N_49556);
xor UO_359 (O_359,N_46174,N_48270);
xnor UO_360 (O_360,N_49756,N_45546);
xnor UO_361 (O_361,N_46846,N_45720);
nand UO_362 (O_362,N_49592,N_48826);
and UO_363 (O_363,N_45929,N_47536);
and UO_364 (O_364,N_46567,N_49846);
and UO_365 (O_365,N_45115,N_49716);
nor UO_366 (O_366,N_46708,N_46228);
nor UO_367 (O_367,N_49115,N_45041);
nand UO_368 (O_368,N_47780,N_47234);
and UO_369 (O_369,N_45734,N_46619);
xor UO_370 (O_370,N_48763,N_49435);
nand UO_371 (O_371,N_49359,N_45189);
and UO_372 (O_372,N_48689,N_46002);
nand UO_373 (O_373,N_48504,N_48919);
or UO_374 (O_374,N_46119,N_46901);
nand UO_375 (O_375,N_49187,N_46865);
nand UO_376 (O_376,N_45795,N_45315);
nor UO_377 (O_377,N_47403,N_47150);
or UO_378 (O_378,N_46200,N_45193);
nand UO_379 (O_379,N_48292,N_47643);
nor UO_380 (O_380,N_48769,N_46726);
nor UO_381 (O_381,N_45090,N_49937);
xnor UO_382 (O_382,N_49262,N_45206);
nand UO_383 (O_383,N_46498,N_47535);
and UO_384 (O_384,N_45692,N_45222);
nor UO_385 (O_385,N_46993,N_48161);
nor UO_386 (O_386,N_49934,N_48471);
nor UO_387 (O_387,N_46971,N_48196);
or UO_388 (O_388,N_48782,N_49074);
nand UO_389 (O_389,N_46221,N_47485);
xor UO_390 (O_390,N_46599,N_47953);
and UO_391 (O_391,N_49021,N_49605);
nand UO_392 (O_392,N_48701,N_45475);
nand UO_393 (O_393,N_45722,N_48673);
nor UO_394 (O_394,N_48343,N_48274);
nand UO_395 (O_395,N_45477,N_47181);
nor UO_396 (O_396,N_47607,N_47443);
xnor UO_397 (O_397,N_47551,N_46935);
or UO_398 (O_398,N_46631,N_46321);
and UO_399 (O_399,N_49214,N_46363);
nor UO_400 (O_400,N_47310,N_46197);
xor UO_401 (O_401,N_46707,N_49365);
xnor UO_402 (O_402,N_49672,N_48688);
nor UO_403 (O_403,N_47425,N_46826);
nand UO_404 (O_404,N_49035,N_48185);
or UO_405 (O_405,N_48604,N_47728);
and UO_406 (O_406,N_45491,N_45229);
and UO_407 (O_407,N_49220,N_45549);
xor UO_408 (O_408,N_47098,N_45499);
nor UO_409 (O_409,N_45297,N_46410);
nand UO_410 (O_410,N_45687,N_46549);
or UO_411 (O_411,N_49636,N_47902);
xor UO_412 (O_412,N_48102,N_47895);
or UO_413 (O_413,N_46145,N_47138);
nor UO_414 (O_414,N_46996,N_46856);
nor UO_415 (O_415,N_45152,N_45758);
or UO_416 (O_416,N_45750,N_49960);
xor UO_417 (O_417,N_46003,N_49260);
or UO_418 (O_418,N_49723,N_45050);
xnor UO_419 (O_419,N_47302,N_47830);
nand UO_420 (O_420,N_46398,N_47210);
xor UO_421 (O_421,N_49231,N_45453);
nand UO_422 (O_422,N_47046,N_45508);
nand UO_423 (O_423,N_46096,N_48842);
and UO_424 (O_424,N_45286,N_49597);
nor UO_425 (O_425,N_45230,N_48459);
xor UO_426 (O_426,N_45328,N_46181);
or UO_427 (O_427,N_47634,N_49647);
xnor UO_428 (O_428,N_49502,N_46941);
and UO_429 (O_429,N_48498,N_47596);
nor UO_430 (O_430,N_46048,N_49737);
and UO_431 (O_431,N_49541,N_49733);
or UO_432 (O_432,N_48569,N_49547);
nor UO_433 (O_433,N_49860,N_48075);
or UO_434 (O_434,N_45579,N_47266);
and UO_435 (O_435,N_45907,N_45957);
and UO_436 (O_436,N_48356,N_46752);
nor UO_437 (O_437,N_47533,N_47103);
and UO_438 (O_438,N_46936,N_49699);
and UO_439 (O_439,N_45134,N_45486);
xor UO_440 (O_440,N_45928,N_46126);
or UO_441 (O_441,N_49518,N_46964);
nor UO_442 (O_442,N_49900,N_47043);
and UO_443 (O_443,N_47053,N_45127);
nand UO_444 (O_444,N_46021,N_48733);
nand UO_445 (O_445,N_45101,N_49505);
and UO_446 (O_446,N_47117,N_46873);
nand UO_447 (O_447,N_47648,N_49394);
and UO_448 (O_448,N_46039,N_48209);
or UO_449 (O_449,N_46274,N_45919);
xnor UO_450 (O_450,N_45876,N_49230);
nand UO_451 (O_451,N_47317,N_49509);
nand UO_452 (O_452,N_49366,N_47013);
nor UO_453 (O_453,N_47814,N_46713);
xnor UO_454 (O_454,N_45241,N_45277);
and UO_455 (O_455,N_45966,N_47142);
and UO_456 (O_456,N_48443,N_47993);
xor UO_457 (O_457,N_45253,N_48401);
nand UO_458 (O_458,N_47174,N_45837);
xor UO_459 (O_459,N_48361,N_47281);
or UO_460 (O_460,N_45846,N_45983);
nand UO_461 (O_461,N_46629,N_49398);
and UO_462 (O_462,N_47282,N_47918);
or UO_463 (O_463,N_46868,N_46404);
xor UO_464 (O_464,N_49309,N_47694);
nand UO_465 (O_465,N_48454,N_48259);
or UO_466 (O_466,N_45849,N_47932);
and UO_467 (O_467,N_47659,N_48005);
and UO_468 (O_468,N_45770,N_49919);
nand UO_469 (O_469,N_47491,N_46372);
xor UO_470 (O_470,N_48366,N_47125);
nor UO_471 (O_471,N_47555,N_47640);
or UO_472 (O_472,N_47440,N_46165);
xor UO_473 (O_473,N_48633,N_45079);
xor UO_474 (O_474,N_48695,N_45025);
nand UO_475 (O_475,N_46802,N_48585);
xnor UO_476 (O_476,N_47359,N_47528);
nor UO_477 (O_477,N_49908,N_48771);
xor UO_478 (O_478,N_48402,N_49283);
and UO_479 (O_479,N_49447,N_46493);
xor UO_480 (O_480,N_47358,N_46773);
and UO_481 (O_481,N_46373,N_48964);
nand UO_482 (O_482,N_49307,N_49897);
nand UO_483 (O_483,N_47526,N_47248);
or UO_484 (O_484,N_45220,N_48649);
xor UO_485 (O_485,N_48592,N_49332);
or UO_486 (O_486,N_47087,N_45700);
nand UO_487 (O_487,N_45408,N_46085);
xnor UO_488 (O_488,N_48834,N_49972);
xor UO_489 (O_489,N_45172,N_45657);
and UO_490 (O_490,N_46673,N_49789);
or UO_491 (O_491,N_46917,N_46331);
nor UO_492 (O_492,N_46451,N_46233);
or UO_493 (O_493,N_45584,N_48021);
nor UO_494 (O_494,N_46056,N_48877);
or UO_495 (O_495,N_48573,N_47265);
or UO_496 (O_496,N_47293,N_48551);
nor UO_497 (O_497,N_47500,N_47263);
and UO_498 (O_498,N_47131,N_49715);
and UO_499 (O_499,N_48195,N_47333);
nor UO_500 (O_500,N_49358,N_49143);
xor UO_501 (O_501,N_47995,N_45143);
nand UO_502 (O_502,N_47072,N_47000);
or UO_503 (O_503,N_48469,N_46424);
or UO_504 (O_504,N_48584,N_47329);
xor UO_505 (O_505,N_48252,N_48074);
and UO_506 (O_506,N_45922,N_45639);
and UO_507 (O_507,N_49807,N_48767);
and UO_508 (O_508,N_47710,N_46129);
xor UO_509 (O_509,N_46324,N_46377);
and UO_510 (O_510,N_46960,N_46108);
nor UO_511 (O_511,N_49427,N_47968);
xor UO_512 (O_512,N_46335,N_49746);
nor UO_513 (O_513,N_47951,N_45685);
nor UO_514 (O_514,N_47798,N_49156);
or UO_515 (O_515,N_46320,N_46303);
and UO_516 (O_516,N_49470,N_47465);
and UO_517 (O_517,N_46926,N_48235);
and UO_518 (O_518,N_45033,N_47852);
and UO_519 (O_519,N_45931,N_48844);
nor UO_520 (O_520,N_45439,N_49958);
nand UO_521 (O_521,N_48833,N_47873);
nand UO_522 (O_522,N_49414,N_48918);
nand UO_523 (O_523,N_47258,N_48043);
xor UO_524 (O_524,N_47209,N_49514);
nand UO_525 (O_525,N_45116,N_48203);
or UO_526 (O_526,N_46161,N_49381);
or UO_527 (O_527,N_49724,N_47867);
nand UO_528 (O_528,N_45965,N_49656);
xor UO_529 (O_529,N_49630,N_46977);
nor UO_530 (O_530,N_45626,N_45741);
and UO_531 (O_531,N_49040,N_45059);
xnor UO_532 (O_532,N_46737,N_45387);
nor UO_533 (O_533,N_45403,N_47474);
and UO_534 (O_534,N_49451,N_48758);
nand UO_535 (O_535,N_49118,N_46249);
or UO_536 (O_536,N_47591,N_45362);
xor UO_537 (O_537,N_48885,N_45535);
and UO_538 (O_538,N_45937,N_45803);
nor UO_539 (O_539,N_47410,N_45162);
nand UO_540 (O_540,N_46422,N_47530);
or UO_541 (O_541,N_49824,N_49729);
and UO_542 (O_542,N_49940,N_48088);
or UO_543 (O_543,N_45029,N_48640);
nor UO_544 (O_544,N_49297,N_45342);
and UO_545 (O_545,N_48904,N_48787);
nor UO_546 (O_546,N_48192,N_49534);
and UO_547 (O_547,N_49382,N_46915);
and UO_548 (O_548,N_49730,N_49421);
xnor UO_549 (O_549,N_47420,N_45924);
nor UO_550 (O_550,N_49742,N_46225);
and UO_551 (O_551,N_45707,N_48666);
nand UO_552 (O_552,N_47758,N_45812);
nor UO_553 (O_553,N_46302,N_49862);
xnor UO_554 (O_554,N_48140,N_49669);
xnor UO_555 (O_555,N_46566,N_47152);
nor UO_556 (O_556,N_45808,N_46771);
and UO_557 (O_557,N_49599,N_48019);
and UO_558 (O_558,N_48117,N_47611);
and UO_559 (O_559,N_46981,N_45105);
or UO_560 (O_560,N_48183,N_45824);
xor UO_561 (O_561,N_47599,N_49924);
xnor UO_562 (O_562,N_49712,N_45232);
or UO_563 (O_563,N_45170,N_45661);
and UO_564 (O_564,N_47136,N_49988);
and UO_565 (O_565,N_48888,N_49520);
nor UO_566 (O_566,N_48827,N_49004);
nand UO_567 (O_567,N_45973,N_47365);
nor UO_568 (O_568,N_47217,N_47532);
and UO_569 (O_569,N_48276,N_45088);
nand UO_570 (O_570,N_46656,N_48762);
and UO_571 (O_571,N_47890,N_47220);
nand UO_572 (O_572,N_45027,N_45529);
or UO_573 (O_573,N_45353,N_47172);
xnor UO_574 (O_574,N_49198,N_47618);
nand UO_575 (O_575,N_46229,N_46061);
nor UO_576 (O_576,N_46539,N_47604);
nor UO_577 (O_577,N_49523,N_46768);
or UO_578 (O_578,N_46973,N_47370);
nor UO_579 (O_579,N_46639,N_46588);
nor UO_580 (O_580,N_49453,N_47559);
nand UO_581 (O_581,N_49100,N_48781);
and UO_582 (O_582,N_45177,N_47567);
nand UO_583 (O_583,N_49843,N_49168);
nand UO_584 (O_584,N_49557,N_45307);
and UO_585 (O_585,N_46254,N_47963);
nor UO_586 (O_586,N_46291,N_47171);
nor UO_587 (O_587,N_46044,N_47973);
nor UO_588 (O_588,N_45208,N_45451);
nor UO_589 (O_589,N_45117,N_45174);
and UO_590 (O_590,N_45295,N_48302);
xnor UO_591 (O_591,N_48938,N_49831);
nand UO_592 (O_592,N_48189,N_46430);
xnor UO_593 (O_593,N_46272,N_45844);
or UO_594 (O_594,N_49663,N_46984);
and UO_595 (O_595,N_49537,N_46607);
xor UO_596 (O_596,N_46876,N_47279);
or UO_597 (O_597,N_47477,N_45274);
and UO_598 (O_598,N_46420,N_46403);
nand UO_599 (O_599,N_48859,N_47754);
nand UO_600 (O_600,N_47770,N_49136);
nor UO_601 (O_601,N_47866,N_48548);
or UO_602 (O_602,N_47502,N_45159);
nand UO_603 (O_603,N_48473,N_46837);
or UO_604 (O_604,N_49489,N_48487);
or UO_605 (O_605,N_48946,N_48094);
nand UO_606 (O_606,N_49274,N_45784);
nand UO_607 (O_607,N_45578,N_45407);
xnor UO_608 (O_608,N_45975,N_46632);
or UO_609 (O_609,N_46111,N_48753);
nor UO_610 (O_610,N_48435,N_48262);
and UO_611 (O_611,N_48403,N_46584);
xnor UO_612 (O_612,N_46281,N_48951);
nand UO_613 (O_613,N_45209,N_46237);
nand UO_614 (O_614,N_45598,N_47987);
xnor UO_615 (O_615,N_45471,N_45345);
or UO_616 (O_616,N_48328,N_46234);
nand UO_617 (O_617,N_48275,N_48817);
xor UO_618 (O_618,N_48679,N_45911);
or UO_619 (O_619,N_45596,N_47433);
xnor UO_620 (O_620,N_47400,N_48407);
or UO_621 (O_621,N_45591,N_48850);
nor UO_622 (O_622,N_45319,N_48352);
and UO_623 (O_623,N_45718,N_48545);
nor UO_624 (O_624,N_47580,N_45343);
nand UO_625 (O_625,N_47861,N_46982);
nor UO_626 (O_626,N_47930,N_47264);
or UO_627 (O_627,N_46081,N_47669);
nor UO_628 (O_628,N_48427,N_45233);
and UO_629 (O_629,N_45468,N_45458);
xor UO_630 (O_630,N_47751,N_47397);
and UO_631 (O_631,N_47330,N_48032);
nand UO_632 (O_632,N_47285,N_47929);
nor UO_633 (O_633,N_47106,N_48325);
xor UO_634 (O_634,N_48194,N_47747);
or UO_635 (O_635,N_45774,N_45284);
nor UO_636 (O_636,N_47899,N_48617);
xor UO_637 (O_637,N_47269,N_47739);
nor UO_638 (O_638,N_46072,N_47822);
xnor UO_639 (O_639,N_47829,N_49969);
nor UO_640 (O_640,N_46681,N_49905);
nor UO_641 (O_641,N_48574,N_45847);
nand UO_642 (O_642,N_48974,N_46440);
or UO_643 (O_643,N_47862,N_45089);
xor UO_644 (O_644,N_46544,N_47026);
and UO_645 (O_645,N_49475,N_46757);
nand UO_646 (O_646,N_48026,N_48567);
nand UO_647 (O_647,N_48227,N_49782);
nand UO_648 (O_648,N_49226,N_49968);
nor UO_649 (O_649,N_47911,N_45076);
or UO_650 (O_650,N_47876,N_48405);
nor UO_651 (O_651,N_47839,N_45607);
or UO_652 (O_652,N_47156,N_46393);
nor UO_653 (O_653,N_47722,N_48897);
or UO_654 (O_654,N_49735,N_49437);
xor UO_655 (O_655,N_46253,N_45921);
or UO_656 (O_656,N_49888,N_46685);
nor UO_657 (O_657,N_49703,N_47429);
or UO_658 (O_658,N_49243,N_46923);
nor UO_659 (O_659,N_48416,N_47154);
nand UO_660 (O_660,N_49861,N_48643);
xnor UO_661 (O_661,N_48702,N_47800);
or UO_662 (O_662,N_47912,N_47863);
and UO_663 (O_663,N_47301,N_49229);
and UO_664 (O_664,N_47743,N_49176);
xnor UO_665 (O_665,N_46835,N_45381);
nand UO_666 (O_666,N_46279,N_47299);
and UO_667 (O_667,N_49490,N_48243);
and UO_668 (O_668,N_48426,N_46686);
nor UO_669 (O_669,N_47539,N_46488);
or UO_670 (O_670,N_45873,N_45990);
and UO_671 (O_671,N_46419,N_47869);
xnor UO_672 (O_672,N_47952,N_49241);
nand UO_673 (O_673,N_49877,N_49345);
or UO_674 (O_674,N_46243,N_46569);
nor UO_675 (O_675,N_49460,N_48909);
or UO_676 (O_676,N_47133,N_46741);
and UO_677 (O_677,N_48731,N_47892);
nor UO_678 (O_678,N_45107,N_49786);
nand UO_679 (O_679,N_47149,N_48950);
nor UO_680 (O_680,N_46214,N_47954);
xnor UO_681 (O_681,N_46339,N_49023);
nand UO_682 (O_682,N_49999,N_45738);
nor UO_683 (O_683,N_47782,N_45100);
nand UO_684 (O_684,N_48544,N_46779);
nor UO_685 (O_685,N_45939,N_45348);
and UO_686 (O_686,N_48712,N_48409);
xnor UO_687 (O_687,N_45506,N_46803);
or UO_688 (O_688,N_45616,N_46814);
nor UO_689 (O_689,N_48451,N_47601);
xor UO_690 (O_690,N_46338,N_49610);
xnor UO_691 (O_691,N_46415,N_45802);
and UO_692 (O_692,N_46104,N_49341);
nor UO_693 (O_693,N_49215,N_48146);
nor UO_694 (O_694,N_48149,N_47510);
or UO_695 (O_695,N_48463,N_45668);
and UO_696 (O_696,N_47200,N_48351);
nand UO_697 (O_697,N_49020,N_45330);
and UO_698 (O_698,N_45615,N_49743);
and UO_699 (O_699,N_48453,N_48141);
nor UO_700 (O_700,N_45565,N_46959);
nor UO_701 (O_701,N_46110,N_45336);
and UO_702 (O_702,N_46127,N_45223);
xnor UO_703 (O_703,N_48532,N_45394);
nand UO_704 (O_704,N_47494,N_45842);
nor UO_705 (O_705,N_49441,N_45494);
and UO_706 (O_706,N_49957,N_49920);
nor UO_707 (O_707,N_48441,N_47088);
and UO_708 (O_708,N_46327,N_45400);
nand UO_709 (O_709,N_45751,N_46041);
xnor UO_710 (O_710,N_45648,N_45935);
nand UO_711 (O_711,N_45332,N_48706);
and UO_712 (O_712,N_46450,N_46118);
nor UO_713 (O_713,N_48754,N_47378);
xnor UO_714 (O_714,N_46574,N_49607);
or UO_715 (O_715,N_45505,N_46099);
and UO_716 (O_716,N_47034,N_45594);
nand UO_717 (O_717,N_46602,N_45329);
nand UO_718 (O_718,N_45454,N_47906);
nand UO_719 (O_719,N_47629,N_46800);
nor UO_720 (O_720,N_47955,N_45762);
nand UO_721 (O_721,N_49640,N_45268);
nor UO_722 (O_722,N_49562,N_48811);
or UO_723 (O_723,N_47720,N_46346);
xnor UO_724 (O_724,N_48123,N_45513);
and UO_725 (O_725,N_49619,N_49581);
and UO_726 (O_726,N_49629,N_48414);
nor UO_727 (O_727,N_49426,N_48512);
xnor UO_728 (O_728,N_47435,N_48034);
xor UO_729 (O_729,N_46563,N_48519);
nand UO_730 (O_730,N_45860,N_45952);
and UO_731 (O_731,N_49104,N_48272);
nor UO_732 (O_732,N_47670,N_49189);
nor UO_733 (O_733,N_49522,N_48713);
xnor UO_734 (O_734,N_46437,N_45947);
xnor UO_735 (O_735,N_45126,N_46674);
xnor UO_736 (O_736,N_45202,N_48870);
xnor UO_737 (O_737,N_46693,N_49895);
and UO_738 (O_738,N_46777,N_48508);
nand UO_739 (O_739,N_46896,N_46494);
xor UO_740 (O_740,N_47186,N_49674);
xnor UO_741 (O_741,N_48119,N_46581);
nor UO_742 (O_742,N_45406,N_46027);
or UO_743 (O_743,N_47649,N_47346);
and UO_744 (O_744,N_45500,N_49906);
nor UO_745 (O_745,N_46943,N_47340);
xor UO_746 (O_746,N_48841,N_49054);
nand UO_747 (O_747,N_47480,N_47727);
xnor UO_748 (O_748,N_47042,N_45125);
or UO_749 (O_749,N_45554,N_48260);
nor UO_750 (O_750,N_47094,N_48038);
xnor UO_751 (O_751,N_45914,N_46698);
or UO_752 (O_752,N_45495,N_45623);
and UO_753 (O_753,N_45150,N_46930);
and UO_754 (O_754,N_46013,N_46252);
or UO_755 (O_755,N_46551,N_45682);
or UO_756 (O_756,N_46655,N_47765);
nand UO_757 (O_757,N_48248,N_48010);
nand UO_758 (O_758,N_46492,N_49342);
xnor UO_759 (O_759,N_47385,N_48928);
and UO_760 (O_760,N_45364,N_45043);
nand UO_761 (O_761,N_45144,N_49551);
or UO_762 (O_762,N_46107,N_45291);
or UO_763 (O_763,N_47511,N_47052);
nand UO_764 (O_764,N_45352,N_47167);
and UO_765 (O_765,N_49706,N_46326);
nor UO_766 (O_766,N_47921,N_47617);
and UO_767 (O_767,N_45369,N_45936);
xor UO_768 (O_768,N_48738,N_46063);
xnor UO_769 (O_769,N_46278,N_47453);
nand UO_770 (O_770,N_47496,N_46723);
and UO_771 (O_771,N_45109,N_45833);
or UO_772 (O_772,N_49668,N_47122);
nor UO_773 (O_773,N_49469,N_46370);
nor UO_774 (O_774,N_46382,N_47382);
or UO_775 (O_775,N_49904,N_45595);
or UO_776 (O_776,N_49657,N_48991);
and UO_777 (O_777,N_48602,N_46675);
nor UO_778 (O_778,N_47236,N_49316);
nand UO_779 (O_779,N_48327,N_48214);
nor UO_780 (O_780,N_49103,N_45052);
nand UO_781 (O_781,N_48802,N_49770);
and UO_782 (O_782,N_49582,N_48428);
xnor UO_783 (O_783,N_46465,N_48225);
xnor UO_784 (O_784,N_47314,N_48294);
and UO_785 (O_785,N_48903,N_49956);
nor UO_786 (O_786,N_48434,N_49380);
nand UO_787 (O_787,N_48036,N_48130);
nand UO_788 (O_788,N_47615,N_46267);
or UO_789 (O_789,N_45334,N_45756);
xnor UO_790 (O_790,N_45178,N_48232);
and UO_791 (O_791,N_45875,N_47123);
nand UO_792 (O_792,N_46392,N_46426);
nor UO_793 (O_793,N_46351,N_47128);
nor UO_794 (O_794,N_45372,N_47926);
nand UO_795 (O_795,N_48160,N_48367);
nand UO_796 (O_796,N_45257,N_46205);
nor UO_797 (O_797,N_49171,N_49688);
xor UO_798 (O_798,N_45891,N_47884);
nor UO_799 (O_799,N_48775,N_49084);
and UO_800 (O_800,N_45219,N_49925);
nor UO_801 (O_801,N_47900,N_48886);
nor UO_802 (O_802,N_49450,N_49211);
nand UO_803 (O_803,N_45768,N_49119);
nand UO_804 (O_804,N_47762,N_46586);
or UO_805 (O_805,N_46471,N_48916);
xor UO_806 (O_806,N_48389,N_49207);
and UO_807 (O_807,N_49650,N_46336);
nor UO_808 (O_808,N_48867,N_46687);
and UO_809 (O_809,N_48475,N_48491);
xnor UO_810 (O_810,N_47177,N_48902);
nor UO_811 (O_811,N_45771,N_49869);
nor UO_812 (O_812,N_47905,N_45603);
nor UO_813 (O_813,N_46764,N_47071);
nor UO_814 (O_814,N_46523,N_47215);
or UO_815 (O_815,N_45961,N_48807);
or UO_816 (O_816,N_45445,N_46231);
nand UO_817 (O_817,N_45577,N_45544);
or UO_818 (O_818,N_49191,N_49780);
and UO_819 (O_819,N_45686,N_45733);
or UO_820 (O_820,N_47473,N_48760);
nand UO_821 (O_821,N_47342,N_45656);
xnor UO_822 (O_822,N_49878,N_49268);
or UO_823 (O_823,N_47837,N_47432);
nand UO_824 (O_824,N_45316,N_45155);
nor UO_825 (O_825,N_47923,N_49714);
and UO_826 (O_826,N_48077,N_47702);
nor UO_827 (O_827,N_47836,N_49094);
xor UO_828 (O_828,N_48070,N_46654);
nor UO_829 (O_829,N_49010,N_46985);
and UO_830 (O_830,N_47356,N_46822);
xnor UO_831 (O_831,N_45299,N_49625);
or UO_832 (O_832,N_47045,N_47457);
nand UO_833 (O_833,N_49530,N_46193);
xor UO_834 (O_834,N_46649,N_47853);
nand UO_835 (O_835,N_45021,N_48156);
and UO_836 (O_836,N_46642,N_45376);
or UO_837 (O_837,N_46762,N_45769);
nor UO_838 (O_838,N_47380,N_46872);
nor UO_839 (O_839,N_47655,N_47778);
nand UO_840 (O_840,N_47713,N_49933);
and UO_841 (O_841,N_47531,N_45550);
nand UO_842 (O_842,N_47840,N_46276);
nor UO_843 (O_843,N_48557,N_49448);
and UO_844 (O_844,N_47663,N_48101);
xnor UO_845 (O_845,N_46646,N_48535);
and UO_846 (O_846,N_49587,N_45294);
or UO_847 (O_847,N_49527,N_48591);
or UO_848 (O_848,N_48107,N_46055);
or UO_849 (O_849,N_45430,N_46195);
nand UO_850 (O_850,N_49602,N_47939);
or UO_851 (O_851,N_46332,N_45462);
nor UO_852 (O_852,N_45515,N_45068);
nor UO_853 (O_853,N_48878,N_48377);
nand UO_854 (O_854,N_45087,N_48699);
or UO_855 (O_855,N_47077,N_47821);
nand UO_856 (O_856,N_45564,N_49529);
and UO_857 (O_857,N_47687,N_48424);
nor UO_858 (O_858,N_46433,N_45995);
nor UO_859 (O_859,N_45318,N_47748);
or UO_860 (O_860,N_49683,N_47159);
nor UO_861 (O_861,N_48956,N_46615);
and UO_862 (O_862,N_47124,N_48601);
xnor UO_863 (O_863,N_47223,N_46057);
or UO_864 (O_864,N_47996,N_46898);
and UO_865 (O_865,N_49393,N_49749);
xor UO_866 (O_866,N_46667,N_46357);
and UO_867 (O_867,N_48957,N_48464);
or UO_868 (O_868,N_49127,N_47893);
nand UO_869 (O_869,N_49014,N_48282);
nor UO_870 (O_870,N_47176,N_45958);
and UO_871 (O_871,N_48206,N_46167);
nor UO_872 (O_872,N_47783,N_48506);
or UO_873 (O_873,N_49468,N_47886);
xnor UO_874 (O_874,N_48210,N_47516);
nor UO_875 (O_875,N_47003,N_48745);
nand UO_876 (O_876,N_48485,N_45748);
and UO_877 (O_877,N_45227,N_46944);
nor UO_878 (O_878,N_45624,N_49898);
nand UO_879 (O_879,N_45872,N_46869);
xor UO_880 (O_880,N_48198,N_46730);
and UO_881 (O_881,N_46785,N_45338);
nor UO_882 (O_882,N_45235,N_48605);
or UO_883 (O_883,N_45238,N_47865);
and UO_884 (O_884,N_48069,N_48676);
nand UO_885 (O_885,N_46308,N_49327);
xor UO_886 (O_886,N_48735,N_49708);
xor UO_887 (O_887,N_46724,N_46788);
or UO_888 (O_888,N_46371,N_48801);
and UO_889 (O_889,N_48795,N_47376);
or UO_890 (O_890,N_49495,N_49855);
and UO_891 (O_891,N_49029,N_46997);
nor UO_892 (O_892,N_48511,N_46628);
xor UO_893 (O_893,N_49109,N_48324);
and UO_894 (O_894,N_45449,N_46296);
xnor UO_895 (O_895,N_45517,N_48819);
xor UO_896 (O_896,N_49131,N_48143);
nand UO_897 (O_897,N_48492,N_48989);
or UO_898 (O_898,N_48992,N_49091);
nor UO_899 (O_899,N_45419,N_45404);
xnor UO_900 (O_900,N_47827,N_45831);
nor UO_901 (O_901,N_46867,N_48559);
nand UO_902 (O_902,N_49296,N_48201);
xnor UO_903 (O_903,N_48114,N_47916);
nor UO_904 (O_904,N_47490,N_49653);
and UO_905 (O_905,N_47941,N_49881);
nand UO_906 (O_906,N_48423,N_46000);
and UO_907 (O_907,N_45840,N_49335);
xnor UO_908 (O_908,N_47155,N_48147);
xor UO_909 (O_909,N_46650,N_45056);
or UO_910 (O_910,N_45962,N_49838);
xor UO_911 (O_911,N_49415,N_49813);
or UO_912 (O_912,N_48607,N_48756);
and UO_913 (O_913,N_45099,N_47462);
and UO_914 (O_914,N_46421,N_46360);
nand UO_915 (O_915,N_48931,N_46946);
xnor UO_916 (O_916,N_48483,N_49627);
nand UO_917 (O_917,N_49785,N_49455);
and UO_918 (O_918,N_48575,N_47109);
nand UO_919 (O_919,N_45146,N_47005);
and UO_920 (O_920,N_46808,N_49034);
xor UO_921 (O_921,N_48929,N_48489);
and UO_922 (O_922,N_48045,N_46819);
and UO_923 (O_923,N_45289,N_45625);
and UO_924 (O_924,N_49397,N_45642);
xor UO_925 (O_925,N_47002,N_49915);
nor UO_926 (O_926,N_47729,N_46924);
nand UO_927 (O_927,N_47288,N_49138);
xor UO_928 (O_928,N_48207,N_46435);
xnor UO_929 (O_929,N_46543,N_46025);
nand UO_930 (O_930,N_45482,N_46236);
or UO_931 (O_931,N_48313,N_46672);
and UO_932 (O_932,N_46045,N_45461);
nand UO_933 (O_933,N_45545,N_46079);
nor UO_934 (O_934,N_49612,N_45270);
or UO_935 (O_935,N_46239,N_49444);
and UO_936 (O_936,N_49006,N_48176);
and UO_937 (O_937,N_47733,N_46853);
nand UO_938 (O_938,N_45669,N_48249);
and UO_939 (O_939,N_45628,N_48962);
and UO_940 (O_940,N_45168,N_49086);
xor UO_941 (O_941,N_45028,N_48749);
and UO_942 (O_942,N_47578,N_47621);
xor UO_943 (O_943,N_47060,N_45045);
nor UO_944 (O_944,N_49833,N_47619);
or UO_945 (O_945,N_47773,N_46929);
nand UO_946 (O_946,N_46579,N_46018);
and UO_947 (O_947,N_46962,N_49019);
xnor UO_948 (O_948,N_46913,N_48211);
and UO_949 (O_949,N_45767,N_47976);
or UO_950 (O_950,N_45064,N_49548);
and UO_951 (O_951,N_48387,N_48611);
or UO_952 (O_952,N_49978,N_49484);
or UO_953 (O_953,N_46173,N_45466);
nor UO_954 (O_954,N_45039,N_45314);
nor UO_955 (O_955,N_49488,N_49528);
xor UO_956 (O_956,N_45874,N_46879);
xnor UO_957 (O_957,N_45698,N_48406);
nor UO_958 (O_958,N_46909,N_45815);
nand UO_959 (O_959,N_48595,N_46159);
or UO_960 (O_960,N_45005,N_45699);
and UO_961 (O_961,N_46524,N_49944);
nand UO_962 (O_962,N_49419,N_45395);
and UO_963 (O_963,N_49330,N_47838);
xor UO_964 (O_964,N_47651,N_47105);
and UO_965 (O_965,N_49821,N_49806);
nor UO_966 (O_966,N_49512,N_46804);
and UO_967 (O_967,N_48949,N_45953);
nor UO_968 (O_968,N_46521,N_47126);
and UO_969 (O_969,N_46199,N_46374);
or UO_970 (O_970,N_45653,N_47864);
nand UO_971 (O_971,N_49464,N_49921);
or UO_972 (O_972,N_48488,N_45672);
nand UO_973 (O_973,N_48538,N_46390);
or UO_974 (O_974,N_47183,N_48497);
xnor UO_975 (O_975,N_45775,N_46644);
nor UO_976 (O_976,N_48908,N_48727);
nand UO_977 (O_977,N_48167,N_46284);
and UO_978 (O_978,N_47100,N_47395);
nand UO_979 (O_979,N_48152,N_49777);
xnor UO_980 (O_980,N_48042,N_47947);
nor UO_981 (O_981,N_48622,N_45627);
nor UO_982 (O_982,N_46515,N_48099);
nand UO_983 (O_983,N_45765,N_49964);
xor UO_984 (O_984,N_48927,N_45501);
or UO_985 (O_985,N_47335,N_48961);
and UO_986 (O_986,N_46269,N_49781);
and UO_987 (O_987,N_45104,N_47820);
xnor UO_988 (O_988,N_45787,N_47016);
and UO_989 (O_989,N_46743,N_47600);
nand UO_990 (O_990,N_45267,N_46530);
nor UO_991 (O_991,N_48180,N_49726);
nand UO_992 (O_992,N_49590,N_46062);
or UO_993 (O_993,N_47482,N_49641);
xor UO_994 (O_994,N_49135,N_47349);
or UO_995 (O_995,N_49546,N_45641);
or UO_996 (O_996,N_47726,N_47712);
or UO_997 (O_997,N_48231,N_47914);
xor UO_998 (O_998,N_48285,N_46058);
xnor UO_999 (O_999,N_46520,N_48969);
nand UO_1000 (O_1000,N_49727,N_47116);
or UO_1001 (O_1001,N_45212,N_49910);
nand UO_1002 (O_1002,N_46400,N_49032);
nand UO_1003 (O_1003,N_49811,N_47842);
xor UO_1004 (O_1004,N_47062,N_45574);
or UO_1005 (O_1005,N_47964,N_48884);
and UO_1006 (O_1006,N_47538,N_49432);
nand UO_1007 (O_1007,N_45537,N_47985);
xor UO_1008 (O_1008,N_46558,N_49251);
and UO_1009 (O_1009,N_48472,N_46829);
nand UO_1010 (O_1010,N_49791,N_45391);
or UO_1011 (O_1011,N_45798,N_46796);
nor UO_1012 (O_1012,N_49815,N_48397);
nand UO_1013 (O_1013,N_46183,N_49456);
or UO_1014 (O_1014,N_47323,N_48664);
and UO_1015 (O_1015,N_47507,N_48540);
nand UO_1016 (O_1016,N_47121,N_49442);
nand UO_1017 (O_1017,N_48516,N_49661);
nor UO_1018 (O_1018,N_49513,N_46556);
nor UO_1019 (O_1019,N_46076,N_49963);
nand UO_1020 (O_1020,N_47079,N_45304);
nand UO_1021 (O_1021,N_46719,N_45988);
and UO_1022 (O_1022,N_45511,N_49146);
or UO_1023 (O_1023,N_48608,N_49745);
nor UO_1024 (O_1024,N_49477,N_45760);
xnor UO_1025 (O_1025,N_45032,N_48752);
nand UO_1026 (O_1026,N_47868,N_49835);
xnor UO_1027 (O_1027,N_47872,N_48565);
nor UO_1028 (O_1028,N_49264,N_45715);
nand UO_1029 (O_1029,N_45925,N_49465);
or UO_1030 (O_1030,N_48665,N_47497);
nand UO_1031 (O_1031,N_46137,N_46292);
and UO_1032 (O_1032,N_46347,N_45030);
xor UO_1033 (O_1033,N_45322,N_48447);
or UO_1034 (O_1034,N_46144,N_48896);
nand UO_1035 (O_1035,N_47622,N_49604);
and UO_1036 (O_1036,N_45035,N_45923);
or UO_1037 (O_1037,N_49613,N_45169);
and UO_1038 (O_1038,N_49805,N_47306);
or UO_1039 (O_1039,N_46189,N_45240);
and UO_1040 (O_1040,N_49333,N_45853);
xnor UO_1041 (O_1041,N_45806,N_48714);
and UO_1042 (O_1042,N_48452,N_47846);
or UO_1043 (O_1043,N_47788,N_48431);
nand UO_1044 (O_1044,N_46484,N_47055);
xor UO_1045 (O_1045,N_48215,N_45048);
xor UO_1046 (O_1046,N_49440,N_45122);
nand UO_1047 (O_1047,N_48996,N_49411);
nand UO_1048 (O_1048,N_49609,N_48293);
xor UO_1049 (O_1049,N_48029,N_49408);
nor UO_1050 (O_1050,N_45999,N_48852);
xor UO_1051 (O_1051,N_45261,N_45930);
nand UO_1052 (O_1052,N_49279,N_47684);
xnor UO_1053 (O_1053,N_46816,N_48718);
xor UO_1054 (O_1054,N_46333,N_45702);
nor UO_1055 (O_1055,N_45793,N_45690);
nor UO_1056 (O_1056,N_47345,N_48794);
nor UO_1057 (O_1057,N_45943,N_48442);
nand UO_1058 (O_1058,N_49966,N_49367);
nor UO_1059 (O_1059,N_46448,N_47623);
or UO_1060 (O_1060,N_47672,N_48046);
xnor UO_1061 (O_1061,N_48765,N_46070);
xor UO_1062 (O_1062,N_49755,N_46215);
nand UO_1063 (O_1063,N_47064,N_48517);
nor UO_1064 (O_1064,N_47948,N_48537);
or UO_1065 (O_1065,N_46022,N_46168);
or UO_1066 (O_1066,N_49157,N_45061);
or UO_1067 (O_1067,N_49236,N_49950);
or UO_1068 (O_1068,N_46598,N_48323);
xnor UO_1069 (O_1069,N_47731,N_46527);
or UO_1070 (O_1070,N_47675,N_49564);
nand UO_1071 (O_1071,N_45671,N_48080);
or UO_1072 (O_1072,N_46585,N_48653);
and UO_1073 (O_1073,N_47620,N_48880);
xnor UO_1074 (O_1074,N_47633,N_45066);
nor UO_1075 (O_1075,N_46306,N_48357);
xor UO_1076 (O_1076,N_47166,N_45380);
or UO_1077 (O_1077,N_49566,N_47324);
nor UO_1078 (O_1078,N_46026,N_48558);
xor UO_1079 (O_1079,N_48571,N_48984);
xor UO_1080 (O_1080,N_45022,N_46452);
nand UO_1081 (O_1081,N_47146,N_46445);
or UO_1082 (O_1082,N_47975,N_48915);
xnor UO_1083 (O_1083,N_46084,N_47858);
or UO_1084 (O_1084,N_47988,N_45077);
and UO_1085 (O_1085,N_48737,N_45167);
nor UO_1086 (O_1086,N_49062,N_46264);
or UO_1087 (O_1087,N_48300,N_47755);
xor UO_1088 (O_1088,N_48087,N_48191);
or UO_1089 (O_1089,N_49395,N_45303);
nand UO_1090 (O_1090,N_49234,N_48821);
or UO_1091 (O_1091,N_49093,N_48148);
and UO_1092 (O_1092,N_46532,N_46187);
nand UO_1093 (O_1093,N_49362,N_45129);
or UO_1094 (O_1094,N_45301,N_47978);
xnor UO_1095 (O_1095,N_49826,N_49741);
xor UO_1096 (O_1096,N_45069,N_47576);
and UO_1097 (O_1097,N_49491,N_47799);
and UO_1098 (O_1098,N_49718,N_47847);
nand UO_1099 (O_1099,N_48412,N_48134);
and UO_1100 (O_1100,N_45351,N_48848);
and UO_1101 (O_1101,N_47904,N_49193);
nand UO_1102 (O_1102,N_49425,N_49946);
nor UO_1103 (O_1103,N_49463,N_46130);
or UO_1104 (O_1104,N_48493,N_46049);
and UO_1105 (O_1105,N_46699,N_49277);
xor UO_1106 (O_1106,N_46836,N_45526);
and UO_1107 (O_1107,N_45934,N_46065);
or UO_1108 (O_1108,N_48741,N_49360);
nor UO_1109 (O_1109,N_48120,N_45528);
or UO_1110 (O_1110,N_49583,N_48008);
nand UO_1111 (O_1111,N_47802,N_48154);
or UO_1112 (O_1112,N_46793,N_48168);
xnor UO_1113 (O_1113,N_45173,N_47095);
nor UO_1114 (O_1114,N_47361,N_45254);
and UO_1115 (O_1115,N_47111,N_46648);
and UO_1116 (O_1116,N_48780,N_49975);
nand UO_1117 (O_1117,N_49132,N_47857);
xnor UO_1118 (O_1118,N_46511,N_47426);
or UO_1119 (O_1119,N_46661,N_47004);
nand UO_1120 (O_1120,N_46071,N_45073);
nor UO_1121 (O_1121,N_46151,N_46499);
xnor UO_1122 (O_1122,N_46224,N_46064);
nor UO_1123 (O_1123,N_46042,N_49938);
nand UO_1124 (O_1124,N_49533,N_48507);
xor UO_1125 (O_1125,N_49142,N_47260);
nor UO_1126 (O_1126,N_47992,N_48100);
or UO_1127 (O_1127,N_45397,N_46874);
xor UO_1128 (O_1128,N_45862,N_46759);
and UO_1129 (O_1129,N_49263,N_48413);
and UO_1130 (O_1130,N_47101,N_47448);
and UO_1131 (O_1131,N_46545,N_46207);
xnor UO_1132 (O_1132,N_47945,N_48380);
nand UO_1133 (O_1133,N_49347,N_45799);
xnor UO_1134 (O_1134,N_49543,N_46744);
or UO_1135 (O_1135,N_48111,N_49987);
nand UO_1136 (O_1136,N_48615,N_46043);
nor UO_1137 (O_1137,N_45103,N_48092);
or UO_1138 (O_1138,N_46206,N_47245);
nand UO_1139 (O_1139,N_46136,N_48830);
xnor UO_1140 (O_1140,N_49175,N_48739);
xor UO_1141 (O_1141,N_49485,N_45674);
or UO_1142 (O_1142,N_47389,N_47417);
xnor UO_1143 (O_1143,N_49899,N_48457);
or UO_1144 (O_1144,N_49545,N_46701);
nor UO_1145 (O_1145,N_48645,N_49139);
and UO_1146 (O_1146,N_47965,N_49401);
xnor UO_1147 (O_1147,N_45583,N_46643);
or UO_1148 (O_1148,N_46314,N_48144);
nor UO_1149 (O_1149,N_45730,N_46140);
and UO_1150 (O_1150,N_48698,N_47240);
and UO_1151 (O_1151,N_48250,N_48440);
xnor UO_1152 (O_1152,N_46645,N_45389);
nand UO_1153 (O_1153,N_47645,N_49667);
or UO_1154 (O_1154,N_45386,N_45207);
or UO_1155 (O_1155,N_45568,N_48770);
nand UO_1156 (O_1156,N_45945,N_45866);
nand UO_1157 (O_1157,N_46204,N_49000);
and UO_1158 (O_1158,N_45344,N_49698);
or UO_1159 (O_1159,N_45618,N_46036);
nand UO_1160 (O_1160,N_48139,N_48006);
nor UO_1161 (O_1161,N_45237,N_49945);
nand UO_1162 (O_1162,N_48384,N_49901);
xor UO_1163 (O_1163,N_47196,N_46304);
and UO_1164 (O_1164,N_48465,N_46659);
nor UO_1165 (O_1165,N_47408,N_49539);
nor UO_1166 (O_1166,N_45480,N_47714);
nand UO_1167 (O_1167,N_45176,N_45300);
nand UO_1168 (O_1168,N_45448,N_45279);
nor UO_1169 (O_1169,N_46428,N_46705);
nor UO_1170 (O_1170,N_46638,N_49902);
or UO_1171 (O_1171,N_45489,N_48972);
nor UO_1172 (O_1172,N_48920,N_46368);
nor UO_1173 (O_1173,N_46995,N_45834);
nand UO_1174 (O_1174,N_46244,N_45673);
nor UO_1175 (O_1175,N_46795,N_48097);
and UO_1176 (O_1176,N_49584,N_49459);
xor UO_1177 (O_1177,N_47806,N_45282);
nand UO_1178 (O_1178,N_45650,N_46847);
and UO_1179 (O_1179,N_46931,N_49059);
or UO_1180 (O_1180,N_49265,N_45666);
or UO_1181 (O_1181,N_46622,N_49885);
or UO_1182 (O_1182,N_47801,N_49199);
xor UO_1183 (O_1183,N_47492,N_47704);
nor UO_1184 (O_1184,N_48386,N_48017);
nor UO_1185 (O_1185,N_47212,N_48365);
or UO_1186 (O_1186,N_47565,N_45604);
nand UO_1187 (O_1187,N_45151,N_46389);
nand UO_1188 (O_1188,N_45779,N_49267);
nor UO_1189 (O_1189,N_47458,N_46030);
nand UO_1190 (O_1190,N_49007,N_45084);
nand UO_1191 (O_1191,N_45080,N_47997);
or UO_1192 (O_1192,N_46417,N_45097);
or UO_1193 (O_1193,N_49254,N_48911);
and UO_1194 (O_1194,N_48954,N_45982);
and UO_1195 (O_1195,N_47843,N_49953);
nand UO_1196 (O_1196,N_48740,N_49569);
or UO_1197 (O_1197,N_49907,N_45467);
and UO_1198 (O_1198,N_47194,N_49417);
nor UO_1199 (O_1199,N_45558,N_47804);
or UO_1200 (O_1200,N_47112,N_47396);
or UO_1201 (O_1201,N_47683,N_48729);
and UO_1202 (O_1202,N_46670,N_46367);
nor UO_1203 (O_1203,N_49368,N_47605);
nand UO_1204 (O_1204,N_45729,N_49575);
and UO_1205 (O_1205,N_49278,N_45373);
nand UO_1206 (O_1206,N_49406,N_46260);
xnor UO_1207 (O_1207,N_48632,N_45991);
or UO_1208 (O_1208,N_46548,N_47874);
and UO_1209 (O_1209,N_48330,N_48800);
nand UO_1210 (O_1210,N_46365,N_47145);
xor UO_1211 (O_1211,N_47630,N_47211);
xnor UO_1212 (O_1212,N_46918,N_49200);
xnor UO_1213 (O_1213,N_48166,N_49232);
nor UO_1214 (O_1214,N_48942,N_46679);
nor UO_1215 (O_1215,N_48177,N_46858);
nor UO_1216 (O_1216,N_49325,N_47808);
or UO_1217 (O_1217,N_46497,N_49312);
xor UO_1218 (O_1218,N_49056,N_47547);
nand UO_1219 (O_1219,N_48341,N_47047);
nor UO_1220 (O_1220,N_49413,N_47373);
and UO_1221 (O_1221,N_47466,N_46769);
or UO_1222 (O_1222,N_49874,N_49622);
nand UO_1223 (O_1223,N_46565,N_45970);
or UO_1224 (O_1224,N_46512,N_45384);
or UO_1225 (O_1225,N_49977,N_46692);
or UO_1226 (O_1226,N_47575,N_48321);
nor UO_1227 (O_1227,N_45444,N_48359);
and UO_1228 (O_1228,N_46573,N_49117);
or UO_1229 (O_1229,N_49246,N_49320);
or UO_1230 (O_1230,N_47326,N_45179);
or UO_1231 (O_1231,N_48131,N_47431);
or UO_1232 (O_1232,N_45509,N_49081);
xor UO_1233 (O_1233,N_45838,N_46812);
nor UO_1234 (O_1234,N_48554,N_47148);
nand UO_1235 (O_1235,N_49511,N_48480);
and UO_1236 (O_1236,N_47207,N_46232);
or UO_1237 (O_1237,N_46555,N_46890);
or UO_1238 (O_1238,N_47920,N_45040);
and UO_1239 (O_1239,N_49428,N_48373);
and UO_1240 (O_1240,N_48082,N_48496);
nand UO_1241 (O_1241,N_48062,N_45753);
or UO_1242 (O_1242,N_46040,N_48641);
or UO_1243 (O_1243,N_48020,N_45612);
and UO_1244 (O_1244,N_46075,N_47897);
nor UO_1245 (O_1245,N_46082,N_45597);
nor UO_1246 (O_1246,N_47708,N_49697);
nand UO_1247 (O_1247,N_45496,N_47337);
or UO_1248 (O_1248,N_46746,N_46916);
xnor UO_1249 (O_1249,N_46240,N_46343);
nand UO_1250 (O_1250,N_48221,N_47742);
xor UO_1251 (O_1251,N_47118,N_49820);
nand UO_1252 (O_1252,N_45142,N_45555);
and UO_1253 (O_1253,N_49552,N_46580);
nand UO_1254 (O_1254,N_48022,N_45306);
and UO_1255 (O_1255,N_47089,N_49646);
or UO_1256 (O_1256,N_45514,N_48450);
and UO_1257 (O_1257,N_45566,N_46091);
or UO_1258 (O_1258,N_47478,N_45667);
nand UO_1259 (O_1259,N_47479,N_45326);
and UO_1260 (O_1260,N_48169,N_45331);
nand UO_1261 (O_1261,N_46460,N_47012);
nand UO_1262 (O_1262,N_45721,N_47129);
nand UO_1263 (O_1263,N_47353,N_46008);
xor UO_1264 (O_1264,N_48722,N_49256);
xnor UO_1265 (O_1265,N_45354,N_49803);
xnor UO_1266 (O_1266,N_46436,N_49594);
nor UO_1267 (O_1267,N_47505,N_48481);
nor UO_1268 (O_1268,N_48590,N_48683);
or UO_1269 (O_1269,N_45556,N_48288);
and UO_1270 (O_1270,N_48858,N_45510);
nor UO_1271 (O_1271,N_47579,N_47044);
nand UO_1272 (O_1272,N_45133,N_45415);
nand UO_1273 (O_1273,N_47553,N_47989);
xor UO_1274 (O_1274,N_49385,N_49645);
xor UO_1275 (O_1275,N_45018,N_48118);
nand UO_1276 (O_1276,N_45814,N_45180);
nor UO_1277 (O_1277,N_45740,N_48432);
nand UO_1278 (O_1278,N_45199,N_47891);
or UO_1279 (O_1279,N_48420,N_47570);
nor UO_1280 (O_1280,N_45382,N_47833);
xor UO_1281 (O_1281,N_49391,N_45092);
nand UO_1282 (O_1282,N_45716,N_45365);
xnor UO_1283 (O_1283,N_48116,N_48503);
nand UO_1284 (O_1284,N_47626,N_46282);
and UO_1285 (O_1285,N_48068,N_49995);
nand UO_1286 (O_1286,N_47498,N_46832);
nand UO_1287 (O_1287,N_49659,N_45948);
or UO_1288 (O_1288,N_48925,N_48164);
nand UO_1289 (O_1289,N_48894,N_48932);
or UO_1290 (O_1290,N_49105,N_47514);
nor UO_1291 (O_1291,N_46150,N_49679);
and UO_1292 (O_1292,N_48868,N_49795);
nor UO_1293 (O_1293,N_46142,N_47674);
nor UO_1294 (O_1294,N_48333,N_45820);
and UO_1295 (O_1295,N_45339,N_47162);
nand UO_1296 (O_1296,N_45723,N_49378);
and UO_1297 (O_1297,N_47959,N_47657);
and UO_1298 (O_1298,N_49092,N_45697);
and UO_1299 (O_1299,N_48603,N_46600);
or UO_1300 (O_1300,N_46031,N_49321);
xor UO_1301 (O_1301,N_48759,N_47010);
xor UO_1302 (O_1302,N_46842,N_45783);
and UO_1303 (O_1303,N_47540,N_47499);
nor UO_1304 (O_1304,N_49772,N_48049);
nand UO_1305 (O_1305,N_47469,N_46691);
nand UO_1306 (O_1306,N_46817,N_45447);
or UO_1307 (O_1307,N_49097,N_46202);
nand UO_1308 (O_1308,N_49774,N_47527);
or UO_1309 (O_1309,N_45166,N_46780);
nor UO_1310 (O_1310,N_46375,N_46344);
xnor UO_1311 (O_1311,N_46007,N_47673);
or UO_1312 (O_1312,N_46870,N_48084);
nand UO_1313 (O_1313,N_49951,N_49064);
xor UO_1314 (O_1314,N_47303,N_46799);
or UO_1315 (O_1315,N_49338,N_48030);
or UO_1316 (O_1316,N_45198,N_48246);
xor UO_1317 (O_1317,N_47592,N_47300);
nor UO_1318 (O_1318,N_49829,N_45309);
xor UO_1319 (O_1319,N_49837,N_47664);
xor UO_1320 (O_1320,N_48347,N_46472);
nand UO_1321 (O_1321,N_49202,N_48290);
nand UO_1322 (O_1322,N_47614,N_49167);
nor UO_1323 (O_1323,N_49651,N_45398);
nor UO_1324 (O_1324,N_46455,N_47934);
or UO_1325 (O_1325,N_45726,N_45110);
nand UO_1326 (O_1326,N_48230,N_45044);
nor UO_1327 (O_1327,N_49303,N_49159);
nand UO_1328 (O_1328,N_46535,N_47797);
and UO_1329 (O_1329,N_49728,N_45446);
xor UO_1330 (O_1330,N_48171,N_48550);
nor UO_1331 (O_1331,N_47736,N_49989);
and UO_1332 (O_1332,N_47093,N_45964);
xnor UO_1333 (O_1333,N_49355,N_46899);
nor UO_1334 (O_1334,N_45926,N_48667);
and UO_1335 (O_1335,N_49400,N_49065);
and UO_1336 (O_1336,N_46094,N_47434);
and UO_1337 (O_1337,N_49340,N_45320);
nor UO_1338 (O_1338,N_46880,N_46476);
and UO_1339 (O_1339,N_46666,N_49868);
nand UO_1340 (O_1340,N_48778,N_45187);
nand UO_1341 (O_1341,N_48524,N_45710);
or UO_1342 (O_1342,N_49244,N_45013);
nand UO_1343 (O_1343,N_49323,N_49377);
or UO_1344 (O_1344,N_45285,N_46298);
and UO_1345 (O_1345,N_45046,N_47936);
xor UO_1346 (O_1346,N_47646,N_46564);
and UO_1347 (O_1347,N_47969,N_49371);
or UO_1348 (O_1348,N_48342,N_45205);
and UO_1349 (O_1349,N_46830,N_45560);
and UO_1350 (O_1350,N_48757,N_49370);
nor UO_1351 (O_1351,N_45994,N_46068);
nor UO_1352 (O_1352,N_46908,N_45732);
nand UO_1353 (O_1353,N_47439,N_46700);
or UO_1354 (O_1354,N_45383,N_46963);
xnor UO_1355 (O_1355,N_49147,N_45742);
xnor UO_1356 (O_1356,N_48630,N_49216);
and UO_1357 (O_1357,N_48937,N_49120);
nor UO_1358 (O_1358,N_49151,N_46983);
xor UO_1359 (O_1359,N_46139,N_47741);
or UO_1360 (O_1360,N_48121,N_49053);
and UO_1361 (O_1361,N_49285,N_48522);
or UO_1362 (O_1362,N_45705,N_47243);
xor UO_1363 (O_1363,N_48199,N_45083);
nand UO_1364 (O_1364,N_47471,N_45852);
xor UO_1365 (O_1365,N_47832,N_45832);
nor UO_1366 (O_1366,N_49178,N_46123);
or UO_1367 (O_1367,N_48484,N_49123);
xnor UO_1368 (O_1368,N_49499,N_46828);
xnor UO_1369 (O_1369,N_46976,N_49286);
nand UO_1370 (O_1370,N_49616,N_45321);
nand UO_1371 (O_1371,N_48218,N_45963);
nor UO_1372 (O_1372,N_45651,N_47205);
and UO_1373 (O_1373,N_48478,N_47405);
and UO_1374 (O_1374,N_48151,N_48979);
nor UO_1375 (O_1375,N_47430,N_45112);
and UO_1376 (O_1376,N_46583,N_49070);
nor UO_1377 (O_1377,N_49050,N_47180);
nor UO_1378 (O_1378,N_49107,N_45676);
nand UO_1379 (O_1379,N_45492,N_49710);
nor UO_1380 (O_1380,N_49331,N_48863);
nand UO_1381 (O_1381,N_47661,N_45450);
and UO_1382 (O_1382,N_47487,N_46547);
or UO_1383 (O_1383,N_49452,N_46255);
xor UO_1384 (O_1384,N_48970,N_49075);
xor UO_1385 (O_1385,N_49558,N_48838);
and UO_1386 (O_1386,N_48502,N_48242);
xnor UO_1387 (O_1387,N_47185,N_47134);
xnor UO_1388 (O_1388,N_46024,N_49886);
nor UO_1389 (O_1389,N_45302,N_45281);
or UO_1390 (O_1390,N_49206,N_45132);
xnor UO_1391 (O_1391,N_47589,N_49273);
nor UO_1392 (O_1392,N_45645,N_46765);
or UO_1393 (O_1393,N_46736,N_48657);
or UO_1394 (O_1394,N_45920,N_48310);
nand UO_1395 (O_1395,N_48239,N_48216);
nor UO_1396 (O_1396,N_47268,N_47569);
xnor UO_1397 (O_1397,N_47308,N_45688);
nand UO_1398 (O_1398,N_46203,N_46037);
nor UO_1399 (O_1399,N_49078,N_49089);
nor UO_1400 (O_1400,N_49955,N_48874);
or UO_1401 (O_1401,N_45522,N_47411);
and UO_1402 (O_1402,N_45654,N_49839);
xor UO_1403 (O_1403,N_46776,N_47825);
and UO_1404 (O_1404,N_46155,N_48360);
nor UO_1405 (O_1405,N_48529,N_45226);
or UO_1406 (O_1406,N_47151,N_48736);
xor UO_1407 (O_1407,N_48287,N_49671);
and UO_1408 (O_1408,N_46798,N_49589);
xnor UO_1409 (O_1409,N_45904,N_45225);
or UO_1410 (O_1410,N_45675,N_47470);
nor UO_1411 (O_1411,N_49759,N_45826);
and UO_1412 (O_1412,N_45234,N_47229);
nand UO_1413 (O_1413,N_47199,N_47232);
nor UO_1414 (O_1414,N_48271,N_46162);
nand UO_1415 (O_1415,N_49106,N_45201);
and UO_1416 (O_1416,N_49298,N_46402);
or UO_1417 (O_1417,N_47813,N_46235);
nand UO_1418 (O_1418,N_46246,N_49003);
nor UO_1419 (O_1419,N_47179,N_49124);
nor UO_1420 (O_1420,N_47815,N_47436);
or UO_1421 (O_1421,N_47450,N_49317);
xor UO_1422 (O_1422,N_46458,N_49854);
xnor UO_1423 (O_1423,N_49573,N_49576);
nor UO_1424 (O_1424,N_46439,N_48670);
or UO_1425 (O_1425,N_49794,N_46486);
nor UO_1426 (O_1426,N_45827,N_49970);
and UO_1427 (O_1427,N_46483,N_46711);
and UO_1428 (O_1428,N_46020,N_45614);
or UO_1429 (O_1429,N_49856,N_45138);
and UO_1430 (O_1430,N_49205,N_47515);
or UO_1431 (O_1431,N_45754,N_48790);
nand UO_1432 (O_1432,N_48779,N_49253);
xnor UO_1433 (O_1433,N_45183,N_47452);
and UO_1434 (O_1434,N_46310,N_48468);
and UO_1435 (O_1435,N_45243,N_49314);
xnor UO_1436 (O_1436,N_48109,N_47375);
nor UO_1437 (O_1437,N_46355,N_45932);
xor UO_1438 (O_1438,N_46160,N_48804);
or UO_1439 (O_1439,N_48777,N_45337);
nand UO_1440 (O_1440,N_47563,N_47120);
and UO_1441 (O_1441,N_47219,N_45985);
nor UO_1442 (O_1442,N_46954,N_49302);
or UO_1443 (O_1443,N_47508,N_49048);
or UO_1444 (O_1444,N_45157,N_47501);
nand UO_1445 (O_1445,N_45363,N_47665);
nor UO_1446 (O_1446,N_47467,N_45764);
nand UO_1447 (O_1447,N_48628,N_48784);
nand UO_1448 (O_1448,N_49289,N_49986);
nor UO_1449 (O_1449,N_45992,N_45635);
nand UO_1450 (O_1450,N_46261,N_48495);
xor UO_1451 (O_1451,N_45835,N_47650);
xnor UO_1452 (O_1452,N_46053,N_45325);
xor UO_1453 (O_1453,N_46792,N_45433);
nand UO_1454 (O_1454,N_49720,N_47158);
xor UO_1455 (O_1455,N_46621,N_47160);
or UO_1456 (O_1456,N_48533,N_49872);
xnor UO_1457 (O_1457,N_49140,N_46994);
nand UO_1458 (O_1458,N_47414,N_48871);
nand UO_1459 (O_1459,N_48971,N_49818);
nor UO_1460 (O_1460,N_46608,N_45766);
nor UO_1461 (O_1461,N_47740,N_45002);
or UO_1462 (O_1462,N_46680,N_45850);
nor UO_1463 (O_1463,N_49593,N_45258);
or UO_1464 (O_1464,N_48547,N_47956);
xnor UO_1465 (O_1465,N_49801,N_49284);
xnor UO_1466 (O_1466,N_49403,N_47090);
or UO_1467 (O_1467,N_48035,N_48052);
and UO_1468 (O_1468,N_49099,N_47039);
and UO_1469 (O_1469,N_49334,N_46134);
nand UO_1470 (O_1470,N_47907,N_47283);
xnor UO_1471 (O_1471,N_49760,N_47449);
nor UO_1472 (O_1472,N_47942,N_47392);
nand UO_1473 (O_1473,N_45981,N_48899);
and UO_1474 (O_1474,N_46050,N_45542);
or UO_1475 (O_1475,N_49328,N_49954);
nor UO_1476 (O_1476,N_48186,N_49550);
nor UO_1477 (O_1477,N_46184,N_49866);
xnor UO_1478 (O_1478,N_48624,N_47325);
or UO_1479 (O_1479,N_47230,N_45094);
nand UO_1480 (O_1480,N_47287,N_48393);
nand UO_1481 (O_1481,N_47459,N_46218);
nand UO_1482 (O_1482,N_49544,N_48175);
xnor UO_1483 (O_1483,N_46245,N_49343);
and UO_1484 (O_1484,N_48586,N_48095);
and UO_1485 (O_1485,N_48284,N_48391);
nand UO_1486 (O_1486,N_49568,N_49867);
xnor UO_1487 (O_1487,N_49194,N_48048);
or UO_1488 (O_1488,N_47541,N_48000);
xnor UO_1489 (O_1489,N_45060,N_49601);
and UO_1490 (O_1490,N_45772,N_47901);
or UO_1491 (O_1491,N_49825,N_45677);
or UO_1492 (O_1492,N_48748,N_47521);
nand UO_1493 (O_1493,N_45986,N_45072);
and UO_1494 (O_1494,N_46950,N_45592);
nor UO_1495 (O_1495,N_49943,N_45023);
nor UO_1496 (O_1496,N_47680,N_49129);
and UO_1497 (O_1497,N_45621,N_49859);
nand UO_1498 (O_1498,N_48301,N_49775);
nor UO_1499 (O_1499,N_48856,N_46932);
nand UO_1500 (O_1500,N_49840,N_48096);
xor UO_1501 (O_1501,N_47493,N_47860);
nand UO_1502 (O_1502,N_48674,N_46578);
nor UO_1503 (O_1503,N_49439,N_48079);
or UO_1504 (O_1504,N_48041,N_49471);
or UO_1505 (O_1505,N_45776,N_47054);
or UO_1506 (O_1506,N_48690,N_45327);
nor UO_1507 (O_1507,N_45971,N_47307);
nand UO_1508 (O_1508,N_48541,N_48247);
nor UO_1509 (O_1509,N_47977,N_45757);
nand UO_1510 (O_1510,N_49765,N_45074);
and UO_1511 (O_1511,N_46903,N_46054);
or UO_1512 (O_1512,N_47796,N_47769);
nand UO_1513 (O_1513,N_47638,N_45388);
xnor UO_1514 (O_1514,N_47027,N_48018);
and UO_1515 (O_1515,N_46991,N_47415);
nor UO_1516 (O_1516,N_46408,N_48976);
and UO_1517 (O_1517,N_48936,N_46120);
nor UO_1518 (O_1518,N_46560,N_49443);
and UO_1519 (O_1519,N_48353,N_48011);
nor UO_1520 (O_1520,N_47178,N_48986);
nand UO_1521 (O_1521,N_47768,N_47719);
and UO_1522 (O_1522,N_46956,N_48329);
nor UO_1523 (O_1523,N_48849,N_45057);
and UO_1524 (O_1524,N_47188,N_45857);
or UO_1525 (O_1525,N_49476,N_47190);
or UO_1526 (O_1526,N_46840,N_47981);
and UO_1527 (O_1527,N_47856,N_46381);
xor UO_1528 (O_1528,N_45221,N_49203);
and UO_1529 (O_1529,N_45898,N_46630);
nor UO_1530 (O_1530,N_48004,N_49600);
nor UO_1531 (O_1531,N_49626,N_48312);
xnor UO_1532 (O_1532,N_46052,N_46309);
and UO_1533 (O_1533,N_47418,N_45478);
xor UO_1534 (O_1534,N_48003,N_45773);
nand UO_1535 (O_1535,N_48869,N_46967);
xor UO_1536 (O_1536,N_49350,N_47584);
nor UO_1537 (O_1537,N_45432,N_46268);
or UO_1538 (O_1538,N_49689,N_47616);
or UO_1539 (O_1539,N_48999,N_48728);
nand UO_1540 (O_1540,N_48162,N_48588);
nand UO_1541 (O_1541,N_49292,N_47550);
and UO_1542 (O_1542,N_48655,N_45098);
and UO_1543 (O_1543,N_48448,N_45796);
nor UO_1544 (O_1544,N_47412,N_45411);
nand UO_1545 (O_1545,N_49591,N_47445);
nand UO_1546 (O_1546,N_46349,N_48265);
xor UO_1547 (O_1547,N_47980,N_49270);
nand UO_1548 (O_1548,N_46456,N_47851);
nor UO_1549 (O_1549,N_45717,N_49030);
xnor UO_1550 (O_1550,N_49507,N_45906);
nor UO_1551 (O_1551,N_46589,N_47760);
or UO_1552 (O_1552,N_46833,N_49858);
xor UO_1553 (O_1553,N_49407,N_47033);
or UO_1554 (O_1554,N_49052,N_46505);
xnor UO_1555 (O_1555,N_48319,N_47568);
or UO_1556 (O_1556,N_49631,N_48315);
and UO_1557 (O_1557,N_45900,N_46323);
and UO_1558 (O_1558,N_47772,N_47069);
or UO_1559 (O_1559,N_47774,N_47635);
xor UO_1560 (O_1560,N_47695,N_48589);
nor UO_1561 (O_1561,N_48112,N_46683);
or UO_1562 (O_1562,N_49773,N_48730);
or UO_1563 (O_1563,N_45293,N_45154);
or UO_1564 (O_1564,N_48085,N_45086);
or UO_1565 (O_1565,N_46540,N_45743);
and UO_1566 (O_1566,N_47785,N_47244);
nand UO_1567 (O_1567,N_47024,N_45051);
xor UO_1568 (O_1568,N_45913,N_47913);
nor UO_1569 (O_1569,N_49572,N_46528);
xnor UO_1570 (O_1570,N_45428,N_46093);
and UO_1571 (O_1571,N_47816,N_47647);
or UO_1572 (O_1572,N_46412,N_45894);
nor UO_1573 (O_1573,N_48582,N_45113);
or UO_1574 (O_1574,N_48056,N_47529);
and UO_1575 (O_1575,N_45217,N_47237);
nor UO_1576 (O_1576,N_49184,N_45600);
and UO_1577 (O_1577,N_48400,N_49747);
nand UO_1578 (O_1578,N_46432,N_47351);
nand UO_1579 (O_1579,N_45744,N_47184);
or UO_1580 (O_1580,N_46247,N_48213);
xnor UO_1581 (O_1581,N_45015,N_47082);
or UO_1582 (O_1582,N_49280,N_45980);
nand UO_1583 (O_1583,N_47056,N_49644);
xor UO_1584 (O_1584,N_49356,N_48809);
nor UO_1585 (O_1585,N_49802,N_49088);
xnor UO_1586 (O_1586,N_48281,N_49166);
and UO_1587 (O_1587,N_45340,N_46745);
nand UO_1588 (O_1588,N_48245,N_48832);
nand UO_1589 (O_1589,N_49182,N_46028);
nor UO_1590 (O_1590,N_49011,N_45622);
or UO_1591 (O_1591,N_45816,N_46843);
or UO_1592 (O_1592,N_47488,N_47732);
xnor UO_1593 (O_1593,N_46809,N_45825);
nand UO_1594 (O_1594,N_49778,N_47518);
nand UO_1595 (O_1595,N_45014,N_47625);
nand UO_1596 (O_1596,N_45194,N_46881);
and UO_1597 (O_1597,N_47050,N_47585);
nand UO_1598 (O_1598,N_47608,N_49585);
and UO_1599 (O_1599,N_48709,N_47723);
nor UO_1600 (O_1600,N_49967,N_47273);
xnor UO_1601 (O_1601,N_48564,N_49102);
nand UO_1602 (O_1602,N_45655,N_49918);
or UO_1603 (O_1603,N_48613,N_48889);
or UO_1604 (O_1604,N_49788,N_45696);
xor UO_1605 (O_1605,N_49294,N_45431);
and UO_1606 (O_1606,N_46603,N_49186);
nand UO_1607 (O_1607,N_48955,N_47803);
nand UO_1608 (O_1608,N_47841,N_45664);
nor UO_1609 (O_1609,N_49352,N_46157);
or UO_1610 (O_1610,N_48570,N_45359);
nor UO_1611 (O_1611,N_47875,N_49183);
xor UO_1612 (O_1612,N_47880,N_47586);
and UO_1613 (O_1613,N_48374,N_46192);
and UO_1614 (O_1614,N_49225,N_48219);
nand UO_1615 (O_1615,N_47915,N_45195);
xor UO_1616 (O_1616,N_48501,N_45896);
and UO_1617 (O_1617,N_46271,N_46914);
xnor UO_1618 (O_1618,N_49252,N_45714);
xnor UO_1619 (O_1619,N_45264,N_45102);
and UO_1620 (O_1620,N_46729,N_45889);
and UO_1621 (O_1621,N_49896,N_46590);
nand UO_1622 (O_1622,N_47348,N_45455);
and UO_1623 (O_1623,N_45997,N_46697);
nand UO_1624 (O_1624,N_46919,N_48845);
nand UO_1625 (O_1625,N_46778,N_48854);
nand UO_1626 (O_1626,N_45536,N_45901);
and UO_1627 (O_1627,N_48960,N_49819);
and UO_1628 (O_1628,N_47703,N_45437);
or UO_1629 (O_1629,N_48629,N_45012);
xor UO_1630 (O_1630,N_45706,N_47332);
nand UO_1631 (O_1631,N_46131,N_45956);
and UO_1632 (O_1632,N_49461,N_48479);
nand UO_1633 (O_1633,N_46714,N_48952);
nand UO_1634 (O_1634,N_46366,N_45438);
nor UO_1635 (O_1635,N_45405,N_47877);
and UO_1636 (O_1636,N_47781,N_47881);
nor UO_1637 (O_1637,N_45474,N_47791);
nand UO_1638 (O_1638,N_49041,N_48345);
nand UO_1639 (O_1639,N_47221,N_45960);
nor UO_1640 (O_1640,N_47261,N_45490);
or UO_1641 (O_1641,N_45256,N_48254);
nand UO_1642 (O_1642,N_48220,N_48014);
or UO_1643 (O_1643,N_47624,N_47545);
xor UO_1644 (O_1644,N_46396,N_49823);
nor UO_1645 (O_1645,N_46287,N_47854);
nand UO_1646 (O_1646,N_47315,N_46180);
and UO_1647 (O_1647,N_45782,N_46825);
nor UO_1648 (O_1648,N_49623,N_48638);
nand UO_1649 (O_1649,N_48823,N_45713);
nor UO_1650 (O_1650,N_47291,N_45186);
nand UO_1651 (O_1651,N_49433,N_46682);
xnor UO_1652 (O_1652,N_48866,N_48901);
and UO_1653 (O_1653,N_46849,N_48933);
nor UO_1654 (O_1654,N_48978,N_46222);
or UO_1655 (O_1655,N_49922,N_47084);
xnor UO_1656 (O_1656,N_46732,N_46534);
or UO_1657 (O_1657,N_47717,N_47031);
or UO_1658 (O_1658,N_49769,N_47850);
or UO_1659 (O_1659,N_47610,N_45093);
nor UO_1660 (O_1660,N_46864,N_48893);
xor UO_1661 (O_1661,N_45148,N_49177);
nor UO_1662 (O_1662,N_49354,N_46479);
xnor UO_1663 (O_1663,N_49438,N_48023);
nor UO_1664 (O_1664,N_46411,N_48822);
and UO_1665 (O_1665,N_47374,N_45464);
nand UO_1666 (O_1666,N_45585,N_47909);
nand UO_1667 (O_1667,N_49066,N_46316);
nand UO_1668 (O_1668,N_47107,N_47409);
xor UO_1669 (O_1669,N_49389,N_46135);
nand UO_1670 (O_1670,N_49516,N_45085);
nand UO_1671 (O_1671,N_47745,N_46702);
nand UO_1672 (O_1672,N_45979,N_45020);
nor UO_1673 (O_1673,N_46399,N_48659);
nand UO_1674 (O_1674,N_46219,N_46889);
xor UO_1675 (O_1675,N_49498,N_49110);
nor UO_1676 (O_1676,N_48734,N_47517);
nand UO_1677 (O_1677,N_49141,N_45786);
nand UO_1678 (O_1678,N_45119,N_47597);
or UO_1679 (O_1679,N_47823,N_48055);
nor UO_1680 (O_1680,N_46317,N_45463);
or UO_1681 (O_1681,N_45882,N_46133);
or UO_1682 (O_1682,N_45763,N_46624);
or UO_1683 (O_1683,N_45887,N_46273);
or UO_1684 (O_1684,N_48223,N_48696);
and UO_1685 (O_1685,N_47557,N_49344);
and UO_1686 (O_1686,N_45745,N_45135);
and UO_1687 (O_1687,N_46782,N_48625);
nor UO_1688 (O_1688,N_49179,N_47318);
and UO_1689 (O_1689,N_49022,N_49409);
or UO_1690 (O_1690,N_47127,N_46100);
and UO_1691 (O_1691,N_49694,N_47549);
xor UO_1692 (O_1692,N_47937,N_45532);
xor UO_1693 (O_1693,N_49923,N_46029);
xnor UO_1694 (O_1694,N_46758,N_45009);
xor UO_1695 (O_1695,N_46447,N_49642);
nor UO_1696 (O_1696,N_47407,N_47182);
xnor UO_1697 (O_1697,N_46961,N_49374);
xor UO_1698 (O_1698,N_45305,N_48467);
nor UO_1699 (O_1699,N_49287,N_48635);
nor UO_1700 (O_1700,N_45440,N_46582);
and UO_1701 (O_1701,N_48510,N_49281);
xnor UO_1702 (O_1702,N_48743,N_46223);
nor UO_1703 (O_1703,N_49044,N_49578);
nor UO_1704 (O_1704,N_48686,N_46606);
nand UO_1705 (O_1705,N_45036,N_49269);
and UO_1706 (O_1706,N_49809,N_46536);
nor UO_1707 (O_1707,N_49929,N_47115);
and UO_1708 (O_1708,N_48197,N_46937);
and UO_1709 (O_1709,N_49519,N_48723);
nor UO_1710 (O_1710,N_48307,N_48609);
or UO_1711 (O_1711,N_49799,N_47065);
xor UO_1712 (O_1712,N_49445,N_47153);
nand UO_1713 (O_1713,N_46216,N_46911);
nand UO_1714 (O_1714,N_46069,N_47327);
xnor UO_1715 (O_1715,N_46663,N_45435);
nand UO_1716 (O_1716,N_48390,N_45429);
nor UO_1717 (O_1717,N_49947,N_45211);
nand UO_1718 (O_1718,N_48610,N_48711);
xor UO_1719 (O_1719,N_47943,N_46859);
nand UO_1720 (O_1720,N_47718,N_48654);
and UO_1721 (O_1721,N_46444,N_46921);
and UO_1722 (O_1722,N_46657,N_48334);
or UO_1723 (O_1723,N_48376,N_48509);
and UO_1724 (O_1724,N_46902,N_48825);
nor UO_1725 (O_1725,N_46158,N_46300);
nand UO_1726 (O_1726,N_47092,N_46694);
nor UO_1727 (O_1727,N_47994,N_45156);
and UO_1728 (O_1728,N_46542,N_48053);
xnor UO_1729 (O_1729,N_49047,N_46513);
nand UO_1730 (O_1730,N_48002,N_48578);
and UO_1731 (O_1731,N_45949,N_49137);
and UO_1732 (O_1732,N_46561,N_47688);
nor UO_1733 (O_1733,N_47971,N_48306);
or UO_1734 (O_1734,N_48460,N_45244);
or UO_1735 (O_1735,N_45950,N_49169);
or UO_1736 (O_1736,N_46934,N_49145);
and UO_1737 (O_1737,N_48369,N_45858);
and UO_1738 (O_1738,N_49073,N_46164);
nand UO_1739 (O_1739,N_49361,N_49363);
or UO_1740 (O_1740,N_49247,N_47928);
nand UO_1741 (O_1741,N_49673,N_47041);
nand UO_1742 (O_1742,N_46077,N_45541);
nand UO_1743 (O_1743,N_48913,N_48308);
nand UO_1744 (O_1744,N_45538,N_46596);
and UO_1745 (O_1745,N_47198,N_47574);
nand UO_1746 (O_1746,N_47706,N_45378);
or UO_1747 (O_1747,N_46912,N_48429);
or UO_1748 (O_1748,N_46684,N_46854);
or UO_1749 (O_1749,N_46122,N_46188);
or UO_1750 (O_1750,N_46518,N_45164);
xor UO_1751 (O_1751,N_46391,N_48847);
nand UO_1752 (O_1752,N_48364,N_45434);
or UO_1753 (O_1753,N_45712,N_45843);
and UO_1754 (O_1754,N_46860,N_48065);
nor UO_1755 (O_1755,N_49322,N_46406);
xnor UO_1756 (O_1756,N_47908,N_49817);
or UO_1757 (O_1757,N_46787,N_48408);
or UO_1758 (O_1758,N_45191,N_46413);
or UO_1759 (O_1759,N_47468,N_45361);
nor UO_1760 (O_1760,N_47364,N_48882);
nand UO_1761 (O_1761,N_47213,N_45246);
nor UO_1762 (O_1762,N_46230,N_49725);
nor UO_1763 (O_1763,N_49063,N_47935);
nand UO_1764 (O_1764,N_47588,N_45606);
nand UO_1765 (O_1765,N_47777,N_46658);
and UO_1766 (O_1766,N_48226,N_48135);
nor UO_1767 (O_1767,N_48717,N_46553);
xnor UO_1768 (O_1768,N_48862,N_49761);
or UO_1769 (O_1769,N_47759,N_48438);
nand UO_1770 (O_1770,N_47113,N_46418);
nand UO_1771 (O_1771,N_48267,N_49300);
and UO_1772 (O_1772,N_48024,N_46299);
nor UO_1773 (O_1773,N_49611,N_49731);
nand UO_1774 (O_1774,N_48103,N_49329);
xnor UO_1775 (O_1775,N_45552,N_49685);
or UO_1776 (O_1776,N_45518,N_49879);
and UO_1777 (O_1777,N_47761,N_49758);
xor UO_1778 (O_1778,N_46087,N_45442);
xnor UO_1779 (O_1779,N_47888,N_46198);
nand UO_1780 (O_1780,N_49503,N_48945);
and UO_1781 (O_1781,N_46283,N_45417);
nand UO_1782 (O_1782,N_46611,N_45047);
or UO_1783 (O_1783,N_49701,N_49515);
nor UO_1784 (O_1784,N_47384,N_47845);
or UO_1785 (O_1785,N_48205,N_47257);
and UO_1786 (O_1786,N_47960,N_45576);
xor UO_1787 (O_1787,N_45038,N_49928);
nand UO_1788 (O_1788,N_48642,N_48562);
xnor UO_1789 (O_1789,N_46461,N_47818);
or UO_1790 (O_1790,N_47456,N_48362);
nor UO_1791 (O_1791,N_45008,N_45643);
or UO_1792 (O_1792,N_47455,N_46735);
xnor UO_1793 (O_1793,N_45275,N_46592);
nor UO_1794 (O_1794,N_47572,N_48914);
nand UO_1795 (O_1795,N_46431,N_45298);
nand UO_1796 (O_1796,N_48820,N_47328);
nor UO_1797 (O_1797,N_48462,N_46978);
nand UO_1798 (O_1798,N_47686,N_45811);
nand UO_1799 (O_1799,N_47347,N_47750);
and UO_1800 (O_1800,N_45781,N_45042);
nand UO_1801 (O_1801,N_46968,N_49060);
nand UO_1802 (O_1802,N_45869,N_48530);
xnor UO_1803 (O_1803,N_49291,N_48188);
xor UO_1804 (O_1804,N_49027,N_47636);
or UO_1805 (O_1805,N_47297,N_46369);
nor UO_1806 (O_1806,N_48552,N_46263);
and UO_1807 (O_1807,N_49620,N_49571);
nand UO_1808 (O_1808,N_46468,N_47015);
and UO_1809 (O_1809,N_49282,N_45807);
and UO_1810 (O_1810,N_47363,N_45260);
nor UO_1811 (O_1811,N_46185,N_46503);
nor UO_1812 (O_1812,N_48370,N_46356);
nor UO_1813 (O_1813,N_47066,N_48705);
and UO_1814 (O_1814,N_49687,N_45055);
and UO_1815 (O_1815,N_46288,N_49994);
nor UO_1816 (O_1816,N_46275,N_47321);
xor UO_1817 (O_1817,N_46883,N_46141);
xnor UO_1818 (O_1818,N_45185,N_48289);
xor UO_1819 (O_1819,N_45647,N_46811);
or UO_1820 (O_1820,N_48261,N_49150);
nor UO_1821 (O_1821,N_45422,N_47986);
nor UO_1822 (O_1822,N_46154,N_49618);
xnor UO_1823 (O_1823,N_45082,N_49271);
and UO_1824 (O_1824,N_47983,N_47239);
and UO_1825 (O_1825,N_47051,N_45617);
and UO_1826 (O_1826,N_48499,N_49213);
nor UO_1827 (O_1827,N_48126,N_46888);
and UO_1828 (O_1828,N_46114,N_45184);
nand UO_1829 (O_1829,N_47083,N_47311);
nand UO_1830 (O_1830,N_48383,N_49998);
xor UO_1831 (O_1831,N_48108,N_46676);
or UO_1832 (O_1832,N_45977,N_47558);
xnor UO_1833 (O_1833,N_48476,N_45000);
or UO_1834 (O_1834,N_45809,N_46362);
nand UO_1835 (O_1835,N_45216,N_47871);
nor UO_1836 (O_1836,N_46387,N_47896);
or UO_1837 (O_1837,N_48421,N_47355);
nand UO_1838 (O_1838,N_47147,N_49883);
nor UO_1839 (O_1839,N_46740,N_49848);
and UO_1840 (O_1840,N_49693,N_48278);
and UO_1841 (O_1841,N_48720,N_45605);
xnor UO_1842 (O_1842,N_46554,N_45003);
and UO_1843 (O_1843,N_47810,N_47421);
nor UO_1844 (O_1844,N_49134,N_49844);
and UO_1845 (O_1845,N_48054,N_48660);
nor UO_1846 (O_1846,N_46605,N_45559);
xor UO_1847 (O_1847,N_47962,N_45902);
and UO_1848 (O_1848,N_46664,N_46522);
and UO_1849 (O_1849,N_47903,N_46731);
or UO_1850 (O_1850,N_45409,N_45942);
and UO_1851 (O_1851,N_49692,N_47336);
xnor UO_1852 (O_1852,N_46998,N_45895);
xor UO_1853 (O_1853,N_49526,N_47187);
or UO_1854 (O_1854,N_46989,N_45210);
and UO_1855 (O_1855,N_46715,N_48646);
and UO_1856 (O_1856,N_45531,N_49072);
or UO_1857 (O_1857,N_48184,N_49894);
and UO_1858 (O_1858,N_46311,N_48129);
and UO_1859 (O_1859,N_47271,N_47406);
nand UO_1860 (O_1860,N_45728,N_46722);
and UO_1861 (O_1861,N_49598,N_47379);
and UO_1862 (O_1862,N_48122,N_49932);
xnor UO_1863 (O_1863,N_45611,N_48583);
and UO_1864 (O_1864,N_47632,N_49658);
xnor UO_1865 (O_1865,N_48855,N_46641);
and UO_1866 (O_1866,N_47309,N_48536);
or UO_1867 (O_1867,N_49349,N_47446);
xor UO_1868 (O_1868,N_49039,N_48350);
and UO_1869 (O_1869,N_49482,N_47715);
and UO_1870 (O_1870,N_45636,N_49154);
xor UO_1871 (O_1871,N_48439,N_46763);
or UO_1872 (O_1872,N_45288,N_48651);
or UO_1873 (O_1873,N_48093,N_45589);
and UO_1874 (O_1874,N_46378,N_48687);
xor UO_1875 (O_1875,N_45120,N_46748);
nand UO_1876 (O_1876,N_46109,N_46988);
or UO_1877 (O_1877,N_47394,N_45165);
nand UO_1878 (O_1878,N_49949,N_46295);
or UO_1879 (O_1879,N_46256,N_47402);
or UO_1880 (O_1880,N_48417,N_47692);
xnor UO_1881 (O_1881,N_49617,N_49196);
nand UO_1882 (O_1882,N_47984,N_45870);
nor UO_1883 (O_1883,N_49912,N_49880);
xnor UO_1884 (O_1884,N_48980,N_48078);
and UO_1885 (O_1885,N_45290,N_47682);
and UO_1886 (O_1886,N_48704,N_45459);
or UO_1887 (O_1887,N_47734,N_47944);
or UO_1888 (O_1888,N_49373,N_48305);
nor UO_1889 (O_1889,N_48237,N_46101);
nor UO_1890 (O_1890,N_46210,N_47272);
and UO_1891 (O_1891,N_49223,N_48236);
nand UO_1892 (O_1892,N_49080,N_45789);
and UO_1893 (O_1893,N_45533,N_45366);
or UO_1894 (O_1894,N_49606,N_47099);
nand UO_1895 (O_1895,N_45001,N_46770);
nor UO_1896 (O_1896,N_49031,N_45367);
or UO_1897 (O_1897,N_48829,N_46871);
xor UO_1898 (O_1898,N_48747,N_48104);
xor UO_1899 (O_1899,N_48298,N_45374);
or UO_1900 (O_1900,N_45649,N_48940);
nand UO_1901 (O_1901,N_49148,N_48064);
nor UO_1902 (O_1902,N_47583,N_48527);
and UO_1903 (O_1903,N_45821,N_45171);
nor UO_1904 (O_1904,N_46990,N_49588);
and UO_1905 (O_1905,N_49122,N_48662);
nor UO_1906 (O_1906,N_47018,N_47250);
nand UO_1907 (O_1907,N_48379,N_49664);
xor UO_1908 (O_1908,N_49404,N_48939);
nand UO_1909 (O_1909,N_47542,N_48015);
nor UO_1910 (O_1910,N_48145,N_46834);
nor UO_1911 (O_1911,N_47922,N_48879);
or UO_1912 (O_1912,N_45629,N_48061);
and UO_1913 (O_1913,N_45613,N_45287);
nor UO_1914 (O_1914,N_46789,N_45951);
and UO_1915 (O_1915,N_46467,N_48098);
xnor UO_1916 (O_1916,N_48637,N_45131);
nor UO_1917 (O_1917,N_45484,N_48707);
xnor UO_1918 (O_1918,N_47137,N_49144);
and UO_1919 (O_1919,N_49098,N_49757);
nand UO_1920 (O_1920,N_45797,N_46533);
and UO_1921 (O_1921,N_46509,N_47140);
and UO_1922 (O_1922,N_49336,N_45323);
and UO_1923 (O_1923,N_45137,N_45308);
nor UO_1924 (O_1924,N_49449,N_48987);
and UO_1925 (O_1925,N_48985,N_47613);
xor UO_1926 (O_1926,N_46190,N_49153);
nor UO_1927 (O_1927,N_45149,N_49580);
and UO_1928 (O_1928,N_49479,N_45644);
or UO_1929 (O_1929,N_49639,N_46277);
and UO_1930 (O_1930,N_49637,N_48286);
or UO_1931 (O_1931,N_46388,N_47566);
xor UO_1932 (O_1932,N_45848,N_45245);
and UO_1933 (O_1933,N_48907,N_46634);
nand UO_1934 (O_1934,N_49677,N_47295);
nand UO_1935 (O_1935,N_46146,N_45711);
or UO_1936 (O_1936,N_48658,N_47752);
xnor UO_1937 (O_1937,N_45976,N_49036);
xnor UO_1938 (O_1938,N_48783,N_46928);
nor UO_1939 (O_1939,N_46176,N_49121);
and UO_1940 (O_1940,N_49643,N_48669);
nor UO_1941 (O_1941,N_46862,N_49108);
or UO_1942 (O_1942,N_49965,N_49614);
or UO_1943 (O_1943,N_46747,N_45563);
nor UO_1944 (O_1944,N_49990,N_45755);
xnor UO_1945 (O_1945,N_48033,N_47678);
nor UO_1946 (O_1946,N_47165,N_49865);
xor UO_1947 (O_1947,N_49985,N_49480);
and UO_1948 (O_1948,N_47014,N_48110);
xor UO_1949 (O_1949,N_47679,N_47201);
nor UO_1950 (O_1950,N_45081,N_47730);
or UO_1951 (O_1951,N_45024,N_47383);
xor UO_1952 (O_1952,N_48318,N_46844);
nor UO_1953 (O_1953,N_46725,N_47472);
nor UO_1954 (O_1954,N_47793,N_46501);
xor UO_1955 (O_1955,N_48255,N_45761);
nand UO_1956 (O_1956,N_48560,N_45347);
or UO_1957 (O_1957,N_47967,N_46756);
xnor UO_1958 (O_1958,N_49648,N_45141);
xnor UO_1959 (O_1959,N_45421,N_46250);
nor UO_1960 (O_1960,N_49276,N_48363);
and UO_1961 (O_1961,N_47917,N_49390);
nor UO_1962 (O_1962,N_45524,N_47422);
xnor UO_1963 (O_1963,N_47135,N_48332);
nand UO_1964 (O_1964,N_45785,N_48317);
nand UO_1965 (O_1965,N_46208,N_46886);
nor UO_1966 (O_1966,N_46462,N_47885);
xnor UO_1967 (O_1967,N_45197,N_46620);
nor UO_1968 (O_1968,N_46861,N_48375);
and UO_1969 (O_1969,N_46438,N_45247);
nand UO_1970 (O_1970,N_48816,N_49796);
nor UO_1971 (O_1971,N_48892,N_46612);
xnor UO_1972 (O_1972,N_49997,N_45123);
nand UO_1973 (O_1973,N_45724,N_46019);
nand UO_1974 (O_1974,N_49233,N_49201);
or UO_1975 (O_1975,N_48612,N_48531);
or UO_1976 (O_1976,N_48742,N_47226);
nand UO_1977 (O_1977,N_48368,N_49652);
xnor UO_1978 (O_1978,N_48241,N_45855);
xnor UO_1979 (O_1979,N_45096,N_49494);
xor UO_1980 (O_1980,N_49752,N_49295);
and UO_1981 (O_1981,N_49852,N_47879);
or UO_1982 (O_1982,N_48277,N_46004);
nor UO_1983 (O_1983,N_47609,N_47401);
or UO_1984 (O_1984,N_47573,N_48910);
and UO_1985 (O_1985,N_48966,N_48700);
xor UO_1986 (O_1986,N_48128,N_48577);
nand UO_1987 (O_1987,N_45908,N_45266);
nor UO_1988 (O_1988,N_49057,N_46073);
nand UO_1989 (O_1989,N_46900,N_46080);
nor UO_1990 (O_1990,N_46945,N_47275);
and UO_1991 (O_1991,N_49559,N_45694);
nor UO_1992 (O_1992,N_47366,N_46541);
nor UO_1993 (O_1993,N_47957,N_47577);
and UO_1994 (O_1994,N_49015,N_46191);
nor UO_1995 (O_1995,N_48371,N_45619);
or UO_1996 (O_1996,N_46481,N_47628);
or UO_1997 (O_1997,N_47950,N_45153);
or UO_1998 (O_1998,N_49863,N_46774);
or UO_1999 (O_1999,N_48668,N_47834);
nand UO_2000 (O_2000,N_49375,N_48968);
and UO_2001 (O_2001,N_48930,N_46179);
and UO_2002 (O_2002,N_48948,N_49808);
nand UO_2003 (O_2003,N_48518,N_47424);
and UO_2004 (O_2004,N_49410,N_47352);
and UO_2005 (O_2005,N_45196,N_48672);
nor UO_2006 (O_2006,N_46015,N_46353);
and UO_2007 (O_2007,N_47030,N_45927);
and UO_2008 (O_2008,N_45570,N_46728);
nand UO_2009 (O_2009,N_47164,N_47387);
nand UO_2010 (O_2010,N_46067,N_45633);
or UO_2011 (O_2011,N_46783,N_45204);
nor UO_2012 (O_2012,N_49058,N_46348);
xor UO_2013 (O_2013,N_45890,N_45139);
and UO_2014 (O_2014,N_48523,N_47509);
and UO_2015 (O_2015,N_47949,N_49939);
nor UO_2016 (O_2016,N_46178,N_46733);
or UO_2017 (O_2017,N_47524,N_49369);
nand UO_2018 (O_2018,N_46609,N_45313);
nor UO_2019 (O_2019,N_47305,N_45249);
nand UO_2020 (O_2020,N_49125,N_45236);
xnor UO_2021 (O_2021,N_47805,N_45678);
nor UO_2022 (O_2022,N_47144,N_45884);
xor UO_2023 (O_2023,N_48840,N_46325);
or UO_2024 (O_2024,N_46337,N_47241);
and UO_2025 (O_2025,N_45801,N_48268);
xor UO_2026 (O_2026,N_49222,N_48165);
xnor UO_2027 (O_2027,N_45371,N_47519);
or UO_2028 (O_2028,N_49095,N_48553);
nor UO_2029 (O_2029,N_46442,N_46074);
xnor UO_2030 (O_2030,N_45670,N_48810);
or UO_2031 (O_2031,N_45070,N_46801);
nor UO_2032 (O_2032,N_46717,N_49069);
or UO_2033 (O_2033,N_45562,N_46754);
xnor UO_2034 (O_2034,N_46845,N_48466);
and UO_2035 (O_2035,N_48204,N_46106);
nand UO_2036 (O_2036,N_49346,N_45968);
or UO_2037 (O_2037,N_45571,N_45719);
nand UO_2038 (O_2038,N_45881,N_46248);
or UO_2039 (O_2039,N_48944,N_46855);
nand UO_2040 (O_2040,N_48113,N_49732);
xor UO_2041 (O_2041,N_48865,N_45360);
or UO_2042 (O_2042,N_49719,N_45547);
nor UO_2043 (O_2043,N_45897,N_45190);
and UO_2044 (O_2044,N_47552,N_46217);
or UO_2045 (O_2045,N_49810,N_49740);
or UO_2046 (O_2046,N_48433,N_46938);
or UO_2047 (O_2047,N_47391,N_49996);
xnor UO_2048 (O_2048,N_49170,N_45652);
and UO_2049 (O_2049,N_49227,N_49797);
or UO_2050 (O_2050,N_49768,N_45498);
nor UO_2051 (O_2051,N_47354,N_49245);
nand UO_2052 (O_2052,N_48067,N_47398);
or UO_2053 (O_2053,N_47543,N_46425);
nor UO_2054 (O_2054,N_45695,N_48394);
and UO_2055 (O_2055,N_46313,N_48864);
and UO_2056 (O_2056,N_46143,N_45124);
nand UO_2057 (O_2057,N_48217,N_47974);
nand UO_2058 (O_2058,N_49257,N_48470);
or UO_2059 (O_2059,N_45460,N_47631);
xnor UO_2060 (O_2060,N_47132,N_46706);
nand UO_2061 (O_2061,N_45037,N_46753);
or UO_2062 (O_2062,N_48808,N_49680);
nor UO_2063 (O_2063,N_48346,N_49563);
xnor UO_2064 (O_2064,N_48788,N_47049);
or UO_2065 (O_2065,N_47228,N_45111);
or UO_2066 (O_2066,N_48514,N_45272);
xnor UO_2067 (O_2067,N_48943,N_46665);
or UO_2068 (O_2068,N_48776,N_47427);
nand UO_2069 (O_2069,N_48125,N_47139);
nand UO_2070 (O_2070,N_48322,N_46290);
xnor UO_2071 (O_2071,N_47277,N_49454);
and UO_2072 (O_2072,N_48182,N_45390);
or UO_2073 (O_2073,N_46386,N_49704);
and UO_2074 (O_2074,N_45886,N_47357);
and UO_2075 (O_2075,N_45423,N_48238);
and UO_2076 (O_2076,N_45599,N_48766);
nand UO_2077 (O_2077,N_45909,N_48792);
xor UO_2078 (O_2078,N_49521,N_49487);
nand UO_2079 (O_2079,N_48106,N_48244);
and UO_2080 (O_2080,N_46750,N_47690);
xnor UO_2081 (O_2081,N_49565,N_47255);
nand UO_2082 (O_2082,N_45263,N_45689);
and UO_2083 (O_2083,N_47377,N_46519);
and UO_2084 (O_2084,N_49655,N_46047);
xnor UO_2085 (O_2085,N_49762,N_45065);
xnor UO_2086 (O_2086,N_48057,N_49038);
nor UO_2087 (O_2087,N_49638,N_46489);
nor UO_2088 (O_2088,N_46163,N_47701);
nor UO_2089 (O_2089,N_46587,N_48142);
or UO_2090 (O_2090,N_49240,N_48066);
or UO_2091 (O_2091,N_47924,N_45818);
nand UO_2092 (O_2092,N_49418,N_46201);
nor UO_2093 (O_2093,N_48410,N_49790);
and UO_2094 (O_2094,N_47504,N_48982);
or UO_2095 (O_2095,N_49853,N_49717);
nor UO_2096 (O_2096,N_47612,N_45620);
nand UO_2097 (O_2097,N_47582,N_49486);
xor UO_2098 (O_2098,N_49930,N_46477);
nor UO_2099 (O_2099,N_46023,N_48685);
nand UO_2100 (O_2100,N_47940,N_45601);
and UO_2101 (O_2101,N_47343,N_48860);
xnor UO_2102 (O_2102,N_48905,N_47520);
nor UO_2103 (O_2103,N_49028,N_47235);
xnor UO_2104 (O_2104,N_48256,N_48222);
xnor UO_2105 (O_2105,N_47606,N_47036);
or UO_2106 (O_2106,N_45470,N_45311);
xnor UO_2107 (O_2107,N_49959,N_47091);
xnor UO_2108 (O_2108,N_46318,N_49353);
xor UO_2109 (O_2109,N_47193,N_49431);
and UO_2110 (O_2110,N_45465,N_49793);
nor UO_2111 (O_2111,N_47506,N_46529);
or UO_2112 (O_2112,N_48619,N_48437);
nor UO_2113 (O_2113,N_48314,N_45609);
or UO_2114 (O_2114,N_49700,N_45839);
nor UO_2115 (O_2115,N_48349,N_45091);
xnor UO_2116 (O_2116,N_49396,N_47554);
nor UO_2117 (O_2117,N_49876,N_46823);
nor UO_2118 (O_2118,N_45539,N_49149);
or UO_2119 (O_2119,N_49372,N_48031);
nor UO_2120 (O_2120,N_46286,N_49500);
and UO_2121 (O_2121,N_46851,N_49219);
xnor UO_2122 (O_2122,N_46212,N_46138);
nor UO_2123 (O_2123,N_45412,N_49991);
and UO_2124 (O_2124,N_47371,N_47523);
or UO_2125 (O_2125,N_48835,N_45892);
xor UO_2126 (O_2126,N_47025,N_46148);
or UO_2127 (O_2127,N_48650,N_49357);
and UO_2128 (O_2128,N_47367,N_46124);
nand UO_2129 (O_2129,N_46340,N_49111);
nand UO_2130 (O_2130,N_46328,N_48600);
nand UO_2131 (O_2131,N_46781,N_48072);
or UO_2132 (O_2132,N_49935,N_47369);
and UO_2133 (O_2133,N_49738,N_49087);
xnor UO_2134 (O_2134,N_48415,N_47870);
nor UO_2135 (O_2135,N_45530,N_48716);
and UO_2136 (O_2136,N_49654,N_47786);
or UO_2137 (O_2137,N_46175,N_45401);
xnor UO_2138 (O_2138,N_47844,N_48751);
nor UO_2139 (O_2139,N_46633,N_47119);
nor UO_2140 (O_2140,N_49061,N_48746);
xor UO_2141 (O_2141,N_49474,N_47350);
or UO_2142 (O_2142,N_47102,N_46469);
or UO_2143 (O_2143,N_48597,N_48708);
xor UO_2144 (O_2144,N_47216,N_47503);
nand UO_2145 (O_2145,N_48812,N_48059);
xnor UO_2146 (O_2146,N_49248,N_46259);
nand UO_2147 (O_2147,N_45910,N_49570);
nor UO_2148 (O_2148,N_45479,N_45026);
and UO_2149 (O_2149,N_49197,N_45865);
nand UO_2150 (O_2150,N_48998,N_45140);
xor UO_2151 (O_2151,N_49560,N_48926);
nor UO_2152 (O_2152,N_45946,N_45736);
nor UO_2153 (O_2153,N_48846,N_47812);
xor UO_2154 (O_2154,N_49492,N_46636);
nand UO_2155 (O_2155,N_46775,N_49553);
or UO_2156 (O_2156,N_48726,N_46059);
and UO_2157 (O_2157,N_47218,N_48309);
nand UO_2158 (O_2158,N_47725,N_48044);
nor UO_2159 (O_2159,N_48789,N_46575);
nor UO_2160 (O_2160,N_49882,N_45067);
and UO_2161 (O_2161,N_48174,N_45637);
or UO_2162 (O_2162,N_47641,N_45693);
xnor UO_2163 (O_2163,N_46651,N_45426);
xor UO_2164 (O_2164,N_49221,N_45879);
or UO_2165 (O_2165,N_47677,N_45830);
and UO_2166 (O_2166,N_45944,N_46066);
xor UO_2167 (O_2167,N_46986,N_47699);
xnor UO_2168 (O_2168,N_47319,N_49164);
and UO_2169 (O_2169,N_47933,N_48772);
nand UO_2170 (O_2170,N_47637,N_49133);
or UO_2171 (O_2171,N_46616,N_48774);
xor UO_2172 (O_2172,N_46470,N_46863);
and UO_2173 (O_2173,N_48656,N_46678);
and UO_2174 (O_2174,N_47393,N_48941);
nand UO_2175 (O_2175,N_46345,N_45888);
nor UO_2176 (O_2176,N_47735,N_48563);
nor UO_2177 (O_2177,N_46010,N_46807);
xnor UO_2178 (O_2178,N_46001,N_48828);
or UO_2179 (O_2179,N_47627,N_48691);
nor UO_2180 (O_2180,N_49851,N_45095);
nor UO_2181 (O_2181,N_49002,N_45472);
nand UO_2182 (O_2182,N_47067,N_49766);
nand UO_2183 (O_2183,N_45006,N_46502);
xor UO_2184 (O_2184,N_45551,N_45357);
nand UO_2185 (O_2185,N_46635,N_45851);
nor UO_2186 (O_2186,N_45399,N_47642);
xnor UO_2187 (O_2187,N_48137,N_47076);
xnor UO_2188 (O_2188,N_45062,N_46805);
xnor UO_2189 (O_2189,N_49682,N_49836);
nand UO_2190 (O_2190,N_47809,N_48684);
or UO_2191 (O_2191,N_46992,N_45638);
xor UO_2192 (O_2192,N_46005,N_45899);
or UO_2193 (O_2193,N_46156,N_45683);
xor UO_2194 (O_2194,N_45984,N_45413);
nand UO_2195 (O_2195,N_46171,N_49830);
or UO_2196 (O_2196,N_45569,N_49828);
xor UO_2197 (O_2197,N_49911,N_49554);
and UO_2198 (O_2198,N_45916,N_46220);
nand UO_2199 (O_2199,N_48399,N_47304);
or UO_2200 (O_2200,N_46429,N_47826);
nor UO_2201 (O_2201,N_47413,N_48127);
and UO_2202 (O_2202,N_48170,N_47195);
nor UO_2203 (O_2203,N_48813,N_45557);
nand UO_2204 (O_2204,N_47339,N_49308);
or UO_2205 (O_2205,N_49691,N_49713);
nor UO_2206 (O_2206,N_49348,N_48335);
and UO_2207 (O_2207,N_46652,N_45516);
and UO_2208 (O_2208,N_48851,N_47484);
nor UO_2209 (O_2209,N_45969,N_48136);
or UO_2210 (O_2210,N_47289,N_49984);
or UO_2211 (O_2211,N_49538,N_45476);
xor UO_2212 (O_2212,N_45561,N_48339);
nand UO_2213 (O_2213,N_46446,N_45010);
or UO_2214 (O_2214,N_49615,N_48786);
nor UO_2215 (O_2215,N_46999,N_47489);
nor UO_2216 (O_2216,N_46397,N_47658);
xnor UO_2217 (O_2217,N_46463,N_47284);
nor UO_2218 (O_2218,N_48258,N_48599);
xnor UO_2219 (O_2219,N_46496,N_45136);
nand UO_2220 (O_2220,N_49624,N_45871);
xor UO_2221 (O_2221,N_45271,N_47059);
nor UO_2222 (O_2222,N_48340,N_45017);
and UO_2223 (O_2223,N_48372,N_46289);
and UO_2224 (O_2224,N_45791,N_49429);
nor UO_2225 (O_2225,N_46514,N_48050);
or UO_2226 (O_2226,N_49875,N_45856);
and UO_2227 (O_2227,N_45276,N_49517);
nand UO_2228 (O_2228,N_45709,N_48791);
or UO_2229 (O_2229,N_49917,N_45368);
nor UO_2230 (O_2230,N_47711,N_47017);
xor UO_2231 (O_2231,N_47061,N_49870);
or UO_2232 (O_2232,N_47561,N_48581);
or UO_2233 (O_2233,N_46453,N_48251);
or UO_2234 (O_2234,N_49666,N_49192);
and UO_2235 (O_2235,N_48411,N_47481);
nor UO_2236 (O_2236,N_47982,N_46721);
nor UO_2237 (O_2237,N_46577,N_49493);
nand UO_2238 (O_2238,N_47689,N_47322);
nand UO_2239 (O_2239,N_47685,N_45996);
nand UO_2240 (O_2240,N_48647,N_47763);
or UO_2241 (O_2241,N_49013,N_49305);
or UO_2242 (O_2242,N_46078,N_45106);
or UO_2243 (O_2243,N_46760,N_48997);
and UO_2244 (O_2244,N_48311,N_45880);
nand UO_2245 (O_2245,N_46033,N_47008);
and UO_2246 (O_2246,N_49798,N_47882);
nor UO_2247 (O_2247,N_48661,N_47070);
nand UO_2248 (O_2248,N_49033,N_48857);
xnor UO_2249 (O_2249,N_49228,N_46395);
nand UO_2250 (O_2250,N_48181,N_47756);
nand UO_2251 (O_2251,N_45868,N_48228);
nor UO_2252 (O_2252,N_45590,N_45011);
and UO_2253 (O_2253,N_45572,N_48983);
nor UO_2254 (O_2254,N_45978,N_49319);
nand UO_2255 (O_2255,N_47667,N_46751);
nor UO_2256 (O_2256,N_46910,N_48058);
and UO_2257 (O_2257,N_46342,N_49739);
xor UO_2258 (O_2258,N_45679,N_49787);
or UO_2259 (O_2259,N_47707,N_46866);
xnor UO_2260 (O_2260,N_45684,N_48138);
xnor UO_2261 (O_2261,N_46266,N_48115);
nand UO_2262 (O_2262,N_45861,N_49012);
xor UO_2263 (O_2263,N_49067,N_49702);
nor UO_2264 (O_2264,N_49628,N_45259);
nand UO_2265 (O_2265,N_49603,N_47811);
and UO_2266 (O_2266,N_46755,N_48744);
nor UO_2267 (O_2267,N_46690,N_45864);
nor UO_2268 (O_2268,N_48273,N_49483);
nor UO_2269 (O_2269,N_46449,N_48304);
nor UO_2270 (O_2270,N_46089,N_46293);
and UO_2271 (O_2271,N_46562,N_46625);
xnor UO_2272 (O_2272,N_49101,N_48973);
xor UO_2273 (O_2273,N_45292,N_46601);
or UO_2274 (O_2274,N_47602,N_49204);
nand UO_2275 (O_2275,N_49458,N_45938);
xnor UO_2276 (O_2276,N_49090,N_46441);
nor UO_2277 (O_2277,N_48295,N_45385);
xor UO_2278 (O_2278,N_45580,N_47372);
nand UO_2279 (O_2279,N_47598,N_48178);
nor UO_2280 (O_2280,N_48047,N_45203);
nor UO_2281 (O_2281,N_49085,N_49272);
or UO_2282 (O_2282,N_46894,N_48229);
or UO_2283 (O_2283,N_45737,N_47253);
nand UO_2284 (O_2284,N_45974,N_47463);
nor UO_2285 (O_2285,N_46824,N_49210);
nor UO_2286 (O_2286,N_49779,N_45940);
nor UO_2287 (O_2287,N_47681,N_47058);
and UO_2288 (O_2288,N_48027,N_48761);
nor UO_2289 (O_2289,N_47662,N_45877);
xor UO_2290 (O_2290,N_47080,N_47292);
xnor UO_2291 (O_2291,N_45822,N_45630);
or UO_2292 (O_2292,N_47749,N_45543);
and UO_2293 (O_2293,N_46884,N_45747);
and UO_2294 (O_2294,N_49387,N_47784);
nand UO_2295 (O_2295,N_47668,N_46334);
xor UO_2296 (O_2296,N_47386,N_49313);
or UO_2297 (O_2297,N_47028,N_49675);
or UO_2298 (O_2298,N_47254,N_46891);
and UO_2299 (O_2299,N_45662,N_46595);
nor UO_2300 (O_2300,N_48556,N_47970);
xnor UO_2301 (O_2301,N_46848,N_49042);
or UO_2302 (O_2302,N_48890,N_48016);
nand UO_2303 (O_2303,N_49979,N_46257);
xor UO_2304 (O_2304,N_48430,N_47280);
xnor UO_2305 (O_2305,N_49009,N_49237);
xnor UO_2306 (O_2306,N_46668,N_47204);
nand UO_2307 (O_2307,N_48081,N_49096);
xnor UO_2308 (O_2308,N_47110,N_48990);
and UO_2309 (O_2309,N_47163,N_45436);
nor UO_2310 (O_2310,N_47334,N_47019);
nor UO_2311 (O_2311,N_49909,N_46709);
nand UO_2312 (O_2312,N_49887,N_48785);
xnor UO_2313 (O_2313,N_48320,N_45054);
nor UO_2314 (O_2314,N_49155,N_47451);
nand UO_2315 (O_2315,N_48089,N_48703);
nand UO_2316 (O_2316,N_48482,N_46797);
and UO_2317 (O_2317,N_45487,N_46895);
or UO_2318 (O_2318,N_46307,N_48715);
or UO_2319 (O_2319,N_45725,N_46480);
and UO_2320 (O_2320,N_48534,N_47169);
xor UO_2321 (O_2321,N_49083,N_46113);
xor UO_2322 (O_2322,N_48425,N_49812);
nand UO_2323 (O_2323,N_45905,N_45163);
xnor UO_2324 (O_2324,N_46095,N_49816);
or UO_2325 (O_2325,N_47404,N_45503);
nor UO_2326 (O_2326,N_46170,N_47246);
xor UO_2327 (O_2327,N_48344,N_48124);
or UO_2328 (O_2328,N_45356,N_45841);
nand UO_2329 (O_2329,N_46060,N_46784);
and UO_2330 (O_2330,N_46211,N_49845);
and UO_2331 (O_2331,N_45941,N_48681);
xnor UO_2332 (O_2332,N_49250,N_47848);
xnor UO_2333 (O_2333,N_45863,N_48934);
or UO_2334 (O_2334,N_48721,N_49649);
xnor UO_2335 (O_2335,N_45727,N_47173);
or UO_2336 (O_2336,N_49055,N_46209);
or UO_2337 (O_2337,N_48872,N_46297);
nand UO_2338 (O_2338,N_49160,N_49212);
nor UO_2339 (O_2339,N_45007,N_48233);
nor UO_2340 (O_2340,N_48486,N_45845);
xor UO_2341 (O_2341,N_48895,N_46925);
nor UO_2342 (O_2342,N_49185,N_48921);
nor UO_2343 (O_2343,N_47652,N_47444);
or UO_2344 (O_2344,N_46034,N_46487);
nor UO_2345 (O_2345,N_46516,N_46322);
xor UO_2346 (O_2346,N_49163,N_46850);
or UO_2347 (O_2347,N_46147,N_49235);
or UO_2348 (O_2348,N_45188,N_47938);
or UO_2349 (O_2349,N_49473,N_47274);
or UO_2350 (O_2350,N_45780,N_45262);
nor UO_2351 (O_2351,N_48525,N_49351);
xnor UO_2352 (O_2352,N_47660,N_47130);
nor UO_2353 (O_2353,N_47057,N_47438);
nor UO_2354 (O_2354,N_46623,N_48623);
and UO_2355 (O_2355,N_45269,N_45792);
nand UO_2356 (O_2356,N_45182,N_46893);
nor UO_2357 (O_2357,N_46970,N_46662);
and UO_2358 (O_2358,N_46820,N_47294);
or UO_2359 (O_2359,N_46115,N_46531);
xnor UO_2360 (O_2360,N_48337,N_49077);
xor UO_2361 (O_2361,N_48839,N_46088);
and UO_2362 (O_2362,N_49992,N_47776);
or UO_2363 (O_2363,N_47191,N_49531);
or UO_2364 (O_2364,N_49068,N_49890);
nor UO_2365 (O_2365,N_45819,N_48861);
or UO_2366 (O_2366,N_45800,N_48958);
nand UO_2367 (O_2367,N_47698,N_46922);
and UO_2368 (O_2368,N_46557,N_49931);
nor UO_2369 (O_2369,N_48594,N_47958);
and UO_2370 (O_2370,N_49376,N_47495);
nor UO_2371 (O_2371,N_47771,N_47331);
nand UO_2372 (O_2372,N_48732,N_45632);
nand UO_2373 (O_2373,N_49242,N_45575);
nand UO_2374 (O_2374,N_49948,N_49497);
xor UO_2375 (O_2375,N_48063,N_46294);
nand UO_2376 (O_2376,N_46821,N_49218);
nand UO_2377 (O_2377,N_49971,N_48818);
nand UO_2378 (O_2378,N_45790,N_49049);
xor UO_2379 (O_2379,N_49993,N_45933);
xnor UO_2380 (O_2380,N_49535,N_47807);
and UO_2381 (O_2381,N_45396,N_45427);
and UO_2382 (O_2382,N_49696,N_49891);
or UO_2383 (O_2383,N_45778,N_47442);
nand UO_2384 (O_2384,N_45031,N_49540);
and UO_2385 (O_2385,N_47744,N_45593);
or UO_2386 (O_2386,N_47247,N_48764);
nand UO_2387 (O_2387,N_48013,N_45416);
nor UO_2388 (O_2388,N_49913,N_47998);
nand UO_2389 (O_2389,N_47697,N_48981);
nor UO_2390 (O_2390,N_47887,N_49467);
and UO_2391 (O_2391,N_48163,N_48009);
nor UO_2392 (O_2392,N_48404,N_46051);
xnor UO_2393 (O_2393,N_46443,N_49293);
or UO_2394 (O_2394,N_46965,N_45379);
nand UO_2395 (O_2395,N_49239,N_48132);
xnor UO_2396 (O_2396,N_49424,N_45456);
xnor UO_2397 (O_2397,N_45250,N_45810);
nand UO_2398 (O_2398,N_46384,N_48083);
nor UO_2399 (O_2399,N_49586,N_48831);
xor UO_2400 (O_2400,N_48837,N_45278);
or UO_2401 (O_2401,N_48692,N_49942);
and UO_2402 (O_2402,N_49711,N_46933);
nor UO_2403 (O_2403,N_48494,N_48815);
nor UO_2404 (O_2404,N_49165,N_45346);
and UO_2405 (O_2405,N_47513,N_47009);
or UO_2406 (O_2406,N_48455,N_49315);
nor UO_2407 (O_2407,N_48395,N_47464);
xnor UO_2408 (O_2408,N_48883,N_45312);
or UO_2409 (O_2409,N_46194,N_48422);
nor UO_2410 (O_2410,N_48520,N_47581);
nand UO_2411 (O_2411,N_47571,N_46376);
nor UO_2412 (O_2412,N_47775,N_48568);
nand UO_2413 (O_2413,N_49690,N_49660);
xor UO_2414 (O_2414,N_47603,N_46046);
xnor UO_2415 (O_2415,N_48634,N_47252);
nand UO_2416 (O_2416,N_45158,N_49430);
and UO_2417 (O_2417,N_47021,N_46464);
nor UO_2418 (O_2418,N_46016,N_48505);
xnor UO_2419 (O_2419,N_46696,N_45317);
nor UO_2420 (O_2420,N_49686,N_48917);
and UO_2421 (O_2421,N_45731,N_45701);
nor UO_2422 (O_2422,N_49542,N_46251);
and UO_2423 (O_2423,N_45214,N_48887);
xor UO_2424 (O_2424,N_49974,N_46285);
nor UO_2425 (O_2425,N_45410,N_49767);
nand UO_2426 (O_2426,N_45181,N_49549);
nand UO_2427 (O_2427,N_48693,N_46358);
nor UO_2428 (O_2428,N_49130,N_45525);
and UO_2429 (O_2429,N_45823,N_46459);
and UO_2430 (O_2430,N_49306,N_48626);
or UO_2431 (O_2431,N_46506,N_49462);
nand UO_2432 (O_2432,N_46610,N_49190);
xnor UO_2433 (O_2433,N_48354,N_46490);
xor UO_2434 (O_2434,N_49076,N_47544);
nand UO_2435 (O_2435,N_48959,N_48663);
and UO_2436 (O_2436,N_45663,N_49676);
nand UO_2437 (O_2437,N_48291,N_48007);
and UO_2438 (O_2438,N_46969,N_45752);
xor UO_2439 (O_2439,N_49018,N_47556);
or UO_2440 (O_2440,N_49217,N_46772);
nand UO_2441 (O_2441,N_49181,N_47512);
nand UO_2442 (O_2442,N_46149,N_45215);
and UO_2443 (O_2443,N_49536,N_46032);
nand UO_2444 (O_2444,N_46121,N_49324);
nor UO_2445 (O_2445,N_46806,N_49927);
nor UO_2446 (O_2446,N_46640,N_49827);
xor UO_2447 (O_2447,N_49736,N_46974);
and UO_2448 (O_2448,N_46383,N_49981);
nand UO_2449 (O_2449,N_48528,N_45878);
nor UO_2450 (O_2450,N_47537,N_48355);
xnor UO_2451 (O_2451,N_46688,N_47298);
nand UO_2452 (O_2452,N_48621,N_49525);
and UO_2453 (O_2453,N_49326,N_47231);
nand UO_2454 (O_2454,N_48796,N_46552);
nand UO_2455 (O_2455,N_47267,N_46738);
or UO_2456 (O_2456,N_47898,N_45805);
xnor UO_2457 (O_2457,N_49017,N_47653);
or UO_2458 (O_2458,N_49567,N_49172);
nand UO_2459 (O_2459,N_46906,N_48153);
nand UO_2460 (O_2460,N_45114,N_45350);
and UO_2461 (O_2461,N_49962,N_45425);
and UO_2462 (O_2462,N_49496,N_46330);
or UO_2463 (O_2463,N_47676,N_46810);
nand UO_2464 (O_2464,N_47654,N_46132);
and UO_2465 (O_2465,N_49822,N_49304);
or UO_2466 (O_2466,N_48398,N_49633);
nand UO_2467 (O_2467,N_45324,N_48843);
xnor UO_2468 (O_2468,N_47560,N_49834);
and UO_2469 (O_2469,N_47233,N_47738);
or UO_2470 (O_2470,N_47594,N_48283);
nor UO_2471 (O_2471,N_45441,N_47208);
or UO_2472 (O_2472,N_48900,N_49238);
xnor UO_2473 (O_2473,N_49209,N_47878);
or UO_2474 (O_2474,N_46897,N_49299);
or UO_2475 (O_2475,N_46841,N_46953);
and UO_2476 (O_2476,N_45019,N_47546);
or UO_2477 (O_2477,N_48593,N_46761);
and UO_2478 (O_2478,N_48798,N_49412);
xnor UO_2479 (O_2479,N_47104,N_48208);
xnor UO_2480 (O_2480,N_47423,N_48202);
or UO_2481 (O_2481,N_47157,N_48836);
nor UO_2482 (O_2482,N_45273,N_49399);
xnor UO_2483 (O_2483,N_47792,N_45993);
nand UO_2484 (O_2484,N_46710,N_46618);
nand UO_2485 (O_2485,N_49596,N_48725);
or UO_2486 (O_2486,N_48671,N_48561);
or UO_2487 (O_2487,N_48257,N_47270);
nand UO_2488 (O_2488,N_47320,N_48618);
nand UO_2489 (O_2489,N_45488,N_49001);
nand UO_2490 (O_2490,N_45817,N_46720);
nand UO_2491 (O_2491,N_47562,N_46153);
and UO_2492 (O_2492,N_48977,N_49045);
or UO_2493 (O_2493,N_47441,N_47242);
and UO_2494 (O_2494,N_49754,N_46885);
nor UO_2495 (O_2495,N_45034,N_48755);
nor UO_2496 (O_2496,N_49678,N_45248);
and UO_2497 (O_2497,N_47085,N_47168);
xnor UO_2498 (O_2498,N_48234,N_46794);
or UO_2499 (O_2499,N_48875,N_48280);
xor UO_2500 (O_2500,N_47900,N_47878);
nand UO_2501 (O_2501,N_46437,N_47753);
nor UO_2502 (O_2502,N_49466,N_49959);
nand UO_2503 (O_2503,N_49117,N_47320);
nand UO_2504 (O_2504,N_45739,N_49831);
and UO_2505 (O_2505,N_49706,N_48302);
or UO_2506 (O_2506,N_49615,N_46447);
or UO_2507 (O_2507,N_48055,N_48991);
xor UO_2508 (O_2508,N_49145,N_49118);
xor UO_2509 (O_2509,N_48833,N_47917);
and UO_2510 (O_2510,N_48457,N_46303);
nand UO_2511 (O_2511,N_48820,N_47438);
or UO_2512 (O_2512,N_49923,N_47140);
nand UO_2513 (O_2513,N_45555,N_48009);
or UO_2514 (O_2514,N_48929,N_47520);
or UO_2515 (O_2515,N_47500,N_49810);
xor UO_2516 (O_2516,N_48338,N_46614);
xnor UO_2517 (O_2517,N_45629,N_49240);
or UO_2518 (O_2518,N_48533,N_46583);
nand UO_2519 (O_2519,N_45340,N_46883);
xor UO_2520 (O_2520,N_46639,N_48883);
and UO_2521 (O_2521,N_49608,N_47441);
or UO_2522 (O_2522,N_49766,N_47751);
nor UO_2523 (O_2523,N_49281,N_48775);
or UO_2524 (O_2524,N_49196,N_47995);
nand UO_2525 (O_2525,N_47853,N_45135);
nand UO_2526 (O_2526,N_45541,N_46851);
or UO_2527 (O_2527,N_47027,N_48805);
nand UO_2528 (O_2528,N_47111,N_47948);
nor UO_2529 (O_2529,N_46786,N_45687);
and UO_2530 (O_2530,N_49076,N_48681);
nor UO_2531 (O_2531,N_46550,N_47378);
nor UO_2532 (O_2532,N_49926,N_46817);
xor UO_2533 (O_2533,N_46824,N_46198);
or UO_2534 (O_2534,N_48589,N_46340);
xnor UO_2535 (O_2535,N_46703,N_48797);
nand UO_2536 (O_2536,N_46259,N_48749);
or UO_2537 (O_2537,N_45606,N_45229);
nor UO_2538 (O_2538,N_46891,N_45072);
and UO_2539 (O_2539,N_46972,N_48792);
or UO_2540 (O_2540,N_47055,N_45493);
xnor UO_2541 (O_2541,N_45882,N_46325);
nor UO_2542 (O_2542,N_46926,N_48075);
nand UO_2543 (O_2543,N_46551,N_45493);
and UO_2544 (O_2544,N_45630,N_49105);
and UO_2545 (O_2545,N_48021,N_47689);
nand UO_2546 (O_2546,N_48311,N_46914);
nor UO_2547 (O_2547,N_46400,N_46599);
xor UO_2548 (O_2548,N_45345,N_49393);
nor UO_2549 (O_2549,N_45148,N_47191);
and UO_2550 (O_2550,N_49686,N_45257);
nand UO_2551 (O_2551,N_46301,N_48908);
nor UO_2552 (O_2552,N_48124,N_48645);
and UO_2553 (O_2553,N_48758,N_48363);
xor UO_2554 (O_2554,N_46516,N_47876);
nand UO_2555 (O_2555,N_46895,N_45832);
and UO_2556 (O_2556,N_46498,N_49012);
nand UO_2557 (O_2557,N_49541,N_46291);
xor UO_2558 (O_2558,N_48277,N_45648);
xor UO_2559 (O_2559,N_46676,N_46612);
xor UO_2560 (O_2560,N_45542,N_46251);
nor UO_2561 (O_2561,N_49357,N_49308);
nor UO_2562 (O_2562,N_49186,N_48799);
or UO_2563 (O_2563,N_47419,N_47423);
nand UO_2564 (O_2564,N_47404,N_48905);
nand UO_2565 (O_2565,N_48807,N_47358);
xnor UO_2566 (O_2566,N_48560,N_49651);
xor UO_2567 (O_2567,N_47743,N_45154);
nor UO_2568 (O_2568,N_45072,N_45609);
xor UO_2569 (O_2569,N_48425,N_47945);
nor UO_2570 (O_2570,N_49724,N_46446);
nand UO_2571 (O_2571,N_49587,N_48258);
or UO_2572 (O_2572,N_45840,N_48401);
nand UO_2573 (O_2573,N_48457,N_48199);
or UO_2574 (O_2574,N_47265,N_47301);
nand UO_2575 (O_2575,N_45599,N_48805);
nand UO_2576 (O_2576,N_49666,N_49802);
nand UO_2577 (O_2577,N_49911,N_47943);
xor UO_2578 (O_2578,N_47076,N_45673);
nand UO_2579 (O_2579,N_46258,N_47609);
nor UO_2580 (O_2580,N_48816,N_49452);
or UO_2581 (O_2581,N_49776,N_49214);
xor UO_2582 (O_2582,N_46204,N_47991);
and UO_2583 (O_2583,N_46269,N_45609);
nand UO_2584 (O_2584,N_48129,N_45973);
or UO_2585 (O_2585,N_45546,N_45371);
xor UO_2586 (O_2586,N_47981,N_49735);
and UO_2587 (O_2587,N_49471,N_47028);
or UO_2588 (O_2588,N_45585,N_46655);
xor UO_2589 (O_2589,N_45070,N_48416);
nor UO_2590 (O_2590,N_48012,N_49556);
xor UO_2591 (O_2591,N_49200,N_48388);
and UO_2592 (O_2592,N_46496,N_46346);
nor UO_2593 (O_2593,N_47085,N_48312);
nand UO_2594 (O_2594,N_49457,N_46619);
xor UO_2595 (O_2595,N_47558,N_49204);
nor UO_2596 (O_2596,N_49749,N_49917);
nor UO_2597 (O_2597,N_46102,N_46299);
and UO_2598 (O_2598,N_49202,N_49506);
nor UO_2599 (O_2599,N_45505,N_49781);
nand UO_2600 (O_2600,N_46081,N_49431);
and UO_2601 (O_2601,N_49657,N_47589);
nand UO_2602 (O_2602,N_48239,N_45671);
nand UO_2603 (O_2603,N_46683,N_48961);
nor UO_2604 (O_2604,N_49241,N_47577);
nand UO_2605 (O_2605,N_48435,N_47972);
and UO_2606 (O_2606,N_49936,N_45274);
xnor UO_2607 (O_2607,N_48403,N_49450);
nor UO_2608 (O_2608,N_46640,N_49368);
or UO_2609 (O_2609,N_49156,N_48196);
nand UO_2610 (O_2610,N_46518,N_48164);
and UO_2611 (O_2611,N_47849,N_47486);
and UO_2612 (O_2612,N_47189,N_49813);
nand UO_2613 (O_2613,N_47390,N_46845);
or UO_2614 (O_2614,N_47778,N_48467);
nor UO_2615 (O_2615,N_49262,N_45345);
nand UO_2616 (O_2616,N_46229,N_47367);
nand UO_2617 (O_2617,N_45632,N_46286);
nand UO_2618 (O_2618,N_46442,N_48371);
nand UO_2619 (O_2619,N_45607,N_46353);
nor UO_2620 (O_2620,N_48713,N_46633);
nand UO_2621 (O_2621,N_46394,N_45910);
nand UO_2622 (O_2622,N_46930,N_48815);
nand UO_2623 (O_2623,N_48254,N_47063);
nand UO_2624 (O_2624,N_45126,N_47682);
xnor UO_2625 (O_2625,N_48453,N_48661);
nand UO_2626 (O_2626,N_45949,N_48494);
nand UO_2627 (O_2627,N_47468,N_45658);
xor UO_2628 (O_2628,N_49394,N_49443);
or UO_2629 (O_2629,N_47875,N_47451);
nor UO_2630 (O_2630,N_45101,N_48570);
nand UO_2631 (O_2631,N_49970,N_49401);
or UO_2632 (O_2632,N_47272,N_45860);
nand UO_2633 (O_2633,N_47996,N_46152);
nor UO_2634 (O_2634,N_45738,N_47947);
nor UO_2635 (O_2635,N_48606,N_47894);
nand UO_2636 (O_2636,N_45191,N_47663);
and UO_2637 (O_2637,N_47591,N_45089);
or UO_2638 (O_2638,N_49964,N_49646);
or UO_2639 (O_2639,N_46608,N_45199);
nor UO_2640 (O_2640,N_48451,N_47688);
nor UO_2641 (O_2641,N_47079,N_47566);
and UO_2642 (O_2642,N_47060,N_49890);
or UO_2643 (O_2643,N_46581,N_47208);
xor UO_2644 (O_2644,N_46627,N_46393);
xor UO_2645 (O_2645,N_47196,N_47320);
or UO_2646 (O_2646,N_48328,N_46731);
and UO_2647 (O_2647,N_49806,N_46834);
and UO_2648 (O_2648,N_49464,N_47123);
nand UO_2649 (O_2649,N_46049,N_46832);
nor UO_2650 (O_2650,N_46105,N_45802);
nor UO_2651 (O_2651,N_48552,N_48251);
nand UO_2652 (O_2652,N_49001,N_47804);
and UO_2653 (O_2653,N_49138,N_47645);
or UO_2654 (O_2654,N_48280,N_49056);
xnor UO_2655 (O_2655,N_47747,N_48259);
nand UO_2656 (O_2656,N_46244,N_48153);
nand UO_2657 (O_2657,N_49687,N_49544);
nand UO_2658 (O_2658,N_46919,N_45633);
and UO_2659 (O_2659,N_45548,N_48283);
or UO_2660 (O_2660,N_48796,N_49665);
and UO_2661 (O_2661,N_45840,N_45133);
nor UO_2662 (O_2662,N_46370,N_49881);
nor UO_2663 (O_2663,N_45900,N_45536);
nand UO_2664 (O_2664,N_49577,N_47172);
nand UO_2665 (O_2665,N_45690,N_47081);
nand UO_2666 (O_2666,N_45752,N_49732);
and UO_2667 (O_2667,N_48279,N_48391);
or UO_2668 (O_2668,N_48564,N_47474);
xnor UO_2669 (O_2669,N_49711,N_47653);
nand UO_2670 (O_2670,N_48423,N_49868);
or UO_2671 (O_2671,N_45698,N_49854);
xor UO_2672 (O_2672,N_48341,N_49995);
nand UO_2673 (O_2673,N_47380,N_46684);
and UO_2674 (O_2674,N_46043,N_48076);
xor UO_2675 (O_2675,N_48694,N_48318);
and UO_2676 (O_2676,N_47702,N_48566);
xnor UO_2677 (O_2677,N_45742,N_48748);
nor UO_2678 (O_2678,N_48058,N_49870);
nand UO_2679 (O_2679,N_48533,N_48902);
nand UO_2680 (O_2680,N_47260,N_47067);
and UO_2681 (O_2681,N_48789,N_46826);
nand UO_2682 (O_2682,N_49040,N_46464);
and UO_2683 (O_2683,N_49467,N_48237);
xnor UO_2684 (O_2684,N_45743,N_46139);
nand UO_2685 (O_2685,N_47005,N_47454);
nor UO_2686 (O_2686,N_49873,N_49461);
xor UO_2687 (O_2687,N_46192,N_46507);
nand UO_2688 (O_2688,N_46438,N_48937);
and UO_2689 (O_2689,N_47670,N_45947);
xnor UO_2690 (O_2690,N_45619,N_47747);
and UO_2691 (O_2691,N_48012,N_46901);
xor UO_2692 (O_2692,N_46016,N_47607);
or UO_2693 (O_2693,N_48990,N_46094);
nand UO_2694 (O_2694,N_45752,N_48489);
nor UO_2695 (O_2695,N_47045,N_48566);
nor UO_2696 (O_2696,N_45743,N_46737);
and UO_2697 (O_2697,N_46997,N_46583);
nand UO_2698 (O_2698,N_49365,N_47879);
xnor UO_2699 (O_2699,N_46930,N_49319);
xor UO_2700 (O_2700,N_45318,N_49593);
or UO_2701 (O_2701,N_47827,N_46729);
or UO_2702 (O_2702,N_48844,N_46786);
nand UO_2703 (O_2703,N_49686,N_47545);
and UO_2704 (O_2704,N_49402,N_45074);
and UO_2705 (O_2705,N_46063,N_48514);
and UO_2706 (O_2706,N_46788,N_47590);
nor UO_2707 (O_2707,N_48524,N_48026);
nor UO_2708 (O_2708,N_49067,N_47039);
nor UO_2709 (O_2709,N_47590,N_46092);
xor UO_2710 (O_2710,N_48146,N_47100);
and UO_2711 (O_2711,N_48974,N_46002);
xor UO_2712 (O_2712,N_48679,N_49135);
and UO_2713 (O_2713,N_47425,N_46561);
nand UO_2714 (O_2714,N_47361,N_47031);
nand UO_2715 (O_2715,N_49705,N_46968);
nand UO_2716 (O_2716,N_47030,N_47017);
nor UO_2717 (O_2717,N_49334,N_45458);
nor UO_2718 (O_2718,N_45220,N_47632);
or UO_2719 (O_2719,N_47758,N_46909);
or UO_2720 (O_2720,N_47103,N_48050);
xor UO_2721 (O_2721,N_47738,N_46711);
or UO_2722 (O_2722,N_47834,N_47010);
nand UO_2723 (O_2723,N_45539,N_49866);
nand UO_2724 (O_2724,N_46509,N_46023);
nor UO_2725 (O_2725,N_46823,N_49329);
nand UO_2726 (O_2726,N_45984,N_48746);
or UO_2727 (O_2727,N_48565,N_49100);
xor UO_2728 (O_2728,N_47307,N_49955);
and UO_2729 (O_2729,N_46056,N_49208);
xor UO_2730 (O_2730,N_48773,N_46405);
nor UO_2731 (O_2731,N_45815,N_45735);
or UO_2732 (O_2732,N_49232,N_46024);
nor UO_2733 (O_2733,N_49434,N_49827);
or UO_2734 (O_2734,N_46981,N_46969);
nand UO_2735 (O_2735,N_48557,N_49915);
nor UO_2736 (O_2736,N_45506,N_47829);
and UO_2737 (O_2737,N_48958,N_49660);
nand UO_2738 (O_2738,N_47430,N_45077);
nand UO_2739 (O_2739,N_47344,N_47688);
or UO_2740 (O_2740,N_48892,N_45923);
xor UO_2741 (O_2741,N_49731,N_49646);
nor UO_2742 (O_2742,N_45447,N_45361);
nand UO_2743 (O_2743,N_49550,N_45686);
xor UO_2744 (O_2744,N_47313,N_48050);
nand UO_2745 (O_2745,N_45365,N_49440);
or UO_2746 (O_2746,N_49232,N_45305);
and UO_2747 (O_2747,N_48042,N_46403);
nor UO_2748 (O_2748,N_47488,N_47001);
or UO_2749 (O_2749,N_49164,N_48098);
xor UO_2750 (O_2750,N_48639,N_45639);
nor UO_2751 (O_2751,N_49140,N_46594);
and UO_2752 (O_2752,N_49366,N_47466);
nor UO_2753 (O_2753,N_49044,N_48175);
or UO_2754 (O_2754,N_45062,N_49137);
nand UO_2755 (O_2755,N_49987,N_49642);
nand UO_2756 (O_2756,N_46065,N_48885);
nor UO_2757 (O_2757,N_46450,N_46816);
nand UO_2758 (O_2758,N_45457,N_49152);
xnor UO_2759 (O_2759,N_45707,N_45968);
and UO_2760 (O_2760,N_49880,N_46087);
nor UO_2761 (O_2761,N_46897,N_48353);
nand UO_2762 (O_2762,N_48769,N_46776);
or UO_2763 (O_2763,N_49113,N_46831);
or UO_2764 (O_2764,N_46670,N_45309);
nand UO_2765 (O_2765,N_45782,N_48973);
and UO_2766 (O_2766,N_45889,N_45454);
nand UO_2767 (O_2767,N_47182,N_47432);
xnor UO_2768 (O_2768,N_46549,N_48353);
nor UO_2769 (O_2769,N_48561,N_46196);
xor UO_2770 (O_2770,N_45987,N_47103);
xor UO_2771 (O_2771,N_48829,N_46204);
or UO_2772 (O_2772,N_49181,N_47473);
nor UO_2773 (O_2773,N_46677,N_48547);
nand UO_2774 (O_2774,N_46333,N_47762);
nor UO_2775 (O_2775,N_46891,N_46315);
nor UO_2776 (O_2776,N_46330,N_48889);
nand UO_2777 (O_2777,N_48957,N_46037);
nand UO_2778 (O_2778,N_45521,N_46905);
nor UO_2779 (O_2779,N_45544,N_46730);
nor UO_2780 (O_2780,N_49556,N_48502);
nor UO_2781 (O_2781,N_47760,N_45230);
nand UO_2782 (O_2782,N_48805,N_45484);
nand UO_2783 (O_2783,N_49272,N_45373);
and UO_2784 (O_2784,N_45425,N_49917);
or UO_2785 (O_2785,N_45237,N_45370);
nor UO_2786 (O_2786,N_48702,N_45679);
and UO_2787 (O_2787,N_46234,N_48967);
nand UO_2788 (O_2788,N_49938,N_48869);
and UO_2789 (O_2789,N_45308,N_45882);
or UO_2790 (O_2790,N_48813,N_47130);
xor UO_2791 (O_2791,N_49677,N_47272);
nand UO_2792 (O_2792,N_45777,N_48953);
and UO_2793 (O_2793,N_48871,N_46742);
or UO_2794 (O_2794,N_45924,N_45136);
nor UO_2795 (O_2795,N_45550,N_46088);
nand UO_2796 (O_2796,N_47023,N_46349);
and UO_2797 (O_2797,N_49232,N_49931);
nor UO_2798 (O_2798,N_46604,N_48492);
xnor UO_2799 (O_2799,N_45272,N_47877);
nand UO_2800 (O_2800,N_48360,N_49759);
nor UO_2801 (O_2801,N_49084,N_48994);
nand UO_2802 (O_2802,N_49574,N_45640);
nand UO_2803 (O_2803,N_45021,N_46044);
nor UO_2804 (O_2804,N_49823,N_49288);
and UO_2805 (O_2805,N_49937,N_48567);
nand UO_2806 (O_2806,N_45795,N_46924);
and UO_2807 (O_2807,N_48978,N_49185);
or UO_2808 (O_2808,N_48410,N_45362);
xnor UO_2809 (O_2809,N_46004,N_47957);
nor UO_2810 (O_2810,N_47449,N_46765);
or UO_2811 (O_2811,N_48597,N_45451);
or UO_2812 (O_2812,N_49335,N_47465);
xor UO_2813 (O_2813,N_47517,N_47800);
nor UO_2814 (O_2814,N_49298,N_48697);
nand UO_2815 (O_2815,N_47133,N_47639);
nor UO_2816 (O_2816,N_47388,N_45684);
xnor UO_2817 (O_2817,N_47585,N_49218);
xor UO_2818 (O_2818,N_45756,N_47211);
nor UO_2819 (O_2819,N_48802,N_48848);
and UO_2820 (O_2820,N_49353,N_47566);
or UO_2821 (O_2821,N_47713,N_46672);
nor UO_2822 (O_2822,N_49576,N_47638);
nor UO_2823 (O_2823,N_48515,N_46508);
and UO_2824 (O_2824,N_48276,N_49092);
xor UO_2825 (O_2825,N_46981,N_47759);
nand UO_2826 (O_2826,N_45168,N_45439);
xor UO_2827 (O_2827,N_45724,N_45068);
xor UO_2828 (O_2828,N_49875,N_49217);
and UO_2829 (O_2829,N_48130,N_47933);
and UO_2830 (O_2830,N_49675,N_49730);
and UO_2831 (O_2831,N_47154,N_48303);
and UO_2832 (O_2832,N_46739,N_46789);
nor UO_2833 (O_2833,N_49821,N_47916);
and UO_2834 (O_2834,N_45539,N_45076);
nand UO_2835 (O_2835,N_48899,N_47829);
nor UO_2836 (O_2836,N_45284,N_46790);
nand UO_2837 (O_2837,N_45276,N_49566);
nand UO_2838 (O_2838,N_49232,N_47904);
xnor UO_2839 (O_2839,N_49423,N_49236);
and UO_2840 (O_2840,N_48666,N_47870);
nor UO_2841 (O_2841,N_49829,N_49874);
and UO_2842 (O_2842,N_45446,N_49780);
or UO_2843 (O_2843,N_47368,N_47428);
nand UO_2844 (O_2844,N_48340,N_46829);
nor UO_2845 (O_2845,N_48286,N_47121);
nand UO_2846 (O_2846,N_46676,N_45021);
nand UO_2847 (O_2847,N_49084,N_49331);
and UO_2848 (O_2848,N_45807,N_47849);
nor UO_2849 (O_2849,N_45316,N_47951);
or UO_2850 (O_2850,N_45368,N_48837);
nand UO_2851 (O_2851,N_48835,N_49175);
nand UO_2852 (O_2852,N_49351,N_46156);
nand UO_2853 (O_2853,N_49287,N_49428);
nor UO_2854 (O_2854,N_47136,N_47500);
and UO_2855 (O_2855,N_45361,N_46087);
nand UO_2856 (O_2856,N_49708,N_45197);
and UO_2857 (O_2857,N_48808,N_49951);
and UO_2858 (O_2858,N_46174,N_45530);
and UO_2859 (O_2859,N_45339,N_45086);
nand UO_2860 (O_2860,N_47352,N_47894);
xor UO_2861 (O_2861,N_46534,N_47357);
nand UO_2862 (O_2862,N_45865,N_47202);
nor UO_2863 (O_2863,N_48827,N_47133);
or UO_2864 (O_2864,N_47347,N_46844);
and UO_2865 (O_2865,N_47669,N_49474);
nor UO_2866 (O_2866,N_47899,N_45479);
or UO_2867 (O_2867,N_48363,N_47509);
and UO_2868 (O_2868,N_48137,N_46243);
nand UO_2869 (O_2869,N_46367,N_47051);
or UO_2870 (O_2870,N_49822,N_48648);
xor UO_2871 (O_2871,N_45678,N_48202);
xor UO_2872 (O_2872,N_47481,N_48839);
nand UO_2873 (O_2873,N_47606,N_46676);
and UO_2874 (O_2874,N_49231,N_49505);
or UO_2875 (O_2875,N_45355,N_48537);
xor UO_2876 (O_2876,N_49500,N_46465);
nand UO_2877 (O_2877,N_48739,N_48055);
or UO_2878 (O_2878,N_49040,N_48189);
nand UO_2879 (O_2879,N_48227,N_47123);
or UO_2880 (O_2880,N_47195,N_49671);
nand UO_2881 (O_2881,N_45279,N_45068);
nor UO_2882 (O_2882,N_48937,N_49731);
nand UO_2883 (O_2883,N_49419,N_49887);
xnor UO_2884 (O_2884,N_47818,N_45573);
nor UO_2885 (O_2885,N_48213,N_48249);
nor UO_2886 (O_2886,N_48756,N_45398);
nand UO_2887 (O_2887,N_46628,N_49811);
nand UO_2888 (O_2888,N_47206,N_49576);
nand UO_2889 (O_2889,N_45368,N_46666);
nand UO_2890 (O_2890,N_45555,N_48045);
xor UO_2891 (O_2891,N_48549,N_49642);
or UO_2892 (O_2892,N_45211,N_49471);
xnor UO_2893 (O_2893,N_45824,N_45810);
and UO_2894 (O_2894,N_45623,N_45967);
nor UO_2895 (O_2895,N_46351,N_46795);
nand UO_2896 (O_2896,N_45936,N_49793);
nor UO_2897 (O_2897,N_45482,N_48114);
or UO_2898 (O_2898,N_48322,N_47739);
and UO_2899 (O_2899,N_46532,N_46339);
and UO_2900 (O_2900,N_49776,N_46682);
and UO_2901 (O_2901,N_49693,N_48797);
nand UO_2902 (O_2902,N_46222,N_45448);
nand UO_2903 (O_2903,N_45795,N_45764);
xor UO_2904 (O_2904,N_49391,N_48047);
or UO_2905 (O_2905,N_48606,N_46009);
or UO_2906 (O_2906,N_47169,N_47667);
or UO_2907 (O_2907,N_46897,N_48992);
xnor UO_2908 (O_2908,N_47407,N_47807);
or UO_2909 (O_2909,N_48669,N_49091);
or UO_2910 (O_2910,N_46033,N_46087);
nand UO_2911 (O_2911,N_46123,N_45525);
and UO_2912 (O_2912,N_48009,N_46955);
and UO_2913 (O_2913,N_48069,N_45212);
xor UO_2914 (O_2914,N_49200,N_45944);
and UO_2915 (O_2915,N_49593,N_46272);
xor UO_2916 (O_2916,N_45154,N_47399);
and UO_2917 (O_2917,N_47338,N_48680);
and UO_2918 (O_2918,N_49320,N_49012);
and UO_2919 (O_2919,N_47645,N_46735);
and UO_2920 (O_2920,N_46166,N_46822);
nand UO_2921 (O_2921,N_46804,N_47091);
and UO_2922 (O_2922,N_49419,N_49148);
and UO_2923 (O_2923,N_45161,N_45106);
nand UO_2924 (O_2924,N_46338,N_47019);
nor UO_2925 (O_2925,N_49013,N_48732);
nand UO_2926 (O_2926,N_48739,N_48037);
nor UO_2927 (O_2927,N_47863,N_49178);
nor UO_2928 (O_2928,N_45551,N_48050);
xor UO_2929 (O_2929,N_48355,N_49137);
nand UO_2930 (O_2930,N_46378,N_46304);
or UO_2931 (O_2931,N_48207,N_49746);
or UO_2932 (O_2932,N_49001,N_47532);
or UO_2933 (O_2933,N_47236,N_48233);
and UO_2934 (O_2934,N_49869,N_45133);
nor UO_2935 (O_2935,N_49942,N_48864);
xnor UO_2936 (O_2936,N_47208,N_48467);
xor UO_2937 (O_2937,N_48493,N_45239);
and UO_2938 (O_2938,N_48983,N_47613);
xor UO_2939 (O_2939,N_49438,N_48673);
nand UO_2940 (O_2940,N_47015,N_48487);
or UO_2941 (O_2941,N_49600,N_45552);
nand UO_2942 (O_2942,N_47352,N_47223);
xnor UO_2943 (O_2943,N_45644,N_48207);
nand UO_2944 (O_2944,N_45427,N_46487);
nand UO_2945 (O_2945,N_46556,N_48256);
and UO_2946 (O_2946,N_47657,N_47167);
or UO_2947 (O_2947,N_46327,N_45958);
nor UO_2948 (O_2948,N_45817,N_48330);
nor UO_2949 (O_2949,N_47880,N_46664);
or UO_2950 (O_2950,N_48757,N_49876);
nor UO_2951 (O_2951,N_45767,N_49176);
xnor UO_2952 (O_2952,N_47279,N_45829);
nor UO_2953 (O_2953,N_45986,N_49674);
nand UO_2954 (O_2954,N_45231,N_49073);
nand UO_2955 (O_2955,N_49356,N_45290);
nand UO_2956 (O_2956,N_45036,N_47875);
xor UO_2957 (O_2957,N_49236,N_49492);
nor UO_2958 (O_2958,N_49060,N_45000);
or UO_2959 (O_2959,N_46974,N_47374);
and UO_2960 (O_2960,N_49227,N_46004);
and UO_2961 (O_2961,N_48197,N_46911);
nand UO_2962 (O_2962,N_46300,N_48238);
nand UO_2963 (O_2963,N_46878,N_45043);
xor UO_2964 (O_2964,N_49209,N_49681);
and UO_2965 (O_2965,N_47065,N_46766);
xor UO_2966 (O_2966,N_47067,N_49041);
or UO_2967 (O_2967,N_45264,N_48119);
or UO_2968 (O_2968,N_48249,N_48351);
or UO_2969 (O_2969,N_48673,N_45107);
nand UO_2970 (O_2970,N_47305,N_45645);
nor UO_2971 (O_2971,N_46538,N_45768);
or UO_2972 (O_2972,N_49495,N_48811);
nand UO_2973 (O_2973,N_47385,N_45954);
nor UO_2974 (O_2974,N_49519,N_46676);
or UO_2975 (O_2975,N_46422,N_48135);
xor UO_2976 (O_2976,N_49529,N_49308);
xor UO_2977 (O_2977,N_47441,N_45550);
xnor UO_2978 (O_2978,N_47384,N_46385);
nand UO_2979 (O_2979,N_48486,N_46749);
or UO_2980 (O_2980,N_49705,N_45082);
nor UO_2981 (O_2981,N_49527,N_46791);
xnor UO_2982 (O_2982,N_48503,N_45157);
nand UO_2983 (O_2983,N_45475,N_46177);
and UO_2984 (O_2984,N_48833,N_47324);
nand UO_2985 (O_2985,N_47495,N_49649);
or UO_2986 (O_2986,N_46212,N_49818);
or UO_2987 (O_2987,N_47927,N_46366);
or UO_2988 (O_2988,N_47253,N_48945);
nor UO_2989 (O_2989,N_47924,N_48748);
nand UO_2990 (O_2990,N_46966,N_46344);
nand UO_2991 (O_2991,N_45196,N_45347);
nor UO_2992 (O_2992,N_46517,N_49039);
nor UO_2993 (O_2993,N_46547,N_48477);
or UO_2994 (O_2994,N_46648,N_47600);
nor UO_2995 (O_2995,N_49606,N_46076);
xor UO_2996 (O_2996,N_46601,N_48406);
xnor UO_2997 (O_2997,N_48069,N_48210);
nand UO_2998 (O_2998,N_49683,N_46024);
and UO_2999 (O_2999,N_46845,N_47570);
nor UO_3000 (O_3000,N_46025,N_49024);
xor UO_3001 (O_3001,N_48162,N_47636);
or UO_3002 (O_3002,N_46697,N_46390);
and UO_3003 (O_3003,N_45289,N_49271);
and UO_3004 (O_3004,N_48363,N_47808);
and UO_3005 (O_3005,N_47563,N_47025);
xnor UO_3006 (O_3006,N_45593,N_47623);
nand UO_3007 (O_3007,N_47752,N_48919);
xor UO_3008 (O_3008,N_45236,N_47960);
or UO_3009 (O_3009,N_49636,N_49466);
xor UO_3010 (O_3010,N_47441,N_49486);
or UO_3011 (O_3011,N_46493,N_48290);
and UO_3012 (O_3012,N_46278,N_47125);
and UO_3013 (O_3013,N_47311,N_49490);
nand UO_3014 (O_3014,N_47563,N_47880);
nand UO_3015 (O_3015,N_47714,N_47657);
and UO_3016 (O_3016,N_45418,N_46441);
nand UO_3017 (O_3017,N_49506,N_49462);
and UO_3018 (O_3018,N_47696,N_45898);
or UO_3019 (O_3019,N_45043,N_45392);
and UO_3020 (O_3020,N_45304,N_46229);
xor UO_3021 (O_3021,N_45735,N_46554);
nand UO_3022 (O_3022,N_46362,N_45816);
xnor UO_3023 (O_3023,N_46684,N_45747);
nand UO_3024 (O_3024,N_47763,N_47239);
nand UO_3025 (O_3025,N_47586,N_45693);
nand UO_3026 (O_3026,N_48087,N_48388);
or UO_3027 (O_3027,N_49290,N_46943);
xnor UO_3028 (O_3028,N_46927,N_45516);
xnor UO_3029 (O_3029,N_49926,N_45224);
nor UO_3030 (O_3030,N_47310,N_48365);
xnor UO_3031 (O_3031,N_47904,N_46080);
xor UO_3032 (O_3032,N_47765,N_45483);
xnor UO_3033 (O_3033,N_49533,N_45887);
and UO_3034 (O_3034,N_46553,N_45862);
and UO_3035 (O_3035,N_45086,N_47077);
or UO_3036 (O_3036,N_49327,N_48456);
and UO_3037 (O_3037,N_48609,N_46961);
xor UO_3038 (O_3038,N_45244,N_48355);
nand UO_3039 (O_3039,N_48194,N_48829);
or UO_3040 (O_3040,N_49667,N_49178);
nor UO_3041 (O_3041,N_49458,N_47277);
or UO_3042 (O_3042,N_49491,N_48281);
nor UO_3043 (O_3043,N_45570,N_46598);
and UO_3044 (O_3044,N_49302,N_45105);
nor UO_3045 (O_3045,N_47077,N_45787);
and UO_3046 (O_3046,N_45401,N_49495);
and UO_3047 (O_3047,N_47577,N_46065);
and UO_3048 (O_3048,N_49061,N_48236);
nor UO_3049 (O_3049,N_48904,N_46015);
nand UO_3050 (O_3050,N_47894,N_48436);
nor UO_3051 (O_3051,N_45552,N_48243);
nor UO_3052 (O_3052,N_49465,N_46863);
nor UO_3053 (O_3053,N_45433,N_47061);
nor UO_3054 (O_3054,N_47676,N_46331);
and UO_3055 (O_3055,N_48770,N_47461);
and UO_3056 (O_3056,N_47374,N_48468);
nor UO_3057 (O_3057,N_49605,N_48077);
nand UO_3058 (O_3058,N_45961,N_49374);
nand UO_3059 (O_3059,N_48374,N_45472);
or UO_3060 (O_3060,N_45333,N_48389);
nor UO_3061 (O_3061,N_49122,N_49859);
or UO_3062 (O_3062,N_46617,N_48800);
nor UO_3063 (O_3063,N_48308,N_49347);
xnor UO_3064 (O_3064,N_49574,N_47400);
nand UO_3065 (O_3065,N_48295,N_48435);
nand UO_3066 (O_3066,N_47934,N_48114);
nor UO_3067 (O_3067,N_47813,N_45804);
nand UO_3068 (O_3068,N_47041,N_45333);
or UO_3069 (O_3069,N_46529,N_47188);
and UO_3070 (O_3070,N_49474,N_45587);
nand UO_3071 (O_3071,N_49768,N_47014);
xor UO_3072 (O_3072,N_47887,N_49776);
nor UO_3073 (O_3073,N_46780,N_47254);
and UO_3074 (O_3074,N_47593,N_46541);
xnor UO_3075 (O_3075,N_47776,N_48507);
nor UO_3076 (O_3076,N_48208,N_48008);
nand UO_3077 (O_3077,N_47471,N_47948);
nor UO_3078 (O_3078,N_49759,N_45153);
nand UO_3079 (O_3079,N_46789,N_46373);
or UO_3080 (O_3080,N_48644,N_48606);
nand UO_3081 (O_3081,N_46245,N_49960);
nor UO_3082 (O_3082,N_48893,N_46402);
or UO_3083 (O_3083,N_46722,N_46903);
xnor UO_3084 (O_3084,N_49137,N_46512);
or UO_3085 (O_3085,N_48967,N_48349);
nand UO_3086 (O_3086,N_46249,N_47671);
nor UO_3087 (O_3087,N_46869,N_48640);
xnor UO_3088 (O_3088,N_46827,N_49195);
or UO_3089 (O_3089,N_48388,N_49212);
nor UO_3090 (O_3090,N_49870,N_48504);
or UO_3091 (O_3091,N_46557,N_45329);
and UO_3092 (O_3092,N_45739,N_49901);
xnor UO_3093 (O_3093,N_49374,N_48092);
xnor UO_3094 (O_3094,N_45749,N_47215);
xor UO_3095 (O_3095,N_49977,N_45394);
and UO_3096 (O_3096,N_47432,N_47662);
nand UO_3097 (O_3097,N_45271,N_47398);
xnor UO_3098 (O_3098,N_47016,N_48831);
nand UO_3099 (O_3099,N_45813,N_47387);
nor UO_3100 (O_3100,N_49254,N_47413);
xnor UO_3101 (O_3101,N_46280,N_46430);
nand UO_3102 (O_3102,N_45745,N_45137);
or UO_3103 (O_3103,N_46858,N_46031);
and UO_3104 (O_3104,N_47543,N_47105);
xor UO_3105 (O_3105,N_46525,N_45754);
nand UO_3106 (O_3106,N_48506,N_48287);
xor UO_3107 (O_3107,N_45173,N_47860);
or UO_3108 (O_3108,N_48933,N_45049);
and UO_3109 (O_3109,N_46803,N_46475);
xnor UO_3110 (O_3110,N_49488,N_48327);
and UO_3111 (O_3111,N_49465,N_48773);
nand UO_3112 (O_3112,N_47067,N_47004);
nor UO_3113 (O_3113,N_45193,N_49331);
or UO_3114 (O_3114,N_47048,N_47348);
nand UO_3115 (O_3115,N_48292,N_48786);
nor UO_3116 (O_3116,N_47724,N_48129);
nand UO_3117 (O_3117,N_49873,N_46674);
nor UO_3118 (O_3118,N_49522,N_46423);
nor UO_3119 (O_3119,N_48267,N_48922);
xor UO_3120 (O_3120,N_48844,N_47869);
or UO_3121 (O_3121,N_45047,N_47021);
nor UO_3122 (O_3122,N_46104,N_46928);
xor UO_3123 (O_3123,N_47588,N_48813);
xor UO_3124 (O_3124,N_46623,N_49438);
and UO_3125 (O_3125,N_45159,N_49762);
nor UO_3126 (O_3126,N_45874,N_45977);
xor UO_3127 (O_3127,N_46040,N_45084);
xor UO_3128 (O_3128,N_46759,N_48908);
or UO_3129 (O_3129,N_46668,N_48799);
and UO_3130 (O_3130,N_45567,N_45886);
nor UO_3131 (O_3131,N_47282,N_47186);
nand UO_3132 (O_3132,N_46754,N_46307);
nor UO_3133 (O_3133,N_45012,N_46371);
nor UO_3134 (O_3134,N_46331,N_48568);
and UO_3135 (O_3135,N_45015,N_46457);
nand UO_3136 (O_3136,N_48662,N_49570);
nor UO_3137 (O_3137,N_45608,N_49755);
and UO_3138 (O_3138,N_45807,N_47494);
xnor UO_3139 (O_3139,N_47486,N_46625);
nor UO_3140 (O_3140,N_49683,N_46788);
or UO_3141 (O_3141,N_46639,N_45897);
nand UO_3142 (O_3142,N_48550,N_46238);
and UO_3143 (O_3143,N_45281,N_49082);
xor UO_3144 (O_3144,N_48311,N_48122);
nand UO_3145 (O_3145,N_48010,N_46109);
or UO_3146 (O_3146,N_46942,N_45888);
or UO_3147 (O_3147,N_49807,N_45857);
nand UO_3148 (O_3148,N_48859,N_48105);
xor UO_3149 (O_3149,N_49069,N_46617);
nor UO_3150 (O_3150,N_45921,N_47692);
and UO_3151 (O_3151,N_46923,N_45312);
nor UO_3152 (O_3152,N_48892,N_49339);
xor UO_3153 (O_3153,N_46255,N_46840);
xor UO_3154 (O_3154,N_49348,N_49905);
or UO_3155 (O_3155,N_48363,N_49695);
nor UO_3156 (O_3156,N_45006,N_48717);
and UO_3157 (O_3157,N_45313,N_46334);
xnor UO_3158 (O_3158,N_45212,N_47066);
nor UO_3159 (O_3159,N_49212,N_49190);
or UO_3160 (O_3160,N_48279,N_49341);
and UO_3161 (O_3161,N_49209,N_47141);
nor UO_3162 (O_3162,N_46026,N_45905);
xor UO_3163 (O_3163,N_48678,N_48085);
or UO_3164 (O_3164,N_47315,N_48266);
nor UO_3165 (O_3165,N_47162,N_47212);
or UO_3166 (O_3166,N_48564,N_49752);
xor UO_3167 (O_3167,N_49943,N_45147);
nor UO_3168 (O_3168,N_47910,N_48264);
nor UO_3169 (O_3169,N_48835,N_47760);
or UO_3170 (O_3170,N_46770,N_46374);
nand UO_3171 (O_3171,N_48456,N_48400);
or UO_3172 (O_3172,N_47937,N_48805);
nor UO_3173 (O_3173,N_49032,N_48520);
nor UO_3174 (O_3174,N_47110,N_46220);
nand UO_3175 (O_3175,N_45555,N_45863);
and UO_3176 (O_3176,N_45445,N_45741);
and UO_3177 (O_3177,N_47940,N_47895);
or UO_3178 (O_3178,N_46739,N_48284);
and UO_3179 (O_3179,N_47335,N_46884);
nor UO_3180 (O_3180,N_49288,N_45614);
xor UO_3181 (O_3181,N_45723,N_49439);
and UO_3182 (O_3182,N_48400,N_49734);
nor UO_3183 (O_3183,N_49034,N_49498);
or UO_3184 (O_3184,N_45035,N_48320);
or UO_3185 (O_3185,N_47287,N_46605);
nor UO_3186 (O_3186,N_48333,N_45942);
and UO_3187 (O_3187,N_45300,N_46441);
nor UO_3188 (O_3188,N_46091,N_48985);
xor UO_3189 (O_3189,N_46998,N_48476);
and UO_3190 (O_3190,N_46026,N_47500);
nor UO_3191 (O_3191,N_47542,N_49922);
xor UO_3192 (O_3192,N_48007,N_46913);
xnor UO_3193 (O_3193,N_45575,N_48680);
nand UO_3194 (O_3194,N_47190,N_47672);
nor UO_3195 (O_3195,N_47037,N_48258);
and UO_3196 (O_3196,N_47397,N_49745);
xnor UO_3197 (O_3197,N_49153,N_48793);
nand UO_3198 (O_3198,N_47883,N_47195);
or UO_3199 (O_3199,N_48957,N_48195);
or UO_3200 (O_3200,N_47605,N_47957);
or UO_3201 (O_3201,N_49092,N_45164);
and UO_3202 (O_3202,N_48717,N_48147);
or UO_3203 (O_3203,N_46610,N_45997);
nand UO_3204 (O_3204,N_49175,N_48135);
nand UO_3205 (O_3205,N_47704,N_46351);
nand UO_3206 (O_3206,N_48197,N_48205);
nor UO_3207 (O_3207,N_48143,N_46668);
nor UO_3208 (O_3208,N_49770,N_46075);
nor UO_3209 (O_3209,N_47195,N_48984);
xor UO_3210 (O_3210,N_49810,N_48876);
nor UO_3211 (O_3211,N_46172,N_48867);
or UO_3212 (O_3212,N_45931,N_46774);
nor UO_3213 (O_3213,N_49097,N_46910);
xor UO_3214 (O_3214,N_47707,N_49093);
nor UO_3215 (O_3215,N_47488,N_48445);
nor UO_3216 (O_3216,N_49987,N_46262);
and UO_3217 (O_3217,N_45238,N_48230);
nor UO_3218 (O_3218,N_48620,N_47015);
xor UO_3219 (O_3219,N_49554,N_48032);
nor UO_3220 (O_3220,N_48112,N_47890);
nand UO_3221 (O_3221,N_49755,N_49001);
or UO_3222 (O_3222,N_47254,N_46564);
and UO_3223 (O_3223,N_48306,N_45754);
xor UO_3224 (O_3224,N_48442,N_49899);
xor UO_3225 (O_3225,N_47954,N_48624);
and UO_3226 (O_3226,N_47171,N_45548);
xor UO_3227 (O_3227,N_47814,N_46400);
xnor UO_3228 (O_3228,N_46460,N_47342);
and UO_3229 (O_3229,N_49751,N_46041);
and UO_3230 (O_3230,N_48604,N_47538);
or UO_3231 (O_3231,N_47541,N_48347);
nor UO_3232 (O_3232,N_46259,N_48605);
and UO_3233 (O_3233,N_46936,N_48085);
xor UO_3234 (O_3234,N_49247,N_46540);
or UO_3235 (O_3235,N_46131,N_45444);
or UO_3236 (O_3236,N_46551,N_49146);
nor UO_3237 (O_3237,N_49858,N_47587);
nand UO_3238 (O_3238,N_47877,N_49367);
nor UO_3239 (O_3239,N_47715,N_47635);
nor UO_3240 (O_3240,N_48437,N_47356);
nor UO_3241 (O_3241,N_45183,N_49412);
or UO_3242 (O_3242,N_45009,N_48673);
or UO_3243 (O_3243,N_47642,N_48469);
or UO_3244 (O_3244,N_49641,N_49721);
and UO_3245 (O_3245,N_46707,N_49137);
nand UO_3246 (O_3246,N_45739,N_47339);
or UO_3247 (O_3247,N_48335,N_48621);
nor UO_3248 (O_3248,N_49216,N_46374);
and UO_3249 (O_3249,N_45677,N_46319);
nand UO_3250 (O_3250,N_46826,N_46232);
or UO_3251 (O_3251,N_46648,N_46359);
or UO_3252 (O_3252,N_47347,N_45577);
and UO_3253 (O_3253,N_47953,N_48306);
and UO_3254 (O_3254,N_49268,N_45238);
and UO_3255 (O_3255,N_49331,N_47055);
and UO_3256 (O_3256,N_47960,N_49304);
and UO_3257 (O_3257,N_48111,N_45687);
or UO_3258 (O_3258,N_46429,N_48249);
xnor UO_3259 (O_3259,N_45784,N_49405);
nor UO_3260 (O_3260,N_45295,N_47113);
and UO_3261 (O_3261,N_46393,N_46305);
or UO_3262 (O_3262,N_49067,N_47724);
xor UO_3263 (O_3263,N_49395,N_45752);
xor UO_3264 (O_3264,N_47261,N_49085);
nand UO_3265 (O_3265,N_46499,N_49475);
xnor UO_3266 (O_3266,N_45954,N_47229);
nor UO_3267 (O_3267,N_46677,N_48616);
nand UO_3268 (O_3268,N_46664,N_46975);
and UO_3269 (O_3269,N_48871,N_48613);
nor UO_3270 (O_3270,N_48773,N_47758);
xor UO_3271 (O_3271,N_47903,N_48927);
xnor UO_3272 (O_3272,N_45312,N_49534);
and UO_3273 (O_3273,N_48751,N_49412);
xnor UO_3274 (O_3274,N_48572,N_47892);
nor UO_3275 (O_3275,N_46866,N_45835);
nand UO_3276 (O_3276,N_49012,N_46544);
xor UO_3277 (O_3277,N_45212,N_48097);
nand UO_3278 (O_3278,N_47873,N_48585);
nor UO_3279 (O_3279,N_46520,N_45167);
nand UO_3280 (O_3280,N_47149,N_48384);
and UO_3281 (O_3281,N_48625,N_49006);
nor UO_3282 (O_3282,N_47819,N_49082);
xor UO_3283 (O_3283,N_45508,N_47820);
and UO_3284 (O_3284,N_49029,N_46183);
and UO_3285 (O_3285,N_49832,N_48929);
and UO_3286 (O_3286,N_48718,N_49974);
or UO_3287 (O_3287,N_49093,N_45557);
nor UO_3288 (O_3288,N_45596,N_48679);
nor UO_3289 (O_3289,N_47419,N_49947);
nor UO_3290 (O_3290,N_45308,N_48147);
xnor UO_3291 (O_3291,N_49392,N_46997);
nand UO_3292 (O_3292,N_47261,N_46395);
xor UO_3293 (O_3293,N_46273,N_47835);
nand UO_3294 (O_3294,N_47741,N_46928);
or UO_3295 (O_3295,N_49997,N_48865);
or UO_3296 (O_3296,N_46637,N_45697);
or UO_3297 (O_3297,N_46669,N_45043);
xnor UO_3298 (O_3298,N_48191,N_49194);
or UO_3299 (O_3299,N_46409,N_48789);
or UO_3300 (O_3300,N_48001,N_45324);
nand UO_3301 (O_3301,N_48233,N_47140);
nor UO_3302 (O_3302,N_47868,N_49137);
or UO_3303 (O_3303,N_45371,N_46951);
nand UO_3304 (O_3304,N_47224,N_46562);
nor UO_3305 (O_3305,N_47910,N_45757);
xor UO_3306 (O_3306,N_48436,N_49892);
or UO_3307 (O_3307,N_49685,N_47859);
nor UO_3308 (O_3308,N_47518,N_47582);
or UO_3309 (O_3309,N_48935,N_48044);
nor UO_3310 (O_3310,N_48397,N_47728);
and UO_3311 (O_3311,N_48648,N_48816);
xnor UO_3312 (O_3312,N_47864,N_48039);
nor UO_3313 (O_3313,N_47650,N_45891);
nand UO_3314 (O_3314,N_45507,N_48542);
and UO_3315 (O_3315,N_47109,N_45571);
nand UO_3316 (O_3316,N_48014,N_48052);
nor UO_3317 (O_3317,N_45915,N_47888);
nand UO_3318 (O_3318,N_47570,N_49173);
xor UO_3319 (O_3319,N_48926,N_45264);
and UO_3320 (O_3320,N_48410,N_46649);
nor UO_3321 (O_3321,N_45155,N_49472);
nor UO_3322 (O_3322,N_49561,N_48402);
or UO_3323 (O_3323,N_47840,N_49424);
nor UO_3324 (O_3324,N_49637,N_47288);
nand UO_3325 (O_3325,N_45456,N_46655);
or UO_3326 (O_3326,N_45954,N_45643);
nand UO_3327 (O_3327,N_46839,N_45512);
xor UO_3328 (O_3328,N_46269,N_48437);
nor UO_3329 (O_3329,N_46622,N_46076);
nor UO_3330 (O_3330,N_45006,N_46382);
nor UO_3331 (O_3331,N_46016,N_49740);
nand UO_3332 (O_3332,N_49743,N_47373);
nor UO_3333 (O_3333,N_48096,N_45012);
xnor UO_3334 (O_3334,N_47513,N_48134);
or UO_3335 (O_3335,N_48656,N_47100);
or UO_3336 (O_3336,N_45002,N_48980);
nand UO_3337 (O_3337,N_49052,N_48198);
xor UO_3338 (O_3338,N_49393,N_49689);
and UO_3339 (O_3339,N_49360,N_45517);
nand UO_3340 (O_3340,N_46512,N_46604);
or UO_3341 (O_3341,N_45263,N_48968);
xor UO_3342 (O_3342,N_48213,N_49814);
and UO_3343 (O_3343,N_47665,N_46590);
nor UO_3344 (O_3344,N_46543,N_47480);
nand UO_3345 (O_3345,N_49410,N_47258);
or UO_3346 (O_3346,N_47204,N_47775);
xor UO_3347 (O_3347,N_45231,N_49688);
and UO_3348 (O_3348,N_45584,N_47484);
and UO_3349 (O_3349,N_48339,N_49325);
nor UO_3350 (O_3350,N_45150,N_47811);
or UO_3351 (O_3351,N_49203,N_47192);
xor UO_3352 (O_3352,N_49925,N_46123);
nand UO_3353 (O_3353,N_47445,N_46051);
xor UO_3354 (O_3354,N_48758,N_49408);
and UO_3355 (O_3355,N_49623,N_46869);
or UO_3356 (O_3356,N_47010,N_48159);
and UO_3357 (O_3357,N_46073,N_48869);
xnor UO_3358 (O_3358,N_48968,N_49129);
or UO_3359 (O_3359,N_47308,N_49975);
nand UO_3360 (O_3360,N_48929,N_48514);
or UO_3361 (O_3361,N_46255,N_45914);
nand UO_3362 (O_3362,N_45747,N_48816);
nand UO_3363 (O_3363,N_46429,N_45325);
or UO_3364 (O_3364,N_45118,N_49911);
and UO_3365 (O_3365,N_45425,N_47006);
xor UO_3366 (O_3366,N_47005,N_49093);
and UO_3367 (O_3367,N_45357,N_49596);
nor UO_3368 (O_3368,N_47543,N_45497);
or UO_3369 (O_3369,N_45015,N_48964);
nand UO_3370 (O_3370,N_48955,N_45227);
nor UO_3371 (O_3371,N_48123,N_47051);
xor UO_3372 (O_3372,N_46505,N_47779);
or UO_3373 (O_3373,N_49241,N_46163);
and UO_3374 (O_3374,N_47409,N_46241);
and UO_3375 (O_3375,N_48081,N_48013);
nand UO_3376 (O_3376,N_46305,N_47244);
and UO_3377 (O_3377,N_46261,N_47954);
and UO_3378 (O_3378,N_45083,N_46310);
nand UO_3379 (O_3379,N_47498,N_46793);
or UO_3380 (O_3380,N_46899,N_49613);
and UO_3381 (O_3381,N_48013,N_48821);
and UO_3382 (O_3382,N_47775,N_48307);
nor UO_3383 (O_3383,N_46895,N_49164);
nor UO_3384 (O_3384,N_47568,N_46567);
or UO_3385 (O_3385,N_46143,N_47517);
and UO_3386 (O_3386,N_46374,N_45830);
and UO_3387 (O_3387,N_46254,N_49428);
and UO_3388 (O_3388,N_46858,N_45585);
xor UO_3389 (O_3389,N_49742,N_49354);
or UO_3390 (O_3390,N_49095,N_48150);
and UO_3391 (O_3391,N_46649,N_47181);
xnor UO_3392 (O_3392,N_48505,N_49890);
and UO_3393 (O_3393,N_45704,N_49141);
nand UO_3394 (O_3394,N_49250,N_49416);
nor UO_3395 (O_3395,N_49065,N_47604);
nand UO_3396 (O_3396,N_45285,N_48117);
and UO_3397 (O_3397,N_46889,N_49382);
nand UO_3398 (O_3398,N_49257,N_47764);
nor UO_3399 (O_3399,N_46764,N_47877);
or UO_3400 (O_3400,N_45039,N_47455);
xnor UO_3401 (O_3401,N_49907,N_46041);
xnor UO_3402 (O_3402,N_48259,N_47745);
nor UO_3403 (O_3403,N_47337,N_47548);
and UO_3404 (O_3404,N_46708,N_46956);
xnor UO_3405 (O_3405,N_45346,N_46542);
nor UO_3406 (O_3406,N_49915,N_46921);
nor UO_3407 (O_3407,N_48597,N_46863);
nand UO_3408 (O_3408,N_49417,N_46608);
or UO_3409 (O_3409,N_46063,N_48452);
nand UO_3410 (O_3410,N_47233,N_49603);
nor UO_3411 (O_3411,N_47342,N_48908);
nand UO_3412 (O_3412,N_46625,N_46787);
nor UO_3413 (O_3413,N_45812,N_45297);
nor UO_3414 (O_3414,N_45453,N_45187);
xnor UO_3415 (O_3415,N_48143,N_49318);
xor UO_3416 (O_3416,N_48104,N_46987);
nor UO_3417 (O_3417,N_49021,N_48303);
and UO_3418 (O_3418,N_45865,N_46522);
nand UO_3419 (O_3419,N_45925,N_49083);
nor UO_3420 (O_3420,N_46194,N_47661);
or UO_3421 (O_3421,N_46835,N_45924);
nand UO_3422 (O_3422,N_46107,N_48906);
and UO_3423 (O_3423,N_46068,N_46777);
nand UO_3424 (O_3424,N_47798,N_48862);
and UO_3425 (O_3425,N_46820,N_47006);
nand UO_3426 (O_3426,N_46563,N_48479);
xnor UO_3427 (O_3427,N_46011,N_46875);
nand UO_3428 (O_3428,N_45751,N_45574);
or UO_3429 (O_3429,N_48188,N_45928);
nand UO_3430 (O_3430,N_47587,N_45079);
and UO_3431 (O_3431,N_46541,N_48829);
xnor UO_3432 (O_3432,N_48494,N_45225);
xnor UO_3433 (O_3433,N_49271,N_49496);
and UO_3434 (O_3434,N_45971,N_48759);
nor UO_3435 (O_3435,N_48289,N_45018);
nand UO_3436 (O_3436,N_47131,N_47756);
or UO_3437 (O_3437,N_46649,N_45656);
nand UO_3438 (O_3438,N_45586,N_48225);
or UO_3439 (O_3439,N_46961,N_45703);
and UO_3440 (O_3440,N_47087,N_49145);
nor UO_3441 (O_3441,N_46290,N_47557);
and UO_3442 (O_3442,N_46400,N_45174);
and UO_3443 (O_3443,N_49465,N_45356);
nor UO_3444 (O_3444,N_45703,N_48036);
nand UO_3445 (O_3445,N_49980,N_47162);
and UO_3446 (O_3446,N_49815,N_47899);
xnor UO_3447 (O_3447,N_45674,N_46709);
nor UO_3448 (O_3448,N_46720,N_48823);
xnor UO_3449 (O_3449,N_46440,N_45143);
xor UO_3450 (O_3450,N_45624,N_46679);
and UO_3451 (O_3451,N_48310,N_45752);
and UO_3452 (O_3452,N_48905,N_45333);
and UO_3453 (O_3453,N_48088,N_47826);
and UO_3454 (O_3454,N_48889,N_47495);
and UO_3455 (O_3455,N_46049,N_49465);
and UO_3456 (O_3456,N_49579,N_48237);
xor UO_3457 (O_3457,N_46607,N_48670);
xor UO_3458 (O_3458,N_45385,N_47478);
nand UO_3459 (O_3459,N_46277,N_48193);
or UO_3460 (O_3460,N_49829,N_47604);
xnor UO_3461 (O_3461,N_47973,N_46823);
nor UO_3462 (O_3462,N_47665,N_49539);
nand UO_3463 (O_3463,N_47125,N_49373);
xnor UO_3464 (O_3464,N_46481,N_47134);
or UO_3465 (O_3465,N_49002,N_49700);
nor UO_3466 (O_3466,N_47353,N_46182);
xnor UO_3467 (O_3467,N_46077,N_49970);
nand UO_3468 (O_3468,N_45560,N_49278);
nand UO_3469 (O_3469,N_49903,N_49079);
nor UO_3470 (O_3470,N_49105,N_49703);
nor UO_3471 (O_3471,N_45138,N_45189);
xor UO_3472 (O_3472,N_48913,N_47590);
nand UO_3473 (O_3473,N_45109,N_45534);
nand UO_3474 (O_3474,N_47207,N_46429);
and UO_3475 (O_3475,N_49451,N_46647);
nor UO_3476 (O_3476,N_49787,N_45011);
or UO_3477 (O_3477,N_46904,N_48447);
nand UO_3478 (O_3478,N_46048,N_46320);
nor UO_3479 (O_3479,N_49420,N_48927);
xor UO_3480 (O_3480,N_45967,N_48472);
or UO_3481 (O_3481,N_47210,N_46619);
xor UO_3482 (O_3482,N_46296,N_48441);
or UO_3483 (O_3483,N_45825,N_46123);
xor UO_3484 (O_3484,N_48904,N_48712);
or UO_3485 (O_3485,N_49475,N_48642);
nand UO_3486 (O_3486,N_47114,N_47529);
or UO_3487 (O_3487,N_47420,N_46237);
or UO_3488 (O_3488,N_49925,N_48093);
xor UO_3489 (O_3489,N_45257,N_48726);
and UO_3490 (O_3490,N_47572,N_48986);
or UO_3491 (O_3491,N_49837,N_45071);
and UO_3492 (O_3492,N_47506,N_49242);
nor UO_3493 (O_3493,N_47201,N_46518);
and UO_3494 (O_3494,N_47823,N_47844);
xnor UO_3495 (O_3495,N_48842,N_47777);
nor UO_3496 (O_3496,N_46920,N_48768);
and UO_3497 (O_3497,N_49646,N_47279);
nand UO_3498 (O_3498,N_45222,N_48074);
nand UO_3499 (O_3499,N_47047,N_46360);
nand UO_3500 (O_3500,N_45370,N_45255);
nand UO_3501 (O_3501,N_49397,N_47278);
and UO_3502 (O_3502,N_48450,N_48458);
nor UO_3503 (O_3503,N_47705,N_45554);
nand UO_3504 (O_3504,N_48534,N_47142);
nor UO_3505 (O_3505,N_45980,N_45319);
and UO_3506 (O_3506,N_47850,N_49874);
or UO_3507 (O_3507,N_47059,N_49443);
xor UO_3508 (O_3508,N_49212,N_49333);
and UO_3509 (O_3509,N_49692,N_46001);
and UO_3510 (O_3510,N_48877,N_46757);
and UO_3511 (O_3511,N_46549,N_45342);
or UO_3512 (O_3512,N_46886,N_48397);
nand UO_3513 (O_3513,N_48859,N_47102);
or UO_3514 (O_3514,N_48851,N_47830);
nor UO_3515 (O_3515,N_45256,N_45199);
nand UO_3516 (O_3516,N_49673,N_45979);
and UO_3517 (O_3517,N_49655,N_49795);
or UO_3518 (O_3518,N_48967,N_49833);
or UO_3519 (O_3519,N_46236,N_49051);
or UO_3520 (O_3520,N_47976,N_49506);
or UO_3521 (O_3521,N_49833,N_47998);
nor UO_3522 (O_3522,N_48849,N_48983);
and UO_3523 (O_3523,N_47697,N_47052);
xor UO_3524 (O_3524,N_45097,N_47593);
and UO_3525 (O_3525,N_47824,N_46889);
and UO_3526 (O_3526,N_45188,N_45087);
and UO_3527 (O_3527,N_49699,N_49576);
nor UO_3528 (O_3528,N_46222,N_46224);
nand UO_3529 (O_3529,N_45522,N_45201);
xor UO_3530 (O_3530,N_45380,N_45112);
and UO_3531 (O_3531,N_47868,N_48893);
and UO_3532 (O_3532,N_46132,N_49371);
nor UO_3533 (O_3533,N_46523,N_49882);
or UO_3534 (O_3534,N_46917,N_48588);
or UO_3535 (O_3535,N_47220,N_47146);
nand UO_3536 (O_3536,N_46888,N_46581);
nand UO_3537 (O_3537,N_49670,N_46165);
nor UO_3538 (O_3538,N_48684,N_46230);
nor UO_3539 (O_3539,N_47958,N_48691);
or UO_3540 (O_3540,N_47129,N_49125);
and UO_3541 (O_3541,N_47657,N_46654);
or UO_3542 (O_3542,N_47603,N_45111);
or UO_3543 (O_3543,N_48148,N_45222);
nand UO_3544 (O_3544,N_49195,N_45990);
and UO_3545 (O_3545,N_46195,N_46285);
nand UO_3546 (O_3546,N_48214,N_45232);
and UO_3547 (O_3547,N_48561,N_47964);
nand UO_3548 (O_3548,N_45168,N_49606);
nand UO_3549 (O_3549,N_49188,N_46320);
nor UO_3550 (O_3550,N_46104,N_45904);
xnor UO_3551 (O_3551,N_49324,N_48208);
xnor UO_3552 (O_3552,N_46863,N_49104);
and UO_3553 (O_3553,N_45956,N_49121);
xnor UO_3554 (O_3554,N_48092,N_48006);
xnor UO_3555 (O_3555,N_46875,N_49293);
nand UO_3556 (O_3556,N_48432,N_46531);
and UO_3557 (O_3557,N_47213,N_45884);
and UO_3558 (O_3558,N_46560,N_47930);
and UO_3559 (O_3559,N_48694,N_47990);
or UO_3560 (O_3560,N_45094,N_48091);
nand UO_3561 (O_3561,N_45359,N_45334);
nand UO_3562 (O_3562,N_48818,N_48536);
nor UO_3563 (O_3563,N_48123,N_46870);
xor UO_3564 (O_3564,N_46258,N_46321);
nor UO_3565 (O_3565,N_46573,N_48304);
xnor UO_3566 (O_3566,N_48282,N_49048);
xnor UO_3567 (O_3567,N_45347,N_48275);
and UO_3568 (O_3568,N_48076,N_45895);
or UO_3569 (O_3569,N_47625,N_48918);
xor UO_3570 (O_3570,N_46715,N_46046);
nor UO_3571 (O_3571,N_49890,N_49349);
and UO_3572 (O_3572,N_48769,N_49192);
or UO_3573 (O_3573,N_47793,N_49409);
or UO_3574 (O_3574,N_49842,N_48645);
or UO_3575 (O_3575,N_45338,N_46344);
and UO_3576 (O_3576,N_48707,N_49347);
nor UO_3577 (O_3577,N_47161,N_46136);
xnor UO_3578 (O_3578,N_47499,N_47613);
or UO_3579 (O_3579,N_45298,N_47570);
nor UO_3580 (O_3580,N_49419,N_45577);
and UO_3581 (O_3581,N_48967,N_48973);
nand UO_3582 (O_3582,N_45372,N_46382);
or UO_3583 (O_3583,N_46074,N_45232);
xor UO_3584 (O_3584,N_47755,N_49706);
xor UO_3585 (O_3585,N_46707,N_46551);
nand UO_3586 (O_3586,N_46391,N_48885);
and UO_3587 (O_3587,N_46858,N_49923);
xor UO_3588 (O_3588,N_46078,N_46737);
xnor UO_3589 (O_3589,N_46860,N_45983);
nor UO_3590 (O_3590,N_48564,N_45471);
and UO_3591 (O_3591,N_48631,N_49655);
xor UO_3592 (O_3592,N_49911,N_45838);
xor UO_3593 (O_3593,N_49975,N_48235);
nor UO_3594 (O_3594,N_47825,N_45568);
and UO_3595 (O_3595,N_47843,N_45929);
nor UO_3596 (O_3596,N_49834,N_46461);
nand UO_3597 (O_3597,N_46423,N_45259);
and UO_3598 (O_3598,N_48907,N_48595);
nor UO_3599 (O_3599,N_49626,N_49977);
nand UO_3600 (O_3600,N_48671,N_45417);
xnor UO_3601 (O_3601,N_46383,N_47911);
and UO_3602 (O_3602,N_49185,N_47519);
nand UO_3603 (O_3603,N_46209,N_47227);
or UO_3604 (O_3604,N_49020,N_49997);
nor UO_3605 (O_3605,N_47121,N_49806);
or UO_3606 (O_3606,N_48345,N_48749);
xnor UO_3607 (O_3607,N_45249,N_47257);
nor UO_3608 (O_3608,N_47995,N_49990);
and UO_3609 (O_3609,N_48324,N_49770);
xor UO_3610 (O_3610,N_49508,N_45781);
xnor UO_3611 (O_3611,N_47703,N_47727);
xnor UO_3612 (O_3612,N_45961,N_46504);
nor UO_3613 (O_3613,N_48679,N_45584);
xnor UO_3614 (O_3614,N_46165,N_47735);
xnor UO_3615 (O_3615,N_46231,N_47036);
nor UO_3616 (O_3616,N_45438,N_49270);
nor UO_3617 (O_3617,N_49255,N_47261);
nand UO_3618 (O_3618,N_45158,N_49063);
nand UO_3619 (O_3619,N_47697,N_48326);
nand UO_3620 (O_3620,N_48937,N_49619);
or UO_3621 (O_3621,N_45413,N_49101);
and UO_3622 (O_3622,N_49122,N_46696);
or UO_3623 (O_3623,N_45912,N_49972);
xnor UO_3624 (O_3624,N_48256,N_49446);
xnor UO_3625 (O_3625,N_45911,N_45336);
nand UO_3626 (O_3626,N_47387,N_46109);
nor UO_3627 (O_3627,N_45297,N_47146);
nor UO_3628 (O_3628,N_45181,N_46602);
or UO_3629 (O_3629,N_49958,N_45138);
xor UO_3630 (O_3630,N_45688,N_49647);
or UO_3631 (O_3631,N_45265,N_49889);
or UO_3632 (O_3632,N_47938,N_48486);
and UO_3633 (O_3633,N_48094,N_49658);
nand UO_3634 (O_3634,N_46654,N_46029);
xnor UO_3635 (O_3635,N_46574,N_46088);
xnor UO_3636 (O_3636,N_48751,N_48284);
xor UO_3637 (O_3637,N_45415,N_49152);
xnor UO_3638 (O_3638,N_46596,N_49813);
nor UO_3639 (O_3639,N_45293,N_47732);
and UO_3640 (O_3640,N_45010,N_47061);
or UO_3641 (O_3641,N_47269,N_48976);
xor UO_3642 (O_3642,N_47887,N_47721);
or UO_3643 (O_3643,N_49251,N_49679);
xor UO_3644 (O_3644,N_48446,N_46541);
nor UO_3645 (O_3645,N_49986,N_48751);
and UO_3646 (O_3646,N_48535,N_49884);
or UO_3647 (O_3647,N_47791,N_45615);
nand UO_3648 (O_3648,N_46632,N_47705);
or UO_3649 (O_3649,N_47408,N_49747);
xor UO_3650 (O_3650,N_49424,N_47942);
nand UO_3651 (O_3651,N_46737,N_48881);
nand UO_3652 (O_3652,N_46661,N_47051);
xnor UO_3653 (O_3653,N_47606,N_47354);
nand UO_3654 (O_3654,N_49555,N_46104);
xor UO_3655 (O_3655,N_48467,N_47989);
or UO_3656 (O_3656,N_46422,N_47088);
or UO_3657 (O_3657,N_45393,N_46843);
xor UO_3658 (O_3658,N_46297,N_48458);
nand UO_3659 (O_3659,N_48178,N_47414);
or UO_3660 (O_3660,N_48438,N_46362);
and UO_3661 (O_3661,N_47581,N_46133);
xor UO_3662 (O_3662,N_46503,N_45918);
and UO_3663 (O_3663,N_49933,N_47549);
and UO_3664 (O_3664,N_45351,N_46658);
xor UO_3665 (O_3665,N_46917,N_49476);
nor UO_3666 (O_3666,N_48928,N_48053);
nand UO_3667 (O_3667,N_47426,N_46345);
or UO_3668 (O_3668,N_49465,N_48118);
nand UO_3669 (O_3669,N_48315,N_47250);
and UO_3670 (O_3670,N_48006,N_46001);
or UO_3671 (O_3671,N_45125,N_48078);
nand UO_3672 (O_3672,N_47805,N_49671);
xnor UO_3673 (O_3673,N_46691,N_47099);
and UO_3674 (O_3674,N_48627,N_46217);
nand UO_3675 (O_3675,N_46578,N_46315);
xor UO_3676 (O_3676,N_49151,N_46628);
and UO_3677 (O_3677,N_47252,N_48991);
or UO_3678 (O_3678,N_45047,N_47144);
xnor UO_3679 (O_3679,N_45154,N_49167);
nor UO_3680 (O_3680,N_48284,N_48474);
xnor UO_3681 (O_3681,N_45688,N_46868);
xor UO_3682 (O_3682,N_46818,N_45454);
or UO_3683 (O_3683,N_45174,N_48091);
nand UO_3684 (O_3684,N_45811,N_49295);
xor UO_3685 (O_3685,N_49306,N_46893);
and UO_3686 (O_3686,N_45479,N_45329);
xnor UO_3687 (O_3687,N_48245,N_47907);
and UO_3688 (O_3688,N_45975,N_48428);
or UO_3689 (O_3689,N_49489,N_49668);
nor UO_3690 (O_3690,N_47792,N_47847);
or UO_3691 (O_3691,N_45501,N_46928);
or UO_3692 (O_3692,N_47639,N_49680);
or UO_3693 (O_3693,N_48478,N_47411);
xor UO_3694 (O_3694,N_48965,N_46239);
nor UO_3695 (O_3695,N_47157,N_49502);
nand UO_3696 (O_3696,N_47564,N_46137);
nor UO_3697 (O_3697,N_48345,N_46594);
and UO_3698 (O_3698,N_47585,N_45043);
or UO_3699 (O_3699,N_48453,N_45817);
or UO_3700 (O_3700,N_47302,N_49540);
and UO_3701 (O_3701,N_45115,N_48783);
or UO_3702 (O_3702,N_45035,N_45784);
xor UO_3703 (O_3703,N_47637,N_46048);
and UO_3704 (O_3704,N_48019,N_49238);
nor UO_3705 (O_3705,N_49061,N_47663);
xor UO_3706 (O_3706,N_49830,N_46872);
nand UO_3707 (O_3707,N_49763,N_46528);
or UO_3708 (O_3708,N_47902,N_48398);
nand UO_3709 (O_3709,N_48665,N_47147);
nand UO_3710 (O_3710,N_48377,N_48957);
xnor UO_3711 (O_3711,N_45899,N_47629);
nand UO_3712 (O_3712,N_49243,N_48952);
and UO_3713 (O_3713,N_48123,N_46979);
and UO_3714 (O_3714,N_48433,N_46941);
nand UO_3715 (O_3715,N_49548,N_45905);
and UO_3716 (O_3716,N_49201,N_49008);
nor UO_3717 (O_3717,N_49926,N_48820);
xor UO_3718 (O_3718,N_45597,N_46228);
nand UO_3719 (O_3719,N_49194,N_47490);
nor UO_3720 (O_3720,N_49256,N_46385);
xor UO_3721 (O_3721,N_48004,N_46932);
or UO_3722 (O_3722,N_45590,N_47671);
and UO_3723 (O_3723,N_49830,N_46286);
xor UO_3724 (O_3724,N_45818,N_46585);
nor UO_3725 (O_3725,N_48864,N_48286);
nand UO_3726 (O_3726,N_45186,N_48856);
xor UO_3727 (O_3727,N_47289,N_49967);
or UO_3728 (O_3728,N_48635,N_45734);
or UO_3729 (O_3729,N_46624,N_45139);
or UO_3730 (O_3730,N_45021,N_45909);
xor UO_3731 (O_3731,N_45450,N_45827);
nor UO_3732 (O_3732,N_48995,N_47499);
nor UO_3733 (O_3733,N_49207,N_48034);
or UO_3734 (O_3734,N_46057,N_47897);
xor UO_3735 (O_3735,N_49600,N_48445);
xor UO_3736 (O_3736,N_48851,N_47973);
nand UO_3737 (O_3737,N_46772,N_48793);
nand UO_3738 (O_3738,N_47531,N_48687);
and UO_3739 (O_3739,N_48106,N_48586);
nand UO_3740 (O_3740,N_47910,N_48068);
xor UO_3741 (O_3741,N_49045,N_45758);
xor UO_3742 (O_3742,N_47507,N_49785);
nor UO_3743 (O_3743,N_46344,N_46462);
xnor UO_3744 (O_3744,N_46035,N_49722);
nor UO_3745 (O_3745,N_48193,N_47118);
nand UO_3746 (O_3746,N_46574,N_46894);
xor UO_3747 (O_3747,N_48634,N_49236);
and UO_3748 (O_3748,N_47884,N_47654);
nor UO_3749 (O_3749,N_46218,N_45789);
xnor UO_3750 (O_3750,N_48299,N_45527);
xnor UO_3751 (O_3751,N_47929,N_46331);
or UO_3752 (O_3752,N_49217,N_46534);
xor UO_3753 (O_3753,N_45682,N_45952);
xor UO_3754 (O_3754,N_45908,N_49059);
nand UO_3755 (O_3755,N_49367,N_48569);
or UO_3756 (O_3756,N_48284,N_49231);
or UO_3757 (O_3757,N_46787,N_47544);
nor UO_3758 (O_3758,N_46514,N_48344);
nand UO_3759 (O_3759,N_46311,N_49284);
nor UO_3760 (O_3760,N_45389,N_45786);
and UO_3761 (O_3761,N_45460,N_45554);
and UO_3762 (O_3762,N_48067,N_48096);
nor UO_3763 (O_3763,N_48171,N_46364);
nand UO_3764 (O_3764,N_46069,N_49970);
nand UO_3765 (O_3765,N_46838,N_49748);
and UO_3766 (O_3766,N_45602,N_47303);
xnor UO_3767 (O_3767,N_48886,N_45751);
nand UO_3768 (O_3768,N_49867,N_46269);
nor UO_3769 (O_3769,N_49590,N_48359);
and UO_3770 (O_3770,N_49109,N_49246);
or UO_3771 (O_3771,N_45182,N_46270);
nand UO_3772 (O_3772,N_49407,N_48582);
nor UO_3773 (O_3773,N_46850,N_49690);
and UO_3774 (O_3774,N_48943,N_47781);
nor UO_3775 (O_3775,N_49703,N_46444);
nor UO_3776 (O_3776,N_47896,N_46835);
or UO_3777 (O_3777,N_48493,N_48441);
nand UO_3778 (O_3778,N_48266,N_49325);
or UO_3779 (O_3779,N_48908,N_46967);
and UO_3780 (O_3780,N_45764,N_48265);
nor UO_3781 (O_3781,N_45215,N_49132);
and UO_3782 (O_3782,N_45199,N_49138);
and UO_3783 (O_3783,N_46972,N_47021);
or UO_3784 (O_3784,N_48142,N_49482);
nand UO_3785 (O_3785,N_45855,N_45582);
nor UO_3786 (O_3786,N_48471,N_47249);
and UO_3787 (O_3787,N_48452,N_46874);
nand UO_3788 (O_3788,N_48363,N_48711);
and UO_3789 (O_3789,N_48885,N_49667);
or UO_3790 (O_3790,N_49496,N_49036);
and UO_3791 (O_3791,N_46858,N_45726);
and UO_3792 (O_3792,N_48732,N_45748);
nand UO_3793 (O_3793,N_48733,N_48155);
nor UO_3794 (O_3794,N_45171,N_46931);
nand UO_3795 (O_3795,N_49382,N_48176);
or UO_3796 (O_3796,N_47277,N_47234);
and UO_3797 (O_3797,N_47029,N_47508);
nor UO_3798 (O_3798,N_48738,N_47131);
nand UO_3799 (O_3799,N_49547,N_47271);
nor UO_3800 (O_3800,N_49799,N_46195);
xor UO_3801 (O_3801,N_46725,N_45578);
xnor UO_3802 (O_3802,N_47031,N_49230);
or UO_3803 (O_3803,N_48696,N_45640);
nand UO_3804 (O_3804,N_48694,N_47561);
or UO_3805 (O_3805,N_49287,N_45924);
nor UO_3806 (O_3806,N_47380,N_45458);
nor UO_3807 (O_3807,N_45297,N_48521);
nor UO_3808 (O_3808,N_48750,N_46359);
nand UO_3809 (O_3809,N_45598,N_48902);
and UO_3810 (O_3810,N_45530,N_46628);
and UO_3811 (O_3811,N_45439,N_47825);
and UO_3812 (O_3812,N_47681,N_49344);
nor UO_3813 (O_3813,N_49843,N_48281);
nand UO_3814 (O_3814,N_47603,N_49841);
and UO_3815 (O_3815,N_49903,N_47534);
and UO_3816 (O_3816,N_47597,N_46398);
or UO_3817 (O_3817,N_46595,N_47832);
xor UO_3818 (O_3818,N_46080,N_49571);
xnor UO_3819 (O_3819,N_49167,N_49787);
nand UO_3820 (O_3820,N_49057,N_49479);
or UO_3821 (O_3821,N_45559,N_46602);
xor UO_3822 (O_3822,N_46453,N_49309);
and UO_3823 (O_3823,N_48988,N_46990);
and UO_3824 (O_3824,N_48811,N_45571);
nor UO_3825 (O_3825,N_45003,N_48965);
xor UO_3826 (O_3826,N_47207,N_47178);
xor UO_3827 (O_3827,N_45385,N_47438);
nand UO_3828 (O_3828,N_48008,N_45056);
nand UO_3829 (O_3829,N_48084,N_47611);
nor UO_3830 (O_3830,N_46009,N_48456);
and UO_3831 (O_3831,N_46969,N_48753);
nor UO_3832 (O_3832,N_45022,N_48310);
xor UO_3833 (O_3833,N_48123,N_46161);
nand UO_3834 (O_3834,N_48587,N_47596);
or UO_3835 (O_3835,N_46216,N_48002);
and UO_3836 (O_3836,N_46799,N_49598);
nor UO_3837 (O_3837,N_47649,N_45855);
nand UO_3838 (O_3838,N_47620,N_49494);
and UO_3839 (O_3839,N_48055,N_47845);
or UO_3840 (O_3840,N_46295,N_47144);
xor UO_3841 (O_3841,N_49825,N_48233);
nor UO_3842 (O_3842,N_48728,N_48360);
xor UO_3843 (O_3843,N_46604,N_45250);
or UO_3844 (O_3844,N_45692,N_47120);
nor UO_3845 (O_3845,N_49322,N_46759);
nand UO_3846 (O_3846,N_48805,N_49435);
or UO_3847 (O_3847,N_46992,N_45528);
and UO_3848 (O_3848,N_49144,N_46799);
and UO_3849 (O_3849,N_45448,N_47806);
xnor UO_3850 (O_3850,N_48509,N_46413);
or UO_3851 (O_3851,N_49628,N_49785);
or UO_3852 (O_3852,N_48181,N_47943);
nor UO_3853 (O_3853,N_45488,N_48282);
or UO_3854 (O_3854,N_47021,N_47375);
nand UO_3855 (O_3855,N_49913,N_45742);
nand UO_3856 (O_3856,N_45707,N_45309);
and UO_3857 (O_3857,N_46467,N_48108);
or UO_3858 (O_3858,N_47774,N_47350);
or UO_3859 (O_3859,N_45088,N_45797);
or UO_3860 (O_3860,N_48485,N_46905);
or UO_3861 (O_3861,N_49949,N_48363);
nor UO_3862 (O_3862,N_49643,N_47983);
nand UO_3863 (O_3863,N_46050,N_48946);
xnor UO_3864 (O_3864,N_46908,N_49435);
and UO_3865 (O_3865,N_48782,N_47669);
and UO_3866 (O_3866,N_45545,N_46077);
xor UO_3867 (O_3867,N_46948,N_47239);
xnor UO_3868 (O_3868,N_49163,N_49365);
nand UO_3869 (O_3869,N_46182,N_45960);
nor UO_3870 (O_3870,N_48788,N_48841);
or UO_3871 (O_3871,N_46756,N_46211);
or UO_3872 (O_3872,N_46082,N_49502);
nand UO_3873 (O_3873,N_47307,N_49640);
or UO_3874 (O_3874,N_46645,N_48960);
nor UO_3875 (O_3875,N_47395,N_48151);
nand UO_3876 (O_3876,N_46192,N_46694);
or UO_3877 (O_3877,N_47909,N_48311);
nor UO_3878 (O_3878,N_46727,N_45550);
nor UO_3879 (O_3879,N_45707,N_45940);
nor UO_3880 (O_3880,N_45756,N_49840);
xor UO_3881 (O_3881,N_46428,N_45657);
nor UO_3882 (O_3882,N_45062,N_47067);
xor UO_3883 (O_3883,N_45447,N_46026);
or UO_3884 (O_3884,N_49344,N_45880);
xnor UO_3885 (O_3885,N_45668,N_46411);
nand UO_3886 (O_3886,N_49662,N_48268);
nand UO_3887 (O_3887,N_49864,N_49805);
nor UO_3888 (O_3888,N_49198,N_49367);
and UO_3889 (O_3889,N_46022,N_49381);
nand UO_3890 (O_3890,N_47158,N_49919);
xnor UO_3891 (O_3891,N_46237,N_46535);
nor UO_3892 (O_3892,N_47267,N_48453);
xnor UO_3893 (O_3893,N_47643,N_46510);
xnor UO_3894 (O_3894,N_46581,N_46677);
nand UO_3895 (O_3895,N_45012,N_49885);
and UO_3896 (O_3896,N_47582,N_48484);
xnor UO_3897 (O_3897,N_47029,N_49168);
nor UO_3898 (O_3898,N_47828,N_48730);
and UO_3899 (O_3899,N_49177,N_49370);
and UO_3900 (O_3900,N_46194,N_45293);
xnor UO_3901 (O_3901,N_47570,N_49619);
xor UO_3902 (O_3902,N_48438,N_48908);
and UO_3903 (O_3903,N_48038,N_45882);
or UO_3904 (O_3904,N_49354,N_45449);
or UO_3905 (O_3905,N_48193,N_47991);
nor UO_3906 (O_3906,N_47183,N_49209);
or UO_3907 (O_3907,N_46847,N_46134);
or UO_3908 (O_3908,N_47443,N_48160);
xnor UO_3909 (O_3909,N_48049,N_47400);
or UO_3910 (O_3910,N_45549,N_48868);
nor UO_3911 (O_3911,N_48934,N_49965);
or UO_3912 (O_3912,N_45240,N_47652);
or UO_3913 (O_3913,N_48139,N_49116);
or UO_3914 (O_3914,N_48692,N_48668);
xor UO_3915 (O_3915,N_47681,N_49921);
nor UO_3916 (O_3916,N_46090,N_49156);
nor UO_3917 (O_3917,N_48965,N_47998);
or UO_3918 (O_3918,N_46081,N_48905);
xnor UO_3919 (O_3919,N_48222,N_46987);
and UO_3920 (O_3920,N_48476,N_47454);
and UO_3921 (O_3921,N_47701,N_48013);
and UO_3922 (O_3922,N_46275,N_47118);
nand UO_3923 (O_3923,N_48538,N_46661);
nand UO_3924 (O_3924,N_48651,N_46262);
nor UO_3925 (O_3925,N_46125,N_45066);
nand UO_3926 (O_3926,N_47767,N_47491);
or UO_3927 (O_3927,N_48619,N_49910);
nand UO_3928 (O_3928,N_45799,N_49901);
nand UO_3929 (O_3929,N_49895,N_47274);
nor UO_3930 (O_3930,N_45471,N_47892);
and UO_3931 (O_3931,N_45175,N_45382);
and UO_3932 (O_3932,N_47894,N_45075);
and UO_3933 (O_3933,N_47156,N_47762);
xor UO_3934 (O_3934,N_49818,N_49159);
xnor UO_3935 (O_3935,N_46791,N_48301);
nand UO_3936 (O_3936,N_45350,N_46013);
nor UO_3937 (O_3937,N_47227,N_49706);
nand UO_3938 (O_3938,N_47801,N_45362);
or UO_3939 (O_3939,N_46826,N_45580);
xnor UO_3940 (O_3940,N_45825,N_45137);
or UO_3941 (O_3941,N_47183,N_48599);
or UO_3942 (O_3942,N_47428,N_46882);
xnor UO_3943 (O_3943,N_46765,N_45001);
and UO_3944 (O_3944,N_48696,N_46889);
or UO_3945 (O_3945,N_49333,N_45170);
or UO_3946 (O_3946,N_47155,N_47059);
nor UO_3947 (O_3947,N_46158,N_46489);
nor UO_3948 (O_3948,N_46973,N_46558);
nand UO_3949 (O_3949,N_45344,N_48731);
and UO_3950 (O_3950,N_48689,N_48789);
nor UO_3951 (O_3951,N_47919,N_46799);
or UO_3952 (O_3952,N_45637,N_48979);
xnor UO_3953 (O_3953,N_48583,N_47911);
and UO_3954 (O_3954,N_47187,N_46132);
or UO_3955 (O_3955,N_45488,N_46497);
nand UO_3956 (O_3956,N_49540,N_47266);
xnor UO_3957 (O_3957,N_48977,N_49208);
or UO_3958 (O_3958,N_46187,N_48866);
nor UO_3959 (O_3959,N_47643,N_48606);
xnor UO_3960 (O_3960,N_45460,N_49134);
xnor UO_3961 (O_3961,N_49364,N_45530);
and UO_3962 (O_3962,N_47272,N_47003);
xor UO_3963 (O_3963,N_45137,N_46277);
nand UO_3964 (O_3964,N_45551,N_49946);
nor UO_3965 (O_3965,N_47053,N_45448);
or UO_3966 (O_3966,N_46231,N_45328);
or UO_3967 (O_3967,N_46403,N_45296);
nand UO_3968 (O_3968,N_46570,N_45454);
xor UO_3969 (O_3969,N_45786,N_48386);
nand UO_3970 (O_3970,N_48569,N_48645);
or UO_3971 (O_3971,N_49318,N_46590);
and UO_3972 (O_3972,N_45750,N_47068);
nor UO_3973 (O_3973,N_47696,N_45429);
or UO_3974 (O_3974,N_46410,N_47706);
or UO_3975 (O_3975,N_46940,N_49639);
or UO_3976 (O_3976,N_49311,N_48052);
xnor UO_3977 (O_3977,N_49391,N_45736);
nand UO_3978 (O_3978,N_49588,N_47531);
nand UO_3979 (O_3979,N_47321,N_47437);
xnor UO_3980 (O_3980,N_47591,N_46363);
and UO_3981 (O_3981,N_49793,N_49207);
nand UO_3982 (O_3982,N_49565,N_47824);
or UO_3983 (O_3983,N_47968,N_49722);
or UO_3984 (O_3984,N_48402,N_48453);
or UO_3985 (O_3985,N_45618,N_48424);
xnor UO_3986 (O_3986,N_48571,N_48813);
nor UO_3987 (O_3987,N_45343,N_46532);
or UO_3988 (O_3988,N_46533,N_45074);
nor UO_3989 (O_3989,N_48786,N_46509);
nand UO_3990 (O_3990,N_49735,N_47156);
or UO_3991 (O_3991,N_46279,N_48946);
or UO_3992 (O_3992,N_48806,N_47899);
nor UO_3993 (O_3993,N_46814,N_48662);
or UO_3994 (O_3994,N_46916,N_45984);
or UO_3995 (O_3995,N_49136,N_48320);
and UO_3996 (O_3996,N_48822,N_45378);
xor UO_3997 (O_3997,N_49209,N_47121);
and UO_3998 (O_3998,N_49954,N_45091);
and UO_3999 (O_3999,N_45565,N_48253);
and UO_4000 (O_4000,N_46795,N_49036);
nor UO_4001 (O_4001,N_48486,N_49661);
or UO_4002 (O_4002,N_47254,N_45255);
or UO_4003 (O_4003,N_49991,N_46427);
nand UO_4004 (O_4004,N_46153,N_48646);
nor UO_4005 (O_4005,N_49370,N_48405);
and UO_4006 (O_4006,N_47511,N_48485);
xor UO_4007 (O_4007,N_47267,N_46052);
nand UO_4008 (O_4008,N_45522,N_46944);
nand UO_4009 (O_4009,N_48837,N_49674);
nor UO_4010 (O_4010,N_49200,N_47199);
or UO_4011 (O_4011,N_49827,N_48308);
or UO_4012 (O_4012,N_46490,N_46010);
nand UO_4013 (O_4013,N_48581,N_47533);
or UO_4014 (O_4014,N_47295,N_45465);
and UO_4015 (O_4015,N_48633,N_46012);
or UO_4016 (O_4016,N_45197,N_47889);
xor UO_4017 (O_4017,N_47886,N_47412);
and UO_4018 (O_4018,N_45502,N_45559);
nand UO_4019 (O_4019,N_49734,N_47756);
nor UO_4020 (O_4020,N_47798,N_49902);
nor UO_4021 (O_4021,N_45647,N_47175);
or UO_4022 (O_4022,N_47810,N_47272);
nor UO_4023 (O_4023,N_45566,N_49818);
nand UO_4024 (O_4024,N_46490,N_49741);
xor UO_4025 (O_4025,N_47196,N_48133);
or UO_4026 (O_4026,N_45947,N_49412);
or UO_4027 (O_4027,N_47434,N_48294);
xnor UO_4028 (O_4028,N_47403,N_47262);
nor UO_4029 (O_4029,N_48646,N_45990);
and UO_4030 (O_4030,N_49282,N_49629);
nor UO_4031 (O_4031,N_45570,N_46002);
nor UO_4032 (O_4032,N_46358,N_46773);
nand UO_4033 (O_4033,N_48507,N_45619);
nand UO_4034 (O_4034,N_47223,N_45561);
xor UO_4035 (O_4035,N_48305,N_48114);
nor UO_4036 (O_4036,N_48051,N_46716);
nor UO_4037 (O_4037,N_47824,N_46364);
nor UO_4038 (O_4038,N_48758,N_48996);
nand UO_4039 (O_4039,N_48439,N_45118);
and UO_4040 (O_4040,N_49282,N_49584);
and UO_4041 (O_4041,N_49850,N_45734);
nand UO_4042 (O_4042,N_48586,N_45903);
or UO_4043 (O_4043,N_47581,N_48592);
and UO_4044 (O_4044,N_49880,N_48960);
and UO_4045 (O_4045,N_49624,N_46495);
nor UO_4046 (O_4046,N_45833,N_47656);
and UO_4047 (O_4047,N_49569,N_47441);
nor UO_4048 (O_4048,N_47476,N_48891);
nor UO_4049 (O_4049,N_49586,N_47764);
xor UO_4050 (O_4050,N_46693,N_48877);
and UO_4051 (O_4051,N_47039,N_46459);
nor UO_4052 (O_4052,N_49469,N_49297);
and UO_4053 (O_4053,N_46214,N_49392);
nor UO_4054 (O_4054,N_49953,N_49601);
nand UO_4055 (O_4055,N_48228,N_47640);
or UO_4056 (O_4056,N_47618,N_49065);
or UO_4057 (O_4057,N_48337,N_46626);
xor UO_4058 (O_4058,N_45088,N_49376);
nor UO_4059 (O_4059,N_47772,N_49788);
and UO_4060 (O_4060,N_46162,N_45359);
nor UO_4061 (O_4061,N_48854,N_45730);
nand UO_4062 (O_4062,N_47993,N_48764);
xor UO_4063 (O_4063,N_49807,N_46203);
and UO_4064 (O_4064,N_46889,N_48356);
nand UO_4065 (O_4065,N_46879,N_46660);
nor UO_4066 (O_4066,N_46783,N_47932);
and UO_4067 (O_4067,N_48029,N_49134);
nor UO_4068 (O_4068,N_48419,N_47733);
or UO_4069 (O_4069,N_48429,N_47687);
and UO_4070 (O_4070,N_45731,N_49995);
nor UO_4071 (O_4071,N_49044,N_46358);
or UO_4072 (O_4072,N_48187,N_45698);
and UO_4073 (O_4073,N_47451,N_48937);
xor UO_4074 (O_4074,N_46800,N_47532);
xor UO_4075 (O_4075,N_47605,N_46339);
nor UO_4076 (O_4076,N_48782,N_48355);
and UO_4077 (O_4077,N_45350,N_49995);
or UO_4078 (O_4078,N_45611,N_48643);
or UO_4079 (O_4079,N_45444,N_45892);
and UO_4080 (O_4080,N_48849,N_46740);
nor UO_4081 (O_4081,N_49268,N_46430);
nor UO_4082 (O_4082,N_49379,N_47101);
nand UO_4083 (O_4083,N_47960,N_45377);
xor UO_4084 (O_4084,N_47055,N_46624);
nand UO_4085 (O_4085,N_46330,N_45255);
and UO_4086 (O_4086,N_49125,N_46698);
nand UO_4087 (O_4087,N_45777,N_48630);
or UO_4088 (O_4088,N_48133,N_49448);
nor UO_4089 (O_4089,N_48650,N_48388);
xor UO_4090 (O_4090,N_49085,N_46739);
nor UO_4091 (O_4091,N_45071,N_46063);
xnor UO_4092 (O_4092,N_46621,N_49101);
nand UO_4093 (O_4093,N_48583,N_45834);
nand UO_4094 (O_4094,N_49511,N_49563);
nand UO_4095 (O_4095,N_47657,N_46328);
and UO_4096 (O_4096,N_47206,N_46179);
and UO_4097 (O_4097,N_45925,N_46876);
or UO_4098 (O_4098,N_49244,N_46270);
xnor UO_4099 (O_4099,N_45121,N_48189);
nand UO_4100 (O_4100,N_47370,N_47719);
and UO_4101 (O_4101,N_45925,N_46956);
or UO_4102 (O_4102,N_47551,N_46508);
xnor UO_4103 (O_4103,N_48351,N_45979);
or UO_4104 (O_4104,N_47711,N_49514);
nand UO_4105 (O_4105,N_47751,N_49740);
xnor UO_4106 (O_4106,N_46015,N_49065);
xnor UO_4107 (O_4107,N_47433,N_47778);
nor UO_4108 (O_4108,N_46542,N_46801);
nand UO_4109 (O_4109,N_46873,N_49357);
and UO_4110 (O_4110,N_46841,N_49189);
and UO_4111 (O_4111,N_46342,N_47026);
xnor UO_4112 (O_4112,N_47781,N_49326);
or UO_4113 (O_4113,N_45346,N_48765);
nand UO_4114 (O_4114,N_49242,N_47509);
and UO_4115 (O_4115,N_46824,N_48467);
xor UO_4116 (O_4116,N_47793,N_49917);
xnor UO_4117 (O_4117,N_47174,N_47849);
nor UO_4118 (O_4118,N_49836,N_46347);
xnor UO_4119 (O_4119,N_46590,N_48299);
xor UO_4120 (O_4120,N_48245,N_49435);
nand UO_4121 (O_4121,N_47851,N_47093);
xnor UO_4122 (O_4122,N_49898,N_48556);
and UO_4123 (O_4123,N_49419,N_49471);
xor UO_4124 (O_4124,N_47842,N_45789);
xnor UO_4125 (O_4125,N_48099,N_46686);
and UO_4126 (O_4126,N_48622,N_48985);
nand UO_4127 (O_4127,N_45155,N_49484);
nor UO_4128 (O_4128,N_49425,N_47221);
nand UO_4129 (O_4129,N_45424,N_48121);
or UO_4130 (O_4130,N_45926,N_47364);
xor UO_4131 (O_4131,N_47320,N_47094);
nand UO_4132 (O_4132,N_47073,N_47027);
xor UO_4133 (O_4133,N_47143,N_46566);
and UO_4134 (O_4134,N_46174,N_45742);
or UO_4135 (O_4135,N_48453,N_48199);
and UO_4136 (O_4136,N_47486,N_47605);
xor UO_4137 (O_4137,N_47496,N_49580);
nor UO_4138 (O_4138,N_46283,N_45567);
or UO_4139 (O_4139,N_46346,N_48004);
and UO_4140 (O_4140,N_45192,N_45814);
nor UO_4141 (O_4141,N_45525,N_47962);
nor UO_4142 (O_4142,N_47560,N_49292);
and UO_4143 (O_4143,N_47709,N_47824);
and UO_4144 (O_4144,N_47551,N_47692);
xnor UO_4145 (O_4145,N_46406,N_47100);
xor UO_4146 (O_4146,N_45381,N_45823);
or UO_4147 (O_4147,N_49732,N_45724);
xnor UO_4148 (O_4148,N_47980,N_49908);
or UO_4149 (O_4149,N_46128,N_48195);
or UO_4150 (O_4150,N_47426,N_48343);
nor UO_4151 (O_4151,N_48636,N_45095);
nor UO_4152 (O_4152,N_46731,N_47234);
and UO_4153 (O_4153,N_46143,N_46276);
xnor UO_4154 (O_4154,N_47295,N_48943);
and UO_4155 (O_4155,N_45649,N_49418);
nand UO_4156 (O_4156,N_49597,N_45523);
and UO_4157 (O_4157,N_46478,N_46282);
and UO_4158 (O_4158,N_49152,N_46111);
xnor UO_4159 (O_4159,N_49495,N_47340);
or UO_4160 (O_4160,N_48323,N_47533);
xor UO_4161 (O_4161,N_48050,N_46289);
nand UO_4162 (O_4162,N_45114,N_48343);
or UO_4163 (O_4163,N_48320,N_45403);
xnor UO_4164 (O_4164,N_48403,N_48427);
or UO_4165 (O_4165,N_47400,N_46501);
nand UO_4166 (O_4166,N_49507,N_48998);
nand UO_4167 (O_4167,N_49879,N_47190);
nand UO_4168 (O_4168,N_49858,N_49002);
or UO_4169 (O_4169,N_47271,N_47371);
xor UO_4170 (O_4170,N_45933,N_46903);
nor UO_4171 (O_4171,N_49796,N_49769);
or UO_4172 (O_4172,N_47393,N_46863);
xor UO_4173 (O_4173,N_45732,N_45025);
nand UO_4174 (O_4174,N_48734,N_49064);
or UO_4175 (O_4175,N_49622,N_49326);
and UO_4176 (O_4176,N_47836,N_48836);
or UO_4177 (O_4177,N_49368,N_48337);
or UO_4178 (O_4178,N_49561,N_46426);
xnor UO_4179 (O_4179,N_49865,N_49403);
and UO_4180 (O_4180,N_46460,N_46916);
xor UO_4181 (O_4181,N_45715,N_48993);
and UO_4182 (O_4182,N_47365,N_45450);
nand UO_4183 (O_4183,N_48217,N_46506);
or UO_4184 (O_4184,N_48300,N_46655);
nor UO_4185 (O_4185,N_47364,N_45632);
and UO_4186 (O_4186,N_48098,N_48000);
nand UO_4187 (O_4187,N_47519,N_49373);
and UO_4188 (O_4188,N_48013,N_48993);
and UO_4189 (O_4189,N_45859,N_45513);
or UO_4190 (O_4190,N_46853,N_46112);
xnor UO_4191 (O_4191,N_49330,N_46795);
and UO_4192 (O_4192,N_48708,N_47262);
nor UO_4193 (O_4193,N_48848,N_45346);
nor UO_4194 (O_4194,N_45013,N_47713);
and UO_4195 (O_4195,N_49127,N_46931);
nand UO_4196 (O_4196,N_45624,N_49290);
xnor UO_4197 (O_4197,N_48286,N_45529);
nand UO_4198 (O_4198,N_47585,N_45861);
or UO_4199 (O_4199,N_45277,N_45930);
nand UO_4200 (O_4200,N_48666,N_49146);
or UO_4201 (O_4201,N_46637,N_47657);
nand UO_4202 (O_4202,N_48059,N_48574);
or UO_4203 (O_4203,N_46352,N_47491);
and UO_4204 (O_4204,N_45069,N_48661);
and UO_4205 (O_4205,N_46143,N_45238);
nand UO_4206 (O_4206,N_49334,N_46376);
nor UO_4207 (O_4207,N_49595,N_45441);
nor UO_4208 (O_4208,N_47809,N_46386);
nor UO_4209 (O_4209,N_45200,N_49825);
xor UO_4210 (O_4210,N_48335,N_48571);
nand UO_4211 (O_4211,N_49615,N_47886);
or UO_4212 (O_4212,N_49005,N_46438);
nand UO_4213 (O_4213,N_48396,N_47148);
or UO_4214 (O_4214,N_45810,N_48232);
nor UO_4215 (O_4215,N_45146,N_48729);
xnor UO_4216 (O_4216,N_47800,N_45062);
nand UO_4217 (O_4217,N_48063,N_46216);
xor UO_4218 (O_4218,N_47103,N_47104);
nor UO_4219 (O_4219,N_45378,N_45687);
and UO_4220 (O_4220,N_45953,N_45022);
nor UO_4221 (O_4221,N_45711,N_48024);
nand UO_4222 (O_4222,N_45672,N_48808);
or UO_4223 (O_4223,N_45867,N_47253);
xor UO_4224 (O_4224,N_46447,N_48617);
or UO_4225 (O_4225,N_48992,N_48545);
and UO_4226 (O_4226,N_45630,N_47284);
nor UO_4227 (O_4227,N_49883,N_45978);
nor UO_4228 (O_4228,N_46733,N_48848);
or UO_4229 (O_4229,N_48904,N_49528);
nor UO_4230 (O_4230,N_47734,N_45171);
nor UO_4231 (O_4231,N_49003,N_48317);
xnor UO_4232 (O_4232,N_47777,N_48840);
or UO_4233 (O_4233,N_47383,N_46201);
nor UO_4234 (O_4234,N_46113,N_45533);
or UO_4235 (O_4235,N_45052,N_47332);
nor UO_4236 (O_4236,N_49483,N_48333);
nand UO_4237 (O_4237,N_45833,N_48642);
nand UO_4238 (O_4238,N_47600,N_48764);
xor UO_4239 (O_4239,N_49289,N_46499);
or UO_4240 (O_4240,N_45841,N_45875);
and UO_4241 (O_4241,N_47724,N_46157);
nand UO_4242 (O_4242,N_49232,N_45179);
or UO_4243 (O_4243,N_46757,N_48610);
and UO_4244 (O_4244,N_46195,N_49703);
or UO_4245 (O_4245,N_45185,N_45046);
nor UO_4246 (O_4246,N_45575,N_49467);
nand UO_4247 (O_4247,N_48752,N_49950);
nor UO_4248 (O_4248,N_48493,N_46046);
nor UO_4249 (O_4249,N_46711,N_49396);
nand UO_4250 (O_4250,N_48130,N_47588);
nor UO_4251 (O_4251,N_45518,N_49256);
xnor UO_4252 (O_4252,N_48456,N_49211);
or UO_4253 (O_4253,N_49851,N_45613);
and UO_4254 (O_4254,N_48288,N_48161);
xnor UO_4255 (O_4255,N_46826,N_46320);
or UO_4256 (O_4256,N_47484,N_48058);
nor UO_4257 (O_4257,N_47044,N_45573);
and UO_4258 (O_4258,N_46526,N_49519);
and UO_4259 (O_4259,N_48989,N_45358);
nand UO_4260 (O_4260,N_48984,N_46408);
and UO_4261 (O_4261,N_48642,N_46526);
nand UO_4262 (O_4262,N_46811,N_49184);
and UO_4263 (O_4263,N_49386,N_46571);
and UO_4264 (O_4264,N_45348,N_49212);
nand UO_4265 (O_4265,N_47820,N_49247);
nor UO_4266 (O_4266,N_49922,N_48583);
or UO_4267 (O_4267,N_47314,N_47249);
xnor UO_4268 (O_4268,N_46255,N_46493);
nor UO_4269 (O_4269,N_48338,N_48276);
xnor UO_4270 (O_4270,N_49705,N_48742);
nor UO_4271 (O_4271,N_48611,N_48478);
and UO_4272 (O_4272,N_49722,N_47080);
nand UO_4273 (O_4273,N_48153,N_48475);
and UO_4274 (O_4274,N_48966,N_48771);
xnor UO_4275 (O_4275,N_48858,N_46083);
or UO_4276 (O_4276,N_48385,N_47155);
or UO_4277 (O_4277,N_48651,N_46972);
or UO_4278 (O_4278,N_45749,N_45438);
or UO_4279 (O_4279,N_48288,N_48191);
or UO_4280 (O_4280,N_48014,N_47129);
and UO_4281 (O_4281,N_48056,N_47987);
nor UO_4282 (O_4282,N_45310,N_45053);
nor UO_4283 (O_4283,N_48424,N_46381);
xor UO_4284 (O_4284,N_49782,N_47512);
and UO_4285 (O_4285,N_46335,N_47927);
and UO_4286 (O_4286,N_48478,N_49874);
and UO_4287 (O_4287,N_48580,N_48678);
nand UO_4288 (O_4288,N_49111,N_47042);
nand UO_4289 (O_4289,N_45526,N_47099);
xnor UO_4290 (O_4290,N_48939,N_46043);
and UO_4291 (O_4291,N_46073,N_49415);
nand UO_4292 (O_4292,N_47036,N_46637);
and UO_4293 (O_4293,N_47568,N_46774);
or UO_4294 (O_4294,N_49347,N_47015);
nand UO_4295 (O_4295,N_48441,N_49822);
or UO_4296 (O_4296,N_47761,N_47402);
nand UO_4297 (O_4297,N_47925,N_49069);
xor UO_4298 (O_4298,N_46146,N_49651);
xor UO_4299 (O_4299,N_49577,N_45893);
nand UO_4300 (O_4300,N_45745,N_45980);
and UO_4301 (O_4301,N_46102,N_45604);
nor UO_4302 (O_4302,N_47080,N_48652);
xor UO_4303 (O_4303,N_48425,N_46735);
xor UO_4304 (O_4304,N_45578,N_45595);
and UO_4305 (O_4305,N_46846,N_45738);
nand UO_4306 (O_4306,N_46097,N_45630);
or UO_4307 (O_4307,N_48393,N_47178);
nor UO_4308 (O_4308,N_49103,N_48241);
and UO_4309 (O_4309,N_47653,N_49947);
and UO_4310 (O_4310,N_47855,N_49229);
nand UO_4311 (O_4311,N_47489,N_46093);
or UO_4312 (O_4312,N_45777,N_47351);
and UO_4313 (O_4313,N_47747,N_49079);
or UO_4314 (O_4314,N_49740,N_49419);
or UO_4315 (O_4315,N_47988,N_47540);
and UO_4316 (O_4316,N_47904,N_48613);
xor UO_4317 (O_4317,N_45682,N_48517);
nand UO_4318 (O_4318,N_47872,N_47980);
nand UO_4319 (O_4319,N_49668,N_48151);
xnor UO_4320 (O_4320,N_46471,N_46300);
and UO_4321 (O_4321,N_48225,N_49674);
nor UO_4322 (O_4322,N_49715,N_49090);
nor UO_4323 (O_4323,N_48280,N_45472);
xor UO_4324 (O_4324,N_49303,N_45058);
nor UO_4325 (O_4325,N_45349,N_49491);
and UO_4326 (O_4326,N_47599,N_46171);
and UO_4327 (O_4327,N_47757,N_46367);
nor UO_4328 (O_4328,N_49640,N_45959);
and UO_4329 (O_4329,N_47095,N_46759);
xnor UO_4330 (O_4330,N_46809,N_47302);
xor UO_4331 (O_4331,N_48936,N_45135);
xnor UO_4332 (O_4332,N_46136,N_48947);
nor UO_4333 (O_4333,N_47972,N_47504);
xor UO_4334 (O_4334,N_47514,N_46427);
and UO_4335 (O_4335,N_46467,N_49248);
xor UO_4336 (O_4336,N_46055,N_46687);
nor UO_4337 (O_4337,N_45939,N_46185);
and UO_4338 (O_4338,N_49442,N_46309);
and UO_4339 (O_4339,N_47619,N_45280);
and UO_4340 (O_4340,N_45556,N_49826);
nor UO_4341 (O_4341,N_48509,N_46531);
nor UO_4342 (O_4342,N_46523,N_49373);
xnor UO_4343 (O_4343,N_45939,N_49726);
and UO_4344 (O_4344,N_49350,N_47814);
nor UO_4345 (O_4345,N_45356,N_49505);
nand UO_4346 (O_4346,N_46677,N_45558);
xnor UO_4347 (O_4347,N_48536,N_46399);
and UO_4348 (O_4348,N_45396,N_49150);
xor UO_4349 (O_4349,N_46146,N_48111);
or UO_4350 (O_4350,N_46463,N_45894);
xnor UO_4351 (O_4351,N_48339,N_45190);
nor UO_4352 (O_4352,N_45761,N_47506);
and UO_4353 (O_4353,N_48707,N_47393);
and UO_4354 (O_4354,N_45298,N_47863);
nor UO_4355 (O_4355,N_47490,N_46706);
nor UO_4356 (O_4356,N_48129,N_46737);
nand UO_4357 (O_4357,N_49734,N_46189);
nand UO_4358 (O_4358,N_48173,N_45915);
xnor UO_4359 (O_4359,N_45648,N_49031);
or UO_4360 (O_4360,N_45547,N_45503);
or UO_4361 (O_4361,N_48228,N_47897);
nand UO_4362 (O_4362,N_49446,N_47343);
or UO_4363 (O_4363,N_46327,N_48524);
or UO_4364 (O_4364,N_49261,N_47707);
nor UO_4365 (O_4365,N_47865,N_45349);
and UO_4366 (O_4366,N_46681,N_47448);
xnor UO_4367 (O_4367,N_48490,N_47323);
nand UO_4368 (O_4368,N_48136,N_46349);
nor UO_4369 (O_4369,N_47164,N_49559);
or UO_4370 (O_4370,N_46926,N_46396);
xor UO_4371 (O_4371,N_49679,N_47568);
and UO_4372 (O_4372,N_46097,N_46165);
or UO_4373 (O_4373,N_47190,N_45257);
and UO_4374 (O_4374,N_48984,N_49837);
xor UO_4375 (O_4375,N_47288,N_46530);
nor UO_4376 (O_4376,N_48630,N_45855);
nor UO_4377 (O_4377,N_46054,N_49048);
xor UO_4378 (O_4378,N_48891,N_48204);
xnor UO_4379 (O_4379,N_49337,N_48143);
and UO_4380 (O_4380,N_46824,N_49463);
nor UO_4381 (O_4381,N_49997,N_48178);
nand UO_4382 (O_4382,N_48456,N_49358);
xor UO_4383 (O_4383,N_49862,N_47810);
nand UO_4384 (O_4384,N_47983,N_46629);
xor UO_4385 (O_4385,N_49404,N_48726);
and UO_4386 (O_4386,N_47890,N_46096);
xor UO_4387 (O_4387,N_46656,N_47959);
or UO_4388 (O_4388,N_46958,N_49628);
nand UO_4389 (O_4389,N_48913,N_49453);
or UO_4390 (O_4390,N_48569,N_47426);
or UO_4391 (O_4391,N_46551,N_48317);
xor UO_4392 (O_4392,N_48591,N_45209);
or UO_4393 (O_4393,N_46766,N_45424);
nor UO_4394 (O_4394,N_46880,N_45363);
and UO_4395 (O_4395,N_47210,N_47697);
nor UO_4396 (O_4396,N_49204,N_48287);
xor UO_4397 (O_4397,N_48410,N_49695);
nor UO_4398 (O_4398,N_45197,N_48050);
nor UO_4399 (O_4399,N_47211,N_49763);
or UO_4400 (O_4400,N_48526,N_48412);
or UO_4401 (O_4401,N_45390,N_46249);
and UO_4402 (O_4402,N_47035,N_47324);
nor UO_4403 (O_4403,N_46487,N_47811);
nand UO_4404 (O_4404,N_47910,N_46447);
or UO_4405 (O_4405,N_45108,N_46122);
nor UO_4406 (O_4406,N_49374,N_48810);
xnor UO_4407 (O_4407,N_46981,N_48719);
or UO_4408 (O_4408,N_49681,N_49751);
nor UO_4409 (O_4409,N_48129,N_48160);
xnor UO_4410 (O_4410,N_48261,N_47188);
nor UO_4411 (O_4411,N_45855,N_49200);
xnor UO_4412 (O_4412,N_45232,N_45254);
nor UO_4413 (O_4413,N_47624,N_47874);
or UO_4414 (O_4414,N_45197,N_47163);
nand UO_4415 (O_4415,N_45687,N_46649);
nand UO_4416 (O_4416,N_47363,N_47046);
and UO_4417 (O_4417,N_45917,N_45939);
and UO_4418 (O_4418,N_48835,N_49141);
nand UO_4419 (O_4419,N_46810,N_46299);
and UO_4420 (O_4420,N_48804,N_47305);
xor UO_4421 (O_4421,N_45862,N_46224);
nand UO_4422 (O_4422,N_45358,N_46081);
or UO_4423 (O_4423,N_48838,N_49748);
xor UO_4424 (O_4424,N_49222,N_45861);
nor UO_4425 (O_4425,N_47890,N_47677);
and UO_4426 (O_4426,N_45427,N_49680);
or UO_4427 (O_4427,N_49269,N_45155);
nand UO_4428 (O_4428,N_49553,N_49209);
and UO_4429 (O_4429,N_45940,N_48029);
xnor UO_4430 (O_4430,N_48649,N_45992);
nand UO_4431 (O_4431,N_45936,N_48794);
and UO_4432 (O_4432,N_47466,N_49648);
nor UO_4433 (O_4433,N_47958,N_48323);
nand UO_4434 (O_4434,N_45445,N_45808);
or UO_4435 (O_4435,N_46207,N_47052);
nand UO_4436 (O_4436,N_45171,N_48964);
or UO_4437 (O_4437,N_45909,N_47420);
and UO_4438 (O_4438,N_49352,N_47421);
nor UO_4439 (O_4439,N_49170,N_48875);
nand UO_4440 (O_4440,N_47299,N_48397);
xor UO_4441 (O_4441,N_46423,N_47023);
and UO_4442 (O_4442,N_48642,N_47285);
and UO_4443 (O_4443,N_45697,N_47871);
or UO_4444 (O_4444,N_48774,N_49501);
and UO_4445 (O_4445,N_46127,N_49435);
nand UO_4446 (O_4446,N_48191,N_45104);
xor UO_4447 (O_4447,N_47578,N_46394);
nand UO_4448 (O_4448,N_45263,N_46730);
xor UO_4449 (O_4449,N_47248,N_46086);
or UO_4450 (O_4450,N_48298,N_45124);
nand UO_4451 (O_4451,N_47652,N_48607);
nor UO_4452 (O_4452,N_46896,N_48856);
or UO_4453 (O_4453,N_45176,N_49854);
or UO_4454 (O_4454,N_48877,N_47839);
and UO_4455 (O_4455,N_45977,N_48889);
and UO_4456 (O_4456,N_46234,N_47813);
and UO_4457 (O_4457,N_46473,N_49565);
xor UO_4458 (O_4458,N_45282,N_48500);
and UO_4459 (O_4459,N_49328,N_46260);
nand UO_4460 (O_4460,N_46424,N_47384);
nand UO_4461 (O_4461,N_47034,N_49136);
xnor UO_4462 (O_4462,N_48747,N_49260);
and UO_4463 (O_4463,N_49750,N_48155);
or UO_4464 (O_4464,N_47792,N_45801);
nor UO_4465 (O_4465,N_48301,N_48042);
nor UO_4466 (O_4466,N_46036,N_47545);
and UO_4467 (O_4467,N_49419,N_45748);
xor UO_4468 (O_4468,N_48689,N_46274);
nand UO_4469 (O_4469,N_47565,N_48407);
and UO_4470 (O_4470,N_45549,N_49004);
xnor UO_4471 (O_4471,N_48744,N_47088);
nor UO_4472 (O_4472,N_48549,N_48834);
xnor UO_4473 (O_4473,N_49221,N_45295);
xor UO_4474 (O_4474,N_48009,N_45235);
nor UO_4475 (O_4475,N_49701,N_46896);
xor UO_4476 (O_4476,N_45607,N_48582);
nand UO_4477 (O_4477,N_45254,N_49673);
or UO_4478 (O_4478,N_45144,N_47440);
or UO_4479 (O_4479,N_45515,N_48873);
or UO_4480 (O_4480,N_45984,N_46885);
xnor UO_4481 (O_4481,N_48997,N_46535);
nand UO_4482 (O_4482,N_46117,N_49641);
and UO_4483 (O_4483,N_49241,N_47431);
or UO_4484 (O_4484,N_48507,N_48176);
nor UO_4485 (O_4485,N_47293,N_47425);
xor UO_4486 (O_4486,N_48655,N_47015);
and UO_4487 (O_4487,N_48578,N_45057);
nor UO_4488 (O_4488,N_47727,N_46902);
and UO_4489 (O_4489,N_47391,N_46366);
and UO_4490 (O_4490,N_46540,N_47235);
xnor UO_4491 (O_4491,N_49420,N_46598);
xor UO_4492 (O_4492,N_46407,N_48721);
or UO_4493 (O_4493,N_47026,N_46326);
xor UO_4494 (O_4494,N_48027,N_46580);
nand UO_4495 (O_4495,N_46424,N_46350);
nand UO_4496 (O_4496,N_46826,N_47122);
and UO_4497 (O_4497,N_49705,N_48435);
nor UO_4498 (O_4498,N_48545,N_45697);
nand UO_4499 (O_4499,N_47198,N_48722);
nand UO_4500 (O_4500,N_48217,N_48781);
or UO_4501 (O_4501,N_48196,N_48182);
nor UO_4502 (O_4502,N_48192,N_46131);
nand UO_4503 (O_4503,N_45767,N_45881);
xnor UO_4504 (O_4504,N_45970,N_45450);
xor UO_4505 (O_4505,N_49481,N_47781);
nor UO_4506 (O_4506,N_45302,N_49870);
xnor UO_4507 (O_4507,N_45002,N_49684);
or UO_4508 (O_4508,N_49895,N_49504);
or UO_4509 (O_4509,N_45771,N_49289);
or UO_4510 (O_4510,N_47028,N_45628);
xnor UO_4511 (O_4511,N_47328,N_47627);
nand UO_4512 (O_4512,N_45036,N_47082);
and UO_4513 (O_4513,N_49524,N_47863);
or UO_4514 (O_4514,N_48183,N_45608);
nor UO_4515 (O_4515,N_45176,N_49117);
nor UO_4516 (O_4516,N_49711,N_49538);
xnor UO_4517 (O_4517,N_45723,N_47375);
or UO_4518 (O_4518,N_47999,N_47946);
nand UO_4519 (O_4519,N_45721,N_48909);
or UO_4520 (O_4520,N_45659,N_49637);
xnor UO_4521 (O_4521,N_49853,N_48048);
nor UO_4522 (O_4522,N_45603,N_46050);
nor UO_4523 (O_4523,N_46609,N_45678);
and UO_4524 (O_4524,N_45280,N_47657);
or UO_4525 (O_4525,N_45386,N_47091);
and UO_4526 (O_4526,N_46430,N_45481);
or UO_4527 (O_4527,N_46424,N_47660);
or UO_4528 (O_4528,N_46664,N_48229);
and UO_4529 (O_4529,N_45578,N_49483);
xnor UO_4530 (O_4530,N_49773,N_49633);
nand UO_4531 (O_4531,N_48474,N_45697);
nor UO_4532 (O_4532,N_45304,N_45642);
and UO_4533 (O_4533,N_47945,N_47301);
and UO_4534 (O_4534,N_47673,N_46958);
or UO_4535 (O_4535,N_49355,N_49654);
and UO_4536 (O_4536,N_47452,N_48144);
xnor UO_4537 (O_4537,N_47149,N_45182);
xnor UO_4538 (O_4538,N_47387,N_46087);
and UO_4539 (O_4539,N_46180,N_48394);
nand UO_4540 (O_4540,N_45794,N_46154);
nand UO_4541 (O_4541,N_46840,N_46480);
xor UO_4542 (O_4542,N_46130,N_46163);
nand UO_4543 (O_4543,N_46744,N_48073);
nand UO_4544 (O_4544,N_45690,N_48421);
or UO_4545 (O_4545,N_46861,N_45476);
or UO_4546 (O_4546,N_48147,N_48645);
and UO_4547 (O_4547,N_49209,N_45452);
xor UO_4548 (O_4548,N_46383,N_49808);
and UO_4549 (O_4549,N_47186,N_48626);
xnor UO_4550 (O_4550,N_46711,N_49326);
nand UO_4551 (O_4551,N_49956,N_46311);
nand UO_4552 (O_4552,N_47151,N_48962);
xor UO_4553 (O_4553,N_45518,N_48522);
nand UO_4554 (O_4554,N_47307,N_49996);
xnor UO_4555 (O_4555,N_48416,N_48411);
nor UO_4556 (O_4556,N_47663,N_45627);
or UO_4557 (O_4557,N_45780,N_47649);
or UO_4558 (O_4558,N_45929,N_47231);
nand UO_4559 (O_4559,N_46667,N_46764);
nor UO_4560 (O_4560,N_48593,N_49837);
and UO_4561 (O_4561,N_45461,N_47150);
nand UO_4562 (O_4562,N_49206,N_45129);
xnor UO_4563 (O_4563,N_49928,N_45762);
nor UO_4564 (O_4564,N_48563,N_47574);
nor UO_4565 (O_4565,N_45046,N_47247);
nor UO_4566 (O_4566,N_48828,N_46722);
xor UO_4567 (O_4567,N_48341,N_48024);
and UO_4568 (O_4568,N_47416,N_48877);
xor UO_4569 (O_4569,N_49281,N_45969);
nor UO_4570 (O_4570,N_49701,N_45817);
nand UO_4571 (O_4571,N_48549,N_47968);
or UO_4572 (O_4572,N_46777,N_47148);
or UO_4573 (O_4573,N_45364,N_49500);
nor UO_4574 (O_4574,N_49930,N_49434);
nor UO_4575 (O_4575,N_47402,N_46892);
nor UO_4576 (O_4576,N_49009,N_48636);
or UO_4577 (O_4577,N_49138,N_49160);
or UO_4578 (O_4578,N_45221,N_47507);
or UO_4579 (O_4579,N_45621,N_47506);
nand UO_4580 (O_4580,N_49864,N_48440);
or UO_4581 (O_4581,N_45126,N_48912);
or UO_4582 (O_4582,N_49714,N_49272);
xor UO_4583 (O_4583,N_46677,N_49816);
and UO_4584 (O_4584,N_46516,N_45944);
and UO_4585 (O_4585,N_48391,N_46858);
or UO_4586 (O_4586,N_47874,N_45717);
and UO_4587 (O_4587,N_49877,N_48533);
nand UO_4588 (O_4588,N_45240,N_49716);
nand UO_4589 (O_4589,N_48977,N_46954);
nor UO_4590 (O_4590,N_49390,N_48589);
xnor UO_4591 (O_4591,N_47823,N_47983);
and UO_4592 (O_4592,N_45308,N_48935);
and UO_4593 (O_4593,N_45473,N_47845);
nor UO_4594 (O_4594,N_45104,N_46253);
nand UO_4595 (O_4595,N_48559,N_47117);
or UO_4596 (O_4596,N_48853,N_46331);
or UO_4597 (O_4597,N_46602,N_45138);
or UO_4598 (O_4598,N_49692,N_46007);
nor UO_4599 (O_4599,N_48695,N_48761);
xnor UO_4600 (O_4600,N_46737,N_45520);
nand UO_4601 (O_4601,N_48517,N_46175);
nand UO_4602 (O_4602,N_46249,N_46914);
or UO_4603 (O_4603,N_45706,N_46343);
or UO_4604 (O_4604,N_47235,N_49683);
and UO_4605 (O_4605,N_45647,N_48134);
nand UO_4606 (O_4606,N_48221,N_47723);
or UO_4607 (O_4607,N_48820,N_46505);
xor UO_4608 (O_4608,N_46631,N_45856);
xnor UO_4609 (O_4609,N_47394,N_45257);
nor UO_4610 (O_4610,N_49082,N_45540);
nor UO_4611 (O_4611,N_45911,N_47689);
nand UO_4612 (O_4612,N_48144,N_45165);
nor UO_4613 (O_4613,N_46939,N_49673);
xor UO_4614 (O_4614,N_49306,N_49009);
and UO_4615 (O_4615,N_45315,N_49416);
or UO_4616 (O_4616,N_48344,N_47038);
nand UO_4617 (O_4617,N_47861,N_47638);
nand UO_4618 (O_4618,N_49269,N_45541);
nand UO_4619 (O_4619,N_48793,N_46699);
xor UO_4620 (O_4620,N_47791,N_48308);
or UO_4621 (O_4621,N_45555,N_48837);
or UO_4622 (O_4622,N_49725,N_46702);
nand UO_4623 (O_4623,N_48156,N_49289);
xor UO_4624 (O_4624,N_46318,N_49924);
nor UO_4625 (O_4625,N_47453,N_49778);
and UO_4626 (O_4626,N_46064,N_48430);
xnor UO_4627 (O_4627,N_45585,N_47837);
and UO_4628 (O_4628,N_47514,N_48343);
nand UO_4629 (O_4629,N_46357,N_49571);
and UO_4630 (O_4630,N_47259,N_46260);
nand UO_4631 (O_4631,N_45827,N_45990);
nand UO_4632 (O_4632,N_48690,N_45762);
xor UO_4633 (O_4633,N_49342,N_47134);
and UO_4634 (O_4634,N_46198,N_45067);
nand UO_4635 (O_4635,N_47088,N_48787);
xnor UO_4636 (O_4636,N_47370,N_48901);
nor UO_4637 (O_4637,N_48307,N_45662);
nand UO_4638 (O_4638,N_47202,N_47395);
or UO_4639 (O_4639,N_47605,N_49984);
xor UO_4640 (O_4640,N_46895,N_46816);
nand UO_4641 (O_4641,N_46993,N_47423);
and UO_4642 (O_4642,N_45389,N_48468);
or UO_4643 (O_4643,N_45420,N_46222);
or UO_4644 (O_4644,N_45985,N_49736);
and UO_4645 (O_4645,N_48030,N_48484);
xor UO_4646 (O_4646,N_48372,N_49088);
and UO_4647 (O_4647,N_45342,N_49294);
xnor UO_4648 (O_4648,N_49150,N_45559);
and UO_4649 (O_4649,N_49003,N_49019);
or UO_4650 (O_4650,N_47099,N_49391);
xor UO_4651 (O_4651,N_49555,N_48795);
or UO_4652 (O_4652,N_48271,N_45884);
and UO_4653 (O_4653,N_48515,N_48120);
xor UO_4654 (O_4654,N_45982,N_47894);
xor UO_4655 (O_4655,N_46342,N_46928);
nand UO_4656 (O_4656,N_48003,N_48558);
and UO_4657 (O_4657,N_49706,N_47568);
xnor UO_4658 (O_4658,N_48639,N_48771);
and UO_4659 (O_4659,N_48233,N_46821);
nor UO_4660 (O_4660,N_48628,N_46045);
xnor UO_4661 (O_4661,N_47858,N_49521);
and UO_4662 (O_4662,N_49045,N_48067);
nor UO_4663 (O_4663,N_47597,N_46335);
and UO_4664 (O_4664,N_45053,N_47383);
nor UO_4665 (O_4665,N_45500,N_45991);
nand UO_4666 (O_4666,N_49144,N_49758);
or UO_4667 (O_4667,N_45739,N_49314);
or UO_4668 (O_4668,N_46233,N_48913);
or UO_4669 (O_4669,N_45723,N_48458);
xnor UO_4670 (O_4670,N_48914,N_46189);
and UO_4671 (O_4671,N_45311,N_47308);
and UO_4672 (O_4672,N_49745,N_49925);
xor UO_4673 (O_4673,N_48753,N_46931);
or UO_4674 (O_4674,N_49798,N_48112);
xor UO_4675 (O_4675,N_49918,N_47696);
or UO_4676 (O_4676,N_48621,N_46435);
nor UO_4677 (O_4677,N_47850,N_45315);
nand UO_4678 (O_4678,N_46018,N_47936);
nor UO_4679 (O_4679,N_49803,N_46870);
nor UO_4680 (O_4680,N_47519,N_45345);
nand UO_4681 (O_4681,N_47050,N_46680);
nor UO_4682 (O_4682,N_47271,N_49656);
xnor UO_4683 (O_4683,N_48160,N_45914);
xor UO_4684 (O_4684,N_46624,N_46356);
xnor UO_4685 (O_4685,N_47133,N_45339);
xor UO_4686 (O_4686,N_45729,N_49549);
nor UO_4687 (O_4687,N_49738,N_48803);
and UO_4688 (O_4688,N_45569,N_45286);
or UO_4689 (O_4689,N_46343,N_46339);
xnor UO_4690 (O_4690,N_46742,N_47900);
nand UO_4691 (O_4691,N_46093,N_49831);
and UO_4692 (O_4692,N_48656,N_49854);
nand UO_4693 (O_4693,N_48353,N_45473);
and UO_4694 (O_4694,N_46695,N_46611);
nand UO_4695 (O_4695,N_48104,N_48879);
xnor UO_4696 (O_4696,N_47745,N_45464);
xnor UO_4697 (O_4697,N_46307,N_47016);
nor UO_4698 (O_4698,N_45673,N_48981);
xnor UO_4699 (O_4699,N_47758,N_45922);
or UO_4700 (O_4700,N_47913,N_48928);
nand UO_4701 (O_4701,N_48013,N_49869);
or UO_4702 (O_4702,N_46616,N_47223);
or UO_4703 (O_4703,N_46776,N_46259);
or UO_4704 (O_4704,N_49623,N_49566);
or UO_4705 (O_4705,N_46428,N_49123);
nor UO_4706 (O_4706,N_46696,N_45201);
or UO_4707 (O_4707,N_47255,N_45399);
and UO_4708 (O_4708,N_47908,N_46676);
nor UO_4709 (O_4709,N_48603,N_47139);
nand UO_4710 (O_4710,N_46472,N_48032);
nand UO_4711 (O_4711,N_47263,N_48201);
xnor UO_4712 (O_4712,N_46279,N_45561);
xnor UO_4713 (O_4713,N_47263,N_45073);
nand UO_4714 (O_4714,N_49339,N_45655);
and UO_4715 (O_4715,N_49911,N_45177);
and UO_4716 (O_4716,N_46338,N_47832);
and UO_4717 (O_4717,N_46646,N_48966);
and UO_4718 (O_4718,N_45019,N_49122);
nand UO_4719 (O_4719,N_46170,N_46313);
or UO_4720 (O_4720,N_47749,N_47547);
nor UO_4721 (O_4721,N_46821,N_47301);
and UO_4722 (O_4722,N_47734,N_47142);
nor UO_4723 (O_4723,N_48801,N_45728);
xnor UO_4724 (O_4724,N_47349,N_45187);
nand UO_4725 (O_4725,N_48364,N_49863);
nand UO_4726 (O_4726,N_47733,N_48864);
or UO_4727 (O_4727,N_45856,N_46174);
xnor UO_4728 (O_4728,N_45125,N_47467);
and UO_4729 (O_4729,N_46225,N_47107);
or UO_4730 (O_4730,N_45645,N_48963);
nand UO_4731 (O_4731,N_47610,N_45653);
or UO_4732 (O_4732,N_49196,N_46242);
or UO_4733 (O_4733,N_46266,N_45228);
nand UO_4734 (O_4734,N_45861,N_48872);
and UO_4735 (O_4735,N_47977,N_46138);
nand UO_4736 (O_4736,N_47980,N_46512);
nor UO_4737 (O_4737,N_48164,N_49010);
nand UO_4738 (O_4738,N_45540,N_47800);
nor UO_4739 (O_4739,N_48806,N_47146);
nor UO_4740 (O_4740,N_47591,N_48713);
xor UO_4741 (O_4741,N_45588,N_46309);
nand UO_4742 (O_4742,N_49854,N_48790);
nor UO_4743 (O_4743,N_46225,N_46251);
nand UO_4744 (O_4744,N_45716,N_49982);
nor UO_4745 (O_4745,N_49465,N_46358);
nand UO_4746 (O_4746,N_47427,N_46602);
xnor UO_4747 (O_4747,N_45867,N_47422);
and UO_4748 (O_4748,N_46104,N_49237);
nor UO_4749 (O_4749,N_47208,N_49075);
nor UO_4750 (O_4750,N_48412,N_46131);
or UO_4751 (O_4751,N_48590,N_46801);
or UO_4752 (O_4752,N_45942,N_46870);
nand UO_4753 (O_4753,N_48498,N_49239);
nor UO_4754 (O_4754,N_47996,N_46154);
nor UO_4755 (O_4755,N_45121,N_47024);
or UO_4756 (O_4756,N_47442,N_47833);
or UO_4757 (O_4757,N_47496,N_49641);
or UO_4758 (O_4758,N_47756,N_47655);
xor UO_4759 (O_4759,N_45128,N_47569);
and UO_4760 (O_4760,N_46980,N_48571);
nor UO_4761 (O_4761,N_46330,N_47059);
or UO_4762 (O_4762,N_46147,N_47926);
xor UO_4763 (O_4763,N_45499,N_48424);
and UO_4764 (O_4764,N_45738,N_46844);
nor UO_4765 (O_4765,N_45740,N_49250);
and UO_4766 (O_4766,N_46524,N_46729);
nor UO_4767 (O_4767,N_48071,N_46252);
and UO_4768 (O_4768,N_49885,N_47389);
nor UO_4769 (O_4769,N_45405,N_46380);
nor UO_4770 (O_4770,N_46759,N_49536);
xnor UO_4771 (O_4771,N_49995,N_47972);
and UO_4772 (O_4772,N_46076,N_46650);
and UO_4773 (O_4773,N_45307,N_48862);
and UO_4774 (O_4774,N_45223,N_48548);
xor UO_4775 (O_4775,N_45896,N_46062);
nand UO_4776 (O_4776,N_46233,N_46936);
or UO_4777 (O_4777,N_48794,N_47124);
nand UO_4778 (O_4778,N_45495,N_45456);
nor UO_4779 (O_4779,N_49768,N_46293);
nor UO_4780 (O_4780,N_46425,N_46287);
xnor UO_4781 (O_4781,N_46262,N_47455);
xnor UO_4782 (O_4782,N_48613,N_48353);
and UO_4783 (O_4783,N_49777,N_45592);
or UO_4784 (O_4784,N_49021,N_49345);
and UO_4785 (O_4785,N_47986,N_45745);
xor UO_4786 (O_4786,N_47313,N_48871);
and UO_4787 (O_4787,N_45285,N_49073);
nand UO_4788 (O_4788,N_46102,N_48659);
or UO_4789 (O_4789,N_47316,N_48371);
xor UO_4790 (O_4790,N_47799,N_48175);
and UO_4791 (O_4791,N_46674,N_45486);
nor UO_4792 (O_4792,N_49076,N_49274);
nand UO_4793 (O_4793,N_47978,N_48213);
nor UO_4794 (O_4794,N_45727,N_46378);
nand UO_4795 (O_4795,N_45853,N_46623);
and UO_4796 (O_4796,N_49308,N_46689);
nor UO_4797 (O_4797,N_48633,N_47856);
nor UO_4798 (O_4798,N_46274,N_45519);
and UO_4799 (O_4799,N_49707,N_47544);
xor UO_4800 (O_4800,N_45586,N_48706);
nor UO_4801 (O_4801,N_45002,N_47874);
nor UO_4802 (O_4802,N_45331,N_48382);
xor UO_4803 (O_4803,N_49529,N_46967);
xnor UO_4804 (O_4804,N_47043,N_48701);
xor UO_4805 (O_4805,N_49931,N_48692);
and UO_4806 (O_4806,N_45320,N_45816);
nand UO_4807 (O_4807,N_47821,N_47656);
nand UO_4808 (O_4808,N_46823,N_46133);
nand UO_4809 (O_4809,N_49993,N_47122);
and UO_4810 (O_4810,N_45478,N_46654);
and UO_4811 (O_4811,N_49117,N_49579);
xnor UO_4812 (O_4812,N_46273,N_47892);
nor UO_4813 (O_4813,N_48840,N_49171);
nor UO_4814 (O_4814,N_47663,N_46043);
or UO_4815 (O_4815,N_49739,N_45903);
and UO_4816 (O_4816,N_49119,N_48901);
or UO_4817 (O_4817,N_48759,N_48063);
nand UO_4818 (O_4818,N_45872,N_49717);
xnor UO_4819 (O_4819,N_48238,N_46683);
and UO_4820 (O_4820,N_45500,N_47225);
and UO_4821 (O_4821,N_45708,N_49388);
or UO_4822 (O_4822,N_48367,N_47927);
nand UO_4823 (O_4823,N_49278,N_47288);
and UO_4824 (O_4824,N_45291,N_46041);
nor UO_4825 (O_4825,N_47089,N_46365);
or UO_4826 (O_4826,N_45276,N_46608);
nand UO_4827 (O_4827,N_45816,N_49695);
or UO_4828 (O_4828,N_45875,N_47849);
and UO_4829 (O_4829,N_47472,N_48536);
xor UO_4830 (O_4830,N_46564,N_45284);
xor UO_4831 (O_4831,N_45194,N_46802);
xor UO_4832 (O_4832,N_46290,N_46580);
nor UO_4833 (O_4833,N_49532,N_45973);
and UO_4834 (O_4834,N_45611,N_49335);
or UO_4835 (O_4835,N_49616,N_45553);
nor UO_4836 (O_4836,N_48913,N_49504);
or UO_4837 (O_4837,N_46762,N_48953);
xor UO_4838 (O_4838,N_45752,N_47400);
nand UO_4839 (O_4839,N_45834,N_49150);
xor UO_4840 (O_4840,N_48176,N_49750);
xor UO_4841 (O_4841,N_48531,N_47845);
nand UO_4842 (O_4842,N_45644,N_45057);
xor UO_4843 (O_4843,N_49288,N_49535);
or UO_4844 (O_4844,N_46671,N_46350);
and UO_4845 (O_4845,N_46813,N_46843);
or UO_4846 (O_4846,N_47622,N_49374);
nand UO_4847 (O_4847,N_46244,N_45500);
nor UO_4848 (O_4848,N_47992,N_45322);
xnor UO_4849 (O_4849,N_48261,N_47424);
xor UO_4850 (O_4850,N_46762,N_47109);
xor UO_4851 (O_4851,N_49991,N_48120);
xnor UO_4852 (O_4852,N_45864,N_48972);
nor UO_4853 (O_4853,N_49025,N_45925);
xor UO_4854 (O_4854,N_49011,N_46862);
nand UO_4855 (O_4855,N_45102,N_48683);
nor UO_4856 (O_4856,N_47229,N_48831);
nand UO_4857 (O_4857,N_45118,N_49859);
nand UO_4858 (O_4858,N_46674,N_45696);
or UO_4859 (O_4859,N_45388,N_47525);
nor UO_4860 (O_4860,N_49975,N_49207);
xor UO_4861 (O_4861,N_49376,N_48420);
xor UO_4862 (O_4862,N_45260,N_49998);
xnor UO_4863 (O_4863,N_47248,N_45515);
xor UO_4864 (O_4864,N_48350,N_49883);
or UO_4865 (O_4865,N_48067,N_45827);
nand UO_4866 (O_4866,N_46992,N_47396);
nor UO_4867 (O_4867,N_45470,N_45353);
or UO_4868 (O_4868,N_46133,N_46328);
nand UO_4869 (O_4869,N_46200,N_49430);
xnor UO_4870 (O_4870,N_49052,N_45475);
nand UO_4871 (O_4871,N_49704,N_46380);
nand UO_4872 (O_4872,N_47586,N_45233);
nor UO_4873 (O_4873,N_49847,N_46544);
nor UO_4874 (O_4874,N_45697,N_47703);
or UO_4875 (O_4875,N_47968,N_46278);
or UO_4876 (O_4876,N_48549,N_47425);
xor UO_4877 (O_4877,N_47417,N_49937);
nand UO_4878 (O_4878,N_49648,N_47397);
nor UO_4879 (O_4879,N_46217,N_49047);
xnor UO_4880 (O_4880,N_45682,N_46585);
nor UO_4881 (O_4881,N_45453,N_48843);
and UO_4882 (O_4882,N_45225,N_47276);
or UO_4883 (O_4883,N_48177,N_47138);
and UO_4884 (O_4884,N_45103,N_45253);
or UO_4885 (O_4885,N_46309,N_46277);
or UO_4886 (O_4886,N_49391,N_47657);
nand UO_4887 (O_4887,N_49947,N_47827);
or UO_4888 (O_4888,N_45309,N_47243);
nor UO_4889 (O_4889,N_45619,N_48997);
nand UO_4890 (O_4890,N_46722,N_47806);
nand UO_4891 (O_4891,N_47646,N_47208);
and UO_4892 (O_4892,N_49606,N_46971);
or UO_4893 (O_4893,N_45235,N_45568);
or UO_4894 (O_4894,N_47755,N_45314);
or UO_4895 (O_4895,N_47202,N_46949);
xnor UO_4896 (O_4896,N_45543,N_46432);
nor UO_4897 (O_4897,N_47360,N_48554);
nor UO_4898 (O_4898,N_47095,N_45071);
nand UO_4899 (O_4899,N_46194,N_47171);
nor UO_4900 (O_4900,N_46852,N_48460);
xor UO_4901 (O_4901,N_45941,N_49478);
nand UO_4902 (O_4902,N_49664,N_47703);
nand UO_4903 (O_4903,N_45173,N_46801);
nand UO_4904 (O_4904,N_46647,N_45298);
nor UO_4905 (O_4905,N_46637,N_46288);
and UO_4906 (O_4906,N_49424,N_49007);
xor UO_4907 (O_4907,N_49296,N_47630);
xor UO_4908 (O_4908,N_46412,N_49112);
nand UO_4909 (O_4909,N_45440,N_48786);
nor UO_4910 (O_4910,N_48863,N_46004);
xor UO_4911 (O_4911,N_47258,N_45350);
nor UO_4912 (O_4912,N_49938,N_46418);
nor UO_4913 (O_4913,N_45775,N_49875);
and UO_4914 (O_4914,N_49153,N_49462);
and UO_4915 (O_4915,N_45456,N_45290);
and UO_4916 (O_4916,N_47988,N_49842);
nand UO_4917 (O_4917,N_49884,N_49213);
nand UO_4918 (O_4918,N_48180,N_45291);
nor UO_4919 (O_4919,N_45774,N_49635);
and UO_4920 (O_4920,N_46702,N_45404);
and UO_4921 (O_4921,N_47022,N_49945);
and UO_4922 (O_4922,N_47257,N_48533);
xor UO_4923 (O_4923,N_46391,N_45521);
nor UO_4924 (O_4924,N_46785,N_47106);
nor UO_4925 (O_4925,N_47080,N_46305);
and UO_4926 (O_4926,N_49709,N_46385);
and UO_4927 (O_4927,N_48006,N_49718);
nand UO_4928 (O_4928,N_49706,N_45505);
xor UO_4929 (O_4929,N_45707,N_48059);
xnor UO_4930 (O_4930,N_47505,N_49190);
or UO_4931 (O_4931,N_45756,N_46765);
nand UO_4932 (O_4932,N_46434,N_45036);
nor UO_4933 (O_4933,N_48781,N_46228);
and UO_4934 (O_4934,N_48350,N_48116);
nor UO_4935 (O_4935,N_49643,N_48281);
xor UO_4936 (O_4936,N_47915,N_47497);
xor UO_4937 (O_4937,N_45501,N_48226);
or UO_4938 (O_4938,N_45735,N_48513);
nand UO_4939 (O_4939,N_49645,N_45291);
nand UO_4940 (O_4940,N_46277,N_46230);
nand UO_4941 (O_4941,N_46356,N_46436);
and UO_4942 (O_4942,N_49298,N_45035);
or UO_4943 (O_4943,N_49044,N_46182);
xnor UO_4944 (O_4944,N_46016,N_47788);
nand UO_4945 (O_4945,N_45475,N_45246);
nor UO_4946 (O_4946,N_47891,N_48863);
or UO_4947 (O_4947,N_45835,N_47192);
nor UO_4948 (O_4948,N_48309,N_45044);
nand UO_4949 (O_4949,N_45720,N_48389);
nand UO_4950 (O_4950,N_48899,N_47403);
nor UO_4951 (O_4951,N_45769,N_47922);
xnor UO_4952 (O_4952,N_46485,N_46994);
nor UO_4953 (O_4953,N_49681,N_49000);
or UO_4954 (O_4954,N_45721,N_47241);
xnor UO_4955 (O_4955,N_45157,N_45782);
nand UO_4956 (O_4956,N_46266,N_48523);
nor UO_4957 (O_4957,N_46600,N_49821);
nand UO_4958 (O_4958,N_46941,N_47017);
nor UO_4959 (O_4959,N_48248,N_46282);
or UO_4960 (O_4960,N_48574,N_46105);
xnor UO_4961 (O_4961,N_45887,N_49355);
nor UO_4962 (O_4962,N_46019,N_45648);
or UO_4963 (O_4963,N_47454,N_46608);
xor UO_4964 (O_4964,N_48000,N_48666);
or UO_4965 (O_4965,N_49701,N_46188);
and UO_4966 (O_4966,N_45291,N_49751);
or UO_4967 (O_4967,N_47445,N_45921);
nor UO_4968 (O_4968,N_45006,N_45108);
nand UO_4969 (O_4969,N_46807,N_49873);
or UO_4970 (O_4970,N_47878,N_48995);
or UO_4971 (O_4971,N_49220,N_46793);
xor UO_4972 (O_4972,N_45658,N_47857);
or UO_4973 (O_4973,N_45462,N_49166);
nand UO_4974 (O_4974,N_45460,N_45633);
and UO_4975 (O_4975,N_47212,N_45349);
nand UO_4976 (O_4976,N_46169,N_48828);
or UO_4977 (O_4977,N_46348,N_46833);
nand UO_4978 (O_4978,N_47739,N_46365);
and UO_4979 (O_4979,N_45678,N_45436);
and UO_4980 (O_4980,N_46872,N_46369);
or UO_4981 (O_4981,N_45543,N_46221);
xor UO_4982 (O_4982,N_49196,N_46262);
xnor UO_4983 (O_4983,N_47381,N_48802);
nand UO_4984 (O_4984,N_49697,N_45450);
or UO_4985 (O_4985,N_48993,N_46022);
nand UO_4986 (O_4986,N_45270,N_46429);
nor UO_4987 (O_4987,N_47713,N_49594);
nor UO_4988 (O_4988,N_45278,N_48425);
nand UO_4989 (O_4989,N_47597,N_45284);
nand UO_4990 (O_4990,N_45593,N_46163);
or UO_4991 (O_4991,N_48644,N_47502);
nand UO_4992 (O_4992,N_47442,N_48905);
nand UO_4993 (O_4993,N_48975,N_47862);
xnor UO_4994 (O_4994,N_49586,N_47207);
xor UO_4995 (O_4995,N_48418,N_47034);
and UO_4996 (O_4996,N_47301,N_48356);
xor UO_4997 (O_4997,N_46456,N_46119);
or UO_4998 (O_4998,N_49613,N_47656);
or UO_4999 (O_4999,N_46549,N_49396);
endmodule