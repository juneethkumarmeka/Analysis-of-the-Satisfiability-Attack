module basic_500_3000_500_50_levels_2xor_5(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_299,In_184);
nor U1 (N_1,In_282,In_131);
xor U2 (N_2,In_170,In_175);
nand U3 (N_3,In_205,In_154);
nor U4 (N_4,In_408,In_393);
or U5 (N_5,In_104,In_114);
xor U6 (N_6,In_49,In_452);
nand U7 (N_7,In_371,In_169);
nor U8 (N_8,In_345,In_223);
and U9 (N_9,In_409,In_117);
nor U10 (N_10,In_256,In_171);
and U11 (N_11,In_362,In_168);
and U12 (N_12,In_332,In_124);
and U13 (N_13,In_304,In_241);
nand U14 (N_14,In_251,In_116);
nor U15 (N_15,In_0,In_340);
nor U16 (N_16,In_388,In_9);
nor U17 (N_17,In_59,In_469);
or U18 (N_18,In_481,In_375);
and U19 (N_19,In_410,In_158);
and U20 (N_20,In_461,In_193);
nand U21 (N_21,In_492,In_383);
nand U22 (N_22,In_425,In_109);
nand U23 (N_23,In_139,In_25);
and U24 (N_24,In_123,In_152);
nand U25 (N_25,In_378,In_216);
nor U26 (N_26,In_192,In_298);
and U27 (N_27,In_384,In_83);
nor U28 (N_28,In_314,In_398);
xor U29 (N_29,In_140,In_277);
or U30 (N_30,In_99,In_15);
or U31 (N_31,In_329,In_115);
or U32 (N_32,In_392,In_402);
or U33 (N_33,In_18,In_111);
nand U34 (N_34,In_422,In_146);
and U35 (N_35,In_235,In_143);
or U36 (N_36,In_27,In_206);
and U37 (N_37,In_194,In_188);
nand U38 (N_38,In_217,In_215);
and U39 (N_39,In_403,In_73);
and U40 (N_40,In_268,In_394);
nand U41 (N_41,In_488,In_252);
or U42 (N_42,In_428,In_407);
or U43 (N_43,In_162,In_261);
or U44 (N_44,In_87,In_13);
nor U45 (N_45,In_301,In_76);
nand U46 (N_46,In_197,In_432);
and U47 (N_47,In_58,In_225);
nand U48 (N_48,In_23,In_210);
or U49 (N_49,In_368,In_449);
nor U50 (N_50,In_453,In_334);
nor U51 (N_51,In_204,In_322);
nor U52 (N_52,In_270,In_212);
nor U53 (N_53,In_344,In_434);
and U54 (N_54,In_433,In_233);
nor U55 (N_55,In_475,In_476);
or U56 (N_56,In_191,In_380);
or U57 (N_57,In_455,In_498);
nand U58 (N_58,In_260,In_63);
xnor U59 (N_59,In_75,In_265);
and U60 (N_60,In_182,In_283);
nor U61 (N_61,In_259,In_324);
nor U62 (N_62,In_36,In_42);
nand U63 (N_63,In_89,In_55);
or U64 (N_64,N_0,In_133);
and U65 (N_65,In_292,In_198);
xnor U66 (N_66,In_451,In_122);
and U67 (N_67,In_77,In_138);
nand U68 (N_68,N_32,In_226);
nand U69 (N_69,In_207,In_155);
nor U70 (N_70,In_297,In_424);
or U71 (N_71,In_132,In_397);
nor U72 (N_72,In_303,In_352);
or U73 (N_73,In_401,In_468);
and U74 (N_74,In_406,In_39);
and U75 (N_75,In_148,In_462);
or U76 (N_76,In_343,In_160);
nor U77 (N_77,In_463,In_134);
nand U78 (N_78,In_214,In_437);
and U79 (N_79,N_31,In_423);
nor U80 (N_80,In_336,In_325);
nand U81 (N_81,In_32,In_163);
nor U82 (N_82,In_319,In_350);
nand U83 (N_83,N_18,In_120);
nand U84 (N_84,In_306,N_21);
and U85 (N_85,In_6,In_430);
or U86 (N_86,In_126,In_12);
nand U87 (N_87,In_480,In_370);
or U88 (N_88,In_274,In_186);
nand U89 (N_89,In_263,In_14);
nor U90 (N_90,In_113,In_189);
nand U91 (N_91,In_180,In_8);
nand U92 (N_92,N_25,In_312);
or U93 (N_93,In_108,In_68);
or U94 (N_94,In_470,In_67);
and U95 (N_95,In_22,In_473);
nand U96 (N_96,In_105,In_267);
or U97 (N_97,In_454,In_436);
and U98 (N_98,In_272,In_294);
nor U99 (N_99,In_440,In_258);
nor U100 (N_100,In_183,In_474);
nor U101 (N_101,In_240,In_78);
or U102 (N_102,N_23,N_39);
and U103 (N_103,In_295,N_19);
nand U104 (N_104,In_17,In_356);
nand U105 (N_105,N_6,In_330);
nor U106 (N_106,In_415,In_245);
nor U107 (N_107,In_307,In_196);
and U108 (N_108,In_444,In_429);
nor U109 (N_109,In_101,In_358);
nand U110 (N_110,In_201,In_121);
or U111 (N_111,In_174,In_351);
nor U112 (N_112,In_244,In_3);
and U113 (N_113,In_161,In_151);
or U114 (N_114,In_46,In_485);
or U115 (N_115,In_222,In_489);
nand U116 (N_116,In_467,In_157);
or U117 (N_117,In_478,In_385);
nor U118 (N_118,N_58,In_218);
and U119 (N_119,In_271,In_30);
nand U120 (N_120,In_70,In_296);
nand U121 (N_121,N_65,N_10);
and U122 (N_122,N_49,N_108);
and U123 (N_123,In_34,In_493);
nand U124 (N_124,In_365,In_56);
and U125 (N_125,N_67,In_439);
xor U126 (N_126,In_106,In_1);
nor U127 (N_127,In_419,In_276);
nand U128 (N_128,In_484,In_400);
xor U129 (N_129,In_107,In_369);
or U130 (N_130,N_2,In_302);
or U131 (N_131,In_389,In_82);
nand U132 (N_132,In_231,In_311);
and U133 (N_133,In_141,N_61);
and U134 (N_134,N_27,In_29);
nand U135 (N_135,N_41,N_35);
or U136 (N_136,In_363,In_327);
and U137 (N_137,N_79,In_497);
and U138 (N_138,In_220,N_97);
or U139 (N_139,In_24,In_458);
nand U140 (N_140,In_127,In_179);
and U141 (N_141,In_257,N_66);
or U142 (N_142,In_224,In_457);
and U143 (N_143,N_26,In_293);
nand U144 (N_144,N_75,N_63);
xnor U145 (N_145,In_431,In_128);
and U146 (N_146,In_208,In_448);
or U147 (N_147,In_234,In_167);
or U148 (N_148,In_178,In_328);
xnor U149 (N_149,N_106,In_487);
or U150 (N_150,In_405,In_66);
xor U151 (N_151,In_95,In_426);
and U152 (N_152,In_118,In_313);
or U153 (N_153,N_107,In_339);
or U154 (N_154,N_17,In_79);
nand U155 (N_155,In_264,N_99);
or U156 (N_156,N_55,In_435);
nor U157 (N_157,N_76,N_93);
nand U158 (N_158,In_442,In_239);
or U159 (N_159,In_181,In_382);
nor U160 (N_160,N_83,In_377);
and U161 (N_161,In_399,N_101);
nor U162 (N_162,In_237,N_29);
and U163 (N_163,In_346,In_69);
nor U164 (N_164,In_414,In_96);
nor U165 (N_165,N_50,In_202);
and U166 (N_166,In_4,In_418);
nor U167 (N_167,In_387,N_37);
nor U168 (N_168,In_413,In_137);
nand U169 (N_169,In_65,In_166);
and U170 (N_170,N_104,In_471);
nor U171 (N_171,N_16,In_43);
and U172 (N_172,In_135,N_62);
nand U173 (N_173,In_342,In_52);
xor U174 (N_174,In_173,In_374);
nand U175 (N_175,In_421,N_46);
nand U176 (N_176,N_68,N_7);
nand U177 (N_177,N_70,In_150);
or U178 (N_178,In_280,In_472);
nand U179 (N_179,In_486,In_110);
and U180 (N_180,N_53,In_255);
or U181 (N_181,In_71,In_200);
and U182 (N_182,N_116,N_12);
and U183 (N_183,In_284,N_144);
nand U184 (N_184,In_367,In_496);
or U185 (N_185,N_56,In_273);
nand U186 (N_186,N_81,In_427);
nand U187 (N_187,In_2,N_168);
nor U188 (N_188,N_91,In_228);
nand U189 (N_189,N_153,In_85);
and U190 (N_190,In_102,In_159);
and U191 (N_191,N_114,In_386);
or U192 (N_192,N_117,N_90);
nand U193 (N_193,In_411,In_112);
nand U194 (N_194,N_176,N_8);
nand U195 (N_195,In_381,In_278);
nor U196 (N_196,In_335,In_460);
or U197 (N_197,In_144,N_177);
nand U198 (N_198,In_221,N_159);
or U199 (N_199,In_262,In_53);
nand U200 (N_200,In_38,N_94);
nand U201 (N_201,N_152,In_129);
or U202 (N_202,In_156,In_395);
nor U203 (N_203,N_129,N_13);
nand U204 (N_204,In_353,N_9);
nand U205 (N_205,N_122,N_133);
and U206 (N_206,In_447,N_34);
nor U207 (N_207,In_147,In_41);
and U208 (N_208,In_310,N_164);
or U209 (N_209,In_373,In_490);
or U210 (N_210,N_4,In_250);
and U211 (N_211,In_81,N_44);
and U212 (N_212,N_14,N_130);
or U213 (N_213,N_64,In_317);
and U214 (N_214,N_125,N_167);
nor U215 (N_215,In_349,In_57);
and U216 (N_216,In_359,In_366);
nand U217 (N_217,In_172,In_323);
nor U218 (N_218,N_98,In_379);
or U219 (N_219,In_50,In_130);
or U220 (N_220,N_60,N_139);
or U221 (N_221,In_318,N_102);
nor U222 (N_222,In_341,N_59);
and U223 (N_223,N_113,N_38);
and U224 (N_224,In_253,N_15);
nor U225 (N_225,N_24,In_26);
and U226 (N_226,N_40,N_84);
and U227 (N_227,N_157,N_178);
nand U228 (N_228,N_140,In_290);
and U229 (N_229,N_128,In_289);
nor U230 (N_230,N_170,N_127);
nand U231 (N_231,N_42,N_110);
nor U232 (N_232,In_227,In_420);
nand U233 (N_233,N_138,N_5);
or U234 (N_234,In_187,In_238);
nand U235 (N_235,In_48,N_149);
nand U236 (N_236,In_176,In_316);
xnor U237 (N_237,In_254,In_499);
nor U238 (N_238,In_438,N_161);
nor U239 (N_239,In_103,In_236);
and U240 (N_240,In_459,In_60);
nand U241 (N_241,In_333,N_218);
nand U242 (N_242,In_5,In_80);
nand U243 (N_243,In_100,N_51);
or U244 (N_244,N_207,In_445);
and U245 (N_245,In_98,N_137);
and U246 (N_246,In_88,In_446);
nand U247 (N_247,In_72,In_7);
nand U248 (N_248,N_215,In_326);
or U249 (N_249,N_85,N_223);
nor U250 (N_250,N_204,In_443);
nor U251 (N_251,N_190,N_226);
nor U252 (N_252,N_88,In_51);
nor U253 (N_253,In_275,N_95);
nand U254 (N_254,N_100,N_3);
or U255 (N_255,N_196,In_153);
or U256 (N_256,N_134,N_169);
and U257 (N_257,N_103,N_112);
and U258 (N_258,In_142,N_172);
or U259 (N_259,N_71,N_235);
nand U260 (N_260,In_47,N_87);
or U261 (N_261,N_118,In_16);
nand U262 (N_262,In_93,In_35);
nor U263 (N_263,N_147,N_74);
or U264 (N_264,N_211,In_40);
or U265 (N_265,In_354,N_151);
nand U266 (N_266,In_33,N_124);
or U267 (N_267,In_269,N_69);
and U268 (N_268,N_145,N_175);
nand U269 (N_269,N_132,N_163);
nand U270 (N_270,In_376,N_160);
nor U271 (N_271,In_199,N_148);
nand U272 (N_272,N_234,In_242);
nand U273 (N_273,In_64,In_315);
and U274 (N_274,In_355,N_187);
and U275 (N_275,In_348,N_185);
and U276 (N_276,In_90,In_494);
or U277 (N_277,N_146,N_220);
and U278 (N_278,In_291,In_19);
nand U279 (N_279,In_203,N_73);
and U280 (N_280,N_72,In_320);
and U281 (N_281,In_248,In_185);
xnor U282 (N_282,In_74,N_231);
or U283 (N_283,In_190,In_465);
or U284 (N_284,N_45,N_126);
or U285 (N_285,N_205,N_221);
nor U286 (N_286,N_80,N_47);
nor U287 (N_287,N_158,In_337);
or U288 (N_288,N_180,N_238);
nor U289 (N_289,N_111,N_119);
nor U290 (N_290,In_308,N_155);
nor U291 (N_291,N_224,N_52);
or U292 (N_292,In_97,In_84);
nand U293 (N_293,N_11,N_188);
nand U294 (N_294,In_396,N_217);
nor U295 (N_295,In_125,In_119);
and U296 (N_296,In_417,N_213);
and U297 (N_297,In_286,N_179);
or U298 (N_298,N_198,N_20);
and U299 (N_299,In_391,In_37);
nor U300 (N_300,N_255,In_219);
nand U301 (N_301,N_232,N_197);
and U302 (N_302,N_120,N_272);
and U303 (N_303,N_216,In_331);
and U304 (N_304,N_251,In_232);
nand U305 (N_305,N_287,In_230);
and U306 (N_306,N_284,In_361);
nor U307 (N_307,N_236,N_194);
or U308 (N_308,In_92,In_229);
nand U309 (N_309,N_293,N_250);
nor U310 (N_310,In_279,N_123);
nand U311 (N_311,N_206,In_136);
nor U312 (N_312,In_28,N_184);
or U313 (N_313,N_253,N_201);
nor U314 (N_314,N_281,In_287);
or U315 (N_315,N_263,In_10);
nor U316 (N_316,N_276,In_321);
and U317 (N_317,N_181,N_259);
nor U318 (N_318,In_357,N_219);
or U319 (N_319,N_182,In_305);
nand U320 (N_320,N_258,N_299);
nor U321 (N_321,In_243,N_135);
nand U322 (N_322,N_252,N_285);
or U323 (N_323,In_94,N_109);
nor U324 (N_324,N_239,N_291);
nor U325 (N_325,N_249,N_278);
xor U326 (N_326,In_412,In_347);
or U327 (N_327,N_229,N_279);
nand U328 (N_328,N_77,N_296);
xnor U329 (N_329,N_22,N_92);
or U330 (N_330,In_11,In_195);
nand U331 (N_331,In_86,N_192);
nor U332 (N_332,N_230,In_456);
and U333 (N_333,N_261,N_193);
xor U334 (N_334,In_246,N_28);
nand U335 (N_335,In_300,N_282);
nand U336 (N_336,N_43,In_209);
and U337 (N_337,N_268,N_86);
and U338 (N_338,In_21,In_213);
or U339 (N_339,In_288,N_30);
or U340 (N_340,N_245,N_96);
nand U341 (N_341,In_62,N_273);
or U342 (N_342,N_150,N_243);
nor U343 (N_343,In_464,N_195);
or U344 (N_344,N_203,N_247);
nor U345 (N_345,N_227,N_121);
nand U346 (N_346,In_309,N_186);
nand U347 (N_347,N_294,N_136);
nor U348 (N_348,N_131,N_244);
or U349 (N_349,N_222,N_228);
nand U350 (N_350,N_280,N_54);
or U351 (N_351,N_48,In_338);
nand U352 (N_352,N_225,N_191);
nor U353 (N_353,N_283,In_360);
or U354 (N_354,N_189,N_265);
and U355 (N_355,In_145,N_199);
nor U356 (N_356,In_372,N_270);
and U357 (N_357,In_482,In_44);
nand U358 (N_358,N_269,In_31);
nor U359 (N_359,N_248,In_285);
nand U360 (N_360,N_82,N_357);
nor U361 (N_361,N_320,N_337);
nand U362 (N_362,N_312,N_156);
nor U363 (N_363,In_450,In_483);
or U364 (N_364,In_477,N_288);
or U365 (N_365,In_54,In_211);
nand U366 (N_366,N_307,N_305);
and U367 (N_367,N_341,In_364);
and U368 (N_368,N_262,N_241);
nor U369 (N_369,N_354,N_302);
nand U370 (N_370,N_313,N_356);
nor U371 (N_371,N_343,N_154);
and U372 (N_372,N_319,N_344);
or U373 (N_373,N_174,N_233);
and U374 (N_374,In_249,N_335);
nand U375 (N_375,N_349,In_20);
nor U376 (N_376,N_297,N_358);
or U377 (N_377,N_331,N_353);
or U378 (N_378,N_200,N_208);
and U379 (N_379,N_183,N_355);
or U380 (N_380,N_214,In_281);
and U381 (N_381,N_289,N_260);
or U382 (N_382,N_105,N_292);
nor U383 (N_383,N_310,N_264);
nor U384 (N_384,N_330,N_317);
or U385 (N_385,N_340,N_33);
nor U386 (N_386,N_266,In_45);
nor U387 (N_387,N_338,N_237);
xnor U388 (N_388,N_304,N_275);
nor U389 (N_389,N_36,N_333);
nand U390 (N_390,N_89,N_209);
xnor U391 (N_391,In_61,In_164);
nand U392 (N_392,N_162,N_141);
nand U393 (N_393,N_315,N_346);
or U394 (N_394,N_274,N_348);
or U395 (N_395,N_303,N_311);
or U396 (N_396,N_306,In_390);
nand U397 (N_397,N_316,N_321);
or U398 (N_398,N_329,N_326);
nor U399 (N_399,N_301,N_298);
and U400 (N_400,N_359,N_336);
and U401 (N_401,N_173,N_256);
nand U402 (N_402,N_339,N_143);
nand U403 (N_403,In_495,N_347);
or U404 (N_404,N_342,N_318);
or U405 (N_405,N_328,N_277);
or U406 (N_406,In_491,N_142);
or U407 (N_407,In_466,In_247);
nor U408 (N_408,In_177,N_1);
nor U409 (N_409,In_149,N_334);
nor U410 (N_410,N_352,N_165);
nor U411 (N_411,In_165,N_309);
or U412 (N_412,N_257,In_266);
and U413 (N_413,N_210,N_327);
nand U414 (N_414,In_441,N_351);
or U415 (N_415,In_479,N_300);
and U416 (N_416,N_115,N_290);
nor U417 (N_417,N_78,N_314);
or U418 (N_418,N_322,N_325);
nor U419 (N_419,N_240,N_242);
nor U420 (N_420,N_407,N_286);
nor U421 (N_421,N_392,N_379);
or U422 (N_422,N_401,N_412);
and U423 (N_423,N_411,N_364);
nand U424 (N_424,N_202,N_380);
or U425 (N_425,N_365,N_400);
or U426 (N_426,N_406,N_308);
and U427 (N_427,N_332,N_410);
or U428 (N_428,N_418,N_383);
or U429 (N_429,N_419,N_171);
nand U430 (N_430,N_369,N_415);
nand U431 (N_431,N_384,N_386);
or U432 (N_432,N_414,N_413);
and U433 (N_433,N_375,N_361);
and U434 (N_434,N_391,N_403);
nor U435 (N_435,N_368,N_373);
nor U436 (N_436,N_363,N_389);
and U437 (N_437,N_377,N_395);
or U438 (N_438,N_362,N_398);
nand U439 (N_439,N_212,N_57);
nor U440 (N_440,In_416,In_91);
nand U441 (N_441,In_404,N_408);
and U442 (N_442,N_393,N_371);
and U443 (N_443,N_374,N_397);
xnor U444 (N_444,N_345,N_372);
and U445 (N_445,N_166,N_366);
nand U446 (N_446,N_396,N_246);
and U447 (N_447,N_409,N_405);
or U448 (N_448,N_385,N_381);
or U449 (N_449,N_388,N_417);
nor U450 (N_450,N_370,N_350);
nand U451 (N_451,N_416,N_390);
nand U452 (N_452,N_323,N_360);
nand U453 (N_453,N_267,N_324);
nor U454 (N_454,N_295,N_254);
and U455 (N_455,N_402,N_387);
nand U456 (N_456,N_404,N_367);
nor U457 (N_457,N_378,N_382);
nor U458 (N_458,N_271,N_394);
and U459 (N_459,N_399,N_376);
and U460 (N_460,N_417,N_246);
nor U461 (N_461,N_372,N_375);
nor U462 (N_462,N_267,N_323);
nor U463 (N_463,N_418,N_360);
or U464 (N_464,N_398,N_402);
nor U465 (N_465,In_91,N_366);
and U466 (N_466,N_377,N_398);
or U467 (N_467,N_166,In_416);
nand U468 (N_468,N_405,N_395);
nor U469 (N_469,N_376,N_373);
nor U470 (N_470,N_286,N_391);
nand U471 (N_471,In_91,N_403);
nand U472 (N_472,N_401,N_286);
nor U473 (N_473,N_391,N_377);
and U474 (N_474,N_419,N_393);
and U475 (N_475,N_365,N_382);
nor U476 (N_476,N_419,N_386);
or U477 (N_477,N_396,In_91);
nor U478 (N_478,N_295,N_373);
or U479 (N_479,N_397,N_371);
nor U480 (N_480,N_426,N_425);
and U481 (N_481,N_462,N_455);
and U482 (N_482,N_431,N_470);
and U483 (N_483,N_460,N_458);
or U484 (N_484,N_466,N_445);
and U485 (N_485,N_437,N_424);
and U486 (N_486,N_434,N_469);
nor U487 (N_487,N_422,N_457);
and U488 (N_488,N_471,N_441);
nand U489 (N_489,N_438,N_474);
and U490 (N_490,N_451,N_475);
nand U491 (N_491,N_468,N_444);
nand U492 (N_492,N_461,N_446);
nor U493 (N_493,N_440,N_436);
nor U494 (N_494,N_427,N_443);
nand U495 (N_495,N_478,N_435);
nor U496 (N_496,N_454,N_449);
or U497 (N_497,N_428,N_453);
nand U498 (N_498,N_433,N_477);
nor U499 (N_499,N_463,N_473);
and U500 (N_500,N_465,N_450);
nand U501 (N_501,N_423,N_447);
and U502 (N_502,N_448,N_472);
and U503 (N_503,N_420,N_456);
or U504 (N_504,N_430,N_432);
or U505 (N_505,N_464,N_421);
or U506 (N_506,N_467,N_439);
nor U507 (N_507,N_429,N_479);
nand U508 (N_508,N_452,N_476);
nand U509 (N_509,N_442,N_459);
nand U510 (N_510,N_442,N_463);
or U511 (N_511,N_463,N_468);
nand U512 (N_512,N_446,N_425);
or U513 (N_513,N_472,N_440);
xor U514 (N_514,N_421,N_474);
and U515 (N_515,N_471,N_449);
and U516 (N_516,N_428,N_462);
and U517 (N_517,N_433,N_421);
and U518 (N_518,N_446,N_441);
or U519 (N_519,N_463,N_458);
nand U520 (N_520,N_463,N_476);
and U521 (N_521,N_461,N_471);
nor U522 (N_522,N_475,N_450);
and U523 (N_523,N_443,N_458);
nor U524 (N_524,N_469,N_436);
and U525 (N_525,N_452,N_473);
nor U526 (N_526,N_475,N_458);
nor U527 (N_527,N_432,N_450);
nor U528 (N_528,N_449,N_433);
nor U529 (N_529,N_451,N_474);
nor U530 (N_530,N_457,N_478);
or U531 (N_531,N_468,N_455);
and U532 (N_532,N_463,N_464);
or U533 (N_533,N_433,N_462);
nor U534 (N_534,N_472,N_439);
xor U535 (N_535,N_460,N_438);
and U536 (N_536,N_439,N_437);
and U537 (N_537,N_452,N_464);
or U538 (N_538,N_467,N_434);
nor U539 (N_539,N_451,N_432);
nor U540 (N_540,N_525,N_519);
nand U541 (N_541,N_511,N_500);
nand U542 (N_542,N_505,N_524);
nand U543 (N_543,N_488,N_491);
nand U544 (N_544,N_508,N_535);
nor U545 (N_545,N_484,N_480);
nor U546 (N_546,N_526,N_536);
or U547 (N_547,N_502,N_496);
or U548 (N_548,N_504,N_522);
xnor U549 (N_549,N_494,N_506);
xor U550 (N_550,N_534,N_492);
nor U551 (N_551,N_538,N_531);
nand U552 (N_552,N_528,N_530);
xnor U553 (N_553,N_529,N_539);
or U554 (N_554,N_490,N_498);
and U555 (N_555,N_513,N_523);
nor U556 (N_556,N_489,N_509);
nand U557 (N_557,N_532,N_518);
nand U558 (N_558,N_486,N_521);
nand U559 (N_559,N_503,N_487);
nand U560 (N_560,N_481,N_482);
and U561 (N_561,N_537,N_495);
nand U562 (N_562,N_520,N_483);
nand U563 (N_563,N_527,N_517);
nand U564 (N_564,N_499,N_533);
or U565 (N_565,N_493,N_485);
or U566 (N_566,N_515,N_512);
nand U567 (N_567,N_514,N_516);
or U568 (N_568,N_510,N_501);
or U569 (N_569,N_507,N_497);
nor U570 (N_570,N_480,N_525);
or U571 (N_571,N_503,N_483);
or U572 (N_572,N_493,N_525);
xnor U573 (N_573,N_495,N_503);
nor U574 (N_574,N_484,N_504);
nor U575 (N_575,N_522,N_514);
and U576 (N_576,N_515,N_513);
nand U577 (N_577,N_509,N_504);
nor U578 (N_578,N_490,N_491);
or U579 (N_579,N_491,N_537);
nand U580 (N_580,N_538,N_503);
nand U581 (N_581,N_518,N_512);
nand U582 (N_582,N_534,N_525);
nand U583 (N_583,N_515,N_521);
xor U584 (N_584,N_490,N_516);
xor U585 (N_585,N_536,N_482);
xor U586 (N_586,N_513,N_535);
and U587 (N_587,N_480,N_539);
or U588 (N_588,N_525,N_522);
nor U589 (N_589,N_533,N_501);
and U590 (N_590,N_526,N_501);
and U591 (N_591,N_526,N_480);
nor U592 (N_592,N_537,N_514);
nand U593 (N_593,N_487,N_504);
nand U594 (N_594,N_535,N_491);
or U595 (N_595,N_509,N_495);
nand U596 (N_596,N_488,N_510);
or U597 (N_597,N_486,N_489);
or U598 (N_598,N_485,N_538);
or U599 (N_599,N_487,N_526);
and U600 (N_600,N_580,N_574);
and U601 (N_601,N_572,N_560);
xnor U602 (N_602,N_595,N_597);
or U603 (N_603,N_584,N_551);
nor U604 (N_604,N_570,N_555);
nand U605 (N_605,N_582,N_553);
nor U606 (N_606,N_554,N_548);
or U607 (N_607,N_545,N_549);
nor U608 (N_608,N_540,N_593);
and U609 (N_609,N_599,N_565);
and U610 (N_610,N_587,N_547);
nand U611 (N_611,N_541,N_571);
and U612 (N_612,N_563,N_569);
nand U613 (N_613,N_546,N_567);
nand U614 (N_614,N_552,N_591);
or U615 (N_615,N_577,N_562);
or U616 (N_616,N_581,N_543);
or U617 (N_617,N_575,N_564);
nor U618 (N_618,N_592,N_550);
nor U619 (N_619,N_594,N_561);
nor U620 (N_620,N_559,N_568);
and U621 (N_621,N_578,N_583);
nand U622 (N_622,N_585,N_596);
or U623 (N_623,N_557,N_556);
and U624 (N_624,N_598,N_544);
nor U625 (N_625,N_558,N_586);
nand U626 (N_626,N_566,N_576);
nand U627 (N_627,N_589,N_579);
nand U628 (N_628,N_588,N_573);
and U629 (N_629,N_542,N_590);
nand U630 (N_630,N_573,N_567);
or U631 (N_631,N_599,N_552);
and U632 (N_632,N_597,N_580);
and U633 (N_633,N_575,N_572);
xnor U634 (N_634,N_596,N_556);
and U635 (N_635,N_554,N_547);
or U636 (N_636,N_551,N_545);
nand U637 (N_637,N_577,N_549);
and U638 (N_638,N_540,N_589);
and U639 (N_639,N_582,N_583);
nor U640 (N_640,N_567,N_540);
or U641 (N_641,N_547,N_540);
and U642 (N_642,N_558,N_552);
and U643 (N_643,N_586,N_553);
nor U644 (N_644,N_598,N_540);
nand U645 (N_645,N_544,N_579);
and U646 (N_646,N_574,N_585);
and U647 (N_647,N_549,N_568);
nand U648 (N_648,N_552,N_544);
nand U649 (N_649,N_589,N_573);
and U650 (N_650,N_592,N_597);
nand U651 (N_651,N_576,N_573);
nand U652 (N_652,N_592,N_548);
nor U653 (N_653,N_588,N_560);
and U654 (N_654,N_568,N_585);
nand U655 (N_655,N_558,N_589);
and U656 (N_656,N_597,N_555);
nor U657 (N_657,N_596,N_558);
and U658 (N_658,N_583,N_565);
nand U659 (N_659,N_551,N_598);
or U660 (N_660,N_617,N_625);
and U661 (N_661,N_654,N_628);
xnor U662 (N_662,N_645,N_600);
and U663 (N_663,N_613,N_649);
nor U664 (N_664,N_641,N_653);
xnor U665 (N_665,N_633,N_607);
nor U666 (N_666,N_626,N_627);
or U667 (N_667,N_623,N_647);
nor U668 (N_668,N_602,N_624);
nor U669 (N_669,N_650,N_639);
or U670 (N_670,N_618,N_642);
nor U671 (N_671,N_611,N_612);
nand U672 (N_672,N_605,N_620);
or U673 (N_673,N_610,N_604);
nand U674 (N_674,N_631,N_606);
nor U675 (N_675,N_616,N_643);
nor U676 (N_676,N_632,N_655);
or U677 (N_677,N_651,N_614);
nand U678 (N_678,N_634,N_656);
or U679 (N_679,N_609,N_603);
or U680 (N_680,N_658,N_622);
and U681 (N_681,N_637,N_636);
and U682 (N_682,N_615,N_659);
and U683 (N_683,N_630,N_601);
nand U684 (N_684,N_608,N_621);
nor U685 (N_685,N_648,N_629);
nor U686 (N_686,N_652,N_646);
xor U687 (N_687,N_640,N_644);
nor U688 (N_688,N_635,N_657);
nor U689 (N_689,N_638,N_619);
nor U690 (N_690,N_617,N_632);
and U691 (N_691,N_611,N_647);
nor U692 (N_692,N_600,N_609);
nor U693 (N_693,N_609,N_608);
and U694 (N_694,N_618,N_650);
nand U695 (N_695,N_641,N_644);
nor U696 (N_696,N_633,N_627);
and U697 (N_697,N_617,N_603);
nor U698 (N_698,N_612,N_614);
nand U699 (N_699,N_644,N_608);
or U700 (N_700,N_625,N_650);
nand U701 (N_701,N_621,N_654);
or U702 (N_702,N_647,N_644);
nor U703 (N_703,N_652,N_614);
nand U704 (N_704,N_630,N_638);
and U705 (N_705,N_639,N_653);
nor U706 (N_706,N_647,N_632);
and U707 (N_707,N_630,N_604);
nor U708 (N_708,N_627,N_615);
and U709 (N_709,N_659,N_628);
or U710 (N_710,N_636,N_653);
nand U711 (N_711,N_636,N_625);
or U712 (N_712,N_650,N_615);
nor U713 (N_713,N_615,N_636);
nand U714 (N_714,N_606,N_607);
or U715 (N_715,N_625,N_607);
nor U716 (N_716,N_639,N_624);
and U717 (N_717,N_609,N_644);
nand U718 (N_718,N_658,N_603);
or U719 (N_719,N_630,N_634);
nand U720 (N_720,N_675,N_695);
and U721 (N_721,N_718,N_668);
nor U722 (N_722,N_713,N_664);
and U723 (N_723,N_678,N_711);
and U724 (N_724,N_673,N_712);
and U725 (N_725,N_686,N_696);
or U726 (N_726,N_683,N_688);
and U727 (N_727,N_717,N_715);
nor U728 (N_728,N_684,N_719);
and U729 (N_729,N_680,N_693);
xnor U730 (N_730,N_679,N_662);
or U731 (N_731,N_671,N_705);
nand U732 (N_732,N_676,N_709);
nor U733 (N_733,N_697,N_665);
nor U734 (N_734,N_708,N_681);
and U735 (N_735,N_682,N_716);
nand U736 (N_736,N_669,N_694);
nand U737 (N_737,N_710,N_660);
nand U738 (N_738,N_714,N_672);
and U739 (N_739,N_670,N_677);
and U740 (N_740,N_690,N_703);
nor U741 (N_741,N_700,N_687);
nand U742 (N_742,N_702,N_689);
nand U743 (N_743,N_699,N_667);
and U744 (N_744,N_674,N_701);
nor U745 (N_745,N_661,N_691);
nand U746 (N_746,N_666,N_704);
nand U747 (N_747,N_663,N_706);
or U748 (N_748,N_698,N_692);
and U749 (N_749,N_685,N_707);
nor U750 (N_750,N_710,N_700);
or U751 (N_751,N_673,N_670);
or U752 (N_752,N_709,N_675);
nand U753 (N_753,N_667,N_686);
nand U754 (N_754,N_669,N_680);
or U755 (N_755,N_699,N_690);
or U756 (N_756,N_668,N_716);
nor U757 (N_757,N_706,N_661);
and U758 (N_758,N_719,N_700);
or U759 (N_759,N_688,N_712);
and U760 (N_760,N_698,N_678);
nor U761 (N_761,N_691,N_707);
and U762 (N_762,N_707,N_660);
and U763 (N_763,N_696,N_666);
nor U764 (N_764,N_715,N_662);
or U765 (N_765,N_698,N_703);
nor U766 (N_766,N_703,N_718);
nand U767 (N_767,N_665,N_675);
nor U768 (N_768,N_670,N_691);
nand U769 (N_769,N_664,N_661);
nor U770 (N_770,N_677,N_719);
or U771 (N_771,N_667,N_715);
nor U772 (N_772,N_677,N_697);
nand U773 (N_773,N_702,N_719);
and U774 (N_774,N_685,N_673);
nand U775 (N_775,N_664,N_702);
xnor U776 (N_776,N_692,N_681);
and U777 (N_777,N_719,N_665);
nand U778 (N_778,N_666,N_684);
or U779 (N_779,N_665,N_684);
nor U780 (N_780,N_731,N_765);
nand U781 (N_781,N_760,N_776);
and U782 (N_782,N_728,N_777);
nand U783 (N_783,N_759,N_774);
nand U784 (N_784,N_779,N_732);
nand U785 (N_785,N_737,N_751);
nand U786 (N_786,N_738,N_739);
or U787 (N_787,N_745,N_758);
nand U788 (N_788,N_742,N_740);
nor U789 (N_789,N_756,N_762);
nand U790 (N_790,N_761,N_734);
and U791 (N_791,N_721,N_766);
and U792 (N_792,N_748,N_764);
nor U793 (N_793,N_729,N_749);
or U794 (N_794,N_726,N_770);
nand U795 (N_795,N_752,N_755);
or U796 (N_796,N_730,N_750);
nor U797 (N_797,N_736,N_746);
and U798 (N_798,N_773,N_735);
nor U799 (N_799,N_733,N_768);
or U800 (N_800,N_725,N_744);
nor U801 (N_801,N_778,N_747);
and U802 (N_802,N_727,N_763);
and U803 (N_803,N_724,N_753);
xnor U804 (N_804,N_769,N_722);
and U805 (N_805,N_771,N_741);
and U806 (N_806,N_767,N_743);
and U807 (N_807,N_775,N_754);
or U808 (N_808,N_720,N_723);
nand U809 (N_809,N_772,N_757);
or U810 (N_810,N_776,N_743);
and U811 (N_811,N_735,N_779);
nor U812 (N_812,N_770,N_757);
nand U813 (N_813,N_746,N_748);
nor U814 (N_814,N_738,N_776);
and U815 (N_815,N_757,N_759);
or U816 (N_816,N_723,N_744);
or U817 (N_817,N_758,N_747);
nor U818 (N_818,N_746,N_727);
nor U819 (N_819,N_779,N_766);
or U820 (N_820,N_778,N_738);
nor U821 (N_821,N_729,N_736);
or U822 (N_822,N_754,N_725);
or U823 (N_823,N_769,N_756);
and U824 (N_824,N_773,N_749);
nand U825 (N_825,N_751,N_728);
or U826 (N_826,N_765,N_724);
or U827 (N_827,N_762,N_777);
or U828 (N_828,N_750,N_729);
nor U829 (N_829,N_745,N_723);
nor U830 (N_830,N_776,N_725);
nand U831 (N_831,N_764,N_758);
nor U832 (N_832,N_731,N_771);
nand U833 (N_833,N_758,N_735);
or U834 (N_834,N_768,N_775);
or U835 (N_835,N_773,N_772);
nor U836 (N_836,N_751,N_736);
nor U837 (N_837,N_745,N_760);
xor U838 (N_838,N_777,N_756);
or U839 (N_839,N_765,N_737);
nor U840 (N_840,N_802,N_799);
nand U841 (N_841,N_836,N_783);
or U842 (N_842,N_793,N_784);
or U843 (N_843,N_822,N_820);
nand U844 (N_844,N_812,N_801);
nor U845 (N_845,N_804,N_794);
nand U846 (N_846,N_814,N_810);
or U847 (N_847,N_823,N_803);
and U848 (N_848,N_797,N_829);
nand U849 (N_849,N_826,N_781);
xnor U850 (N_850,N_834,N_837);
or U851 (N_851,N_786,N_787);
and U852 (N_852,N_805,N_791);
and U853 (N_853,N_798,N_830);
nor U854 (N_854,N_825,N_785);
or U855 (N_855,N_813,N_780);
nor U856 (N_856,N_832,N_806);
nor U857 (N_857,N_807,N_835);
or U858 (N_858,N_816,N_796);
or U859 (N_859,N_800,N_790);
or U860 (N_860,N_827,N_833);
or U861 (N_861,N_811,N_789);
or U862 (N_862,N_831,N_792);
nor U863 (N_863,N_819,N_795);
nand U864 (N_864,N_788,N_808);
nand U865 (N_865,N_824,N_838);
or U866 (N_866,N_839,N_818);
nor U867 (N_867,N_809,N_828);
xor U868 (N_868,N_782,N_821);
or U869 (N_869,N_815,N_817);
nand U870 (N_870,N_825,N_793);
or U871 (N_871,N_786,N_785);
and U872 (N_872,N_816,N_834);
nor U873 (N_873,N_803,N_836);
or U874 (N_874,N_823,N_791);
or U875 (N_875,N_780,N_835);
or U876 (N_876,N_786,N_783);
nor U877 (N_877,N_782,N_806);
nor U878 (N_878,N_808,N_796);
and U879 (N_879,N_822,N_796);
or U880 (N_880,N_827,N_837);
nor U881 (N_881,N_817,N_796);
nand U882 (N_882,N_782,N_780);
nor U883 (N_883,N_826,N_780);
xor U884 (N_884,N_839,N_800);
or U885 (N_885,N_838,N_819);
and U886 (N_886,N_797,N_798);
nand U887 (N_887,N_803,N_792);
and U888 (N_888,N_826,N_806);
and U889 (N_889,N_799,N_821);
nor U890 (N_890,N_836,N_827);
nand U891 (N_891,N_826,N_785);
or U892 (N_892,N_795,N_815);
nor U893 (N_893,N_792,N_836);
nor U894 (N_894,N_835,N_790);
nand U895 (N_895,N_807,N_803);
nand U896 (N_896,N_837,N_793);
nand U897 (N_897,N_784,N_791);
or U898 (N_898,N_832,N_798);
and U899 (N_899,N_838,N_802);
or U900 (N_900,N_850,N_860);
nand U901 (N_901,N_878,N_888);
nand U902 (N_902,N_891,N_847);
nor U903 (N_903,N_898,N_842);
and U904 (N_904,N_897,N_876);
and U905 (N_905,N_874,N_872);
nor U906 (N_906,N_892,N_883);
nor U907 (N_907,N_873,N_882);
or U908 (N_908,N_875,N_852);
or U909 (N_909,N_853,N_856);
or U910 (N_910,N_866,N_893);
nand U911 (N_911,N_849,N_863);
nor U912 (N_912,N_858,N_884);
nand U913 (N_913,N_896,N_846);
and U914 (N_914,N_861,N_854);
nor U915 (N_915,N_843,N_885);
nand U916 (N_916,N_845,N_886);
and U917 (N_917,N_864,N_857);
or U918 (N_918,N_865,N_879);
and U919 (N_919,N_894,N_889);
and U920 (N_920,N_890,N_862);
nand U921 (N_921,N_869,N_871);
and U922 (N_922,N_870,N_867);
and U923 (N_923,N_841,N_844);
nand U924 (N_924,N_851,N_880);
nor U925 (N_925,N_887,N_899);
nor U926 (N_926,N_848,N_859);
nand U927 (N_927,N_877,N_895);
xor U928 (N_928,N_881,N_855);
and U929 (N_929,N_840,N_868);
or U930 (N_930,N_883,N_890);
and U931 (N_931,N_876,N_862);
nor U932 (N_932,N_883,N_881);
nand U933 (N_933,N_898,N_887);
nand U934 (N_934,N_857,N_843);
or U935 (N_935,N_898,N_873);
or U936 (N_936,N_853,N_878);
nand U937 (N_937,N_888,N_890);
and U938 (N_938,N_840,N_853);
nand U939 (N_939,N_896,N_871);
nor U940 (N_940,N_867,N_842);
nand U941 (N_941,N_887,N_860);
or U942 (N_942,N_874,N_868);
nor U943 (N_943,N_874,N_889);
or U944 (N_944,N_858,N_855);
or U945 (N_945,N_861,N_864);
nand U946 (N_946,N_847,N_855);
nand U947 (N_947,N_890,N_894);
and U948 (N_948,N_892,N_879);
nand U949 (N_949,N_891,N_853);
nor U950 (N_950,N_854,N_870);
or U951 (N_951,N_845,N_876);
or U952 (N_952,N_852,N_872);
and U953 (N_953,N_847,N_857);
and U954 (N_954,N_850,N_877);
or U955 (N_955,N_886,N_869);
nand U956 (N_956,N_846,N_855);
nand U957 (N_957,N_879,N_876);
nor U958 (N_958,N_887,N_897);
and U959 (N_959,N_847,N_895);
or U960 (N_960,N_944,N_905);
or U961 (N_961,N_913,N_920);
nand U962 (N_962,N_947,N_927);
nand U963 (N_963,N_949,N_934);
and U964 (N_964,N_953,N_921);
nor U965 (N_965,N_929,N_945);
nand U966 (N_966,N_906,N_924);
and U967 (N_967,N_938,N_935);
nand U968 (N_968,N_908,N_917);
nor U969 (N_969,N_951,N_903);
nor U970 (N_970,N_954,N_943);
and U971 (N_971,N_932,N_955);
nor U972 (N_972,N_912,N_958);
nand U973 (N_973,N_939,N_941);
or U974 (N_974,N_936,N_957);
or U975 (N_975,N_914,N_942);
nand U976 (N_976,N_952,N_901);
and U977 (N_977,N_911,N_948);
nor U978 (N_978,N_946,N_915);
nand U979 (N_979,N_950,N_959);
nor U980 (N_980,N_922,N_918);
or U981 (N_981,N_940,N_931);
or U982 (N_982,N_923,N_956);
and U983 (N_983,N_904,N_926);
and U984 (N_984,N_925,N_928);
nor U985 (N_985,N_907,N_937);
nand U986 (N_986,N_910,N_916);
and U987 (N_987,N_930,N_919);
nand U988 (N_988,N_902,N_909);
or U989 (N_989,N_900,N_933);
or U990 (N_990,N_929,N_954);
or U991 (N_991,N_946,N_907);
nand U992 (N_992,N_925,N_954);
or U993 (N_993,N_952,N_916);
nor U994 (N_994,N_905,N_955);
and U995 (N_995,N_906,N_915);
nand U996 (N_996,N_910,N_954);
and U997 (N_997,N_953,N_951);
and U998 (N_998,N_944,N_938);
or U999 (N_999,N_947,N_913);
or U1000 (N_1000,N_953,N_944);
nor U1001 (N_1001,N_930,N_953);
and U1002 (N_1002,N_934,N_956);
xor U1003 (N_1003,N_934,N_953);
and U1004 (N_1004,N_959,N_955);
nor U1005 (N_1005,N_902,N_908);
nand U1006 (N_1006,N_944,N_955);
nand U1007 (N_1007,N_908,N_901);
nand U1008 (N_1008,N_909,N_903);
nor U1009 (N_1009,N_900,N_909);
and U1010 (N_1010,N_957,N_951);
or U1011 (N_1011,N_942,N_930);
nand U1012 (N_1012,N_935,N_921);
and U1013 (N_1013,N_944,N_919);
and U1014 (N_1014,N_925,N_936);
and U1015 (N_1015,N_946,N_926);
nand U1016 (N_1016,N_959,N_937);
nand U1017 (N_1017,N_950,N_933);
nor U1018 (N_1018,N_923,N_945);
or U1019 (N_1019,N_949,N_902);
nand U1020 (N_1020,N_961,N_960);
and U1021 (N_1021,N_1002,N_997);
nor U1022 (N_1022,N_1004,N_1000);
nor U1023 (N_1023,N_973,N_1001);
and U1024 (N_1024,N_968,N_1012);
and U1025 (N_1025,N_980,N_1019);
or U1026 (N_1026,N_967,N_989);
nand U1027 (N_1027,N_981,N_1014);
nor U1028 (N_1028,N_976,N_998);
or U1029 (N_1029,N_1017,N_964);
and U1030 (N_1030,N_982,N_984);
nand U1031 (N_1031,N_983,N_1009);
nor U1032 (N_1032,N_993,N_977);
nor U1033 (N_1033,N_1015,N_1007);
and U1034 (N_1034,N_995,N_966);
nor U1035 (N_1035,N_999,N_969);
nand U1036 (N_1036,N_986,N_971);
and U1037 (N_1037,N_988,N_990);
and U1038 (N_1038,N_1018,N_970);
and U1039 (N_1039,N_975,N_1006);
nor U1040 (N_1040,N_996,N_1016);
nor U1041 (N_1041,N_1005,N_979);
nor U1042 (N_1042,N_974,N_1010);
or U1043 (N_1043,N_994,N_1008);
nand U1044 (N_1044,N_962,N_972);
and U1045 (N_1045,N_987,N_978);
or U1046 (N_1046,N_985,N_992);
nand U1047 (N_1047,N_963,N_991);
nand U1048 (N_1048,N_965,N_1003);
and U1049 (N_1049,N_1013,N_1011);
nand U1050 (N_1050,N_1000,N_966);
nor U1051 (N_1051,N_1014,N_962);
or U1052 (N_1052,N_1014,N_1015);
or U1053 (N_1053,N_1012,N_967);
and U1054 (N_1054,N_1018,N_1017);
or U1055 (N_1055,N_1000,N_981);
xor U1056 (N_1056,N_985,N_1004);
nand U1057 (N_1057,N_976,N_977);
and U1058 (N_1058,N_1015,N_965);
and U1059 (N_1059,N_983,N_991);
nor U1060 (N_1060,N_962,N_1016);
and U1061 (N_1061,N_1010,N_965);
and U1062 (N_1062,N_963,N_974);
or U1063 (N_1063,N_991,N_994);
nor U1064 (N_1064,N_973,N_962);
and U1065 (N_1065,N_1015,N_994);
xor U1066 (N_1066,N_1014,N_1016);
and U1067 (N_1067,N_1002,N_1015);
and U1068 (N_1068,N_992,N_1013);
and U1069 (N_1069,N_989,N_962);
nor U1070 (N_1070,N_990,N_974);
nand U1071 (N_1071,N_1011,N_987);
nor U1072 (N_1072,N_991,N_1018);
nand U1073 (N_1073,N_1009,N_974);
and U1074 (N_1074,N_987,N_983);
nand U1075 (N_1075,N_968,N_997);
nor U1076 (N_1076,N_1007,N_969);
nor U1077 (N_1077,N_1001,N_1016);
nand U1078 (N_1078,N_992,N_987);
and U1079 (N_1079,N_1014,N_969);
nor U1080 (N_1080,N_1048,N_1046);
or U1081 (N_1081,N_1037,N_1068);
and U1082 (N_1082,N_1066,N_1033);
or U1083 (N_1083,N_1027,N_1022);
nand U1084 (N_1084,N_1059,N_1035);
nor U1085 (N_1085,N_1040,N_1050);
nand U1086 (N_1086,N_1062,N_1071);
nor U1087 (N_1087,N_1065,N_1063);
nand U1088 (N_1088,N_1038,N_1024);
and U1089 (N_1089,N_1070,N_1052);
or U1090 (N_1090,N_1075,N_1061);
xnor U1091 (N_1091,N_1045,N_1028);
nor U1092 (N_1092,N_1030,N_1051);
nor U1093 (N_1093,N_1056,N_1029);
nor U1094 (N_1094,N_1072,N_1042);
or U1095 (N_1095,N_1054,N_1025);
or U1096 (N_1096,N_1023,N_1064);
nor U1097 (N_1097,N_1020,N_1057);
and U1098 (N_1098,N_1060,N_1036);
and U1099 (N_1099,N_1047,N_1044);
nor U1100 (N_1100,N_1049,N_1078);
nor U1101 (N_1101,N_1073,N_1076);
nor U1102 (N_1102,N_1041,N_1053);
nor U1103 (N_1103,N_1077,N_1039);
or U1104 (N_1104,N_1034,N_1031);
or U1105 (N_1105,N_1055,N_1067);
nor U1106 (N_1106,N_1069,N_1043);
and U1107 (N_1107,N_1058,N_1021);
nand U1108 (N_1108,N_1032,N_1074);
or U1109 (N_1109,N_1079,N_1026);
nand U1110 (N_1110,N_1051,N_1074);
or U1111 (N_1111,N_1033,N_1024);
or U1112 (N_1112,N_1043,N_1063);
or U1113 (N_1113,N_1061,N_1056);
nor U1114 (N_1114,N_1061,N_1038);
nor U1115 (N_1115,N_1059,N_1055);
nor U1116 (N_1116,N_1037,N_1051);
nor U1117 (N_1117,N_1072,N_1076);
or U1118 (N_1118,N_1029,N_1028);
nand U1119 (N_1119,N_1057,N_1079);
xnor U1120 (N_1120,N_1032,N_1025);
nor U1121 (N_1121,N_1071,N_1065);
or U1122 (N_1122,N_1056,N_1032);
and U1123 (N_1123,N_1044,N_1031);
or U1124 (N_1124,N_1032,N_1038);
nand U1125 (N_1125,N_1055,N_1050);
nor U1126 (N_1126,N_1030,N_1046);
or U1127 (N_1127,N_1030,N_1058);
nand U1128 (N_1128,N_1077,N_1042);
nor U1129 (N_1129,N_1078,N_1058);
nor U1130 (N_1130,N_1023,N_1043);
or U1131 (N_1131,N_1025,N_1035);
nand U1132 (N_1132,N_1059,N_1043);
and U1133 (N_1133,N_1028,N_1038);
xnor U1134 (N_1134,N_1078,N_1035);
and U1135 (N_1135,N_1076,N_1036);
nand U1136 (N_1136,N_1064,N_1069);
and U1137 (N_1137,N_1043,N_1062);
or U1138 (N_1138,N_1032,N_1049);
nand U1139 (N_1139,N_1051,N_1064);
nand U1140 (N_1140,N_1098,N_1123);
nand U1141 (N_1141,N_1132,N_1110);
and U1142 (N_1142,N_1101,N_1102);
nor U1143 (N_1143,N_1100,N_1087);
or U1144 (N_1144,N_1127,N_1105);
or U1145 (N_1145,N_1113,N_1107);
nor U1146 (N_1146,N_1097,N_1085);
nand U1147 (N_1147,N_1086,N_1115);
and U1148 (N_1148,N_1121,N_1134);
and U1149 (N_1149,N_1139,N_1091);
or U1150 (N_1150,N_1120,N_1095);
and U1151 (N_1151,N_1090,N_1135);
or U1152 (N_1152,N_1088,N_1083);
or U1153 (N_1153,N_1124,N_1108);
and U1154 (N_1154,N_1131,N_1126);
or U1155 (N_1155,N_1080,N_1116);
nor U1156 (N_1156,N_1081,N_1112);
nand U1157 (N_1157,N_1099,N_1092);
nand U1158 (N_1158,N_1122,N_1118);
nand U1159 (N_1159,N_1093,N_1103);
or U1160 (N_1160,N_1109,N_1136);
nor U1161 (N_1161,N_1117,N_1104);
or U1162 (N_1162,N_1082,N_1129);
nand U1163 (N_1163,N_1094,N_1096);
nand U1164 (N_1164,N_1084,N_1133);
nand U1165 (N_1165,N_1111,N_1138);
nand U1166 (N_1166,N_1137,N_1128);
and U1167 (N_1167,N_1106,N_1089);
xor U1168 (N_1168,N_1119,N_1114);
nand U1169 (N_1169,N_1130,N_1125);
nand U1170 (N_1170,N_1105,N_1111);
nor U1171 (N_1171,N_1139,N_1081);
or U1172 (N_1172,N_1098,N_1082);
or U1173 (N_1173,N_1138,N_1119);
nor U1174 (N_1174,N_1139,N_1106);
or U1175 (N_1175,N_1110,N_1108);
or U1176 (N_1176,N_1095,N_1136);
or U1177 (N_1177,N_1113,N_1118);
and U1178 (N_1178,N_1102,N_1099);
nand U1179 (N_1179,N_1091,N_1138);
and U1180 (N_1180,N_1109,N_1119);
nor U1181 (N_1181,N_1080,N_1123);
or U1182 (N_1182,N_1093,N_1135);
nor U1183 (N_1183,N_1099,N_1086);
or U1184 (N_1184,N_1093,N_1125);
xnor U1185 (N_1185,N_1108,N_1111);
or U1186 (N_1186,N_1135,N_1138);
nand U1187 (N_1187,N_1134,N_1086);
nor U1188 (N_1188,N_1103,N_1094);
nand U1189 (N_1189,N_1127,N_1132);
or U1190 (N_1190,N_1122,N_1121);
nand U1191 (N_1191,N_1110,N_1111);
or U1192 (N_1192,N_1096,N_1101);
and U1193 (N_1193,N_1121,N_1094);
and U1194 (N_1194,N_1119,N_1136);
nor U1195 (N_1195,N_1109,N_1085);
nand U1196 (N_1196,N_1125,N_1108);
and U1197 (N_1197,N_1137,N_1100);
nand U1198 (N_1198,N_1084,N_1134);
and U1199 (N_1199,N_1135,N_1082);
nand U1200 (N_1200,N_1146,N_1173);
and U1201 (N_1201,N_1163,N_1181);
or U1202 (N_1202,N_1148,N_1140);
nand U1203 (N_1203,N_1151,N_1195);
or U1204 (N_1204,N_1144,N_1157);
xor U1205 (N_1205,N_1165,N_1159);
nor U1206 (N_1206,N_1186,N_1197);
or U1207 (N_1207,N_1169,N_1149);
or U1208 (N_1208,N_1188,N_1193);
or U1209 (N_1209,N_1199,N_1168);
nor U1210 (N_1210,N_1166,N_1187);
nand U1211 (N_1211,N_1191,N_1198);
and U1212 (N_1212,N_1171,N_1179);
nand U1213 (N_1213,N_1194,N_1177);
or U1214 (N_1214,N_1189,N_1190);
and U1215 (N_1215,N_1172,N_1180);
and U1216 (N_1216,N_1156,N_1160);
nor U1217 (N_1217,N_1143,N_1158);
nand U1218 (N_1218,N_1162,N_1152);
nor U1219 (N_1219,N_1184,N_1175);
nor U1220 (N_1220,N_1192,N_1147);
and U1221 (N_1221,N_1178,N_1196);
and U1222 (N_1222,N_1174,N_1176);
or U1223 (N_1223,N_1170,N_1183);
and U1224 (N_1224,N_1154,N_1182);
nor U1225 (N_1225,N_1164,N_1142);
nor U1226 (N_1226,N_1145,N_1153);
or U1227 (N_1227,N_1155,N_1141);
nor U1228 (N_1228,N_1167,N_1161);
and U1229 (N_1229,N_1185,N_1150);
or U1230 (N_1230,N_1143,N_1184);
xor U1231 (N_1231,N_1140,N_1163);
nor U1232 (N_1232,N_1165,N_1187);
nand U1233 (N_1233,N_1184,N_1155);
and U1234 (N_1234,N_1164,N_1157);
nor U1235 (N_1235,N_1167,N_1182);
nand U1236 (N_1236,N_1147,N_1170);
and U1237 (N_1237,N_1166,N_1151);
nand U1238 (N_1238,N_1194,N_1172);
or U1239 (N_1239,N_1141,N_1178);
nor U1240 (N_1240,N_1164,N_1160);
nor U1241 (N_1241,N_1168,N_1172);
nor U1242 (N_1242,N_1191,N_1196);
or U1243 (N_1243,N_1143,N_1153);
and U1244 (N_1244,N_1155,N_1181);
or U1245 (N_1245,N_1171,N_1143);
or U1246 (N_1246,N_1182,N_1180);
and U1247 (N_1247,N_1148,N_1156);
nor U1248 (N_1248,N_1187,N_1179);
nand U1249 (N_1249,N_1158,N_1157);
nor U1250 (N_1250,N_1162,N_1182);
nand U1251 (N_1251,N_1191,N_1185);
xor U1252 (N_1252,N_1158,N_1175);
or U1253 (N_1253,N_1175,N_1173);
or U1254 (N_1254,N_1186,N_1176);
or U1255 (N_1255,N_1172,N_1145);
nand U1256 (N_1256,N_1181,N_1144);
or U1257 (N_1257,N_1161,N_1183);
nand U1258 (N_1258,N_1199,N_1163);
nand U1259 (N_1259,N_1144,N_1175);
and U1260 (N_1260,N_1228,N_1258);
nand U1261 (N_1261,N_1214,N_1200);
nor U1262 (N_1262,N_1211,N_1247);
nand U1263 (N_1263,N_1234,N_1236);
or U1264 (N_1264,N_1210,N_1225);
or U1265 (N_1265,N_1242,N_1215);
or U1266 (N_1266,N_1237,N_1233);
nor U1267 (N_1267,N_1235,N_1259);
and U1268 (N_1268,N_1220,N_1240);
nand U1269 (N_1269,N_1222,N_1218);
nand U1270 (N_1270,N_1253,N_1206);
nor U1271 (N_1271,N_1232,N_1213);
nor U1272 (N_1272,N_1216,N_1241);
and U1273 (N_1273,N_1251,N_1255);
nor U1274 (N_1274,N_1202,N_1250);
or U1275 (N_1275,N_1203,N_1224);
nor U1276 (N_1276,N_1249,N_1238);
and U1277 (N_1277,N_1207,N_1205);
and U1278 (N_1278,N_1227,N_1254);
and U1279 (N_1279,N_1223,N_1221);
and U1280 (N_1280,N_1204,N_1201);
or U1281 (N_1281,N_1226,N_1212);
or U1282 (N_1282,N_1217,N_1231);
nand U1283 (N_1283,N_1245,N_1256);
nand U1284 (N_1284,N_1209,N_1248);
nor U1285 (N_1285,N_1257,N_1252);
xor U1286 (N_1286,N_1244,N_1219);
or U1287 (N_1287,N_1246,N_1243);
or U1288 (N_1288,N_1239,N_1230);
nor U1289 (N_1289,N_1208,N_1229);
nor U1290 (N_1290,N_1216,N_1212);
or U1291 (N_1291,N_1233,N_1225);
or U1292 (N_1292,N_1250,N_1207);
and U1293 (N_1293,N_1259,N_1240);
nor U1294 (N_1294,N_1204,N_1219);
nand U1295 (N_1295,N_1249,N_1213);
and U1296 (N_1296,N_1233,N_1242);
and U1297 (N_1297,N_1225,N_1203);
nor U1298 (N_1298,N_1213,N_1227);
or U1299 (N_1299,N_1259,N_1242);
nand U1300 (N_1300,N_1235,N_1240);
nand U1301 (N_1301,N_1217,N_1244);
or U1302 (N_1302,N_1259,N_1239);
nand U1303 (N_1303,N_1234,N_1230);
or U1304 (N_1304,N_1247,N_1238);
and U1305 (N_1305,N_1208,N_1244);
nor U1306 (N_1306,N_1217,N_1247);
nand U1307 (N_1307,N_1211,N_1243);
nor U1308 (N_1308,N_1233,N_1208);
nand U1309 (N_1309,N_1224,N_1220);
or U1310 (N_1310,N_1245,N_1210);
nor U1311 (N_1311,N_1255,N_1252);
nor U1312 (N_1312,N_1219,N_1214);
nand U1313 (N_1313,N_1203,N_1206);
xnor U1314 (N_1314,N_1208,N_1235);
or U1315 (N_1315,N_1215,N_1209);
nor U1316 (N_1316,N_1213,N_1253);
nor U1317 (N_1317,N_1207,N_1230);
or U1318 (N_1318,N_1250,N_1234);
nor U1319 (N_1319,N_1223,N_1218);
and U1320 (N_1320,N_1264,N_1310);
nand U1321 (N_1321,N_1269,N_1303);
nand U1322 (N_1322,N_1272,N_1274);
nor U1323 (N_1323,N_1277,N_1291);
or U1324 (N_1324,N_1275,N_1305);
or U1325 (N_1325,N_1295,N_1287);
nor U1326 (N_1326,N_1286,N_1282);
or U1327 (N_1327,N_1319,N_1288);
nand U1328 (N_1328,N_1266,N_1297);
and U1329 (N_1329,N_1278,N_1315);
nor U1330 (N_1330,N_1284,N_1308);
and U1331 (N_1331,N_1317,N_1265);
nand U1332 (N_1332,N_1267,N_1281);
and U1333 (N_1333,N_1314,N_1268);
nor U1334 (N_1334,N_1307,N_1293);
nand U1335 (N_1335,N_1311,N_1271);
nor U1336 (N_1336,N_1273,N_1283);
nand U1337 (N_1337,N_1292,N_1300);
and U1338 (N_1338,N_1289,N_1261);
or U1339 (N_1339,N_1263,N_1306);
or U1340 (N_1340,N_1312,N_1313);
or U1341 (N_1341,N_1304,N_1299);
nor U1342 (N_1342,N_1298,N_1279);
nand U1343 (N_1343,N_1280,N_1285);
and U1344 (N_1344,N_1262,N_1294);
and U1345 (N_1345,N_1316,N_1301);
or U1346 (N_1346,N_1260,N_1290);
and U1347 (N_1347,N_1302,N_1318);
or U1348 (N_1348,N_1276,N_1270);
and U1349 (N_1349,N_1309,N_1296);
nor U1350 (N_1350,N_1273,N_1280);
nand U1351 (N_1351,N_1287,N_1313);
and U1352 (N_1352,N_1290,N_1265);
nor U1353 (N_1353,N_1279,N_1300);
xnor U1354 (N_1354,N_1307,N_1272);
and U1355 (N_1355,N_1297,N_1284);
nand U1356 (N_1356,N_1312,N_1314);
and U1357 (N_1357,N_1312,N_1303);
and U1358 (N_1358,N_1276,N_1278);
nor U1359 (N_1359,N_1309,N_1314);
and U1360 (N_1360,N_1309,N_1270);
nor U1361 (N_1361,N_1302,N_1274);
and U1362 (N_1362,N_1275,N_1260);
and U1363 (N_1363,N_1270,N_1277);
or U1364 (N_1364,N_1264,N_1276);
nor U1365 (N_1365,N_1311,N_1261);
nand U1366 (N_1366,N_1271,N_1261);
nand U1367 (N_1367,N_1292,N_1272);
nand U1368 (N_1368,N_1286,N_1262);
and U1369 (N_1369,N_1292,N_1277);
or U1370 (N_1370,N_1278,N_1293);
nor U1371 (N_1371,N_1268,N_1282);
or U1372 (N_1372,N_1300,N_1267);
or U1373 (N_1373,N_1313,N_1309);
or U1374 (N_1374,N_1261,N_1299);
nor U1375 (N_1375,N_1266,N_1294);
nor U1376 (N_1376,N_1275,N_1263);
nor U1377 (N_1377,N_1288,N_1293);
or U1378 (N_1378,N_1293,N_1315);
nand U1379 (N_1379,N_1284,N_1275);
or U1380 (N_1380,N_1370,N_1368);
or U1381 (N_1381,N_1330,N_1363);
and U1382 (N_1382,N_1357,N_1356);
nand U1383 (N_1383,N_1339,N_1372);
and U1384 (N_1384,N_1350,N_1353);
nand U1385 (N_1385,N_1343,N_1348);
nor U1386 (N_1386,N_1347,N_1352);
nor U1387 (N_1387,N_1375,N_1334);
and U1388 (N_1388,N_1336,N_1324);
nor U1389 (N_1389,N_1361,N_1323);
and U1390 (N_1390,N_1367,N_1364);
nand U1391 (N_1391,N_1340,N_1329);
and U1392 (N_1392,N_1355,N_1365);
or U1393 (N_1393,N_1335,N_1354);
and U1394 (N_1394,N_1362,N_1321);
nor U1395 (N_1395,N_1337,N_1320);
nand U1396 (N_1396,N_1351,N_1333);
nor U1397 (N_1397,N_1374,N_1345);
xnor U1398 (N_1398,N_1371,N_1373);
nand U1399 (N_1399,N_1360,N_1359);
or U1400 (N_1400,N_1366,N_1322);
and U1401 (N_1401,N_1338,N_1349);
or U1402 (N_1402,N_1377,N_1328);
and U1403 (N_1403,N_1332,N_1376);
xnor U1404 (N_1404,N_1341,N_1378);
nor U1405 (N_1405,N_1358,N_1344);
and U1406 (N_1406,N_1326,N_1327);
and U1407 (N_1407,N_1369,N_1342);
or U1408 (N_1408,N_1346,N_1325);
or U1409 (N_1409,N_1331,N_1379);
or U1410 (N_1410,N_1339,N_1357);
or U1411 (N_1411,N_1354,N_1349);
or U1412 (N_1412,N_1375,N_1329);
or U1413 (N_1413,N_1357,N_1320);
nand U1414 (N_1414,N_1369,N_1346);
and U1415 (N_1415,N_1342,N_1374);
nand U1416 (N_1416,N_1361,N_1364);
and U1417 (N_1417,N_1365,N_1338);
and U1418 (N_1418,N_1320,N_1378);
or U1419 (N_1419,N_1373,N_1330);
and U1420 (N_1420,N_1372,N_1348);
or U1421 (N_1421,N_1342,N_1336);
nand U1422 (N_1422,N_1378,N_1342);
nor U1423 (N_1423,N_1328,N_1371);
or U1424 (N_1424,N_1320,N_1348);
nand U1425 (N_1425,N_1323,N_1354);
nor U1426 (N_1426,N_1348,N_1358);
nor U1427 (N_1427,N_1371,N_1330);
xnor U1428 (N_1428,N_1378,N_1351);
nor U1429 (N_1429,N_1339,N_1338);
nor U1430 (N_1430,N_1339,N_1362);
nor U1431 (N_1431,N_1321,N_1331);
and U1432 (N_1432,N_1363,N_1372);
nor U1433 (N_1433,N_1361,N_1339);
nand U1434 (N_1434,N_1337,N_1321);
and U1435 (N_1435,N_1366,N_1350);
xnor U1436 (N_1436,N_1368,N_1361);
and U1437 (N_1437,N_1357,N_1334);
xnor U1438 (N_1438,N_1365,N_1362);
nand U1439 (N_1439,N_1341,N_1348);
nand U1440 (N_1440,N_1407,N_1437);
nor U1441 (N_1441,N_1409,N_1403);
nand U1442 (N_1442,N_1384,N_1383);
or U1443 (N_1443,N_1423,N_1387);
and U1444 (N_1444,N_1392,N_1404);
nand U1445 (N_1445,N_1410,N_1411);
or U1446 (N_1446,N_1434,N_1412);
or U1447 (N_1447,N_1414,N_1395);
and U1448 (N_1448,N_1432,N_1430);
xnor U1449 (N_1449,N_1408,N_1426);
nand U1450 (N_1450,N_1381,N_1431);
or U1451 (N_1451,N_1401,N_1391);
or U1452 (N_1452,N_1424,N_1402);
nor U1453 (N_1453,N_1405,N_1422);
or U1454 (N_1454,N_1386,N_1419);
and U1455 (N_1455,N_1425,N_1398);
nor U1456 (N_1456,N_1421,N_1389);
or U1457 (N_1457,N_1390,N_1406);
or U1458 (N_1458,N_1427,N_1385);
or U1459 (N_1459,N_1435,N_1418);
and U1460 (N_1460,N_1388,N_1380);
nor U1461 (N_1461,N_1413,N_1439);
or U1462 (N_1462,N_1400,N_1415);
or U1463 (N_1463,N_1429,N_1382);
nand U1464 (N_1464,N_1399,N_1396);
nor U1465 (N_1465,N_1428,N_1394);
nand U1466 (N_1466,N_1393,N_1436);
or U1467 (N_1467,N_1397,N_1438);
nor U1468 (N_1468,N_1416,N_1433);
nand U1469 (N_1469,N_1417,N_1420);
and U1470 (N_1470,N_1404,N_1399);
or U1471 (N_1471,N_1382,N_1412);
and U1472 (N_1472,N_1382,N_1413);
and U1473 (N_1473,N_1439,N_1381);
nand U1474 (N_1474,N_1390,N_1428);
and U1475 (N_1475,N_1439,N_1405);
nor U1476 (N_1476,N_1402,N_1380);
nand U1477 (N_1477,N_1402,N_1407);
nor U1478 (N_1478,N_1382,N_1414);
nor U1479 (N_1479,N_1384,N_1410);
and U1480 (N_1480,N_1398,N_1429);
nand U1481 (N_1481,N_1391,N_1389);
and U1482 (N_1482,N_1431,N_1410);
nor U1483 (N_1483,N_1380,N_1413);
and U1484 (N_1484,N_1402,N_1385);
and U1485 (N_1485,N_1431,N_1411);
nand U1486 (N_1486,N_1414,N_1398);
nor U1487 (N_1487,N_1437,N_1428);
or U1488 (N_1488,N_1423,N_1391);
or U1489 (N_1489,N_1428,N_1384);
or U1490 (N_1490,N_1402,N_1408);
or U1491 (N_1491,N_1418,N_1395);
and U1492 (N_1492,N_1403,N_1388);
or U1493 (N_1493,N_1395,N_1425);
nand U1494 (N_1494,N_1435,N_1429);
nor U1495 (N_1495,N_1435,N_1421);
nand U1496 (N_1496,N_1420,N_1397);
or U1497 (N_1497,N_1408,N_1418);
nor U1498 (N_1498,N_1398,N_1391);
nor U1499 (N_1499,N_1416,N_1384);
or U1500 (N_1500,N_1446,N_1465);
and U1501 (N_1501,N_1447,N_1492);
and U1502 (N_1502,N_1493,N_1485);
nand U1503 (N_1503,N_1441,N_1451);
nor U1504 (N_1504,N_1498,N_1470);
nand U1505 (N_1505,N_1442,N_1483);
or U1506 (N_1506,N_1486,N_1478);
and U1507 (N_1507,N_1491,N_1489);
or U1508 (N_1508,N_1454,N_1496);
nand U1509 (N_1509,N_1448,N_1482);
nand U1510 (N_1510,N_1484,N_1449);
nand U1511 (N_1511,N_1461,N_1444);
or U1512 (N_1512,N_1453,N_1488);
nor U1513 (N_1513,N_1481,N_1445);
nor U1514 (N_1514,N_1463,N_1487);
nor U1515 (N_1515,N_1490,N_1452);
and U1516 (N_1516,N_1462,N_1499);
nor U1517 (N_1517,N_1459,N_1468);
nand U1518 (N_1518,N_1456,N_1443);
or U1519 (N_1519,N_1476,N_1497);
xor U1520 (N_1520,N_1477,N_1455);
and U1521 (N_1521,N_1458,N_1475);
or U1522 (N_1522,N_1472,N_1474);
nor U1523 (N_1523,N_1450,N_1460);
nor U1524 (N_1524,N_1467,N_1473);
nor U1525 (N_1525,N_1469,N_1494);
nor U1526 (N_1526,N_1471,N_1479);
or U1527 (N_1527,N_1440,N_1457);
or U1528 (N_1528,N_1466,N_1495);
nor U1529 (N_1529,N_1480,N_1464);
nand U1530 (N_1530,N_1452,N_1466);
and U1531 (N_1531,N_1455,N_1469);
and U1532 (N_1532,N_1458,N_1486);
or U1533 (N_1533,N_1477,N_1459);
xor U1534 (N_1534,N_1446,N_1443);
or U1535 (N_1535,N_1477,N_1499);
and U1536 (N_1536,N_1444,N_1440);
nand U1537 (N_1537,N_1476,N_1480);
nor U1538 (N_1538,N_1466,N_1456);
nand U1539 (N_1539,N_1455,N_1445);
nand U1540 (N_1540,N_1479,N_1445);
and U1541 (N_1541,N_1444,N_1445);
nor U1542 (N_1542,N_1493,N_1472);
and U1543 (N_1543,N_1446,N_1481);
nand U1544 (N_1544,N_1495,N_1494);
nand U1545 (N_1545,N_1468,N_1490);
nor U1546 (N_1546,N_1474,N_1484);
nor U1547 (N_1547,N_1449,N_1480);
nor U1548 (N_1548,N_1460,N_1441);
xor U1549 (N_1549,N_1450,N_1462);
nor U1550 (N_1550,N_1449,N_1485);
and U1551 (N_1551,N_1469,N_1450);
nor U1552 (N_1552,N_1442,N_1445);
nor U1553 (N_1553,N_1465,N_1455);
or U1554 (N_1554,N_1460,N_1465);
nand U1555 (N_1555,N_1496,N_1443);
or U1556 (N_1556,N_1457,N_1480);
and U1557 (N_1557,N_1440,N_1482);
nand U1558 (N_1558,N_1450,N_1480);
nor U1559 (N_1559,N_1456,N_1499);
or U1560 (N_1560,N_1512,N_1523);
and U1561 (N_1561,N_1504,N_1553);
or U1562 (N_1562,N_1510,N_1539);
and U1563 (N_1563,N_1527,N_1524);
nor U1564 (N_1564,N_1516,N_1517);
nor U1565 (N_1565,N_1505,N_1546);
nor U1566 (N_1566,N_1548,N_1514);
and U1567 (N_1567,N_1531,N_1543);
nand U1568 (N_1568,N_1530,N_1511);
and U1569 (N_1569,N_1532,N_1515);
or U1570 (N_1570,N_1547,N_1555);
and U1571 (N_1571,N_1521,N_1501);
and U1572 (N_1572,N_1529,N_1526);
and U1573 (N_1573,N_1544,N_1519);
or U1574 (N_1574,N_1503,N_1533);
nand U1575 (N_1575,N_1535,N_1520);
nand U1576 (N_1576,N_1540,N_1513);
or U1577 (N_1577,N_1550,N_1525);
and U1578 (N_1578,N_1518,N_1554);
nand U1579 (N_1579,N_1522,N_1551);
or U1580 (N_1580,N_1506,N_1558);
or U1581 (N_1581,N_1538,N_1509);
nand U1582 (N_1582,N_1502,N_1500);
and U1583 (N_1583,N_1541,N_1528);
and U1584 (N_1584,N_1552,N_1537);
and U1585 (N_1585,N_1542,N_1557);
nor U1586 (N_1586,N_1556,N_1536);
nand U1587 (N_1587,N_1549,N_1507);
and U1588 (N_1588,N_1559,N_1534);
nor U1589 (N_1589,N_1508,N_1545);
nand U1590 (N_1590,N_1559,N_1556);
or U1591 (N_1591,N_1512,N_1526);
and U1592 (N_1592,N_1530,N_1516);
and U1593 (N_1593,N_1527,N_1550);
and U1594 (N_1594,N_1501,N_1554);
nor U1595 (N_1595,N_1525,N_1512);
nand U1596 (N_1596,N_1555,N_1504);
nand U1597 (N_1597,N_1558,N_1523);
or U1598 (N_1598,N_1537,N_1500);
or U1599 (N_1599,N_1517,N_1543);
or U1600 (N_1600,N_1516,N_1533);
nor U1601 (N_1601,N_1512,N_1502);
nor U1602 (N_1602,N_1538,N_1527);
nand U1603 (N_1603,N_1514,N_1508);
and U1604 (N_1604,N_1535,N_1508);
nand U1605 (N_1605,N_1546,N_1551);
and U1606 (N_1606,N_1555,N_1518);
and U1607 (N_1607,N_1527,N_1506);
or U1608 (N_1608,N_1537,N_1524);
nand U1609 (N_1609,N_1555,N_1557);
and U1610 (N_1610,N_1510,N_1527);
nand U1611 (N_1611,N_1514,N_1515);
or U1612 (N_1612,N_1524,N_1558);
and U1613 (N_1613,N_1504,N_1558);
nor U1614 (N_1614,N_1556,N_1528);
nand U1615 (N_1615,N_1506,N_1500);
xnor U1616 (N_1616,N_1548,N_1550);
nand U1617 (N_1617,N_1509,N_1558);
nand U1618 (N_1618,N_1533,N_1529);
nand U1619 (N_1619,N_1546,N_1545);
and U1620 (N_1620,N_1577,N_1604);
nand U1621 (N_1621,N_1591,N_1576);
or U1622 (N_1622,N_1578,N_1600);
nor U1623 (N_1623,N_1564,N_1562);
nand U1624 (N_1624,N_1613,N_1573);
and U1625 (N_1625,N_1584,N_1616);
nor U1626 (N_1626,N_1575,N_1595);
nand U1627 (N_1627,N_1614,N_1618);
and U1628 (N_1628,N_1572,N_1587);
nor U1629 (N_1629,N_1615,N_1592);
or U1630 (N_1630,N_1594,N_1561);
nor U1631 (N_1631,N_1571,N_1581);
or U1632 (N_1632,N_1606,N_1609);
or U1633 (N_1633,N_1588,N_1603);
or U1634 (N_1634,N_1590,N_1607);
and U1635 (N_1635,N_1566,N_1611);
and U1636 (N_1636,N_1593,N_1570);
or U1637 (N_1637,N_1596,N_1569);
nor U1638 (N_1638,N_1586,N_1574);
nand U1639 (N_1639,N_1568,N_1563);
or U1640 (N_1640,N_1567,N_1585);
nor U1641 (N_1641,N_1617,N_1598);
nand U1642 (N_1642,N_1619,N_1579);
nand U1643 (N_1643,N_1565,N_1560);
and U1644 (N_1644,N_1602,N_1612);
or U1645 (N_1645,N_1608,N_1597);
nand U1646 (N_1646,N_1589,N_1580);
nor U1647 (N_1647,N_1599,N_1610);
nor U1648 (N_1648,N_1582,N_1583);
and U1649 (N_1649,N_1605,N_1601);
nand U1650 (N_1650,N_1573,N_1611);
or U1651 (N_1651,N_1613,N_1601);
nor U1652 (N_1652,N_1612,N_1597);
and U1653 (N_1653,N_1569,N_1583);
and U1654 (N_1654,N_1605,N_1591);
or U1655 (N_1655,N_1603,N_1615);
and U1656 (N_1656,N_1582,N_1585);
nand U1657 (N_1657,N_1576,N_1614);
or U1658 (N_1658,N_1567,N_1595);
and U1659 (N_1659,N_1586,N_1577);
nand U1660 (N_1660,N_1580,N_1593);
or U1661 (N_1661,N_1591,N_1574);
nor U1662 (N_1662,N_1599,N_1573);
nor U1663 (N_1663,N_1568,N_1605);
nand U1664 (N_1664,N_1576,N_1599);
and U1665 (N_1665,N_1614,N_1582);
nand U1666 (N_1666,N_1602,N_1575);
and U1667 (N_1667,N_1574,N_1597);
and U1668 (N_1668,N_1583,N_1588);
nand U1669 (N_1669,N_1598,N_1581);
and U1670 (N_1670,N_1599,N_1605);
and U1671 (N_1671,N_1590,N_1617);
or U1672 (N_1672,N_1589,N_1591);
or U1673 (N_1673,N_1614,N_1603);
nor U1674 (N_1674,N_1567,N_1571);
nor U1675 (N_1675,N_1611,N_1600);
nor U1676 (N_1676,N_1588,N_1587);
nor U1677 (N_1677,N_1617,N_1567);
and U1678 (N_1678,N_1571,N_1596);
or U1679 (N_1679,N_1593,N_1575);
and U1680 (N_1680,N_1677,N_1649);
and U1681 (N_1681,N_1636,N_1660);
and U1682 (N_1682,N_1628,N_1656);
nand U1683 (N_1683,N_1650,N_1674);
or U1684 (N_1684,N_1676,N_1666);
nor U1685 (N_1685,N_1642,N_1661);
or U1686 (N_1686,N_1626,N_1652);
nand U1687 (N_1687,N_1663,N_1655);
nand U1688 (N_1688,N_1673,N_1658);
nor U1689 (N_1689,N_1621,N_1669);
or U1690 (N_1690,N_1633,N_1664);
nand U1691 (N_1691,N_1647,N_1641);
nand U1692 (N_1692,N_1665,N_1635);
xnor U1693 (N_1693,N_1639,N_1625);
nand U1694 (N_1694,N_1645,N_1627);
xnor U1695 (N_1695,N_1653,N_1644);
xnor U1696 (N_1696,N_1657,N_1679);
nand U1697 (N_1697,N_1630,N_1624);
nor U1698 (N_1698,N_1622,N_1668);
and U1699 (N_1699,N_1643,N_1629);
and U1700 (N_1700,N_1638,N_1675);
nand U1701 (N_1701,N_1631,N_1637);
nand U1702 (N_1702,N_1654,N_1620);
nand U1703 (N_1703,N_1640,N_1634);
nand U1704 (N_1704,N_1632,N_1623);
nor U1705 (N_1705,N_1678,N_1670);
nor U1706 (N_1706,N_1646,N_1659);
nand U1707 (N_1707,N_1662,N_1651);
nand U1708 (N_1708,N_1671,N_1672);
and U1709 (N_1709,N_1648,N_1667);
nand U1710 (N_1710,N_1645,N_1677);
nand U1711 (N_1711,N_1650,N_1627);
nand U1712 (N_1712,N_1679,N_1643);
or U1713 (N_1713,N_1632,N_1643);
or U1714 (N_1714,N_1656,N_1630);
nand U1715 (N_1715,N_1650,N_1651);
or U1716 (N_1716,N_1640,N_1671);
nand U1717 (N_1717,N_1662,N_1656);
nor U1718 (N_1718,N_1645,N_1652);
or U1719 (N_1719,N_1654,N_1645);
nand U1720 (N_1720,N_1672,N_1640);
or U1721 (N_1721,N_1624,N_1646);
and U1722 (N_1722,N_1668,N_1623);
and U1723 (N_1723,N_1658,N_1640);
and U1724 (N_1724,N_1668,N_1624);
or U1725 (N_1725,N_1643,N_1677);
nand U1726 (N_1726,N_1635,N_1663);
xor U1727 (N_1727,N_1626,N_1647);
or U1728 (N_1728,N_1660,N_1663);
and U1729 (N_1729,N_1646,N_1647);
nand U1730 (N_1730,N_1632,N_1668);
or U1731 (N_1731,N_1667,N_1669);
or U1732 (N_1732,N_1658,N_1662);
nor U1733 (N_1733,N_1630,N_1640);
or U1734 (N_1734,N_1644,N_1624);
and U1735 (N_1735,N_1657,N_1649);
nor U1736 (N_1736,N_1628,N_1621);
or U1737 (N_1737,N_1661,N_1667);
nand U1738 (N_1738,N_1627,N_1640);
nor U1739 (N_1739,N_1655,N_1652);
and U1740 (N_1740,N_1716,N_1718);
nor U1741 (N_1741,N_1694,N_1728);
nor U1742 (N_1742,N_1703,N_1724);
nor U1743 (N_1743,N_1708,N_1702);
nand U1744 (N_1744,N_1693,N_1733);
nand U1745 (N_1745,N_1687,N_1723);
or U1746 (N_1746,N_1690,N_1699);
nor U1747 (N_1747,N_1732,N_1706);
or U1748 (N_1748,N_1695,N_1684);
nor U1749 (N_1749,N_1700,N_1726);
and U1750 (N_1750,N_1686,N_1707);
nand U1751 (N_1751,N_1709,N_1717);
and U1752 (N_1752,N_1688,N_1736);
or U1753 (N_1753,N_1701,N_1681);
or U1754 (N_1754,N_1720,N_1691);
xnor U1755 (N_1755,N_1725,N_1713);
or U1756 (N_1756,N_1731,N_1689);
nor U1757 (N_1757,N_1696,N_1738);
nor U1758 (N_1758,N_1722,N_1685);
and U1759 (N_1759,N_1680,N_1715);
or U1760 (N_1760,N_1729,N_1730);
or U1761 (N_1761,N_1735,N_1682);
nor U1762 (N_1762,N_1739,N_1719);
nand U1763 (N_1763,N_1721,N_1714);
and U1764 (N_1764,N_1698,N_1710);
nor U1765 (N_1765,N_1727,N_1712);
nand U1766 (N_1766,N_1711,N_1705);
nor U1767 (N_1767,N_1734,N_1737);
or U1768 (N_1768,N_1704,N_1683);
or U1769 (N_1769,N_1692,N_1697);
nor U1770 (N_1770,N_1723,N_1716);
nand U1771 (N_1771,N_1736,N_1685);
and U1772 (N_1772,N_1721,N_1686);
and U1773 (N_1773,N_1687,N_1728);
or U1774 (N_1774,N_1708,N_1697);
nand U1775 (N_1775,N_1717,N_1712);
and U1776 (N_1776,N_1714,N_1724);
or U1777 (N_1777,N_1714,N_1711);
and U1778 (N_1778,N_1681,N_1714);
xnor U1779 (N_1779,N_1739,N_1690);
nor U1780 (N_1780,N_1685,N_1708);
and U1781 (N_1781,N_1689,N_1697);
nand U1782 (N_1782,N_1715,N_1706);
xor U1783 (N_1783,N_1697,N_1704);
or U1784 (N_1784,N_1726,N_1683);
nand U1785 (N_1785,N_1702,N_1681);
and U1786 (N_1786,N_1726,N_1689);
xnor U1787 (N_1787,N_1708,N_1738);
and U1788 (N_1788,N_1737,N_1738);
nor U1789 (N_1789,N_1723,N_1708);
and U1790 (N_1790,N_1702,N_1695);
or U1791 (N_1791,N_1686,N_1711);
or U1792 (N_1792,N_1733,N_1686);
nor U1793 (N_1793,N_1694,N_1726);
or U1794 (N_1794,N_1703,N_1699);
or U1795 (N_1795,N_1683,N_1705);
nor U1796 (N_1796,N_1724,N_1730);
or U1797 (N_1797,N_1738,N_1680);
nor U1798 (N_1798,N_1698,N_1718);
nand U1799 (N_1799,N_1714,N_1734);
nand U1800 (N_1800,N_1746,N_1754);
and U1801 (N_1801,N_1748,N_1785);
and U1802 (N_1802,N_1788,N_1797);
nand U1803 (N_1803,N_1749,N_1796);
or U1804 (N_1804,N_1765,N_1751);
nor U1805 (N_1805,N_1758,N_1756);
and U1806 (N_1806,N_1787,N_1782);
or U1807 (N_1807,N_1742,N_1790);
or U1808 (N_1808,N_1743,N_1741);
or U1809 (N_1809,N_1763,N_1745);
nor U1810 (N_1810,N_1759,N_1783);
nor U1811 (N_1811,N_1773,N_1757);
nand U1812 (N_1812,N_1771,N_1791);
nor U1813 (N_1813,N_1781,N_1761);
and U1814 (N_1814,N_1755,N_1768);
or U1815 (N_1815,N_1752,N_1740);
and U1816 (N_1816,N_1760,N_1795);
nor U1817 (N_1817,N_1793,N_1753);
or U1818 (N_1818,N_1764,N_1780);
and U1819 (N_1819,N_1799,N_1775);
or U1820 (N_1820,N_1762,N_1798);
nor U1821 (N_1821,N_1772,N_1774);
nand U1822 (N_1822,N_1794,N_1778);
and U1823 (N_1823,N_1792,N_1784);
nor U1824 (N_1824,N_1769,N_1747);
and U1825 (N_1825,N_1767,N_1750);
or U1826 (N_1826,N_1776,N_1786);
nand U1827 (N_1827,N_1770,N_1777);
nor U1828 (N_1828,N_1766,N_1744);
nand U1829 (N_1829,N_1779,N_1789);
and U1830 (N_1830,N_1744,N_1760);
and U1831 (N_1831,N_1760,N_1764);
nor U1832 (N_1832,N_1777,N_1792);
nand U1833 (N_1833,N_1791,N_1745);
nand U1834 (N_1834,N_1787,N_1764);
nor U1835 (N_1835,N_1770,N_1799);
or U1836 (N_1836,N_1763,N_1772);
nor U1837 (N_1837,N_1770,N_1767);
and U1838 (N_1838,N_1769,N_1742);
or U1839 (N_1839,N_1742,N_1757);
nand U1840 (N_1840,N_1745,N_1741);
nand U1841 (N_1841,N_1763,N_1776);
nand U1842 (N_1842,N_1764,N_1773);
nor U1843 (N_1843,N_1771,N_1784);
nor U1844 (N_1844,N_1797,N_1768);
or U1845 (N_1845,N_1747,N_1751);
and U1846 (N_1846,N_1785,N_1789);
and U1847 (N_1847,N_1791,N_1755);
or U1848 (N_1848,N_1758,N_1750);
or U1849 (N_1849,N_1748,N_1794);
and U1850 (N_1850,N_1757,N_1772);
nor U1851 (N_1851,N_1761,N_1754);
and U1852 (N_1852,N_1755,N_1745);
and U1853 (N_1853,N_1770,N_1787);
or U1854 (N_1854,N_1773,N_1786);
nand U1855 (N_1855,N_1768,N_1748);
nand U1856 (N_1856,N_1767,N_1778);
or U1857 (N_1857,N_1757,N_1789);
xor U1858 (N_1858,N_1747,N_1785);
nand U1859 (N_1859,N_1781,N_1795);
nand U1860 (N_1860,N_1857,N_1801);
nor U1861 (N_1861,N_1838,N_1837);
or U1862 (N_1862,N_1819,N_1842);
or U1863 (N_1863,N_1804,N_1805);
or U1864 (N_1864,N_1828,N_1849);
and U1865 (N_1865,N_1813,N_1847);
and U1866 (N_1866,N_1846,N_1852);
or U1867 (N_1867,N_1803,N_1811);
nor U1868 (N_1868,N_1831,N_1839);
and U1869 (N_1869,N_1825,N_1844);
or U1870 (N_1870,N_1818,N_1823);
and U1871 (N_1871,N_1821,N_1817);
or U1872 (N_1872,N_1830,N_1824);
or U1873 (N_1873,N_1822,N_1806);
and U1874 (N_1874,N_1826,N_1845);
nand U1875 (N_1875,N_1835,N_1808);
and U1876 (N_1876,N_1851,N_1843);
nor U1877 (N_1877,N_1815,N_1848);
nor U1878 (N_1878,N_1859,N_1800);
nor U1879 (N_1879,N_1816,N_1858);
and U1880 (N_1880,N_1809,N_1856);
nor U1881 (N_1881,N_1812,N_1850);
nor U1882 (N_1882,N_1854,N_1832);
nand U1883 (N_1883,N_1802,N_1836);
and U1884 (N_1884,N_1829,N_1807);
or U1885 (N_1885,N_1820,N_1841);
nand U1886 (N_1886,N_1814,N_1834);
or U1887 (N_1887,N_1827,N_1833);
nor U1888 (N_1888,N_1810,N_1855);
nor U1889 (N_1889,N_1853,N_1840);
nor U1890 (N_1890,N_1804,N_1838);
and U1891 (N_1891,N_1855,N_1842);
nor U1892 (N_1892,N_1839,N_1852);
or U1893 (N_1893,N_1815,N_1826);
or U1894 (N_1894,N_1851,N_1813);
nand U1895 (N_1895,N_1825,N_1829);
and U1896 (N_1896,N_1809,N_1833);
nor U1897 (N_1897,N_1848,N_1810);
and U1898 (N_1898,N_1818,N_1833);
or U1899 (N_1899,N_1859,N_1830);
nor U1900 (N_1900,N_1821,N_1846);
nor U1901 (N_1901,N_1805,N_1854);
nor U1902 (N_1902,N_1822,N_1803);
and U1903 (N_1903,N_1859,N_1833);
or U1904 (N_1904,N_1852,N_1824);
nand U1905 (N_1905,N_1801,N_1834);
or U1906 (N_1906,N_1821,N_1848);
nand U1907 (N_1907,N_1822,N_1812);
or U1908 (N_1908,N_1841,N_1854);
nor U1909 (N_1909,N_1848,N_1802);
and U1910 (N_1910,N_1821,N_1859);
or U1911 (N_1911,N_1842,N_1834);
nor U1912 (N_1912,N_1830,N_1819);
or U1913 (N_1913,N_1823,N_1847);
and U1914 (N_1914,N_1825,N_1814);
and U1915 (N_1915,N_1828,N_1846);
nor U1916 (N_1916,N_1859,N_1849);
and U1917 (N_1917,N_1826,N_1831);
and U1918 (N_1918,N_1812,N_1807);
and U1919 (N_1919,N_1851,N_1831);
or U1920 (N_1920,N_1869,N_1864);
or U1921 (N_1921,N_1872,N_1902);
nor U1922 (N_1922,N_1880,N_1916);
and U1923 (N_1923,N_1882,N_1899);
or U1924 (N_1924,N_1877,N_1879);
or U1925 (N_1925,N_1918,N_1884);
xnor U1926 (N_1926,N_1863,N_1905);
and U1927 (N_1927,N_1890,N_1894);
nor U1928 (N_1928,N_1900,N_1910);
nand U1929 (N_1929,N_1909,N_1871);
nand U1930 (N_1930,N_1895,N_1913);
nor U1931 (N_1931,N_1891,N_1912);
or U1932 (N_1932,N_1887,N_1917);
and U1933 (N_1933,N_1875,N_1886);
and U1934 (N_1934,N_1873,N_1898);
and U1935 (N_1935,N_1881,N_1906);
nor U1936 (N_1936,N_1893,N_1885);
or U1937 (N_1937,N_1904,N_1876);
or U1938 (N_1938,N_1889,N_1874);
and U1939 (N_1939,N_1907,N_1870);
or U1940 (N_1940,N_1866,N_1892);
or U1941 (N_1941,N_1911,N_1908);
and U1942 (N_1942,N_1897,N_1865);
or U1943 (N_1943,N_1868,N_1901);
or U1944 (N_1944,N_1867,N_1888);
or U1945 (N_1945,N_1896,N_1861);
nor U1946 (N_1946,N_1860,N_1915);
or U1947 (N_1947,N_1914,N_1883);
or U1948 (N_1948,N_1862,N_1903);
nand U1949 (N_1949,N_1878,N_1919);
or U1950 (N_1950,N_1906,N_1876);
nor U1951 (N_1951,N_1917,N_1871);
nand U1952 (N_1952,N_1875,N_1901);
or U1953 (N_1953,N_1890,N_1896);
and U1954 (N_1954,N_1867,N_1899);
or U1955 (N_1955,N_1908,N_1861);
and U1956 (N_1956,N_1914,N_1861);
nand U1957 (N_1957,N_1860,N_1899);
nor U1958 (N_1958,N_1888,N_1899);
nor U1959 (N_1959,N_1912,N_1888);
and U1960 (N_1960,N_1893,N_1901);
or U1961 (N_1961,N_1886,N_1910);
or U1962 (N_1962,N_1877,N_1880);
or U1963 (N_1963,N_1886,N_1891);
or U1964 (N_1964,N_1874,N_1903);
nand U1965 (N_1965,N_1867,N_1895);
and U1966 (N_1966,N_1867,N_1889);
nor U1967 (N_1967,N_1870,N_1901);
nor U1968 (N_1968,N_1862,N_1911);
or U1969 (N_1969,N_1891,N_1880);
and U1970 (N_1970,N_1911,N_1885);
nor U1971 (N_1971,N_1861,N_1874);
or U1972 (N_1972,N_1868,N_1888);
or U1973 (N_1973,N_1877,N_1884);
nor U1974 (N_1974,N_1915,N_1872);
or U1975 (N_1975,N_1872,N_1917);
and U1976 (N_1976,N_1868,N_1897);
nor U1977 (N_1977,N_1917,N_1867);
nor U1978 (N_1978,N_1871,N_1890);
or U1979 (N_1979,N_1871,N_1872);
and U1980 (N_1980,N_1937,N_1928);
nand U1981 (N_1981,N_1966,N_1927);
and U1982 (N_1982,N_1933,N_1977);
or U1983 (N_1983,N_1969,N_1957);
nor U1984 (N_1984,N_1944,N_1955);
nand U1985 (N_1985,N_1922,N_1923);
nor U1986 (N_1986,N_1956,N_1968);
and U1987 (N_1987,N_1954,N_1963);
nand U1988 (N_1988,N_1949,N_1939);
or U1989 (N_1989,N_1967,N_1972);
or U1990 (N_1990,N_1935,N_1920);
nor U1991 (N_1991,N_1941,N_1930);
nand U1992 (N_1992,N_1960,N_1952);
or U1993 (N_1993,N_1946,N_1932);
nor U1994 (N_1994,N_1940,N_1961);
nand U1995 (N_1995,N_1974,N_1962);
nor U1996 (N_1996,N_1965,N_1943);
and U1997 (N_1997,N_1925,N_1948);
or U1998 (N_1998,N_1945,N_1973);
and U1999 (N_1999,N_1929,N_1931);
and U2000 (N_2000,N_1934,N_1921);
nor U2001 (N_2001,N_1971,N_1951);
nand U2002 (N_2002,N_1942,N_1938);
nand U2003 (N_2003,N_1979,N_1975);
nor U2004 (N_2004,N_1970,N_1964);
nor U2005 (N_2005,N_1936,N_1958);
nand U2006 (N_2006,N_1947,N_1953);
nand U2007 (N_2007,N_1978,N_1976);
or U2008 (N_2008,N_1926,N_1959);
nor U2009 (N_2009,N_1924,N_1950);
or U2010 (N_2010,N_1974,N_1950);
nor U2011 (N_2011,N_1956,N_1955);
nand U2012 (N_2012,N_1975,N_1966);
or U2013 (N_2013,N_1957,N_1930);
nand U2014 (N_2014,N_1935,N_1922);
nor U2015 (N_2015,N_1979,N_1956);
and U2016 (N_2016,N_1947,N_1928);
nor U2017 (N_2017,N_1928,N_1964);
or U2018 (N_2018,N_1942,N_1929);
nor U2019 (N_2019,N_1939,N_1976);
and U2020 (N_2020,N_1938,N_1963);
nor U2021 (N_2021,N_1945,N_1929);
and U2022 (N_2022,N_1960,N_1966);
and U2023 (N_2023,N_1922,N_1948);
nand U2024 (N_2024,N_1926,N_1976);
or U2025 (N_2025,N_1968,N_1940);
or U2026 (N_2026,N_1959,N_1949);
nor U2027 (N_2027,N_1976,N_1973);
and U2028 (N_2028,N_1964,N_1920);
nor U2029 (N_2029,N_1968,N_1979);
nand U2030 (N_2030,N_1970,N_1937);
nand U2031 (N_2031,N_1973,N_1940);
or U2032 (N_2032,N_1940,N_1921);
and U2033 (N_2033,N_1935,N_1970);
nor U2034 (N_2034,N_1967,N_1955);
and U2035 (N_2035,N_1943,N_1951);
or U2036 (N_2036,N_1940,N_1927);
nor U2037 (N_2037,N_1929,N_1947);
nand U2038 (N_2038,N_1934,N_1965);
and U2039 (N_2039,N_1925,N_1968);
and U2040 (N_2040,N_2007,N_2030);
and U2041 (N_2041,N_1987,N_2022);
nand U2042 (N_2042,N_2027,N_2036);
or U2043 (N_2043,N_2011,N_1989);
and U2044 (N_2044,N_2039,N_1999);
nand U2045 (N_2045,N_2033,N_2019);
and U2046 (N_2046,N_2023,N_2035);
nor U2047 (N_2047,N_2002,N_1988);
and U2048 (N_2048,N_1984,N_1994);
and U2049 (N_2049,N_2018,N_1998);
and U2050 (N_2050,N_1993,N_1997);
nor U2051 (N_2051,N_2032,N_2038);
nand U2052 (N_2052,N_1982,N_2029);
nor U2053 (N_2053,N_2013,N_2021);
or U2054 (N_2054,N_2010,N_1996);
nand U2055 (N_2055,N_2003,N_1985);
or U2056 (N_2056,N_2020,N_2037);
nand U2057 (N_2057,N_2026,N_2009);
and U2058 (N_2058,N_2000,N_2014);
nand U2059 (N_2059,N_2031,N_1981);
or U2060 (N_2060,N_2024,N_2004);
and U2061 (N_2061,N_1983,N_2034);
or U2062 (N_2062,N_2016,N_1986);
nor U2063 (N_2063,N_2015,N_2008);
xor U2064 (N_2064,N_1991,N_1992);
nand U2065 (N_2065,N_2017,N_2005);
nor U2066 (N_2066,N_2012,N_1980);
nand U2067 (N_2067,N_2006,N_2001);
or U2068 (N_2068,N_2025,N_1990);
nor U2069 (N_2069,N_1995,N_2028);
and U2070 (N_2070,N_1981,N_2016);
and U2071 (N_2071,N_1991,N_2017);
nor U2072 (N_2072,N_1995,N_2020);
nand U2073 (N_2073,N_2036,N_1987);
nand U2074 (N_2074,N_2006,N_2026);
nor U2075 (N_2075,N_2016,N_2015);
or U2076 (N_2076,N_2029,N_1993);
and U2077 (N_2077,N_1986,N_1985);
or U2078 (N_2078,N_1994,N_2027);
nand U2079 (N_2079,N_1990,N_2011);
nor U2080 (N_2080,N_2035,N_2013);
nor U2081 (N_2081,N_2003,N_2006);
and U2082 (N_2082,N_2034,N_1999);
and U2083 (N_2083,N_2028,N_2029);
or U2084 (N_2084,N_2026,N_2034);
nand U2085 (N_2085,N_2009,N_1998);
and U2086 (N_2086,N_1986,N_1982);
and U2087 (N_2087,N_1996,N_2005);
and U2088 (N_2088,N_1985,N_2034);
or U2089 (N_2089,N_2025,N_2033);
and U2090 (N_2090,N_1994,N_2002);
or U2091 (N_2091,N_2011,N_1995);
xor U2092 (N_2092,N_2038,N_2010);
nor U2093 (N_2093,N_2032,N_2037);
and U2094 (N_2094,N_2000,N_1982);
nor U2095 (N_2095,N_2018,N_2029);
xnor U2096 (N_2096,N_2030,N_1992);
nand U2097 (N_2097,N_2007,N_2000);
or U2098 (N_2098,N_2014,N_2026);
nor U2099 (N_2099,N_1999,N_2031);
or U2100 (N_2100,N_2061,N_2065);
nand U2101 (N_2101,N_2095,N_2040);
nor U2102 (N_2102,N_2062,N_2052);
or U2103 (N_2103,N_2093,N_2086);
nor U2104 (N_2104,N_2048,N_2078);
and U2105 (N_2105,N_2057,N_2077);
xor U2106 (N_2106,N_2064,N_2092);
nor U2107 (N_2107,N_2050,N_2084);
or U2108 (N_2108,N_2081,N_2041);
and U2109 (N_2109,N_2045,N_2071);
or U2110 (N_2110,N_2066,N_2067);
nor U2111 (N_2111,N_2051,N_2094);
nor U2112 (N_2112,N_2080,N_2089);
or U2113 (N_2113,N_2072,N_2096);
or U2114 (N_2114,N_2070,N_2083);
nor U2115 (N_2115,N_2063,N_2069);
or U2116 (N_2116,N_2049,N_2044);
nand U2117 (N_2117,N_2068,N_2099);
nand U2118 (N_2118,N_2091,N_2055);
nand U2119 (N_2119,N_2087,N_2079);
nand U2120 (N_2120,N_2053,N_2090);
nor U2121 (N_2121,N_2054,N_2073);
and U2122 (N_2122,N_2059,N_2058);
nor U2123 (N_2123,N_2047,N_2097);
and U2124 (N_2124,N_2074,N_2088);
xnor U2125 (N_2125,N_2043,N_2075);
nand U2126 (N_2126,N_2042,N_2085);
nor U2127 (N_2127,N_2060,N_2046);
nor U2128 (N_2128,N_2098,N_2056);
nor U2129 (N_2129,N_2082,N_2076);
or U2130 (N_2130,N_2043,N_2057);
nor U2131 (N_2131,N_2071,N_2057);
or U2132 (N_2132,N_2066,N_2077);
and U2133 (N_2133,N_2042,N_2046);
or U2134 (N_2134,N_2074,N_2097);
nand U2135 (N_2135,N_2057,N_2081);
or U2136 (N_2136,N_2042,N_2078);
nand U2137 (N_2137,N_2081,N_2046);
nand U2138 (N_2138,N_2099,N_2067);
xnor U2139 (N_2139,N_2092,N_2097);
or U2140 (N_2140,N_2075,N_2066);
or U2141 (N_2141,N_2083,N_2065);
and U2142 (N_2142,N_2094,N_2075);
nand U2143 (N_2143,N_2068,N_2042);
nor U2144 (N_2144,N_2074,N_2071);
nand U2145 (N_2145,N_2090,N_2062);
or U2146 (N_2146,N_2071,N_2099);
nor U2147 (N_2147,N_2078,N_2082);
nand U2148 (N_2148,N_2086,N_2057);
and U2149 (N_2149,N_2059,N_2071);
nand U2150 (N_2150,N_2097,N_2050);
nand U2151 (N_2151,N_2068,N_2085);
nand U2152 (N_2152,N_2088,N_2069);
nor U2153 (N_2153,N_2052,N_2041);
or U2154 (N_2154,N_2092,N_2087);
nand U2155 (N_2155,N_2091,N_2060);
and U2156 (N_2156,N_2044,N_2062);
nand U2157 (N_2157,N_2060,N_2074);
or U2158 (N_2158,N_2062,N_2084);
or U2159 (N_2159,N_2096,N_2079);
nor U2160 (N_2160,N_2112,N_2152);
and U2161 (N_2161,N_2107,N_2106);
xnor U2162 (N_2162,N_2148,N_2133);
and U2163 (N_2163,N_2124,N_2109);
nand U2164 (N_2164,N_2121,N_2117);
nand U2165 (N_2165,N_2120,N_2111);
nand U2166 (N_2166,N_2108,N_2140);
nor U2167 (N_2167,N_2144,N_2126);
or U2168 (N_2168,N_2116,N_2142);
xnor U2169 (N_2169,N_2123,N_2115);
xor U2170 (N_2170,N_2105,N_2128);
nor U2171 (N_2171,N_2157,N_2129);
or U2172 (N_2172,N_2134,N_2127);
and U2173 (N_2173,N_2122,N_2143);
and U2174 (N_2174,N_2132,N_2138);
and U2175 (N_2175,N_2154,N_2159);
nor U2176 (N_2176,N_2113,N_2118);
or U2177 (N_2177,N_2125,N_2139);
nor U2178 (N_2178,N_2151,N_2137);
nand U2179 (N_2179,N_2130,N_2136);
nand U2180 (N_2180,N_2103,N_2146);
nand U2181 (N_2181,N_2141,N_2153);
nand U2182 (N_2182,N_2131,N_2155);
or U2183 (N_2183,N_2158,N_2114);
nand U2184 (N_2184,N_2147,N_2156);
and U2185 (N_2185,N_2149,N_2102);
and U2186 (N_2186,N_2100,N_2104);
and U2187 (N_2187,N_2150,N_2110);
nor U2188 (N_2188,N_2101,N_2119);
xor U2189 (N_2189,N_2135,N_2145);
and U2190 (N_2190,N_2100,N_2126);
or U2191 (N_2191,N_2126,N_2121);
and U2192 (N_2192,N_2103,N_2117);
nor U2193 (N_2193,N_2107,N_2145);
nor U2194 (N_2194,N_2123,N_2122);
nor U2195 (N_2195,N_2115,N_2112);
or U2196 (N_2196,N_2149,N_2142);
nand U2197 (N_2197,N_2138,N_2129);
nor U2198 (N_2198,N_2102,N_2159);
and U2199 (N_2199,N_2102,N_2142);
nor U2200 (N_2200,N_2122,N_2129);
and U2201 (N_2201,N_2153,N_2149);
or U2202 (N_2202,N_2145,N_2127);
or U2203 (N_2203,N_2135,N_2156);
and U2204 (N_2204,N_2154,N_2120);
nand U2205 (N_2205,N_2129,N_2135);
nor U2206 (N_2206,N_2155,N_2126);
and U2207 (N_2207,N_2103,N_2123);
nor U2208 (N_2208,N_2131,N_2112);
nand U2209 (N_2209,N_2129,N_2143);
or U2210 (N_2210,N_2157,N_2142);
and U2211 (N_2211,N_2153,N_2144);
or U2212 (N_2212,N_2154,N_2111);
xnor U2213 (N_2213,N_2131,N_2136);
nor U2214 (N_2214,N_2130,N_2109);
and U2215 (N_2215,N_2106,N_2135);
and U2216 (N_2216,N_2136,N_2129);
and U2217 (N_2217,N_2138,N_2143);
or U2218 (N_2218,N_2123,N_2135);
nand U2219 (N_2219,N_2126,N_2152);
or U2220 (N_2220,N_2175,N_2160);
nand U2221 (N_2221,N_2182,N_2206);
or U2222 (N_2222,N_2202,N_2218);
nand U2223 (N_2223,N_2167,N_2191);
and U2224 (N_2224,N_2181,N_2165);
xnor U2225 (N_2225,N_2207,N_2163);
and U2226 (N_2226,N_2192,N_2170);
nand U2227 (N_2227,N_2174,N_2214);
nand U2228 (N_2228,N_2186,N_2194);
or U2229 (N_2229,N_2193,N_2180);
nor U2230 (N_2230,N_2213,N_2184);
or U2231 (N_2231,N_2173,N_2187);
nand U2232 (N_2232,N_2161,N_2201);
nor U2233 (N_2233,N_2204,N_2189);
or U2234 (N_2234,N_2169,N_2166);
nand U2235 (N_2235,N_2176,N_2208);
nand U2236 (N_2236,N_2200,N_2183);
or U2237 (N_2237,N_2162,N_2199);
nand U2238 (N_2238,N_2209,N_2177);
and U2239 (N_2239,N_2185,N_2195);
nand U2240 (N_2240,N_2217,N_2196);
and U2241 (N_2241,N_2172,N_2216);
nor U2242 (N_2242,N_2164,N_2210);
nor U2243 (N_2243,N_2219,N_2203);
xor U2244 (N_2244,N_2168,N_2190);
nand U2245 (N_2245,N_2205,N_2212);
or U2246 (N_2246,N_2198,N_2179);
nor U2247 (N_2247,N_2215,N_2188);
or U2248 (N_2248,N_2211,N_2178);
or U2249 (N_2249,N_2171,N_2197);
nand U2250 (N_2250,N_2197,N_2200);
nand U2251 (N_2251,N_2213,N_2204);
and U2252 (N_2252,N_2168,N_2196);
nor U2253 (N_2253,N_2205,N_2202);
or U2254 (N_2254,N_2182,N_2208);
or U2255 (N_2255,N_2169,N_2200);
and U2256 (N_2256,N_2173,N_2172);
nand U2257 (N_2257,N_2187,N_2169);
or U2258 (N_2258,N_2167,N_2171);
or U2259 (N_2259,N_2182,N_2168);
and U2260 (N_2260,N_2180,N_2214);
xnor U2261 (N_2261,N_2187,N_2188);
or U2262 (N_2262,N_2214,N_2216);
nand U2263 (N_2263,N_2170,N_2175);
xor U2264 (N_2264,N_2217,N_2175);
nor U2265 (N_2265,N_2212,N_2188);
nor U2266 (N_2266,N_2206,N_2194);
nor U2267 (N_2267,N_2182,N_2165);
and U2268 (N_2268,N_2184,N_2182);
nand U2269 (N_2269,N_2192,N_2213);
and U2270 (N_2270,N_2189,N_2182);
nand U2271 (N_2271,N_2183,N_2194);
nand U2272 (N_2272,N_2161,N_2170);
or U2273 (N_2273,N_2204,N_2191);
or U2274 (N_2274,N_2181,N_2176);
or U2275 (N_2275,N_2172,N_2160);
and U2276 (N_2276,N_2160,N_2212);
and U2277 (N_2277,N_2178,N_2172);
and U2278 (N_2278,N_2207,N_2200);
or U2279 (N_2279,N_2187,N_2172);
or U2280 (N_2280,N_2258,N_2274);
or U2281 (N_2281,N_2257,N_2236);
nor U2282 (N_2282,N_2233,N_2265);
and U2283 (N_2283,N_2238,N_2264);
nand U2284 (N_2284,N_2247,N_2271);
and U2285 (N_2285,N_2250,N_2249);
nand U2286 (N_2286,N_2246,N_2256);
and U2287 (N_2287,N_2253,N_2251);
nand U2288 (N_2288,N_2228,N_2227);
and U2289 (N_2289,N_2259,N_2273);
nand U2290 (N_2290,N_2268,N_2275);
xor U2291 (N_2291,N_2267,N_2254);
xnor U2292 (N_2292,N_2220,N_2272);
and U2293 (N_2293,N_2239,N_2261);
or U2294 (N_2294,N_2276,N_2252);
xor U2295 (N_2295,N_2240,N_2255);
nor U2296 (N_2296,N_2278,N_2245);
nand U2297 (N_2297,N_2237,N_2221);
nor U2298 (N_2298,N_2222,N_2263);
nand U2299 (N_2299,N_2235,N_2231);
or U2300 (N_2300,N_2223,N_2243);
nand U2301 (N_2301,N_2226,N_2229);
nand U2302 (N_2302,N_2230,N_2277);
and U2303 (N_2303,N_2232,N_2260);
nand U2304 (N_2304,N_2234,N_2244);
nor U2305 (N_2305,N_2270,N_2241);
nor U2306 (N_2306,N_2224,N_2242);
or U2307 (N_2307,N_2262,N_2266);
nand U2308 (N_2308,N_2279,N_2269);
nor U2309 (N_2309,N_2225,N_2248);
or U2310 (N_2310,N_2233,N_2230);
or U2311 (N_2311,N_2236,N_2279);
and U2312 (N_2312,N_2232,N_2266);
nand U2313 (N_2313,N_2274,N_2231);
xor U2314 (N_2314,N_2247,N_2233);
nor U2315 (N_2315,N_2272,N_2258);
nor U2316 (N_2316,N_2249,N_2223);
nand U2317 (N_2317,N_2272,N_2273);
and U2318 (N_2318,N_2279,N_2276);
nor U2319 (N_2319,N_2257,N_2222);
nand U2320 (N_2320,N_2254,N_2239);
or U2321 (N_2321,N_2249,N_2252);
nand U2322 (N_2322,N_2252,N_2227);
or U2323 (N_2323,N_2242,N_2221);
nand U2324 (N_2324,N_2224,N_2236);
and U2325 (N_2325,N_2257,N_2221);
nor U2326 (N_2326,N_2227,N_2236);
or U2327 (N_2327,N_2273,N_2221);
or U2328 (N_2328,N_2246,N_2251);
nor U2329 (N_2329,N_2223,N_2226);
nor U2330 (N_2330,N_2232,N_2259);
and U2331 (N_2331,N_2225,N_2220);
or U2332 (N_2332,N_2248,N_2265);
or U2333 (N_2333,N_2254,N_2231);
nor U2334 (N_2334,N_2245,N_2255);
or U2335 (N_2335,N_2234,N_2225);
and U2336 (N_2336,N_2243,N_2240);
or U2337 (N_2337,N_2234,N_2256);
and U2338 (N_2338,N_2266,N_2252);
nand U2339 (N_2339,N_2241,N_2237);
nor U2340 (N_2340,N_2326,N_2318);
nor U2341 (N_2341,N_2295,N_2308);
or U2342 (N_2342,N_2306,N_2319);
nand U2343 (N_2343,N_2324,N_2290);
or U2344 (N_2344,N_2285,N_2315);
and U2345 (N_2345,N_2333,N_2304);
or U2346 (N_2346,N_2288,N_2312);
or U2347 (N_2347,N_2314,N_2300);
or U2348 (N_2348,N_2331,N_2296);
and U2349 (N_2349,N_2320,N_2298);
xor U2350 (N_2350,N_2284,N_2283);
nor U2351 (N_2351,N_2328,N_2286);
nand U2352 (N_2352,N_2281,N_2307);
and U2353 (N_2353,N_2301,N_2303);
or U2354 (N_2354,N_2310,N_2321);
nor U2355 (N_2355,N_2287,N_2280);
and U2356 (N_2356,N_2332,N_2313);
and U2357 (N_2357,N_2322,N_2338);
and U2358 (N_2358,N_2311,N_2335);
nor U2359 (N_2359,N_2299,N_2291);
nor U2360 (N_2360,N_2294,N_2305);
or U2361 (N_2361,N_2302,N_2297);
nand U2362 (N_2362,N_2330,N_2337);
or U2363 (N_2363,N_2282,N_2334);
nand U2364 (N_2364,N_2292,N_2293);
and U2365 (N_2365,N_2309,N_2325);
or U2366 (N_2366,N_2289,N_2336);
and U2367 (N_2367,N_2327,N_2317);
nor U2368 (N_2368,N_2339,N_2316);
or U2369 (N_2369,N_2323,N_2329);
and U2370 (N_2370,N_2287,N_2311);
or U2371 (N_2371,N_2290,N_2287);
or U2372 (N_2372,N_2291,N_2282);
and U2373 (N_2373,N_2292,N_2323);
or U2374 (N_2374,N_2317,N_2315);
and U2375 (N_2375,N_2336,N_2298);
nor U2376 (N_2376,N_2332,N_2315);
nand U2377 (N_2377,N_2314,N_2335);
nand U2378 (N_2378,N_2284,N_2333);
nand U2379 (N_2379,N_2310,N_2289);
nand U2380 (N_2380,N_2310,N_2285);
nand U2381 (N_2381,N_2282,N_2317);
nor U2382 (N_2382,N_2288,N_2322);
or U2383 (N_2383,N_2323,N_2339);
nor U2384 (N_2384,N_2322,N_2321);
nand U2385 (N_2385,N_2280,N_2309);
and U2386 (N_2386,N_2285,N_2295);
and U2387 (N_2387,N_2330,N_2315);
nand U2388 (N_2388,N_2335,N_2288);
or U2389 (N_2389,N_2302,N_2326);
nor U2390 (N_2390,N_2297,N_2291);
or U2391 (N_2391,N_2311,N_2292);
or U2392 (N_2392,N_2331,N_2293);
nand U2393 (N_2393,N_2334,N_2304);
nand U2394 (N_2394,N_2302,N_2303);
or U2395 (N_2395,N_2314,N_2326);
or U2396 (N_2396,N_2292,N_2319);
nor U2397 (N_2397,N_2285,N_2303);
or U2398 (N_2398,N_2314,N_2315);
or U2399 (N_2399,N_2305,N_2320);
nand U2400 (N_2400,N_2386,N_2356);
or U2401 (N_2401,N_2343,N_2352);
nor U2402 (N_2402,N_2397,N_2366);
or U2403 (N_2403,N_2360,N_2382);
and U2404 (N_2404,N_2381,N_2383);
or U2405 (N_2405,N_2374,N_2398);
nand U2406 (N_2406,N_2377,N_2373);
nor U2407 (N_2407,N_2384,N_2362);
nand U2408 (N_2408,N_2393,N_2368);
nor U2409 (N_2409,N_2378,N_2376);
nor U2410 (N_2410,N_2353,N_2396);
nor U2411 (N_2411,N_2385,N_2371);
nand U2412 (N_2412,N_2387,N_2344);
nor U2413 (N_2413,N_2375,N_2367);
nor U2414 (N_2414,N_2369,N_2363);
and U2415 (N_2415,N_2342,N_2390);
nor U2416 (N_2416,N_2394,N_2341);
and U2417 (N_2417,N_2348,N_2351);
nand U2418 (N_2418,N_2391,N_2361);
nor U2419 (N_2419,N_2379,N_2372);
nor U2420 (N_2420,N_2388,N_2340);
nor U2421 (N_2421,N_2395,N_2365);
and U2422 (N_2422,N_2354,N_2392);
nand U2423 (N_2423,N_2389,N_2358);
and U2424 (N_2424,N_2399,N_2349);
xnor U2425 (N_2425,N_2364,N_2359);
and U2426 (N_2426,N_2355,N_2347);
or U2427 (N_2427,N_2350,N_2345);
or U2428 (N_2428,N_2346,N_2380);
nor U2429 (N_2429,N_2357,N_2370);
nand U2430 (N_2430,N_2344,N_2346);
and U2431 (N_2431,N_2372,N_2352);
nor U2432 (N_2432,N_2371,N_2381);
or U2433 (N_2433,N_2379,N_2373);
or U2434 (N_2434,N_2363,N_2350);
or U2435 (N_2435,N_2360,N_2374);
nand U2436 (N_2436,N_2355,N_2392);
nand U2437 (N_2437,N_2386,N_2385);
nor U2438 (N_2438,N_2346,N_2379);
or U2439 (N_2439,N_2348,N_2388);
nor U2440 (N_2440,N_2340,N_2394);
nand U2441 (N_2441,N_2369,N_2355);
and U2442 (N_2442,N_2356,N_2352);
xnor U2443 (N_2443,N_2355,N_2372);
nor U2444 (N_2444,N_2343,N_2358);
and U2445 (N_2445,N_2385,N_2377);
and U2446 (N_2446,N_2378,N_2347);
nor U2447 (N_2447,N_2382,N_2381);
or U2448 (N_2448,N_2376,N_2341);
and U2449 (N_2449,N_2340,N_2382);
nor U2450 (N_2450,N_2391,N_2370);
and U2451 (N_2451,N_2346,N_2347);
or U2452 (N_2452,N_2368,N_2341);
nor U2453 (N_2453,N_2354,N_2364);
or U2454 (N_2454,N_2347,N_2369);
nor U2455 (N_2455,N_2381,N_2395);
nand U2456 (N_2456,N_2379,N_2382);
nand U2457 (N_2457,N_2360,N_2381);
or U2458 (N_2458,N_2397,N_2379);
nor U2459 (N_2459,N_2384,N_2396);
or U2460 (N_2460,N_2416,N_2407);
or U2461 (N_2461,N_2401,N_2409);
nor U2462 (N_2462,N_2434,N_2423);
and U2463 (N_2463,N_2415,N_2436);
nand U2464 (N_2464,N_2458,N_2410);
and U2465 (N_2465,N_2430,N_2448);
nand U2466 (N_2466,N_2452,N_2425);
and U2467 (N_2467,N_2444,N_2412);
nor U2468 (N_2468,N_2441,N_2428);
or U2469 (N_2469,N_2404,N_2414);
nand U2470 (N_2470,N_2455,N_2402);
and U2471 (N_2471,N_2459,N_2403);
nor U2472 (N_2472,N_2438,N_2451);
or U2473 (N_2473,N_2426,N_2446);
nor U2474 (N_2474,N_2429,N_2447);
or U2475 (N_2475,N_2420,N_2453);
and U2476 (N_2476,N_2400,N_2442);
or U2477 (N_2477,N_2418,N_2421);
and U2478 (N_2478,N_2443,N_2454);
nor U2479 (N_2479,N_2449,N_2433);
nor U2480 (N_2480,N_2417,N_2419);
and U2481 (N_2481,N_2408,N_2427);
xnor U2482 (N_2482,N_2450,N_2424);
or U2483 (N_2483,N_2431,N_2440);
and U2484 (N_2484,N_2411,N_2435);
or U2485 (N_2485,N_2457,N_2413);
and U2486 (N_2486,N_2406,N_2405);
nor U2487 (N_2487,N_2422,N_2439);
and U2488 (N_2488,N_2456,N_2437);
nor U2489 (N_2489,N_2432,N_2445);
nand U2490 (N_2490,N_2442,N_2402);
nor U2491 (N_2491,N_2447,N_2407);
nor U2492 (N_2492,N_2427,N_2438);
or U2493 (N_2493,N_2418,N_2431);
nor U2494 (N_2494,N_2454,N_2427);
or U2495 (N_2495,N_2401,N_2443);
nand U2496 (N_2496,N_2410,N_2435);
or U2497 (N_2497,N_2416,N_2420);
nand U2498 (N_2498,N_2427,N_2418);
and U2499 (N_2499,N_2436,N_2425);
or U2500 (N_2500,N_2434,N_2442);
nor U2501 (N_2501,N_2400,N_2453);
nand U2502 (N_2502,N_2422,N_2423);
or U2503 (N_2503,N_2404,N_2400);
and U2504 (N_2504,N_2424,N_2438);
and U2505 (N_2505,N_2440,N_2427);
or U2506 (N_2506,N_2424,N_2419);
nor U2507 (N_2507,N_2431,N_2439);
nor U2508 (N_2508,N_2439,N_2417);
nor U2509 (N_2509,N_2426,N_2435);
or U2510 (N_2510,N_2425,N_2456);
or U2511 (N_2511,N_2419,N_2411);
and U2512 (N_2512,N_2440,N_2426);
nor U2513 (N_2513,N_2402,N_2438);
and U2514 (N_2514,N_2414,N_2416);
or U2515 (N_2515,N_2401,N_2412);
nor U2516 (N_2516,N_2416,N_2404);
or U2517 (N_2517,N_2456,N_2417);
or U2518 (N_2518,N_2437,N_2449);
or U2519 (N_2519,N_2426,N_2431);
nand U2520 (N_2520,N_2493,N_2497);
or U2521 (N_2521,N_2491,N_2475);
nor U2522 (N_2522,N_2509,N_2465);
and U2523 (N_2523,N_2514,N_2473);
nor U2524 (N_2524,N_2495,N_2517);
or U2525 (N_2525,N_2503,N_2488);
and U2526 (N_2526,N_2513,N_2484);
nand U2527 (N_2527,N_2505,N_2501);
and U2528 (N_2528,N_2468,N_2510);
nor U2529 (N_2529,N_2511,N_2472);
nand U2530 (N_2530,N_2481,N_2460);
nand U2531 (N_2531,N_2504,N_2463);
nor U2532 (N_2532,N_2479,N_2518);
or U2533 (N_2533,N_2496,N_2461);
and U2534 (N_2534,N_2487,N_2486);
or U2535 (N_2535,N_2519,N_2482);
and U2536 (N_2536,N_2508,N_2470);
or U2537 (N_2537,N_2477,N_2467);
or U2538 (N_2538,N_2474,N_2490);
nand U2539 (N_2539,N_2469,N_2480);
and U2540 (N_2540,N_2476,N_2464);
or U2541 (N_2541,N_2489,N_2462);
nand U2542 (N_2542,N_2471,N_2498);
nor U2543 (N_2543,N_2494,N_2492);
and U2544 (N_2544,N_2478,N_2485);
nand U2545 (N_2545,N_2515,N_2506);
nand U2546 (N_2546,N_2516,N_2500);
and U2547 (N_2547,N_2502,N_2483);
and U2548 (N_2548,N_2507,N_2512);
nor U2549 (N_2549,N_2466,N_2499);
or U2550 (N_2550,N_2491,N_2515);
nor U2551 (N_2551,N_2469,N_2474);
and U2552 (N_2552,N_2480,N_2518);
nor U2553 (N_2553,N_2462,N_2511);
or U2554 (N_2554,N_2510,N_2499);
nand U2555 (N_2555,N_2500,N_2505);
nor U2556 (N_2556,N_2471,N_2462);
nor U2557 (N_2557,N_2519,N_2476);
nor U2558 (N_2558,N_2501,N_2500);
nand U2559 (N_2559,N_2506,N_2469);
nor U2560 (N_2560,N_2517,N_2507);
nand U2561 (N_2561,N_2499,N_2511);
nor U2562 (N_2562,N_2512,N_2501);
or U2563 (N_2563,N_2460,N_2503);
nor U2564 (N_2564,N_2506,N_2482);
and U2565 (N_2565,N_2477,N_2503);
and U2566 (N_2566,N_2501,N_2479);
or U2567 (N_2567,N_2513,N_2505);
or U2568 (N_2568,N_2499,N_2488);
or U2569 (N_2569,N_2514,N_2482);
nor U2570 (N_2570,N_2514,N_2465);
and U2571 (N_2571,N_2504,N_2508);
nand U2572 (N_2572,N_2509,N_2516);
nor U2573 (N_2573,N_2519,N_2470);
and U2574 (N_2574,N_2508,N_2484);
nor U2575 (N_2575,N_2506,N_2505);
or U2576 (N_2576,N_2474,N_2519);
or U2577 (N_2577,N_2519,N_2477);
nand U2578 (N_2578,N_2467,N_2512);
and U2579 (N_2579,N_2500,N_2519);
xnor U2580 (N_2580,N_2552,N_2538);
and U2581 (N_2581,N_2547,N_2550);
nor U2582 (N_2582,N_2543,N_2546);
nor U2583 (N_2583,N_2534,N_2535);
xor U2584 (N_2584,N_2548,N_2561);
and U2585 (N_2585,N_2523,N_2560);
nor U2586 (N_2586,N_2574,N_2540);
or U2587 (N_2587,N_2568,N_2542);
and U2588 (N_2588,N_2544,N_2576);
and U2589 (N_2589,N_2579,N_2533);
or U2590 (N_2590,N_2539,N_2532);
nor U2591 (N_2591,N_2520,N_2571);
and U2592 (N_2592,N_2551,N_2573);
or U2593 (N_2593,N_2549,N_2555);
nand U2594 (N_2594,N_2570,N_2558);
and U2595 (N_2595,N_2529,N_2572);
nor U2596 (N_2596,N_2556,N_2528);
nand U2597 (N_2597,N_2578,N_2545);
and U2598 (N_2598,N_2566,N_2527);
or U2599 (N_2599,N_2524,N_2531);
or U2600 (N_2600,N_2565,N_2559);
or U2601 (N_2601,N_2541,N_2537);
nand U2602 (N_2602,N_2569,N_2557);
nand U2603 (N_2603,N_2563,N_2525);
nor U2604 (N_2604,N_2553,N_2564);
nand U2605 (N_2605,N_2526,N_2536);
or U2606 (N_2606,N_2530,N_2521);
or U2607 (N_2607,N_2554,N_2575);
nand U2608 (N_2608,N_2577,N_2522);
or U2609 (N_2609,N_2562,N_2567);
nor U2610 (N_2610,N_2522,N_2534);
nand U2611 (N_2611,N_2558,N_2577);
nor U2612 (N_2612,N_2551,N_2522);
and U2613 (N_2613,N_2568,N_2528);
nor U2614 (N_2614,N_2569,N_2552);
nand U2615 (N_2615,N_2554,N_2563);
or U2616 (N_2616,N_2527,N_2532);
xnor U2617 (N_2617,N_2550,N_2548);
and U2618 (N_2618,N_2565,N_2544);
nor U2619 (N_2619,N_2561,N_2541);
nor U2620 (N_2620,N_2541,N_2568);
or U2621 (N_2621,N_2525,N_2544);
nor U2622 (N_2622,N_2549,N_2521);
nor U2623 (N_2623,N_2551,N_2576);
nor U2624 (N_2624,N_2548,N_2538);
or U2625 (N_2625,N_2554,N_2522);
nor U2626 (N_2626,N_2544,N_2527);
nor U2627 (N_2627,N_2575,N_2576);
and U2628 (N_2628,N_2539,N_2550);
or U2629 (N_2629,N_2565,N_2573);
and U2630 (N_2630,N_2524,N_2526);
nor U2631 (N_2631,N_2533,N_2559);
nand U2632 (N_2632,N_2542,N_2545);
or U2633 (N_2633,N_2525,N_2528);
nand U2634 (N_2634,N_2554,N_2577);
nand U2635 (N_2635,N_2556,N_2534);
nor U2636 (N_2636,N_2569,N_2576);
or U2637 (N_2637,N_2537,N_2578);
nand U2638 (N_2638,N_2547,N_2579);
nand U2639 (N_2639,N_2578,N_2551);
xor U2640 (N_2640,N_2606,N_2586);
nor U2641 (N_2641,N_2582,N_2604);
nor U2642 (N_2642,N_2588,N_2614);
nor U2643 (N_2643,N_2584,N_2630);
nand U2644 (N_2644,N_2629,N_2591);
nor U2645 (N_2645,N_2608,N_2627);
and U2646 (N_2646,N_2628,N_2607);
nand U2647 (N_2647,N_2599,N_2621);
and U2648 (N_2648,N_2638,N_2635);
nor U2649 (N_2649,N_2590,N_2592);
nand U2650 (N_2650,N_2633,N_2611);
nor U2651 (N_2651,N_2622,N_2637);
nor U2652 (N_2652,N_2639,N_2589);
or U2653 (N_2653,N_2618,N_2615);
nor U2654 (N_2654,N_2623,N_2602);
nand U2655 (N_2655,N_2612,N_2617);
nand U2656 (N_2656,N_2620,N_2587);
nor U2657 (N_2657,N_2636,N_2624);
nor U2658 (N_2658,N_2595,N_2613);
nand U2659 (N_2659,N_2610,N_2593);
nand U2660 (N_2660,N_2631,N_2603);
nor U2661 (N_2661,N_2616,N_2580);
nor U2662 (N_2662,N_2634,N_2601);
nand U2663 (N_2663,N_2598,N_2583);
nand U2664 (N_2664,N_2596,N_2619);
or U2665 (N_2665,N_2625,N_2600);
or U2666 (N_2666,N_2632,N_2605);
nand U2667 (N_2667,N_2594,N_2609);
nand U2668 (N_2668,N_2597,N_2581);
nand U2669 (N_2669,N_2626,N_2585);
or U2670 (N_2670,N_2630,N_2580);
nand U2671 (N_2671,N_2622,N_2585);
or U2672 (N_2672,N_2604,N_2580);
and U2673 (N_2673,N_2605,N_2639);
nor U2674 (N_2674,N_2624,N_2635);
or U2675 (N_2675,N_2588,N_2628);
nand U2676 (N_2676,N_2631,N_2609);
or U2677 (N_2677,N_2582,N_2623);
nor U2678 (N_2678,N_2583,N_2629);
nand U2679 (N_2679,N_2616,N_2619);
nor U2680 (N_2680,N_2610,N_2604);
nand U2681 (N_2681,N_2602,N_2590);
nor U2682 (N_2682,N_2603,N_2627);
xor U2683 (N_2683,N_2625,N_2595);
and U2684 (N_2684,N_2585,N_2597);
nand U2685 (N_2685,N_2612,N_2633);
and U2686 (N_2686,N_2614,N_2605);
nand U2687 (N_2687,N_2630,N_2632);
and U2688 (N_2688,N_2583,N_2621);
nand U2689 (N_2689,N_2580,N_2615);
nand U2690 (N_2690,N_2625,N_2624);
or U2691 (N_2691,N_2635,N_2617);
and U2692 (N_2692,N_2614,N_2604);
nor U2693 (N_2693,N_2617,N_2632);
nor U2694 (N_2694,N_2602,N_2589);
nor U2695 (N_2695,N_2615,N_2635);
nor U2696 (N_2696,N_2582,N_2611);
nor U2697 (N_2697,N_2589,N_2626);
nor U2698 (N_2698,N_2639,N_2584);
or U2699 (N_2699,N_2595,N_2626);
nand U2700 (N_2700,N_2681,N_2663);
or U2701 (N_2701,N_2680,N_2653);
or U2702 (N_2702,N_2684,N_2686);
nor U2703 (N_2703,N_2692,N_2674);
nor U2704 (N_2704,N_2647,N_2654);
nor U2705 (N_2705,N_2691,N_2696);
nor U2706 (N_2706,N_2651,N_2649);
nor U2707 (N_2707,N_2671,N_2669);
nor U2708 (N_2708,N_2685,N_2656);
nor U2709 (N_2709,N_2645,N_2670);
or U2710 (N_2710,N_2678,N_2679);
nand U2711 (N_2711,N_2640,N_2659);
nor U2712 (N_2712,N_2666,N_2676);
nor U2713 (N_2713,N_2689,N_2695);
nor U2714 (N_2714,N_2662,N_2668);
nand U2715 (N_2715,N_2672,N_2644);
nor U2716 (N_2716,N_2675,N_2665);
nand U2717 (N_2717,N_2655,N_2646);
or U2718 (N_2718,N_2641,N_2657);
and U2719 (N_2719,N_2673,N_2652);
and U2720 (N_2720,N_2694,N_2642);
nand U2721 (N_2721,N_2683,N_2693);
nand U2722 (N_2722,N_2688,N_2660);
nand U2723 (N_2723,N_2699,N_2690);
nor U2724 (N_2724,N_2697,N_2682);
and U2725 (N_2725,N_2658,N_2664);
or U2726 (N_2726,N_2648,N_2677);
nor U2727 (N_2727,N_2698,N_2650);
xor U2728 (N_2728,N_2667,N_2643);
nor U2729 (N_2729,N_2661,N_2687);
nand U2730 (N_2730,N_2643,N_2660);
or U2731 (N_2731,N_2669,N_2664);
and U2732 (N_2732,N_2665,N_2658);
and U2733 (N_2733,N_2675,N_2669);
and U2734 (N_2734,N_2661,N_2663);
nor U2735 (N_2735,N_2696,N_2642);
xnor U2736 (N_2736,N_2683,N_2649);
nand U2737 (N_2737,N_2643,N_2664);
and U2738 (N_2738,N_2652,N_2655);
nor U2739 (N_2739,N_2678,N_2695);
and U2740 (N_2740,N_2648,N_2649);
nand U2741 (N_2741,N_2655,N_2687);
nor U2742 (N_2742,N_2658,N_2648);
and U2743 (N_2743,N_2657,N_2677);
and U2744 (N_2744,N_2682,N_2681);
and U2745 (N_2745,N_2670,N_2695);
nor U2746 (N_2746,N_2693,N_2664);
or U2747 (N_2747,N_2654,N_2649);
nor U2748 (N_2748,N_2640,N_2686);
and U2749 (N_2749,N_2696,N_2665);
nor U2750 (N_2750,N_2692,N_2651);
or U2751 (N_2751,N_2673,N_2666);
xor U2752 (N_2752,N_2650,N_2694);
nand U2753 (N_2753,N_2652,N_2662);
and U2754 (N_2754,N_2686,N_2687);
nand U2755 (N_2755,N_2653,N_2693);
and U2756 (N_2756,N_2657,N_2667);
nand U2757 (N_2757,N_2642,N_2659);
or U2758 (N_2758,N_2667,N_2651);
nand U2759 (N_2759,N_2678,N_2683);
and U2760 (N_2760,N_2726,N_2712);
xor U2761 (N_2761,N_2737,N_2750);
or U2762 (N_2762,N_2704,N_2727);
nor U2763 (N_2763,N_2720,N_2758);
nor U2764 (N_2764,N_2710,N_2746);
nor U2765 (N_2765,N_2738,N_2748);
and U2766 (N_2766,N_2741,N_2753);
and U2767 (N_2767,N_2715,N_2723);
nor U2768 (N_2768,N_2749,N_2754);
and U2769 (N_2769,N_2755,N_2744);
and U2770 (N_2770,N_2732,N_2745);
nand U2771 (N_2771,N_2703,N_2759);
nand U2772 (N_2772,N_2740,N_2743);
or U2773 (N_2773,N_2721,N_2709);
nand U2774 (N_2774,N_2739,N_2756);
and U2775 (N_2775,N_2716,N_2708);
and U2776 (N_2776,N_2714,N_2700);
or U2777 (N_2777,N_2701,N_2729);
and U2778 (N_2778,N_2730,N_2736);
or U2779 (N_2779,N_2719,N_2724);
nand U2780 (N_2780,N_2757,N_2713);
or U2781 (N_2781,N_2742,N_2707);
nor U2782 (N_2782,N_2711,N_2706);
nand U2783 (N_2783,N_2734,N_2717);
and U2784 (N_2784,N_2722,N_2752);
or U2785 (N_2785,N_2728,N_2731);
nand U2786 (N_2786,N_2747,N_2735);
and U2787 (N_2787,N_2751,N_2718);
or U2788 (N_2788,N_2702,N_2733);
and U2789 (N_2789,N_2725,N_2705);
or U2790 (N_2790,N_2717,N_2754);
nand U2791 (N_2791,N_2717,N_2711);
or U2792 (N_2792,N_2705,N_2742);
nor U2793 (N_2793,N_2732,N_2726);
or U2794 (N_2794,N_2736,N_2729);
nor U2795 (N_2795,N_2753,N_2740);
nand U2796 (N_2796,N_2718,N_2721);
or U2797 (N_2797,N_2733,N_2704);
or U2798 (N_2798,N_2727,N_2734);
xnor U2799 (N_2799,N_2726,N_2713);
or U2800 (N_2800,N_2716,N_2711);
or U2801 (N_2801,N_2709,N_2745);
nand U2802 (N_2802,N_2739,N_2726);
nor U2803 (N_2803,N_2758,N_2715);
and U2804 (N_2804,N_2751,N_2747);
or U2805 (N_2805,N_2705,N_2723);
or U2806 (N_2806,N_2728,N_2717);
or U2807 (N_2807,N_2727,N_2726);
or U2808 (N_2808,N_2727,N_2723);
and U2809 (N_2809,N_2752,N_2751);
or U2810 (N_2810,N_2700,N_2755);
or U2811 (N_2811,N_2718,N_2740);
or U2812 (N_2812,N_2739,N_2718);
nand U2813 (N_2813,N_2727,N_2749);
or U2814 (N_2814,N_2719,N_2737);
and U2815 (N_2815,N_2747,N_2728);
nor U2816 (N_2816,N_2757,N_2752);
nor U2817 (N_2817,N_2718,N_2703);
nor U2818 (N_2818,N_2758,N_2750);
or U2819 (N_2819,N_2725,N_2749);
nor U2820 (N_2820,N_2815,N_2780);
nor U2821 (N_2821,N_2779,N_2785);
and U2822 (N_2822,N_2802,N_2818);
or U2823 (N_2823,N_2761,N_2816);
or U2824 (N_2824,N_2799,N_2792);
nor U2825 (N_2825,N_2776,N_2817);
or U2826 (N_2826,N_2782,N_2764);
or U2827 (N_2827,N_2784,N_2768);
nor U2828 (N_2828,N_2805,N_2806);
nor U2829 (N_2829,N_2781,N_2774);
nand U2830 (N_2830,N_2787,N_2803);
and U2831 (N_2831,N_2814,N_2765);
nor U2832 (N_2832,N_2794,N_2793);
nand U2833 (N_2833,N_2771,N_2807);
or U2834 (N_2834,N_2813,N_2801);
and U2835 (N_2835,N_2796,N_2783);
and U2836 (N_2836,N_2808,N_2791);
and U2837 (N_2837,N_2795,N_2790);
nor U2838 (N_2838,N_2769,N_2810);
and U2839 (N_2839,N_2778,N_2819);
or U2840 (N_2840,N_2777,N_2773);
or U2841 (N_2841,N_2788,N_2762);
nand U2842 (N_2842,N_2789,N_2770);
nand U2843 (N_2843,N_2775,N_2800);
or U2844 (N_2844,N_2811,N_2767);
nor U2845 (N_2845,N_2812,N_2786);
nor U2846 (N_2846,N_2772,N_2763);
xor U2847 (N_2847,N_2797,N_2760);
and U2848 (N_2848,N_2804,N_2798);
or U2849 (N_2849,N_2809,N_2766);
and U2850 (N_2850,N_2770,N_2783);
nor U2851 (N_2851,N_2798,N_2787);
xnor U2852 (N_2852,N_2777,N_2788);
and U2853 (N_2853,N_2774,N_2767);
nor U2854 (N_2854,N_2794,N_2765);
or U2855 (N_2855,N_2799,N_2805);
nor U2856 (N_2856,N_2801,N_2788);
nor U2857 (N_2857,N_2817,N_2819);
or U2858 (N_2858,N_2763,N_2802);
or U2859 (N_2859,N_2801,N_2784);
or U2860 (N_2860,N_2772,N_2777);
xnor U2861 (N_2861,N_2791,N_2805);
or U2862 (N_2862,N_2803,N_2805);
nand U2863 (N_2863,N_2784,N_2783);
or U2864 (N_2864,N_2810,N_2811);
or U2865 (N_2865,N_2780,N_2792);
nand U2866 (N_2866,N_2772,N_2765);
nand U2867 (N_2867,N_2775,N_2767);
and U2868 (N_2868,N_2790,N_2770);
and U2869 (N_2869,N_2781,N_2797);
nor U2870 (N_2870,N_2808,N_2811);
nand U2871 (N_2871,N_2799,N_2762);
and U2872 (N_2872,N_2818,N_2781);
nor U2873 (N_2873,N_2777,N_2796);
nor U2874 (N_2874,N_2804,N_2782);
nor U2875 (N_2875,N_2781,N_2788);
nor U2876 (N_2876,N_2763,N_2804);
or U2877 (N_2877,N_2816,N_2818);
and U2878 (N_2878,N_2787,N_2813);
and U2879 (N_2879,N_2805,N_2781);
nand U2880 (N_2880,N_2853,N_2828);
nand U2881 (N_2881,N_2825,N_2871);
or U2882 (N_2882,N_2852,N_2870);
or U2883 (N_2883,N_2868,N_2831);
nor U2884 (N_2884,N_2849,N_2839);
nand U2885 (N_2885,N_2840,N_2843);
nor U2886 (N_2886,N_2848,N_2838);
and U2887 (N_2887,N_2846,N_2877);
nand U2888 (N_2888,N_2830,N_2872);
or U2889 (N_2889,N_2858,N_2821);
and U2890 (N_2890,N_2820,N_2842);
nand U2891 (N_2891,N_2855,N_2867);
or U2892 (N_2892,N_2835,N_2860);
and U2893 (N_2893,N_2844,N_2841);
nand U2894 (N_2894,N_2833,N_2869);
and U2895 (N_2895,N_2854,N_2879);
or U2896 (N_2896,N_2823,N_2878);
or U2897 (N_2897,N_2856,N_2826);
or U2898 (N_2898,N_2864,N_2857);
and U2899 (N_2899,N_2874,N_2832);
nor U2900 (N_2900,N_2861,N_2847);
nor U2901 (N_2901,N_2859,N_2827);
or U2902 (N_2902,N_2837,N_2836);
or U2903 (N_2903,N_2822,N_2873);
or U2904 (N_2904,N_2865,N_2834);
or U2905 (N_2905,N_2866,N_2845);
nand U2906 (N_2906,N_2862,N_2824);
or U2907 (N_2907,N_2875,N_2850);
nor U2908 (N_2908,N_2851,N_2876);
xnor U2909 (N_2909,N_2829,N_2863);
and U2910 (N_2910,N_2861,N_2877);
or U2911 (N_2911,N_2828,N_2876);
nand U2912 (N_2912,N_2875,N_2874);
or U2913 (N_2913,N_2871,N_2863);
and U2914 (N_2914,N_2859,N_2861);
and U2915 (N_2915,N_2865,N_2859);
or U2916 (N_2916,N_2876,N_2845);
and U2917 (N_2917,N_2835,N_2870);
or U2918 (N_2918,N_2848,N_2851);
or U2919 (N_2919,N_2821,N_2856);
or U2920 (N_2920,N_2873,N_2820);
and U2921 (N_2921,N_2833,N_2844);
and U2922 (N_2922,N_2864,N_2874);
or U2923 (N_2923,N_2830,N_2849);
or U2924 (N_2924,N_2838,N_2874);
and U2925 (N_2925,N_2840,N_2823);
or U2926 (N_2926,N_2820,N_2851);
nor U2927 (N_2927,N_2821,N_2849);
nor U2928 (N_2928,N_2857,N_2854);
and U2929 (N_2929,N_2822,N_2869);
nand U2930 (N_2930,N_2821,N_2865);
and U2931 (N_2931,N_2872,N_2877);
or U2932 (N_2932,N_2855,N_2849);
and U2933 (N_2933,N_2849,N_2853);
nor U2934 (N_2934,N_2858,N_2830);
xnor U2935 (N_2935,N_2876,N_2824);
or U2936 (N_2936,N_2840,N_2866);
and U2937 (N_2937,N_2824,N_2828);
or U2938 (N_2938,N_2831,N_2872);
nand U2939 (N_2939,N_2827,N_2831);
or U2940 (N_2940,N_2887,N_2898);
nand U2941 (N_2941,N_2889,N_2905);
nand U2942 (N_2942,N_2920,N_2934);
or U2943 (N_2943,N_2918,N_2882);
nor U2944 (N_2944,N_2910,N_2911);
nand U2945 (N_2945,N_2886,N_2915);
nand U2946 (N_2946,N_2880,N_2881);
nand U2947 (N_2947,N_2925,N_2913);
nand U2948 (N_2948,N_2909,N_2931);
or U2949 (N_2949,N_2899,N_2895);
or U2950 (N_2950,N_2906,N_2885);
nor U2951 (N_2951,N_2908,N_2939);
nand U2952 (N_2952,N_2907,N_2903);
nand U2953 (N_2953,N_2935,N_2916);
nand U2954 (N_2954,N_2891,N_2921);
nand U2955 (N_2955,N_2897,N_2933);
and U2956 (N_2956,N_2892,N_2904);
and U2957 (N_2957,N_2923,N_2936);
or U2958 (N_2958,N_2926,N_2930);
or U2959 (N_2959,N_2929,N_2893);
xnor U2960 (N_2960,N_2922,N_2884);
and U2961 (N_2961,N_2928,N_2888);
nand U2962 (N_2962,N_2912,N_2894);
nand U2963 (N_2963,N_2919,N_2938);
and U2964 (N_2964,N_2900,N_2902);
or U2965 (N_2965,N_2896,N_2883);
nor U2966 (N_2966,N_2914,N_2890);
nand U2967 (N_2967,N_2937,N_2927);
or U2968 (N_2968,N_2924,N_2932);
nand U2969 (N_2969,N_2901,N_2917);
nor U2970 (N_2970,N_2909,N_2893);
and U2971 (N_2971,N_2920,N_2887);
nand U2972 (N_2972,N_2900,N_2929);
or U2973 (N_2973,N_2889,N_2935);
or U2974 (N_2974,N_2880,N_2895);
nor U2975 (N_2975,N_2901,N_2888);
or U2976 (N_2976,N_2896,N_2887);
and U2977 (N_2977,N_2920,N_2882);
and U2978 (N_2978,N_2884,N_2904);
nor U2979 (N_2979,N_2932,N_2933);
nor U2980 (N_2980,N_2915,N_2927);
and U2981 (N_2981,N_2911,N_2893);
and U2982 (N_2982,N_2930,N_2903);
and U2983 (N_2983,N_2885,N_2907);
nand U2984 (N_2984,N_2917,N_2928);
or U2985 (N_2985,N_2926,N_2933);
nand U2986 (N_2986,N_2924,N_2914);
and U2987 (N_2987,N_2882,N_2905);
or U2988 (N_2988,N_2935,N_2888);
nand U2989 (N_2989,N_2883,N_2937);
xnor U2990 (N_2990,N_2937,N_2915);
nand U2991 (N_2991,N_2890,N_2897);
and U2992 (N_2992,N_2939,N_2931);
and U2993 (N_2993,N_2893,N_2916);
or U2994 (N_2994,N_2899,N_2911);
or U2995 (N_2995,N_2908,N_2892);
nand U2996 (N_2996,N_2916,N_2904);
or U2997 (N_2997,N_2881,N_2906);
xor U2998 (N_2998,N_2909,N_2895);
or U2999 (N_2999,N_2930,N_2931);
nand UO_0 (O_0,N_2962,N_2963);
xor UO_1 (O_1,N_2997,N_2947);
nand UO_2 (O_2,N_2984,N_2978);
nor UO_3 (O_3,N_2987,N_2969);
nor UO_4 (O_4,N_2956,N_2966);
nor UO_5 (O_5,N_2976,N_2958);
nor UO_6 (O_6,N_2943,N_2975);
nand UO_7 (O_7,N_2946,N_2942);
nand UO_8 (O_8,N_2979,N_2993);
and UO_9 (O_9,N_2988,N_2971);
or UO_10 (O_10,N_2985,N_2989);
or UO_11 (O_11,N_2990,N_2998);
nand UO_12 (O_12,N_2948,N_2957);
or UO_13 (O_13,N_2961,N_2944);
nor UO_14 (O_14,N_2945,N_2982);
nand UO_15 (O_15,N_2953,N_2968);
nor UO_16 (O_16,N_2967,N_2991);
and UO_17 (O_17,N_2970,N_2959);
nand UO_18 (O_18,N_2983,N_2972);
and UO_19 (O_19,N_2980,N_2986);
nand UO_20 (O_20,N_2949,N_2952);
or UO_21 (O_21,N_2994,N_2940);
nand UO_22 (O_22,N_2951,N_2999);
nor UO_23 (O_23,N_2950,N_2973);
nand UO_24 (O_24,N_2995,N_2941);
nor UO_25 (O_25,N_2981,N_2954);
or UO_26 (O_26,N_2964,N_2977);
nand UO_27 (O_27,N_2965,N_2992);
nor UO_28 (O_28,N_2974,N_2960);
xor UO_29 (O_29,N_2996,N_2955);
nor UO_30 (O_30,N_2947,N_2962);
nor UO_31 (O_31,N_2983,N_2943);
nor UO_32 (O_32,N_2993,N_2982);
nand UO_33 (O_33,N_2974,N_2981);
and UO_34 (O_34,N_2986,N_2948);
nand UO_35 (O_35,N_2992,N_2962);
nand UO_36 (O_36,N_2971,N_2960);
nor UO_37 (O_37,N_2997,N_2999);
xnor UO_38 (O_38,N_2952,N_2974);
or UO_39 (O_39,N_2977,N_2960);
and UO_40 (O_40,N_2985,N_2963);
nand UO_41 (O_41,N_2951,N_2985);
nand UO_42 (O_42,N_2963,N_2953);
nor UO_43 (O_43,N_2947,N_2948);
and UO_44 (O_44,N_2944,N_2977);
nor UO_45 (O_45,N_2987,N_2946);
or UO_46 (O_46,N_2957,N_2979);
or UO_47 (O_47,N_2988,N_2942);
nor UO_48 (O_48,N_2966,N_2990);
nor UO_49 (O_49,N_2963,N_2997);
nor UO_50 (O_50,N_2997,N_2979);
nand UO_51 (O_51,N_2961,N_2996);
or UO_52 (O_52,N_2988,N_2947);
nor UO_53 (O_53,N_2978,N_2995);
and UO_54 (O_54,N_2994,N_2973);
nand UO_55 (O_55,N_2964,N_2955);
or UO_56 (O_56,N_2988,N_2983);
and UO_57 (O_57,N_2969,N_2976);
xor UO_58 (O_58,N_2971,N_2955);
and UO_59 (O_59,N_2954,N_2994);
or UO_60 (O_60,N_2991,N_2971);
nor UO_61 (O_61,N_2972,N_2952);
nand UO_62 (O_62,N_2950,N_2975);
or UO_63 (O_63,N_2960,N_2997);
or UO_64 (O_64,N_2970,N_2993);
nor UO_65 (O_65,N_2955,N_2944);
nor UO_66 (O_66,N_2997,N_2953);
or UO_67 (O_67,N_2947,N_2977);
and UO_68 (O_68,N_2946,N_2992);
nor UO_69 (O_69,N_2977,N_2941);
xor UO_70 (O_70,N_2974,N_2945);
nand UO_71 (O_71,N_2989,N_2992);
nor UO_72 (O_72,N_2969,N_2999);
nand UO_73 (O_73,N_2942,N_2993);
and UO_74 (O_74,N_2943,N_2966);
nand UO_75 (O_75,N_2947,N_2995);
or UO_76 (O_76,N_2987,N_2996);
nand UO_77 (O_77,N_2996,N_2986);
and UO_78 (O_78,N_2951,N_2995);
nand UO_79 (O_79,N_2941,N_2998);
or UO_80 (O_80,N_2984,N_2971);
and UO_81 (O_81,N_2999,N_2940);
nor UO_82 (O_82,N_2996,N_2953);
nand UO_83 (O_83,N_2974,N_2991);
nor UO_84 (O_84,N_2951,N_2943);
or UO_85 (O_85,N_2983,N_2950);
nor UO_86 (O_86,N_2999,N_2970);
nor UO_87 (O_87,N_2977,N_2945);
nand UO_88 (O_88,N_2978,N_2983);
or UO_89 (O_89,N_2959,N_2991);
or UO_90 (O_90,N_2975,N_2967);
or UO_91 (O_91,N_2997,N_2978);
nor UO_92 (O_92,N_2988,N_2986);
and UO_93 (O_93,N_2978,N_2945);
and UO_94 (O_94,N_2981,N_2957);
or UO_95 (O_95,N_2946,N_2970);
xnor UO_96 (O_96,N_2941,N_2951);
and UO_97 (O_97,N_2971,N_2956);
nand UO_98 (O_98,N_2969,N_2958);
nand UO_99 (O_99,N_2999,N_2947);
nand UO_100 (O_100,N_2977,N_2955);
nand UO_101 (O_101,N_2999,N_2961);
or UO_102 (O_102,N_2968,N_2948);
xor UO_103 (O_103,N_2949,N_2950);
nand UO_104 (O_104,N_2988,N_2985);
or UO_105 (O_105,N_2981,N_2958);
nand UO_106 (O_106,N_2987,N_2992);
or UO_107 (O_107,N_2946,N_2957);
nand UO_108 (O_108,N_2996,N_2995);
nand UO_109 (O_109,N_2977,N_2987);
or UO_110 (O_110,N_2974,N_2977);
nor UO_111 (O_111,N_2998,N_2985);
nand UO_112 (O_112,N_2940,N_2981);
and UO_113 (O_113,N_2972,N_2967);
nand UO_114 (O_114,N_2957,N_2964);
nor UO_115 (O_115,N_2951,N_2961);
nand UO_116 (O_116,N_2983,N_2960);
and UO_117 (O_117,N_2985,N_2984);
nand UO_118 (O_118,N_2954,N_2948);
nand UO_119 (O_119,N_2998,N_2944);
nand UO_120 (O_120,N_2944,N_2989);
nand UO_121 (O_121,N_2953,N_2954);
or UO_122 (O_122,N_2989,N_2959);
nand UO_123 (O_123,N_2996,N_2990);
or UO_124 (O_124,N_2992,N_2967);
nand UO_125 (O_125,N_2943,N_2970);
nand UO_126 (O_126,N_2957,N_2980);
nand UO_127 (O_127,N_2984,N_2941);
nor UO_128 (O_128,N_2981,N_2945);
nand UO_129 (O_129,N_2985,N_2954);
and UO_130 (O_130,N_2976,N_2950);
and UO_131 (O_131,N_2944,N_2973);
xor UO_132 (O_132,N_2964,N_2987);
and UO_133 (O_133,N_2991,N_2966);
nor UO_134 (O_134,N_2959,N_2956);
or UO_135 (O_135,N_2956,N_2945);
and UO_136 (O_136,N_2952,N_2975);
nand UO_137 (O_137,N_2940,N_2948);
nor UO_138 (O_138,N_2946,N_2964);
nor UO_139 (O_139,N_2950,N_2957);
or UO_140 (O_140,N_2952,N_2958);
nor UO_141 (O_141,N_2985,N_2943);
and UO_142 (O_142,N_2985,N_2959);
nand UO_143 (O_143,N_2968,N_2942);
nand UO_144 (O_144,N_2984,N_2952);
nor UO_145 (O_145,N_2993,N_2986);
and UO_146 (O_146,N_2966,N_2953);
or UO_147 (O_147,N_2957,N_2978);
or UO_148 (O_148,N_2949,N_2974);
nor UO_149 (O_149,N_2958,N_2961);
or UO_150 (O_150,N_2957,N_2960);
nand UO_151 (O_151,N_2942,N_2960);
nor UO_152 (O_152,N_2999,N_2946);
nand UO_153 (O_153,N_2999,N_2956);
xor UO_154 (O_154,N_2983,N_2941);
nor UO_155 (O_155,N_2972,N_2949);
or UO_156 (O_156,N_2951,N_2980);
nand UO_157 (O_157,N_2975,N_2968);
nor UO_158 (O_158,N_2988,N_2976);
nand UO_159 (O_159,N_2942,N_2955);
nand UO_160 (O_160,N_2991,N_2949);
and UO_161 (O_161,N_2962,N_2949);
nor UO_162 (O_162,N_2978,N_2970);
or UO_163 (O_163,N_2948,N_2994);
nand UO_164 (O_164,N_2983,N_2973);
nand UO_165 (O_165,N_2976,N_2996);
and UO_166 (O_166,N_2961,N_2962);
or UO_167 (O_167,N_2942,N_2961);
nor UO_168 (O_168,N_2959,N_2984);
nor UO_169 (O_169,N_2959,N_2975);
nor UO_170 (O_170,N_2987,N_2968);
nor UO_171 (O_171,N_2946,N_2983);
and UO_172 (O_172,N_2983,N_2959);
nor UO_173 (O_173,N_2990,N_2989);
nor UO_174 (O_174,N_2974,N_2978);
nor UO_175 (O_175,N_2952,N_2964);
or UO_176 (O_176,N_2947,N_2958);
nand UO_177 (O_177,N_2988,N_2964);
nand UO_178 (O_178,N_2959,N_2980);
nor UO_179 (O_179,N_2979,N_2973);
nor UO_180 (O_180,N_2955,N_2992);
xor UO_181 (O_181,N_2965,N_2986);
and UO_182 (O_182,N_2989,N_2953);
or UO_183 (O_183,N_2962,N_2946);
nand UO_184 (O_184,N_2957,N_2973);
nand UO_185 (O_185,N_2988,N_2966);
nand UO_186 (O_186,N_2944,N_2978);
and UO_187 (O_187,N_2995,N_2962);
nand UO_188 (O_188,N_2971,N_2957);
and UO_189 (O_189,N_2957,N_2943);
nand UO_190 (O_190,N_2989,N_2982);
or UO_191 (O_191,N_2987,N_2950);
nor UO_192 (O_192,N_2959,N_2945);
and UO_193 (O_193,N_2942,N_2997);
nand UO_194 (O_194,N_2944,N_2974);
or UO_195 (O_195,N_2963,N_2970);
nor UO_196 (O_196,N_2983,N_2981);
nor UO_197 (O_197,N_2982,N_2962);
nand UO_198 (O_198,N_2947,N_2985);
or UO_199 (O_199,N_2968,N_2969);
nor UO_200 (O_200,N_2994,N_2987);
or UO_201 (O_201,N_2967,N_2961);
nor UO_202 (O_202,N_2986,N_2971);
and UO_203 (O_203,N_2974,N_2995);
nor UO_204 (O_204,N_2969,N_2942);
or UO_205 (O_205,N_2999,N_2996);
and UO_206 (O_206,N_2982,N_2959);
nand UO_207 (O_207,N_2964,N_2990);
or UO_208 (O_208,N_2970,N_2940);
xor UO_209 (O_209,N_2952,N_2979);
nand UO_210 (O_210,N_2965,N_2954);
nor UO_211 (O_211,N_2968,N_2960);
or UO_212 (O_212,N_2960,N_2943);
and UO_213 (O_213,N_2981,N_2943);
or UO_214 (O_214,N_2965,N_2990);
nand UO_215 (O_215,N_2953,N_2983);
nor UO_216 (O_216,N_2985,N_2961);
or UO_217 (O_217,N_2959,N_2968);
nor UO_218 (O_218,N_2969,N_2996);
and UO_219 (O_219,N_2983,N_2944);
nand UO_220 (O_220,N_2996,N_2950);
and UO_221 (O_221,N_2946,N_2945);
nor UO_222 (O_222,N_2965,N_2958);
nand UO_223 (O_223,N_2968,N_2947);
or UO_224 (O_224,N_2994,N_2972);
nand UO_225 (O_225,N_2944,N_2981);
xnor UO_226 (O_226,N_2971,N_2941);
nand UO_227 (O_227,N_2974,N_2958);
and UO_228 (O_228,N_2968,N_2951);
and UO_229 (O_229,N_2952,N_2976);
nor UO_230 (O_230,N_2992,N_2970);
nor UO_231 (O_231,N_2965,N_2978);
nor UO_232 (O_232,N_2998,N_2976);
and UO_233 (O_233,N_2955,N_2993);
or UO_234 (O_234,N_2972,N_2974);
nor UO_235 (O_235,N_2978,N_2940);
or UO_236 (O_236,N_2978,N_2952);
nor UO_237 (O_237,N_2974,N_2982);
nand UO_238 (O_238,N_2982,N_2998);
nand UO_239 (O_239,N_2980,N_2979);
and UO_240 (O_240,N_2971,N_2990);
and UO_241 (O_241,N_2974,N_2954);
or UO_242 (O_242,N_2989,N_2943);
nor UO_243 (O_243,N_2992,N_2999);
nor UO_244 (O_244,N_2995,N_2950);
nor UO_245 (O_245,N_2951,N_2990);
nand UO_246 (O_246,N_2941,N_2981);
or UO_247 (O_247,N_2954,N_2959);
or UO_248 (O_248,N_2994,N_2985);
nor UO_249 (O_249,N_2987,N_2999);
and UO_250 (O_250,N_2948,N_2952);
nand UO_251 (O_251,N_2983,N_2967);
and UO_252 (O_252,N_2988,N_2959);
nand UO_253 (O_253,N_2951,N_2986);
nor UO_254 (O_254,N_2989,N_2984);
and UO_255 (O_255,N_2940,N_2990);
nand UO_256 (O_256,N_2967,N_2956);
and UO_257 (O_257,N_2977,N_2995);
and UO_258 (O_258,N_2957,N_2940);
nor UO_259 (O_259,N_2987,N_2960);
or UO_260 (O_260,N_2980,N_2966);
nand UO_261 (O_261,N_2985,N_2981);
nor UO_262 (O_262,N_2945,N_2997);
and UO_263 (O_263,N_2990,N_2995);
or UO_264 (O_264,N_2968,N_2940);
xor UO_265 (O_265,N_2982,N_2951);
nor UO_266 (O_266,N_2971,N_2989);
and UO_267 (O_267,N_2940,N_2977);
nand UO_268 (O_268,N_2941,N_2992);
nor UO_269 (O_269,N_2947,N_2969);
or UO_270 (O_270,N_2985,N_2990);
and UO_271 (O_271,N_2980,N_2942);
and UO_272 (O_272,N_2991,N_2947);
or UO_273 (O_273,N_2941,N_2950);
nand UO_274 (O_274,N_2953,N_2975);
or UO_275 (O_275,N_2989,N_2949);
and UO_276 (O_276,N_2946,N_2944);
or UO_277 (O_277,N_2958,N_2946);
or UO_278 (O_278,N_2995,N_2987);
and UO_279 (O_279,N_2991,N_2961);
nor UO_280 (O_280,N_2960,N_2992);
nor UO_281 (O_281,N_2971,N_2958);
and UO_282 (O_282,N_2966,N_2946);
and UO_283 (O_283,N_2986,N_2981);
nand UO_284 (O_284,N_2982,N_2970);
xnor UO_285 (O_285,N_2953,N_2992);
nor UO_286 (O_286,N_2943,N_2987);
or UO_287 (O_287,N_2993,N_2990);
nor UO_288 (O_288,N_2980,N_2963);
nand UO_289 (O_289,N_2980,N_2972);
nand UO_290 (O_290,N_2985,N_2957);
nand UO_291 (O_291,N_2953,N_2952);
and UO_292 (O_292,N_2969,N_2977);
or UO_293 (O_293,N_2992,N_2957);
or UO_294 (O_294,N_2956,N_2983);
nand UO_295 (O_295,N_2998,N_2977);
and UO_296 (O_296,N_2963,N_2968);
or UO_297 (O_297,N_2963,N_2949);
nor UO_298 (O_298,N_2983,N_2979);
nor UO_299 (O_299,N_2977,N_2981);
and UO_300 (O_300,N_2979,N_2984);
or UO_301 (O_301,N_2993,N_2964);
nand UO_302 (O_302,N_2975,N_2976);
and UO_303 (O_303,N_2957,N_2965);
or UO_304 (O_304,N_2985,N_2958);
or UO_305 (O_305,N_2968,N_2950);
nand UO_306 (O_306,N_2969,N_2974);
or UO_307 (O_307,N_2958,N_2948);
or UO_308 (O_308,N_2955,N_2946);
and UO_309 (O_309,N_2940,N_2984);
and UO_310 (O_310,N_2981,N_2987);
and UO_311 (O_311,N_2948,N_2951);
and UO_312 (O_312,N_2993,N_2972);
nor UO_313 (O_313,N_2986,N_2973);
nand UO_314 (O_314,N_2956,N_2957);
nand UO_315 (O_315,N_2967,N_2946);
or UO_316 (O_316,N_2954,N_2957);
or UO_317 (O_317,N_2949,N_2992);
nand UO_318 (O_318,N_2943,N_2947);
or UO_319 (O_319,N_2964,N_2962);
nor UO_320 (O_320,N_2944,N_2966);
nor UO_321 (O_321,N_2940,N_2950);
nand UO_322 (O_322,N_2979,N_2995);
or UO_323 (O_323,N_2986,N_2955);
or UO_324 (O_324,N_2950,N_2967);
or UO_325 (O_325,N_2981,N_2956);
or UO_326 (O_326,N_2959,N_2953);
or UO_327 (O_327,N_2973,N_2984);
and UO_328 (O_328,N_2987,N_2955);
or UO_329 (O_329,N_2973,N_2996);
nor UO_330 (O_330,N_2941,N_2969);
nand UO_331 (O_331,N_2999,N_2949);
or UO_332 (O_332,N_2948,N_2993);
nor UO_333 (O_333,N_2950,N_2992);
or UO_334 (O_334,N_2982,N_2960);
nor UO_335 (O_335,N_2954,N_2992);
nor UO_336 (O_336,N_2958,N_2989);
or UO_337 (O_337,N_2986,N_2997);
or UO_338 (O_338,N_2949,N_2978);
or UO_339 (O_339,N_2984,N_2967);
and UO_340 (O_340,N_2950,N_2956);
and UO_341 (O_341,N_2971,N_2961);
nor UO_342 (O_342,N_2966,N_2967);
nor UO_343 (O_343,N_2952,N_2981);
nand UO_344 (O_344,N_2986,N_2959);
nor UO_345 (O_345,N_2990,N_2956);
nor UO_346 (O_346,N_2979,N_2956);
and UO_347 (O_347,N_2956,N_2996);
or UO_348 (O_348,N_2978,N_2972);
or UO_349 (O_349,N_2986,N_2972);
or UO_350 (O_350,N_2978,N_2973);
nand UO_351 (O_351,N_2965,N_2972);
or UO_352 (O_352,N_2954,N_2983);
xor UO_353 (O_353,N_2941,N_2957);
nor UO_354 (O_354,N_2953,N_2964);
nor UO_355 (O_355,N_2942,N_2956);
nand UO_356 (O_356,N_2999,N_2990);
nand UO_357 (O_357,N_2966,N_2970);
nand UO_358 (O_358,N_2994,N_2964);
nand UO_359 (O_359,N_2961,N_2970);
nand UO_360 (O_360,N_2954,N_2963);
and UO_361 (O_361,N_2985,N_2969);
or UO_362 (O_362,N_2997,N_2944);
nand UO_363 (O_363,N_2974,N_2959);
nand UO_364 (O_364,N_2979,N_2981);
nand UO_365 (O_365,N_2958,N_2951);
nor UO_366 (O_366,N_2984,N_2954);
nor UO_367 (O_367,N_2998,N_2992);
and UO_368 (O_368,N_2962,N_2980);
or UO_369 (O_369,N_2969,N_2984);
nor UO_370 (O_370,N_2970,N_2958);
or UO_371 (O_371,N_2969,N_2991);
and UO_372 (O_372,N_2989,N_2942);
nand UO_373 (O_373,N_2957,N_2951);
nor UO_374 (O_374,N_2996,N_2962);
nand UO_375 (O_375,N_2965,N_2980);
and UO_376 (O_376,N_2967,N_2968);
or UO_377 (O_377,N_2958,N_2968);
and UO_378 (O_378,N_2945,N_2996);
and UO_379 (O_379,N_2964,N_2942);
nor UO_380 (O_380,N_2953,N_2976);
nand UO_381 (O_381,N_2985,N_2960);
or UO_382 (O_382,N_2990,N_2973);
and UO_383 (O_383,N_2944,N_2980);
nand UO_384 (O_384,N_2984,N_2949);
nor UO_385 (O_385,N_2960,N_2954);
nor UO_386 (O_386,N_2947,N_2975);
nand UO_387 (O_387,N_2944,N_2950);
nand UO_388 (O_388,N_2990,N_2972);
nand UO_389 (O_389,N_2951,N_2964);
nor UO_390 (O_390,N_2956,N_2976);
nor UO_391 (O_391,N_2991,N_2950);
nor UO_392 (O_392,N_2944,N_2984);
and UO_393 (O_393,N_2942,N_2972);
nor UO_394 (O_394,N_2942,N_2967);
nor UO_395 (O_395,N_2958,N_2990);
and UO_396 (O_396,N_2942,N_2971);
nor UO_397 (O_397,N_2945,N_2987);
and UO_398 (O_398,N_2948,N_2941);
or UO_399 (O_399,N_2952,N_2973);
or UO_400 (O_400,N_2972,N_2992);
and UO_401 (O_401,N_2963,N_2978);
or UO_402 (O_402,N_2980,N_2945);
nand UO_403 (O_403,N_2969,N_2951);
or UO_404 (O_404,N_2982,N_2966);
xor UO_405 (O_405,N_2962,N_2940);
nand UO_406 (O_406,N_2947,N_2946);
nand UO_407 (O_407,N_2965,N_2942);
and UO_408 (O_408,N_2989,N_2964);
xnor UO_409 (O_409,N_2980,N_2997);
and UO_410 (O_410,N_2977,N_2991);
nor UO_411 (O_411,N_2961,N_2963);
nor UO_412 (O_412,N_2981,N_2976);
nand UO_413 (O_413,N_2963,N_2956);
nand UO_414 (O_414,N_2966,N_2983);
xnor UO_415 (O_415,N_2976,N_2949);
nor UO_416 (O_416,N_2948,N_2955);
nor UO_417 (O_417,N_2987,N_2978);
or UO_418 (O_418,N_2961,N_2940);
xnor UO_419 (O_419,N_2945,N_2961);
nand UO_420 (O_420,N_2989,N_2951);
or UO_421 (O_421,N_2950,N_2985);
nor UO_422 (O_422,N_2967,N_2987);
and UO_423 (O_423,N_2971,N_2980);
nor UO_424 (O_424,N_2952,N_2947);
and UO_425 (O_425,N_2950,N_2970);
nand UO_426 (O_426,N_2999,N_2953);
nor UO_427 (O_427,N_2947,N_2978);
nor UO_428 (O_428,N_2967,N_2960);
nand UO_429 (O_429,N_2991,N_2993);
or UO_430 (O_430,N_2994,N_2967);
nor UO_431 (O_431,N_2942,N_2953);
nand UO_432 (O_432,N_2988,N_2984);
nand UO_433 (O_433,N_2956,N_2962);
or UO_434 (O_434,N_2942,N_2958);
nand UO_435 (O_435,N_2971,N_2951);
nand UO_436 (O_436,N_2940,N_2973);
and UO_437 (O_437,N_2993,N_2980);
nor UO_438 (O_438,N_2942,N_2940);
nor UO_439 (O_439,N_2956,N_2998);
and UO_440 (O_440,N_2983,N_2985);
nor UO_441 (O_441,N_2941,N_2979);
and UO_442 (O_442,N_2949,N_2965);
and UO_443 (O_443,N_2976,N_2957);
and UO_444 (O_444,N_2943,N_2946);
and UO_445 (O_445,N_2947,N_2971);
nor UO_446 (O_446,N_2998,N_2972);
and UO_447 (O_447,N_2954,N_2956);
or UO_448 (O_448,N_2988,N_2951);
nand UO_449 (O_449,N_2954,N_2975);
nand UO_450 (O_450,N_2940,N_2972);
nor UO_451 (O_451,N_2986,N_2974);
and UO_452 (O_452,N_2965,N_2946);
or UO_453 (O_453,N_2981,N_2965);
nor UO_454 (O_454,N_2994,N_2952);
or UO_455 (O_455,N_2961,N_2997);
or UO_456 (O_456,N_2946,N_2976);
and UO_457 (O_457,N_2966,N_2978);
and UO_458 (O_458,N_2987,N_2973);
nand UO_459 (O_459,N_2955,N_2994);
nand UO_460 (O_460,N_2943,N_2996);
nor UO_461 (O_461,N_2973,N_2999);
nand UO_462 (O_462,N_2985,N_2964);
or UO_463 (O_463,N_2982,N_2954);
or UO_464 (O_464,N_2990,N_2980);
nor UO_465 (O_465,N_2983,N_2997);
and UO_466 (O_466,N_2991,N_2958);
nand UO_467 (O_467,N_2982,N_2975);
nor UO_468 (O_468,N_2963,N_2984);
nand UO_469 (O_469,N_2983,N_2947);
nand UO_470 (O_470,N_2940,N_2949);
nor UO_471 (O_471,N_2995,N_2966);
nor UO_472 (O_472,N_2949,N_2994);
nand UO_473 (O_473,N_2991,N_2973);
nand UO_474 (O_474,N_2951,N_2944);
nand UO_475 (O_475,N_2967,N_2948);
or UO_476 (O_476,N_2992,N_2943);
or UO_477 (O_477,N_2942,N_2950);
or UO_478 (O_478,N_2980,N_2983);
or UO_479 (O_479,N_2954,N_2943);
or UO_480 (O_480,N_2975,N_2951);
nor UO_481 (O_481,N_2940,N_2964);
nor UO_482 (O_482,N_2974,N_2976);
nand UO_483 (O_483,N_2952,N_2990);
and UO_484 (O_484,N_2979,N_2964);
or UO_485 (O_485,N_2970,N_2994);
nor UO_486 (O_486,N_2948,N_2977);
or UO_487 (O_487,N_2979,N_2972);
or UO_488 (O_488,N_2996,N_2967);
nor UO_489 (O_489,N_2957,N_2983);
nor UO_490 (O_490,N_2968,N_2962);
or UO_491 (O_491,N_2986,N_2957);
and UO_492 (O_492,N_2965,N_2993);
nor UO_493 (O_493,N_2953,N_2956);
nor UO_494 (O_494,N_2954,N_2946);
and UO_495 (O_495,N_2993,N_2958);
nand UO_496 (O_496,N_2949,N_2987);
and UO_497 (O_497,N_2949,N_2981);
and UO_498 (O_498,N_2987,N_2956);
nor UO_499 (O_499,N_2981,N_2959);
endmodule