module basic_500_3000_500_3_levels_1xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_453,In_439);
or U1 (N_1,In_466,In_250);
nand U2 (N_2,In_127,In_361);
nor U3 (N_3,In_224,In_0);
and U4 (N_4,In_99,In_151);
and U5 (N_5,In_420,In_273);
nor U6 (N_6,In_186,In_155);
or U7 (N_7,In_221,In_342);
nor U8 (N_8,In_67,In_440);
or U9 (N_9,In_109,In_122);
or U10 (N_10,In_33,In_265);
nor U11 (N_11,In_391,In_1);
or U12 (N_12,In_264,In_278);
nand U13 (N_13,In_362,In_302);
or U14 (N_14,In_415,In_102);
or U15 (N_15,In_179,In_73);
nor U16 (N_16,In_66,In_86);
nor U17 (N_17,In_484,In_424);
or U18 (N_18,In_245,In_171);
or U19 (N_19,In_54,In_492);
or U20 (N_20,In_57,In_84);
or U21 (N_21,In_108,In_296);
and U22 (N_22,In_293,In_305);
or U23 (N_23,In_287,In_412);
and U24 (N_24,In_358,In_206);
nor U25 (N_25,In_456,In_344);
nor U26 (N_26,In_208,In_71);
nor U27 (N_27,In_238,In_353);
or U28 (N_28,In_397,In_24);
or U29 (N_29,In_133,In_350);
or U30 (N_30,In_365,In_5);
or U31 (N_31,In_85,In_100);
or U32 (N_32,In_387,In_450);
and U33 (N_33,In_58,In_315);
and U34 (N_34,In_269,In_392);
nor U35 (N_35,In_113,In_174);
and U36 (N_36,In_438,In_8);
or U37 (N_37,In_129,In_246);
nand U38 (N_38,In_432,In_312);
or U39 (N_39,In_385,In_301);
nor U40 (N_40,In_96,In_21);
nor U41 (N_41,In_212,In_360);
and U42 (N_42,In_409,In_316);
nand U43 (N_43,In_156,In_338);
nand U44 (N_44,In_430,In_346);
nor U45 (N_45,In_343,In_395);
or U46 (N_46,In_259,In_261);
nand U47 (N_47,In_46,In_134);
or U48 (N_48,In_390,In_45);
nor U49 (N_49,In_427,In_354);
nand U50 (N_50,In_126,In_419);
and U51 (N_51,In_281,In_486);
nor U52 (N_52,In_447,In_410);
nor U53 (N_53,In_497,In_159);
nand U54 (N_54,In_405,In_407);
nor U55 (N_55,In_28,In_325);
nor U56 (N_56,In_203,In_334);
or U57 (N_57,In_388,In_393);
and U58 (N_58,In_496,In_426);
nor U59 (N_59,In_42,In_148);
and U60 (N_60,In_123,In_163);
nor U61 (N_61,In_394,In_51);
xor U62 (N_62,In_313,In_421);
or U63 (N_63,In_48,In_91);
nor U64 (N_64,In_194,In_181);
and U65 (N_65,In_472,In_105);
and U66 (N_66,In_168,In_76);
and U67 (N_67,In_90,In_452);
or U68 (N_68,In_317,In_470);
nand U69 (N_69,In_490,In_229);
and U70 (N_70,In_256,In_26);
or U71 (N_71,In_161,In_382);
nand U72 (N_72,In_364,In_23);
nand U73 (N_73,In_411,In_363);
nor U74 (N_74,In_272,In_49);
and U75 (N_75,In_384,In_266);
or U76 (N_76,In_72,In_132);
or U77 (N_77,In_286,In_489);
and U78 (N_78,In_199,In_477);
and U79 (N_79,In_60,In_241);
and U80 (N_80,In_95,In_173);
and U81 (N_81,In_31,In_308);
nor U82 (N_82,In_217,In_14);
or U83 (N_83,In_220,In_219);
and U84 (N_84,In_368,In_422);
and U85 (N_85,In_299,In_143);
and U86 (N_86,In_119,In_82);
or U87 (N_87,In_396,In_169);
and U88 (N_88,In_298,In_330);
nor U89 (N_89,In_383,In_189);
and U90 (N_90,In_16,In_11);
nand U91 (N_91,In_9,In_240);
and U92 (N_92,In_192,In_205);
nand U93 (N_93,In_112,In_116);
nor U94 (N_94,In_243,In_494);
or U95 (N_95,In_59,In_323);
or U96 (N_96,In_307,In_32);
nand U97 (N_97,In_337,In_235);
or U98 (N_98,In_107,In_333);
or U99 (N_99,In_137,In_157);
nand U100 (N_100,In_47,In_38);
nor U101 (N_101,In_320,In_445);
nor U102 (N_102,In_321,In_30);
nor U103 (N_103,In_247,In_190);
nor U104 (N_104,In_294,In_239);
or U105 (N_105,In_120,In_418);
nor U106 (N_106,In_331,In_252);
and U107 (N_107,In_288,In_69);
and U108 (N_108,In_372,In_7);
and U109 (N_109,In_202,In_423);
nand U110 (N_110,In_340,In_341);
nand U111 (N_111,In_454,In_399);
nor U112 (N_112,In_487,In_275);
nor U113 (N_113,In_480,In_175);
and U114 (N_114,In_25,In_34);
or U115 (N_115,In_77,In_3);
nor U116 (N_116,In_193,In_429);
nor U117 (N_117,In_43,In_416);
nand U118 (N_118,In_366,In_311);
nand U119 (N_119,In_81,In_306);
and U120 (N_120,In_22,In_130);
nand U121 (N_121,In_483,In_79);
and U122 (N_122,In_460,In_6);
nor U123 (N_123,In_242,In_117);
or U124 (N_124,In_431,In_128);
nand U125 (N_125,In_65,In_162);
and U126 (N_126,In_19,In_160);
nor U127 (N_127,In_377,In_324);
nor U128 (N_128,In_441,In_428);
and U129 (N_129,In_282,In_200);
nor U130 (N_130,In_491,In_40);
nor U131 (N_131,In_18,In_425);
nor U132 (N_132,In_61,In_178);
and U133 (N_133,In_124,In_17);
nor U134 (N_134,In_121,In_404);
nand U135 (N_135,In_12,In_446);
nand U136 (N_136,In_141,In_356);
nor U137 (N_137,In_231,In_253);
nand U138 (N_138,In_267,In_443);
nand U139 (N_139,In_164,In_255);
and U140 (N_140,In_166,In_2);
and U141 (N_141,In_499,In_335);
or U142 (N_142,In_111,In_464);
and U143 (N_143,In_214,In_131);
nand U144 (N_144,In_244,In_187);
nand U145 (N_145,In_101,In_336);
or U146 (N_146,In_234,In_165);
nand U147 (N_147,In_39,In_92);
or U148 (N_148,In_359,In_257);
nor U149 (N_149,In_370,In_115);
nor U150 (N_150,In_152,In_262);
nor U151 (N_151,In_196,In_218);
nor U152 (N_152,In_468,In_52);
nor U153 (N_153,In_44,In_13);
nor U154 (N_154,In_106,In_185);
nor U155 (N_155,In_145,In_433);
and U156 (N_156,In_20,In_222);
or U157 (N_157,In_318,In_74);
nor U158 (N_158,In_345,In_482);
nand U159 (N_159,In_332,In_118);
and U160 (N_160,In_457,In_451);
or U161 (N_161,In_94,In_455);
nor U162 (N_162,In_283,In_103);
nor U163 (N_163,In_211,In_413);
nor U164 (N_164,In_326,In_310);
nand U165 (N_165,In_437,In_41);
nor U166 (N_166,In_373,In_210);
or U167 (N_167,In_50,In_260);
nand U168 (N_168,In_488,In_4);
nor U169 (N_169,In_36,In_53);
and U170 (N_170,In_314,In_436);
or U171 (N_171,In_300,In_322);
nor U172 (N_172,In_458,In_276);
and U173 (N_173,In_474,In_328);
or U174 (N_174,In_435,In_434);
or U175 (N_175,In_184,In_64);
or U176 (N_176,In_70,In_291);
and U177 (N_177,In_198,In_402);
nand U178 (N_178,In_467,In_417);
and U179 (N_179,In_62,In_97);
and U180 (N_180,In_449,In_195);
or U181 (N_181,In_476,In_297);
nor U182 (N_182,In_380,In_459);
nand U183 (N_183,In_478,In_149);
and U184 (N_184,In_191,In_254);
nor U185 (N_185,In_237,In_248);
nor U186 (N_186,In_140,In_147);
nand U187 (N_187,In_270,In_56);
or U188 (N_188,In_183,In_158);
nor U189 (N_189,In_233,In_227);
nand U190 (N_190,In_292,In_498);
nand U191 (N_191,In_369,In_87);
xnor U192 (N_192,In_136,In_448);
nand U193 (N_193,In_35,In_172);
or U194 (N_194,In_274,In_479);
nor U195 (N_195,In_357,In_68);
nand U196 (N_196,In_280,In_375);
nand U197 (N_197,In_493,In_277);
or U198 (N_198,In_406,In_327);
and U199 (N_199,In_379,In_176);
and U200 (N_200,In_88,In_376);
or U201 (N_201,In_347,In_125);
and U202 (N_202,In_444,In_93);
nor U203 (N_203,In_495,In_304);
nor U204 (N_204,In_263,In_230);
nor U205 (N_205,In_400,In_27);
nand U206 (N_206,In_177,In_351);
or U207 (N_207,In_371,In_290);
nor U208 (N_208,In_374,In_188);
or U209 (N_209,In_398,In_228);
or U210 (N_210,In_75,In_139);
nand U211 (N_211,In_110,In_207);
nand U212 (N_212,In_461,In_10);
nor U213 (N_213,In_98,In_89);
or U214 (N_214,In_401,In_268);
nand U215 (N_215,In_349,In_170);
or U216 (N_216,In_209,In_462);
or U217 (N_217,In_226,In_232);
nand U218 (N_218,In_180,In_150);
nand U219 (N_219,In_348,In_329);
nand U220 (N_220,In_469,In_271);
and U221 (N_221,In_142,In_37);
and U222 (N_222,In_167,In_197);
and U223 (N_223,In_114,In_463);
or U224 (N_224,In_309,In_485);
or U225 (N_225,In_146,In_144);
nand U226 (N_226,In_471,In_475);
or U227 (N_227,In_442,In_204);
nor U228 (N_228,In_481,In_182);
and U229 (N_229,In_319,In_153);
and U230 (N_230,In_389,In_83);
and U231 (N_231,In_289,In_225);
and U232 (N_232,In_78,In_213);
or U233 (N_233,In_63,In_473);
and U234 (N_234,In_279,In_414);
nand U235 (N_235,In_154,In_258);
or U236 (N_236,In_352,In_355);
or U237 (N_237,In_339,In_249);
and U238 (N_238,In_80,In_216);
and U239 (N_239,In_285,In_386);
or U240 (N_240,In_251,In_236);
and U241 (N_241,In_104,In_284);
nor U242 (N_242,In_15,In_378);
or U243 (N_243,In_138,In_403);
or U244 (N_244,In_223,In_55);
nand U245 (N_245,In_215,In_201);
nor U246 (N_246,In_295,In_465);
and U247 (N_247,In_135,In_381);
or U248 (N_248,In_303,In_367);
or U249 (N_249,In_29,In_408);
or U250 (N_250,In_324,In_253);
nor U251 (N_251,In_416,In_369);
nor U252 (N_252,In_128,In_376);
nor U253 (N_253,In_378,In_360);
xor U254 (N_254,In_417,In_355);
nor U255 (N_255,In_205,In_263);
nand U256 (N_256,In_216,In_441);
and U257 (N_257,In_254,In_186);
or U258 (N_258,In_348,In_136);
and U259 (N_259,In_3,In_496);
nand U260 (N_260,In_127,In_414);
or U261 (N_261,In_152,In_153);
or U262 (N_262,In_462,In_135);
nor U263 (N_263,In_299,In_185);
and U264 (N_264,In_116,In_392);
or U265 (N_265,In_52,In_215);
nand U266 (N_266,In_43,In_208);
or U267 (N_267,In_147,In_195);
and U268 (N_268,In_415,In_20);
or U269 (N_269,In_3,In_288);
nand U270 (N_270,In_246,In_465);
nand U271 (N_271,In_79,In_181);
and U272 (N_272,In_382,In_278);
xor U273 (N_273,In_44,In_86);
or U274 (N_274,In_396,In_287);
or U275 (N_275,In_221,In_409);
or U276 (N_276,In_455,In_112);
and U277 (N_277,In_190,In_104);
or U278 (N_278,In_444,In_87);
or U279 (N_279,In_495,In_130);
and U280 (N_280,In_16,In_497);
nand U281 (N_281,In_240,In_346);
or U282 (N_282,In_101,In_93);
and U283 (N_283,In_481,In_136);
nor U284 (N_284,In_85,In_411);
nor U285 (N_285,In_482,In_199);
nand U286 (N_286,In_279,In_209);
nor U287 (N_287,In_153,In_159);
nor U288 (N_288,In_489,In_27);
nor U289 (N_289,In_65,In_412);
nand U290 (N_290,In_417,In_159);
and U291 (N_291,In_363,In_100);
nor U292 (N_292,In_296,In_12);
nand U293 (N_293,In_221,In_255);
and U294 (N_294,In_80,In_305);
nor U295 (N_295,In_484,In_20);
and U296 (N_296,In_162,In_214);
nor U297 (N_297,In_478,In_433);
and U298 (N_298,In_54,In_471);
and U299 (N_299,In_272,In_144);
or U300 (N_300,In_70,In_64);
nand U301 (N_301,In_132,In_265);
and U302 (N_302,In_445,In_126);
and U303 (N_303,In_288,In_70);
and U304 (N_304,In_399,In_475);
nor U305 (N_305,In_220,In_282);
nand U306 (N_306,In_425,In_311);
nor U307 (N_307,In_465,In_129);
or U308 (N_308,In_424,In_113);
and U309 (N_309,In_379,In_326);
nand U310 (N_310,In_369,In_190);
and U311 (N_311,In_230,In_455);
nor U312 (N_312,In_333,In_211);
or U313 (N_313,In_304,In_158);
or U314 (N_314,In_43,In_349);
nor U315 (N_315,In_400,In_489);
nand U316 (N_316,In_244,In_146);
and U317 (N_317,In_186,In_101);
nand U318 (N_318,In_329,In_54);
or U319 (N_319,In_492,In_309);
or U320 (N_320,In_237,In_83);
nor U321 (N_321,In_497,In_327);
nand U322 (N_322,In_380,In_202);
nor U323 (N_323,In_312,In_329);
nor U324 (N_324,In_306,In_159);
and U325 (N_325,In_262,In_17);
nand U326 (N_326,In_183,In_311);
or U327 (N_327,In_198,In_319);
nor U328 (N_328,In_130,In_93);
or U329 (N_329,In_181,In_453);
nor U330 (N_330,In_257,In_26);
nor U331 (N_331,In_240,In_219);
or U332 (N_332,In_408,In_484);
and U333 (N_333,In_420,In_36);
nand U334 (N_334,In_40,In_360);
and U335 (N_335,In_10,In_55);
or U336 (N_336,In_172,In_160);
and U337 (N_337,In_195,In_310);
nor U338 (N_338,In_199,In_391);
and U339 (N_339,In_209,In_489);
or U340 (N_340,In_236,In_302);
nor U341 (N_341,In_433,In_80);
nand U342 (N_342,In_290,In_291);
or U343 (N_343,In_196,In_301);
nand U344 (N_344,In_332,In_257);
or U345 (N_345,In_134,In_404);
and U346 (N_346,In_378,In_77);
or U347 (N_347,In_145,In_377);
nand U348 (N_348,In_136,In_241);
nand U349 (N_349,In_182,In_459);
nand U350 (N_350,In_343,In_419);
or U351 (N_351,In_285,In_416);
nor U352 (N_352,In_455,In_405);
nand U353 (N_353,In_238,In_400);
nor U354 (N_354,In_297,In_175);
or U355 (N_355,In_407,In_119);
and U356 (N_356,In_170,In_45);
nor U357 (N_357,In_408,In_335);
nor U358 (N_358,In_360,In_284);
nor U359 (N_359,In_242,In_218);
nand U360 (N_360,In_75,In_275);
nand U361 (N_361,In_217,In_132);
and U362 (N_362,In_437,In_127);
nand U363 (N_363,In_106,In_34);
nand U364 (N_364,In_188,In_184);
and U365 (N_365,In_325,In_422);
nand U366 (N_366,In_371,In_115);
nor U367 (N_367,In_269,In_233);
and U368 (N_368,In_7,In_253);
and U369 (N_369,In_441,In_20);
nor U370 (N_370,In_158,In_479);
and U371 (N_371,In_496,In_173);
nand U372 (N_372,In_407,In_411);
nand U373 (N_373,In_388,In_215);
nor U374 (N_374,In_493,In_217);
nand U375 (N_375,In_479,In_240);
nand U376 (N_376,In_412,In_372);
nor U377 (N_377,In_5,In_7);
and U378 (N_378,In_456,In_123);
and U379 (N_379,In_187,In_77);
nand U380 (N_380,In_417,In_345);
or U381 (N_381,In_314,In_161);
and U382 (N_382,In_311,In_22);
nor U383 (N_383,In_133,In_78);
or U384 (N_384,In_361,In_142);
or U385 (N_385,In_417,In_379);
or U386 (N_386,In_217,In_382);
and U387 (N_387,In_115,In_48);
or U388 (N_388,In_342,In_328);
nor U389 (N_389,In_389,In_443);
and U390 (N_390,In_3,In_186);
nand U391 (N_391,In_82,In_275);
nor U392 (N_392,In_261,In_294);
nor U393 (N_393,In_379,In_60);
nor U394 (N_394,In_67,In_4);
nor U395 (N_395,In_259,In_41);
nor U396 (N_396,In_148,In_369);
nor U397 (N_397,In_481,In_458);
and U398 (N_398,In_22,In_127);
nand U399 (N_399,In_380,In_295);
and U400 (N_400,In_350,In_410);
nand U401 (N_401,In_123,In_31);
and U402 (N_402,In_483,In_460);
nand U403 (N_403,In_252,In_401);
nand U404 (N_404,In_105,In_22);
and U405 (N_405,In_112,In_208);
or U406 (N_406,In_193,In_247);
or U407 (N_407,In_312,In_203);
and U408 (N_408,In_450,In_247);
nand U409 (N_409,In_363,In_351);
or U410 (N_410,In_426,In_153);
or U411 (N_411,In_483,In_211);
or U412 (N_412,In_347,In_291);
or U413 (N_413,In_298,In_487);
or U414 (N_414,In_324,In_471);
or U415 (N_415,In_209,In_253);
or U416 (N_416,In_460,In_324);
or U417 (N_417,In_357,In_268);
nor U418 (N_418,In_340,In_203);
or U419 (N_419,In_207,In_462);
or U420 (N_420,In_147,In_27);
xnor U421 (N_421,In_215,In_344);
and U422 (N_422,In_41,In_169);
and U423 (N_423,In_260,In_395);
or U424 (N_424,In_282,In_218);
or U425 (N_425,In_126,In_72);
or U426 (N_426,In_233,In_398);
or U427 (N_427,In_60,In_339);
nand U428 (N_428,In_384,In_322);
and U429 (N_429,In_257,In_389);
nand U430 (N_430,In_45,In_112);
and U431 (N_431,In_369,In_375);
or U432 (N_432,In_247,In_30);
or U433 (N_433,In_499,In_300);
nand U434 (N_434,In_149,In_7);
nor U435 (N_435,In_381,In_85);
or U436 (N_436,In_377,In_374);
or U437 (N_437,In_351,In_34);
or U438 (N_438,In_116,In_292);
nor U439 (N_439,In_60,In_232);
nand U440 (N_440,In_122,In_313);
and U441 (N_441,In_82,In_153);
and U442 (N_442,In_485,In_124);
nand U443 (N_443,In_137,In_162);
nor U444 (N_444,In_159,In_60);
nand U445 (N_445,In_138,In_440);
nand U446 (N_446,In_437,In_156);
nand U447 (N_447,In_404,In_438);
nand U448 (N_448,In_99,In_361);
and U449 (N_449,In_162,In_377);
nor U450 (N_450,In_422,In_138);
or U451 (N_451,In_139,In_174);
or U452 (N_452,In_28,In_421);
or U453 (N_453,In_357,In_52);
nand U454 (N_454,In_440,In_142);
nor U455 (N_455,In_232,In_177);
and U456 (N_456,In_348,In_38);
or U457 (N_457,In_307,In_193);
nand U458 (N_458,In_325,In_367);
or U459 (N_459,In_188,In_291);
nor U460 (N_460,In_273,In_51);
nand U461 (N_461,In_337,In_316);
nand U462 (N_462,In_215,In_351);
and U463 (N_463,In_161,In_52);
nor U464 (N_464,In_467,In_481);
nor U465 (N_465,In_278,In_454);
and U466 (N_466,In_45,In_381);
or U467 (N_467,In_497,In_422);
nand U468 (N_468,In_49,In_255);
nand U469 (N_469,In_256,In_320);
and U470 (N_470,In_446,In_277);
and U471 (N_471,In_203,In_246);
nand U472 (N_472,In_324,In_466);
or U473 (N_473,In_216,In_49);
and U474 (N_474,In_78,In_455);
or U475 (N_475,In_100,In_135);
or U476 (N_476,In_449,In_328);
nor U477 (N_477,In_331,In_40);
nand U478 (N_478,In_111,In_223);
nor U479 (N_479,In_239,In_236);
or U480 (N_480,In_376,In_268);
or U481 (N_481,In_210,In_362);
nand U482 (N_482,In_206,In_425);
and U483 (N_483,In_146,In_405);
xnor U484 (N_484,In_45,In_442);
and U485 (N_485,In_459,In_206);
nand U486 (N_486,In_376,In_119);
and U487 (N_487,In_141,In_373);
nor U488 (N_488,In_296,In_444);
nor U489 (N_489,In_346,In_11);
nor U490 (N_490,In_466,In_190);
nand U491 (N_491,In_413,In_66);
nor U492 (N_492,In_116,In_418);
nand U493 (N_493,In_351,In_247);
or U494 (N_494,In_140,In_115);
nand U495 (N_495,In_52,In_279);
nor U496 (N_496,In_168,In_167);
or U497 (N_497,In_11,In_447);
or U498 (N_498,In_92,In_333);
nor U499 (N_499,In_386,In_345);
or U500 (N_500,In_236,In_207);
xnor U501 (N_501,In_54,In_206);
nand U502 (N_502,In_326,In_354);
nor U503 (N_503,In_199,In_490);
and U504 (N_504,In_247,In_311);
and U505 (N_505,In_320,In_448);
nand U506 (N_506,In_232,In_157);
nor U507 (N_507,In_98,In_224);
and U508 (N_508,In_468,In_343);
and U509 (N_509,In_115,In_301);
nand U510 (N_510,In_108,In_268);
nor U511 (N_511,In_314,In_30);
nor U512 (N_512,In_308,In_413);
nand U513 (N_513,In_107,In_20);
nand U514 (N_514,In_75,In_98);
and U515 (N_515,In_151,In_475);
or U516 (N_516,In_485,In_288);
nor U517 (N_517,In_12,In_165);
nor U518 (N_518,In_145,In_355);
nor U519 (N_519,In_458,In_443);
or U520 (N_520,In_257,In_439);
and U521 (N_521,In_449,In_347);
and U522 (N_522,In_60,In_213);
nor U523 (N_523,In_463,In_354);
and U524 (N_524,In_330,In_131);
nor U525 (N_525,In_10,In_495);
or U526 (N_526,In_127,In_3);
and U527 (N_527,In_166,In_109);
nand U528 (N_528,In_137,In_254);
nand U529 (N_529,In_487,In_301);
and U530 (N_530,In_300,In_424);
or U531 (N_531,In_129,In_254);
and U532 (N_532,In_460,In_315);
and U533 (N_533,In_487,In_363);
and U534 (N_534,In_163,In_173);
nor U535 (N_535,In_392,In_329);
and U536 (N_536,In_186,In_386);
and U537 (N_537,In_364,In_77);
or U538 (N_538,In_452,In_439);
or U539 (N_539,In_231,In_247);
nor U540 (N_540,In_289,In_222);
nor U541 (N_541,In_365,In_136);
nand U542 (N_542,In_326,In_469);
and U543 (N_543,In_167,In_458);
nor U544 (N_544,In_421,In_241);
nand U545 (N_545,In_66,In_455);
or U546 (N_546,In_274,In_281);
and U547 (N_547,In_87,In_400);
nand U548 (N_548,In_4,In_33);
and U549 (N_549,In_346,In_99);
nor U550 (N_550,In_123,In_433);
nand U551 (N_551,In_53,In_472);
and U552 (N_552,In_487,In_314);
nor U553 (N_553,In_140,In_466);
nand U554 (N_554,In_180,In_269);
and U555 (N_555,In_190,In_197);
and U556 (N_556,In_446,In_360);
nor U557 (N_557,In_341,In_312);
nand U558 (N_558,In_342,In_242);
nand U559 (N_559,In_15,In_325);
or U560 (N_560,In_295,In_338);
nand U561 (N_561,In_368,In_249);
and U562 (N_562,In_287,In_368);
nand U563 (N_563,In_390,In_269);
nor U564 (N_564,In_358,In_480);
or U565 (N_565,In_154,In_69);
nor U566 (N_566,In_444,In_68);
nand U567 (N_567,In_364,In_300);
or U568 (N_568,In_1,In_410);
nor U569 (N_569,In_80,In_112);
nor U570 (N_570,In_390,In_279);
and U571 (N_571,In_29,In_92);
nand U572 (N_572,In_462,In_108);
and U573 (N_573,In_62,In_86);
or U574 (N_574,In_417,In_357);
nand U575 (N_575,In_61,In_265);
or U576 (N_576,In_263,In_343);
nand U577 (N_577,In_376,In_47);
nor U578 (N_578,In_486,In_170);
and U579 (N_579,In_117,In_386);
or U580 (N_580,In_184,In_325);
nor U581 (N_581,In_245,In_265);
nor U582 (N_582,In_484,In_324);
or U583 (N_583,In_70,In_102);
nand U584 (N_584,In_79,In_24);
and U585 (N_585,In_312,In_442);
or U586 (N_586,In_382,In_406);
nand U587 (N_587,In_261,In_80);
or U588 (N_588,In_159,In_32);
or U589 (N_589,In_66,In_105);
nand U590 (N_590,In_263,In_131);
and U591 (N_591,In_439,In_228);
nor U592 (N_592,In_217,In_44);
nor U593 (N_593,In_474,In_382);
or U594 (N_594,In_105,In_345);
or U595 (N_595,In_346,In_145);
or U596 (N_596,In_207,In_337);
and U597 (N_597,In_106,In_256);
nor U598 (N_598,In_326,In_125);
nor U599 (N_599,In_44,In_274);
and U600 (N_600,In_23,In_176);
nand U601 (N_601,In_213,In_260);
and U602 (N_602,In_144,In_410);
xnor U603 (N_603,In_52,In_450);
nor U604 (N_604,In_457,In_57);
nand U605 (N_605,In_367,In_112);
or U606 (N_606,In_46,In_401);
nor U607 (N_607,In_364,In_138);
nor U608 (N_608,In_8,In_74);
nand U609 (N_609,In_278,In_221);
xnor U610 (N_610,In_399,In_412);
nor U611 (N_611,In_2,In_104);
nand U612 (N_612,In_372,In_403);
nor U613 (N_613,In_91,In_269);
nor U614 (N_614,In_42,In_163);
nor U615 (N_615,In_276,In_385);
nand U616 (N_616,In_460,In_346);
and U617 (N_617,In_470,In_401);
and U618 (N_618,In_351,In_226);
and U619 (N_619,In_138,In_320);
or U620 (N_620,In_319,In_427);
nand U621 (N_621,In_447,In_418);
or U622 (N_622,In_309,In_97);
and U623 (N_623,In_4,In_487);
and U624 (N_624,In_417,In_269);
and U625 (N_625,In_469,In_47);
nor U626 (N_626,In_200,In_487);
or U627 (N_627,In_201,In_245);
nand U628 (N_628,In_363,In_68);
nand U629 (N_629,In_313,In_468);
and U630 (N_630,In_3,In_72);
nand U631 (N_631,In_273,In_70);
nor U632 (N_632,In_246,In_187);
nor U633 (N_633,In_55,In_382);
nor U634 (N_634,In_124,In_413);
xor U635 (N_635,In_341,In_441);
nand U636 (N_636,In_170,In_247);
nand U637 (N_637,In_108,In_337);
or U638 (N_638,In_416,In_244);
and U639 (N_639,In_154,In_361);
or U640 (N_640,In_275,In_154);
nor U641 (N_641,In_325,In_59);
nor U642 (N_642,In_281,In_369);
nor U643 (N_643,In_285,In_88);
and U644 (N_644,In_413,In_162);
nand U645 (N_645,In_305,In_492);
nor U646 (N_646,In_488,In_290);
nand U647 (N_647,In_327,In_243);
nand U648 (N_648,In_371,In_13);
nor U649 (N_649,In_77,In_300);
nand U650 (N_650,In_434,In_328);
and U651 (N_651,In_480,In_303);
nand U652 (N_652,In_169,In_354);
nand U653 (N_653,In_214,In_320);
or U654 (N_654,In_121,In_234);
nor U655 (N_655,In_93,In_91);
nand U656 (N_656,In_439,In_422);
nor U657 (N_657,In_376,In_136);
or U658 (N_658,In_80,In_49);
nor U659 (N_659,In_326,In_485);
and U660 (N_660,In_39,In_64);
nor U661 (N_661,In_29,In_493);
and U662 (N_662,In_391,In_418);
and U663 (N_663,In_166,In_286);
and U664 (N_664,In_484,In_225);
nand U665 (N_665,In_427,In_204);
nand U666 (N_666,In_252,In_211);
nand U667 (N_667,In_37,In_416);
and U668 (N_668,In_241,In_7);
and U669 (N_669,In_436,In_440);
or U670 (N_670,In_21,In_170);
or U671 (N_671,In_95,In_499);
and U672 (N_672,In_368,In_188);
nor U673 (N_673,In_320,In_362);
nor U674 (N_674,In_464,In_99);
and U675 (N_675,In_322,In_337);
or U676 (N_676,In_492,In_198);
nor U677 (N_677,In_18,In_105);
and U678 (N_678,In_160,In_103);
and U679 (N_679,In_333,In_41);
nand U680 (N_680,In_301,In_43);
nand U681 (N_681,In_465,In_390);
or U682 (N_682,In_15,In_459);
xnor U683 (N_683,In_87,In_476);
or U684 (N_684,In_459,In_404);
or U685 (N_685,In_499,In_313);
and U686 (N_686,In_231,In_66);
nor U687 (N_687,In_432,In_284);
and U688 (N_688,In_446,In_395);
or U689 (N_689,In_22,In_378);
or U690 (N_690,In_473,In_13);
nor U691 (N_691,In_487,In_55);
or U692 (N_692,In_148,In_74);
and U693 (N_693,In_197,In_70);
nor U694 (N_694,In_196,In_393);
nand U695 (N_695,In_279,In_263);
or U696 (N_696,In_420,In_89);
nand U697 (N_697,In_446,In_376);
and U698 (N_698,In_210,In_134);
nand U699 (N_699,In_271,In_141);
and U700 (N_700,In_381,In_138);
nand U701 (N_701,In_347,In_355);
and U702 (N_702,In_354,In_117);
nand U703 (N_703,In_394,In_341);
or U704 (N_704,In_275,In_32);
nand U705 (N_705,In_182,In_397);
or U706 (N_706,In_246,In_403);
and U707 (N_707,In_446,In_80);
nor U708 (N_708,In_268,In_296);
or U709 (N_709,In_259,In_407);
and U710 (N_710,In_132,In_220);
and U711 (N_711,In_380,In_150);
or U712 (N_712,In_171,In_423);
or U713 (N_713,In_425,In_342);
and U714 (N_714,In_306,In_264);
and U715 (N_715,In_128,In_51);
nor U716 (N_716,In_243,In_292);
or U717 (N_717,In_234,In_362);
nor U718 (N_718,In_401,In_56);
nand U719 (N_719,In_25,In_123);
or U720 (N_720,In_197,In_253);
nand U721 (N_721,In_133,In_256);
nor U722 (N_722,In_285,In_126);
or U723 (N_723,In_64,In_111);
or U724 (N_724,In_490,In_114);
and U725 (N_725,In_323,In_128);
and U726 (N_726,In_289,In_382);
and U727 (N_727,In_40,In_202);
and U728 (N_728,In_445,In_427);
nor U729 (N_729,In_194,In_48);
nor U730 (N_730,In_52,In_395);
nand U731 (N_731,In_310,In_142);
nand U732 (N_732,In_182,In_83);
nor U733 (N_733,In_0,In_294);
nor U734 (N_734,In_457,In_123);
and U735 (N_735,In_272,In_252);
nor U736 (N_736,In_269,In_149);
and U737 (N_737,In_116,In_80);
or U738 (N_738,In_268,In_448);
and U739 (N_739,In_117,In_311);
nand U740 (N_740,In_134,In_278);
or U741 (N_741,In_200,In_337);
nor U742 (N_742,In_441,In_473);
nor U743 (N_743,In_82,In_91);
nor U744 (N_744,In_9,In_449);
nor U745 (N_745,In_68,In_259);
nor U746 (N_746,In_239,In_438);
and U747 (N_747,In_71,In_117);
nor U748 (N_748,In_411,In_312);
or U749 (N_749,In_178,In_45);
or U750 (N_750,In_354,In_15);
nor U751 (N_751,In_442,In_371);
or U752 (N_752,In_258,In_415);
nand U753 (N_753,In_270,In_3);
nand U754 (N_754,In_411,In_175);
nand U755 (N_755,In_65,In_295);
nor U756 (N_756,In_37,In_250);
and U757 (N_757,In_383,In_144);
nor U758 (N_758,In_408,In_364);
and U759 (N_759,In_195,In_114);
nor U760 (N_760,In_74,In_48);
or U761 (N_761,In_176,In_234);
and U762 (N_762,In_297,In_454);
or U763 (N_763,In_149,In_119);
and U764 (N_764,In_295,In_247);
nor U765 (N_765,In_461,In_442);
nor U766 (N_766,In_379,In_80);
nand U767 (N_767,In_402,In_73);
and U768 (N_768,In_137,In_10);
or U769 (N_769,In_297,In_355);
and U770 (N_770,In_178,In_356);
and U771 (N_771,In_426,In_17);
nand U772 (N_772,In_491,In_5);
and U773 (N_773,In_33,In_166);
and U774 (N_774,In_368,In_384);
nor U775 (N_775,In_195,In_408);
or U776 (N_776,In_222,In_113);
nor U777 (N_777,In_112,In_354);
nand U778 (N_778,In_166,In_127);
nand U779 (N_779,In_426,In_335);
nor U780 (N_780,In_115,In_87);
nand U781 (N_781,In_62,In_349);
or U782 (N_782,In_71,In_423);
nor U783 (N_783,In_89,In_491);
nand U784 (N_784,In_358,In_360);
nor U785 (N_785,In_19,In_405);
nand U786 (N_786,In_316,In_38);
nor U787 (N_787,In_482,In_305);
or U788 (N_788,In_339,In_456);
nand U789 (N_789,In_134,In_167);
or U790 (N_790,In_153,In_116);
or U791 (N_791,In_31,In_392);
or U792 (N_792,In_119,In_293);
and U793 (N_793,In_228,In_239);
or U794 (N_794,In_440,In_423);
nand U795 (N_795,In_161,In_365);
nor U796 (N_796,In_386,In_89);
and U797 (N_797,In_257,In_295);
nor U798 (N_798,In_322,In_423);
or U799 (N_799,In_2,In_72);
or U800 (N_800,In_98,In_378);
nor U801 (N_801,In_56,In_143);
nor U802 (N_802,In_232,In_20);
or U803 (N_803,In_164,In_296);
and U804 (N_804,In_17,In_352);
and U805 (N_805,In_223,In_221);
nor U806 (N_806,In_371,In_243);
and U807 (N_807,In_466,In_420);
nand U808 (N_808,In_125,In_203);
and U809 (N_809,In_457,In_287);
nor U810 (N_810,In_386,In_300);
and U811 (N_811,In_130,In_79);
nor U812 (N_812,In_484,In_343);
nor U813 (N_813,In_440,In_70);
xnor U814 (N_814,In_112,In_254);
nor U815 (N_815,In_496,In_11);
nor U816 (N_816,In_167,In_476);
nor U817 (N_817,In_150,In_383);
nor U818 (N_818,In_194,In_14);
nor U819 (N_819,In_401,In_231);
or U820 (N_820,In_192,In_466);
and U821 (N_821,In_361,In_434);
or U822 (N_822,In_475,In_324);
and U823 (N_823,In_37,In_404);
or U824 (N_824,In_241,In_329);
or U825 (N_825,In_43,In_493);
nand U826 (N_826,In_397,In_453);
nor U827 (N_827,In_299,In_178);
or U828 (N_828,In_10,In_342);
and U829 (N_829,In_131,In_467);
nor U830 (N_830,In_50,In_46);
xnor U831 (N_831,In_66,In_474);
or U832 (N_832,In_234,In_410);
nand U833 (N_833,In_180,In_340);
or U834 (N_834,In_462,In_168);
nand U835 (N_835,In_470,In_262);
and U836 (N_836,In_382,In_266);
nand U837 (N_837,In_471,In_356);
and U838 (N_838,In_208,In_247);
nand U839 (N_839,In_498,In_158);
nand U840 (N_840,In_304,In_314);
or U841 (N_841,In_31,In_145);
or U842 (N_842,In_231,In_23);
nand U843 (N_843,In_379,In_361);
and U844 (N_844,In_12,In_56);
nor U845 (N_845,In_401,In_468);
or U846 (N_846,In_406,In_331);
nand U847 (N_847,In_325,In_338);
nor U848 (N_848,In_330,In_143);
and U849 (N_849,In_412,In_239);
nor U850 (N_850,In_136,In_296);
nor U851 (N_851,In_370,In_91);
nor U852 (N_852,In_205,In_127);
nor U853 (N_853,In_347,In_156);
or U854 (N_854,In_8,In_309);
nand U855 (N_855,In_314,In_276);
xnor U856 (N_856,In_484,In_18);
nand U857 (N_857,In_153,In_351);
or U858 (N_858,In_295,In_260);
and U859 (N_859,In_60,In_454);
nor U860 (N_860,In_157,In_28);
nor U861 (N_861,In_103,In_179);
nor U862 (N_862,In_136,In_425);
nor U863 (N_863,In_483,In_329);
or U864 (N_864,In_92,In_491);
nor U865 (N_865,In_347,In_264);
nor U866 (N_866,In_497,In_289);
or U867 (N_867,In_241,In_349);
nor U868 (N_868,In_249,In_235);
and U869 (N_869,In_395,In_407);
and U870 (N_870,In_385,In_168);
nand U871 (N_871,In_413,In_202);
or U872 (N_872,In_369,In_186);
nor U873 (N_873,In_430,In_89);
and U874 (N_874,In_207,In_133);
and U875 (N_875,In_257,In_40);
nor U876 (N_876,In_194,In_493);
nand U877 (N_877,In_443,In_466);
nand U878 (N_878,In_383,In_467);
nand U879 (N_879,In_376,In_358);
nor U880 (N_880,In_309,In_299);
nand U881 (N_881,In_451,In_4);
nor U882 (N_882,In_291,In_54);
nor U883 (N_883,In_117,In_432);
and U884 (N_884,In_116,In_79);
and U885 (N_885,In_154,In_232);
or U886 (N_886,In_302,In_73);
nor U887 (N_887,In_327,In_269);
nand U888 (N_888,In_248,In_341);
nor U889 (N_889,In_232,In_29);
nand U890 (N_890,In_360,In_171);
and U891 (N_891,In_416,In_374);
or U892 (N_892,In_350,In_138);
nor U893 (N_893,In_92,In_492);
nand U894 (N_894,In_55,In_145);
nand U895 (N_895,In_184,In_469);
or U896 (N_896,In_363,In_52);
or U897 (N_897,In_274,In_193);
nand U898 (N_898,In_245,In_163);
or U899 (N_899,In_422,In_29);
or U900 (N_900,In_275,In_81);
or U901 (N_901,In_257,In_334);
xor U902 (N_902,In_168,In_307);
and U903 (N_903,In_334,In_48);
nand U904 (N_904,In_149,In_103);
nor U905 (N_905,In_31,In_69);
or U906 (N_906,In_495,In_443);
nand U907 (N_907,In_247,In_270);
or U908 (N_908,In_146,In_130);
nand U909 (N_909,In_54,In_411);
and U910 (N_910,In_474,In_273);
nor U911 (N_911,In_488,In_446);
nand U912 (N_912,In_26,In_314);
nand U913 (N_913,In_412,In_244);
nor U914 (N_914,In_458,In_146);
nor U915 (N_915,In_145,In_6);
nor U916 (N_916,In_114,In_78);
nand U917 (N_917,In_90,In_422);
nor U918 (N_918,In_423,In_416);
or U919 (N_919,In_475,In_90);
nor U920 (N_920,In_432,In_209);
or U921 (N_921,In_10,In_438);
or U922 (N_922,In_102,In_30);
or U923 (N_923,In_125,In_254);
nor U924 (N_924,In_381,In_456);
nand U925 (N_925,In_261,In_192);
nand U926 (N_926,In_170,In_442);
or U927 (N_927,In_243,In_87);
or U928 (N_928,In_456,In_406);
and U929 (N_929,In_30,In_112);
nor U930 (N_930,In_390,In_240);
nor U931 (N_931,In_167,In_207);
nand U932 (N_932,In_28,In_292);
or U933 (N_933,In_391,In_136);
or U934 (N_934,In_76,In_82);
nand U935 (N_935,In_391,In_135);
nor U936 (N_936,In_359,In_404);
and U937 (N_937,In_88,In_463);
and U938 (N_938,In_107,In_148);
nand U939 (N_939,In_475,In_321);
and U940 (N_940,In_53,In_296);
and U941 (N_941,In_481,In_242);
nand U942 (N_942,In_310,In_396);
or U943 (N_943,In_429,In_343);
nand U944 (N_944,In_440,In_497);
or U945 (N_945,In_246,In_199);
nor U946 (N_946,In_445,In_418);
nand U947 (N_947,In_324,In_286);
nand U948 (N_948,In_389,In_65);
and U949 (N_949,In_129,In_2);
nor U950 (N_950,In_34,In_353);
nand U951 (N_951,In_228,In_250);
or U952 (N_952,In_309,In_369);
and U953 (N_953,In_237,In_252);
nand U954 (N_954,In_241,In_351);
and U955 (N_955,In_219,In_145);
and U956 (N_956,In_314,In_271);
or U957 (N_957,In_494,In_12);
and U958 (N_958,In_347,In_489);
nor U959 (N_959,In_406,In_407);
nor U960 (N_960,In_25,In_467);
or U961 (N_961,In_60,In_334);
or U962 (N_962,In_37,In_3);
nor U963 (N_963,In_258,In_114);
or U964 (N_964,In_435,In_40);
nand U965 (N_965,In_114,In_443);
or U966 (N_966,In_384,In_255);
nand U967 (N_967,In_5,In_132);
and U968 (N_968,In_27,In_334);
nand U969 (N_969,In_472,In_171);
nand U970 (N_970,In_352,In_132);
or U971 (N_971,In_430,In_78);
nor U972 (N_972,In_142,In_170);
or U973 (N_973,In_314,In_441);
nor U974 (N_974,In_341,In_349);
and U975 (N_975,In_341,In_101);
nand U976 (N_976,In_331,In_239);
or U977 (N_977,In_195,In_296);
and U978 (N_978,In_138,In_287);
and U979 (N_979,In_36,In_357);
or U980 (N_980,In_469,In_445);
and U981 (N_981,In_291,In_342);
and U982 (N_982,In_220,In_98);
nor U983 (N_983,In_31,In_192);
or U984 (N_984,In_258,In_28);
and U985 (N_985,In_491,In_387);
and U986 (N_986,In_31,In_56);
nor U987 (N_987,In_356,In_2);
nand U988 (N_988,In_68,In_478);
nand U989 (N_989,In_491,In_496);
nor U990 (N_990,In_499,In_241);
or U991 (N_991,In_74,In_365);
or U992 (N_992,In_343,In_210);
and U993 (N_993,In_181,In_51);
or U994 (N_994,In_101,In_384);
nor U995 (N_995,In_307,In_452);
and U996 (N_996,In_292,In_123);
xor U997 (N_997,In_273,In_423);
nor U998 (N_998,In_170,In_51);
or U999 (N_999,In_479,In_307);
nand U1000 (N_1000,N_451,N_478);
or U1001 (N_1001,N_593,N_261);
and U1002 (N_1002,N_707,N_165);
and U1003 (N_1003,N_872,N_610);
nand U1004 (N_1004,N_7,N_268);
or U1005 (N_1005,N_605,N_699);
or U1006 (N_1006,N_555,N_4);
or U1007 (N_1007,N_295,N_603);
and U1008 (N_1008,N_221,N_586);
and U1009 (N_1009,N_401,N_568);
nor U1010 (N_1010,N_829,N_766);
nand U1011 (N_1011,N_904,N_823);
nand U1012 (N_1012,N_937,N_456);
and U1013 (N_1013,N_855,N_570);
nor U1014 (N_1014,N_387,N_717);
and U1015 (N_1015,N_772,N_687);
nand U1016 (N_1016,N_417,N_513);
nor U1017 (N_1017,N_312,N_956);
nand U1018 (N_1018,N_260,N_645);
nor U1019 (N_1019,N_34,N_712);
nor U1020 (N_1020,N_669,N_868);
and U1021 (N_1021,N_444,N_6);
or U1022 (N_1022,N_472,N_196);
or U1023 (N_1023,N_147,N_854);
or U1024 (N_1024,N_507,N_75);
nor U1025 (N_1025,N_942,N_198);
nor U1026 (N_1026,N_627,N_109);
or U1027 (N_1027,N_266,N_479);
or U1028 (N_1028,N_858,N_382);
nor U1029 (N_1029,N_683,N_670);
nand U1030 (N_1030,N_602,N_174);
nor U1031 (N_1031,N_53,N_822);
nor U1032 (N_1032,N_424,N_771);
or U1033 (N_1033,N_103,N_0);
and U1034 (N_1034,N_769,N_230);
nand U1035 (N_1035,N_265,N_613);
nor U1036 (N_1036,N_969,N_350);
or U1037 (N_1037,N_125,N_962);
nor U1038 (N_1038,N_947,N_519);
nand U1039 (N_1039,N_517,N_463);
and U1040 (N_1040,N_970,N_142);
and U1041 (N_1041,N_911,N_963);
and U1042 (N_1042,N_764,N_921);
or U1043 (N_1043,N_723,N_191);
nor U1044 (N_1044,N_274,N_425);
and U1045 (N_1045,N_55,N_696);
nand U1046 (N_1046,N_497,N_841);
and U1047 (N_1047,N_359,N_280);
and U1048 (N_1048,N_17,N_888);
or U1049 (N_1049,N_214,N_227);
and U1050 (N_1050,N_657,N_83);
and U1051 (N_1051,N_704,N_930);
or U1052 (N_1052,N_975,N_892);
or U1053 (N_1053,N_659,N_887);
or U1054 (N_1054,N_621,N_572);
or U1055 (N_1055,N_524,N_453);
and U1056 (N_1056,N_495,N_189);
or U1057 (N_1057,N_640,N_84);
nand U1058 (N_1058,N_733,N_418);
nand U1059 (N_1059,N_158,N_656);
nor U1060 (N_1060,N_991,N_779);
nand U1061 (N_1061,N_556,N_340);
nand U1062 (N_1062,N_716,N_59);
or U1063 (N_1063,N_20,N_420);
nand U1064 (N_1064,N_817,N_306);
nand U1065 (N_1065,N_315,N_363);
nor U1066 (N_1066,N_408,N_334);
or U1067 (N_1067,N_619,N_541);
and U1068 (N_1068,N_743,N_511);
and U1069 (N_1069,N_554,N_152);
and U1070 (N_1070,N_238,N_532);
and U1071 (N_1071,N_200,N_70);
and U1072 (N_1072,N_967,N_338);
nor U1073 (N_1073,N_12,N_161);
or U1074 (N_1074,N_215,N_212);
and U1075 (N_1075,N_972,N_201);
or U1076 (N_1076,N_940,N_86);
nand U1077 (N_1077,N_71,N_959);
nor U1078 (N_1078,N_977,N_600);
nand U1079 (N_1079,N_432,N_992);
or U1080 (N_1080,N_430,N_692);
or U1081 (N_1081,N_129,N_759);
and U1082 (N_1082,N_375,N_611);
and U1083 (N_1083,N_643,N_121);
nand U1084 (N_1084,N_286,N_440);
nor U1085 (N_1085,N_435,N_477);
nand U1086 (N_1086,N_585,N_861);
nor U1087 (N_1087,N_285,N_148);
nand U1088 (N_1088,N_303,N_933);
and U1089 (N_1089,N_1,N_879);
and U1090 (N_1090,N_410,N_51);
nor U1091 (N_1091,N_800,N_849);
nand U1092 (N_1092,N_386,N_481);
nor U1093 (N_1093,N_976,N_445);
nor U1094 (N_1094,N_377,N_442);
or U1095 (N_1095,N_92,N_316);
nand U1096 (N_1096,N_753,N_912);
nand U1097 (N_1097,N_691,N_458);
nand U1098 (N_1098,N_313,N_354);
nand U1099 (N_1099,N_528,N_885);
and U1100 (N_1100,N_379,N_837);
nand U1101 (N_1101,N_383,N_981);
nand U1102 (N_1102,N_851,N_647);
nand U1103 (N_1103,N_796,N_546);
or U1104 (N_1104,N_918,N_697);
or U1105 (N_1105,N_839,N_80);
or U1106 (N_1106,N_913,N_179);
and U1107 (N_1107,N_317,N_391);
and U1108 (N_1108,N_182,N_811);
and U1109 (N_1109,N_90,N_865);
nand U1110 (N_1110,N_795,N_628);
and U1111 (N_1111,N_690,N_655);
nor U1112 (N_1112,N_449,N_762);
or U1113 (N_1113,N_884,N_203);
xnor U1114 (N_1114,N_906,N_510);
nor U1115 (N_1115,N_738,N_231);
nand U1116 (N_1116,N_798,N_832);
and U1117 (N_1117,N_701,N_140);
nor U1118 (N_1118,N_237,N_816);
and U1119 (N_1119,N_686,N_380);
and U1120 (N_1120,N_407,N_873);
nand U1121 (N_1121,N_422,N_480);
nor U1122 (N_1122,N_256,N_708);
or U1123 (N_1123,N_351,N_789);
and U1124 (N_1124,N_111,N_715);
nor U1125 (N_1125,N_565,N_150);
and U1126 (N_1126,N_490,N_136);
nand U1127 (N_1127,N_939,N_289);
or U1128 (N_1128,N_803,N_15);
nand U1129 (N_1129,N_986,N_642);
nand U1130 (N_1130,N_396,N_287);
or U1131 (N_1131,N_979,N_130);
and U1132 (N_1132,N_877,N_676);
nand U1133 (N_1133,N_801,N_909);
nor U1134 (N_1134,N_763,N_91);
nand U1135 (N_1135,N_277,N_199);
nand U1136 (N_1136,N_624,N_551);
or U1137 (N_1137,N_902,N_830);
or U1138 (N_1138,N_290,N_580);
or U1139 (N_1139,N_443,N_649);
nor U1140 (N_1140,N_100,N_677);
or U1141 (N_1141,N_587,N_333);
xor U1142 (N_1142,N_702,N_890);
nor U1143 (N_1143,N_331,N_998);
nand U1144 (N_1144,N_573,N_505);
nand U1145 (N_1145,N_438,N_133);
and U1146 (N_1146,N_362,N_36);
nand U1147 (N_1147,N_745,N_127);
or U1148 (N_1148,N_104,N_465);
nand U1149 (N_1149,N_767,N_31);
nand U1150 (N_1150,N_826,N_297);
or U1151 (N_1151,N_709,N_93);
and U1152 (N_1152,N_978,N_67);
nand U1153 (N_1153,N_328,N_689);
nand U1154 (N_1154,N_819,N_559);
or U1155 (N_1155,N_654,N_557);
nand U1156 (N_1156,N_954,N_705);
and U1157 (N_1157,N_255,N_840);
and U1158 (N_1158,N_482,N_920);
or U1159 (N_1159,N_989,N_378);
or U1160 (N_1160,N_469,N_343);
nand U1161 (N_1161,N_175,N_239);
nand U1162 (N_1162,N_48,N_700);
and U1163 (N_1163,N_758,N_97);
or U1164 (N_1164,N_739,N_321);
or U1165 (N_1165,N_827,N_953);
or U1166 (N_1166,N_590,N_935);
nor U1167 (N_1167,N_539,N_852);
nand U1168 (N_1168,N_373,N_208);
and U1169 (N_1169,N_352,N_60);
or U1170 (N_1170,N_644,N_155);
nand U1171 (N_1171,N_115,N_648);
nand U1172 (N_1172,N_320,N_123);
or U1173 (N_1173,N_264,N_102);
nor U1174 (N_1174,N_732,N_188);
or U1175 (N_1175,N_89,N_671);
and U1176 (N_1176,N_951,N_825);
and U1177 (N_1177,N_542,N_908);
nor U1178 (N_1178,N_845,N_869);
or U1179 (N_1179,N_411,N_398);
or U1180 (N_1180,N_901,N_294);
nand U1181 (N_1181,N_730,N_184);
and U1182 (N_1182,N_850,N_974);
or U1183 (N_1183,N_368,N_522);
or U1184 (N_1184,N_578,N_774);
and U1185 (N_1185,N_964,N_18);
nand U1186 (N_1186,N_982,N_842);
nand U1187 (N_1187,N_710,N_462);
nor U1188 (N_1188,N_925,N_405);
or U1189 (N_1189,N_612,N_952);
nand U1190 (N_1190,N_126,N_240);
and U1191 (N_1191,N_518,N_857);
and U1192 (N_1192,N_157,N_646);
nand U1193 (N_1193,N_735,N_33);
and U1194 (N_1194,N_948,N_38);
and U1195 (N_1195,N_170,N_786);
nand U1196 (N_1196,N_564,N_509);
and U1197 (N_1197,N_630,N_193);
nor U1198 (N_1198,N_584,N_162);
nor U1199 (N_1199,N_186,N_69);
or U1200 (N_1200,N_698,N_566);
nand U1201 (N_1201,N_299,N_665);
nand U1202 (N_1202,N_381,N_178);
nand U1203 (N_1203,N_545,N_454);
and U1204 (N_1204,N_897,N_523);
nor U1205 (N_1205,N_82,N_750);
or U1206 (N_1206,N_117,N_813);
and U1207 (N_1207,N_356,N_579);
or U1208 (N_1208,N_838,N_537);
nor U1209 (N_1209,N_599,N_258);
or U1210 (N_1210,N_429,N_618);
nor U1211 (N_1211,N_428,N_997);
nand U1212 (N_1212,N_987,N_291);
nand U1213 (N_1213,N_747,N_775);
nor U1214 (N_1214,N_348,N_641);
nand U1215 (N_1215,N_29,N_607);
xor U1216 (N_1216,N_335,N_263);
nand U1217 (N_1217,N_250,N_344);
and U1218 (N_1218,N_202,N_792);
nor U1219 (N_1219,N_606,N_326);
and U1220 (N_1220,N_146,N_714);
and U1221 (N_1221,N_931,N_304);
nor U1222 (N_1222,N_168,N_608);
nor U1223 (N_1223,N_965,N_390);
nor U1224 (N_1224,N_864,N_151);
nand U1225 (N_1225,N_577,N_110);
and U1226 (N_1226,N_980,N_504);
and U1227 (N_1227,N_571,N_544);
or U1228 (N_1228,N_720,N_828);
nand U1229 (N_1229,N_112,N_156);
nor U1230 (N_1230,N_63,N_601);
nand U1231 (N_1231,N_558,N_369);
nand U1232 (N_1232,N_399,N_164);
or U1233 (N_1233,N_549,N_28);
nor U1234 (N_1234,N_216,N_211);
nor U1235 (N_1235,N_5,N_736);
nor U1236 (N_1236,N_583,N_222);
or U1237 (N_1237,N_985,N_76);
nand U1238 (N_1238,N_724,N_388);
or U1239 (N_1239,N_251,N_706);
nor U1240 (N_1240,N_574,N_693);
and U1241 (N_1241,N_791,N_744);
nor U1242 (N_1242,N_961,N_530);
and U1243 (N_1243,N_740,N_153);
nand U1244 (N_1244,N_85,N_971);
or U1245 (N_1245,N_722,N_248);
nor U1246 (N_1246,N_468,N_397);
nor U1247 (N_1247,N_922,N_787);
and U1248 (N_1248,N_596,N_298);
nand U1249 (N_1249,N_903,N_984);
nand U1250 (N_1250,N_353,N_149);
nand U1251 (N_1251,N_875,N_415);
or U1252 (N_1252,N_225,N_489);
and U1253 (N_1253,N_794,N_536);
or U1254 (N_1254,N_144,N_821);
nand U1255 (N_1255,N_124,N_760);
nor U1256 (N_1256,N_259,N_543);
and U1257 (N_1257,N_50,N_272);
and U1258 (N_1258,N_421,N_664);
and U1259 (N_1259,N_808,N_412);
nand U1260 (N_1260,N_404,N_72);
or U1261 (N_1261,N_361,N_302);
nor U1262 (N_1262,N_177,N_941);
or U1263 (N_1263,N_946,N_651);
nor U1264 (N_1264,N_242,N_355);
or U1265 (N_1265,N_820,N_731);
nor U1266 (N_1266,N_400,N_11);
nor U1267 (N_1267,N_135,N_322);
or U1268 (N_1268,N_847,N_553);
nand U1269 (N_1269,N_521,N_673);
nor U1270 (N_1270,N_217,N_834);
nand U1271 (N_1271,N_662,N_950);
nand U1272 (N_1272,N_436,N_923);
nor U1273 (N_1273,N_282,N_815);
nor U1274 (N_1274,N_278,N_32);
nor U1275 (N_1275,N_721,N_23);
and U1276 (N_1276,N_450,N_540);
nor U1277 (N_1277,N_484,N_765);
nor U1278 (N_1278,N_171,N_681);
or U1279 (N_1279,N_195,N_737);
or U1280 (N_1280,N_853,N_209);
nand U1281 (N_1281,N_276,N_128);
and U1282 (N_1282,N_94,N_741);
nand U1283 (N_1283,N_515,N_314);
or U1284 (N_1284,N_52,N_488);
nand U1285 (N_1285,N_748,N_205);
nor U1286 (N_1286,N_384,N_812);
or U1287 (N_1287,N_228,N_672);
nand U1288 (N_1288,N_439,N_99);
and U1289 (N_1289,N_269,N_414);
nor U1290 (N_1290,N_249,N_635);
nand U1291 (N_1291,N_860,N_183);
and U1292 (N_1292,N_374,N_30);
or U1293 (N_1293,N_141,N_896);
nand U1294 (N_1294,N_863,N_403);
nand U1295 (N_1295,N_360,N_300);
nand U1296 (N_1296,N_273,N_21);
or U1297 (N_1297,N_675,N_219);
or U1298 (N_1298,N_43,N_13);
and U1299 (N_1299,N_999,N_653);
nor U1300 (N_1300,N_27,N_19);
and U1301 (N_1301,N_527,N_496);
or U1302 (N_1302,N_270,N_756);
and U1303 (N_1303,N_433,N_726);
and U1304 (N_1304,N_491,N_471);
xnor U1305 (N_1305,N_207,N_871);
or U1306 (N_1306,N_336,N_770);
or U1307 (N_1307,N_292,N_402);
nand U1308 (N_1308,N_729,N_325);
nand U1309 (N_1309,N_636,N_218);
nor U1310 (N_1310,N_134,N_241);
nand U1311 (N_1311,N_244,N_16);
xor U1312 (N_1312,N_392,N_475);
nor U1313 (N_1313,N_810,N_79);
or U1314 (N_1314,N_995,N_169);
nor U1315 (N_1315,N_45,N_595);
nor U1316 (N_1316,N_473,N_327);
and U1317 (N_1317,N_910,N_660);
or U1318 (N_1318,N_878,N_234);
nor U1319 (N_1319,N_78,N_512);
nor U1320 (N_1320,N_894,N_154);
nor U1321 (N_1321,N_223,N_685);
nor U1322 (N_1322,N_460,N_139);
nor U1323 (N_1323,N_591,N_889);
nor U1324 (N_1324,N_167,N_550);
nor U1325 (N_1325,N_876,N_113);
and U1326 (N_1326,N_781,N_98);
and U1327 (N_1327,N_552,N_968);
nand U1328 (N_1328,N_874,N_220);
and U1329 (N_1329,N_594,N_926);
nand U1330 (N_1330,N_680,N_395);
and U1331 (N_1331,N_917,N_684);
or U1332 (N_1332,N_859,N_65);
xor U1333 (N_1333,N_275,N_499);
nand U1334 (N_1334,N_245,N_132);
nand U1335 (N_1335,N_2,N_243);
and U1336 (N_1336,N_58,N_301);
nor U1337 (N_1337,N_500,N_597);
or U1338 (N_1338,N_609,N_347);
nand U1339 (N_1339,N_163,N_486);
nand U1340 (N_1340,N_634,N_831);
nand U1341 (N_1341,N_49,N_576);
nand U1342 (N_1342,N_131,N_994);
and U1343 (N_1343,N_806,N_824);
nor U1344 (N_1344,N_73,N_725);
and U1345 (N_1345,N_87,N_24);
and U1346 (N_1346,N_213,N_915);
and U1347 (N_1347,N_802,N_966);
nor U1348 (N_1348,N_41,N_844);
nand U1349 (N_1349,N_604,N_120);
nand U1350 (N_1350,N_589,N_26);
nand U1351 (N_1351,N_711,N_626);
nand U1352 (N_1352,N_284,N_105);
nand U1353 (N_1353,N_508,N_311);
or U1354 (N_1354,N_784,N_40);
nor U1355 (N_1355,N_814,N_797);
nor U1356 (N_1356,N_310,N_254);
nor U1357 (N_1357,N_780,N_62);
nor U1358 (N_1358,N_835,N_502);
nand U1359 (N_1359,N_881,N_159);
nand U1360 (N_1360,N_166,N_569);
or U1361 (N_1361,N_533,N_592);
nor U1362 (N_1362,N_101,N_916);
nand U1363 (N_1363,N_307,N_341);
or U1364 (N_1364,N_777,N_474);
and U1365 (N_1365,N_682,N_487);
nand U1366 (N_1366,N_498,N_703);
nor U1367 (N_1367,N_520,N_788);
or U1368 (N_1368,N_883,N_927);
nand U1369 (N_1369,N_668,N_192);
nand U1370 (N_1370,N_437,N_932);
nor U1371 (N_1371,N_357,N_617);
nand U1372 (N_1372,N_406,N_66);
and U1373 (N_1373,N_547,N_581);
nand U1374 (N_1374,N_160,N_534);
and U1375 (N_1375,N_293,N_247);
nor U1376 (N_1376,N_843,N_81);
and U1377 (N_1377,N_658,N_623);
nor U1378 (N_1378,N_394,N_434);
nand U1379 (N_1379,N_663,N_281);
nor U1380 (N_1380,N_993,N_799);
nor U1381 (N_1381,N_616,N_560);
nand U1382 (N_1382,N_983,N_856);
nand U1383 (N_1383,N_538,N_516);
or U1384 (N_1384,N_919,N_924);
or U1385 (N_1385,N_77,N_719);
nor U1386 (N_1386,N_620,N_452);
nor U1387 (N_1387,N_324,N_431);
nor U1388 (N_1388,N_9,N_426);
and U1389 (N_1389,N_185,N_204);
or U1390 (N_1390,N_253,N_562);
or U1391 (N_1391,N_943,N_905);
nor U1392 (N_1392,N_667,N_308);
nor U1393 (N_1393,N_470,N_914);
xor U1394 (N_1394,N_389,N_106);
or U1395 (N_1395,N_413,N_37);
or U1396 (N_1396,N_305,N_68);
nand U1397 (N_1397,N_337,N_900);
or U1398 (N_1398,N_107,N_323);
nor U1399 (N_1399,N_661,N_805);
nand U1400 (N_1400,N_46,N_329);
nand U1401 (N_1401,N_793,N_118);
or U1402 (N_1402,N_61,N_768);
nor U1403 (N_1403,N_531,N_678);
and U1404 (N_1404,N_370,N_393);
nor U1405 (N_1405,N_476,N_448);
and U1406 (N_1406,N_776,N_749);
or U1407 (N_1407,N_346,N_688);
nand U1408 (N_1408,N_575,N_514);
nand U1409 (N_1409,N_694,N_74);
or U1410 (N_1410,N_582,N_427);
or U1411 (N_1411,N_232,N_752);
and U1412 (N_1412,N_833,N_330);
nor U1413 (N_1413,N_928,N_734);
nand U1414 (N_1414,N_371,N_862);
nor U1415 (N_1415,N_455,N_419);
nand U1416 (N_1416,N_973,N_267);
nor U1417 (N_1417,N_358,N_116);
or U1418 (N_1418,N_467,N_934);
and U1419 (N_1419,N_446,N_54);
nor U1420 (N_1420,N_345,N_907);
nand U1421 (N_1421,N_235,N_886);
nor U1422 (N_1422,N_296,N_773);
nor U1423 (N_1423,N_367,N_631);
nand U1424 (N_1424,N_493,N_197);
nand U1425 (N_1425,N_880,N_181);
nand U1426 (N_1426,N_790,N_464);
nand U1427 (N_1427,N_990,N_746);
nand U1428 (N_1428,N_409,N_526);
nor U1429 (N_1429,N_441,N_638);
or U1430 (N_1430,N_893,N_818);
or U1431 (N_1431,N_870,N_588);
and U1432 (N_1432,N_180,N_271);
or U1433 (N_1433,N_751,N_761);
nor U1434 (N_1434,N_25,N_246);
nand U1435 (N_1435,N_283,N_728);
nor U1436 (N_1436,N_137,N_996);
and U1437 (N_1437,N_332,N_364);
nor U1438 (N_1438,N_561,N_755);
nor U1439 (N_1439,N_57,N_176);
nand U1440 (N_1440,N_461,N_957);
and U1441 (N_1441,N_944,N_342);
and U1442 (N_1442,N_349,N_108);
nor U1443 (N_1443,N_194,N_309);
nand U1444 (N_1444,N_757,N_742);
and U1445 (N_1445,N_206,N_506);
and U1446 (N_1446,N_233,N_936);
nor U1447 (N_1447,N_882,N_958);
nand U1448 (N_1448,N_548,N_718);
xor U1449 (N_1449,N_42,N_891);
nor U1450 (N_1450,N_633,N_567);
nor U1451 (N_1451,N_494,N_713);
nand U1452 (N_1452,N_114,N_423);
nand U1453 (N_1453,N_319,N_88);
or U1454 (N_1454,N_848,N_938);
or U1455 (N_1455,N_372,N_376);
nand U1456 (N_1456,N_754,N_598);
nand U1457 (N_1457,N_945,N_836);
nor U1458 (N_1458,N_318,N_252);
nor U1459 (N_1459,N_172,N_563);
and U1460 (N_1460,N_679,N_190);
nand U1461 (N_1461,N_695,N_727);
and U1462 (N_1462,N_898,N_529);
and U1463 (N_1463,N_666,N_22);
nand U1464 (N_1464,N_95,N_39);
nand U1465 (N_1465,N_366,N_288);
nor U1466 (N_1466,N_143,N_778);
and U1467 (N_1467,N_614,N_122);
nor U1468 (N_1468,N_14,N_785);
nand U1469 (N_1469,N_960,N_629);
nand U1470 (N_1470,N_236,N_47);
and U1471 (N_1471,N_96,N_622);
nand U1472 (N_1472,N_809,N_929);
or U1473 (N_1473,N_459,N_485);
and U1474 (N_1474,N_525,N_257);
nand U1475 (N_1475,N_365,N_949);
nand U1476 (N_1476,N_138,N_899);
nor U1477 (N_1477,N_501,N_173);
nor U1478 (N_1478,N_279,N_483);
and U1479 (N_1479,N_262,N_625);
nor U1480 (N_1480,N_535,N_639);
and U1481 (N_1481,N_650,N_895);
nand U1482 (N_1482,N_226,N_637);
xnor U1483 (N_1483,N_652,N_210);
nor U1484 (N_1484,N_447,N_35);
and U1485 (N_1485,N_866,N_988);
nor U1486 (N_1486,N_145,N_804);
nand U1487 (N_1487,N_466,N_846);
or U1488 (N_1488,N_44,N_229);
and U1489 (N_1489,N_503,N_3);
and U1490 (N_1490,N_10,N_64);
and U1491 (N_1491,N_416,N_807);
and U1492 (N_1492,N_782,N_492);
nand U1493 (N_1493,N_187,N_632);
or U1494 (N_1494,N_955,N_339);
and U1495 (N_1495,N_224,N_783);
nand U1496 (N_1496,N_8,N_867);
or U1497 (N_1497,N_119,N_457);
and U1498 (N_1498,N_385,N_674);
and U1499 (N_1499,N_615,N_56);
nor U1500 (N_1500,N_771,N_631);
nand U1501 (N_1501,N_367,N_185);
nand U1502 (N_1502,N_341,N_247);
and U1503 (N_1503,N_177,N_615);
and U1504 (N_1504,N_847,N_438);
nand U1505 (N_1505,N_948,N_657);
and U1506 (N_1506,N_950,N_493);
nor U1507 (N_1507,N_224,N_280);
and U1508 (N_1508,N_247,N_766);
or U1509 (N_1509,N_167,N_596);
nand U1510 (N_1510,N_370,N_466);
or U1511 (N_1511,N_998,N_412);
nand U1512 (N_1512,N_306,N_315);
or U1513 (N_1513,N_371,N_805);
and U1514 (N_1514,N_396,N_84);
or U1515 (N_1515,N_223,N_473);
nor U1516 (N_1516,N_71,N_533);
nor U1517 (N_1517,N_267,N_825);
nand U1518 (N_1518,N_894,N_782);
and U1519 (N_1519,N_867,N_844);
and U1520 (N_1520,N_456,N_733);
or U1521 (N_1521,N_501,N_991);
and U1522 (N_1522,N_543,N_317);
nand U1523 (N_1523,N_666,N_423);
nand U1524 (N_1524,N_953,N_293);
nor U1525 (N_1525,N_767,N_491);
nor U1526 (N_1526,N_977,N_996);
and U1527 (N_1527,N_262,N_793);
nor U1528 (N_1528,N_463,N_553);
nand U1529 (N_1529,N_329,N_638);
and U1530 (N_1530,N_571,N_244);
and U1531 (N_1531,N_46,N_867);
and U1532 (N_1532,N_191,N_662);
nand U1533 (N_1533,N_448,N_509);
nor U1534 (N_1534,N_867,N_462);
nor U1535 (N_1535,N_203,N_579);
nand U1536 (N_1536,N_325,N_480);
nor U1537 (N_1537,N_976,N_189);
and U1538 (N_1538,N_983,N_375);
nor U1539 (N_1539,N_772,N_303);
or U1540 (N_1540,N_460,N_283);
nor U1541 (N_1541,N_23,N_698);
nor U1542 (N_1542,N_44,N_450);
nand U1543 (N_1543,N_423,N_785);
nand U1544 (N_1544,N_658,N_699);
and U1545 (N_1545,N_592,N_850);
nor U1546 (N_1546,N_461,N_40);
nand U1547 (N_1547,N_778,N_655);
nand U1548 (N_1548,N_410,N_195);
or U1549 (N_1549,N_120,N_719);
nand U1550 (N_1550,N_829,N_563);
or U1551 (N_1551,N_589,N_387);
or U1552 (N_1552,N_632,N_732);
nor U1553 (N_1553,N_825,N_780);
nor U1554 (N_1554,N_347,N_258);
and U1555 (N_1555,N_207,N_834);
and U1556 (N_1556,N_44,N_40);
and U1557 (N_1557,N_175,N_70);
nand U1558 (N_1558,N_344,N_309);
or U1559 (N_1559,N_685,N_88);
nor U1560 (N_1560,N_333,N_167);
nand U1561 (N_1561,N_344,N_130);
nor U1562 (N_1562,N_345,N_980);
nor U1563 (N_1563,N_439,N_761);
nand U1564 (N_1564,N_295,N_399);
nor U1565 (N_1565,N_561,N_427);
and U1566 (N_1566,N_730,N_359);
or U1567 (N_1567,N_776,N_82);
nand U1568 (N_1568,N_878,N_383);
and U1569 (N_1569,N_331,N_906);
and U1570 (N_1570,N_330,N_144);
and U1571 (N_1571,N_509,N_270);
or U1572 (N_1572,N_203,N_260);
nor U1573 (N_1573,N_41,N_8);
nor U1574 (N_1574,N_559,N_993);
or U1575 (N_1575,N_811,N_539);
or U1576 (N_1576,N_755,N_67);
nand U1577 (N_1577,N_484,N_327);
and U1578 (N_1578,N_366,N_755);
nor U1579 (N_1579,N_155,N_160);
nor U1580 (N_1580,N_726,N_920);
nand U1581 (N_1581,N_672,N_121);
nor U1582 (N_1582,N_278,N_187);
or U1583 (N_1583,N_990,N_103);
nor U1584 (N_1584,N_885,N_477);
nor U1585 (N_1585,N_808,N_205);
xnor U1586 (N_1586,N_787,N_401);
and U1587 (N_1587,N_176,N_390);
and U1588 (N_1588,N_293,N_193);
nor U1589 (N_1589,N_991,N_545);
and U1590 (N_1590,N_151,N_449);
and U1591 (N_1591,N_688,N_315);
and U1592 (N_1592,N_856,N_752);
or U1593 (N_1593,N_402,N_577);
and U1594 (N_1594,N_877,N_650);
nand U1595 (N_1595,N_316,N_356);
nor U1596 (N_1596,N_855,N_652);
nor U1597 (N_1597,N_400,N_27);
or U1598 (N_1598,N_478,N_713);
and U1599 (N_1599,N_941,N_185);
nor U1600 (N_1600,N_719,N_747);
and U1601 (N_1601,N_882,N_557);
nand U1602 (N_1602,N_809,N_465);
nand U1603 (N_1603,N_43,N_116);
nor U1604 (N_1604,N_326,N_173);
xor U1605 (N_1605,N_335,N_234);
nor U1606 (N_1606,N_907,N_17);
or U1607 (N_1607,N_478,N_916);
or U1608 (N_1608,N_121,N_269);
nand U1609 (N_1609,N_824,N_686);
xor U1610 (N_1610,N_758,N_5);
or U1611 (N_1611,N_537,N_915);
or U1612 (N_1612,N_271,N_109);
nor U1613 (N_1613,N_743,N_116);
and U1614 (N_1614,N_481,N_40);
nand U1615 (N_1615,N_888,N_325);
or U1616 (N_1616,N_131,N_48);
or U1617 (N_1617,N_723,N_860);
nor U1618 (N_1618,N_969,N_616);
nor U1619 (N_1619,N_172,N_51);
and U1620 (N_1620,N_939,N_378);
nand U1621 (N_1621,N_700,N_704);
nor U1622 (N_1622,N_673,N_881);
or U1623 (N_1623,N_936,N_962);
nand U1624 (N_1624,N_224,N_447);
and U1625 (N_1625,N_551,N_774);
or U1626 (N_1626,N_586,N_3);
or U1627 (N_1627,N_890,N_664);
nor U1628 (N_1628,N_822,N_918);
nor U1629 (N_1629,N_568,N_915);
nor U1630 (N_1630,N_1,N_140);
nand U1631 (N_1631,N_882,N_413);
and U1632 (N_1632,N_516,N_361);
nand U1633 (N_1633,N_574,N_75);
and U1634 (N_1634,N_834,N_887);
or U1635 (N_1635,N_137,N_813);
nor U1636 (N_1636,N_177,N_709);
and U1637 (N_1637,N_138,N_227);
and U1638 (N_1638,N_535,N_206);
and U1639 (N_1639,N_563,N_24);
and U1640 (N_1640,N_157,N_350);
nand U1641 (N_1641,N_554,N_580);
and U1642 (N_1642,N_135,N_659);
nor U1643 (N_1643,N_586,N_492);
and U1644 (N_1644,N_246,N_157);
nand U1645 (N_1645,N_922,N_203);
or U1646 (N_1646,N_204,N_980);
nand U1647 (N_1647,N_969,N_935);
nand U1648 (N_1648,N_317,N_998);
nand U1649 (N_1649,N_946,N_71);
and U1650 (N_1650,N_575,N_779);
and U1651 (N_1651,N_255,N_766);
nand U1652 (N_1652,N_345,N_401);
and U1653 (N_1653,N_581,N_726);
nand U1654 (N_1654,N_15,N_150);
and U1655 (N_1655,N_7,N_892);
nand U1656 (N_1656,N_258,N_647);
nand U1657 (N_1657,N_542,N_497);
or U1658 (N_1658,N_602,N_502);
nor U1659 (N_1659,N_577,N_476);
and U1660 (N_1660,N_853,N_354);
and U1661 (N_1661,N_522,N_872);
and U1662 (N_1662,N_903,N_250);
nand U1663 (N_1663,N_512,N_956);
nand U1664 (N_1664,N_486,N_157);
and U1665 (N_1665,N_6,N_479);
and U1666 (N_1666,N_852,N_870);
nand U1667 (N_1667,N_194,N_305);
nand U1668 (N_1668,N_699,N_453);
and U1669 (N_1669,N_491,N_536);
nand U1670 (N_1670,N_3,N_455);
nor U1671 (N_1671,N_258,N_995);
or U1672 (N_1672,N_202,N_366);
and U1673 (N_1673,N_806,N_766);
nor U1674 (N_1674,N_713,N_551);
or U1675 (N_1675,N_102,N_477);
and U1676 (N_1676,N_45,N_29);
nand U1677 (N_1677,N_209,N_76);
and U1678 (N_1678,N_996,N_767);
and U1679 (N_1679,N_424,N_825);
nor U1680 (N_1680,N_143,N_75);
and U1681 (N_1681,N_354,N_584);
nor U1682 (N_1682,N_524,N_273);
nand U1683 (N_1683,N_708,N_340);
nor U1684 (N_1684,N_961,N_540);
or U1685 (N_1685,N_276,N_683);
nor U1686 (N_1686,N_590,N_112);
or U1687 (N_1687,N_132,N_823);
and U1688 (N_1688,N_821,N_415);
or U1689 (N_1689,N_22,N_837);
nand U1690 (N_1690,N_243,N_129);
and U1691 (N_1691,N_315,N_23);
nor U1692 (N_1692,N_315,N_241);
nand U1693 (N_1693,N_831,N_904);
nor U1694 (N_1694,N_588,N_339);
and U1695 (N_1695,N_768,N_826);
nand U1696 (N_1696,N_64,N_251);
or U1697 (N_1697,N_126,N_844);
and U1698 (N_1698,N_14,N_611);
nand U1699 (N_1699,N_570,N_812);
and U1700 (N_1700,N_578,N_728);
or U1701 (N_1701,N_189,N_211);
nand U1702 (N_1702,N_4,N_649);
and U1703 (N_1703,N_938,N_160);
nand U1704 (N_1704,N_157,N_346);
and U1705 (N_1705,N_886,N_106);
nand U1706 (N_1706,N_345,N_951);
or U1707 (N_1707,N_836,N_735);
nor U1708 (N_1708,N_265,N_323);
nor U1709 (N_1709,N_719,N_565);
nand U1710 (N_1710,N_281,N_841);
nand U1711 (N_1711,N_672,N_929);
or U1712 (N_1712,N_532,N_542);
nor U1713 (N_1713,N_529,N_849);
nand U1714 (N_1714,N_93,N_844);
nand U1715 (N_1715,N_857,N_563);
nand U1716 (N_1716,N_552,N_929);
or U1717 (N_1717,N_4,N_13);
nor U1718 (N_1718,N_728,N_241);
and U1719 (N_1719,N_360,N_729);
nand U1720 (N_1720,N_110,N_346);
nand U1721 (N_1721,N_13,N_805);
or U1722 (N_1722,N_121,N_827);
nand U1723 (N_1723,N_918,N_153);
or U1724 (N_1724,N_886,N_523);
nand U1725 (N_1725,N_12,N_643);
or U1726 (N_1726,N_266,N_670);
or U1727 (N_1727,N_733,N_887);
nand U1728 (N_1728,N_926,N_837);
or U1729 (N_1729,N_586,N_102);
nand U1730 (N_1730,N_874,N_376);
and U1731 (N_1731,N_638,N_832);
and U1732 (N_1732,N_582,N_543);
nor U1733 (N_1733,N_772,N_76);
nand U1734 (N_1734,N_918,N_885);
nand U1735 (N_1735,N_543,N_70);
or U1736 (N_1736,N_775,N_412);
or U1737 (N_1737,N_631,N_803);
or U1738 (N_1738,N_938,N_344);
or U1739 (N_1739,N_48,N_339);
nand U1740 (N_1740,N_680,N_327);
or U1741 (N_1741,N_748,N_231);
or U1742 (N_1742,N_450,N_914);
or U1743 (N_1743,N_65,N_958);
nand U1744 (N_1744,N_377,N_300);
or U1745 (N_1745,N_72,N_957);
nand U1746 (N_1746,N_388,N_318);
nor U1747 (N_1747,N_904,N_957);
or U1748 (N_1748,N_199,N_497);
nor U1749 (N_1749,N_234,N_333);
or U1750 (N_1750,N_560,N_257);
nor U1751 (N_1751,N_634,N_952);
or U1752 (N_1752,N_374,N_712);
or U1753 (N_1753,N_323,N_57);
nand U1754 (N_1754,N_815,N_792);
or U1755 (N_1755,N_284,N_739);
nand U1756 (N_1756,N_895,N_682);
or U1757 (N_1757,N_859,N_320);
nand U1758 (N_1758,N_948,N_62);
or U1759 (N_1759,N_11,N_654);
nand U1760 (N_1760,N_720,N_952);
or U1761 (N_1761,N_370,N_519);
and U1762 (N_1762,N_209,N_602);
nor U1763 (N_1763,N_38,N_105);
xor U1764 (N_1764,N_278,N_608);
or U1765 (N_1765,N_478,N_96);
or U1766 (N_1766,N_420,N_14);
nor U1767 (N_1767,N_170,N_908);
or U1768 (N_1768,N_136,N_776);
and U1769 (N_1769,N_28,N_790);
and U1770 (N_1770,N_963,N_478);
nor U1771 (N_1771,N_847,N_393);
and U1772 (N_1772,N_27,N_452);
or U1773 (N_1773,N_770,N_360);
or U1774 (N_1774,N_216,N_734);
or U1775 (N_1775,N_731,N_822);
or U1776 (N_1776,N_806,N_897);
and U1777 (N_1777,N_985,N_841);
and U1778 (N_1778,N_436,N_581);
or U1779 (N_1779,N_445,N_134);
or U1780 (N_1780,N_346,N_119);
nor U1781 (N_1781,N_613,N_120);
nor U1782 (N_1782,N_441,N_19);
nand U1783 (N_1783,N_497,N_753);
and U1784 (N_1784,N_31,N_296);
or U1785 (N_1785,N_901,N_742);
nor U1786 (N_1786,N_916,N_497);
or U1787 (N_1787,N_67,N_521);
and U1788 (N_1788,N_970,N_732);
or U1789 (N_1789,N_163,N_238);
or U1790 (N_1790,N_907,N_513);
nand U1791 (N_1791,N_729,N_688);
or U1792 (N_1792,N_492,N_914);
nor U1793 (N_1793,N_513,N_634);
or U1794 (N_1794,N_811,N_984);
nor U1795 (N_1795,N_879,N_722);
or U1796 (N_1796,N_634,N_297);
nand U1797 (N_1797,N_682,N_777);
and U1798 (N_1798,N_958,N_608);
and U1799 (N_1799,N_564,N_767);
and U1800 (N_1800,N_988,N_771);
nand U1801 (N_1801,N_485,N_364);
nor U1802 (N_1802,N_128,N_100);
or U1803 (N_1803,N_914,N_861);
and U1804 (N_1804,N_143,N_198);
nand U1805 (N_1805,N_811,N_524);
and U1806 (N_1806,N_993,N_828);
nand U1807 (N_1807,N_44,N_213);
nand U1808 (N_1808,N_534,N_791);
or U1809 (N_1809,N_194,N_457);
nor U1810 (N_1810,N_562,N_593);
and U1811 (N_1811,N_594,N_916);
nor U1812 (N_1812,N_79,N_520);
and U1813 (N_1813,N_211,N_428);
and U1814 (N_1814,N_281,N_762);
nand U1815 (N_1815,N_144,N_437);
nand U1816 (N_1816,N_547,N_812);
nand U1817 (N_1817,N_475,N_447);
nand U1818 (N_1818,N_934,N_594);
nand U1819 (N_1819,N_946,N_377);
and U1820 (N_1820,N_99,N_614);
or U1821 (N_1821,N_166,N_466);
nor U1822 (N_1822,N_564,N_189);
or U1823 (N_1823,N_728,N_432);
and U1824 (N_1824,N_62,N_905);
and U1825 (N_1825,N_833,N_23);
nor U1826 (N_1826,N_395,N_70);
or U1827 (N_1827,N_508,N_140);
or U1828 (N_1828,N_253,N_933);
and U1829 (N_1829,N_270,N_440);
or U1830 (N_1830,N_40,N_135);
nand U1831 (N_1831,N_591,N_746);
nand U1832 (N_1832,N_151,N_730);
nand U1833 (N_1833,N_889,N_193);
or U1834 (N_1834,N_547,N_485);
nand U1835 (N_1835,N_846,N_103);
nand U1836 (N_1836,N_593,N_772);
or U1837 (N_1837,N_160,N_192);
and U1838 (N_1838,N_463,N_611);
nand U1839 (N_1839,N_582,N_314);
nand U1840 (N_1840,N_55,N_797);
nor U1841 (N_1841,N_844,N_359);
nand U1842 (N_1842,N_287,N_375);
or U1843 (N_1843,N_951,N_323);
nor U1844 (N_1844,N_352,N_10);
nand U1845 (N_1845,N_989,N_894);
nor U1846 (N_1846,N_135,N_831);
nand U1847 (N_1847,N_807,N_463);
nand U1848 (N_1848,N_861,N_876);
or U1849 (N_1849,N_133,N_491);
nor U1850 (N_1850,N_288,N_341);
nand U1851 (N_1851,N_907,N_996);
nor U1852 (N_1852,N_382,N_574);
nor U1853 (N_1853,N_492,N_975);
nor U1854 (N_1854,N_419,N_64);
or U1855 (N_1855,N_9,N_243);
nor U1856 (N_1856,N_39,N_424);
and U1857 (N_1857,N_290,N_407);
nand U1858 (N_1858,N_622,N_375);
nand U1859 (N_1859,N_926,N_176);
and U1860 (N_1860,N_322,N_779);
or U1861 (N_1861,N_297,N_864);
or U1862 (N_1862,N_283,N_190);
nor U1863 (N_1863,N_968,N_789);
or U1864 (N_1864,N_762,N_771);
or U1865 (N_1865,N_7,N_52);
and U1866 (N_1866,N_609,N_421);
nand U1867 (N_1867,N_803,N_110);
and U1868 (N_1868,N_177,N_855);
nor U1869 (N_1869,N_339,N_275);
or U1870 (N_1870,N_522,N_293);
nor U1871 (N_1871,N_993,N_75);
nor U1872 (N_1872,N_752,N_52);
nor U1873 (N_1873,N_744,N_837);
nor U1874 (N_1874,N_535,N_920);
nor U1875 (N_1875,N_370,N_974);
nor U1876 (N_1876,N_425,N_408);
or U1877 (N_1877,N_824,N_432);
and U1878 (N_1878,N_833,N_437);
nor U1879 (N_1879,N_787,N_597);
or U1880 (N_1880,N_877,N_189);
and U1881 (N_1881,N_183,N_766);
nand U1882 (N_1882,N_561,N_870);
and U1883 (N_1883,N_214,N_202);
nand U1884 (N_1884,N_153,N_603);
nor U1885 (N_1885,N_591,N_260);
and U1886 (N_1886,N_605,N_907);
or U1887 (N_1887,N_82,N_79);
and U1888 (N_1888,N_605,N_54);
and U1889 (N_1889,N_967,N_977);
nor U1890 (N_1890,N_298,N_259);
nor U1891 (N_1891,N_549,N_811);
nand U1892 (N_1892,N_517,N_817);
nor U1893 (N_1893,N_663,N_35);
or U1894 (N_1894,N_716,N_193);
or U1895 (N_1895,N_282,N_287);
nand U1896 (N_1896,N_880,N_404);
nor U1897 (N_1897,N_653,N_576);
nand U1898 (N_1898,N_220,N_861);
or U1899 (N_1899,N_650,N_804);
and U1900 (N_1900,N_668,N_441);
nor U1901 (N_1901,N_709,N_32);
nor U1902 (N_1902,N_394,N_329);
or U1903 (N_1903,N_137,N_805);
xor U1904 (N_1904,N_731,N_536);
or U1905 (N_1905,N_341,N_280);
nor U1906 (N_1906,N_518,N_321);
nand U1907 (N_1907,N_938,N_351);
nand U1908 (N_1908,N_855,N_179);
nor U1909 (N_1909,N_32,N_341);
nor U1910 (N_1910,N_250,N_366);
nor U1911 (N_1911,N_73,N_191);
nand U1912 (N_1912,N_29,N_755);
and U1913 (N_1913,N_62,N_789);
nand U1914 (N_1914,N_17,N_820);
nand U1915 (N_1915,N_52,N_718);
nor U1916 (N_1916,N_656,N_483);
nand U1917 (N_1917,N_165,N_240);
nand U1918 (N_1918,N_980,N_857);
or U1919 (N_1919,N_567,N_411);
and U1920 (N_1920,N_470,N_887);
or U1921 (N_1921,N_759,N_283);
or U1922 (N_1922,N_240,N_286);
nand U1923 (N_1923,N_393,N_507);
nand U1924 (N_1924,N_832,N_875);
nand U1925 (N_1925,N_659,N_564);
or U1926 (N_1926,N_232,N_490);
or U1927 (N_1927,N_681,N_457);
or U1928 (N_1928,N_610,N_512);
nand U1929 (N_1929,N_325,N_338);
or U1930 (N_1930,N_273,N_831);
nand U1931 (N_1931,N_518,N_297);
and U1932 (N_1932,N_250,N_320);
and U1933 (N_1933,N_396,N_316);
nand U1934 (N_1934,N_118,N_479);
nor U1935 (N_1935,N_246,N_329);
and U1936 (N_1936,N_745,N_271);
and U1937 (N_1937,N_325,N_844);
xor U1938 (N_1938,N_14,N_910);
nor U1939 (N_1939,N_997,N_667);
nor U1940 (N_1940,N_445,N_914);
or U1941 (N_1941,N_140,N_666);
nor U1942 (N_1942,N_599,N_323);
nor U1943 (N_1943,N_571,N_856);
nand U1944 (N_1944,N_869,N_102);
and U1945 (N_1945,N_624,N_864);
or U1946 (N_1946,N_67,N_610);
and U1947 (N_1947,N_19,N_379);
nand U1948 (N_1948,N_692,N_310);
or U1949 (N_1949,N_282,N_187);
or U1950 (N_1950,N_999,N_522);
nor U1951 (N_1951,N_368,N_885);
or U1952 (N_1952,N_437,N_543);
or U1953 (N_1953,N_972,N_200);
nand U1954 (N_1954,N_545,N_697);
nand U1955 (N_1955,N_921,N_53);
nor U1956 (N_1956,N_281,N_519);
or U1957 (N_1957,N_381,N_621);
nand U1958 (N_1958,N_966,N_604);
and U1959 (N_1959,N_633,N_582);
nor U1960 (N_1960,N_524,N_105);
nand U1961 (N_1961,N_520,N_869);
and U1962 (N_1962,N_16,N_589);
and U1963 (N_1963,N_272,N_523);
nor U1964 (N_1964,N_865,N_441);
nand U1965 (N_1965,N_573,N_409);
or U1966 (N_1966,N_87,N_695);
nand U1967 (N_1967,N_981,N_289);
nand U1968 (N_1968,N_567,N_911);
nand U1969 (N_1969,N_762,N_102);
nor U1970 (N_1970,N_94,N_401);
and U1971 (N_1971,N_896,N_671);
nand U1972 (N_1972,N_745,N_975);
nor U1973 (N_1973,N_412,N_435);
nand U1974 (N_1974,N_913,N_572);
nand U1975 (N_1975,N_989,N_213);
nand U1976 (N_1976,N_803,N_99);
or U1977 (N_1977,N_439,N_853);
nor U1978 (N_1978,N_731,N_830);
or U1979 (N_1979,N_383,N_168);
or U1980 (N_1980,N_56,N_672);
nor U1981 (N_1981,N_670,N_125);
or U1982 (N_1982,N_989,N_920);
and U1983 (N_1983,N_32,N_981);
or U1984 (N_1984,N_896,N_366);
nor U1985 (N_1985,N_779,N_482);
and U1986 (N_1986,N_534,N_302);
xnor U1987 (N_1987,N_410,N_644);
nor U1988 (N_1988,N_110,N_988);
nand U1989 (N_1989,N_514,N_16);
and U1990 (N_1990,N_459,N_683);
nand U1991 (N_1991,N_290,N_695);
or U1992 (N_1992,N_156,N_460);
or U1993 (N_1993,N_838,N_920);
and U1994 (N_1994,N_762,N_835);
or U1995 (N_1995,N_838,N_697);
and U1996 (N_1996,N_408,N_282);
and U1997 (N_1997,N_454,N_357);
nand U1998 (N_1998,N_634,N_792);
or U1999 (N_1999,N_807,N_75);
nand U2000 (N_2000,N_1348,N_1420);
nor U2001 (N_2001,N_1300,N_1819);
nor U2002 (N_2002,N_1567,N_1979);
and U2003 (N_2003,N_1579,N_1385);
nand U2004 (N_2004,N_1112,N_1738);
and U2005 (N_2005,N_1524,N_1386);
or U2006 (N_2006,N_1731,N_1423);
nand U2007 (N_2007,N_1742,N_1690);
or U2008 (N_2008,N_1971,N_1261);
and U2009 (N_2009,N_1628,N_1243);
nor U2010 (N_2010,N_1719,N_1970);
or U2011 (N_2011,N_1236,N_1611);
and U2012 (N_2012,N_1590,N_1571);
or U2013 (N_2013,N_1996,N_1411);
and U2014 (N_2014,N_1522,N_1600);
and U2015 (N_2015,N_1500,N_1052);
nand U2016 (N_2016,N_1637,N_1589);
and U2017 (N_2017,N_1340,N_1418);
xor U2018 (N_2018,N_1463,N_1679);
nor U2019 (N_2019,N_1059,N_1426);
and U2020 (N_2020,N_1908,N_1836);
nor U2021 (N_2021,N_1472,N_1337);
or U2022 (N_2022,N_1678,N_1911);
or U2023 (N_2023,N_1098,N_1271);
nor U2024 (N_2024,N_1498,N_1976);
or U2025 (N_2025,N_1393,N_1978);
nor U2026 (N_2026,N_1294,N_1718);
nand U2027 (N_2027,N_1026,N_1379);
and U2028 (N_2028,N_1495,N_1083);
and U2029 (N_2029,N_1964,N_1159);
nor U2030 (N_2030,N_1754,N_1278);
or U2031 (N_2031,N_1072,N_1661);
nand U2032 (N_2032,N_1684,N_1111);
nand U2033 (N_2033,N_1366,N_1410);
nor U2034 (N_2034,N_1959,N_1615);
or U2035 (N_2035,N_1141,N_1503);
nand U2036 (N_2036,N_1006,N_1541);
or U2037 (N_2037,N_1889,N_1621);
or U2038 (N_2038,N_1239,N_1943);
and U2039 (N_2039,N_1794,N_1296);
or U2040 (N_2040,N_1178,N_1228);
and U2041 (N_2041,N_1080,N_1057);
and U2042 (N_2042,N_1322,N_1939);
nand U2043 (N_2043,N_1127,N_1413);
and U2044 (N_2044,N_1848,N_1707);
and U2045 (N_2045,N_1131,N_1377);
or U2046 (N_2046,N_1174,N_1598);
nand U2047 (N_2047,N_1055,N_1345);
and U2048 (N_2048,N_1103,N_1396);
or U2049 (N_2049,N_1428,N_1431);
xor U2050 (N_2050,N_1370,N_1099);
and U2051 (N_2051,N_1948,N_1408);
or U2052 (N_2052,N_1267,N_1722);
and U2053 (N_2053,N_1042,N_1643);
nor U2054 (N_2054,N_1019,N_1710);
nor U2055 (N_2055,N_1788,N_1311);
or U2056 (N_2056,N_1597,N_1434);
nor U2057 (N_2057,N_1186,N_1049);
and U2058 (N_2058,N_1115,N_1768);
nand U2059 (N_2059,N_1818,N_1549);
nor U2060 (N_2060,N_1693,N_1044);
nand U2061 (N_2061,N_1384,N_1121);
nand U2062 (N_2062,N_1323,N_1817);
or U2063 (N_2063,N_1835,N_1721);
and U2064 (N_2064,N_1785,N_1803);
nor U2065 (N_2065,N_1381,N_1068);
xor U2066 (N_2066,N_1724,N_1190);
or U2067 (N_2067,N_1744,N_1601);
xor U2068 (N_2068,N_1977,N_1649);
or U2069 (N_2069,N_1605,N_1997);
and U2070 (N_2070,N_1667,N_1596);
nand U2071 (N_2071,N_1451,N_1839);
nand U2072 (N_2072,N_1953,N_1716);
or U2073 (N_2073,N_1856,N_1189);
or U2074 (N_2074,N_1318,N_1406);
or U2075 (N_2075,N_1488,N_1985);
or U2076 (N_2076,N_1930,N_1945);
or U2077 (N_2077,N_1346,N_1904);
or U2078 (N_2078,N_1150,N_1181);
and U2079 (N_2079,N_1466,N_1851);
nand U2080 (N_2080,N_1266,N_1265);
nor U2081 (N_2081,N_1609,N_1039);
and U2082 (N_2082,N_1101,N_1833);
nor U2083 (N_2083,N_1898,N_1882);
or U2084 (N_2084,N_1796,N_1002);
and U2085 (N_2085,N_1433,N_1805);
nand U2086 (N_2086,N_1392,N_1850);
or U2087 (N_2087,N_1879,N_1367);
nor U2088 (N_2088,N_1060,N_1260);
or U2089 (N_2089,N_1588,N_1975);
or U2090 (N_2090,N_1653,N_1214);
or U2091 (N_2091,N_1497,N_1914);
nand U2092 (N_2092,N_1523,N_1696);
nor U2093 (N_2093,N_1921,N_1051);
nand U2094 (N_2094,N_1585,N_1246);
and U2095 (N_2095,N_1264,N_1496);
and U2096 (N_2096,N_1187,N_1883);
and U2097 (N_2097,N_1148,N_1515);
nand U2098 (N_2098,N_1425,N_1586);
and U2099 (N_2099,N_1702,N_1761);
and U2100 (N_2100,N_1587,N_1258);
nor U2101 (N_2101,N_1618,N_1041);
nor U2102 (N_2102,N_1046,N_1217);
nand U2103 (N_2103,N_1884,N_1666);
and U2104 (N_2104,N_1896,N_1226);
nand U2105 (N_2105,N_1096,N_1212);
and U2106 (N_2106,N_1215,N_1000);
or U2107 (N_2107,N_1140,N_1765);
or U2108 (N_2108,N_1281,N_1946);
nand U2109 (N_2109,N_1673,N_1030);
nor U2110 (N_2110,N_1151,N_1309);
or U2111 (N_2111,N_1631,N_1619);
or U2112 (N_2112,N_1102,N_1224);
or U2113 (N_2113,N_1903,N_1745);
nand U2114 (N_2114,N_1739,N_1574);
and U2115 (N_2115,N_1545,N_1824);
nand U2116 (N_2116,N_1550,N_1638);
nor U2117 (N_2117,N_1280,N_1004);
or U2118 (N_2118,N_1772,N_1158);
nand U2119 (N_2119,N_1357,N_1798);
or U2120 (N_2120,N_1407,N_1437);
nor U2121 (N_2121,N_1380,N_1779);
nor U2122 (N_2122,N_1421,N_1025);
nor U2123 (N_2123,N_1270,N_1614);
nor U2124 (N_2124,N_1447,N_1485);
and U2125 (N_2125,N_1194,N_1610);
and U2126 (N_2126,N_1209,N_1699);
and U2127 (N_2127,N_1035,N_1519);
nand U2128 (N_2128,N_1837,N_1474);
or U2129 (N_2129,N_1078,N_1747);
and U2130 (N_2130,N_1165,N_1446);
nand U2131 (N_2131,N_1917,N_1064);
or U2132 (N_2132,N_1320,N_1100);
nand U2133 (N_2133,N_1893,N_1166);
and U2134 (N_2134,N_1480,N_1992);
and U2135 (N_2135,N_1016,N_1641);
nor U2136 (N_2136,N_1462,N_1179);
nor U2137 (N_2137,N_1729,N_1458);
nand U2138 (N_2138,N_1277,N_1771);
and U2139 (N_2139,N_1843,N_1577);
nand U2140 (N_2140,N_1352,N_1409);
or U2141 (N_2141,N_1169,N_1010);
and U2142 (N_2142,N_1302,N_1469);
and U2143 (N_2143,N_1775,N_1027);
or U2144 (N_2144,N_1897,N_1198);
and U2145 (N_2145,N_1074,N_1132);
or U2146 (N_2146,N_1725,N_1560);
nand U2147 (N_2147,N_1698,N_1923);
nor U2148 (N_2148,N_1534,N_1336);
or U2149 (N_2149,N_1966,N_1412);
nor U2150 (N_2150,N_1252,N_1024);
nand U2151 (N_2151,N_1350,N_1509);
nor U2152 (N_2152,N_1654,N_1555);
nor U2153 (N_2153,N_1402,N_1138);
and U2154 (N_2154,N_1162,N_1543);
nand U2155 (N_2155,N_1814,N_1758);
and U2156 (N_2156,N_1863,N_1616);
nand U2157 (N_2157,N_1720,N_1872);
and U2158 (N_2158,N_1234,N_1564);
or U2159 (N_2159,N_1812,N_1191);
nand U2160 (N_2160,N_1144,N_1070);
nor U2161 (N_2161,N_1008,N_1196);
or U2162 (N_2162,N_1944,N_1094);
nand U2163 (N_2163,N_1235,N_1691);
and U2164 (N_2164,N_1416,N_1983);
nor U2165 (N_2165,N_1134,N_1629);
nand U2166 (N_2166,N_1206,N_1632);
nand U2167 (N_2167,N_1283,N_1043);
nand U2168 (N_2168,N_1774,N_1401);
nor U2169 (N_2169,N_1688,N_1561);
or U2170 (N_2170,N_1343,N_1382);
and U2171 (N_2171,N_1624,N_1275);
nor U2172 (N_2172,N_1659,N_1700);
nand U2173 (N_2173,N_1442,N_1295);
or U2174 (N_2174,N_1968,N_1082);
and U2175 (N_2175,N_1544,N_1730);
xor U2176 (N_2176,N_1973,N_1118);
or U2177 (N_2177,N_1439,N_1071);
and U2178 (N_2178,N_1201,N_1886);
nand U2179 (N_2179,N_1200,N_1031);
or U2180 (N_2180,N_1777,N_1827);
or U2181 (N_2181,N_1334,N_1636);
and U2182 (N_2182,N_1237,N_1445);
nand U2183 (N_2183,N_1395,N_1987);
or U2184 (N_2184,N_1737,N_1712);
nand U2185 (N_2185,N_1332,N_1387);
nor U2186 (N_2186,N_1823,N_1962);
nor U2187 (N_2187,N_1864,N_1360);
nor U2188 (N_2188,N_1706,N_1483);
or U2189 (N_2189,N_1205,N_1842);
and U2190 (N_2190,N_1783,N_1630);
or U2191 (N_2191,N_1905,N_1368);
and U2192 (N_2192,N_1374,N_1108);
nor U2193 (N_2193,N_1161,N_1313);
and U2194 (N_2194,N_1885,N_1486);
and U2195 (N_2195,N_1849,N_1967);
xnor U2196 (N_2196,N_1665,N_1981);
or U2197 (N_2197,N_1202,N_1167);
nor U2198 (N_2198,N_1723,N_1029);
nor U2199 (N_2199,N_1928,N_1834);
and U2200 (N_2200,N_1607,N_1372);
or U2201 (N_2201,N_1963,N_1473);
and U2202 (N_2202,N_1881,N_1816);
nor U2203 (N_2203,N_1222,N_1454);
or U2204 (N_2204,N_1860,N_1135);
or U2205 (N_2205,N_1566,N_1089);
nor U2206 (N_2206,N_1859,N_1419);
or U2207 (N_2207,N_1792,N_1219);
or U2208 (N_2208,N_1404,N_1751);
nand U2209 (N_2209,N_1648,N_1084);
nor U2210 (N_2210,N_1652,N_1701);
nor U2211 (N_2211,N_1553,N_1284);
xnor U2212 (N_2212,N_1133,N_1356);
or U2213 (N_2213,N_1853,N_1766);
or U2214 (N_2214,N_1536,N_1552);
and U2215 (N_2215,N_1291,N_1347);
nand U2216 (N_2216,N_1517,N_1117);
or U2217 (N_2217,N_1991,N_1199);
or U2218 (N_2218,N_1079,N_1282);
and U2219 (N_2219,N_1533,N_1949);
or U2220 (N_2220,N_1880,N_1931);
and U2221 (N_2221,N_1890,N_1399);
and U2222 (N_2222,N_1233,N_1811);
nor U2223 (N_2223,N_1502,N_1906);
or U2224 (N_2224,N_1061,N_1163);
nand U2225 (N_2225,N_1520,N_1625);
or U2226 (N_2226,N_1770,N_1829);
and U2227 (N_2227,N_1476,N_1021);
or U2228 (N_2228,N_1984,N_1822);
nand U2229 (N_2229,N_1505,N_1542);
nand U2230 (N_2230,N_1173,N_1875);
or U2231 (N_2231,N_1565,N_1405);
nand U2232 (N_2232,N_1986,N_1918);
and U2233 (N_2233,N_1527,N_1867);
nor U2234 (N_2234,N_1249,N_1218);
nor U2235 (N_2235,N_1869,N_1335);
and U2236 (N_2236,N_1290,N_1556);
and U2237 (N_2237,N_1989,N_1965);
nor U2238 (N_2238,N_1168,N_1952);
nor U2239 (N_2239,N_1941,N_1557);
and U2240 (N_2240,N_1806,N_1248);
nor U2241 (N_2241,N_1353,N_1714);
and U2242 (N_2242,N_1563,N_1105);
xor U2243 (N_2243,N_1109,N_1171);
or U2244 (N_2244,N_1225,N_1364);
nand U2245 (N_2245,N_1398,N_1862);
or U2246 (N_2246,N_1414,N_1477);
or U2247 (N_2247,N_1531,N_1339);
or U2248 (N_2248,N_1184,N_1781);
nand U2249 (N_2249,N_1899,N_1014);
nand U2250 (N_2250,N_1680,N_1922);
nand U2251 (N_2251,N_1866,N_1358);
or U2252 (N_2252,N_1307,N_1286);
and U2253 (N_2253,N_1958,N_1241);
nand U2254 (N_2254,N_1086,N_1067);
nand U2255 (N_2255,N_1435,N_1110);
and U2256 (N_2256,N_1034,N_1521);
nor U2257 (N_2257,N_1308,N_1593);
and U2258 (N_2258,N_1066,N_1773);
nor U2259 (N_2259,N_1204,N_1732);
and U2260 (N_2260,N_1668,N_1164);
nand U2261 (N_2261,N_1499,N_1924);
nor U2262 (N_2262,N_1037,N_1230);
nand U2263 (N_2263,N_1655,N_1040);
nor U2264 (N_2264,N_1644,N_1940);
nand U2265 (N_2265,N_1316,N_1810);
nor U2266 (N_2266,N_1907,N_1790);
or U2267 (N_2267,N_1936,N_1023);
and U2268 (N_2268,N_1430,N_1182);
and U2269 (N_2269,N_1033,N_1136);
and U2270 (N_2270,N_1018,N_1925);
nor U2271 (N_2271,N_1532,N_1207);
and U2272 (N_2272,N_1954,N_1292);
or U2273 (N_2273,N_1617,N_1942);
or U2274 (N_2274,N_1444,N_1633);
or U2275 (N_2275,N_1324,N_1247);
and U2276 (N_2276,N_1888,N_1211);
nor U2277 (N_2277,N_1326,N_1464);
nand U2278 (N_2278,N_1494,N_1578);
or U2279 (N_2279,N_1916,N_1003);
or U2280 (N_2280,N_1487,N_1203);
or U2281 (N_2281,N_1139,N_1394);
nand U2282 (N_2282,N_1511,N_1288);
nor U2283 (N_2283,N_1481,N_1053);
or U2284 (N_2284,N_1076,N_1764);
nor U2285 (N_2285,N_1310,N_1746);
nor U2286 (N_2286,N_1341,N_1547);
nor U2287 (N_2287,N_1180,N_1333);
and U2288 (N_2288,N_1220,N_1852);
or U2289 (N_2289,N_1767,N_1756);
nor U2290 (N_2290,N_1753,N_1915);
nand U2291 (N_2291,N_1622,N_1955);
or U2292 (N_2292,N_1263,N_1459);
nand U2293 (N_2293,N_1902,N_1581);
and U2294 (N_2294,N_1383,N_1492);
and U2295 (N_2295,N_1778,N_1170);
nand U2296 (N_2296,N_1254,N_1646);
nand U2297 (N_2297,N_1047,N_1675);
nand U2298 (N_2298,N_1325,N_1569);
nand U2299 (N_2299,N_1583,N_1512);
nor U2300 (N_2300,N_1734,N_1048);
nor U2301 (N_2301,N_1826,N_1528);
nor U2302 (N_2302,N_1461,N_1735);
and U2303 (N_2303,N_1130,N_1453);
nand U2304 (N_2304,N_1452,N_1830);
or U2305 (N_2305,N_1301,N_1969);
or U2306 (N_2306,N_1257,N_1328);
nand U2307 (N_2307,N_1149,N_1450);
or U2308 (N_2308,N_1892,N_1660);
or U2309 (N_2309,N_1640,N_1672);
nor U2310 (N_2310,N_1752,N_1855);
nor U2311 (N_2311,N_1603,N_1650);
nand U2312 (N_2312,N_1670,N_1259);
nand U2313 (N_2313,N_1208,N_1663);
nand U2314 (N_2314,N_1832,N_1397);
nor U2315 (N_2315,N_1865,N_1327);
nand U2316 (N_2316,N_1363,N_1821);
nor U2317 (N_2317,N_1359,N_1013);
and U2318 (N_2318,N_1113,N_1216);
xnor U2319 (N_2319,N_1988,N_1009);
nor U2320 (N_2320,N_1484,N_1238);
nand U2321 (N_2321,N_1825,N_1093);
nand U2322 (N_2322,N_1657,N_1841);
nor U2323 (N_2323,N_1620,N_1901);
nor U2324 (N_2324,N_1961,N_1256);
nor U2325 (N_2325,N_1119,N_1362);
and U2326 (N_2326,N_1314,N_1268);
or U2327 (N_2327,N_1990,N_1602);
nand U2328 (N_2328,N_1526,N_1197);
and U2329 (N_2329,N_1683,N_1800);
nor U2330 (N_2330,N_1075,N_1592);
and U2331 (N_2331,N_1175,N_1791);
and U2332 (N_2332,N_1920,N_1786);
or U2333 (N_2333,N_1627,N_1831);
nor U2334 (N_2334,N_1145,N_1994);
and U2335 (N_2335,N_1365,N_1465);
nand U2336 (N_2336,N_1676,N_1424);
or U2337 (N_2337,N_1479,N_1999);
and U2338 (N_2338,N_1176,N_1183);
and U2339 (N_2339,N_1116,N_1692);
nand U2340 (N_2340,N_1262,N_1015);
and U2341 (N_2341,N_1489,N_1507);
and U2342 (N_2342,N_1669,N_1594);
nand U2343 (N_2343,N_1020,N_1705);
nor U2344 (N_2344,N_1681,N_1926);
or U2345 (N_2345,N_1441,N_1974);
or U2346 (N_2346,N_1107,N_1289);
or U2347 (N_2347,N_1674,N_1980);
or U2348 (N_2348,N_1580,N_1717);
or U2349 (N_2349,N_1595,N_1354);
nand U2350 (N_2350,N_1330,N_1715);
nor U2351 (N_2351,N_1645,N_1784);
xor U2352 (N_2352,N_1287,N_1285);
nor U2353 (N_2353,N_1575,N_1912);
nor U2354 (N_2354,N_1874,N_1799);
nand U2355 (N_2355,N_1956,N_1378);
nand U2356 (N_2356,N_1312,N_1240);
or U2357 (N_2357,N_1123,N_1537);
nor U2358 (N_2358,N_1146,N_1934);
nor U2359 (N_2359,N_1584,N_1389);
or U2360 (N_2360,N_1795,N_1455);
nor U2361 (N_2361,N_1844,N_1514);
and U2362 (N_2362,N_1697,N_1315);
nand U2363 (N_2363,N_1001,N_1376);
and U2364 (N_2364,N_1104,N_1937);
nand U2365 (N_2365,N_1085,N_1114);
and U2366 (N_2366,N_1022,N_1913);
and U2367 (N_2367,N_1960,N_1662);
or U2368 (N_2368,N_1467,N_1909);
and U2369 (N_2369,N_1160,N_1443);
or U2370 (N_2370,N_1876,N_1172);
and U2371 (N_2371,N_1137,N_1255);
and U2372 (N_2372,N_1910,N_1375);
or U2373 (N_2373,N_1687,N_1736);
or U2374 (N_2374,N_1828,N_1551);
nand U2375 (N_2375,N_1713,N_1570);
and U2376 (N_2376,N_1599,N_1143);
and U2377 (N_2377,N_1846,N_1838);
and U2378 (N_2378,N_1355,N_1935);
or U2379 (N_2379,N_1427,N_1656);
nand U2380 (N_2380,N_1279,N_1193);
nand U2381 (N_2381,N_1576,N_1436);
nand U2382 (N_2382,N_1728,N_1868);
nor U2383 (N_2383,N_1518,N_1342);
nor U2384 (N_2384,N_1642,N_1005);
and U2385 (N_2385,N_1504,N_1007);
and U2386 (N_2386,N_1801,N_1482);
or U2387 (N_2387,N_1932,N_1535);
nor U2388 (N_2388,N_1877,N_1417);
nor U2389 (N_2389,N_1854,N_1478);
or U2390 (N_2390,N_1077,N_1153);
nor U2391 (N_2391,N_1741,N_1231);
nand U2392 (N_2392,N_1686,N_1344);
and U2393 (N_2393,N_1092,N_1032);
or U2394 (N_2394,N_1703,N_1470);
and U2395 (N_2395,N_1815,N_1269);
nor U2396 (N_2396,N_1709,N_1303);
and U2397 (N_2397,N_1623,N_1229);
or U2398 (N_2398,N_1120,N_1604);
or U2399 (N_2399,N_1582,N_1319);
and U2400 (N_2400,N_1530,N_1797);
nand U2401 (N_2401,N_1708,N_1250);
nor U2402 (N_2402,N_1177,N_1506);
or U2403 (N_2403,N_1608,N_1878);
nor U2404 (N_2404,N_1185,N_1919);
or U2405 (N_2405,N_1572,N_1242);
and U2406 (N_2406,N_1449,N_1529);
and U2407 (N_2407,N_1769,N_1900);
nor U2408 (N_2408,N_1210,N_1634);
nand U2409 (N_2409,N_1142,N_1847);
and U2410 (N_2410,N_1195,N_1087);
nand U2411 (N_2411,N_1244,N_1251);
and U2412 (N_2412,N_1490,N_1927);
nor U2413 (N_2413,N_1065,N_1689);
or U2414 (N_2414,N_1998,N_1647);
nor U2415 (N_2415,N_1651,N_1017);
nand U2416 (N_2416,N_1857,N_1743);
nand U2417 (N_2417,N_1331,N_1391);
nor U2418 (N_2418,N_1272,N_1128);
nor U2419 (N_2419,N_1058,N_1403);
and U2420 (N_2420,N_1147,N_1887);
nor U2421 (N_2421,N_1090,N_1062);
or U2422 (N_2422,N_1993,N_1274);
or U2423 (N_2423,N_1568,N_1245);
nor U2424 (N_2424,N_1063,N_1606);
and U2425 (N_2425,N_1704,N_1694);
nand U2426 (N_2426,N_1789,N_1759);
nor U2427 (N_2427,N_1298,N_1038);
or U2428 (N_2428,N_1432,N_1972);
or U2429 (N_2429,N_1213,N_1011);
nand U2430 (N_2430,N_1124,N_1685);
nor U2431 (N_2431,N_1122,N_1106);
or U2432 (N_2432,N_1510,N_1513);
or U2433 (N_2433,N_1317,N_1929);
nor U2434 (N_2434,N_1152,N_1304);
and U2435 (N_2435,N_1891,N_1540);
nand U2436 (N_2436,N_1299,N_1351);
nand U2437 (N_2437,N_1858,N_1400);
nor U2438 (N_2438,N_1804,N_1097);
xor U2439 (N_2439,N_1081,N_1373);
nand U2440 (N_2440,N_1012,N_1757);
and U2441 (N_2441,N_1626,N_1760);
and U2442 (N_2442,N_1776,N_1369);
nand U2443 (N_2443,N_1305,N_1129);
or U2444 (N_2444,N_1126,N_1695);
or U2445 (N_2445,N_1156,N_1297);
nor U2446 (N_2446,N_1493,N_1782);
nand U2447 (N_2447,N_1733,N_1820);
nand U2448 (N_2448,N_1740,N_1448);
or U2449 (N_2449,N_1371,N_1787);
nand U2450 (N_2450,N_1950,N_1188);
nand U2451 (N_2451,N_1861,N_1471);
or U2452 (N_2452,N_1808,N_1045);
nor U2453 (N_2453,N_1809,N_1415);
nand U2454 (N_2454,N_1711,N_1613);
and U2455 (N_2455,N_1125,N_1306);
or U2456 (N_2456,N_1329,N_1573);
nand U2457 (N_2457,N_1460,N_1361);
nor U2458 (N_2458,N_1054,N_1845);
nand U2459 (N_2459,N_1028,N_1755);
nor U2460 (N_2460,N_1762,N_1501);
or U2461 (N_2461,N_1349,N_1321);
nand U2462 (N_2462,N_1276,N_1840);
nor U2463 (N_2463,N_1982,N_1390);
and U2464 (N_2464,N_1995,N_1095);
nand U2465 (N_2465,N_1056,N_1951);
nand U2466 (N_2466,N_1894,N_1548);
and U2467 (N_2467,N_1895,N_1591);
nand U2468 (N_2468,N_1793,N_1525);
or U2469 (N_2469,N_1677,N_1223);
nor U2470 (N_2470,N_1438,N_1508);
nor U2471 (N_2471,N_1807,N_1457);
and U2472 (N_2472,N_1870,N_1873);
nand U2473 (N_2473,N_1154,N_1073);
nand U2474 (N_2474,N_1273,N_1538);
and U2475 (N_2475,N_1658,N_1748);
and U2476 (N_2476,N_1682,N_1468);
nand U2477 (N_2477,N_1491,N_1947);
nand U2478 (N_2478,N_1664,N_1639);
or U2479 (N_2479,N_1539,N_1422);
and U2480 (N_2480,N_1227,N_1088);
or U2481 (N_2481,N_1232,N_1763);
nor U2482 (N_2482,N_1155,N_1456);
or U2483 (N_2483,N_1871,N_1727);
nor U2484 (N_2484,N_1802,N_1293);
nand U2485 (N_2485,N_1388,N_1671);
nand U2486 (N_2486,N_1440,N_1157);
nand U2487 (N_2487,N_1338,N_1475);
and U2488 (N_2488,N_1635,N_1558);
or U2489 (N_2489,N_1516,N_1559);
or U2490 (N_2490,N_1957,N_1562);
nand U2491 (N_2491,N_1749,N_1780);
nor U2492 (N_2492,N_1554,N_1813);
nand U2493 (N_2493,N_1546,N_1726);
or U2494 (N_2494,N_1091,N_1429);
nand U2495 (N_2495,N_1938,N_1221);
or U2496 (N_2496,N_1050,N_1036);
nor U2497 (N_2497,N_1750,N_1192);
nand U2498 (N_2498,N_1069,N_1612);
and U2499 (N_2499,N_1933,N_1253);
or U2500 (N_2500,N_1547,N_1762);
nor U2501 (N_2501,N_1788,N_1982);
nor U2502 (N_2502,N_1830,N_1884);
and U2503 (N_2503,N_1295,N_1024);
nand U2504 (N_2504,N_1140,N_1122);
and U2505 (N_2505,N_1640,N_1202);
nor U2506 (N_2506,N_1977,N_1429);
and U2507 (N_2507,N_1517,N_1337);
and U2508 (N_2508,N_1408,N_1562);
nor U2509 (N_2509,N_1121,N_1342);
nand U2510 (N_2510,N_1612,N_1934);
and U2511 (N_2511,N_1332,N_1271);
or U2512 (N_2512,N_1817,N_1925);
nand U2513 (N_2513,N_1789,N_1175);
or U2514 (N_2514,N_1062,N_1427);
nor U2515 (N_2515,N_1717,N_1443);
and U2516 (N_2516,N_1308,N_1312);
or U2517 (N_2517,N_1520,N_1698);
and U2518 (N_2518,N_1660,N_1297);
or U2519 (N_2519,N_1444,N_1705);
nor U2520 (N_2520,N_1804,N_1583);
or U2521 (N_2521,N_1729,N_1149);
nor U2522 (N_2522,N_1130,N_1895);
nor U2523 (N_2523,N_1893,N_1090);
or U2524 (N_2524,N_1153,N_1407);
nor U2525 (N_2525,N_1870,N_1356);
nor U2526 (N_2526,N_1481,N_1472);
or U2527 (N_2527,N_1816,N_1013);
nor U2528 (N_2528,N_1423,N_1337);
or U2529 (N_2529,N_1548,N_1056);
nor U2530 (N_2530,N_1745,N_1615);
and U2531 (N_2531,N_1243,N_1737);
and U2532 (N_2532,N_1207,N_1746);
or U2533 (N_2533,N_1673,N_1598);
and U2534 (N_2534,N_1956,N_1735);
nand U2535 (N_2535,N_1259,N_1694);
and U2536 (N_2536,N_1236,N_1061);
nor U2537 (N_2537,N_1346,N_1492);
nand U2538 (N_2538,N_1476,N_1303);
nand U2539 (N_2539,N_1119,N_1639);
nand U2540 (N_2540,N_1698,N_1423);
and U2541 (N_2541,N_1101,N_1394);
nand U2542 (N_2542,N_1070,N_1315);
and U2543 (N_2543,N_1204,N_1645);
nor U2544 (N_2544,N_1900,N_1951);
or U2545 (N_2545,N_1402,N_1653);
nand U2546 (N_2546,N_1120,N_1258);
nand U2547 (N_2547,N_1191,N_1531);
or U2548 (N_2548,N_1239,N_1023);
nand U2549 (N_2549,N_1772,N_1999);
or U2550 (N_2550,N_1523,N_1341);
and U2551 (N_2551,N_1475,N_1047);
and U2552 (N_2552,N_1122,N_1764);
nor U2553 (N_2553,N_1890,N_1699);
nand U2554 (N_2554,N_1661,N_1240);
nand U2555 (N_2555,N_1801,N_1464);
nand U2556 (N_2556,N_1266,N_1747);
nor U2557 (N_2557,N_1809,N_1839);
nand U2558 (N_2558,N_1912,N_1966);
nand U2559 (N_2559,N_1732,N_1796);
and U2560 (N_2560,N_1821,N_1090);
and U2561 (N_2561,N_1762,N_1671);
nor U2562 (N_2562,N_1984,N_1751);
and U2563 (N_2563,N_1586,N_1203);
or U2564 (N_2564,N_1966,N_1811);
and U2565 (N_2565,N_1554,N_1132);
and U2566 (N_2566,N_1289,N_1819);
nor U2567 (N_2567,N_1711,N_1621);
and U2568 (N_2568,N_1710,N_1316);
nand U2569 (N_2569,N_1889,N_1509);
nand U2570 (N_2570,N_1833,N_1359);
and U2571 (N_2571,N_1849,N_1105);
and U2572 (N_2572,N_1298,N_1081);
nand U2573 (N_2573,N_1547,N_1857);
xor U2574 (N_2574,N_1041,N_1182);
or U2575 (N_2575,N_1710,N_1699);
nor U2576 (N_2576,N_1052,N_1653);
nand U2577 (N_2577,N_1486,N_1132);
nand U2578 (N_2578,N_1912,N_1851);
or U2579 (N_2579,N_1086,N_1581);
and U2580 (N_2580,N_1545,N_1722);
nand U2581 (N_2581,N_1171,N_1122);
nor U2582 (N_2582,N_1522,N_1523);
nor U2583 (N_2583,N_1955,N_1330);
and U2584 (N_2584,N_1468,N_1982);
and U2585 (N_2585,N_1200,N_1824);
or U2586 (N_2586,N_1706,N_1710);
nand U2587 (N_2587,N_1013,N_1050);
nor U2588 (N_2588,N_1714,N_1029);
nor U2589 (N_2589,N_1205,N_1042);
nor U2590 (N_2590,N_1971,N_1241);
and U2591 (N_2591,N_1851,N_1066);
and U2592 (N_2592,N_1188,N_1527);
nand U2593 (N_2593,N_1157,N_1306);
or U2594 (N_2594,N_1539,N_1810);
and U2595 (N_2595,N_1629,N_1882);
or U2596 (N_2596,N_1900,N_1145);
nand U2597 (N_2597,N_1637,N_1449);
or U2598 (N_2598,N_1114,N_1258);
nor U2599 (N_2599,N_1842,N_1807);
nand U2600 (N_2600,N_1911,N_1061);
or U2601 (N_2601,N_1922,N_1410);
nand U2602 (N_2602,N_1675,N_1686);
nand U2603 (N_2603,N_1282,N_1799);
and U2604 (N_2604,N_1656,N_1046);
nand U2605 (N_2605,N_1413,N_1571);
or U2606 (N_2606,N_1010,N_1009);
or U2607 (N_2607,N_1468,N_1562);
and U2608 (N_2608,N_1405,N_1957);
or U2609 (N_2609,N_1265,N_1780);
or U2610 (N_2610,N_1208,N_1946);
nor U2611 (N_2611,N_1322,N_1515);
or U2612 (N_2612,N_1186,N_1558);
nor U2613 (N_2613,N_1523,N_1867);
nor U2614 (N_2614,N_1596,N_1021);
nand U2615 (N_2615,N_1920,N_1224);
and U2616 (N_2616,N_1019,N_1280);
or U2617 (N_2617,N_1977,N_1794);
nand U2618 (N_2618,N_1061,N_1923);
or U2619 (N_2619,N_1219,N_1750);
nand U2620 (N_2620,N_1747,N_1905);
or U2621 (N_2621,N_1849,N_1685);
and U2622 (N_2622,N_1798,N_1789);
or U2623 (N_2623,N_1411,N_1242);
nand U2624 (N_2624,N_1687,N_1121);
and U2625 (N_2625,N_1121,N_1205);
and U2626 (N_2626,N_1945,N_1815);
nand U2627 (N_2627,N_1397,N_1286);
and U2628 (N_2628,N_1552,N_1086);
xor U2629 (N_2629,N_1453,N_1086);
or U2630 (N_2630,N_1684,N_1058);
nand U2631 (N_2631,N_1325,N_1848);
and U2632 (N_2632,N_1091,N_1297);
nand U2633 (N_2633,N_1558,N_1308);
nor U2634 (N_2634,N_1477,N_1526);
and U2635 (N_2635,N_1443,N_1390);
and U2636 (N_2636,N_1968,N_1896);
and U2637 (N_2637,N_1928,N_1157);
or U2638 (N_2638,N_1378,N_1647);
nor U2639 (N_2639,N_1826,N_1798);
nand U2640 (N_2640,N_1854,N_1313);
nor U2641 (N_2641,N_1921,N_1945);
nand U2642 (N_2642,N_1874,N_1515);
or U2643 (N_2643,N_1779,N_1702);
and U2644 (N_2644,N_1683,N_1783);
nor U2645 (N_2645,N_1377,N_1349);
and U2646 (N_2646,N_1228,N_1060);
or U2647 (N_2647,N_1131,N_1640);
or U2648 (N_2648,N_1615,N_1718);
nor U2649 (N_2649,N_1178,N_1278);
or U2650 (N_2650,N_1266,N_1561);
nand U2651 (N_2651,N_1484,N_1787);
nor U2652 (N_2652,N_1308,N_1182);
nor U2653 (N_2653,N_1121,N_1760);
nor U2654 (N_2654,N_1387,N_1296);
or U2655 (N_2655,N_1534,N_1881);
nand U2656 (N_2656,N_1182,N_1596);
nor U2657 (N_2657,N_1606,N_1527);
and U2658 (N_2658,N_1831,N_1077);
and U2659 (N_2659,N_1051,N_1763);
nand U2660 (N_2660,N_1052,N_1896);
or U2661 (N_2661,N_1769,N_1782);
nor U2662 (N_2662,N_1262,N_1541);
nor U2663 (N_2663,N_1732,N_1438);
and U2664 (N_2664,N_1397,N_1413);
nor U2665 (N_2665,N_1462,N_1230);
or U2666 (N_2666,N_1715,N_1043);
nand U2667 (N_2667,N_1695,N_1128);
nand U2668 (N_2668,N_1826,N_1835);
nor U2669 (N_2669,N_1782,N_1647);
and U2670 (N_2670,N_1860,N_1682);
nand U2671 (N_2671,N_1992,N_1368);
or U2672 (N_2672,N_1421,N_1793);
or U2673 (N_2673,N_1963,N_1874);
or U2674 (N_2674,N_1042,N_1924);
nor U2675 (N_2675,N_1571,N_1223);
or U2676 (N_2676,N_1861,N_1381);
nand U2677 (N_2677,N_1813,N_1199);
nand U2678 (N_2678,N_1810,N_1459);
and U2679 (N_2679,N_1199,N_1474);
nor U2680 (N_2680,N_1570,N_1559);
nand U2681 (N_2681,N_1594,N_1217);
and U2682 (N_2682,N_1470,N_1485);
and U2683 (N_2683,N_1287,N_1017);
nor U2684 (N_2684,N_1663,N_1881);
or U2685 (N_2685,N_1834,N_1085);
and U2686 (N_2686,N_1352,N_1419);
nor U2687 (N_2687,N_1343,N_1193);
and U2688 (N_2688,N_1170,N_1088);
nor U2689 (N_2689,N_1213,N_1064);
nand U2690 (N_2690,N_1802,N_1638);
and U2691 (N_2691,N_1520,N_1649);
nor U2692 (N_2692,N_1841,N_1415);
and U2693 (N_2693,N_1462,N_1433);
or U2694 (N_2694,N_1383,N_1522);
nor U2695 (N_2695,N_1944,N_1763);
or U2696 (N_2696,N_1559,N_1031);
nor U2697 (N_2697,N_1545,N_1050);
and U2698 (N_2698,N_1591,N_1576);
and U2699 (N_2699,N_1126,N_1102);
nor U2700 (N_2700,N_1989,N_1395);
nand U2701 (N_2701,N_1841,N_1699);
nor U2702 (N_2702,N_1847,N_1536);
nand U2703 (N_2703,N_1629,N_1421);
and U2704 (N_2704,N_1564,N_1728);
nand U2705 (N_2705,N_1681,N_1639);
or U2706 (N_2706,N_1002,N_1345);
and U2707 (N_2707,N_1255,N_1062);
and U2708 (N_2708,N_1208,N_1280);
nor U2709 (N_2709,N_1965,N_1617);
and U2710 (N_2710,N_1306,N_1393);
nand U2711 (N_2711,N_1717,N_1739);
nand U2712 (N_2712,N_1032,N_1588);
nand U2713 (N_2713,N_1791,N_1910);
and U2714 (N_2714,N_1240,N_1556);
and U2715 (N_2715,N_1751,N_1903);
and U2716 (N_2716,N_1112,N_1697);
and U2717 (N_2717,N_1228,N_1244);
nand U2718 (N_2718,N_1383,N_1984);
or U2719 (N_2719,N_1040,N_1175);
nor U2720 (N_2720,N_1387,N_1830);
nor U2721 (N_2721,N_1480,N_1991);
nor U2722 (N_2722,N_1864,N_1389);
nor U2723 (N_2723,N_1210,N_1691);
or U2724 (N_2724,N_1134,N_1304);
and U2725 (N_2725,N_1240,N_1647);
or U2726 (N_2726,N_1859,N_1290);
nand U2727 (N_2727,N_1578,N_1469);
and U2728 (N_2728,N_1985,N_1286);
nand U2729 (N_2729,N_1815,N_1217);
and U2730 (N_2730,N_1391,N_1334);
and U2731 (N_2731,N_1159,N_1452);
nand U2732 (N_2732,N_1711,N_1415);
or U2733 (N_2733,N_1855,N_1614);
and U2734 (N_2734,N_1103,N_1359);
or U2735 (N_2735,N_1363,N_1933);
and U2736 (N_2736,N_1561,N_1992);
nand U2737 (N_2737,N_1591,N_1038);
nor U2738 (N_2738,N_1551,N_1124);
nor U2739 (N_2739,N_1351,N_1011);
nor U2740 (N_2740,N_1620,N_1248);
nand U2741 (N_2741,N_1306,N_1418);
nand U2742 (N_2742,N_1295,N_1485);
or U2743 (N_2743,N_1494,N_1901);
nand U2744 (N_2744,N_1373,N_1276);
or U2745 (N_2745,N_1247,N_1439);
or U2746 (N_2746,N_1021,N_1376);
nor U2747 (N_2747,N_1382,N_1389);
nand U2748 (N_2748,N_1844,N_1300);
nor U2749 (N_2749,N_1809,N_1930);
or U2750 (N_2750,N_1437,N_1520);
or U2751 (N_2751,N_1830,N_1770);
and U2752 (N_2752,N_1458,N_1482);
nand U2753 (N_2753,N_1924,N_1462);
nor U2754 (N_2754,N_1208,N_1811);
nor U2755 (N_2755,N_1059,N_1488);
or U2756 (N_2756,N_1631,N_1101);
nor U2757 (N_2757,N_1225,N_1493);
nand U2758 (N_2758,N_1931,N_1905);
or U2759 (N_2759,N_1834,N_1111);
or U2760 (N_2760,N_1782,N_1054);
or U2761 (N_2761,N_1408,N_1551);
nand U2762 (N_2762,N_1499,N_1669);
and U2763 (N_2763,N_1635,N_1818);
nor U2764 (N_2764,N_1203,N_1095);
or U2765 (N_2765,N_1516,N_1818);
or U2766 (N_2766,N_1009,N_1338);
nand U2767 (N_2767,N_1266,N_1500);
nor U2768 (N_2768,N_1740,N_1142);
nand U2769 (N_2769,N_1525,N_1405);
or U2770 (N_2770,N_1281,N_1310);
nor U2771 (N_2771,N_1729,N_1933);
and U2772 (N_2772,N_1096,N_1377);
and U2773 (N_2773,N_1358,N_1141);
nand U2774 (N_2774,N_1933,N_1306);
nor U2775 (N_2775,N_1308,N_1575);
or U2776 (N_2776,N_1660,N_1960);
nor U2777 (N_2777,N_1844,N_1460);
and U2778 (N_2778,N_1848,N_1201);
nor U2779 (N_2779,N_1055,N_1597);
xor U2780 (N_2780,N_1918,N_1849);
and U2781 (N_2781,N_1206,N_1968);
and U2782 (N_2782,N_1195,N_1265);
nand U2783 (N_2783,N_1321,N_1097);
nand U2784 (N_2784,N_1432,N_1943);
or U2785 (N_2785,N_1982,N_1831);
or U2786 (N_2786,N_1028,N_1925);
nand U2787 (N_2787,N_1548,N_1252);
nand U2788 (N_2788,N_1910,N_1337);
nand U2789 (N_2789,N_1024,N_1555);
nor U2790 (N_2790,N_1912,N_1627);
nand U2791 (N_2791,N_1864,N_1980);
and U2792 (N_2792,N_1225,N_1330);
nor U2793 (N_2793,N_1800,N_1614);
or U2794 (N_2794,N_1008,N_1776);
nand U2795 (N_2795,N_1286,N_1782);
nand U2796 (N_2796,N_1351,N_1438);
nand U2797 (N_2797,N_1012,N_1374);
and U2798 (N_2798,N_1651,N_1397);
and U2799 (N_2799,N_1235,N_1057);
nor U2800 (N_2800,N_1929,N_1549);
and U2801 (N_2801,N_1598,N_1752);
nor U2802 (N_2802,N_1337,N_1140);
nand U2803 (N_2803,N_1842,N_1556);
or U2804 (N_2804,N_1147,N_1725);
nand U2805 (N_2805,N_1637,N_1907);
and U2806 (N_2806,N_1563,N_1410);
or U2807 (N_2807,N_1846,N_1720);
and U2808 (N_2808,N_1396,N_1573);
or U2809 (N_2809,N_1049,N_1880);
nor U2810 (N_2810,N_1022,N_1679);
or U2811 (N_2811,N_1572,N_1353);
nor U2812 (N_2812,N_1168,N_1684);
nor U2813 (N_2813,N_1645,N_1104);
nand U2814 (N_2814,N_1486,N_1639);
nand U2815 (N_2815,N_1288,N_1877);
and U2816 (N_2816,N_1725,N_1708);
or U2817 (N_2817,N_1177,N_1926);
xor U2818 (N_2818,N_1770,N_1955);
and U2819 (N_2819,N_1007,N_1575);
or U2820 (N_2820,N_1382,N_1804);
or U2821 (N_2821,N_1926,N_1768);
and U2822 (N_2822,N_1137,N_1368);
or U2823 (N_2823,N_1572,N_1487);
or U2824 (N_2824,N_1544,N_1036);
and U2825 (N_2825,N_1142,N_1164);
nand U2826 (N_2826,N_1431,N_1159);
nand U2827 (N_2827,N_1716,N_1328);
and U2828 (N_2828,N_1526,N_1870);
and U2829 (N_2829,N_1474,N_1100);
nand U2830 (N_2830,N_1998,N_1089);
or U2831 (N_2831,N_1488,N_1239);
nand U2832 (N_2832,N_1911,N_1976);
nand U2833 (N_2833,N_1854,N_1229);
or U2834 (N_2834,N_1534,N_1849);
nor U2835 (N_2835,N_1735,N_1592);
xor U2836 (N_2836,N_1908,N_1308);
nor U2837 (N_2837,N_1813,N_1642);
nor U2838 (N_2838,N_1085,N_1134);
or U2839 (N_2839,N_1062,N_1423);
and U2840 (N_2840,N_1904,N_1271);
and U2841 (N_2841,N_1521,N_1738);
or U2842 (N_2842,N_1064,N_1378);
nor U2843 (N_2843,N_1226,N_1619);
and U2844 (N_2844,N_1971,N_1697);
nor U2845 (N_2845,N_1548,N_1608);
nor U2846 (N_2846,N_1215,N_1199);
and U2847 (N_2847,N_1834,N_1835);
or U2848 (N_2848,N_1145,N_1752);
or U2849 (N_2849,N_1752,N_1151);
nor U2850 (N_2850,N_1385,N_1530);
nor U2851 (N_2851,N_1199,N_1462);
or U2852 (N_2852,N_1512,N_1504);
and U2853 (N_2853,N_1229,N_1434);
nor U2854 (N_2854,N_1305,N_1919);
or U2855 (N_2855,N_1516,N_1132);
nand U2856 (N_2856,N_1669,N_1331);
and U2857 (N_2857,N_1236,N_1969);
nor U2858 (N_2858,N_1051,N_1035);
and U2859 (N_2859,N_1350,N_1933);
nor U2860 (N_2860,N_1212,N_1422);
or U2861 (N_2861,N_1285,N_1085);
or U2862 (N_2862,N_1777,N_1498);
or U2863 (N_2863,N_1642,N_1790);
or U2864 (N_2864,N_1255,N_1837);
and U2865 (N_2865,N_1769,N_1209);
nor U2866 (N_2866,N_1909,N_1361);
nor U2867 (N_2867,N_1535,N_1256);
nor U2868 (N_2868,N_1657,N_1594);
and U2869 (N_2869,N_1116,N_1810);
nand U2870 (N_2870,N_1073,N_1831);
nand U2871 (N_2871,N_1085,N_1409);
and U2872 (N_2872,N_1680,N_1980);
nand U2873 (N_2873,N_1156,N_1355);
nor U2874 (N_2874,N_1104,N_1465);
nand U2875 (N_2875,N_1647,N_1755);
nor U2876 (N_2876,N_1275,N_1102);
and U2877 (N_2877,N_1342,N_1679);
nand U2878 (N_2878,N_1477,N_1517);
and U2879 (N_2879,N_1989,N_1013);
and U2880 (N_2880,N_1694,N_1797);
nor U2881 (N_2881,N_1820,N_1540);
nand U2882 (N_2882,N_1021,N_1003);
or U2883 (N_2883,N_1128,N_1677);
and U2884 (N_2884,N_1972,N_1979);
nor U2885 (N_2885,N_1796,N_1755);
nor U2886 (N_2886,N_1847,N_1106);
nand U2887 (N_2887,N_1432,N_1023);
or U2888 (N_2888,N_1058,N_1517);
and U2889 (N_2889,N_1950,N_1916);
or U2890 (N_2890,N_1587,N_1627);
nand U2891 (N_2891,N_1090,N_1141);
and U2892 (N_2892,N_1500,N_1703);
nor U2893 (N_2893,N_1082,N_1530);
and U2894 (N_2894,N_1513,N_1525);
nand U2895 (N_2895,N_1014,N_1336);
nand U2896 (N_2896,N_1149,N_1212);
or U2897 (N_2897,N_1442,N_1123);
or U2898 (N_2898,N_1285,N_1587);
and U2899 (N_2899,N_1244,N_1064);
or U2900 (N_2900,N_1835,N_1745);
xnor U2901 (N_2901,N_1773,N_1546);
nand U2902 (N_2902,N_1884,N_1592);
nor U2903 (N_2903,N_1819,N_1429);
or U2904 (N_2904,N_1721,N_1833);
or U2905 (N_2905,N_1637,N_1305);
nor U2906 (N_2906,N_1708,N_1490);
or U2907 (N_2907,N_1046,N_1153);
or U2908 (N_2908,N_1760,N_1447);
and U2909 (N_2909,N_1138,N_1172);
nor U2910 (N_2910,N_1871,N_1425);
or U2911 (N_2911,N_1828,N_1112);
nor U2912 (N_2912,N_1282,N_1747);
nand U2913 (N_2913,N_1022,N_1081);
nor U2914 (N_2914,N_1881,N_1538);
nor U2915 (N_2915,N_1771,N_1349);
nor U2916 (N_2916,N_1466,N_1526);
and U2917 (N_2917,N_1534,N_1003);
and U2918 (N_2918,N_1541,N_1111);
or U2919 (N_2919,N_1450,N_1318);
and U2920 (N_2920,N_1000,N_1763);
or U2921 (N_2921,N_1929,N_1556);
and U2922 (N_2922,N_1054,N_1015);
nand U2923 (N_2923,N_1140,N_1735);
and U2924 (N_2924,N_1941,N_1172);
or U2925 (N_2925,N_1270,N_1921);
or U2926 (N_2926,N_1081,N_1932);
and U2927 (N_2927,N_1206,N_1687);
nand U2928 (N_2928,N_1688,N_1803);
or U2929 (N_2929,N_1169,N_1767);
and U2930 (N_2930,N_1727,N_1779);
or U2931 (N_2931,N_1665,N_1952);
or U2932 (N_2932,N_1896,N_1580);
nand U2933 (N_2933,N_1433,N_1499);
and U2934 (N_2934,N_1680,N_1888);
nor U2935 (N_2935,N_1917,N_1092);
or U2936 (N_2936,N_1424,N_1498);
and U2937 (N_2937,N_1827,N_1991);
or U2938 (N_2938,N_1081,N_1177);
or U2939 (N_2939,N_1017,N_1697);
nor U2940 (N_2940,N_1776,N_1855);
or U2941 (N_2941,N_1993,N_1179);
nand U2942 (N_2942,N_1917,N_1892);
nand U2943 (N_2943,N_1972,N_1580);
or U2944 (N_2944,N_1460,N_1402);
nand U2945 (N_2945,N_1404,N_1451);
or U2946 (N_2946,N_1833,N_1391);
nand U2947 (N_2947,N_1558,N_1994);
nor U2948 (N_2948,N_1115,N_1275);
and U2949 (N_2949,N_1651,N_1385);
nand U2950 (N_2950,N_1601,N_1202);
and U2951 (N_2951,N_1001,N_1266);
nand U2952 (N_2952,N_1910,N_1390);
and U2953 (N_2953,N_1525,N_1748);
or U2954 (N_2954,N_1949,N_1444);
nor U2955 (N_2955,N_1899,N_1921);
nand U2956 (N_2956,N_1520,N_1183);
nand U2957 (N_2957,N_1790,N_1718);
or U2958 (N_2958,N_1878,N_1715);
nand U2959 (N_2959,N_1422,N_1297);
or U2960 (N_2960,N_1543,N_1246);
or U2961 (N_2961,N_1109,N_1676);
and U2962 (N_2962,N_1721,N_1240);
and U2963 (N_2963,N_1811,N_1293);
and U2964 (N_2964,N_1090,N_1960);
nor U2965 (N_2965,N_1334,N_1207);
nor U2966 (N_2966,N_1325,N_1506);
nor U2967 (N_2967,N_1142,N_1596);
or U2968 (N_2968,N_1123,N_1379);
nand U2969 (N_2969,N_1380,N_1024);
nor U2970 (N_2970,N_1444,N_1723);
or U2971 (N_2971,N_1454,N_1354);
nand U2972 (N_2972,N_1666,N_1624);
nand U2973 (N_2973,N_1122,N_1687);
nand U2974 (N_2974,N_1781,N_1215);
and U2975 (N_2975,N_1278,N_1562);
nor U2976 (N_2976,N_1293,N_1154);
or U2977 (N_2977,N_1192,N_1933);
nand U2978 (N_2978,N_1918,N_1996);
and U2979 (N_2979,N_1178,N_1964);
or U2980 (N_2980,N_1969,N_1296);
xnor U2981 (N_2981,N_1757,N_1167);
and U2982 (N_2982,N_1132,N_1582);
nor U2983 (N_2983,N_1450,N_1316);
or U2984 (N_2984,N_1199,N_1621);
or U2985 (N_2985,N_1511,N_1561);
nor U2986 (N_2986,N_1802,N_1866);
and U2987 (N_2987,N_1185,N_1718);
nor U2988 (N_2988,N_1498,N_1693);
nor U2989 (N_2989,N_1761,N_1000);
or U2990 (N_2990,N_1598,N_1878);
nand U2991 (N_2991,N_1189,N_1474);
nor U2992 (N_2992,N_1178,N_1223);
xnor U2993 (N_2993,N_1926,N_1350);
nand U2994 (N_2994,N_1834,N_1976);
and U2995 (N_2995,N_1703,N_1936);
and U2996 (N_2996,N_1914,N_1113);
nor U2997 (N_2997,N_1284,N_1375);
or U2998 (N_2998,N_1555,N_1174);
nand U2999 (N_2999,N_1011,N_1241);
nand UO_0 (O_0,N_2234,N_2991);
and UO_1 (O_1,N_2866,N_2454);
and UO_2 (O_2,N_2335,N_2878);
nand UO_3 (O_3,N_2474,N_2941);
and UO_4 (O_4,N_2802,N_2357);
or UO_5 (O_5,N_2914,N_2536);
or UO_6 (O_6,N_2289,N_2537);
or UO_7 (O_7,N_2705,N_2530);
nand UO_8 (O_8,N_2689,N_2475);
nor UO_9 (O_9,N_2328,N_2861);
or UO_10 (O_10,N_2130,N_2112);
nor UO_11 (O_11,N_2815,N_2937);
nand UO_12 (O_12,N_2459,N_2901);
and UO_13 (O_13,N_2392,N_2293);
or UO_14 (O_14,N_2143,N_2166);
or UO_15 (O_15,N_2349,N_2133);
nor UO_16 (O_16,N_2822,N_2152);
or UO_17 (O_17,N_2642,N_2033);
nor UO_18 (O_18,N_2498,N_2850);
nor UO_19 (O_19,N_2927,N_2180);
or UO_20 (O_20,N_2731,N_2630);
or UO_21 (O_21,N_2207,N_2363);
nand UO_22 (O_22,N_2424,N_2750);
nand UO_23 (O_23,N_2742,N_2585);
nand UO_24 (O_24,N_2471,N_2535);
nand UO_25 (O_25,N_2276,N_2626);
and UO_26 (O_26,N_2001,N_2285);
and UO_27 (O_27,N_2528,N_2496);
or UO_28 (O_28,N_2990,N_2087);
and UO_29 (O_29,N_2519,N_2681);
and UO_30 (O_30,N_2075,N_2716);
and UO_31 (O_31,N_2090,N_2604);
nand UO_32 (O_32,N_2921,N_2608);
nand UO_33 (O_33,N_2910,N_2957);
or UO_34 (O_34,N_2402,N_2377);
or UO_35 (O_35,N_2557,N_2317);
nand UO_36 (O_36,N_2504,N_2398);
and UO_37 (O_37,N_2186,N_2659);
or UO_38 (O_38,N_2366,N_2623);
or UO_39 (O_39,N_2146,N_2666);
nand UO_40 (O_40,N_2987,N_2477);
nand UO_41 (O_41,N_2397,N_2575);
or UO_42 (O_42,N_2789,N_2939);
or UO_43 (O_43,N_2230,N_2974);
nand UO_44 (O_44,N_2124,N_2325);
or UO_45 (O_45,N_2416,N_2027);
nand UO_46 (O_46,N_2120,N_2997);
and UO_47 (O_47,N_2999,N_2661);
or UO_48 (O_48,N_2687,N_2645);
nor UO_49 (O_49,N_2396,N_2839);
nor UO_50 (O_50,N_2610,N_2988);
and UO_51 (O_51,N_2707,N_2523);
or UO_52 (O_52,N_2801,N_2669);
nand UO_53 (O_53,N_2151,N_2805);
nor UO_54 (O_54,N_2011,N_2653);
or UO_55 (O_55,N_2488,N_2235);
and UO_56 (O_56,N_2930,N_2270);
or UO_57 (O_57,N_2702,N_2036);
or UO_58 (O_58,N_2310,N_2029);
and UO_59 (O_59,N_2521,N_2158);
and UO_60 (O_60,N_2017,N_2843);
or UO_61 (O_61,N_2899,N_2970);
nor UO_62 (O_62,N_2732,N_2177);
nand UO_63 (O_63,N_2190,N_2852);
and UO_64 (O_64,N_2749,N_2332);
or UO_65 (O_65,N_2923,N_2596);
nand UO_66 (O_66,N_2863,N_2563);
or UO_67 (O_67,N_2404,N_2426);
nand UO_68 (O_68,N_2294,N_2381);
nand UO_69 (O_69,N_2055,N_2409);
and UO_70 (O_70,N_2943,N_2217);
nor UO_71 (O_71,N_2612,N_2356);
or UO_72 (O_72,N_2111,N_2358);
nand UO_73 (O_73,N_2338,N_2347);
or UO_74 (O_74,N_2628,N_2600);
and UO_75 (O_75,N_2007,N_2127);
and UO_76 (O_76,N_2204,N_2751);
nor UO_77 (O_77,N_2261,N_2136);
nand UO_78 (O_78,N_2083,N_2110);
nor UO_79 (O_79,N_2460,N_2492);
nor UO_80 (O_80,N_2466,N_2214);
or UO_81 (O_81,N_2713,N_2387);
nor UO_82 (O_82,N_2942,N_2532);
or UO_83 (O_83,N_2539,N_2425);
nand UO_84 (O_84,N_2674,N_2697);
nand UO_85 (O_85,N_2983,N_2300);
or UO_86 (O_86,N_2044,N_2076);
nor UO_87 (O_87,N_2516,N_2208);
or UO_88 (O_88,N_2021,N_2609);
nand UO_89 (O_89,N_2820,N_2710);
and UO_90 (O_90,N_2003,N_2547);
and UO_91 (O_91,N_2922,N_2148);
nor UO_92 (O_92,N_2336,N_2643);
or UO_93 (O_93,N_2531,N_2868);
and UO_94 (O_94,N_2159,N_2961);
or UO_95 (O_95,N_2566,N_2485);
and UO_96 (O_96,N_2810,N_2018);
or UO_97 (O_97,N_2388,N_2156);
and UO_98 (O_98,N_2541,N_2342);
nand UO_99 (O_99,N_2389,N_2995);
or UO_100 (O_100,N_2655,N_2147);
and UO_101 (O_101,N_2854,N_2509);
and UO_102 (O_102,N_2581,N_2828);
nand UO_103 (O_103,N_2144,N_2238);
or UO_104 (O_104,N_2793,N_2639);
nand UO_105 (O_105,N_2950,N_2114);
or UO_106 (O_106,N_2685,N_2520);
nor UO_107 (O_107,N_2340,N_2501);
and UO_108 (O_108,N_2161,N_2200);
nor UO_109 (O_109,N_2369,N_2879);
and UO_110 (O_110,N_2020,N_2095);
nor UO_111 (O_111,N_2502,N_2318);
and UO_112 (O_112,N_2002,N_2976);
and UO_113 (O_113,N_2675,N_2853);
and UO_114 (O_114,N_2179,N_2719);
nand UO_115 (O_115,N_2272,N_2137);
or UO_116 (O_116,N_2503,N_2320);
and UO_117 (O_117,N_2614,N_2327);
or UO_118 (O_118,N_2533,N_2678);
nand UO_119 (O_119,N_2924,N_2589);
nand UO_120 (O_120,N_2082,N_2763);
nor UO_121 (O_121,N_2042,N_2032);
nand UO_122 (O_122,N_2684,N_2829);
nand UO_123 (O_123,N_2876,N_2907);
nand UO_124 (O_124,N_2920,N_2592);
or UO_125 (O_125,N_2522,N_2712);
nand UO_126 (O_126,N_2479,N_2091);
nor UO_127 (O_127,N_2915,N_2184);
nand UO_128 (O_128,N_2804,N_2119);
or UO_129 (O_129,N_2182,N_2965);
nor UO_130 (O_130,N_2478,N_2054);
or UO_131 (O_131,N_2844,N_2051);
nor UO_132 (O_132,N_2275,N_2025);
and UO_133 (O_133,N_2679,N_2255);
or UO_134 (O_134,N_2438,N_2631);
or UO_135 (O_135,N_2237,N_2613);
nor UO_136 (O_136,N_2252,N_2633);
and UO_137 (O_137,N_2641,N_2744);
nand UO_138 (O_138,N_2004,N_2405);
nor UO_139 (O_139,N_2295,N_2725);
nor UO_140 (O_140,N_2692,N_2005);
and UO_141 (O_141,N_2445,N_2231);
or UO_142 (O_142,N_2418,N_2491);
nor UO_143 (O_143,N_2066,N_2619);
nor UO_144 (O_144,N_2071,N_2383);
and UO_145 (O_145,N_2931,N_2181);
nor UO_146 (O_146,N_2785,N_2851);
or UO_147 (O_147,N_2380,N_2164);
nand UO_148 (O_148,N_2354,N_2824);
or UO_149 (O_149,N_2078,N_2059);
or UO_150 (O_150,N_2470,N_2896);
nand UO_151 (O_151,N_2220,N_2508);
or UO_152 (O_152,N_2319,N_2656);
nand UO_153 (O_153,N_2061,N_2169);
and UO_154 (O_154,N_2529,N_2215);
nor UO_155 (O_155,N_2000,N_2193);
nand UO_156 (O_156,N_2873,N_2093);
and UO_157 (O_157,N_2913,N_2359);
or UO_158 (O_158,N_2654,N_2188);
nand UO_159 (O_159,N_2772,N_2728);
nor UO_160 (O_160,N_2212,N_2154);
nand UO_161 (O_161,N_2086,N_2287);
nand UO_162 (O_162,N_2467,N_2792);
or UO_163 (O_163,N_2350,N_2780);
nand UO_164 (O_164,N_2781,N_2885);
nor UO_165 (O_165,N_2374,N_2009);
or UO_166 (O_166,N_2830,N_2089);
nor UO_167 (O_167,N_2651,N_2216);
nor UO_168 (O_168,N_2831,N_2764);
nor UO_169 (O_169,N_2567,N_2218);
or UO_170 (O_170,N_2473,N_2788);
or UO_171 (O_171,N_2761,N_2098);
nand UO_172 (O_172,N_2281,N_2172);
and UO_173 (O_173,N_2891,N_2233);
nor UO_174 (O_174,N_2371,N_2736);
and UO_175 (O_175,N_2715,N_2813);
nand UO_176 (O_176,N_2209,N_2867);
and UO_177 (O_177,N_2875,N_2149);
or UO_178 (O_178,N_2433,N_2883);
and UO_179 (O_179,N_2232,N_2448);
and UO_180 (O_180,N_2065,N_2431);
nand UO_181 (O_181,N_2219,N_2814);
or UO_182 (O_182,N_2480,N_2067);
nor UO_183 (O_183,N_2056,N_2578);
nand UO_184 (O_184,N_2518,N_2576);
or UO_185 (O_185,N_2379,N_2259);
nor UO_186 (O_186,N_2583,N_2511);
nor UO_187 (O_187,N_2443,N_2045);
or UO_188 (O_188,N_2419,N_2352);
xor UO_189 (O_189,N_2227,N_2741);
nand UO_190 (O_190,N_2570,N_2420);
and UO_191 (O_191,N_2131,N_2265);
and UO_192 (O_192,N_2128,N_2399);
nand UO_193 (O_193,N_2205,N_2629);
nand UO_194 (O_194,N_2390,N_2979);
nor UO_195 (O_195,N_2249,N_2267);
and UO_196 (O_196,N_2301,N_2006);
nand UO_197 (O_197,N_2198,N_2196);
nor UO_198 (O_198,N_2436,N_2577);
nand UO_199 (O_199,N_2401,N_2334);
and UO_200 (O_200,N_2616,N_2437);
nand UO_201 (O_201,N_2393,N_2429);
nand UO_202 (O_202,N_2283,N_2947);
or UO_203 (O_203,N_2412,N_2554);
or UO_204 (O_204,N_2959,N_2562);
or UO_205 (O_205,N_2224,N_2746);
nand UO_206 (O_206,N_2934,N_2415);
and UO_207 (O_207,N_2010,N_2928);
or UO_208 (O_208,N_2862,N_2245);
or UO_209 (O_209,N_2263,N_2620);
nand UO_210 (O_210,N_2348,N_2672);
and UO_211 (O_211,N_2439,N_2680);
nand UO_212 (O_212,N_2842,N_2493);
and UO_213 (O_213,N_2700,N_2070);
and UO_214 (O_214,N_2375,N_2253);
or UO_215 (O_215,N_2135,N_2632);
nand UO_216 (O_216,N_2989,N_2601);
or UO_217 (O_217,N_2428,N_2919);
or UO_218 (O_218,N_2819,N_2786);
or UO_219 (O_219,N_2647,N_2973);
nor UO_220 (O_220,N_2298,N_2667);
nand UO_221 (O_221,N_2704,N_2838);
or UO_222 (O_222,N_2201,N_2247);
nor UO_223 (O_223,N_2775,N_2549);
and UO_224 (O_224,N_2050,N_2948);
and UO_225 (O_225,N_2463,N_2622);
and UO_226 (O_226,N_2037,N_2895);
nor UO_227 (O_227,N_2625,N_2297);
nor UO_228 (O_228,N_2484,N_2964);
or UO_229 (O_229,N_2057,N_2903);
nor UO_230 (O_230,N_2755,N_2676);
nor UO_231 (O_231,N_2892,N_2548);
and UO_232 (O_232,N_2422,N_2580);
or UO_233 (O_233,N_2703,N_2902);
or UO_234 (O_234,N_2307,N_2243);
nand UO_235 (O_235,N_2456,N_2229);
nor UO_236 (O_236,N_2514,N_2933);
or UO_237 (O_237,N_2228,N_2175);
nor UO_238 (O_238,N_2462,N_2063);
or UO_239 (O_239,N_2818,N_2579);
or UO_240 (O_240,N_2798,N_2553);
and UO_241 (O_241,N_2041,N_2992);
or UO_242 (O_242,N_2753,N_2362);
or UO_243 (O_243,N_2121,N_2869);
nor UO_244 (O_244,N_2729,N_2808);
nand UO_245 (O_245,N_2617,N_2835);
nand UO_246 (O_246,N_2960,N_2650);
and UO_247 (O_247,N_2291,N_2039);
or UO_248 (O_248,N_2395,N_2150);
or UO_249 (O_249,N_2968,N_2925);
nor UO_250 (O_250,N_2202,N_2823);
or UO_251 (O_251,N_2752,N_2160);
and UO_252 (O_252,N_2627,N_2115);
nor UO_253 (O_253,N_2178,N_2026);
nand UO_254 (O_254,N_2926,N_2453);
and UO_255 (O_255,N_2062,N_2945);
and UO_256 (O_256,N_2351,N_2183);
or UO_257 (O_257,N_2837,N_2337);
and UO_258 (O_258,N_2315,N_2646);
or UO_259 (O_259,N_2884,N_2497);
nand UO_260 (O_260,N_2889,N_2394);
nand UO_261 (O_261,N_2203,N_2652);
nand UO_262 (O_262,N_2391,N_2993);
and UO_263 (O_263,N_2546,N_2094);
nor UO_264 (O_264,N_2047,N_2806);
nor UO_265 (O_265,N_2157,N_2048);
xor UO_266 (O_266,N_2542,N_2308);
and UO_267 (O_267,N_2584,N_2386);
and UO_268 (O_268,N_2413,N_2104);
or UO_269 (O_269,N_2225,N_2597);
and UO_270 (O_270,N_2917,N_2944);
or UO_271 (O_271,N_2260,N_2985);
nand UO_272 (O_272,N_2880,N_2423);
and UO_273 (O_273,N_2552,N_2013);
and UO_274 (O_274,N_2735,N_2545);
and UO_275 (O_275,N_2803,N_2743);
or UO_276 (O_276,N_2897,N_2043);
or UO_277 (O_277,N_2540,N_2199);
or UO_278 (O_278,N_2754,N_2440);
nand UO_279 (O_279,N_2640,N_2882);
nand UO_280 (O_280,N_2058,N_2723);
nand UO_281 (O_281,N_2333,N_2206);
and UO_282 (O_282,N_2101,N_2777);
and UO_283 (O_283,N_2904,N_2257);
or UO_284 (O_284,N_2686,N_2079);
and UO_285 (O_285,N_2197,N_2872);
or UO_286 (O_286,N_2611,N_2773);
or UO_287 (O_287,N_2572,N_2194);
and UO_288 (O_288,N_2586,N_2140);
nand UO_289 (O_289,N_2299,N_2012);
nor UO_290 (O_290,N_2527,N_2343);
and UO_291 (O_291,N_2117,N_2860);
nand UO_292 (O_292,N_2008,N_2417);
nor UO_293 (O_293,N_2015,N_2469);
nor UO_294 (O_294,N_2796,N_2367);
and UO_295 (O_295,N_2911,N_2797);
and UO_296 (O_296,N_2370,N_2077);
nor UO_297 (O_297,N_2345,N_2962);
nand UO_298 (O_298,N_2740,N_2072);
or UO_299 (O_299,N_2734,N_2145);
and UO_300 (O_300,N_2022,N_2538);
nand UO_301 (O_301,N_2846,N_2408);
nand UO_302 (O_302,N_2765,N_2384);
nor UO_303 (O_303,N_2014,N_2324);
or UO_304 (O_304,N_2167,N_2305);
or UO_305 (O_305,N_2168,N_2946);
nor UO_306 (O_306,N_2449,N_2967);
nand UO_307 (O_307,N_2840,N_2176);
nor UO_308 (O_308,N_2069,N_2099);
and UO_309 (O_309,N_2118,N_2770);
and UO_310 (O_310,N_2932,N_2778);
and UO_311 (O_311,N_2634,N_2649);
nand UO_312 (O_312,N_2938,N_2721);
or UO_313 (O_313,N_2302,N_2747);
and UO_314 (O_314,N_2598,N_2331);
and UO_315 (O_315,N_2564,N_2816);
or UO_316 (O_316,N_2123,N_2929);
nor UO_317 (O_317,N_2784,N_2790);
nand UO_318 (O_318,N_2845,N_2918);
nor UO_319 (O_319,N_2053,N_2155);
nor UO_320 (O_320,N_2126,N_2284);
and UO_321 (O_321,N_2660,N_2452);
nor UO_322 (O_322,N_2574,N_2500);
and UO_323 (O_323,N_2906,N_2241);
nand UO_324 (O_324,N_2556,N_2142);
nor UO_325 (O_325,N_2870,N_2936);
nor UO_326 (O_326,N_2971,N_2407);
or UO_327 (O_327,N_2483,N_2256);
nand UO_328 (O_328,N_2213,N_2558);
nor UO_329 (O_329,N_2210,N_2951);
nand UO_330 (O_330,N_2986,N_2759);
and UO_331 (O_331,N_2534,N_2739);
xnor UO_332 (O_332,N_2323,N_2636);
nor UO_333 (O_333,N_2834,N_2096);
nand UO_334 (O_334,N_2637,N_2688);
nand UO_335 (O_335,N_2254,N_2016);
and UO_336 (O_336,N_2092,N_2696);
nand UO_337 (O_337,N_2344,N_2693);
or UO_338 (O_338,N_2403,N_2368);
nor UO_339 (O_339,N_2410,N_2264);
and UO_340 (O_340,N_2956,N_2758);
nor UO_341 (O_341,N_2515,N_2174);
nor UO_342 (O_342,N_2490,N_2455);
and UO_343 (O_343,N_2242,N_2355);
and UO_344 (O_344,N_2624,N_2821);
nor UO_345 (O_345,N_2849,N_2321);
or UO_346 (O_346,N_2841,N_2836);
or UO_347 (O_347,N_2827,N_2106);
or UO_348 (O_348,N_2060,N_2271);
and UO_349 (O_349,N_2881,N_2125);
or UO_350 (O_350,N_2288,N_2116);
and UO_351 (O_351,N_2720,N_2958);
or UO_352 (O_352,N_2046,N_2594);
and UO_353 (O_353,N_2486,N_2664);
or UO_354 (O_354,N_2165,N_2809);
and UO_355 (O_355,N_2191,N_2952);
nor UO_356 (O_356,N_2769,N_2030);
nand UO_357 (O_357,N_2024,N_2465);
and UO_358 (O_358,N_2185,N_2372);
and UO_359 (O_359,N_2665,N_2141);
nand UO_360 (O_360,N_2748,N_2282);
and UO_361 (O_361,N_2832,N_2107);
or UO_362 (O_362,N_2329,N_2468);
and UO_363 (O_363,N_2857,N_2544);
and UO_364 (O_364,N_2888,N_2767);
nand UO_365 (O_365,N_2565,N_2691);
nor UO_366 (O_366,N_2129,N_2593);
nand UO_367 (O_367,N_2273,N_2442);
nand UO_368 (O_368,N_2718,N_2701);
or UO_369 (O_369,N_2373,N_2262);
nor UO_370 (O_370,N_2346,N_2618);
and UO_371 (O_371,N_2524,N_2411);
nor UO_372 (O_372,N_2361,N_2727);
nand UO_373 (O_373,N_2977,N_2434);
and UO_374 (O_374,N_2239,N_2311);
or UO_375 (O_375,N_2447,N_2122);
and UO_376 (O_376,N_2304,N_2766);
nand UO_377 (O_377,N_2683,N_2031);
and UO_378 (O_378,N_2108,N_2595);
and UO_379 (O_379,N_2673,N_2481);
or UO_380 (O_380,N_2886,N_2573);
or UO_381 (O_381,N_2560,N_2153);
nor UO_382 (O_382,N_2341,N_2457);
nand UO_383 (O_383,N_2621,N_2994);
or UO_384 (O_384,N_2280,N_2035);
and UO_385 (O_385,N_2762,N_2313);
or UO_386 (O_386,N_2482,N_2049);
nand UO_387 (O_387,N_2286,N_2756);
nand UO_388 (O_388,N_2935,N_2817);
and UO_389 (O_389,N_2605,N_2427);
nand UO_390 (O_390,N_2084,N_2028);
and UO_391 (O_391,N_2550,N_2677);
nor UO_392 (O_392,N_2312,N_2464);
nand UO_393 (O_393,N_2858,N_2097);
and UO_394 (O_394,N_2494,N_2978);
or UO_395 (O_395,N_2714,N_2435);
or UO_396 (O_396,N_2774,N_2446);
and UO_397 (O_397,N_2450,N_2864);
nand UO_398 (O_398,N_2171,N_2258);
nor UO_399 (O_399,N_2812,N_2757);
and UO_400 (O_400,N_2266,N_2848);
or UO_401 (O_401,N_2559,N_2737);
and UO_402 (O_402,N_2246,N_2080);
or UO_403 (O_403,N_2698,N_2795);
nor UO_404 (O_404,N_2587,N_2695);
nand UO_405 (O_405,N_2635,N_2364);
xor UO_406 (O_406,N_2745,N_2360);
or UO_407 (O_407,N_2268,N_2980);
nor UO_408 (O_408,N_2510,N_2874);
nand UO_409 (O_409,N_2800,N_2314);
nand UO_410 (O_410,N_2706,N_2353);
nor UO_411 (O_411,N_2162,N_2525);
nor UO_412 (O_412,N_2517,N_2571);
or UO_413 (O_413,N_2890,N_2251);
or UO_414 (O_414,N_2908,N_2406);
nand UO_415 (O_415,N_2339,N_2476);
or UO_416 (O_416,N_2984,N_2195);
or UO_417 (O_417,N_2682,N_2551);
nor UO_418 (O_418,N_2421,N_2222);
nand UO_419 (O_419,N_2138,N_2783);
or UO_420 (O_420,N_2590,N_2776);
or UO_421 (O_421,N_2717,N_2441);
and UO_422 (O_422,N_2940,N_2724);
or UO_423 (O_423,N_2506,N_2859);
nand UO_424 (O_424,N_2513,N_2290);
nand UO_425 (O_425,N_2708,N_2430);
or UO_426 (O_426,N_2807,N_2699);
nand UO_427 (O_427,N_2900,N_2733);
nand UO_428 (O_428,N_2998,N_2909);
nor UO_429 (O_429,N_2606,N_2211);
or UO_430 (O_430,N_2969,N_2771);
and UO_431 (O_431,N_2134,N_2170);
nor UO_432 (O_432,N_2690,N_2192);
and UO_433 (O_433,N_2223,N_2221);
nand UO_434 (O_434,N_2444,N_2244);
or UO_435 (O_435,N_2236,N_2955);
or UO_436 (O_436,N_2966,N_2599);
nand UO_437 (O_437,N_2414,N_2489);
or UO_438 (O_438,N_2949,N_2972);
nor UO_439 (O_439,N_2694,N_2113);
or UO_440 (O_440,N_2451,N_2898);
and UO_441 (O_441,N_2088,N_2068);
and UO_442 (O_442,N_2378,N_2274);
and UO_443 (O_443,N_2109,N_2543);
and UO_444 (O_444,N_2316,N_2582);
and UO_445 (O_445,N_2278,N_2472);
or UO_446 (O_446,N_2825,N_2309);
nand UO_447 (O_447,N_2499,N_2400);
nor UO_448 (O_448,N_2975,N_2607);
nand UO_449 (O_449,N_2730,N_2382);
xnor UO_450 (O_450,N_2603,N_2306);
and UO_451 (O_451,N_2105,N_2982);
nand UO_452 (O_452,N_2663,N_2658);
nor UO_453 (O_453,N_2038,N_2877);
nand UO_454 (O_454,N_2040,N_2782);
nand UO_455 (O_455,N_2760,N_2102);
and UO_456 (O_456,N_2487,N_2826);
nor UO_457 (O_457,N_2100,N_2561);
nor UO_458 (O_458,N_2953,N_2894);
nand UO_459 (O_459,N_2905,N_2495);
and UO_460 (O_460,N_2505,N_2139);
nor UO_461 (O_461,N_2248,N_2322);
and UO_462 (O_462,N_2023,N_2799);
or UO_463 (O_463,N_2555,N_2779);
or UO_464 (O_464,N_2512,N_2670);
or UO_465 (O_465,N_2326,N_2189);
or UO_466 (O_466,N_2996,N_2657);
and UO_467 (O_467,N_2791,N_2292);
and UO_468 (O_468,N_2615,N_2648);
or UO_469 (O_469,N_2064,N_2981);
xor UO_470 (O_470,N_2833,N_2073);
nand UO_471 (O_471,N_2074,N_2269);
nor UO_472 (O_472,N_2296,N_2602);
or UO_473 (O_473,N_2726,N_2668);
or UO_474 (O_474,N_2085,N_2526);
nand UO_475 (O_475,N_2591,N_2507);
or UO_476 (O_476,N_2855,N_2240);
nand UO_477 (O_477,N_2787,N_2279);
xnor UO_478 (O_478,N_2385,N_2638);
nand UO_479 (O_479,N_2871,N_2963);
and UO_480 (O_480,N_2226,N_2738);
nor UO_481 (O_481,N_2365,N_2768);
or UO_482 (O_482,N_2458,N_2811);
and UO_483 (O_483,N_2330,N_2865);
nand UO_484 (O_484,N_2432,N_2916);
and UO_485 (O_485,N_2912,N_2887);
nand UO_486 (O_486,N_2794,N_2569);
or UO_487 (O_487,N_2052,N_2856);
nand UO_488 (O_488,N_2893,N_2709);
nor UO_489 (O_489,N_2644,N_2034);
and UO_490 (O_490,N_2132,N_2954);
nand UO_491 (O_491,N_2847,N_2461);
and UO_492 (O_492,N_2103,N_2568);
nand UO_493 (O_493,N_2303,N_2250);
xnor UO_494 (O_494,N_2019,N_2711);
nor UO_495 (O_495,N_2187,N_2376);
and UO_496 (O_496,N_2662,N_2163);
and UO_497 (O_497,N_2722,N_2173);
or UO_498 (O_498,N_2671,N_2588);
or UO_499 (O_499,N_2277,N_2081);
endmodule