module basic_750_5000_1000_2_levels_1xor_4(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2502,N_2503,N_2504,N_2506,N_2507,N_2508,N_2510,N_2511,N_2512,N_2513,N_2514,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2572,N_2574,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2591,N_2592,N_2593,N_2595,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2609,N_2610,N_2611,N_2612,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2639,N_2640,N_2643,N_2648,N_2649,N_2650,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2664,N_2665,N_2666,N_2667,N_2670,N_2671,N_2672,N_2674,N_2675,N_2676,N_2677,N_2678,N_2680,N_2682,N_2683,N_2684,N_2685,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2715,N_2716,N_2717,N_2719,N_2721,N_2722,N_2723,N_2724,N_2726,N_2727,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2745,N_2746,N_2748,N_2753,N_2755,N_2756,N_2758,N_2759,N_2760,N_2762,N_2764,N_2765,N_2767,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2777,N_2779,N_2780,N_2781,N_2782,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2792,N_2793,N_2795,N_2796,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2806,N_2807,N_2808,N_2810,N_2811,N_2812,N_2813,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2835,N_2836,N_2839,N_2840,N_2842,N_2843,N_2844,N_2845,N_2847,N_2848,N_2850,N_2852,N_2854,N_2856,N_2857,N_2859,N_2860,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2883,N_2888,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2902,N_2904,N_2905,N_2906,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2922,N_2924,N_2926,N_2927,N_2928,N_2929,N_2930,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2939,N_2940,N_2941,N_2944,N_2945,N_2946,N_2948,N_2949,N_2950,N_2951,N_2952,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2965,N_2967,N_2968,N_2969,N_2970,N_2972,N_2978,N_2980,N_2981,N_2982,N_2983,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3015,N_3016,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3027,N_3028,N_3029,N_3030,N_3031,N_3033,N_3034,N_3039,N_3040,N_3041,N_3042,N_3044,N_3045,N_3046,N_3047,N_3049,N_3050,N_3051,N_3052,N_3053,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3078,N_3081,N_3083,N_3084,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3096,N_3098,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3107,N_3108,N_3109,N_3110,N_3111,N_3114,N_3115,N_3116,N_3118,N_3120,N_3122,N_3123,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3133,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3145,N_3146,N_3148,N_3149,N_3150,N_3152,N_3153,N_3154,N_3158,N_3159,N_3161,N_3162,N_3163,N_3164,N_3165,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3174,N_3175,N_3176,N_3177,N_3178,N_3180,N_3181,N_3182,N_3183,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3211,N_3212,N_3213,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3237,N_3238,N_3239,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3256,N_3257,N_3259,N_3260,N_3261,N_3262,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3279,N_3280,N_3281,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3291,N_3292,N_3293,N_3294,N_3296,N_3298,N_3300,N_3301,N_3303,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3328,N_3329,N_3330,N_3331,N_3332,N_3335,N_3336,N_3337,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3347,N_3348,N_3349,N_3350,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3394,N_3395,N_3396,N_3397,N_3398,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3407,N_3408,N_3409,N_3411,N_3412,N_3415,N_3416,N_3417,N_3418,N_3421,N_3422,N_3423,N_3425,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3434,N_3436,N_3437,N_3438,N_3440,N_3441,N_3442,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3456,N_3457,N_3458,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3478,N_3479,N_3481,N_3483,N_3484,N_3486,N_3487,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3517,N_3518,N_3519,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3535,N_3538,N_3539,N_3540,N_3542,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3552,N_3553,N_3554,N_3555,N_3557,N_3558,N_3559,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3592,N_3593,N_3594,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3612,N_3614,N_3616,N_3617,N_3618,N_3619,N_3620,N_3623,N_3624,N_3625,N_3627,N_3629,N_3630,N_3631,N_3632,N_3633,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3643,N_3644,N_3646,N_3648,N_3649,N_3650,N_3652,N_3653,N_3654,N_3655,N_3657,N_3658,N_3659,N_3660,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3669,N_3670,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3680,N_3682,N_3683,N_3686,N_3687,N_3688,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3704,N_3705,N_3706,N_3707,N_3708,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3720,N_3721,N_3722,N_3723,N_3724,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3748,N_3750,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3760,N_3761,N_3762,N_3763,N_3765,N_3766,N_3767,N_3769,N_3770,N_3771,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3781,N_3782,N_3783,N_3784,N_3785,N_3787,N_3788,N_3790,N_3791,N_3792,N_3793,N_3796,N_3797,N_3798,N_3799,N_3800,N_3802,N_3803,N_3805,N_3806,N_3807,N_3808,N_3809,N_3811,N_3812,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3823,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3837,N_3838,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3851,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3861,N_3863,N_3864,N_3865,N_3866,N_3867,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3879,N_3881,N_3882,N_3883,N_3885,N_3887,N_3888,N_3889,N_3890,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3904,N_3905,N_3906,N_3907,N_3909,N_3910,N_3911,N_3913,N_3914,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3925,N_3926,N_3927,N_3932,N_3933,N_3935,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3969,N_3970,N_3972,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4006,N_4007,N_4008,N_4009,N_4010,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4038,N_4039,N_4040,N_4041,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4073,N_4074,N_4075,N_4077,N_4078,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4089,N_4090,N_4091,N_4093,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4104,N_4106,N_4108,N_4109,N_4111,N_4112,N_4113,N_4115,N_4116,N_4117,N_4118,N_4120,N_4121,N_4122,N_4124,N_4125,N_4126,N_4127,N_4128,N_4131,N_4134,N_4135,N_4137,N_4138,N_4139,N_4142,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4151,N_4153,N_4154,N_4155,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4193,N_4194,N_4195,N_4196,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4238,N_4239,N_4241,N_4242,N_4243,N_4245,N_4246,N_4248,N_4249,N_4250,N_4251,N_4253,N_4254,N_4256,N_4257,N_4258,N_4259,N_4260,N_4263,N_4265,N_4266,N_4267,N_4269,N_4270,N_4273,N_4274,N_4275,N_4276,N_4277,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4287,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4308,N_4309,N_4310,N_4311,N_4312,N_4314,N_4317,N_4318,N_4319,N_4320,N_4321,N_4323,N_4325,N_4326,N_4327,N_4328,N_4329,N_4331,N_4333,N_4334,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4353,N_4354,N_4355,N_4356,N_4357,N_4359,N_4360,N_4361,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4377,N_4378,N_4379,N_4382,N_4384,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4400,N_4401,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4411,N_4412,N_4413,N_4414,N_4415,N_4417,N_4418,N_4419,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4428,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4456,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4480,N_4482,N_4485,N_4487,N_4488,N_4489,N_4491,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4510,N_4511,N_4513,N_4514,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4532,N_4533,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4550,N_4551,N_4552,N_4553,N_4554,N_4556,N_4557,N_4558,N_4559,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4575,N_4576,N_4577,N_4579,N_4580,N_4581,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4591,N_4592,N_4593,N_4595,N_4596,N_4597,N_4600,N_4601,N_4602,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4621,N_4623,N_4624,N_4625,N_4627,N_4628,N_4629,N_4630,N_4631,N_4633,N_4634,N_4635,N_4637,N_4638,N_4639,N_4641,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4652,N_4653,N_4655,N_4656,N_4657,N_4658,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4670,N_4671,N_4672,N_4673,N_4674,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4708,N_4709,N_4710,N_4711,N_4712,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4774,N_4776,N_4777,N_4778,N_4779,N_4780,N_4782,N_4784,N_4786,N_4787,N_4789,N_4790,N_4791,N_4792,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4813,N_4815,N_4816,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4838,N_4839,N_4841,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4868,N_4869,N_4872,N_4874,N_4875,N_4876,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4901,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4919,N_4920,N_4921,N_4922,N_4923,N_4925,N_4926,N_4927,N_4929,N_4930,N_4931,N_4932,N_4934,N_4935,N_4937,N_4938,N_4939,N_4940,N_4942,N_4943,N_4944,N_4945,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4996,N_4998,N_4999;
nand U0 (N_0,In_61,In_183);
nor U1 (N_1,In_224,In_419);
and U2 (N_2,In_401,In_89);
or U3 (N_3,In_362,In_473);
or U4 (N_4,In_3,In_51);
nand U5 (N_5,In_37,In_454);
and U6 (N_6,In_319,In_619);
nor U7 (N_7,In_602,In_153);
and U8 (N_8,In_110,In_517);
xnor U9 (N_9,In_239,In_451);
and U10 (N_10,In_625,In_570);
or U11 (N_11,In_68,In_450);
nor U12 (N_12,In_680,In_485);
nand U13 (N_13,In_399,In_283);
nand U14 (N_14,In_242,In_638);
and U15 (N_15,In_18,In_585);
nand U16 (N_16,In_115,In_346);
nand U17 (N_17,In_17,In_439);
and U18 (N_18,In_371,In_344);
and U19 (N_19,In_112,In_216);
nand U20 (N_20,In_238,In_103);
or U21 (N_21,In_578,In_706);
nor U22 (N_22,In_181,In_489);
and U23 (N_23,In_222,In_257);
or U24 (N_24,In_11,In_174);
xnor U25 (N_25,In_562,In_219);
nor U26 (N_26,In_210,In_65);
nand U27 (N_27,In_526,In_46);
nand U28 (N_28,In_621,In_298);
nand U29 (N_29,In_447,In_465);
or U30 (N_30,In_415,In_47);
or U31 (N_31,In_540,In_285);
nor U32 (N_32,In_329,In_354);
nor U33 (N_33,In_8,In_280);
or U34 (N_34,In_220,In_566);
or U35 (N_35,In_295,In_207);
and U36 (N_36,In_708,In_171);
xnor U37 (N_37,In_116,In_406);
or U38 (N_38,In_700,In_312);
and U39 (N_39,In_507,In_311);
and U40 (N_40,In_471,In_350);
and U41 (N_41,In_626,In_321);
nand U42 (N_42,In_133,In_263);
or U43 (N_43,In_552,In_452);
nor U44 (N_44,In_376,In_327);
nand U45 (N_45,In_16,In_460);
or U46 (N_46,In_577,In_728);
or U47 (N_47,In_688,In_237);
and U48 (N_48,In_564,In_482);
nand U49 (N_49,In_109,In_325);
and U50 (N_50,In_78,In_208);
nor U51 (N_51,In_330,In_685);
nor U52 (N_52,In_179,In_256);
or U53 (N_53,In_666,In_333);
or U54 (N_54,In_521,In_90);
and U55 (N_55,In_52,In_611);
and U56 (N_56,In_710,In_353);
and U57 (N_57,In_199,In_259);
and U58 (N_58,In_593,In_313);
or U59 (N_59,In_273,In_212);
or U60 (N_60,In_387,In_424);
nand U61 (N_61,In_433,In_122);
and U62 (N_62,In_294,In_572);
or U63 (N_63,In_206,In_410);
and U64 (N_64,In_262,In_217);
or U65 (N_65,In_745,In_48);
or U66 (N_66,In_718,In_504);
or U67 (N_67,In_658,In_200);
or U68 (N_68,In_605,In_495);
nor U69 (N_69,In_691,In_701);
or U70 (N_70,In_98,In_719);
nand U71 (N_71,In_240,In_36);
xnor U72 (N_72,In_286,In_185);
or U73 (N_73,In_443,In_738);
or U74 (N_74,In_165,In_339);
nor U75 (N_75,In_15,In_25);
or U76 (N_76,In_129,In_631);
nor U77 (N_77,In_277,In_628);
nand U78 (N_78,In_657,In_723);
or U79 (N_79,In_522,In_104);
nand U80 (N_80,In_656,In_557);
nor U81 (N_81,In_411,In_587);
and U82 (N_82,In_31,In_622);
nor U83 (N_83,In_385,In_43);
nor U84 (N_84,In_612,In_309);
nand U85 (N_85,In_24,In_147);
or U86 (N_86,In_484,In_202);
and U87 (N_87,In_448,In_535);
or U88 (N_88,In_250,In_449);
nand U89 (N_89,In_323,In_604);
xnor U90 (N_90,In_740,In_429);
nor U91 (N_91,In_696,In_393);
or U92 (N_92,In_1,In_427);
and U93 (N_93,In_609,In_440);
and U94 (N_94,In_378,In_154);
or U95 (N_95,In_359,In_170);
nor U96 (N_96,In_500,In_82);
nor U97 (N_97,In_223,In_157);
or U98 (N_98,In_81,In_610);
nand U99 (N_99,In_374,In_391);
or U100 (N_100,In_95,In_652);
and U101 (N_101,In_404,In_35);
and U102 (N_102,In_230,In_514);
and U103 (N_103,In_101,In_388);
nand U104 (N_104,In_458,In_138);
xnor U105 (N_105,In_469,In_508);
nand U106 (N_106,In_152,In_275);
or U107 (N_107,In_664,In_727);
nand U108 (N_108,In_445,In_532);
nor U109 (N_109,In_413,In_107);
nand U110 (N_110,In_747,In_124);
and U111 (N_111,In_204,In_180);
and U112 (N_112,In_169,In_647);
and U113 (N_113,In_697,In_57);
or U114 (N_114,In_714,In_398);
or U115 (N_115,In_466,In_588);
nand U116 (N_116,In_530,In_364);
nor U117 (N_117,In_34,In_307);
nor U118 (N_118,In_118,In_251);
nor U119 (N_119,In_264,In_117);
nor U120 (N_120,In_426,In_565);
nor U121 (N_121,In_474,In_352);
nand U122 (N_122,In_435,In_357);
nand U123 (N_123,In_648,In_113);
nor U124 (N_124,In_580,In_175);
nor U125 (N_125,In_258,In_446);
nor U126 (N_126,In_505,In_608);
nor U127 (N_127,In_316,In_487);
or U128 (N_128,In_67,In_528);
nor U129 (N_129,In_66,In_269);
nand U130 (N_130,In_707,In_550);
nor U131 (N_131,In_100,In_299);
nor U132 (N_132,In_252,In_58);
nand U133 (N_133,In_228,In_246);
xor U134 (N_134,In_637,In_151);
nor U135 (N_135,In_53,In_335);
and U136 (N_136,In_742,In_544);
or U137 (N_137,In_434,In_501);
or U138 (N_138,In_235,In_599);
and U139 (N_139,In_709,In_108);
and U140 (N_140,In_197,In_131);
or U141 (N_141,In_589,In_689);
nand U142 (N_142,In_41,In_372);
or U143 (N_143,In_662,In_59);
and U144 (N_144,In_88,In_678);
or U145 (N_145,In_623,In_29);
nand U146 (N_146,In_649,In_699);
and U147 (N_147,In_60,In_724);
and U148 (N_148,In_314,In_653);
and U149 (N_149,In_145,In_291);
nor U150 (N_150,In_6,In_392);
nand U151 (N_151,In_54,In_615);
and U152 (N_152,In_177,In_594);
and U153 (N_153,In_375,In_584);
xor U154 (N_154,In_83,In_39);
or U155 (N_155,In_492,In_726);
nand U156 (N_156,In_620,In_351);
nand U157 (N_157,In_201,In_749);
nand U158 (N_158,In_496,In_674);
nand U159 (N_159,In_468,In_693);
nor U160 (N_160,In_56,In_360);
nor U161 (N_161,In_293,In_571);
and U162 (N_162,In_568,In_64);
or U163 (N_163,In_270,In_455);
nand U164 (N_164,In_274,In_545);
nor U165 (N_165,In_193,In_28);
or U166 (N_166,In_560,In_698);
or U167 (N_167,In_336,In_267);
nand U168 (N_168,In_310,In_265);
and U169 (N_169,In_515,In_255);
or U170 (N_170,In_337,In_472);
and U171 (N_171,In_630,In_245);
nor U172 (N_172,In_345,In_554);
nor U173 (N_173,In_318,In_10);
nor U174 (N_174,In_462,In_72);
nand U175 (N_175,In_334,In_198);
and U176 (N_176,In_475,In_290);
nand U177 (N_177,In_533,In_668);
and U178 (N_178,In_422,In_397);
and U179 (N_179,In_178,In_559);
or U180 (N_180,In_470,In_73);
and U181 (N_181,In_272,In_244);
nor U182 (N_182,In_420,In_695);
xor U183 (N_183,In_494,In_320);
or U184 (N_184,In_45,In_386);
and U185 (N_185,In_643,In_687);
nor U186 (N_186,In_677,In_137);
nor U187 (N_187,In_590,In_93);
nor U188 (N_188,In_21,In_644);
or U189 (N_189,In_720,In_69);
and U190 (N_190,In_195,In_407);
nand U191 (N_191,In_624,In_87);
and U192 (N_192,In_736,In_479);
or U193 (N_193,In_191,In_158);
nand U194 (N_194,In_159,In_326);
and U195 (N_195,In_384,In_729);
nor U196 (N_196,In_205,In_671);
or U197 (N_197,In_261,In_534);
or U198 (N_198,In_414,In_498);
nor U199 (N_199,In_132,In_84);
nor U200 (N_200,In_490,In_324);
nand U201 (N_201,In_189,In_79);
and U202 (N_202,In_600,In_9);
and U203 (N_203,In_85,In_349);
or U204 (N_204,In_97,In_548);
or U205 (N_205,In_213,In_614);
nor U206 (N_206,In_395,In_305);
nand U207 (N_207,In_308,In_70);
or U208 (N_208,In_394,In_513);
or U209 (N_209,In_128,In_231);
nand U210 (N_210,In_527,In_659);
or U211 (N_211,In_425,In_144);
nand U212 (N_212,In_381,In_338);
or U213 (N_213,In_493,In_176);
and U214 (N_214,In_13,In_403);
and U215 (N_215,In_77,In_168);
or U216 (N_216,In_681,In_423);
nor U217 (N_217,In_408,In_187);
or U218 (N_218,In_497,In_721);
or U219 (N_219,In_667,In_591);
nor U220 (N_220,In_597,In_106);
and U221 (N_221,In_412,In_182);
and U222 (N_222,In_567,In_303);
nand U223 (N_223,In_221,In_188);
or U224 (N_224,In_289,In_725);
nand U225 (N_225,In_711,In_369);
or U226 (N_226,In_276,In_739);
nor U227 (N_227,In_682,In_607);
or U228 (N_228,In_30,In_102);
or U229 (N_229,In_486,In_86);
nand U230 (N_230,In_531,In_746);
or U231 (N_231,In_120,In_543);
and U232 (N_232,In_389,In_382);
or U233 (N_233,In_190,In_260);
or U234 (N_234,In_601,In_617);
and U235 (N_235,In_478,In_576);
and U236 (N_236,In_71,In_488);
nand U237 (N_237,In_91,In_121);
or U238 (N_238,In_672,In_156);
and U239 (N_239,In_524,In_33);
and U240 (N_240,In_126,In_733);
or U241 (N_241,In_430,In_322);
and U242 (N_242,In_379,In_483);
xnor U243 (N_243,In_75,In_538);
or U244 (N_244,In_511,In_111);
and U245 (N_245,In_315,In_537);
and U246 (N_246,In_227,In_341);
or U247 (N_247,In_661,In_287);
or U248 (N_248,In_186,In_373);
or U249 (N_249,In_5,In_744);
or U250 (N_250,In_347,In_49);
nand U251 (N_251,In_491,In_639);
and U252 (N_252,In_139,In_119);
or U253 (N_253,In_301,In_634);
nor U254 (N_254,In_225,In_266);
nand U255 (N_255,In_99,In_380);
or U256 (N_256,In_467,In_400);
xor U257 (N_257,In_383,In_402);
or U258 (N_258,In_140,In_660);
nand U259 (N_259,In_651,In_510);
nor U260 (N_260,In_163,In_670);
or U261 (N_261,In_236,In_343);
and U262 (N_262,In_583,In_509);
or U263 (N_263,In_282,In_632);
or U264 (N_264,In_172,In_2);
xor U265 (N_265,In_683,In_92);
nand U266 (N_266,In_713,In_271);
nand U267 (N_267,In_141,In_722);
or U268 (N_268,In_123,In_536);
and U269 (N_269,In_355,In_457);
nor U270 (N_270,In_14,In_167);
or U271 (N_271,In_367,In_731);
nor U272 (N_272,In_22,In_686);
and U273 (N_273,In_253,In_542);
nand U274 (N_274,In_692,In_541);
nor U275 (N_275,In_248,In_748);
nor U276 (N_276,In_629,In_569);
nand U277 (N_277,In_421,In_241);
or U278 (N_278,In_23,In_300);
nor U279 (N_279,In_641,In_431);
nand U280 (N_280,In_50,In_476);
and U281 (N_281,In_125,In_438);
nor U282 (N_282,In_32,In_716);
nand U283 (N_283,In_645,In_613);
nand U284 (N_284,In_636,In_409);
and U285 (N_285,In_684,In_646);
and U286 (N_286,In_616,In_563);
or U287 (N_287,In_436,In_42);
nand U288 (N_288,In_20,In_377);
and U289 (N_289,In_214,In_456);
nand U290 (N_290,In_80,In_665);
and U291 (N_291,In_342,In_592);
or U292 (N_292,In_734,In_650);
nand U293 (N_293,In_302,In_676);
nand U294 (N_294,In_161,In_633);
or U295 (N_295,In_55,In_136);
or U296 (N_296,In_365,In_390);
nand U297 (N_297,In_243,In_441);
and U298 (N_298,In_453,In_94);
nand U299 (N_299,In_673,In_627);
and U300 (N_300,In_477,In_209);
or U301 (N_301,In_574,In_503);
or U302 (N_302,In_12,In_297);
or U303 (N_303,In_558,In_268);
nor U304 (N_304,In_328,In_194);
or U305 (N_305,In_366,In_553);
nor U306 (N_306,In_595,In_26);
or U307 (N_307,In_361,In_135);
nor U308 (N_308,In_155,In_704);
and U309 (N_309,In_368,In_655);
or U310 (N_310,In_164,In_654);
and U311 (N_311,In_428,In_288);
nand U312 (N_312,In_292,In_596);
nand U313 (N_313,In_506,In_481);
or U314 (N_314,In_735,In_418);
nor U315 (N_315,In_598,In_586);
nand U316 (N_316,In_203,In_520);
and U317 (N_317,In_134,In_279);
and U318 (N_318,In_730,In_743);
or U319 (N_319,In_281,In_127);
nand U320 (N_320,In_226,In_499);
nand U321 (N_321,In_254,In_249);
or U322 (N_322,In_442,In_705);
nand U323 (N_323,In_7,In_675);
or U324 (N_324,In_40,In_332);
and U325 (N_325,In_459,In_546);
or U326 (N_326,In_192,In_306);
and U327 (N_327,In_732,In_148);
or U328 (N_328,In_27,In_444);
nand U329 (N_329,In_166,In_464);
nand U330 (N_330,In_396,In_150);
nor U331 (N_331,In_370,In_74);
nor U332 (N_332,In_19,In_603);
and U333 (N_333,In_502,In_556);
or U334 (N_334,In_173,In_44);
nand U335 (N_335,In_215,In_76);
nor U336 (N_336,In_523,In_38);
and U337 (N_337,In_582,In_284);
and U338 (N_338,In_317,In_715);
and U339 (N_339,In_142,In_331);
and U340 (N_340,In_278,In_463);
and U341 (N_341,In_551,In_184);
nand U342 (N_342,In_561,In_196);
nor U343 (N_343,In_547,In_694);
and U344 (N_344,In_663,In_233);
and U345 (N_345,In_149,In_356);
nor U346 (N_346,In_0,In_737);
nand U347 (N_347,In_512,In_416);
nand U348 (N_348,In_146,In_635);
or U349 (N_349,In_579,In_96);
nand U350 (N_350,In_348,In_304);
nand U351 (N_351,In_437,In_702);
nand U352 (N_352,In_229,In_690);
nand U353 (N_353,In_234,In_575);
and U354 (N_354,In_62,In_105);
and U355 (N_355,In_518,In_679);
nand U356 (N_356,In_480,In_4);
nor U357 (N_357,In_63,In_549);
and U358 (N_358,In_211,In_555);
nor U359 (N_359,In_461,In_640);
and U360 (N_360,In_218,In_405);
nand U361 (N_361,In_296,In_581);
and U362 (N_362,In_717,In_130);
nand U363 (N_363,In_539,In_232);
and U364 (N_364,In_358,In_642);
nor U365 (N_365,In_712,In_432);
and U366 (N_366,In_525,In_519);
or U367 (N_367,In_247,In_669);
or U368 (N_368,In_162,In_160);
and U369 (N_369,In_573,In_340);
and U370 (N_370,In_114,In_703);
or U371 (N_371,In_143,In_741);
nand U372 (N_372,In_618,In_529);
and U373 (N_373,In_417,In_516);
nand U374 (N_374,In_363,In_606);
and U375 (N_375,In_101,In_651);
nand U376 (N_376,In_297,In_221);
or U377 (N_377,In_31,In_260);
nand U378 (N_378,In_174,In_500);
nor U379 (N_379,In_292,In_66);
and U380 (N_380,In_296,In_611);
nor U381 (N_381,In_295,In_569);
and U382 (N_382,In_29,In_105);
and U383 (N_383,In_349,In_27);
or U384 (N_384,In_457,In_539);
nand U385 (N_385,In_741,In_619);
and U386 (N_386,In_738,In_489);
nand U387 (N_387,In_363,In_575);
nor U388 (N_388,In_195,In_348);
nor U389 (N_389,In_670,In_314);
and U390 (N_390,In_582,In_690);
and U391 (N_391,In_108,In_676);
nor U392 (N_392,In_640,In_705);
and U393 (N_393,In_645,In_406);
nor U394 (N_394,In_327,In_388);
nand U395 (N_395,In_631,In_264);
nand U396 (N_396,In_102,In_268);
or U397 (N_397,In_243,In_456);
nand U398 (N_398,In_472,In_718);
nor U399 (N_399,In_55,In_307);
xnor U400 (N_400,In_525,In_518);
or U401 (N_401,In_384,In_340);
nand U402 (N_402,In_192,In_421);
nor U403 (N_403,In_601,In_162);
nor U404 (N_404,In_72,In_46);
nand U405 (N_405,In_535,In_37);
or U406 (N_406,In_731,In_327);
or U407 (N_407,In_139,In_150);
nand U408 (N_408,In_207,In_503);
nor U409 (N_409,In_646,In_355);
nand U410 (N_410,In_529,In_534);
nor U411 (N_411,In_658,In_414);
or U412 (N_412,In_484,In_13);
and U413 (N_413,In_612,In_75);
nor U414 (N_414,In_398,In_414);
and U415 (N_415,In_33,In_6);
and U416 (N_416,In_686,In_284);
or U417 (N_417,In_708,In_232);
and U418 (N_418,In_499,In_203);
or U419 (N_419,In_289,In_599);
nand U420 (N_420,In_269,In_444);
nor U421 (N_421,In_544,In_355);
nor U422 (N_422,In_556,In_499);
or U423 (N_423,In_574,In_141);
nand U424 (N_424,In_491,In_649);
or U425 (N_425,In_263,In_734);
nor U426 (N_426,In_326,In_445);
nor U427 (N_427,In_421,In_425);
or U428 (N_428,In_542,In_448);
nor U429 (N_429,In_538,In_158);
nand U430 (N_430,In_444,In_368);
xnor U431 (N_431,In_410,In_27);
nand U432 (N_432,In_676,In_400);
nand U433 (N_433,In_219,In_386);
or U434 (N_434,In_446,In_102);
nor U435 (N_435,In_468,In_451);
nor U436 (N_436,In_716,In_171);
nand U437 (N_437,In_690,In_443);
nand U438 (N_438,In_254,In_699);
or U439 (N_439,In_687,In_491);
nor U440 (N_440,In_127,In_132);
nor U441 (N_441,In_664,In_142);
nand U442 (N_442,In_98,In_607);
and U443 (N_443,In_30,In_172);
nand U444 (N_444,In_722,In_78);
or U445 (N_445,In_262,In_745);
and U446 (N_446,In_566,In_369);
nand U447 (N_447,In_583,In_184);
nand U448 (N_448,In_54,In_584);
nor U449 (N_449,In_194,In_428);
nand U450 (N_450,In_157,In_249);
nor U451 (N_451,In_439,In_615);
nor U452 (N_452,In_224,In_68);
nand U453 (N_453,In_18,In_214);
and U454 (N_454,In_683,In_679);
and U455 (N_455,In_347,In_21);
or U456 (N_456,In_622,In_10);
nand U457 (N_457,In_372,In_480);
xor U458 (N_458,In_40,In_4);
nor U459 (N_459,In_706,In_84);
nand U460 (N_460,In_97,In_637);
and U461 (N_461,In_626,In_109);
or U462 (N_462,In_299,In_546);
nor U463 (N_463,In_62,In_148);
nand U464 (N_464,In_118,In_218);
or U465 (N_465,In_675,In_409);
and U466 (N_466,In_56,In_630);
and U467 (N_467,In_648,In_613);
nor U468 (N_468,In_493,In_382);
nor U469 (N_469,In_316,In_90);
nand U470 (N_470,In_62,In_662);
and U471 (N_471,In_389,In_673);
nor U472 (N_472,In_725,In_685);
nand U473 (N_473,In_281,In_384);
or U474 (N_474,In_566,In_93);
nand U475 (N_475,In_80,In_710);
nand U476 (N_476,In_241,In_447);
and U477 (N_477,In_623,In_397);
and U478 (N_478,In_438,In_22);
and U479 (N_479,In_219,In_202);
and U480 (N_480,In_90,In_287);
or U481 (N_481,In_471,In_137);
nand U482 (N_482,In_104,In_333);
nand U483 (N_483,In_604,In_60);
nand U484 (N_484,In_70,In_748);
nand U485 (N_485,In_84,In_599);
and U486 (N_486,In_627,In_747);
or U487 (N_487,In_368,In_356);
nor U488 (N_488,In_85,In_153);
and U489 (N_489,In_330,In_506);
and U490 (N_490,In_610,In_188);
nand U491 (N_491,In_223,In_138);
or U492 (N_492,In_298,In_322);
or U493 (N_493,In_674,In_26);
nand U494 (N_494,In_60,In_422);
nor U495 (N_495,In_147,In_740);
nor U496 (N_496,In_194,In_329);
nand U497 (N_497,In_559,In_177);
nor U498 (N_498,In_144,In_107);
or U499 (N_499,In_180,In_107);
and U500 (N_500,In_376,In_222);
and U501 (N_501,In_121,In_160);
nor U502 (N_502,In_43,In_279);
nor U503 (N_503,In_367,In_72);
or U504 (N_504,In_720,In_40);
nor U505 (N_505,In_447,In_155);
xnor U506 (N_506,In_478,In_511);
and U507 (N_507,In_45,In_619);
or U508 (N_508,In_697,In_394);
nor U509 (N_509,In_171,In_242);
nand U510 (N_510,In_571,In_693);
or U511 (N_511,In_675,In_329);
or U512 (N_512,In_738,In_115);
nor U513 (N_513,In_530,In_586);
and U514 (N_514,In_524,In_194);
xnor U515 (N_515,In_288,In_711);
nand U516 (N_516,In_212,In_282);
or U517 (N_517,In_251,In_41);
nand U518 (N_518,In_567,In_82);
xor U519 (N_519,In_567,In_215);
nor U520 (N_520,In_244,In_112);
or U521 (N_521,In_579,In_260);
nor U522 (N_522,In_137,In_574);
nor U523 (N_523,In_564,In_271);
nor U524 (N_524,In_689,In_189);
and U525 (N_525,In_272,In_270);
nor U526 (N_526,In_245,In_36);
and U527 (N_527,In_505,In_484);
or U528 (N_528,In_371,In_513);
and U529 (N_529,In_577,In_294);
and U530 (N_530,In_148,In_338);
nor U531 (N_531,In_592,In_150);
and U532 (N_532,In_463,In_500);
nor U533 (N_533,In_503,In_488);
nor U534 (N_534,In_416,In_79);
or U535 (N_535,In_720,In_234);
nor U536 (N_536,In_238,In_447);
nand U537 (N_537,In_296,In_470);
or U538 (N_538,In_50,In_309);
nor U539 (N_539,In_546,In_198);
nor U540 (N_540,In_341,In_569);
xor U541 (N_541,In_529,In_383);
or U542 (N_542,In_535,In_153);
nor U543 (N_543,In_275,In_308);
or U544 (N_544,In_269,In_441);
nand U545 (N_545,In_500,In_98);
nand U546 (N_546,In_117,In_166);
and U547 (N_547,In_480,In_7);
nand U548 (N_548,In_490,In_395);
or U549 (N_549,In_493,In_113);
or U550 (N_550,In_723,In_686);
nor U551 (N_551,In_441,In_55);
and U552 (N_552,In_131,In_65);
or U553 (N_553,In_59,In_199);
and U554 (N_554,In_439,In_556);
nor U555 (N_555,In_735,In_420);
or U556 (N_556,In_198,In_589);
and U557 (N_557,In_62,In_93);
and U558 (N_558,In_672,In_52);
nand U559 (N_559,In_365,In_199);
and U560 (N_560,In_494,In_327);
nor U561 (N_561,In_716,In_341);
and U562 (N_562,In_671,In_173);
or U563 (N_563,In_463,In_324);
nor U564 (N_564,In_248,In_716);
or U565 (N_565,In_174,In_316);
and U566 (N_566,In_184,In_378);
nor U567 (N_567,In_187,In_569);
nor U568 (N_568,In_232,In_44);
and U569 (N_569,In_574,In_195);
and U570 (N_570,In_450,In_729);
or U571 (N_571,In_724,In_198);
nor U572 (N_572,In_146,In_503);
nor U573 (N_573,In_364,In_244);
nor U574 (N_574,In_255,In_72);
and U575 (N_575,In_23,In_421);
and U576 (N_576,In_199,In_285);
and U577 (N_577,In_616,In_510);
nor U578 (N_578,In_298,In_257);
nand U579 (N_579,In_214,In_181);
nor U580 (N_580,In_204,In_144);
or U581 (N_581,In_603,In_18);
nand U582 (N_582,In_618,In_98);
nand U583 (N_583,In_705,In_630);
or U584 (N_584,In_349,In_151);
nand U585 (N_585,In_656,In_713);
nand U586 (N_586,In_24,In_94);
nand U587 (N_587,In_39,In_297);
nand U588 (N_588,In_22,In_143);
nand U589 (N_589,In_431,In_65);
nand U590 (N_590,In_594,In_361);
nand U591 (N_591,In_170,In_409);
or U592 (N_592,In_12,In_714);
or U593 (N_593,In_182,In_366);
nor U594 (N_594,In_246,In_661);
nor U595 (N_595,In_294,In_543);
nand U596 (N_596,In_580,In_97);
or U597 (N_597,In_658,In_205);
nand U598 (N_598,In_502,In_712);
nor U599 (N_599,In_322,In_338);
nor U600 (N_600,In_650,In_186);
or U601 (N_601,In_208,In_362);
and U602 (N_602,In_576,In_152);
nor U603 (N_603,In_513,In_169);
nor U604 (N_604,In_564,In_719);
nand U605 (N_605,In_385,In_481);
nor U606 (N_606,In_481,In_729);
nand U607 (N_607,In_135,In_631);
nand U608 (N_608,In_295,In_711);
and U609 (N_609,In_695,In_739);
nor U610 (N_610,In_401,In_395);
nor U611 (N_611,In_670,In_351);
and U612 (N_612,In_241,In_730);
nor U613 (N_613,In_102,In_587);
and U614 (N_614,In_209,In_238);
and U615 (N_615,In_113,In_92);
or U616 (N_616,In_614,In_528);
and U617 (N_617,In_665,In_286);
or U618 (N_618,In_742,In_313);
or U619 (N_619,In_548,In_306);
nor U620 (N_620,In_518,In_106);
or U621 (N_621,In_56,In_327);
nor U622 (N_622,In_383,In_274);
or U623 (N_623,In_162,In_134);
and U624 (N_624,In_688,In_676);
or U625 (N_625,In_317,In_14);
nor U626 (N_626,In_42,In_102);
or U627 (N_627,In_540,In_729);
or U628 (N_628,In_114,In_542);
nor U629 (N_629,In_742,In_219);
nor U630 (N_630,In_479,In_417);
or U631 (N_631,In_95,In_203);
or U632 (N_632,In_354,In_104);
nand U633 (N_633,In_651,In_247);
nand U634 (N_634,In_621,In_314);
nand U635 (N_635,In_653,In_40);
nor U636 (N_636,In_319,In_70);
nor U637 (N_637,In_325,In_419);
nand U638 (N_638,In_358,In_649);
nor U639 (N_639,In_185,In_335);
nor U640 (N_640,In_535,In_292);
xor U641 (N_641,In_305,In_722);
and U642 (N_642,In_641,In_533);
nand U643 (N_643,In_310,In_175);
and U644 (N_644,In_711,In_464);
and U645 (N_645,In_442,In_201);
nand U646 (N_646,In_526,In_476);
nand U647 (N_647,In_402,In_567);
and U648 (N_648,In_598,In_579);
nor U649 (N_649,In_645,In_625);
and U650 (N_650,In_456,In_609);
nor U651 (N_651,In_285,In_717);
or U652 (N_652,In_254,In_618);
and U653 (N_653,In_367,In_51);
and U654 (N_654,In_192,In_697);
nor U655 (N_655,In_21,In_630);
nand U656 (N_656,In_693,In_317);
nand U657 (N_657,In_367,In_405);
and U658 (N_658,In_293,In_705);
and U659 (N_659,In_565,In_223);
and U660 (N_660,In_155,In_365);
nand U661 (N_661,In_436,In_290);
nor U662 (N_662,In_470,In_443);
and U663 (N_663,In_601,In_346);
and U664 (N_664,In_656,In_112);
and U665 (N_665,In_46,In_293);
nand U666 (N_666,In_156,In_198);
and U667 (N_667,In_143,In_7);
nand U668 (N_668,In_534,In_710);
nand U669 (N_669,In_76,In_139);
nor U670 (N_670,In_444,In_318);
nor U671 (N_671,In_34,In_442);
or U672 (N_672,In_579,In_591);
nand U673 (N_673,In_361,In_716);
nor U674 (N_674,In_196,In_233);
and U675 (N_675,In_79,In_433);
nor U676 (N_676,In_563,In_396);
nor U677 (N_677,In_579,In_640);
or U678 (N_678,In_503,In_608);
or U679 (N_679,In_182,In_32);
and U680 (N_680,In_51,In_718);
and U681 (N_681,In_50,In_179);
nor U682 (N_682,In_577,In_13);
nand U683 (N_683,In_344,In_349);
and U684 (N_684,In_91,In_546);
and U685 (N_685,In_637,In_117);
nand U686 (N_686,In_480,In_257);
nand U687 (N_687,In_650,In_612);
and U688 (N_688,In_417,In_263);
nand U689 (N_689,In_739,In_126);
and U690 (N_690,In_409,In_647);
or U691 (N_691,In_607,In_377);
and U692 (N_692,In_229,In_559);
nor U693 (N_693,In_280,In_636);
or U694 (N_694,In_21,In_181);
nor U695 (N_695,In_469,In_370);
or U696 (N_696,In_108,In_302);
and U697 (N_697,In_726,In_654);
or U698 (N_698,In_41,In_565);
nand U699 (N_699,In_276,In_587);
or U700 (N_700,In_443,In_510);
and U701 (N_701,In_54,In_161);
and U702 (N_702,In_228,In_328);
and U703 (N_703,In_62,In_607);
and U704 (N_704,In_71,In_371);
or U705 (N_705,In_524,In_282);
and U706 (N_706,In_395,In_566);
or U707 (N_707,In_348,In_713);
nor U708 (N_708,In_224,In_556);
nand U709 (N_709,In_543,In_734);
and U710 (N_710,In_461,In_436);
and U711 (N_711,In_624,In_302);
nand U712 (N_712,In_170,In_215);
and U713 (N_713,In_496,In_335);
nor U714 (N_714,In_537,In_355);
and U715 (N_715,In_501,In_168);
nand U716 (N_716,In_160,In_230);
nand U717 (N_717,In_294,In_656);
nor U718 (N_718,In_473,In_329);
nor U719 (N_719,In_201,In_70);
or U720 (N_720,In_375,In_627);
nand U721 (N_721,In_138,In_713);
xnor U722 (N_722,In_554,In_577);
nand U723 (N_723,In_189,In_667);
nor U724 (N_724,In_553,In_359);
nor U725 (N_725,In_532,In_605);
nand U726 (N_726,In_14,In_199);
and U727 (N_727,In_218,In_446);
and U728 (N_728,In_682,In_217);
nand U729 (N_729,In_586,In_251);
or U730 (N_730,In_422,In_289);
nor U731 (N_731,In_675,In_628);
and U732 (N_732,In_305,In_220);
or U733 (N_733,In_115,In_146);
and U734 (N_734,In_687,In_461);
and U735 (N_735,In_443,In_22);
nand U736 (N_736,In_259,In_302);
or U737 (N_737,In_521,In_391);
nor U738 (N_738,In_734,In_59);
nand U739 (N_739,In_344,In_46);
and U740 (N_740,In_321,In_359);
or U741 (N_741,In_635,In_280);
and U742 (N_742,In_677,In_666);
nor U743 (N_743,In_10,In_141);
nand U744 (N_744,In_306,In_491);
nor U745 (N_745,In_60,In_304);
or U746 (N_746,In_273,In_548);
and U747 (N_747,In_138,In_520);
nor U748 (N_748,In_551,In_689);
nor U749 (N_749,In_517,In_391);
nand U750 (N_750,In_345,In_670);
and U751 (N_751,In_382,In_373);
nor U752 (N_752,In_68,In_532);
nor U753 (N_753,In_431,In_484);
or U754 (N_754,In_298,In_444);
and U755 (N_755,In_189,In_402);
and U756 (N_756,In_286,In_184);
and U757 (N_757,In_53,In_35);
nand U758 (N_758,In_218,In_8);
nand U759 (N_759,In_257,In_594);
and U760 (N_760,In_291,In_524);
nor U761 (N_761,In_370,In_602);
and U762 (N_762,In_601,In_217);
and U763 (N_763,In_585,In_735);
nand U764 (N_764,In_136,In_37);
or U765 (N_765,In_307,In_96);
or U766 (N_766,In_314,In_233);
nand U767 (N_767,In_224,In_564);
nand U768 (N_768,In_727,In_259);
nor U769 (N_769,In_478,In_639);
and U770 (N_770,In_510,In_726);
nor U771 (N_771,In_327,In_126);
nand U772 (N_772,In_651,In_370);
nor U773 (N_773,In_362,In_251);
and U774 (N_774,In_137,In_443);
or U775 (N_775,In_61,In_409);
and U776 (N_776,In_396,In_452);
or U777 (N_777,In_60,In_453);
or U778 (N_778,In_631,In_488);
or U779 (N_779,In_120,In_401);
and U780 (N_780,In_27,In_274);
and U781 (N_781,In_589,In_358);
nor U782 (N_782,In_466,In_23);
nor U783 (N_783,In_315,In_744);
and U784 (N_784,In_510,In_225);
nand U785 (N_785,In_526,In_1);
and U786 (N_786,In_654,In_561);
nor U787 (N_787,In_74,In_636);
and U788 (N_788,In_708,In_526);
or U789 (N_789,In_715,In_530);
nand U790 (N_790,In_449,In_225);
nor U791 (N_791,In_224,In_607);
nand U792 (N_792,In_278,In_564);
nor U793 (N_793,In_549,In_562);
nor U794 (N_794,In_259,In_682);
and U795 (N_795,In_550,In_321);
and U796 (N_796,In_72,In_571);
nor U797 (N_797,In_437,In_252);
nor U798 (N_798,In_76,In_503);
nand U799 (N_799,In_668,In_540);
or U800 (N_800,In_140,In_225);
nand U801 (N_801,In_88,In_283);
or U802 (N_802,In_242,In_361);
or U803 (N_803,In_87,In_636);
nand U804 (N_804,In_145,In_373);
and U805 (N_805,In_411,In_303);
nor U806 (N_806,In_562,In_598);
nand U807 (N_807,In_602,In_189);
nor U808 (N_808,In_375,In_492);
nor U809 (N_809,In_661,In_393);
or U810 (N_810,In_632,In_424);
nor U811 (N_811,In_206,In_239);
xnor U812 (N_812,In_500,In_575);
and U813 (N_813,In_31,In_104);
nor U814 (N_814,In_673,In_223);
nor U815 (N_815,In_511,In_725);
and U816 (N_816,In_684,In_687);
nand U817 (N_817,In_731,In_407);
or U818 (N_818,In_505,In_119);
nand U819 (N_819,In_695,In_702);
or U820 (N_820,In_534,In_307);
and U821 (N_821,In_91,In_285);
nand U822 (N_822,In_189,In_94);
and U823 (N_823,In_275,In_408);
or U824 (N_824,In_444,In_154);
and U825 (N_825,In_380,In_111);
and U826 (N_826,In_585,In_88);
and U827 (N_827,In_312,In_519);
nor U828 (N_828,In_105,In_295);
nor U829 (N_829,In_216,In_671);
nand U830 (N_830,In_222,In_691);
nor U831 (N_831,In_326,In_217);
or U832 (N_832,In_175,In_350);
and U833 (N_833,In_569,In_685);
and U834 (N_834,In_414,In_470);
and U835 (N_835,In_164,In_231);
nor U836 (N_836,In_375,In_629);
or U837 (N_837,In_520,In_301);
nand U838 (N_838,In_208,In_293);
and U839 (N_839,In_656,In_554);
nand U840 (N_840,In_366,In_538);
xnor U841 (N_841,In_236,In_340);
nand U842 (N_842,In_434,In_725);
nand U843 (N_843,In_499,In_377);
and U844 (N_844,In_504,In_150);
or U845 (N_845,In_656,In_183);
and U846 (N_846,In_629,In_194);
nand U847 (N_847,In_219,In_360);
or U848 (N_848,In_569,In_672);
nor U849 (N_849,In_101,In_467);
nand U850 (N_850,In_336,In_201);
and U851 (N_851,In_283,In_158);
nor U852 (N_852,In_671,In_10);
nand U853 (N_853,In_183,In_737);
and U854 (N_854,In_227,In_684);
nor U855 (N_855,In_137,In_460);
nand U856 (N_856,In_226,In_182);
nand U857 (N_857,In_298,In_644);
nand U858 (N_858,In_707,In_339);
nor U859 (N_859,In_553,In_93);
nand U860 (N_860,In_41,In_711);
nand U861 (N_861,In_258,In_262);
nor U862 (N_862,In_208,In_183);
or U863 (N_863,In_635,In_674);
nand U864 (N_864,In_124,In_511);
and U865 (N_865,In_389,In_177);
or U866 (N_866,In_323,In_369);
or U867 (N_867,In_439,In_54);
nand U868 (N_868,In_69,In_253);
and U869 (N_869,In_175,In_204);
and U870 (N_870,In_524,In_492);
and U871 (N_871,In_607,In_622);
nand U872 (N_872,In_153,In_347);
nor U873 (N_873,In_584,In_555);
and U874 (N_874,In_485,In_338);
nor U875 (N_875,In_350,In_212);
or U876 (N_876,In_251,In_238);
and U877 (N_877,In_337,In_428);
and U878 (N_878,In_658,In_441);
nand U879 (N_879,In_123,In_221);
nand U880 (N_880,In_218,In_157);
and U881 (N_881,In_622,In_720);
and U882 (N_882,In_566,In_50);
or U883 (N_883,In_331,In_571);
or U884 (N_884,In_727,In_629);
or U885 (N_885,In_564,In_357);
and U886 (N_886,In_436,In_413);
or U887 (N_887,In_440,In_553);
nand U888 (N_888,In_492,In_119);
nor U889 (N_889,In_476,In_230);
nor U890 (N_890,In_582,In_154);
nor U891 (N_891,In_250,In_156);
nand U892 (N_892,In_184,In_226);
nand U893 (N_893,In_719,In_332);
and U894 (N_894,In_7,In_132);
or U895 (N_895,In_339,In_713);
or U896 (N_896,In_61,In_415);
nand U897 (N_897,In_710,In_228);
nand U898 (N_898,In_478,In_58);
nor U899 (N_899,In_238,In_62);
or U900 (N_900,In_628,In_264);
nor U901 (N_901,In_639,In_600);
nand U902 (N_902,In_280,In_649);
nand U903 (N_903,In_274,In_596);
nor U904 (N_904,In_215,In_651);
and U905 (N_905,In_557,In_361);
and U906 (N_906,In_351,In_232);
or U907 (N_907,In_488,In_246);
or U908 (N_908,In_588,In_673);
and U909 (N_909,In_352,In_147);
nand U910 (N_910,In_116,In_263);
xor U911 (N_911,In_454,In_550);
or U912 (N_912,In_205,In_333);
nor U913 (N_913,In_302,In_524);
nor U914 (N_914,In_372,In_352);
nor U915 (N_915,In_535,In_484);
and U916 (N_916,In_153,In_134);
nor U917 (N_917,In_104,In_723);
nand U918 (N_918,In_682,In_128);
and U919 (N_919,In_641,In_298);
nand U920 (N_920,In_167,In_494);
and U921 (N_921,In_489,In_409);
and U922 (N_922,In_55,In_697);
nand U923 (N_923,In_100,In_374);
nor U924 (N_924,In_359,In_592);
or U925 (N_925,In_179,In_302);
nand U926 (N_926,In_186,In_360);
nand U927 (N_927,In_509,In_732);
and U928 (N_928,In_219,In_727);
nand U929 (N_929,In_558,In_516);
or U930 (N_930,In_678,In_545);
nor U931 (N_931,In_406,In_13);
and U932 (N_932,In_153,In_696);
and U933 (N_933,In_166,In_17);
nand U934 (N_934,In_0,In_699);
or U935 (N_935,In_717,In_539);
or U936 (N_936,In_368,In_486);
nor U937 (N_937,In_198,In_540);
and U938 (N_938,In_602,In_16);
nand U939 (N_939,In_354,In_491);
nor U940 (N_940,In_602,In_303);
or U941 (N_941,In_321,In_646);
nor U942 (N_942,In_160,In_386);
nor U943 (N_943,In_425,In_248);
or U944 (N_944,In_366,In_387);
and U945 (N_945,In_443,In_703);
nor U946 (N_946,In_511,In_82);
nor U947 (N_947,In_659,In_571);
nor U948 (N_948,In_659,In_153);
or U949 (N_949,In_496,In_633);
nor U950 (N_950,In_303,In_589);
or U951 (N_951,In_210,In_622);
or U952 (N_952,In_184,In_616);
nor U953 (N_953,In_330,In_621);
nand U954 (N_954,In_173,In_657);
or U955 (N_955,In_256,In_730);
nor U956 (N_956,In_483,In_662);
nor U957 (N_957,In_549,In_680);
nor U958 (N_958,In_722,In_378);
and U959 (N_959,In_238,In_455);
and U960 (N_960,In_306,In_10);
nor U961 (N_961,In_146,In_119);
or U962 (N_962,In_315,In_19);
nor U963 (N_963,In_430,In_212);
or U964 (N_964,In_702,In_735);
or U965 (N_965,In_652,In_78);
nor U966 (N_966,In_626,In_640);
or U967 (N_967,In_320,In_395);
or U968 (N_968,In_623,In_743);
nand U969 (N_969,In_303,In_643);
or U970 (N_970,In_28,In_727);
nand U971 (N_971,In_657,In_440);
or U972 (N_972,In_206,In_168);
and U973 (N_973,In_279,In_531);
and U974 (N_974,In_571,In_700);
and U975 (N_975,In_256,In_403);
nand U976 (N_976,In_166,In_431);
nor U977 (N_977,In_208,In_51);
nor U978 (N_978,In_304,In_674);
or U979 (N_979,In_426,In_676);
nand U980 (N_980,In_55,In_164);
xnor U981 (N_981,In_675,In_739);
or U982 (N_982,In_449,In_689);
and U983 (N_983,In_283,In_742);
nand U984 (N_984,In_165,In_178);
or U985 (N_985,In_556,In_164);
nand U986 (N_986,In_539,In_523);
or U987 (N_987,In_432,In_338);
or U988 (N_988,In_737,In_273);
and U989 (N_989,In_480,In_629);
and U990 (N_990,In_193,In_249);
and U991 (N_991,In_655,In_422);
and U992 (N_992,In_261,In_450);
and U993 (N_993,In_492,In_505);
nand U994 (N_994,In_616,In_737);
or U995 (N_995,In_368,In_421);
and U996 (N_996,In_597,In_537);
and U997 (N_997,In_509,In_95);
nor U998 (N_998,In_337,In_675);
and U999 (N_999,In_212,In_647);
or U1000 (N_1000,In_228,In_300);
nand U1001 (N_1001,In_120,In_362);
nand U1002 (N_1002,In_568,In_340);
and U1003 (N_1003,In_599,In_589);
or U1004 (N_1004,In_248,In_260);
nand U1005 (N_1005,In_555,In_108);
and U1006 (N_1006,In_42,In_129);
or U1007 (N_1007,In_269,In_738);
and U1008 (N_1008,In_742,In_661);
nand U1009 (N_1009,In_264,In_576);
nand U1010 (N_1010,In_22,In_402);
nand U1011 (N_1011,In_290,In_155);
or U1012 (N_1012,In_492,In_620);
nor U1013 (N_1013,In_539,In_465);
nor U1014 (N_1014,In_212,In_476);
and U1015 (N_1015,In_490,In_322);
nand U1016 (N_1016,In_542,In_99);
and U1017 (N_1017,In_128,In_158);
nand U1018 (N_1018,In_173,In_606);
nand U1019 (N_1019,In_411,In_105);
or U1020 (N_1020,In_720,In_717);
or U1021 (N_1021,In_624,In_257);
nor U1022 (N_1022,In_536,In_555);
and U1023 (N_1023,In_591,In_632);
or U1024 (N_1024,In_645,In_286);
nor U1025 (N_1025,In_68,In_432);
or U1026 (N_1026,In_409,In_448);
or U1027 (N_1027,In_450,In_216);
nor U1028 (N_1028,In_481,In_44);
or U1029 (N_1029,In_551,In_32);
and U1030 (N_1030,In_393,In_213);
nor U1031 (N_1031,In_628,In_77);
and U1032 (N_1032,In_513,In_640);
or U1033 (N_1033,In_450,In_556);
nor U1034 (N_1034,In_622,In_110);
nand U1035 (N_1035,In_496,In_171);
or U1036 (N_1036,In_122,In_395);
or U1037 (N_1037,In_386,In_727);
nor U1038 (N_1038,In_454,In_674);
nor U1039 (N_1039,In_372,In_626);
nand U1040 (N_1040,In_248,In_120);
and U1041 (N_1041,In_96,In_385);
or U1042 (N_1042,In_50,In_231);
and U1043 (N_1043,In_193,In_671);
and U1044 (N_1044,In_419,In_249);
or U1045 (N_1045,In_322,In_381);
or U1046 (N_1046,In_489,In_25);
nand U1047 (N_1047,In_42,In_28);
or U1048 (N_1048,In_74,In_544);
nand U1049 (N_1049,In_477,In_523);
or U1050 (N_1050,In_705,In_487);
and U1051 (N_1051,In_321,In_502);
or U1052 (N_1052,In_444,In_357);
or U1053 (N_1053,In_232,In_35);
nand U1054 (N_1054,In_151,In_28);
and U1055 (N_1055,In_557,In_535);
nand U1056 (N_1056,In_94,In_267);
nor U1057 (N_1057,In_13,In_568);
or U1058 (N_1058,In_551,In_484);
and U1059 (N_1059,In_684,In_397);
nand U1060 (N_1060,In_135,In_263);
or U1061 (N_1061,In_247,In_28);
nand U1062 (N_1062,In_123,In_405);
and U1063 (N_1063,In_157,In_728);
or U1064 (N_1064,In_319,In_342);
or U1065 (N_1065,In_156,In_710);
or U1066 (N_1066,In_576,In_516);
nor U1067 (N_1067,In_2,In_749);
nand U1068 (N_1068,In_76,In_417);
nor U1069 (N_1069,In_201,In_288);
nor U1070 (N_1070,In_629,In_378);
nand U1071 (N_1071,In_213,In_419);
nand U1072 (N_1072,In_522,In_21);
or U1073 (N_1073,In_394,In_694);
nor U1074 (N_1074,In_731,In_412);
and U1075 (N_1075,In_256,In_142);
nor U1076 (N_1076,In_460,In_382);
nor U1077 (N_1077,In_152,In_347);
or U1078 (N_1078,In_64,In_246);
xor U1079 (N_1079,In_578,In_291);
nand U1080 (N_1080,In_519,In_58);
nor U1081 (N_1081,In_264,In_309);
nor U1082 (N_1082,In_610,In_559);
nand U1083 (N_1083,In_255,In_179);
nor U1084 (N_1084,In_57,In_489);
nand U1085 (N_1085,In_192,In_177);
or U1086 (N_1086,In_167,In_446);
nand U1087 (N_1087,In_537,In_602);
and U1088 (N_1088,In_187,In_148);
and U1089 (N_1089,In_202,In_599);
or U1090 (N_1090,In_146,In_725);
nor U1091 (N_1091,In_83,In_511);
and U1092 (N_1092,In_79,In_375);
or U1093 (N_1093,In_129,In_36);
and U1094 (N_1094,In_737,In_418);
and U1095 (N_1095,In_283,In_243);
nor U1096 (N_1096,In_596,In_114);
nor U1097 (N_1097,In_643,In_115);
nand U1098 (N_1098,In_143,In_295);
nor U1099 (N_1099,In_573,In_739);
and U1100 (N_1100,In_503,In_554);
nor U1101 (N_1101,In_337,In_435);
nor U1102 (N_1102,In_698,In_670);
nand U1103 (N_1103,In_356,In_455);
nor U1104 (N_1104,In_32,In_345);
nor U1105 (N_1105,In_426,In_183);
nand U1106 (N_1106,In_697,In_232);
nor U1107 (N_1107,In_296,In_293);
and U1108 (N_1108,In_492,In_208);
and U1109 (N_1109,In_652,In_336);
and U1110 (N_1110,In_342,In_504);
nand U1111 (N_1111,In_245,In_548);
nor U1112 (N_1112,In_596,In_599);
nor U1113 (N_1113,In_93,In_272);
nor U1114 (N_1114,In_55,In_181);
nor U1115 (N_1115,In_84,In_372);
and U1116 (N_1116,In_261,In_415);
nor U1117 (N_1117,In_507,In_651);
or U1118 (N_1118,In_469,In_414);
nand U1119 (N_1119,In_399,In_629);
nand U1120 (N_1120,In_385,In_600);
nor U1121 (N_1121,In_740,In_20);
and U1122 (N_1122,In_476,In_195);
nand U1123 (N_1123,In_456,In_184);
or U1124 (N_1124,In_477,In_355);
nor U1125 (N_1125,In_533,In_645);
nor U1126 (N_1126,In_227,In_164);
xor U1127 (N_1127,In_397,In_464);
and U1128 (N_1128,In_395,In_399);
and U1129 (N_1129,In_71,In_35);
and U1130 (N_1130,In_37,In_177);
nand U1131 (N_1131,In_315,In_510);
nand U1132 (N_1132,In_1,In_320);
nor U1133 (N_1133,In_205,In_224);
nand U1134 (N_1134,In_334,In_651);
nand U1135 (N_1135,In_265,In_229);
nor U1136 (N_1136,In_42,In_200);
or U1137 (N_1137,In_469,In_304);
and U1138 (N_1138,In_629,In_743);
nor U1139 (N_1139,In_494,In_631);
or U1140 (N_1140,In_211,In_177);
nor U1141 (N_1141,In_538,In_460);
nand U1142 (N_1142,In_273,In_106);
or U1143 (N_1143,In_317,In_341);
or U1144 (N_1144,In_310,In_467);
or U1145 (N_1145,In_265,In_613);
and U1146 (N_1146,In_226,In_514);
or U1147 (N_1147,In_623,In_679);
nand U1148 (N_1148,In_259,In_694);
and U1149 (N_1149,In_48,In_634);
and U1150 (N_1150,In_508,In_332);
nor U1151 (N_1151,In_310,In_687);
nand U1152 (N_1152,In_301,In_354);
nand U1153 (N_1153,In_123,In_368);
nand U1154 (N_1154,In_598,In_317);
nor U1155 (N_1155,In_420,In_626);
or U1156 (N_1156,In_608,In_159);
xor U1157 (N_1157,In_467,In_30);
or U1158 (N_1158,In_530,In_348);
nor U1159 (N_1159,In_429,In_72);
nand U1160 (N_1160,In_75,In_351);
and U1161 (N_1161,In_590,In_477);
or U1162 (N_1162,In_356,In_476);
nand U1163 (N_1163,In_545,In_558);
or U1164 (N_1164,In_665,In_79);
nor U1165 (N_1165,In_103,In_534);
and U1166 (N_1166,In_43,In_622);
or U1167 (N_1167,In_450,In_383);
nand U1168 (N_1168,In_696,In_189);
nand U1169 (N_1169,In_537,In_443);
nand U1170 (N_1170,In_194,In_68);
nor U1171 (N_1171,In_354,In_163);
or U1172 (N_1172,In_364,In_543);
and U1173 (N_1173,In_520,In_563);
nor U1174 (N_1174,In_89,In_388);
and U1175 (N_1175,In_539,In_373);
nand U1176 (N_1176,In_13,In_203);
and U1177 (N_1177,In_278,In_591);
nand U1178 (N_1178,In_667,In_24);
or U1179 (N_1179,In_522,In_426);
nand U1180 (N_1180,In_601,In_1);
nor U1181 (N_1181,In_404,In_176);
nor U1182 (N_1182,In_342,In_464);
nor U1183 (N_1183,In_664,In_179);
nor U1184 (N_1184,In_224,In_155);
nand U1185 (N_1185,In_495,In_216);
or U1186 (N_1186,In_238,In_74);
or U1187 (N_1187,In_262,In_57);
nor U1188 (N_1188,In_172,In_399);
and U1189 (N_1189,In_588,In_106);
and U1190 (N_1190,In_699,In_193);
and U1191 (N_1191,In_452,In_549);
nor U1192 (N_1192,In_93,In_497);
nand U1193 (N_1193,In_337,In_90);
nand U1194 (N_1194,In_74,In_623);
or U1195 (N_1195,In_264,In_616);
and U1196 (N_1196,In_525,In_473);
and U1197 (N_1197,In_586,In_181);
nor U1198 (N_1198,In_552,In_359);
nand U1199 (N_1199,In_290,In_309);
nand U1200 (N_1200,In_162,In_264);
nor U1201 (N_1201,In_10,In_385);
and U1202 (N_1202,In_380,In_142);
nor U1203 (N_1203,In_202,In_738);
or U1204 (N_1204,In_399,In_358);
and U1205 (N_1205,In_403,In_392);
or U1206 (N_1206,In_520,In_719);
or U1207 (N_1207,In_683,In_308);
and U1208 (N_1208,In_657,In_293);
nor U1209 (N_1209,In_662,In_537);
nor U1210 (N_1210,In_350,In_515);
nor U1211 (N_1211,In_701,In_273);
and U1212 (N_1212,In_414,In_748);
nor U1213 (N_1213,In_656,In_106);
nand U1214 (N_1214,In_666,In_146);
nand U1215 (N_1215,In_361,In_339);
nor U1216 (N_1216,In_6,In_420);
nor U1217 (N_1217,In_185,In_747);
nor U1218 (N_1218,In_554,In_140);
nand U1219 (N_1219,In_109,In_582);
nand U1220 (N_1220,In_45,In_280);
and U1221 (N_1221,In_145,In_586);
nor U1222 (N_1222,In_453,In_317);
and U1223 (N_1223,In_605,In_542);
nand U1224 (N_1224,In_110,In_523);
or U1225 (N_1225,In_90,In_584);
or U1226 (N_1226,In_280,In_618);
and U1227 (N_1227,In_473,In_160);
and U1228 (N_1228,In_720,In_715);
nand U1229 (N_1229,In_377,In_342);
or U1230 (N_1230,In_433,In_698);
nor U1231 (N_1231,In_629,In_426);
or U1232 (N_1232,In_292,In_108);
or U1233 (N_1233,In_416,In_340);
or U1234 (N_1234,In_235,In_206);
nor U1235 (N_1235,In_382,In_464);
and U1236 (N_1236,In_143,In_505);
and U1237 (N_1237,In_354,In_4);
nor U1238 (N_1238,In_313,In_249);
and U1239 (N_1239,In_652,In_285);
and U1240 (N_1240,In_460,In_285);
nor U1241 (N_1241,In_112,In_71);
nor U1242 (N_1242,In_575,In_196);
and U1243 (N_1243,In_436,In_740);
nor U1244 (N_1244,In_717,In_133);
and U1245 (N_1245,In_147,In_691);
or U1246 (N_1246,In_535,In_552);
nand U1247 (N_1247,In_536,In_605);
and U1248 (N_1248,In_481,In_389);
nor U1249 (N_1249,In_398,In_406);
nand U1250 (N_1250,In_226,In_382);
nor U1251 (N_1251,In_290,In_419);
and U1252 (N_1252,In_49,In_230);
nor U1253 (N_1253,In_208,In_748);
and U1254 (N_1254,In_127,In_72);
nand U1255 (N_1255,In_570,In_154);
and U1256 (N_1256,In_576,In_66);
nor U1257 (N_1257,In_326,In_680);
or U1258 (N_1258,In_378,In_55);
or U1259 (N_1259,In_319,In_660);
nor U1260 (N_1260,In_649,In_565);
or U1261 (N_1261,In_236,In_589);
and U1262 (N_1262,In_327,In_54);
and U1263 (N_1263,In_94,In_574);
nor U1264 (N_1264,In_364,In_532);
and U1265 (N_1265,In_257,In_11);
and U1266 (N_1266,In_709,In_112);
or U1267 (N_1267,In_255,In_143);
or U1268 (N_1268,In_180,In_684);
and U1269 (N_1269,In_728,In_444);
nor U1270 (N_1270,In_557,In_439);
nand U1271 (N_1271,In_581,In_689);
or U1272 (N_1272,In_458,In_303);
or U1273 (N_1273,In_245,In_373);
nand U1274 (N_1274,In_633,In_725);
nor U1275 (N_1275,In_129,In_199);
nor U1276 (N_1276,In_195,In_705);
and U1277 (N_1277,In_288,In_300);
or U1278 (N_1278,In_323,In_298);
and U1279 (N_1279,In_192,In_89);
or U1280 (N_1280,In_506,In_179);
nor U1281 (N_1281,In_92,In_724);
nor U1282 (N_1282,In_575,In_416);
or U1283 (N_1283,In_394,In_75);
or U1284 (N_1284,In_613,In_98);
nor U1285 (N_1285,In_721,In_149);
nand U1286 (N_1286,In_66,In_557);
nand U1287 (N_1287,In_507,In_190);
or U1288 (N_1288,In_182,In_313);
nor U1289 (N_1289,In_618,In_682);
nor U1290 (N_1290,In_560,In_332);
nand U1291 (N_1291,In_471,In_740);
nand U1292 (N_1292,In_429,In_5);
and U1293 (N_1293,In_29,In_229);
or U1294 (N_1294,In_91,In_597);
and U1295 (N_1295,In_549,In_133);
and U1296 (N_1296,In_181,In_15);
nor U1297 (N_1297,In_373,In_666);
nand U1298 (N_1298,In_719,In_615);
and U1299 (N_1299,In_291,In_163);
nand U1300 (N_1300,In_211,In_688);
and U1301 (N_1301,In_252,In_492);
nand U1302 (N_1302,In_726,In_383);
nor U1303 (N_1303,In_94,In_176);
nor U1304 (N_1304,In_330,In_92);
or U1305 (N_1305,In_173,In_179);
and U1306 (N_1306,In_119,In_124);
nand U1307 (N_1307,In_191,In_479);
and U1308 (N_1308,In_555,In_654);
and U1309 (N_1309,In_584,In_382);
nor U1310 (N_1310,In_562,In_332);
nand U1311 (N_1311,In_158,In_638);
nand U1312 (N_1312,In_87,In_204);
or U1313 (N_1313,In_619,In_601);
nor U1314 (N_1314,In_329,In_435);
nand U1315 (N_1315,In_522,In_137);
or U1316 (N_1316,In_695,In_230);
or U1317 (N_1317,In_50,In_555);
nand U1318 (N_1318,In_530,In_742);
nand U1319 (N_1319,In_291,In_48);
nand U1320 (N_1320,In_377,In_646);
and U1321 (N_1321,In_388,In_531);
and U1322 (N_1322,In_124,In_713);
nor U1323 (N_1323,In_170,In_523);
nand U1324 (N_1324,In_467,In_32);
nand U1325 (N_1325,In_59,In_5);
nand U1326 (N_1326,In_116,In_108);
nor U1327 (N_1327,In_179,In_203);
nand U1328 (N_1328,In_428,In_313);
nand U1329 (N_1329,In_184,In_620);
nand U1330 (N_1330,In_116,In_685);
nor U1331 (N_1331,In_481,In_361);
or U1332 (N_1332,In_176,In_4);
nor U1333 (N_1333,In_592,In_482);
and U1334 (N_1334,In_63,In_630);
nor U1335 (N_1335,In_378,In_149);
nand U1336 (N_1336,In_266,In_0);
xnor U1337 (N_1337,In_497,In_581);
nand U1338 (N_1338,In_674,In_157);
xor U1339 (N_1339,In_674,In_553);
or U1340 (N_1340,In_21,In_619);
and U1341 (N_1341,In_264,In_672);
or U1342 (N_1342,In_531,In_257);
or U1343 (N_1343,In_295,In_697);
nor U1344 (N_1344,In_360,In_454);
nand U1345 (N_1345,In_464,In_254);
nor U1346 (N_1346,In_24,In_680);
nor U1347 (N_1347,In_426,In_481);
and U1348 (N_1348,In_614,In_664);
nand U1349 (N_1349,In_541,In_672);
and U1350 (N_1350,In_719,In_472);
nor U1351 (N_1351,In_665,In_652);
or U1352 (N_1352,In_720,In_31);
or U1353 (N_1353,In_475,In_698);
nand U1354 (N_1354,In_85,In_329);
nand U1355 (N_1355,In_235,In_308);
nor U1356 (N_1356,In_659,In_713);
nor U1357 (N_1357,In_732,In_203);
nor U1358 (N_1358,In_611,In_408);
and U1359 (N_1359,In_727,In_630);
or U1360 (N_1360,In_626,In_308);
nand U1361 (N_1361,In_156,In_342);
and U1362 (N_1362,In_52,In_237);
nor U1363 (N_1363,In_67,In_735);
or U1364 (N_1364,In_581,In_257);
nand U1365 (N_1365,In_171,In_281);
nor U1366 (N_1366,In_39,In_391);
nand U1367 (N_1367,In_361,In_369);
nor U1368 (N_1368,In_44,In_24);
and U1369 (N_1369,In_392,In_361);
nor U1370 (N_1370,In_10,In_515);
nor U1371 (N_1371,In_456,In_167);
nor U1372 (N_1372,In_399,In_713);
and U1373 (N_1373,In_211,In_152);
or U1374 (N_1374,In_611,In_332);
or U1375 (N_1375,In_305,In_500);
nor U1376 (N_1376,In_505,In_583);
nor U1377 (N_1377,In_703,In_91);
nand U1378 (N_1378,In_436,In_134);
nand U1379 (N_1379,In_734,In_683);
nor U1380 (N_1380,In_153,In_619);
nor U1381 (N_1381,In_498,In_511);
nand U1382 (N_1382,In_392,In_587);
nor U1383 (N_1383,In_387,In_364);
and U1384 (N_1384,In_181,In_297);
nand U1385 (N_1385,In_474,In_508);
and U1386 (N_1386,In_535,In_273);
or U1387 (N_1387,In_588,In_88);
or U1388 (N_1388,In_488,In_685);
and U1389 (N_1389,In_670,In_465);
nand U1390 (N_1390,In_458,In_606);
or U1391 (N_1391,In_258,In_274);
nor U1392 (N_1392,In_198,In_271);
nor U1393 (N_1393,In_570,In_507);
nand U1394 (N_1394,In_538,In_674);
and U1395 (N_1395,In_614,In_197);
nor U1396 (N_1396,In_651,In_198);
and U1397 (N_1397,In_155,In_664);
and U1398 (N_1398,In_458,In_523);
xor U1399 (N_1399,In_736,In_647);
or U1400 (N_1400,In_386,In_587);
and U1401 (N_1401,In_647,In_531);
xor U1402 (N_1402,In_495,In_176);
nor U1403 (N_1403,In_87,In_48);
nand U1404 (N_1404,In_600,In_387);
nand U1405 (N_1405,In_499,In_697);
and U1406 (N_1406,In_569,In_257);
or U1407 (N_1407,In_110,In_658);
and U1408 (N_1408,In_675,In_308);
or U1409 (N_1409,In_230,In_91);
or U1410 (N_1410,In_249,In_588);
nor U1411 (N_1411,In_684,In_241);
or U1412 (N_1412,In_444,In_553);
nor U1413 (N_1413,In_154,In_652);
or U1414 (N_1414,In_435,In_338);
or U1415 (N_1415,In_544,In_597);
nor U1416 (N_1416,In_416,In_315);
and U1417 (N_1417,In_199,In_559);
nand U1418 (N_1418,In_744,In_134);
nand U1419 (N_1419,In_680,In_628);
xnor U1420 (N_1420,In_89,In_550);
nand U1421 (N_1421,In_11,In_328);
nor U1422 (N_1422,In_355,In_714);
nor U1423 (N_1423,In_256,In_164);
or U1424 (N_1424,In_199,In_331);
or U1425 (N_1425,In_73,In_229);
nand U1426 (N_1426,In_329,In_500);
or U1427 (N_1427,In_199,In_102);
or U1428 (N_1428,In_664,In_403);
nor U1429 (N_1429,In_572,In_341);
or U1430 (N_1430,In_569,In_510);
and U1431 (N_1431,In_497,In_29);
and U1432 (N_1432,In_443,In_86);
or U1433 (N_1433,In_109,In_111);
nor U1434 (N_1434,In_596,In_230);
nor U1435 (N_1435,In_400,In_583);
or U1436 (N_1436,In_54,In_83);
nor U1437 (N_1437,In_422,In_445);
nand U1438 (N_1438,In_498,In_692);
nand U1439 (N_1439,In_586,In_130);
and U1440 (N_1440,In_167,In_144);
or U1441 (N_1441,In_174,In_577);
nand U1442 (N_1442,In_676,In_439);
or U1443 (N_1443,In_611,In_409);
or U1444 (N_1444,In_629,In_442);
or U1445 (N_1445,In_450,In_262);
and U1446 (N_1446,In_677,In_300);
nor U1447 (N_1447,In_660,In_626);
and U1448 (N_1448,In_94,In_76);
and U1449 (N_1449,In_214,In_3);
nand U1450 (N_1450,In_563,In_62);
nand U1451 (N_1451,In_724,In_645);
or U1452 (N_1452,In_507,In_696);
nor U1453 (N_1453,In_92,In_118);
and U1454 (N_1454,In_385,In_352);
or U1455 (N_1455,In_383,In_655);
nor U1456 (N_1456,In_728,In_297);
nand U1457 (N_1457,In_287,In_377);
nand U1458 (N_1458,In_576,In_575);
nand U1459 (N_1459,In_669,In_301);
or U1460 (N_1460,In_610,In_603);
nand U1461 (N_1461,In_487,In_717);
and U1462 (N_1462,In_525,In_490);
nor U1463 (N_1463,In_667,In_97);
and U1464 (N_1464,In_199,In_608);
nand U1465 (N_1465,In_368,In_553);
nand U1466 (N_1466,In_584,In_43);
nand U1467 (N_1467,In_350,In_122);
or U1468 (N_1468,In_215,In_656);
and U1469 (N_1469,In_242,In_24);
or U1470 (N_1470,In_723,In_253);
nor U1471 (N_1471,In_249,In_621);
or U1472 (N_1472,In_393,In_68);
nand U1473 (N_1473,In_470,In_348);
nand U1474 (N_1474,In_253,In_614);
and U1475 (N_1475,In_212,In_363);
nor U1476 (N_1476,In_479,In_561);
nand U1477 (N_1477,In_483,In_719);
or U1478 (N_1478,In_363,In_731);
and U1479 (N_1479,In_405,In_574);
nor U1480 (N_1480,In_747,In_24);
nand U1481 (N_1481,In_89,In_598);
nand U1482 (N_1482,In_671,In_18);
or U1483 (N_1483,In_714,In_404);
and U1484 (N_1484,In_36,In_25);
nor U1485 (N_1485,In_590,In_450);
nor U1486 (N_1486,In_230,In_265);
or U1487 (N_1487,In_743,In_497);
nor U1488 (N_1488,In_637,In_654);
and U1489 (N_1489,In_174,In_253);
or U1490 (N_1490,In_441,In_286);
nor U1491 (N_1491,In_29,In_530);
and U1492 (N_1492,In_408,In_28);
nor U1493 (N_1493,In_199,In_639);
nand U1494 (N_1494,In_563,In_452);
and U1495 (N_1495,In_129,In_206);
and U1496 (N_1496,In_544,In_363);
nor U1497 (N_1497,In_594,In_343);
nor U1498 (N_1498,In_141,In_151);
nand U1499 (N_1499,In_602,In_111);
or U1500 (N_1500,In_381,In_134);
nor U1501 (N_1501,In_721,In_746);
or U1502 (N_1502,In_71,In_397);
nor U1503 (N_1503,In_101,In_165);
or U1504 (N_1504,In_727,In_551);
or U1505 (N_1505,In_345,In_504);
and U1506 (N_1506,In_169,In_591);
nand U1507 (N_1507,In_703,In_279);
or U1508 (N_1508,In_105,In_153);
or U1509 (N_1509,In_132,In_317);
nor U1510 (N_1510,In_447,In_351);
nor U1511 (N_1511,In_747,In_35);
and U1512 (N_1512,In_527,In_213);
nand U1513 (N_1513,In_332,In_13);
and U1514 (N_1514,In_729,In_488);
or U1515 (N_1515,In_234,In_722);
nand U1516 (N_1516,In_562,In_342);
nor U1517 (N_1517,In_122,In_525);
nand U1518 (N_1518,In_16,In_466);
and U1519 (N_1519,In_713,In_12);
nand U1520 (N_1520,In_85,In_486);
nand U1521 (N_1521,In_576,In_683);
or U1522 (N_1522,In_393,In_169);
xnor U1523 (N_1523,In_364,In_118);
nand U1524 (N_1524,In_218,In_111);
nand U1525 (N_1525,In_30,In_97);
nor U1526 (N_1526,In_582,In_128);
and U1527 (N_1527,In_497,In_528);
nand U1528 (N_1528,In_233,In_131);
and U1529 (N_1529,In_682,In_22);
or U1530 (N_1530,In_650,In_343);
nand U1531 (N_1531,In_42,In_622);
nand U1532 (N_1532,In_674,In_413);
nand U1533 (N_1533,In_609,In_603);
nor U1534 (N_1534,In_98,In_185);
xnor U1535 (N_1535,In_103,In_415);
nand U1536 (N_1536,In_48,In_284);
or U1537 (N_1537,In_458,In_175);
and U1538 (N_1538,In_718,In_723);
nor U1539 (N_1539,In_242,In_175);
and U1540 (N_1540,In_111,In_173);
or U1541 (N_1541,In_20,In_371);
nor U1542 (N_1542,In_660,In_318);
nand U1543 (N_1543,In_520,In_356);
nor U1544 (N_1544,In_705,In_652);
nand U1545 (N_1545,In_559,In_227);
or U1546 (N_1546,In_491,In_82);
and U1547 (N_1547,In_157,In_566);
and U1548 (N_1548,In_152,In_138);
or U1549 (N_1549,In_510,In_37);
or U1550 (N_1550,In_248,In_488);
nor U1551 (N_1551,In_380,In_33);
nor U1552 (N_1552,In_578,In_233);
or U1553 (N_1553,In_546,In_548);
nor U1554 (N_1554,In_677,In_628);
nor U1555 (N_1555,In_702,In_402);
and U1556 (N_1556,In_611,In_658);
or U1557 (N_1557,In_550,In_669);
and U1558 (N_1558,In_350,In_52);
nand U1559 (N_1559,In_76,In_267);
nand U1560 (N_1560,In_494,In_12);
or U1561 (N_1561,In_676,In_39);
nand U1562 (N_1562,In_678,In_105);
or U1563 (N_1563,In_306,In_556);
and U1564 (N_1564,In_407,In_718);
and U1565 (N_1565,In_187,In_573);
and U1566 (N_1566,In_23,In_282);
nor U1567 (N_1567,In_555,In_39);
nand U1568 (N_1568,In_686,In_566);
nor U1569 (N_1569,In_511,In_193);
and U1570 (N_1570,In_737,In_37);
or U1571 (N_1571,In_466,In_181);
and U1572 (N_1572,In_165,In_680);
nor U1573 (N_1573,In_374,In_339);
and U1574 (N_1574,In_713,In_382);
nor U1575 (N_1575,In_147,In_175);
or U1576 (N_1576,In_663,In_300);
and U1577 (N_1577,In_520,In_36);
or U1578 (N_1578,In_194,In_720);
or U1579 (N_1579,In_546,In_708);
nor U1580 (N_1580,In_12,In_734);
or U1581 (N_1581,In_688,In_461);
and U1582 (N_1582,In_686,In_203);
and U1583 (N_1583,In_242,In_111);
and U1584 (N_1584,In_573,In_13);
or U1585 (N_1585,In_359,In_9);
and U1586 (N_1586,In_234,In_561);
and U1587 (N_1587,In_159,In_173);
nand U1588 (N_1588,In_61,In_335);
nor U1589 (N_1589,In_302,In_636);
nand U1590 (N_1590,In_173,In_555);
nor U1591 (N_1591,In_199,In_206);
or U1592 (N_1592,In_217,In_714);
and U1593 (N_1593,In_157,In_362);
nor U1594 (N_1594,In_127,In_698);
nand U1595 (N_1595,In_203,In_233);
nand U1596 (N_1596,In_387,In_699);
xor U1597 (N_1597,In_45,In_302);
or U1598 (N_1598,In_406,In_655);
and U1599 (N_1599,In_483,In_228);
nor U1600 (N_1600,In_564,In_3);
and U1601 (N_1601,In_530,In_127);
nor U1602 (N_1602,In_293,In_446);
nand U1603 (N_1603,In_369,In_33);
nand U1604 (N_1604,In_247,In_742);
nand U1605 (N_1605,In_577,In_236);
or U1606 (N_1606,In_20,In_623);
nor U1607 (N_1607,In_408,In_229);
and U1608 (N_1608,In_597,In_327);
and U1609 (N_1609,In_576,In_585);
nand U1610 (N_1610,In_64,In_388);
and U1611 (N_1611,In_630,In_48);
nor U1612 (N_1612,In_119,In_713);
or U1613 (N_1613,In_599,In_236);
nand U1614 (N_1614,In_279,In_643);
nand U1615 (N_1615,In_397,In_637);
or U1616 (N_1616,In_719,In_26);
nor U1617 (N_1617,In_233,In_617);
nor U1618 (N_1618,In_381,In_97);
or U1619 (N_1619,In_359,In_616);
nor U1620 (N_1620,In_371,In_347);
nand U1621 (N_1621,In_550,In_150);
nor U1622 (N_1622,In_40,In_661);
or U1623 (N_1623,In_281,In_70);
or U1624 (N_1624,In_59,In_714);
nand U1625 (N_1625,In_148,In_628);
or U1626 (N_1626,In_256,In_360);
nor U1627 (N_1627,In_681,In_239);
nand U1628 (N_1628,In_408,In_431);
nand U1629 (N_1629,In_327,In_665);
nor U1630 (N_1630,In_155,In_462);
or U1631 (N_1631,In_120,In_561);
nand U1632 (N_1632,In_737,In_495);
and U1633 (N_1633,In_698,In_25);
nand U1634 (N_1634,In_245,In_579);
nand U1635 (N_1635,In_654,In_238);
or U1636 (N_1636,In_48,In_614);
nor U1637 (N_1637,In_714,In_358);
nor U1638 (N_1638,In_32,In_195);
nor U1639 (N_1639,In_580,In_117);
nand U1640 (N_1640,In_628,In_218);
nand U1641 (N_1641,In_96,In_526);
or U1642 (N_1642,In_174,In_586);
or U1643 (N_1643,In_386,In_255);
nor U1644 (N_1644,In_139,In_411);
nor U1645 (N_1645,In_376,In_663);
and U1646 (N_1646,In_207,In_53);
nand U1647 (N_1647,In_562,In_724);
or U1648 (N_1648,In_603,In_601);
nor U1649 (N_1649,In_107,In_667);
and U1650 (N_1650,In_490,In_133);
nor U1651 (N_1651,In_327,In_158);
or U1652 (N_1652,In_642,In_418);
nor U1653 (N_1653,In_505,In_411);
or U1654 (N_1654,In_306,In_661);
and U1655 (N_1655,In_110,In_612);
and U1656 (N_1656,In_76,In_591);
or U1657 (N_1657,In_532,In_721);
nand U1658 (N_1658,In_242,In_661);
nand U1659 (N_1659,In_76,In_587);
and U1660 (N_1660,In_222,In_19);
nor U1661 (N_1661,In_547,In_454);
nand U1662 (N_1662,In_440,In_642);
or U1663 (N_1663,In_619,In_678);
or U1664 (N_1664,In_653,In_652);
nor U1665 (N_1665,In_607,In_102);
nor U1666 (N_1666,In_237,In_207);
and U1667 (N_1667,In_283,In_209);
and U1668 (N_1668,In_210,In_428);
or U1669 (N_1669,In_387,In_620);
nor U1670 (N_1670,In_456,In_619);
nor U1671 (N_1671,In_154,In_327);
nand U1672 (N_1672,In_266,In_4);
nor U1673 (N_1673,In_13,In_110);
nor U1674 (N_1674,In_294,In_95);
or U1675 (N_1675,In_335,In_705);
and U1676 (N_1676,In_451,In_163);
nand U1677 (N_1677,In_123,In_245);
and U1678 (N_1678,In_284,In_297);
nor U1679 (N_1679,In_134,In_306);
and U1680 (N_1680,In_147,In_8);
and U1681 (N_1681,In_632,In_232);
nor U1682 (N_1682,In_606,In_451);
nor U1683 (N_1683,In_456,In_202);
and U1684 (N_1684,In_546,In_480);
nor U1685 (N_1685,In_543,In_156);
nand U1686 (N_1686,In_107,In_427);
and U1687 (N_1687,In_414,In_54);
nor U1688 (N_1688,In_592,In_391);
nand U1689 (N_1689,In_259,In_658);
and U1690 (N_1690,In_223,In_63);
nand U1691 (N_1691,In_629,In_61);
and U1692 (N_1692,In_434,In_311);
nor U1693 (N_1693,In_642,In_447);
nor U1694 (N_1694,In_190,In_211);
nand U1695 (N_1695,In_674,In_38);
nor U1696 (N_1696,In_271,In_173);
or U1697 (N_1697,In_124,In_189);
nor U1698 (N_1698,In_132,In_509);
or U1699 (N_1699,In_672,In_248);
nand U1700 (N_1700,In_494,In_279);
nand U1701 (N_1701,In_189,In_376);
or U1702 (N_1702,In_535,In_396);
and U1703 (N_1703,In_223,In_613);
nor U1704 (N_1704,In_611,In_568);
or U1705 (N_1705,In_377,In_483);
nand U1706 (N_1706,In_221,In_533);
nor U1707 (N_1707,In_696,In_540);
or U1708 (N_1708,In_19,In_273);
and U1709 (N_1709,In_660,In_410);
or U1710 (N_1710,In_746,In_72);
and U1711 (N_1711,In_197,In_173);
nand U1712 (N_1712,In_566,In_54);
nand U1713 (N_1713,In_455,In_129);
nand U1714 (N_1714,In_67,In_668);
nand U1715 (N_1715,In_137,In_538);
nor U1716 (N_1716,In_686,In_114);
and U1717 (N_1717,In_308,In_483);
or U1718 (N_1718,In_100,In_73);
and U1719 (N_1719,In_117,In_203);
or U1720 (N_1720,In_592,In_305);
and U1721 (N_1721,In_464,In_503);
nand U1722 (N_1722,In_396,In_362);
and U1723 (N_1723,In_169,In_128);
and U1724 (N_1724,In_101,In_479);
nand U1725 (N_1725,In_245,In_514);
or U1726 (N_1726,In_599,In_314);
and U1727 (N_1727,In_283,In_593);
nor U1728 (N_1728,In_632,In_128);
nor U1729 (N_1729,In_260,In_614);
or U1730 (N_1730,In_595,In_93);
or U1731 (N_1731,In_65,In_653);
and U1732 (N_1732,In_139,In_573);
or U1733 (N_1733,In_234,In_50);
and U1734 (N_1734,In_434,In_44);
nand U1735 (N_1735,In_520,In_371);
nand U1736 (N_1736,In_632,In_198);
and U1737 (N_1737,In_180,In_235);
nand U1738 (N_1738,In_207,In_62);
and U1739 (N_1739,In_347,In_645);
or U1740 (N_1740,In_258,In_537);
nor U1741 (N_1741,In_611,In_131);
nor U1742 (N_1742,In_574,In_90);
xnor U1743 (N_1743,In_432,In_236);
and U1744 (N_1744,In_166,In_328);
nor U1745 (N_1745,In_579,In_72);
xnor U1746 (N_1746,In_215,In_195);
and U1747 (N_1747,In_136,In_79);
nand U1748 (N_1748,In_477,In_392);
and U1749 (N_1749,In_650,In_434);
and U1750 (N_1750,In_607,In_10);
nand U1751 (N_1751,In_599,In_741);
nor U1752 (N_1752,In_709,In_692);
nand U1753 (N_1753,In_460,In_86);
nor U1754 (N_1754,In_543,In_299);
nor U1755 (N_1755,In_740,In_317);
and U1756 (N_1756,In_732,In_634);
nand U1757 (N_1757,In_375,In_543);
nor U1758 (N_1758,In_161,In_749);
and U1759 (N_1759,In_748,In_282);
or U1760 (N_1760,In_349,In_738);
or U1761 (N_1761,In_225,In_644);
and U1762 (N_1762,In_622,In_181);
nor U1763 (N_1763,In_394,In_66);
nor U1764 (N_1764,In_243,In_176);
nand U1765 (N_1765,In_238,In_647);
nor U1766 (N_1766,In_215,In_359);
nand U1767 (N_1767,In_630,In_715);
nor U1768 (N_1768,In_613,In_31);
nor U1769 (N_1769,In_374,In_45);
or U1770 (N_1770,In_711,In_402);
and U1771 (N_1771,In_697,In_238);
nand U1772 (N_1772,In_688,In_518);
or U1773 (N_1773,In_697,In_28);
xnor U1774 (N_1774,In_201,In_554);
or U1775 (N_1775,In_449,In_169);
nand U1776 (N_1776,In_177,In_487);
nor U1777 (N_1777,In_601,In_306);
nor U1778 (N_1778,In_141,In_105);
and U1779 (N_1779,In_22,In_457);
nand U1780 (N_1780,In_387,In_300);
nor U1781 (N_1781,In_543,In_537);
nand U1782 (N_1782,In_455,In_296);
or U1783 (N_1783,In_372,In_560);
and U1784 (N_1784,In_207,In_228);
nor U1785 (N_1785,In_22,In_60);
nor U1786 (N_1786,In_402,In_145);
nor U1787 (N_1787,In_306,In_466);
and U1788 (N_1788,In_116,In_598);
or U1789 (N_1789,In_20,In_723);
nand U1790 (N_1790,In_353,In_121);
nor U1791 (N_1791,In_139,In_249);
nor U1792 (N_1792,In_284,In_424);
or U1793 (N_1793,In_400,In_748);
or U1794 (N_1794,In_250,In_686);
nor U1795 (N_1795,In_529,In_452);
nand U1796 (N_1796,In_14,In_417);
and U1797 (N_1797,In_164,In_682);
and U1798 (N_1798,In_599,In_555);
nor U1799 (N_1799,In_142,In_622);
and U1800 (N_1800,In_152,In_431);
nand U1801 (N_1801,In_507,In_409);
nand U1802 (N_1802,In_137,In_231);
and U1803 (N_1803,In_26,In_342);
nor U1804 (N_1804,In_151,In_278);
xor U1805 (N_1805,In_627,In_660);
nor U1806 (N_1806,In_305,In_449);
and U1807 (N_1807,In_532,In_633);
nand U1808 (N_1808,In_0,In_107);
nor U1809 (N_1809,In_673,In_616);
nand U1810 (N_1810,In_721,In_139);
nand U1811 (N_1811,In_313,In_276);
nor U1812 (N_1812,In_349,In_546);
and U1813 (N_1813,In_220,In_415);
nand U1814 (N_1814,In_704,In_181);
xor U1815 (N_1815,In_99,In_487);
or U1816 (N_1816,In_517,In_705);
and U1817 (N_1817,In_7,In_425);
and U1818 (N_1818,In_85,In_643);
nor U1819 (N_1819,In_270,In_6);
nand U1820 (N_1820,In_378,In_301);
and U1821 (N_1821,In_90,In_159);
nor U1822 (N_1822,In_735,In_292);
xor U1823 (N_1823,In_88,In_687);
or U1824 (N_1824,In_188,In_607);
or U1825 (N_1825,In_51,In_416);
nor U1826 (N_1826,In_283,In_356);
and U1827 (N_1827,In_150,In_121);
or U1828 (N_1828,In_530,In_328);
or U1829 (N_1829,In_12,In_518);
nor U1830 (N_1830,In_652,In_628);
nor U1831 (N_1831,In_504,In_466);
nor U1832 (N_1832,In_127,In_446);
and U1833 (N_1833,In_404,In_472);
nor U1834 (N_1834,In_39,In_226);
or U1835 (N_1835,In_256,In_606);
or U1836 (N_1836,In_347,In_278);
nor U1837 (N_1837,In_164,In_652);
or U1838 (N_1838,In_565,In_306);
nand U1839 (N_1839,In_625,In_293);
nand U1840 (N_1840,In_243,In_724);
and U1841 (N_1841,In_369,In_379);
nand U1842 (N_1842,In_130,In_640);
nor U1843 (N_1843,In_518,In_354);
and U1844 (N_1844,In_145,In_175);
nand U1845 (N_1845,In_170,In_387);
nand U1846 (N_1846,In_134,In_206);
xor U1847 (N_1847,In_515,In_184);
nand U1848 (N_1848,In_381,In_38);
nor U1849 (N_1849,In_600,In_133);
nor U1850 (N_1850,In_639,In_156);
or U1851 (N_1851,In_652,In_158);
nor U1852 (N_1852,In_20,In_461);
or U1853 (N_1853,In_712,In_277);
or U1854 (N_1854,In_350,In_579);
nor U1855 (N_1855,In_477,In_678);
or U1856 (N_1856,In_245,In_293);
or U1857 (N_1857,In_341,In_49);
or U1858 (N_1858,In_278,In_269);
and U1859 (N_1859,In_445,In_86);
nand U1860 (N_1860,In_45,In_62);
nor U1861 (N_1861,In_646,In_526);
nand U1862 (N_1862,In_295,In_651);
nand U1863 (N_1863,In_36,In_15);
nand U1864 (N_1864,In_268,In_62);
nand U1865 (N_1865,In_427,In_244);
nand U1866 (N_1866,In_676,In_529);
nand U1867 (N_1867,In_45,In_75);
and U1868 (N_1868,In_519,In_713);
nand U1869 (N_1869,In_122,In_133);
or U1870 (N_1870,In_365,In_496);
nor U1871 (N_1871,In_193,In_330);
nand U1872 (N_1872,In_242,In_280);
nor U1873 (N_1873,In_283,In_23);
or U1874 (N_1874,In_24,In_480);
nor U1875 (N_1875,In_134,In_734);
nand U1876 (N_1876,In_45,In_404);
or U1877 (N_1877,In_394,In_97);
or U1878 (N_1878,In_64,In_532);
nand U1879 (N_1879,In_669,In_503);
and U1880 (N_1880,In_384,In_662);
or U1881 (N_1881,In_459,In_207);
or U1882 (N_1882,In_203,In_426);
or U1883 (N_1883,In_737,In_666);
and U1884 (N_1884,In_462,In_618);
and U1885 (N_1885,In_422,In_570);
nor U1886 (N_1886,In_503,In_117);
nor U1887 (N_1887,In_299,In_689);
nor U1888 (N_1888,In_715,In_508);
nand U1889 (N_1889,In_679,In_155);
nand U1890 (N_1890,In_344,In_456);
xnor U1891 (N_1891,In_537,In_730);
or U1892 (N_1892,In_705,In_379);
nor U1893 (N_1893,In_331,In_117);
nand U1894 (N_1894,In_672,In_582);
nand U1895 (N_1895,In_194,In_518);
nor U1896 (N_1896,In_676,In_183);
and U1897 (N_1897,In_459,In_293);
and U1898 (N_1898,In_216,In_355);
nand U1899 (N_1899,In_625,In_224);
and U1900 (N_1900,In_41,In_128);
and U1901 (N_1901,In_394,In_485);
and U1902 (N_1902,In_135,In_301);
nand U1903 (N_1903,In_217,In_541);
and U1904 (N_1904,In_388,In_528);
or U1905 (N_1905,In_20,In_734);
nand U1906 (N_1906,In_27,In_247);
or U1907 (N_1907,In_141,In_653);
nand U1908 (N_1908,In_395,In_522);
nor U1909 (N_1909,In_475,In_674);
or U1910 (N_1910,In_196,In_745);
and U1911 (N_1911,In_417,In_13);
or U1912 (N_1912,In_624,In_513);
nand U1913 (N_1913,In_309,In_695);
and U1914 (N_1914,In_624,In_281);
nor U1915 (N_1915,In_129,In_334);
nand U1916 (N_1916,In_434,In_581);
nor U1917 (N_1917,In_637,In_425);
or U1918 (N_1918,In_166,In_679);
nand U1919 (N_1919,In_105,In_252);
or U1920 (N_1920,In_379,In_411);
and U1921 (N_1921,In_579,In_218);
nor U1922 (N_1922,In_529,In_638);
nand U1923 (N_1923,In_170,In_707);
xor U1924 (N_1924,In_684,In_51);
and U1925 (N_1925,In_687,In_564);
and U1926 (N_1926,In_621,In_453);
or U1927 (N_1927,In_564,In_597);
nand U1928 (N_1928,In_462,In_500);
nand U1929 (N_1929,In_592,In_516);
nor U1930 (N_1930,In_546,In_175);
nand U1931 (N_1931,In_147,In_85);
nand U1932 (N_1932,In_681,In_688);
nor U1933 (N_1933,In_572,In_716);
and U1934 (N_1934,In_117,In_308);
nor U1935 (N_1935,In_376,In_25);
nor U1936 (N_1936,In_203,In_93);
or U1937 (N_1937,In_643,In_11);
and U1938 (N_1938,In_594,In_602);
nand U1939 (N_1939,In_606,In_322);
nor U1940 (N_1940,In_74,In_424);
nand U1941 (N_1941,In_553,In_648);
or U1942 (N_1942,In_371,In_10);
nor U1943 (N_1943,In_539,In_161);
nand U1944 (N_1944,In_437,In_294);
or U1945 (N_1945,In_368,In_149);
or U1946 (N_1946,In_449,In_232);
nand U1947 (N_1947,In_310,In_348);
and U1948 (N_1948,In_713,In_24);
and U1949 (N_1949,In_166,In_240);
or U1950 (N_1950,In_601,In_523);
or U1951 (N_1951,In_372,In_87);
or U1952 (N_1952,In_703,In_97);
and U1953 (N_1953,In_648,In_271);
nand U1954 (N_1954,In_257,In_186);
and U1955 (N_1955,In_579,In_520);
nor U1956 (N_1956,In_429,In_123);
nand U1957 (N_1957,In_433,In_38);
nand U1958 (N_1958,In_130,In_258);
or U1959 (N_1959,In_719,In_517);
or U1960 (N_1960,In_593,In_122);
nand U1961 (N_1961,In_746,In_257);
nor U1962 (N_1962,In_51,In_370);
nand U1963 (N_1963,In_110,In_122);
nand U1964 (N_1964,In_727,In_744);
nor U1965 (N_1965,In_542,In_664);
nand U1966 (N_1966,In_708,In_488);
or U1967 (N_1967,In_233,In_417);
xnor U1968 (N_1968,In_193,In_677);
and U1969 (N_1969,In_47,In_447);
nand U1970 (N_1970,In_304,In_163);
nand U1971 (N_1971,In_336,In_272);
nor U1972 (N_1972,In_527,In_181);
nand U1973 (N_1973,In_38,In_174);
or U1974 (N_1974,In_96,In_580);
and U1975 (N_1975,In_193,In_648);
and U1976 (N_1976,In_709,In_217);
or U1977 (N_1977,In_424,In_478);
nor U1978 (N_1978,In_525,In_641);
nor U1979 (N_1979,In_209,In_598);
or U1980 (N_1980,In_103,In_412);
nor U1981 (N_1981,In_420,In_731);
or U1982 (N_1982,In_105,In_463);
nor U1983 (N_1983,In_307,In_645);
and U1984 (N_1984,In_397,In_411);
nand U1985 (N_1985,In_348,In_711);
or U1986 (N_1986,In_409,In_332);
nand U1987 (N_1987,In_421,In_686);
or U1988 (N_1988,In_566,In_71);
nand U1989 (N_1989,In_44,In_734);
or U1990 (N_1990,In_659,In_672);
nor U1991 (N_1991,In_156,In_194);
and U1992 (N_1992,In_270,In_34);
nand U1993 (N_1993,In_501,In_125);
nand U1994 (N_1994,In_458,In_612);
nor U1995 (N_1995,In_579,In_532);
nand U1996 (N_1996,In_699,In_587);
nor U1997 (N_1997,In_531,In_592);
nand U1998 (N_1998,In_235,In_297);
or U1999 (N_1999,In_632,In_122);
or U2000 (N_2000,In_445,In_271);
nor U2001 (N_2001,In_152,In_514);
or U2002 (N_2002,In_514,In_522);
nand U2003 (N_2003,In_509,In_255);
nor U2004 (N_2004,In_423,In_209);
and U2005 (N_2005,In_496,In_508);
nor U2006 (N_2006,In_470,In_482);
nor U2007 (N_2007,In_483,In_660);
and U2008 (N_2008,In_33,In_408);
or U2009 (N_2009,In_482,In_109);
nor U2010 (N_2010,In_46,In_388);
nor U2011 (N_2011,In_568,In_418);
and U2012 (N_2012,In_569,In_545);
or U2013 (N_2013,In_571,In_462);
nor U2014 (N_2014,In_64,In_552);
and U2015 (N_2015,In_40,In_320);
or U2016 (N_2016,In_370,In_137);
and U2017 (N_2017,In_233,In_206);
or U2018 (N_2018,In_115,In_687);
nor U2019 (N_2019,In_147,In_686);
or U2020 (N_2020,In_567,In_686);
or U2021 (N_2021,In_375,In_23);
or U2022 (N_2022,In_383,In_116);
nor U2023 (N_2023,In_378,In_352);
or U2024 (N_2024,In_296,In_558);
nor U2025 (N_2025,In_190,In_344);
nor U2026 (N_2026,In_663,In_433);
or U2027 (N_2027,In_462,In_661);
nand U2028 (N_2028,In_376,In_172);
nor U2029 (N_2029,In_161,In_129);
or U2030 (N_2030,In_561,In_299);
nand U2031 (N_2031,In_558,In_133);
and U2032 (N_2032,In_583,In_14);
nand U2033 (N_2033,In_616,In_708);
nor U2034 (N_2034,In_517,In_204);
and U2035 (N_2035,In_198,In_728);
or U2036 (N_2036,In_332,In_360);
or U2037 (N_2037,In_316,In_550);
nor U2038 (N_2038,In_655,In_646);
nor U2039 (N_2039,In_585,In_622);
or U2040 (N_2040,In_368,In_192);
or U2041 (N_2041,In_92,In_81);
nand U2042 (N_2042,In_233,In_443);
nor U2043 (N_2043,In_489,In_502);
or U2044 (N_2044,In_87,In_31);
and U2045 (N_2045,In_162,In_407);
nor U2046 (N_2046,In_384,In_586);
and U2047 (N_2047,In_559,In_284);
or U2048 (N_2048,In_475,In_616);
nor U2049 (N_2049,In_299,In_583);
nand U2050 (N_2050,In_284,In_17);
nand U2051 (N_2051,In_77,In_245);
or U2052 (N_2052,In_499,In_478);
nor U2053 (N_2053,In_447,In_258);
nor U2054 (N_2054,In_678,In_390);
or U2055 (N_2055,In_427,In_688);
nor U2056 (N_2056,In_645,In_610);
nor U2057 (N_2057,In_652,In_75);
xor U2058 (N_2058,In_480,In_337);
or U2059 (N_2059,In_515,In_442);
nand U2060 (N_2060,In_193,In_160);
nor U2061 (N_2061,In_521,In_106);
nor U2062 (N_2062,In_34,In_511);
nor U2063 (N_2063,In_396,In_32);
xor U2064 (N_2064,In_539,In_203);
nor U2065 (N_2065,In_623,In_566);
nor U2066 (N_2066,In_711,In_476);
and U2067 (N_2067,In_201,In_572);
nand U2068 (N_2068,In_480,In_99);
nor U2069 (N_2069,In_110,In_465);
or U2070 (N_2070,In_395,In_13);
or U2071 (N_2071,In_505,In_648);
and U2072 (N_2072,In_614,In_391);
and U2073 (N_2073,In_37,In_369);
nor U2074 (N_2074,In_439,In_312);
or U2075 (N_2075,In_423,In_306);
nor U2076 (N_2076,In_317,In_589);
nand U2077 (N_2077,In_741,In_523);
nor U2078 (N_2078,In_443,In_226);
or U2079 (N_2079,In_462,In_518);
or U2080 (N_2080,In_179,In_186);
xnor U2081 (N_2081,In_571,In_742);
nor U2082 (N_2082,In_78,In_549);
nand U2083 (N_2083,In_432,In_218);
and U2084 (N_2084,In_417,In_505);
and U2085 (N_2085,In_422,In_478);
and U2086 (N_2086,In_49,In_482);
or U2087 (N_2087,In_721,In_710);
nor U2088 (N_2088,In_257,In_535);
nand U2089 (N_2089,In_122,In_131);
nor U2090 (N_2090,In_607,In_641);
xnor U2091 (N_2091,In_727,In_514);
or U2092 (N_2092,In_74,In_167);
nand U2093 (N_2093,In_394,In_317);
or U2094 (N_2094,In_719,In_745);
or U2095 (N_2095,In_434,In_117);
nand U2096 (N_2096,In_382,In_263);
nor U2097 (N_2097,In_521,In_86);
and U2098 (N_2098,In_670,In_129);
nand U2099 (N_2099,In_427,In_439);
and U2100 (N_2100,In_238,In_404);
and U2101 (N_2101,In_678,In_719);
nor U2102 (N_2102,In_564,In_89);
and U2103 (N_2103,In_170,In_325);
or U2104 (N_2104,In_257,In_233);
and U2105 (N_2105,In_273,In_608);
nor U2106 (N_2106,In_18,In_458);
and U2107 (N_2107,In_174,In_219);
and U2108 (N_2108,In_598,In_557);
or U2109 (N_2109,In_105,In_442);
nand U2110 (N_2110,In_698,In_234);
or U2111 (N_2111,In_139,In_390);
nor U2112 (N_2112,In_394,In_350);
and U2113 (N_2113,In_106,In_249);
nor U2114 (N_2114,In_738,In_151);
and U2115 (N_2115,In_108,In_448);
nor U2116 (N_2116,In_156,In_423);
nor U2117 (N_2117,In_122,In_648);
nor U2118 (N_2118,In_169,In_25);
or U2119 (N_2119,In_18,In_208);
and U2120 (N_2120,In_118,In_563);
and U2121 (N_2121,In_514,In_254);
nor U2122 (N_2122,In_315,In_242);
or U2123 (N_2123,In_58,In_514);
and U2124 (N_2124,In_139,In_237);
nor U2125 (N_2125,In_20,In_145);
and U2126 (N_2126,In_128,In_566);
nor U2127 (N_2127,In_519,In_83);
and U2128 (N_2128,In_229,In_258);
and U2129 (N_2129,In_246,In_501);
nand U2130 (N_2130,In_187,In_575);
or U2131 (N_2131,In_231,In_529);
and U2132 (N_2132,In_84,In_419);
and U2133 (N_2133,In_263,In_106);
nor U2134 (N_2134,In_270,In_435);
nor U2135 (N_2135,In_690,In_472);
nand U2136 (N_2136,In_564,In_253);
and U2137 (N_2137,In_22,In_470);
nand U2138 (N_2138,In_382,In_390);
or U2139 (N_2139,In_236,In_179);
nor U2140 (N_2140,In_187,In_110);
nand U2141 (N_2141,In_165,In_14);
and U2142 (N_2142,In_79,In_744);
and U2143 (N_2143,In_43,In_388);
and U2144 (N_2144,In_325,In_575);
nand U2145 (N_2145,In_5,In_676);
or U2146 (N_2146,In_190,In_683);
nor U2147 (N_2147,In_612,In_652);
nand U2148 (N_2148,In_603,In_632);
or U2149 (N_2149,In_665,In_303);
or U2150 (N_2150,In_433,In_538);
and U2151 (N_2151,In_500,In_489);
and U2152 (N_2152,In_402,In_73);
nand U2153 (N_2153,In_189,In_664);
or U2154 (N_2154,In_585,In_247);
nor U2155 (N_2155,In_224,In_223);
nand U2156 (N_2156,In_352,In_595);
or U2157 (N_2157,In_155,In_698);
and U2158 (N_2158,In_366,In_130);
nand U2159 (N_2159,In_642,In_137);
nand U2160 (N_2160,In_220,In_498);
nand U2161 (N_2161,In_248,In_266);
or U2162 (N_2162,In_198,In_290);
or U2163 (N_2163,In_75,In_434);
nor U2164 (N_2164,In_637,In_585);
nand U2165 (N_2165,In_564,In_49);
nand U2166 (N_2166,In_394,In_6);
or U2167 (N_2167,In_681,In_377);
and U2168 (N_2168,In_592,In_553);
nor U2169 (N_2169,In_187,In_197);
or U2170 (N_2170,In_611,In_266);
nor U2171 (N_2171,In_90,In_452);
nor U2172 (N_2172,In_363,In_56);
and U2173 (N_2173,In_121,In_259);
or U2174 (N_2174,In_374,In_291);
nand U2175 (N_2175,In_335,In_659);
and U2176 (N_2176,In_306,In_588);
nand U2177 (N_2177,In_438,In_284);
or U2178 (N_2178,In_407,In_256);
or U2179 (N_2179,In_479,In_223);
or U2180 (N_2180,In_116,In_533);
nor U2181 (N_2181,In_190,In_508);
nand U2182 (N_2182,In_398,In_21);
and U2183 (N_2183,In_64,In_432);
and U2184 (N_2184,In_263,In_463);
and U2185 (N_2185,In_337,In_553);
and U2186 (N_2186,In_127,In_348);
nand U2187 (N_2187,In_207,In_375);
and U2188 (N_2188,In_266,In_136);
and U2189 (N_2189,In_613,In_588);
or U2190 (N_2190,In_703,In_129);
nand U2191 (N_2191,In_63,In_404);
nor U2192 (N_2192,In_201,In_747);
or U2193 (N_2193,In_236,In_3);
or U2194 (N_2194,In_243,In_742);
and U2195 (N_2195,In_108,In_175);
nor U2196 (N_2196,In_0,In_605);
and U2197 (N_2197,In_413,In_489);
nand U2198 (N_2198,In_342,In_638);
nand U2199 (N_2199,In_612,In_628);
and U2200 (N_2200,In_94,In_352);
nor U2201 (N_2201,In_443,In_34);
or U2202 (N_2202,In_48,In_17);
nor U2203 (N_2203,In_734,In_459);
or U2204 (N_2204,In_680,In_10);
nor U2205 (N_2205,In_496,In_259);
and U2206 (N_2206,In_658,In_151);
nand U2207 (N_2207,In_733,In_697);
and U2208 (N_2208,In_459,In_505);
nand U2209 (N_2209,In_352,In_367);
or U2210 (N_2210,In_356,In_495);
nand U2211 (N_2211,In_607,In_222);
and U2212 (N_2212,In_112,In_91);
nand U2213 (N_2213,In_739,In_498);
and U2214 (N_2214,In_17,In_213);
nor U2215 (N_2215,In_435,In_444);
nand U2216 (N_2216,In_378,In_542);
or U2217 (N_2217,In_370,In_738);
or U2218 (N_2218,In_60,In_310);
and U2219 (N_2219,In_239,In_324);
and U2220 (N_2220,In_201,In_598);
nor U2221 (N_2221,In_481,In_11);
and U2222 (N_2222,In_564,In_244);
or U2223 (N_2223,In_691,In_329);
and U2224 (N_2224,In_720,In_48);
nand U2225 (N_2225,In_530,In_689);
or U2226 (N_2226,In_432,In_472);
nor U2227 (N_2227,In_481,In_631);
nand U2228 (N_2228,In_326,In_362);
nand U2229 (N_2229,In_420,In_432);
nand U2230 (N_2230,In_273,In_141);
or U2231 (N_2231,In_729,In_683);
nor U2232 (N_2232,In_210,In_276);
nand U2233 (N_2233,In_337,In_488);
or U2234 (N_2234,In_554,In_334);
nand U2235 (N_2235,In_470,In_630);
and U2236 (N_2236,In_469,In_584);
or U2237 (N_2237,In_616,In_601);
and U2238 (N_2238,In_40,In_601);
nand U2239 (N_2239,In_637,In_88);
or U2240 (N_2240,In_295,In_150);
nand U2241 (N_2241,In_704,In_457);
or U2242 (N_2242,In_525,In_708);
nor U2243 (N_2243,In_261,In_564);
nor U2244 (N_2244,In_347,In_492);
nor U2245 (N_2245,In_277,In_211);
nor U2246 (N_2246,In_505,In_528);
and U2247 (N_2247,In_457,In_637);
nand U2248 (N_2248,In_127,In_353);
nor U2249 (N_2249,In_319,In_279);
or U2250 (N_2250,In_348,In_66);
nor U2251 (N_2251,In_592,In_249);
xor U2252 (N_2252,In_683,In_420);
nand U2253 (N_2253,In_713,In_653);
and U2254 (N_2254,In_83,In_249);
and U2255 (N_2255,In_464,In_600);
and U2256 (N_2256,In_325,In_498);
nand U2257 (N_2257,In_600,In_432);
nand U2258 (N_2258,In_163,In_473);
nand U2259 (N_2259,In_122,In_84);
nor U2260 (N_2260,In_729,In_83);
nand U2261 (N_2261,In_493,In_256);
nand U2262 (N_2262,In_210,In_570);
and U2263 (N_2263,In_421,In_659);
and U2264 (N_2264,In_86,In_297);
and U2265 (N_2265,In_517,In_399);
or U2266 (N_2266,In_243,In_102);
nor U2267 (N_2267,In_382,In_327);
and U2268 (N_2268,In_443,In_480);
nand U2269 (N_2269,In_685,In_378);
or U2270 (N_2270,In_13,In_415);
and U2271 (N_2271,In_712,In_714);
nor U2272 (N_2272,In_7,In_420);
nand U2273 (N_2273,In_90,In_437);
nand U2274 (N_2274,In_701,In_181);
or U2275 (N_2275,In_4,In_28);
and U2276 (N_2276,In_298,In_264);
and U2277 (N_2277,In_370,In_504);
and U2278 (N_2278,In_399,In_299);
nor U2279 (N_2279,In_92,In_102);
and U2280 (N_2280,In_429,In_193);
or U2281 (N_2281,In_480,In_118);
nor U2282 (N_2282,In_623,In_218);
nand U2283 (N_2283,In_484,In_603);
nor U2284 (N_2284,In_564,In_594);
nand U2285 (N_2285,In_676,In_405);
nand U2286 (N_2286,In_703,In_39);
or U2287 (N_2287,In_59,In_424);
nor U2288 (N_2288,In_570,In_666);
and U2289 (N_2289,In_716,In_517);
nor U2290 (N_2290,In_455,In_211);
nand U2291 (N_2291,In_255,In_99);
and U2292 (N_2292,In_403,In_161);
nor U2293 (N_2293,In_539,In_331);
nor U2294 (N_2294,In_704,In_333);
and U2295 (N_2295,In_129,In_312);
nand U2296 (N_2296,In_677,In_184);
nand U2297 (N_2297,In_552,In_529);
or U2298 (N_2298,In_74,In_18);
nor U2299 (N_2299,In_646,In_573);
nand U2300 (N_2300,In_31,In_283);
nor U2301 (N_2301,In_745,In_303);
or U2302 (N_2302,In_560,In_35);
nand U2303 (N_2303,In_46,In_674);
or U2304 (N_2304,In_14,In_126);
or U2305 (N_2305,In_187,In_436);
nor U2306 (N_2306,In_480,In_304);
or U2307 (N_2307,In_503,In_6);
nor U2308 (N_2308,In_508,In_583);
nand U2309 (N_2309,In_245,In_380);
or U2310 (N_2310,In_335,In_325);
nand U2311 (N_2311,In_612,In_422);
or U2312 (N_2312,In_672,In_151);
nor U2313 (N_2313,In_474,In_168);
and U2314 (N_2314,In_688,In_471);
or U2315 (N_2315,In_715,In_43);
and U2316 (N_2316,In_663,In_684);
or U2317 (N_2317,In_255,In_167);
nand U2318 (N_2318,In_721,In_78);
xor U2319 (N_2319,In_579,In_435);
nor U2320 (N_2320,In_60,In_744);
nand U2321 (N_2321,In_356,In_594);
nor U2322 (N_2322,In_535,In_233);
nand U2323 (N_2323,In_375,In_494);
or U2324 (N_2324,In_30,In_504);
nand U2325 (N_2325,In_613,In_682);
and U2326 (N_2326,In_479,In_39);
xnor U2327 (N_2327,In_448,In_149);
nor U2328 (N_2328,In_204,In_320);
nor U2329 (N_2329,In_8,In_87);
or U2330 (N_2330,In_731,In_25);
nand U2331 (N_2331,In_627,In_723);
or U2332 (N_2332,In_425,In_266);
or U2333 (N_2333,In_669,In_163);
nor U2334 (N_2334,In_265,In_514);
and U2335 (N_2335,In_326,In_316);
and U2336 (N_2336,In_578,In_262);
and U2337 (N_2337,In_595,In_18);
and U2338 (N_2338,In_388,In_353);
or U2339 (N_2339,In_81,In_110);
nand U2340 (N_2340,In_77,In_92);
nand U2341 (N_2341,In_163,In_338);
and U2342 (N_2342,In_382,In_683);
nand U2343 (N_2343,In_329,In_281);
and U2344 (N_2344,In_413,In_311);
or U2345 (N_2345,In_20,In_195);
nand U2346 (N_2346,In_246,In_266);
and U2347 (N_2347,In_3,In_73);
and U2348 (N_2348,In_425,In_707);
nand U2349 (N_2349,In_599,In_346);
or U2350 (N_2350,In_720,In_700);
or U2351 (N_2351,In_574,In_17);
nand U2352 (N_2352,In_476,In_297);
or U2353 (N_2353,In_623,In_192);
and U2354 (N_2354,In_120,In_18);
and U2355 (N_2355,In_475,In_175);
and U2356 (N_2356,In_88,In_622);
and U2357 (N_2357,In_565,In_323);
nand U2358 (N_2358,In_547,In_452);
nor U2359 (N_2359,In_572,In_446);
nor U2360 (N_2360,In_197,In_321);
and U2361 (N_2361,In_133,In_560);
and U2362 (N_2362,In_435,In_229);
and U2363 (N_2363,In_145,In_636);
nor U2364 (N_2364,In_525,In_160);
and U2365 (N_2365,In_181,In_230);
nor U2366 (N_2366,In_534,In_148);
and U2367 (N_2367,In_45,In_176);
and U2368 (N_2368,In_241,In_178);
or U2369 (N_2369,In_606,In_219);
nand U2370 (N_2370,In_104,In_43);
or U2371 (N_2371,In_249,In_452);
and U2372 (N_2372,In_400,In_222);
nor U2373 (N_2373,In_136,In_196);
nand U2374 (N_2374,In_698,In_107);
or U2375 (N_2375,In_353,In_500);
or U2376 (N_2376,In_91,In_98);
nor U2377 (N_2377,In_119,In_223);
nor U2378 (N_2378,In_88,In_656);
or U2379 (N_2379,In_728,In_98);
or U2380 (N_2380,In_461,In_649);
or U2381 (N_2381,In_99,In_690);
nand U2382 (N_2382,In_651,In_18);
nor U2383 (N_2383,In_219,In_465);
and U2384 (N_2384,In_83,In_176);
nand U2385 (N_2385,In_625,In_66);
nor U2386 (N_2386,In_63,In_143);
and U2387 (N_2387,In_518,In_314);
nor U2388 (N_2388,In_352,In_148);
and U2389 (N_2389,In_259,In_590);
nand U2390 (N_2390,In_488,In_31);
nor U2391 (N_2391,In_305,In_61);
nand U2392 (N_2392,In_593,In_429);
nand U2393 (N_2393,In_648,In_77);
or U2394 (N_2394,In_451,In_244);
nand U2395 (N_2395,In_615,In_96);
nand U2396 (N_2396,In_5,In_417);
and U2397 (N_2397,In_642,In_66);
nor U2398 (N_2398,In_14,In_210);
nor U2399 (N_2399,In_85,In_500);
nor U2400 (N_2400,In_626,In_100);
nor U2401 (N_2401,In_130,In_704);
and U2402 (N_2402,In_178,In_251);
nand U2403 (N_2403,In_97,In_430);
and U2404 (N_2404,In_484,In_738);
nand U2405 (N_2405,In_727,In_446);
and U2406 (N_2406,In_702,In_29);
nand U2407 (N_2407,In_35,In_76);
nand U2408 (N_2408,In_737,In_293);
nor U2409 (N_2409,In_113,In_412);
or U2410 (N_2410,In_589,In_401);
xnor U2411 (N_2411,In_681,In_189);
and U2412 (N_2412,In_341,In_310);
nor U2413 (N_2413,In_71,In_628);
nand U2414 (N_2414,In_109,In_635);
nor U2415 (N_2415,In_219,In_661);
or U2416 (N_2416,In_589,In_222);
or U2417 (N_2417,In_396,In_257);
or U2418 (N_2418,In_683,In_61);
nor U2419 (N_2419,In_188,In_111);
and U2420 (N_2420,In_201,In_413);
or U2421 (N_2421,In_71,In_400);
or U2422 (N_2422,In_550,In_16);
nand U2423 (N_2423,In_230,In_128);
and U2424 (N_2424,In_281,In_134);
and U2425 (N_2425,In_616,In_122);
and U2426 (N_2426,In_366,In_473);
nor U2427 (N_2427,In_335,In_75);
or U2428 (N_2428,In_314,In_141);
nor U2429 (N_2429,In_481,In_156);
or U2430 (N_2430,In_653,In_548);
or U2431 (N_2431,In_223,In_346);
and U2432 (N_2432,In_11,In_707);
or U2433 (N_2433,In_177,In_376);
and U2434 (N_2434,In_494,In_374);
nor U2435 (N_2435,In_164,In_9);
nand U2436 (N_2436,In_675,In_76);
nor U2437 (N_2437,In_438,In_683);
nand U2438 (N_2438,In_409,In_284);
xnor U2439 (N_2439,In_484,In_454);
and U2440 (N_2440,In_48,In_245);
or U2441 (N_2441,In_123,In_515);
or U2442 (N_2442,In_490,In_413);
nor U2443 (N_2443,In_346,In_83);
nor U2444 (N_2444,In_621,In_242);
and U2445 (N_2445,In_239,In_347);
nor U2446 (N_2446,In_463,In_390);
and U2447 (N_2447,In_160,In_24);
nand U2448 (N_2448,In_56,In_724);
nor U2449 (N_2449,In_362,In_512);
nand U2450 (N_2450,In_81,In_511);
and U2451 (N_2451,In_606,In_358);
nor U2452 (N_2452,In_527,In_691);
nor U2453 (N_2453,In_582,In_205);
nand U2454 (N_2454,In_345,In_209);
nor U2455 (N_2455,In_224,In_536);
and U2456 (N_2456,In_601,In_284);
and U2457 (N_2457,In_236,In_193);
nand U2458 (N_2458,In_10,In_443);
nand U2459 (N_2459,In_192,In_563);
or U2460 (N_2460,In_579,In_377);
and U2461 (N_2461,In_292,In_687);
nor U2462 (N_2462,In_654,In_187);
nand U2463 (N_2463,In_136,In_413);
nor U2464 (N_2464,In_709,In_175);
nor U2465 (N_2465,In_697,In_604);
nand U2466 (N_2466,In_91,In_254);
and U2467 (N_2467,In_286,In_50);
or U2468 (N_2468,In_589,In_104);
nand U2469 (N_2469,In_257,In_57);
nor U2470 (N_2470,In_207,In_586);
and U2471 (N_2471,In_190,In_596);
and U2472 (N_2472,In_378,In_280);
or U2473 (N_2473,In_86,In_450);
and U2474 (N_2474,In_491,In_95);
nor U2475 (N_2475,In_653,In_541);
nor U2476 (N_2476,In_377,In_168);
or U2477 (N_2477,In_597,In_416);
nor U2478 (N_2478,In_445,In_456);
and U2479 (N_2479,In_344,In_8);
nor U2480 (N_2480,In_728,In_349);
nor U2481 (N_2481,In_708,In_261);
and U2482 (N_2482,In_154,In_418);
or U2483 (N_2483,In_129,In_408);
or U2484 (N_2484,In_575,In_322);
nor U2485 (N_2485,In_543,In_37);
nand U2486 (N_2486,In_460,In_436);
or U2487 (N_2487,In_153,In_90);
xor U2488 (N_2488,In_213,In_2);
and U2489 (N_2489,In_339,In_60);
nor U2490 (N_2490,In_304,In_69);
nand U2491 (N_2491,In_259,In_613);
nor U2492 (N_2492,In_710,In_46);
or U2493 (N_2493,In_470,In_422);
nor U2494 (N_2494,In_181,In_659);
nor U2495 (N_2495,In_298,In_560);
nor U2496 (N_2496,In_91,In_51);
or U2497 (N_2497,In_713,In_163);
nand U2498 (N_2498,In_646,In_451);
nand U2499 (N_2499,In_491,In_317);
xnor U2500 (N_2500,N_296,N_1874);
nand U2501 (N_2501,N_1324,N_2388);
nand U2502 (N_2502,N_415,N_2092);
nor U2503 (N_2503,N_459,N_1191);
nand U2504 (N_2504,N_309,N_504);
nor U2505 (N_2505,N_2219,N_1077);
or U2506 (N_2506,N_1108,N_878);
nor U2507 (N_2507,N_351,N_38);
nor U2508 (N_2508,N_1850,N_2425);
and U2509 (N_2509,N_905,N_1312);
and U2510 (N_2510,N_1884,N_236);
and U2511 (N_2511,N_791,N_397);
nor U2512 (N_2512,N_961,N_1728);
nor U2513 (N_2513,N_2022,N_740);
and U2514 (N_2514,N_1352,N_1970);
or U2515 (N_2515,N_1896,N_1437);
or U2516 (N_2516,N_2147,N_1630);
nand U2517 (N_2517,N_2046,N_2368);
nor U2518 (N_2518,N_411,N_124);
and U2519 (N_2519,N_1286,N_175);
or U2520 (N_2520,N_1549,N_1729);
and U2521 (N_2521,N_508,N_10);
or U2522 (N_2522,N_63,N_538);
nand U2523 (N_2523,N_171,N_42);
xor U2524 (N_2524,N_1488,N_1635);
xor U2525 (N_2525,N_409,N_1112);
or U2526 (N_2526,N_1989,N_2261);
or U2527 (N_2527,N_938,N_325);
nor U2528 (N_2528,N_807,N_2314);
or U2529 (N_2529,N_2376,N_2190);
and U2530 (N_2530,N_161,N_1861);
nand U2531 (N_2531,N_1341,N_975);
nand U2532 (N_2532,N_1291,N_2077);
nor U2533 (N_2533,N_55,N_378);
or U2534 (N_2534,N_1535,N_1941);
and U2535 (N_2535,N_796,N_1492);
and U2536 (N_2536,N_1576,N_1351);
nand U2537 (N_2537,N_1052,N_652);
and U2538 (N_2538,N_1822,N_1785);
and U2539 (N_2539,N_448,N_2372);
nor U2540 (N_2540,N_453,N_748);
nand U2541 (N_2541,N_491,N_637);
nor U2542 (N_2542,N_2484,N_2167);
nand U2543 (N_2543,N_1115,N_1181);
nor U2544 (N_2544,N_385,N_1424);
nor U2545 (N_2545,N_1900,N_1154);
nand U2546 (N_2546,N_2402,N_2462);
nor U2547 (N_2547,N_565,N_1128);
nand U2548 (N_2548,N_1261,N_692);
nor U2549 (N_2549,N_2341,N_1219);
or U2550 (N_2550,N_2440,N_473);
nor U2551 (N_2551,N_853,N_2315);
nand U2552 (N_2552,N_8,N_1572);
or U2553 (N_2553,N_1302,N_726);
or U2554 (N_2554,N_1264,N_2416);
nand U2555 (N_2555,N_836,N_224);
or U2556 (N_2556,N_737,N_1195);
nor U2557 (N_2557,N_300,N_166);
nand U2558 (N_2558,N_29,N_2450);
or U2559 (N_2559,N_2241,N_1168);
nand U2560 (N_2560,N_629,N_139);
and U2561 (N_2561,N_984,N_1918);
nand U2562 (N_2562,N_222,N_380);
or U2563 (N_2563,N_1189,N_2481);
nor U2564 (N_2564,N_1068,N_1173);
and U2565 (N_2565,N_607,N_188);
and U2566 (N_2566,N_1706,N_1987);
and U2567 (N_2567,N_874,N_214);
nand U2568 (N_2568,N_1338,N_1840);
and U2569 (N_2569,N_698,N_2039);
or U2570 (N_2570,N_183,N_90);
or U2571 (N_2571,N_1771,N_2061);
nand U2572 (N_2572,N_2199,N_1726);
nand U2573 (N_2573,N_1369,N_1982);
and U2574 (N_2574,N_290,N_2047);
xnor U2575 (N_2575,N_690,N_2187);
nand U2576 (N_2576,N_1463,N_1713);
xor U2577 (N_2577,N_2268,N_1122);
nand U2578 (N_2578,N_919,N_1548);
or U2579 (N_2579,N_1618,N_2359);
nor U2580 (N_2580,N_1749,N_2114);
nand U2581 (N_2581,N_108,N_1304);
or U2582 (N_2582,N_924,N_1760);
or U2583 (N_2583,N_1695,N_2082);
and U2584 (N_2584,N_1927,N_2421);
and U2585 (N_2585,N_1015,N_2037);
or U2586 (N_2586,N_2446,N_24);
and U2587 (N_2587,N_2374,N_1791);
and U2588 (N_2588,N_1085,N_1620);
nor U2589 (N_2589,N_2439,N_2206);
or U2590 (N_2590,N_1082,N_2493);
and U2591 (N_2591,N_1190,N_1866);
and U2592 (N_2592,N_2191,N_2363);
nor U2593 (N_2593,N_923,N_136);
nor U2594 (N_2594,N_318,N_1904);
and U2595 (N_2595,N_948,N_1836);
nor U2596 (N_2596,N_2429,N_903);
nand U2597 (N_2597,N_1089,N_733);
nand U2598 (N_2598,N_2379,N_1563);
nand U2599 (N_2599,N_277,N_1722);
nand U2600 (N_2600,N_2348,N_1881);
and U2601 (N_2601,N_408,N_254);
nand U2602 (N_2602,N_2021,N_1409);
nand U2603 (N_2603,N_1731,N_1010);
nor U2604 (N_2604,N_1715,N_1960);
and U2605 (N_2605,N_455,N_479);
and U2606 (N_2606,N_799,N_238);
nand U2607 (N_2607,N_729,N_346);
nand U2608 (N_2608,N_1503,N_2267);
and U2609 (N_2609,N_1738,N_1757);
nand U2610 (N_2610,N_1188,N_2119);
or U2611 (N_2611,N_1638,N_2140);
and U2612 (N_2612,N_123,N_876);
nand U2613 (N_2613,N_1629,N_360);
nand U2614 (N_2614,N_78,N_2005);
nand U2615 (N_2615,N_1151,N_304);
or U2616 (N_2616,N_574,N_2085);
nor U2617 (N_2617,N_1837,N_1676);
nor U2618 (N_2618,N_1924,N_977);
nand U2619 (N_2619,N_2016,N_1353);
nand U2620 (N_2620,N_1327,N_1251);
and U2621 (N_2621,N_1395,N_1121);
and U2622 (N_2622,N_1499,N_1818);
nand U2623 (N_2623,N_2424,N_429);
nor U2624 (N_2624,N_2338,N_140);
nand U2625 (N_2625,N_1509,N_1185);
or U2626 (N_2626,N_598,N_410);
nor U2627 (N_2627,N_601,N_2161);
nand U2628 (N_2628,N_1273,N_1864);
and U2629 (N_2629,N_1136,N_332);
or U2630 (N_2630,N_2101,N_520);
xnor U2631 (N_2631,N_592,N_1457);
and U2632 (N_2632,N_1475,N_114);
or U2633 (N_2633,N_2098,N_1510);
and U2634 (N_2634,N_452,N_1674);
nand U2635 (N_2635,N_1092,N_1293);
nor U2636 (N_2636,N_165,N_744);
and U2637 (N_2637,N_1320,N_723);
nand U2638 (N_2638,N_2130,N_1746);
nand U2639 (N_2639,N_2320,N_1875);
xor U2640 (N_2640,N_1282,N_2304);
and U2641 (N_2641,N_1685,N_2323);
or U2642 (N_2642,N_2216,N_105);
or U2643 (N_2643,N_787,N_1595);
nand U2644 (N_2644,N_2486,N_2316);
nand U2645 (N_2645,N_1116,N_1290);
nand U2646 (N_2646,N_1751,N_967);
nand U2647 (N_2647,N_1249,N_1625);
nor U2648 (N_2648,N_329,N_347);
and U2649 (N_2649,N_912,N_344);
and U2650 (N_2650,N_638,N_311);
nand U2651 (N_2651,N_2298,N_1410);
nor U2652 (N_2652,N_827,N_1741);
nand U2653 (N_2653,N_1235,N_635);
nor U2654 (N_2654,N_1654,N_1484);
or U2655 (N_2655,N_1607,N_87);
and U2656 (N_2656,N_2122,N_2185);
nor U2657 (N_2657,N_2257,N_1642);
and U2658 (N_2658,N_252,N_441);
and U2659 (N_2659,N_2043,N_482);
or U2660 (N_2660,N_1171,N_2074);
nor U2661 (N_2661,N_2394,N_2398);
nor U2662 (N_2662,N_1428,N_2070);
nand U2663 (N_2663,N_467,N_1664);
and U2664 (N_2664,N_642,N_2303);
or U2665 (N_2665,N_471,N_1035);
and U2666 (N_2666,N_1434,N_900);
or U2667 (N_2667,N_1794,N_1801);
or U2668 (N_2668,N_1453,N_391);
and U2669 (N_2669,N_417,N_1627);
or U2670 (N_2670,N_1833,N_297);
nand U2671 (N_2671,N_1473,N_321);
nand U2672 (N_2672,N_138,N_851);
nand U2673 (N_2673,N_208,N_669);
and U2674 (N_2674,N_686,N_2286);
nor U2675 (N_2675,N_2210,N_1272);
nand U2676 (N_2676,N_1634,N_1949);
nor U2677 (N_2677,N_1955,N_627);
or U2678 (N_2678,N_1003,N_1455);
nand U2679 (N_2679,N_1934,N_272);
or U2680 (N_2680,N_1540,N_187);
nor U2681 (N_2681,N_22,N_317);
or U2682 (N_2682,N_783,N_2221);
nand U2683 (N_2683,N_798,N_2136);
and U2684 (N_2684,N_1311,N_256);
or U2685 (N_2685,N_1610,N_2271);
and U2686 (N_2686,N_2020,N_602);
nand U2687 (N_2687,N_1187,N_440);
nor U2688 (N_2688,N_267,N_1787);
nand U2689 (N_2689,N_894,N_566);
and U2690 (N_2690,N_2213,N_1065);
nand U2691 (N_2691,N_357,N_469);
nor U2692 (N_2692,N_530,N_819);
and U2693 (N_2693,N_1464,N_929);
nand U2694 (N_2694,N_1201,N_1521);
and U2695 (N_2695,N_1469,N_1977);
nand U2696 (N_2696,N_1919,N_197);
nor U2697 (N_2697,N_1231,N_1343);
nor U2698 (N_2698,N_1640,N_1334);
nand U2699 (N_2699,N_1470,N_94);
nor U2700 (N_2700,N_913,N_562);
nor U2701 (N_2701,N_1846,N_680);
nor U2702 (N_2702,N_625,N_115);
and U2703 (N_2703,N_863,N_199);
nand U2704 (N_2704,N_2002,N_1339);
and U2705 (N_2705,N_1933,N_835);
nand U2706 (N_2706,N_2109,N_2365);
and U2707 (N_2707,N_1662,N_1124);
nor U2708 (N_2708,N_1018,N_1360);
nor U2709 (N_2709,N_1717,N_1332);
nand U2710 (N_2710,N_1347,N_618);
nor U2711 (N_2711,N_2311,N_1345);
or U2712 (N_2712,N_728,N_2053);
nand U2713 (N_2713,N_1700,N_595);
and U2714 (N_2714,N_1669,N_763);
or U2715 (N_2715,N_1718,N_1930);
and U2716 (N_2716,N_61,N_275);
and U2717 (N_2717,N_1340,N_2204);
nor U2718 (N_2718,N_2103,N_2292);
and U2719 (N_2719,N_922,N_2285);
or U2720 (N_2720,N_2117,N_1914);
nor U2721 (N_2721,N_387,N_2473);
and U2722 (N_2722,N_1845,N_1598);
and U2723 (N_2723,N_586,N_969);
or U2724 (N_2724,N_72,N_1416);
or U2725 (N_2725,N_785,N_1587);
and U2726 (N_2726,N_1218,N_2050);
nor U2727 (N_2727,N_2351,N_591);
nand U2728 (N_2728,N_1232,N_1023);
or U2729 (N_2729,N_615,N_2015);
nand U2730 (N_2730,N_2313,N_1276);
xor U2731 (N_2731,N_1009,N_964);
or U2732 (N_2732,N_892,N_192);
nor U2733 (N_2733,N_67,N_31);
nor U2734 (N_2734,N_872,N_1140);
and U2735 (N_2735,N_456,N_978);
or U2736 (N_2736,N_2243,N_493);
nor U2737 (N_2737,N_2404,N_1910);
and U2738 (N_2738,N_323,N_789);
and U2739 (N_2739,N_1995,N_769);
or U2740 (N_2740,N_1940,N_2356);
nor U2741 (N_2741,N_462,N_1752);
and U2742 (N_2742,N_1800,N_997);
xor U2743 (N_2743,N_2225,N_877);
or U2744 (N_2744,N_1579,N_2203);
nor U2745 (N_2745,N_1570,N_69);
nand U2746 (N_2746,N_676,N_1011);
and U2747 (N_2747,N_849,N_1078);
xnor U2748 (N_2748,N_2346,N_1091);
or U2749 (N_2749,N_1277,N_678);
nor U2750 (N_2750,N_416,N_255);
nor U2751 (N_2751,N_1274,N_164);
nor U2752 (N_2752,N_613,N_1971);
nor U2753 (N_2753,N_128,N_1830);
or U2754 (N_2754,N_143,N_1867);
nand U2755 (N_2755,N_710,N_2115);
or U2756 (N_2756,N_1271,N_291);
nor U2757 (N_2757,N_1820,N_2399);
nor U2758 (N_2758,N_279,N_965);
nor U2759 (N_2759,N_492,N_389);
nand U2760 (N_2760,N_376,N_1908);
nand U2761 (N_2761,N_881,N_2383);
nand U2762 (N_2762,N_1043,N_2441);
and U2763 (N_2763,N_1478,N_1139);
and U2764 (N_2764,N_589,N_741);
and U2765 (N_2765,N_1532,N_264);
nand U2766 (N_2766,N_20,N_281);
nand U2767 (N_2767,N_1725,N_1421);
or U2768 (N_2768,N_1034,N_2266);
or U2769 (N_2769,N_65,N_1044);
nor U2770 (N_2770,N_1692,N_1902);
nor U2771 (N_2771,N_213,N_1056);
nand U2772 (N_2772,N_1436,N_2017);
nand U2773 (N_2773,N_1118,N_1883);
or U2774 (N_2774,N_1593,N_730);
nand U2775 (N_2775,N_2168,N_1710);
nor U2776 (N_2776,N_1193,N_2469);
or U2777 (N_2777,N_1542,N_982);
and U2778 (N_2778,N_1066,N_1917);
nor U2779 (N_2779,N_2062,N_112);
or U2780 (N_2780,N_767,N_1423);
or U2781 (N_2781,N_246,N_1240);
or U2782 (N_2782,N_372,N_1979);
nand U2783 (N_2783,N_1659,N_821);
and U2784 (N_2784,N_1967,N_1497);
or U2785 (N_2785,N_887,N_298);
or U2786 (N_2786,N_2192,N_424);
and U2787 (N_2787,N_1747,N_612);
or U2788 (N_2788,N_2222,N_1182);
and U2789 (N_2789,N_1086,N_1204);
nor U2790 (N_2790,N_694,N_1442);
or U2791 (N_2791,N_1515,N_1821);
and U2792 (N_2792,N_834,N_910);
nand U2793 (N_2793,N_1809,N_289);
nand U2794 (N_2794,N_1631,N_994);
nand U2795 (N_2795,N_1100,N_1916);
nand U2796 (N_2796,N_1999,N_2143);
nor U2797 (N_2797,N_37,N_2463);
and U2798 (N_2798,N_228,N_1247);
and U2799 (N_2799,N_2453,N_280);
and U2800 (N_2800,N_1458,N_708);
and U2801 (N_2801,N_759,N_914);
and U2802 (N_2802,N_2418,N_2459);
nor U2803 (N_2803,N_2094,N_477);
or U2804 (N_2804,N_1922,N_2112);
and U2805 (N_2805,N_2400,N_1899);
or U2806 (N_2806,N_16,N_1885);
and U2807 (N_2807,N_801,N_830);
and U2808 (N_2808,N_1694,N_181);
nor U2809 (N_2809,N_1359,N_2477);
and U2810 (N_2810,N_2309,N_1407);
nor U2811 (N_2811,N_1248,N_1117);
nor U2812 (N_2812,N_1348,N_691);
or U2813 (N_2813,N_1993,N_1445);
nor U2814 (N_2814,N_1106,N_2442);
and U2815 (N_2815,N_2054,N_671);
nor U2816 (N_2816,N_1931,N_2322);
and U2817 (N_2817,N_2460,N_163);
nor U2818 (N_2818,N_1690,N_616);
nand U2819 (N_2819,N_711,N_1641);
and U2820 (N_2820,N_369,N_2051);
and U2821 (N_2821,N_2283,N_995);
nor U2822 (N_2822,N_365,N_2024);
and U2823 (N_2823,N_1807,N_689);
and U2824 (N_2824,N_1723,N_1712);
nand U2825 (N_2825,N_817,N_1498);
or U2826 (N_2826,N_1857,N_1903);
nand U2827 (N_2827,N_1965,N_2457);
and U2828 (N_2828,N_749,N_1397);
and U2829 (N_2829,N_2164,N_1948);
and U2830 (N_2830,N_1546,N_1824);
nand U2831 (N_2831,N_1553,N_1768);
nor U2832 (N_2832,N_1390,N_1557);
nand U2833 (N_2833,N_2288,N_2166);
or U2834 (N_2834,N_1321,N_2010);
nand U2835 (N_2835,N_1853,N_1670);
and U2836 (N_2836,N_1365,N_303);
and U2837 (N_2837,N_1701,N_2260);
nor U2838 (N_2838,N_2128,N_987);
nand U2839 (N_2839,N_582,N_1370);
nor U2840 (N_2840,N_1755,N_1525);
nor U2841 (N_2841,N_1580,N_2263);
nor U2842 (N_2842,N_621,N_33);
or U2843 (N_2843,N_1594,N_2342);
nand U2844 (N_2844,N_2234,N_925);
or U2845 (N_2845,N_266,N_2397);
nand U2846 (N_2846,N_859,N_1012);
or U2847 (N_2847,N_1789,N_936);
nor U2848 (N_2848,N_648,N_1870);
and U2849 (N_2849,N_1137,N_521);
nor U2850 (N_2850,N_82,N_824);
nand U2851 (N_2851,N_406,N_340);
nor U2852 (N_2852,N_1573,N_662);
and U2853 (N_2853,N_2480,N_1259);
and U2854 (N_2854,N_2104,N_1648);
xor U2855 (N_2855,N_273,N_1632);
nor U2856 (N_2856,N_624,N_2254);
nor U2857 (N_2857,N_1336,N_1149);
nand U2858 (N_2858,N_1939,N_2297);
and U2859 (N_2859,N_839,N_1678);
nand U2860 (N_2860,N_237,N_433);
or U2861 (N_2861,N_156,N_927);
and U2862 (N_2862,N_867,N_295);
nor U2863 (N_2863,N_1501,N_696);
nand U2864 (N_2864,N_1319,N_498);
or U2865 (N_2865,N_947,N_517);
nand U2866 (N_2866,N_412,N_2034);
nand U2867 (N_2867,N_257,N_949);
and U2868 (N_2868,N_262,N_363);
nor U2869 (N_2869,N_2134,N_2401);
and U2870 (N_2870,N_1220,N_2148);
nor U2871 (N_2871,N_1871,N_575);
nor U2872 (N_2872,N_420,N_77);
nor U2873 (N_2873,N_2223,N_2264);
or U2874 (N_2874,N_971,N_2300);
nor U2875 (N_2875,N_1699,N_2326);
nand U2876 (N_2876,N_402,N_945);
or U2877 (N_2877,N_714,N_720);
nand U2878 (N_2878,N_1687,N_893);
and U2879 (N_2879,N_1257,N_2253);
nor U2880 (N_2880,N_1780,N_675);
and U2881 (N_2881,N_782,N_1008);
nor U2882 (N_2882,N_431,N_2090);
nand U2883 (N_2883,N_2375,N_1819);
and U2884 (N_2884,N_2279,N_1443);
or U2885 (N_2885,N_382,N_11);
and U2886 (N_2886,N_988,N_1138);
nand U2887 (N_2887,N_2494,N_1224);
and U2888 (N_2888,N_2454,N_778);
or U2889 (N_2889,N_1762,N_245);
and U2890 (N_2890,N_2217,N_2328);
or U2891 (N_2891,N_470,N_1180);
nor U2892 (N_2892,N_797,N_2159);
nand U2893 (N_2893,N_223,N_2118);
nor U2894 (N_2894,N_59,N_707);
or U2895 (N_2895,N_644,N_49);
or U2896 (N_2896,N_2412,N_1486);
or U2897 (N_2897,N_1055,N_1668);
nor U2898 (N_2898,N_1493,N_904);
nor U2899 (N_2899,N_1230,N_1774);
nor U2900 (N_2900,N_1465,N_486);
nand U2901 (N_2901,N_1646,N_784);
and U2902 (N_2902,N_1511,N_812);
and U2903 (N_2903,N_1911,N_2042);
or U2904 (N_2904,N_511,N_147);
nor U2905 (N_2905,N_942,N_1992);
nand U2906 (N_2906,N_556,N_1878);
nor U2907 (N_2907,N_917,N_1028);
nand U2908 (N_2908,N_1730,N_2371);
nor U2909 (N_2909,N_2093,N_1682);
or U2910 (N_2910,N_219,N_1179);
or U2911 (N_2911,N_1560,N_1462);
nand U2912 (N_2912,N_559,N_1776);
or U2913 (N_2913,N_2478,N_57);
nand U2914 (N_2914,N_432,N_1408);
and U2915 (N_2915,N_2152,N_2174);
nor U2916 (N_2916,N_64,N_2182);
or U2917 (N_2917,N_1221,N_1344);
nand U2918 (N_2918,N_980,N_1425);
and U2919 (N_2919,N_2445,N_202);
nand U2920 (N_2920,N_954,N_674);
nand U2921 (N_2921,N_972,N_916);
or U2922 (N_2922,N_2242,N_259);
nor U2923 (N_2923,N_1773,N_1355);
nor U2924 (N_2924,N_2492,N_1036);
or U2925 (N_2925,N_585,N_2321);
and U2926 (N_2926,N_225,N_684);
nor U2927 (N_2927,N_1759,N_974);
and U2928 (N_2928,N_1309,N_1412);
and U2929 (N_2929,N_1838,N_702);
and U2930 (N_2930,N_2487,N_557);
nor U2931 (N_2931,N_466,N_1790);
or U2932 (N_2932,N_1767,N_144);
nor U2933 (N_2933,N_1326,N_753);
and U2934 (N_2934,N_717,N_823);
or U2935 (N_2935,N_1337,N_2052);
and U2936 (N_2936,N_1050,N_2461);
and U2937 (N_2937,N_1125,N_2087);
nand U2938 (N_2938,N_1508,N_102);
nor U2939 (N_2939,N_2330,N_1988);
nand U2940 (N_2940,N_73,N_436);
and U2941 (N_2941,N_2198,N_1766);
or U2942 (N_2942,N_1422,N_1539);
nor U2943 (N_2943,N_1667,N_1385);
and U2944 (N_2944,N_1169,N_2048);
and U2945 (N_2945,N_777,N_292);
and U2946 (N_2946,N_345,N_647);
nor U2947 (N_2947,N_1526,N_1313);
nand U2948 (N_2948,N_7,N_1719);
xnor U2949 (N_2949,N_240,N_1920);
or U2950 (N_2950,N_1556,N_2405);
and U2951 (N_2951,N_1087,N_2296);
nor U2952 (N_2952,N_1447,N_896);
nor U2953 (N_2953,N_1483,N_26);
and U2954 (N_2954,N_1624,N_1841);
nand U2955 (N_2955,N_32,N_1996);
and U2956 (N_2956,N_715,N_600);
and U2957 (N_2957,N_1574,N_1049);
nor U2958 (N_2958,N_1227,N_2235);
and U2959 (N_2959,N_560,N_2137);
or U2960 (N_2960,N_172,N_746);
or U2961 (N_2961,N_1175,N_943);
and U2962 (N_2962,N_48,N_885);
nand U2963 (N_2963,N_1450,N_1020);
or U2964 (N_2964,N_818,N_1333);
nor U2965 (N_2965,N_198,N_1957);
nor U2966 (N_2966,N_921,N_2102);
nor U2967 (N_2967,N_307,N_1517);
nand U2968 (N_2968,N_1656,N_952);
and U2969 (N_2969,N_2110,N_203);
nand U2970 (N_2970,N_1157,N_434);
and U2971 (N_2971,N_1358,N_1196);
nor U2972 (N_2972,N_1242,N_1148);
and U2973 (N_2973,N_1782,N_577);
or U2974 (N_2974,N_2007,N_1879);
and U2975 (N_2975,N_1817,N_109);
nand U2976 (N_2976,N_2436,N_2443);
or U2977 (N_2977,N_2170,N_846);
nand U2978 (N_2978,N_1950,N_40);
and U2979 (N_2979,N_1680,N_1233);
and U2980 (N_2980,N_1225,N_1016);
nand U2981 (N_2981,N_447,N_1889);
and U2982 (N_2982,N_705,N_488);
and U2983 (N_2983,N_1522,N_731);
and U2984 (N_2984,N_1859,N_831);
and U2985 (N_2985,N_2369,N_1211);
nand U2986 (N_2986,N_1742,N_1119);
nand U2987 (N_2987,N_472,N_1804);
or U2988 (N_2988,N_709,N_2332);
nor U2989 (N_2989,N_568,N_2458);
nand U2990 (N_2990,N_1222,N_693);
and U2991 (N_2991,N_654,N_771);
and U2992 (N_2992,N_656,N_636);
or U2993 (N_2993,N_883,N_1243);
and U2994 (N_2994,N_2265,N_985);
nor U2995 (N_2995,N_1946,N_401);
or U2996 (N_2996,N_1544,N_908);
nor U2997 (N_2997,N_2003,N_788);
nor U2998 (N_2998,N_185,N_2239);
and U2999 (N_2999,N_107,N_2428);
or U3000 (N_3000,N_2224,N_2189);
and U3001 (N_3001,N_324,N_113);
or U3002 (N_3002,N_1798,N_806);
nand U3003 (N_3003,N_999,N_747);
nand U3004 (N_3004,N_842,N_1460);
nand U3005 (N_3005,N_1200,N_1494);
or U3006 (N_3006,N_1585,N_1854);
nor U3007 (N_3007,N_944,N_1482);
nand U3008 (N_3008,N_1868,N_1547);
nor U3009 (N_3009,N_1714,N_1566);
or U3010 (N_3010,N_71,N_1452);
nand U3011 (N_3011,N_2284,N_1349);
or U3012 (N_3012,N_734,N_840);
nand U3013 (N_3013,N_581,N_1392);
nor U3014 (N_3014,N_500,N_131);
and U3015 (N_3015,N_2000,N_1578);
or U3016 (N_3016,N_1166,N_1006);
nor U3017 (N_3017,N_1551,N_1612);
and U3018 (N_3018,N_1213,N_2269);
or U3019 (N_3019,N_1058,N_2331);
or U3020 (N_3020,N_2419,N_2032);
nand U3021 (N_3021,N_1802,N_1652);
nor U3022 (N_3022,N_2333,N_308);
nor U3023 (N_3023,N_1644,N_992);
nand U3024 (N_3024,N_122,N_152);
nor U3025 (N_3025,N_739,N_56);
and U3026 (N_3026,N_1863,N_1827);
or U3027 (N_3027,N_706,N_1178);
and U3028 (N_3028,N_542,N_204);
nand U3029 (N_3029,N_1250,N_233);
nor U3030 (N_3030,N_398,N_169);
or U3031 (N_3031,N_1912,N_18);
and U3032 (N_3032,N_2361,N_1103);
or U3033 (N_3033,N_1026,N_1301);
or U3034 (N_3034,N_718,N_1698);
nor U3035 (N_3035,N_803,N_926);
or U3036 (N_3036,N_177,N_2012);
and U3037 (N_3037,N_1167,N_328);
nor U3038 (N_3038,N_1490,N_1356);
nor U3039 (N_3039,N_1451,N_512);
or U3040 (N_3040,N_2476,N_1586);
or U3041 (N_3041,N_811,N_231);
nand U3042 (N_3042,N_1316,N_1703);
nor U3043 (N_3043,N_1500,N_2081);
and U3044 (N_3044,N_2420,N_35);
nor U3045 (N_3045,N_2362,N_1582);
and U3046 (N_3046,N_1133,N_735);
or U3047 (N_3047,N_1454,N_1377);
nand U3048 (N_3048,N_549,N_426);
nand U3049 (N_3049,N_770,N_386);
nand U3050 (N_3050,N_721,N_572);
nand U3051 (N_3051,N_173,N_2151);
or U3052 (N_3052,N_132,N_2408);
and U3053 (N_3053,N_2350,N_826);
and U3054 (N_3054,N_953,N_2045);
nor U3055 (N_3055,N_146,N_54);
or U3056 (N_3056,N_1686,N_1727);
nand U3057 (N_3057,N_868,N_1278);
nor U3058 (N_3058,N_1888,N_2277);
and U3059 (N_3059,N_825,N_2238);
nand U3060 (N_3060,N_2100,N_1584);
or U3061 (N_3061,N_2160,N_1696);
nor U3062 (N_3062,N_1506,N_1898);
and U3063 (N_3063,N_23,N_653);
nand U3064 (N_3064,N_1354,N_976);
nand U3065 (N_3065,N_1805,N_1890);
nand U3066 (N_3066,N_320,N_632);
or U3067 (N_3067,N_760,N_2448);
or U3068 (N_3068,N_766,N_776);
nor U3069 (N_3069,N_1985,N_76);
nor U3070 (N_3070,N_1849,N_2030);
or U3071 (N_3071,N_1083,N_2067);
and U3072 (N_3072,N_1502,N_1387);
nor U3073 (N_3073,N_200,N_2305);
or U3074 (N_3074,N_2139,N_2275);
nand U3075 (N_3075,N_2088,N_814);
and U3076 (N_3076,N_1808,N_1516);
nand U3077 (N_3077,N_736,N_1983);
nand U3078 (N_3078,N_2025,N_1843);
nor U3079 (N_3079,N_1440,N_489);
nand U3080 (N_3080,N_2212,N_2466);
nor U3081 (N_3081,N_1990,N_142);
or U3082 (N_3082,N_2135,N_1037);
or U3083 (N_3083,N_2273,N_902);
or U3084 (N_3084,N_2096,N_518);
or U3085 (N_3085,N_781,N_792);
or U3086 (N_3086,N_606,N_1937);
nor U3087 (N_3087,N_1894,N_350);
nor U3088 (N_3088,N_1057,N_1255);
nor U3089 (N_3089,N_155,N_2410);
and U3090 (N_3090,N_590,N_117);
and U3091 (N_3091,N_2497,N_119);
or U3092 (N_3092,N_1367,N_2019);
or U3093 (N_3093,N_438,N_2126);
nor U3094 (N_3094,N_339,N_2073);
or U3095 (N_3095,N_1705,N_1262);
nor U3096 (N_3096,N_1842,N_1310);
or U3097 (N_3097,N_1129,N_879);
and U3098 (N_3098,N_75,N_700);
and U3099 (N_3099,N_1897,N_435);
or U3100 (N_3100,N_1079,N_1238);
and U3101 (N_3101,N_51,N_804);
or U3102 (N_3102,N_1073,N_422);
nor U3103 (N_3103,N_2465,N_523);
nor U3104 (N_3104,N_2479,N_2083);
and U3105 (N_3105,N_1024,N_2385);
nor U3106 (N_3106,N_1658,N_1707);
or U3107 (N_3107,N_1275,N_1192);
or U3108 (N_3108,N_1318,N_2378);
and U3109 (N_3109,N_683,N_4);
nand U3110 (N_3110,N_2072,N_419);
and U3111 (N_3111,N_2380,N_151);
or U3112 (N_3112,N_2044,N_1444);
nor U3113 (N_3113,N_1909,N_430);
and U3114 (N_3114,N_940,N_1779);
nor U3115 (N_3115,N_1953,N_768);
nand U3116 (N_3116,N_1972,N_239);
or U3117 (N_3117,N_882,N_1285);
nand U3118 (N_3118,N_2438,N_2214);
and U3119 (N_3119,N_460,N_121);
or U3120 (N_3120,N_861,N_127);
and U3121 (N_3121,N_2195,N_1609);
nand U3122 (N_3122,N_1524,N_1675);
nor U3123 (N_3123,N_1184,N_561);
and U3124 (N_3124,N_599,N_191);
and U3125 (N_3125,N_180,N_1513);
or U3126 (N_3126,N_584,N_1872);
and U3127 (N_3127,N_2364,N_487);
and U3128 (N_3128,N_209,N_1431);
nor U3129 (N_3129,N_1683,N_468);
nand U3130 (N_3130,N_1141,N_2040);
nor U3131 (N_3131,N_2411,N_1155);
nand U3132 (N_3132,N_659,N_1216);
and U3133 (N_3133,N_1380,N_1404);
nand U3134 (N_3134,N_1554,N_2142);
or U3135 (N_3135,N_2123,N_1076);
nand U3136 (N_3136,N_2360,N_745);
nor U3137 (N_3137,N_1418,N_1880);
nand U3138 (N_3138,N_21,N_1740);
and U3139 (N_3139,N_352,N_888);
nor U3140 (N_3140,N_780,N_1697);
nand U3141 (N_3141,N_920,N_1401);
nor U3142 (N_3142,N_25,N_1778);
nor U3143 (N_3143,N_1212,N_545);
nor U3144 (N_3144,N_100,N_552);
or U3145 (N_3145,N_1756,N_1721);
and U3146 (N_3146,N_665,N_305);
nor U3147 (N_3147,N_1514,N_388);
or U3148 (N_3148,N_44,N_1758);
or U3149 (N_3149,N_1734,N_525);
or U3150 (N_3150,N_1681,N_941);
and U3151 (N_3151,N_1429,N_1280);
nand U3152 (N_3152,N_1399,N_442);
nor U3153 (N_3153,N_1229,N_1031);
nand U3154 (N_3154,N_62,N_2184);
nor U3155 (N_3155,N_1411,N_1733);
and U3156 (N_3156,N_1799,N_413);
nand U3157 (N_3157,N_1709,N_3);
and U3158 (N_3158,N_2011,N_2156);
and U3159 (N_3159,N_1307,N_393);
and U3160 (N_3160,N_2488,N_564);
or U3161 (N_3161,N_2357,N_1583);
and U3162 (N_3162,N_286,N_2490);
and U3163 (N_3163,N_1393,N_2437);
and U3164 (N_3164,N_1060,N_764);
or U3165 (N_3165,N_1263,N_1764);
or U3166 (N_3166,N_1704,N_2125);
or U3167 (N_3167,N_1852,N_319);
and U3168 (N_3168,N_2395,N_2409);
and U3169 (N_3169,N_97,N_1025);
and U3170 (N_3170,N_1002,N_314);
and U3171 (N_3171,N_1265,N_2208);
nand U3172 (N_3172,N_2023,N_2069);
nor U3173 (N_3173,N_2150,N_1368);
and U3174 (N_3174,N_1538,N_1724);
and U3175 (N_3175,N_1384,N_162);
nor U3176 (N_3176,N_154,N_129);
nand U3177 (N_3177,N_293,N_1565);
nor U3178 (N_3178,N_847,N_400);
nand U3179 (N_3179,N_66,N_27);
or U3180 (N_3180,N_15,N_1070);
nor U3181 (N_3181,N_588,N_1426);
nand U3182 (N_3182,N_567,N_404);
nor U3183 (N_3183,N_1732,N_174);
or U3184 (N_3184,N_1936,N_445);
nor U3185 (N_3185,N_1763,N_178);
and U3186 (N_3186,N_1205,N_1022);
and U3187 (N_3187,N_554,N_333);
nand U3188 (N_3188,N_2145,N_1665);
nor U3189 (N_3189,N_1329,N_587);
and U3190 (N_3190,N_250,N_1969);
and U3191 (N_3191,N_2317,N_1645);
or U3192 (N_3192,N_2294,N_2089);
or U3193 (N_3193,N_1533,N_935);
nor U3194 (N_3194,N_951,N_1300);
or U3195 (N_3195,N_2,N_2175);
and U3196 (N_3196,N_533,N_1381);
nor U3197 (N_3197,N_1379,N_1643);
and U3198 (N_3198,N_1559,N_1750);
or U3199 (N_3199,N_857,N_2033);
and U3200 (N_3200,N_1986,N_1788);
and U3201 (N_3201,N_757,N_1661);
nor U3202 (N_3202,N_270,N_983);
nand U3203 (N_3203,N_2299,N_95);
nand U3204 (N_3204,N_810,N_1882);
nand U3205 (N_3205,N_2422,N_1600);
or U3206 (N_3206,N_2470,N_2447);
nand U3207 (N_3207,N_93,N_955);
xor U3208 (N_3208,N_2059,N_593);
or U3209 (N_3209,N_2307,N_1951);
and U3210 (N_3210,N_1541,N_1215);
and U3211 (N_3211,N_150,N_1374);
and U3212 (N_3212,N_125,N_1305);
nand U3213 (N_3213,N_2455,N_1603);
or U3214 (N_3214,N_534,N_1711);
nand U3215 (N_3215,N_2163,N_1000);
nor U3216 (N_3216,N_1816,N_510);
or U3217 (N_3217,N_1507,N_800);
and U3218 (N_3218,N_218,N_1651);
and U3219 (N_3219,N_608,N_956);
or U3220 (N_3220,N_522,N_248);
or U3221 (N_3221,N_1350,N_2382);
or U3222 (N_3222,N_1736,N_1966);
nor U3223 (N_3223,N_1688,N_1014);
or U3224 (N_3224,N_1062,N_1657);
or U3225 (N_3225,N_2390,N_2336);
or U3226 (N_3226,N_1973,N_1446);
xor U3227 (N_3227,N_2041,N_2430);
and U3228 (N_3228,N_1217,N_53);
nand U3229 (N_3229,N_1810,N_2353);
or U3230 (N_3230,N_2324,N_1131);
xor U3231 (N_3231,N_722,N_2339);
nand U3232 (N_3232,N_957,N_243);
and U3233 (N_3233,N_889,N_1869);
or U3234 (N_3234,N_1288,N_828);
nor U3235 (N_3235,N_215,N_2251);
nand U3236 (N_3236,N_623,N_2282);
or U3237 (N_3237,N_1555,N_230);
nor U3238 (N_3238,N_341,N_2280);
or U3239 (N_3239,N_1147,N_2132);
and U3240 (N_3240,N_931,N_41);
nor U3241 (N_3241,N_2080,N_1793);
and U3242 (N_3242,N_253,N_1376);
nor U3243 (N_3243,N_2202,N_1803);
nor U3244 (N_3244,N_703,N_193);
nor U3245 (N_3245,N_2258,N_750);
nor U3246 (N_3246,N_229,N_2289);
or U3247 (N_3247,N_205,N_2031);
and U3248 (N_3248,N_45,N_2434);
nor U3249 (N_3249,N_1944,N_148);
nor U3250 (N_3250,N_1832,N_1156);
nand U3251 (N_3251,N_47,N_1633);
nor U3252 (N_3252,N_1479,N_1921);
and U3253 (N_3253,N_1765,N_979);
nor U3254 (N_3254,N_1592,N_1649);
and U3255 (N_3255,N_337,N_2335);
xor U3256 (N_3256,N_1873,N_2173);
and U3257 (N_3257,N_379,N_1815);
and U3258 (N_3258,N_1001,N_370);
or U3259 (N_3259,N_195,N_149);
and U3260 (N_3260,N_2377,N_667);
nor U3261 (N_3261,N_349,N_2370);
nand U3262 (N_3262,N_499,N_2188);
and U3263 (N_3263,N_579,N_930);
and U3264 (N_3264,N_312,N_484);
or U3265 (N_3265,N_1581,N_1847);
nor U3266 (N_3266,N_425,N_1405);
nand U3267 (N_3267,N_1984,N_1472);
and U3268 (N_3268,N_2427,N_1906);
nor U3269 (N_3269,N_1162,N_2075);
or U3270 (N_3270,N_2318,N_540);
and U3271 (N_3271,N_2149,N_390);
and U3272 (N_3272,N_1476,N_110);
nand U3273 (N_3273,N_2272,N_514);
or U3274 (N_3274,N_217,N_526);
nor U3275 (N_3275,N_2352,N_1860);
nor U3276 (N_3276,N_92,N_232);
nand U3277 (N_3277,N_1877,N_2475);
nor U3278 (N_3278,N_490,N_6);
and U3279 (N_3279,N_1505,N_2349);
or U3280 (N_3280,N_2068,N_2111);
nand U3281 (N_3281,N_695,N_362);
nand U3282 (N_3282,N_1461,N_1158);
and U3283 (N_3283,N_1363,N_515);
and U3284 (N_3284,N_179,N_1956);
or U3285 (N_3285,N_1033,N_1102);
and U3286 (N_3286,N_302,N_1716);
and U3287 (N_3287,N_2129,N_1456);
nor U3288 (N_3288,N_1223,N_1061);
nand U3289 (N_3289,N_666,N_2244);
and U3290 (N_3290,N_260,N_2347);
nor U3291 (N_3291,N_30,N_1239);
nor U3292 (N_3292,N_553,N_1954);
or U3293 (N_3293,N_697,N_907);
nor U3294 (N_3294,N_1606,N_2354);
and U3295 (N_3295,N_1938,N_915);
or U3296 (N_3296,N_2306,N_1386);
nor U3297 (N_3297,N_196,N_83);
or U3298 (N_3298,N_1637,N_1150);
and U3299 (N_3299,N_134,N_1396);
and U3300 (N_3300,N_1769,N_1614);
nand U3301 (N_3301,N_485,N_313);
nand U3302 (N_3302,N_1375,N_713);
or U3303 (N_3303,N_1754,N_1047);
or U3304 (N_3304,N_189,N_353);
and U3305 (N_3305,N_2491,N_1622);
and U3306 (N_3306,N_1295,N_153);
and U3307 (N_3307,N_84,N_679);
and U3308 (N_3308,N_381,N_1080);
and U3309 (N_3309,N_2146,N_70);
or U3310 (N_3310,N_1528,N_2403);
and U3311 (N_3311,N_497,N_330);
and U3312 (N_3312,N_461,N_2274);
nand U3313 (N_3313,N_1744,N_829);
or U3314 (N_3314,N_2169,N_960);
or U3315 (N_3315,N_1905,N_2113);
nor U3316 (N_3316,N_1045,N_516);
and U3317 (N_3317,N_664,N_96);
and U3318 (N_3318,N_1038,N_480);
and U3319 (N_3319,N_1346,N_2496);
nor U3320 (N_3320,N_444,N_399);
nor U3321 (N_3321,N_354,N_1258);
or U3322 (N_3322,N_578,N_170);
and U3323 (N_3323,N_1406,N_220);
nor U3324 (N_3324,N_89,N_1477);
nor U3325 (N_3325,N_645,N_1013);
nand U3326 (N_3326,N_970,N_869);
nand U3327 (N_3327,N_610,N_909);
nand U3328 (N_3328,N_1737,N_1174);
nand U3329 (N_3329,N_1172,N_1177);
nand U3330 (N_3330,N_405,N_1543);
nand U3331 (N_3331,N_19,N_1702);
or U3332 (N_3332,N_682,N_2417);
or U3333 (N_3333,N_802,N_809);
nor U3334 (N_3334,N_1605,N_541);
or U3335 (N_3335,N_509,N_1096);
nor U3336 (N_3336,N_315,N_1527);
nand U3337 (N_3337,N_1270,N_604);
nor U3338 (N_3338,N_285,N_546);
or U3339 (N_3339,N_167,N_594);
or U3340 (N_3340,N_1739,N_2343);
nor U3341 (N_3341,N_1371,N_1099);
or U3342 (N_3342,N_701,N_2064);
nor U3343 (N_3343,N_2063,N_855);
nor U3344 (N_3344,N_1226,N_725);
and U3345 (N_3345,N_899,N_539);
and U3346 (N_3346,N_86,N_583);
nor U3347 (N_3347,N_617,N_528);
nand U3348 (N_3348,N_1126,N_2200);
nand U3349 (N_3349,N_437,N_641);
nor U3350 (N_3350,N_2392,N_2180);
and U3351 (N_3351,N_427,N_1653);
nor U3352 (N_3352,N_2026,N_1382);
xor U3353 (N_3353,N_201,N_1448);
nand U3354 (N_3354,N_901,N_1279);
nor U3355 (N_3355,N_1292,N_865);
or U3356 (N_3356,N_454,N_1046);
nand U3357 (N_3357,N_464,N_1266);
nand U3358 (N_3358,N_963,N_1677);
and U3359 (N_3359,N_60,N_822);
and U3360 (N_3360,N_1134,N_1958);
or U3361 (N_3361,N_182,N_449);
and U3362 (N_3362,N_342,N_384);
or U3363 (N_3363,N_2099,N_1186);
and U3364 (N_3364,N_1604,N_98);
or U3365 (N_3365,N_331,N_1209);
nand U3366 (N_3366,N_1784,N_1330);
nor U3367 (N_3367,N_1032,N_1591);
and U3368 (N_3368,N_1362,N_672);
nor U3369 (N_3369,N_1254,N_571);
nand U3370 (N_3370,N_1161,N_1391);
and U3371 (N_3371,N_2367,N_355);
nor U3372 (N_3372,N_1417,N_348);
xor U3373 (N_3373,N_2232,N_1439);
or U3374 (N_3374,N_1655,N_866);
xor U3375 (N_3375,N_959,N_981);
and U3376 (N_3376,N_2464,N_407);
or U3377 (N_3377,N_1795,N_1289);
or U3378 (N_3378,N_1929,N_294);
nor U3379 (N_3379,N_1994,N_2108);
nor U3380 (N_3380,N_2227,N_1893);
nor U3381 (N_3381,N_1781,N_310);
or U3382 (N_3382,N_1775,N_1673);
nor U3383 (N_3383,N_2406,N_1588);
or U3384 (N_3384,N_2262,N_2290);
nand U3385 (N_3385,N_1474,N_338);
or U3386 (N_3386,N_1611,N_765);
nand U3387 (N_3387,N_2240,N_1735);
nand U3388 (N_3388,N_2008,N_1901);
or U3389 (N_3389,N_2183,N_373);
xor U3390 (N_3390,N_336,N_2386);
nor U3391 (N_3391,N_2177,N_2474);
nand U3392 (N_3392,N_596,N_966);
or U3393 (N_3393,N_265,N_1135);
or U3394 (N_3394,N_2312,N_1159);
nor U3395 (N_3395,N_1962,N_221);
nor U3396 (N_3396,N_284,N_1252);
nand U3397 (N_3397,N_210,N_2358);
nand U3398 (N_3398,N_1123,N_2218);
nor U3399 (N_3399,N_870,N_1577);
or U3400 (N_3400,N_263,N_474);
nand U3401 (N_3401,N_2482,N_630);
or U3402 (N_3402,N_428,N_626);
and U3403 (N_3403,N_1708,N_536);
and U3404 (N_3404,N_2121,N_1357);
and U3405 (N_3405,N_1299,N_1831);
or U3406 (N_3406,N_2049,N_996);
nand U3407 (N_3407,N_1449,N_2193);
nand U3408 (N_3408,N_249,N_2107);
and U3409 (N_3409,N_212,N_864);
nor U3410 (N_3410,N_1928,N_1862);
xnor U3411 (N_3411,N_990,N_1796);
or U3412 (N_3412,N_14,N_368);
nor U3413 (N_3413,N_1415,N_1403);
nand U3414 (N_3414,N_793,N_481);
nand U3415 (N_3415,N_1626,N_1414);
and U3416 (N_3416,N_242,N_1164);
and U3417 (N_3417,N_234,N_2215);
or U3418 (N_3418,N_2176,N_184);
or U3419 (N_3419,N_1317,N_423);
nor U3420 (N_3420,N_1923,N_986);
or U3421 (N_3421,N_326,N_754);
nand U3422 (N_3422,N_1435,N_327);
and U3423 (N_3423,N_1550,N_1964);
nand U3424 (N_3424,N_1072,N_1978);
nor U3425 (N_3425,N_2246,N_2467);
nand U3426 (N_3426,N_928,N_946);
and U3427 (N_3427,N_1963,N_2211);
or U3428 (N_3428,N_772,N_120);
nand U3429 (N_3429,N_1051,N_5);
nor U3430 (N_3430,N_2036,N_1389);
and U3431 (N_3431,N_794,N_506);
or U3432 (N_3432,N_343,N_68);
and U3433 (N_3433,N_2131,N_501);
nand U3434 (N_3434,N_2340,N_137);
nand U3435 (N_3435,N_2186,N_663);
nor U3436 (N_3436,N_159,N_1615);
nand U3437 (N_3437,N_168,N_446);
nand U3438 (N_3438,N_1628,N_43);
or U3439 (N_3439,N_1113,N_1081);
nand U3440 (N_3440,N_1074,N_738);
and U3441 (N_3441,N_2485,N_547);
or U3442 (N_3442,N_439,N_1745);
or U3443 (N_3443,N_1926,N_235);
nand U3444 (N_3444,N_890,N_28);
nor U3445 (N_3445,N_2471,N_2278);
or U3446 (N_3446,N_34,N_2157);
nor U3447 (N_3447,N_775,N_158);
nor U3448 (N_3448,N_301,N_1256);
nor U3449 (N_3449,N_135,N_1042);
nand U3450 (N_3450,N_2197,N_1146);
nand U3451 (N_3451,N_2058,N_1892);
nand U3452 (N_3452,N_1398,N_1976);
and U3453 (N_3453,N_145,N_443);
nor U3454 (N_3454,N_704,N_2116);
nand U3455 (N_3455,N_1153,N_856);
nand U3456 (N_3456,N_1895,N_2138);
nor U3457 (N_3457,N_786,N_716);
nor U3458 (N_3458,N_2079,N_1487);
nor U3459 (N_3459,N_2423,N_1597);
and U3460 (N_3460,N_1915,N_570);
nand U3461 (N_3461,N_1504,N_860);
or U3462 (N_3462,N_2179,N_1427);
nand U3463 (N_3463,N_850,N_1120);
nor U3464 (N_3464,N_1886,N_845);
nor U3465 (N_3465,N_287,N_269);
and U3466 (N_3466,N_1998,N_1599);
nor U3467 (N_3467,N_858,N_283);
or U3468 (N_3468,N_1244,N_2028);
nand U3469 (N_3469,N_2325,N_1991);
nand U3470 (N_3470,N_1029,N_278);
nand U3471 (N_3471,N_1770,N_1361);
or U3472 (N_3472,N_756,N_1623);
nand U3473 (N_3473,N_605,N_507);
or U3474 (N_3474,N_2301,N_1019);
and U3475 (N_3475,N_2432,N_2281);
or U3476 (N_3476,N_958,N_2414);
nand U3477 (N_3477,N_2209,N_1856);
nand U3478 (N_3478,N_603,N_773);
and U3479 (N_3479,N_1485,N_418);
nor U3480 (N_3480,N_1378,N_762);
and U3481 (N_3481,N_268,N_1518);
and U3482 (N_3482,N_1132,N_998);
and U3483 (N_3483,N_421,N_1030);
and U3484 (N_3484,N_1059,N_1101);
and U3485 (N_3485,N_50,N_622);
or U3486 (N_3486,N_1281,N_2327);
nor U3487 (N_3487,N_133,N_1021);
and U3488 (N_3488,N_2196,N_609);
nand U3489 (N_3489,N_1144,N_2334);
and U3490 (N_3490,N_2018,N_2250);
and U3491 (N_3491,N_2237,N_186);
and U3492 (N_3492,N_2105,N_2248);
nand U3493 (N_3493,N_226,N_1531);
nand U3494 (N_3494,N_126,N_2456);
and U3495 (N_3495,N_2124,N_640);
nor U3496 (N_3496,N_1772,N_1253);
nand U3497 (N_3497,N_934,N_1194);
nand U3498 (N_3498,N_1468,N_130);
and U3499 (N_3499,N_1105,N_1660);
nand U3500 (N_3500,N_1537,N_1084);
nor U3501 (N_3501,N_2391,N_1214);
or U3502 (N_3502,N_555,N_465);
and U3503 (N_3503,N_2498,N_673);
nand U3504 (N_3504,N_1210,N_1303);
and U3505 (N_3505,N_1679,N_937);
nor U3506 (N_3506,N_274,N_2344);
or U3507 (N_3507,N_2270,N_1163);
and U3508 (N_3508,N_176,N_742);
nor U3509 (N_3509,N_752,N_103);
or U3510 (N_3510,N_573,N_743);
nand U3511 (N_3511,N_2172,N_1373);
nor U3512 (N_3512,N_1943,N_1636);
and U3513 (N_3513,N_1571,N_1981);
or U3514 (N_3514,N_2293,N_1466);
nor U3515 (N_3515,N_1942,N_513);
or U3516 (N_3516,N_1590,N_2144);
or U3517 (N_3517,N_1287,N_2231);
nand U3518 (N_3518,N_2431,N_527);
nand U3519 (N_3519,N_1430,N_519);
or U3520 (N_3520,N_106,N_1663);
nand U3521 (N_3521,N_1575,N_1165);
or U3522 (N_3522,N_207,N_1974);
nand U3523 (N_3523,N_1792,N_576);
or U3524 (N_3524,N_1027,N_837);
nor U3525 (N_3525,N_620,N_1331);
nor U3526 (N_3526,N_681,N_2207);
and U3527 (N_3527,N_1,N_1413);
or U3528 (N_3528,N_458,N_2444);
or U3529 (N_3529,N_670,N_875);
or U3530 (N_3530,N_2065,N_2229);
nand U3531 (N_3531,N_1438,N_841);
or U3532 (N_3532,N_244,N_1441);
nand U3533 (N_3533,N_862,N_1143);
or U3534 (N_3534,N_2295,N_104);
and U3535 (N_3535,N_1569,N_1858);
or U3536 (N_3536,N_2155,N_2106);
and U3537 (N_3537,N_2141,N_1420);
or U3538 (N_3538,N_1608,N_1459);
and U3539 (N_3539,N_451,N_2095);
nand U3540 (N_3540,N_276,N_2287);
or U3541 (N_3541,N_1306,N_1237);
or U3542 (N_3542,N_1402,N_1825);
and U3543 (N_3543,N_1284,N_1206);
and U3544 (N_3544,N_227,N_688);
nand U3545 (N_3545,N_611,N_1552);
or U3546 (N_3546,N_1005,N_1308);
nand U3547 (N_3547,N_463,N_1152);
or U3548 (N_3548,N_1114,N_1907);
nor U3549 (N_3549,N_396,N_1071);
nor U3550 (N_3550,N_2396,N_2162);
or U3551 (N_3551,N_871,N_99);
or U3552 (N_3552,N_677,N_1865);
nor U3553 (N_3553,N_251,N_1589);
and U3554 (N_3554,N_2407,N_299);
and U3555 (N_3555,N_643,N_1689);
nand U3556 (N_3556,N_2056,N_12);
or U3557 (N_3557,N_1761,N_1568);
nand U3558 (N_3558,N_91,N_1063);
and U3559 (N_3559,N_639,N_1814);
nand U3560 (N_3560,N_1260,N_2055);
or U3561 (N_3561,N_1098,N_1672);
or U3562 (N_3562,N_2468,N_2006);
nand U3563 (N_3563,N_2384,N_1198);
nand U3564 (N_3564,N_1283,N_1480);
and U3565 (N_3565,N_1372,N_1753);
or U3566 (N_3566,N_1891,N_80);
nor U3567 (N_3567,N_1621,N_2252);
nand U3568 (N_3568,N_0,N_932);
or U3569 (N_3569,N_52,N_1596);
or U3570 (N_3570,N_271,N_1269);
nand U3571 (N_3571,N_1601,N_658);
or U3572 (N_3572,N_633,N_1296);
or U3573 (N_3573,N_918,N_790);
nor U3574 (N_3574,N_1797,N_1777);
and U3575 (N_3575,N_2001,N_1811);
nand U3576 (N_3576,N_1952,N_1130);
or U3577 (N_3577,N_39,N_1433);
nand U3578 (N_3578,N_897,N_2194);
or U3579 (N_3579,N_503,N_101);
and U3580 (N_3580,N_36,N_1007);
nand U3581 (N_3581,N_288,N_1512);
nor U3582 (N_3582,N_247,N_1197);
or U3583 (N_3583,N_367,N_687);
and U3584 (N_3584,N_211,N_1323);
or U3585 (N_3585,N_1564,N_2236);
nand U3586 (N_3586,N_1975,N_1935);
and U3587 (N_3587,N_392,N_1267);
nand U3588 (N_3588,N_1110,N_2256);
nor U3589 (N_3589,N_1602,N_450);
or U3590 (N_3590,N_1383,N_1094);
or U3591 (N_3591,N_2291,N_685);
and U3592 (N_3592,N_1471,N_1127);
or U3593 (N_3593,N_1834,N_1666);
nor U3594 (N_3594,N_655,N_496);
nor U3595 (N_3595,N_719,N_383);
or U3596 (N_3596,N_1961,N_1684);
nand U3597 (N_3597,N_1054,N_1298);
or U3598 (N_3598,N_1616,N_46);
or U3599 (N_3599,N_2389,N_634);
nor U3600 (N_3600,N_2014,N_2181);
nor U3601 (N_3601,N_661,N_2329);
and U3602 (N_3602,N_524,N_1199);
and U3603 (N_3603,N_1491,N_2413);
and U3604 (N_3604,N_1997,N_628);
nor U3605 (N_3605,N_2201,N_111);
nor U3606 (N_3606,N_1647,N_2226);
or U3607 (N_3607,N_1064,N_316);
or U3608 (N_3608,N_1481,N_306);
and U3609 (N_3609,N_1322,N_1228);
and U3610 (N_3610,N_1090,N_1268);
nand U3611 (N_3611,N_2415,N_668);
nand U3612 (N_3612,N_241,N_2451);
nor U3613 (N_3613,N_1806,N_2452);
and U3614 (N_3614,N_619,N_116);
and U3615 (N_3615,N_2153,N_544);
nand U3616 (N_3616,N_2276,N_1839);
nand U3617 (N_3617,N_1246,N_805);
nand U3618 (N_3618,N_1203,N_1783);
nor U3619 (N_3619,N_1489,N_1245);
nand U3620 (N_3620,N_2435,N_1617);
nand U3621 (N_3621,N_1558,N_1812);
nand U3622 (N_3622,N_1234,N_2495);
nand U3623 (N_3623,N_1176,N_2233);
nor U3624 (N_3624,N_1040,N_1851);
nand U3625 (N_3625,N_1053,N_991);
nand U3626 (N_3626,N_1980,N_478);
nand U3627 (N_3627,N_2499,N_190);
nor U3628 (N_3628,N_650,N_1342);
or U3629 (N_3629,N_933,N_2086);
or U3630 (N_3630,N_261,N_1142);
nand U3631 (N_3631,N_1495,N_374);
and U3632 (N_3632,N_2259,N_1748);
nand U3633 (N_3633,N_2127,N_85);
nand U3634 (N_3634,N_813,N_1650);
or U3635 (N_3635,N_898,N_993);
or U3636 (N_3636,N_2205,N_1075);
nand U3637 (N_3637,N_495,N_712);
nor U3638 (N_3638,N_779,N_651);
and U3639 (N_3639,N_2310,N_206);
and U3640 (N_3640,N_2057,N_1968);
nand U3641 (N_3641,N_334,N_660);
and U3642 (N_3642,N_548,N_2154);
and U3643 (N_3643,N_1561,N_843);
nand U3644 (N_3644,N_1545,N_1876);
nand U3645 (N_3645,N_2091,N_1041);
and U3646 (N_3646,N_74,N_2004);
nor U3647 (N_3647,N_1529,N_580);
nor U3648 (N_3648,N_873,N_356);
nor U3649 (N_3649,N_558,N_973);
nor U3650 (N_3650,N_377,N_157);
and U3651 (N_3651,N_1530,N_1743);
or U3652 (N_3652,N_844,N_751);
or U3653 (N_3653,N_216,N_1364);
and U3654 (N_3654,N_141,N_1207);
or U3655 (N_3655,N_2071,N_1109);
or U3656 (N_3656,N_1314,N_1828);
nor U3657 (N_3657,N_2245,N_2228);
and U3658 (N_3658,N_989,N_657);
nor U3659 (N_3659,N_2381,N_2337);
nor U3660 (N_3660,N_2035,N_1107);
nor U3661 (N_3661,N_358,N_1236);
nand U3662 (N_3662,N_950,N_815);
and U3663 (N_3663,N_457,N_335);
or U3664 (N_3664,N_1202,N_1925);
nand U3665 (N_3665,N_2060,N_550);
and U3666 (N_3666,N_1241,N_1325);
nand U3667 (N_3667,N_1613,N_1097);
nor U3668 (N_3668,N_939,N_475);
nor U3669 (N_3669,N_17,N_88);
and U3670 (N_3670,N_1388,N_1534);
and U3671 (N_3671,N_1959,N_531);
and U3672 (N_3672,N_2366,N_2120);
nand U3673 (N_3673,N_395,N_2489);
and U3674 (N_3674,N_1520,N_727);
nand U3675 (N_3675,N_761,N_569);
or U3676 (N_3676,N_359,N_1720);
or U3677 (N_3677,N_1067,N_1536);
nor U3678 (N_3678,N_2426,N_848);
and U3679 (N_3679,N_1093,N_1855);
or U3680 (N_3680,N_2355,N_1913);
and U3681 (N_3681,N_258,N_2171);
and U3682 (N_3682,N_375,N_631);
and U3683 (N_3683,N_854,N_833);
nand U3684 (N_3684,N_2029,N_1366);
and U3685 (N_3685,N_2027,N_1017);
or U3686 (N_3686,N_774,N_2220);
nor U3687 (N_3687,N_282,N_2066);
or U3688 (N_3688,N_1639,N_2013);
nand U3689 (N_3689,N_79,N_2302);
or U3690 (N_3690,N_1945,N_2178);
nor U3691 (N_3691,N_1835,N_820);
nor U3692 (N_3692,N_838,N_2009);
and U3693 (N_3693,N_483,N_886);
nand U3694 (N_3694,N_1786,N_1069);
nand U3695 (N_3695,N_1519,N_880);
and U3696 (N_3696,N_160,N_9);
nor U3697 (N_3697,N_2308,N_1315);
nor U3698 (N_3698,N_532,N_2158);
or U3699 (N_3699,N_962,N_2078);
nand U3700 (N_3700,N_1813,N_732);
and U3701 (N_3701,N_758,N_1328);
and U3702 (N_3702,N_1294,N_1039);
and U3703 (N_3703,N_2393,N_1170);
nor U3704 (N_3704,N_1562,N_884);
nand U3705 (N_3705,N_194,N_13);
xor U3706 (N_3706,N_494,N_394);
nor U3707 (N_3707,N_755,N_1160);
or U3708 (N_3708,N_1567,N_2373);
or U3709 (N_3709,N_906,N_1335);
nor U3710 (N_3710,N_2449,N_403);
nor U3711 (N_3711,N_2249,N_2387);
or U3712 (N_3712,N_1111,N_699);
nor U3713 (N_3713,N_2319,N_1823);
xnor U3714 (N_3714,N_2038,N_1691);
nand U3715 (N_3715,N_1183,N_1826);
and U3716 (N_3716,N_795,N_1095);
and U3717 (N_3717,N_1887,N_2483);
or U3718 (N_3718,N_1932,N_1400);
or U3719 (N_3719,N_81,N_2472);
nor U3720 (N_3720,N_476,N_2433);
or U3721 (N_3721,N_597,N_911);
or U3722 (N_3722,N_535,N_361);
nor U3723 (N_3723,N_2255,N_563);
and U3724 (N_3724,N_1208,N_2345);
or U3725 (N_3725,N_1523,N_2076);
and U3726 (N_3726,N_2084,N_646);
nand U3727 (N_3727,N_1947,N_1048);
nand U3728 (N_3728,N_1394,N_649);
nand U3729 (N_3729,N_322,N_1145);
and U3730 (N_3730,N_1104,N_371);
nand U3731 (N_3731,N_537,N_1829);
or U3732 (N_3732,N_118,N_1004);
nand U3733 (N_3733,N_2165,N_551);
and U3734 (N_3734,N_364,N_891);
or U3735 (N_3735,N_1671,N_1297);
or U3736 (N_3736,N_1619,N_1844);
or U3737 (N_3737,N_414,N_2097);
or U3738 (N_3738,N_852,N_366);
or U3739 (N_3739,N_2247,N_816);
and U3740 (N_3740,N_543,N_614);
nand U3741 (N_3741,N_895,N_1848);
or U3742 (N_3742,N_58,N_505);
and U3743 (N_3743,N_808,N_832);
nor U3744 (N_3744,N_1467,N_2230);
and U3745 (N_3745,N_529,N_1419);
or U3746 (N_3746,N_502,N_724);
nand U3747 (N_3747,N_1432,N_1088);
nand U3748 (N_3748,N_2133,N_968);
nor U3749 (N_3749,N_1693,N_1496);
nor U3750 (N_3750,N_2247,N_1235);
nor U3751 (N_3751,N_195,N_1807);
or U3752 (N_3752,N_1780,N_1099);
and U3753 (N_3753,N_1338,N_1436);
nand U3754 (N_3754,N_172,N_2432);
nor U3755 (N_3755,N_2233,N_652);
nor U3756 (N_3756,N_229,N_2442);
nand U3757 (N_3757,N_1200,N_2236);
and U3758 (N_3758,N_1015,N_2230);
nand U3759 (N_3759,N_1041,N_1663);
or U3760 (N_3760,N_1410,N_1015);
nor U3761 (N_3761,N_2249,N_2401);
or U3762 (N_3762,N_2086,N_1654);
nand U3763 (N_3763,N_267,N_1564);
nor U3764 (N_3764,N_99,N_2122);
or U3765 (N_3765,N_89,N_53);
and U3766 (N_3766,N_396,N_115);
nor U3767 (N_3767,N_388,N_1173);
nand U3768 (N_3768,N_1411,N_559);
nor U3769 (N_3769,N_1094,N_90);
nand U3770 (N_3770,N_37,N_807);
and U3771 (N_3771,N_309,N_408);
or U3772 (N_3772,N_670,N_2189);
nand U3773 (N_3773,N_1345,N_1632);
nand U3774 (N_3774,N_2382,N_2370);
or U3775 (N_3775,N_1016,N_2276);
or U3776 (N_3776,N_1679,N_2110);
nand U3777 (N_3777,N_617,N_899);
and U3778 (N_3778,N_18,N_2134);
nor U3779 (N_3779,N_2079,N_595);
or U3780 (N_3780,N_1041,N_2128);
or U3781 (N_3781,N_1062,N_1468);
nor U3782 (N_3782,N_2037,N_503);
or U3783 (N_3783,N_2106,N_1531);
or U3784 (N_3784,N_1628,N_787);
nand U3785 (N_3785,N_1307,N_1937);
and U3786 (N_3786,N_897,N_1928);
nand U3787 (N_3787,N_265,N_703);
nand U3788 (N_3788,N_1653,N_631);
nor U3789 (N_3789,N_857,N_1759);
nand U3790 (N_3790,N_2,N_2137);
and U3791 (N_3791,N_455,N_319);
and U3792 (N_3792,N_1314,N_1298);
nor U3793 (N_3793,N_2436,N_1923);
and U3794 (N_3794,N_1984,N_2130);
nor U3795 (N_3795,N_376,N_116);
or U3796 (N_3796,N_771,N_2494);
nor U3797 (N_3797,N_1134,N_698);
nor U3798 (N_3798,N_1966,N_730);
or U3799 (N_3799,N_2398,N_1497);
or U3800 (N_3800,N_2447,N_1490);
and U3801 (N_3801,N_1244,N_1224);
and U3802 (N_3802,N_1712,N_74);
nor U3803 (N_3803,N_1835,N_2477);
nand U3804 (N_3804,N_906,N_195);
and U3805 (N_3805,N_233,N_2457);
and U3806 (N_3806,N_2180,N_1116);
and U3807 (N_3807,N_2326,N_2115);
or U3808 (N_3808,N_705,N_2412);
or U3809 (N_3809,N_1474,N_1299);
nand U3810 (N_3810,N_190,N_2414);
nand U3811 (N_3811,N_1035,N_209);
or U3812 (N_3812,N_2314,N_1093);
or U3813 (N_3813,N_2028,N_1776);
and U3814 (N_3814,N_2011,N_25);
or U3815 (N_3815,N_2481,N_1127);
or U3816 (N_3816,N_969,N_1006);
nand U3817 (N_3817,N_524,N_1684);
and U3818 (N_3818,N_2349,N_211);
nand U3819 (N_3819,N_755,N_1014);
and U3820 (N_3820,N_623,N_1111);
or U3821 (N_3821,N_2483,N_30);
nor U3822 (N_3822,N_777,N_2302);
and U3823 (N_3823,N_1123,N_88);
nor U3824 (N_3824,N_1485,N_813);
nor U3825 (N_3825,N_1040,N_2496);
or U3826 (N_3826,N_1173,N_1648);
or U3827 (N_3827,N_68,N_119);
and U3828 (N_3828,N_435,N_79);
nand U3829 (N_3829,N_2279,N_530);
nand U3830 (N_3830,N_306,N_568);
and U3831 (N_3831,N_1713,N_1774);
nor U3832 (N_3832,N_1631,N_1106);
and U3833 (N_3833,N_687,N_648);
and U3834 (N_3834,N_1805,N_380);
nand U3835 (N_3835,N_1610,N_1779);
and U3836 (N_3836,N_1838,N_1768);
nand U3837 (N_3837,N_669,N_495);
and U3838 (N_3838,N_1217,N_684);
nand U3839 (N_3839,N_715,N_560);
nand U3840 (N_3840,N_958,N_1998);
nor U3841 (N_3841,N_64,N_1198);
or U3842 (N_3842,N_442,N_981);
nor U3843 (N_3843,N_10,N_142);
and U3844 (N_3844,N_1003,N_580);
nand U3845 (N_3845,N_175,N_580);
or U3846 (N_3846,N_1314,N_596);
nor U3847 (N_3847,N_1800,N_588);
or U3848 (N_3848,N_1527,N_755);
nor U3849 (N_3849,N_581,N_395);
and U3850 (N_3850,N_2206,N_99);
and U3851 (N_3851,N_1847,N_1460);
nor U3852 (N_3852,N_1524,N_1853);
or U3853 (N_3853,N_1108,N_1144);
and U3854 (N_3854,N_1650,N_286);
nand U3855 (N_3855,N_1288,N_1969);
or U3856 (N_3856,N_501,N_608);
or U3857 (N_3857,N_616,N_224);
nand U3858 (N_3858,N_1914,N_1339);
nand U3859 (N_3859,N_1113,N_698);
nand U3860 (N_3860,N_1552,N_2423);
or U3861 (N_3861,N_1134,N_1178);
or U3862 (N_3862,N_679,N_2341);
or U3863 (N_3863,N_1590,N_1214);
and U3864 (N_3864,N_1386,N_10);
nor U3865 (N_3865,N_471,N_1927);
or U3866 (N_3866,N_766,N_2047);
nor U3867 (N_3867,N_471,N_2162);
nand U3868 (N_3868,N_2317,N_1434);
and U3869 (N_3869,N_2430,N_1639);
nand U3870 (N_3870,N_1028,N_830);
and U3871 (N_3871,N_2403,N_1436);
nand U3872 (N_3872,N_2311,N_2318);
nand U3873 (N_3873,N_1366,N_2372);
nand U3874 (N_3874,N_1683,N_1977);
and U3875 (N_3875,N_1404,N_509);
nand U3876 (N_3876,N_1085,N_1789);
nor U3877 (N_3877,N_204,N_782);
nand U3878 (N_3878,N_186,N_2031);
or U3879 (N_3879,N_1553,N_1152);
nand U3880 (N_3880,N_2096,N_424);
nor U3881 (N_3881,N_2279,N_609);
or U3882 (N_3882,N_1795,N_188);
or U3883 (N_3883,N_2242,N_1591);
and U3884 (N_3884,N_2197,N_1034);
nor U3885 (N_3885,N_1322,N_205);
or U3886 (N_3886,N_323,N_450);
or U3887 (N_3887,N_868,N_1208);
or U3888 (N_3888,N_647,N_1916);
nor U3889 (N_3889,N_2091,N_1674);
and U3890 (N_3890,N_1612,N_954);
nand U3891 (N_3891,N_1414,N_1316);
or U3892 (N_3892,N_1415,N_1486);
nor U3893 (N_3893,N_201,N_2004);
or U3894 (N_3894,N_1392,N_528);
or U3895 (N_3895,N_1845,N_2377);
or U3896 (N_3896,N_1124,N_1148);
nor U3897 (N_3897,N_2064,N_1787);
and U3898 (N_3898,N_420,N_993);
and U3899 (N_3899,N_1456,N_186);
nor U3900 (N_3900,N_511,N_1596);
and U3901 (N_3901,N_2206,N_1747);
and U3902 (N_3902,N_2203,N_1906);
nor U3903 (N_3903,N_1961,N_393);
nand U3904 (N_3904,N_151,N_2312);
and U3905 (N_3905,N_2306,N_1853);
and U3906 (N_3906,N_15,N_994);
nor U3907 (N_3907,N_2034,N_378);
and U3908 (N_3908,N_1209,N_342);
nor U3909 (N_3909,N_1925,N_1159);
nor U3910 (N_3910,N_267,N_231);
and U3911 (N_3911,N_319,N_1745);
and U3912 (N_3912,N_411,N_2157);
nor U3913 (N_3913,N_467,N_1922);
or U3914 (N_3914,N_2186,N_1405);
nor U3915 (N_3915,N_2021,N_1427);
and U3916 (N_3916,N_802,N_1277);
nand U3917 (N_3917,N_194,N_2149);
or U3918 (N_3918,N_123,N_1892);
and U3919 (N_3919,N_675,N_1508);
and U3920 (N_3920,N_1662,N_1210);
or U3921 (N_3921,N_1926,N_2096);
or U3922 (N_3922,N_149,N_2307);
or U3923 (N_3923,N_919,N_310);
or U3924 (N_3924,N_878,N_1312);
and U3925 (N_3925,N_1359,N_1775);
and U3926 (N_3926,N_644,N_180);
or U3927 (N_3927,N_1988,N_858);
nor U3928 (N_3928,N_1501,N_1685);
or U3929 (N_3929,N_570,N_395);
nand U3930 (N_3930,N_1890,N_1509);
or U3931 (N_3931,N_611,N_293);
nor U3932 (N_3932,N_134,N_1974);
or U3933 (N_3933,N_859,N_2340);
and U3934 (N_3934,N_1953,N_1823);
nor U3935 (N_3935,N_853,N_1836);
nor U3936 (N_3936,N_1266,N_1131);
nand U3937 (N_3937,N_10,N_1047);
or U3938 (N_3938,N_646,N_878);
nand U3939 (N_3939,N_1405,N_680);
nor U3940 (N_3940,N_1509,N_1636);
nor U3941 (N_3941,N_1017,N_926);
or U3942 (N_3942,N_308,N_164);
nor U3943 (N_3943,N_1142,N_1084);
and U3944 (N_3944,N_542,N_1575);
nand U3945 (N_3945,N_1888,N_194);
or U3946 (N_3946,N_141,N_1280);
nor U3947 (N_3947,N_218,N_941);
nor U3948 (N_3948,N_541,N_608);
nor U3949 (N_3949,N_557,N_894);
and U3950 (N_3950,N_1740,N_1475);
and U3951 (N_3951,N_849,N_221);
nor U3952 (N_3952,N_1500,N_1087);
nor U3953 (N_3953,N_1869,N_2346);
nand U3954 (N_3954,N_1621,N_1213);
nor U3955 (N_3955,N_925,N_1947);
and U3956 (N_3956,N_854,N_2045);
nor U3957 (N_3957,N_2163,N_525);
nor U3958 (N_3958,N_2213,N_74);
and U3959 (N_3959,N_1282,N_838);
or U3960 (N_3960,N_674,N_122);
and U3961 (N_3961,N_197,N_1939);
and U3962 (N_3962,N_1824,N_1185);
and U3963 (N_3963,N_389,N_1949);
and U3964 (N_3964,N_1510,N_871);
and U3965 (N_3965,N_1036,N_2266);
xor U3966 (N_3966,N_517,N_39);
nand U3967 (N_3967,N_461,N_635);
or U3968 (N_3968,N_1174,N_2465);
or U3969 (N_3969,N_1482,N_898);
nand U3970 (N_3970,N_355,N_1585);
and U3971 (N_3971,N_1433,N_1652);
or U3972 (N_3972,N_992,N_2364);
nor U3973 (N_3973,N_1880,N_1007);
nor U3974 (N_3974,N_1688,N_1109);
nand U3975 (N_3975,N_2400,N_1169);
nor U3976 (N_3976,N_1137,N_790);
or U3977 (N_3977,N_794,N_1556);
nand U3978 (N_3978,N_1383,N_1423);
nand U3979 (N_3979,N_83,N_121);
nand U3980 (N_3980,N_2204,N_1481);
xor U3981 (N_3981,N_170,N_435);
and U3982 (N_3982,N_412,N_769);
nand U3983 (N_3983,N_1234,N_1405);
nor U3984 (N_3984,N_2450,N_1254);
or U3985 (N_3985,N_452,N_1525);
and U3986 (N_3986,N_2260,N_161);
nor U3987 (N_3987,N_1068,N_1722);
nand U3988 (N_3988,N_1420,N_1814);
nand U3989 (N_3989,N_1430,N_297);
nand U3990 (N_3990,N_132,N_990);
nor U3991 (N_3991,N_2377,N_1864);
or U3992 (N_3992,N_2266,N_2449);
nor U3993 (N_3993,N_540,N_1486);
and U3994 (N_3994,N_1873,N_1770);
nor U3995 (N_3995,N_2295,N_1841);
and U3996 (N_3996,N_3,N_1570);
nor U3997 (N_3997,N_1337,N_1890);
nand U3998 (N_3998,N_5,N_2135);
nor U3999 (N_3999,N_1024,N_1725);
nor U4000 (N_4000,N_787,N_649);
and U4001 (N_4001,N_835,N_2032);
nand U4002 (N_4002,N_1265,N_411);
nand U4003 (N_4003,N_1959,N_453);
and U4004 (N_4004,N_1063,N_1416);
nand U4005 (N_4005,N_127,N_64);
nand U4006 (N_4006,N_971,N_1679);
nand U4007 (N_4007,N_2168,N_106);
or U4008 (N_4008,N_2418,N_1543);
nor U4009 (N_4009,N_2394,N_1247);
nand U4010 (N_4010,N_1844,N_1157);
and U4011 (N_4011,N_1141,N_2388);
and U4012 (N_4012,N_600,N_1849);
or U4013 (N_4013,N_266,N_17);
nand U4014 (N_4014,N_1517,N_270);
nand U4015 (N_4015,N_1199,N_553);
nand U4016 (N_4016,N_2037,N_122);
nor U4017 (N_4017,N_867,N_1612);
nand U4018 (N_4018,N_647,N_2421);
or U4019 (N_4019,N_1514,N_2197);
and U4020 (N_4020,N_2211,N_212);
nor U4021 (N_4021,N_1935,N_2041);
or U4022 (N_4022,N_1756,N_969);
or U4023 (N_4023,N_1735,N_2266);
and U4024 (N_4024,N_1169,N_566);
nand U4025 (N_4025,N_549,N_1109);
or U4026 (N_4026,N_1354,N_2497);
nor U4027 (N_4027,N_1413,N_764);
or U4028 (N_4028,N_671,N_213);
or U4029 (N_4029,N_2296,N_323);
nor U4030 (N_4030,N_13,N_39);
or U4031 (N_4031,N_2173,N_1069);
and U4032 (N_4032,N_1072,N_1539);
and U4033 (N_4033,N_2059,N_179);
nand U4034 (N_4034,N_1987,N_1398);
nand U4035 (N_4035,N_1286,N_1746);
nor U4036 (N_4036,N_1096,N_1868);
nand U4037 (N_4037,N_682,N_2296);
or U4038 (N_4038,N_2417,N_634);
or U4039 (N_4039,N_1016,N_2079);
or U4040 (N_4040,N_937,N_514);
or U4041 (N_4041,N_1717,N_1996);
and U4042 (N_4042,N_2046,N_2385);
or U4043 (N_4043,N_1655,N_1199);
and U4044 (N_4044,N_2250,N_574);
and U4045 (N_4045,N_1426,N_1904);
nand U4046 (N_4046,N_626,N_97);
nor U4047 (N_4047,N_1907,N_2457);
or U4048 (N_4048,N_1948,N_1258);
nor U4049 (N_4049,N_244,N_2170);
nand U4050 (N_4050,N_1710,N_1207);
nor U4051 (N_4051,N_847,N_288);
nand U4052 (N_4052,N_1228,N_672);
or U4053 (N_4053,N_1579,N_193);
or U4054 (N_4054,N_1989,N_2294);
nor U4055 (N_4055,N_456,N_1569);
or U4056 (N_4056,N_646,N_1650);
or U4057 (N_4057,N_1904,N_298);
nor U4058 (N_4058,N_2369,N_2436);
and U4059 (N_4059,N_522,N_481);
nand U4060 (N_4060,N_2441,N_251);
nor U4061 (N_4061,N_574,N_617);
nand U4062 (N_4062,N_2226,N_604);
nand U4063 (N_4063,N_111,N_589);
or U4064 (N_4064,N_1179,N_933);
nand U4065 (N_4065,N_1079,N_707);
or U4066 (N_4066,N_2400,N_1843);
and U4067 (N_4067,N_1079,N_1338);
or U4068 (N_4068,N_656,N_1463);
and U4069 (N_4069,N_2210,N_1115);
or U4070 (N_4070,N_1522,N_1866);
nor U4071 (N_4071,N_1820,N_210);
and U4072 (N_4072,N_1234,N_620);
nor U4073 (N_4073,N_1179,N_1967);
nor U4074 (N_4074,N_2488,N_15);
or U4075 (N_4075,N_730,N_1332);
nand U4076 (N_4076,N_1588,N_632);
and U4077 (N_4077,N_1609,N_1068);
nand U4078 (N_4078,N_2072,N_2364);
nand U4079 (N_4079,N_324,N_2309);
and U4080 (N_4080,N_1616,N_220);
nor U4081 (N_4081,N_1600,N_643);
nand U4082 (N_4082,N_1557,N_2049);
or U4083 (N_4083,N_713,N_102);
and U4084 (N_4084,N_432,N_1492);
and U4085 (N_4085,N_426,N_1193);
nand U4086 (N_4086,N_254,N_1120);
and U4087 (N_4087,N_2100,N_1587);
nor U4088 (N_4088,N_11,N_847);
and U4089 (N_4089,N_1804,N_2297);
nand U4090 (N_4090,N_770,N_331);
and U4091 (N_4091,N_1577,N_1987);
nor U4092 (N_4092,N_2127,N_1117);
nand U4093 (N_4093,N_163,N_1902);
nor U4094 (N_4094,N_1539,N_974);
and U4095 (N_4095,N_2124,N_1156);
and U4096 (N_4096,N_285,N_1595);
or U4097 (N_4097,N_817,N_692);
and U4098 (N_4098,N_133,N_631);
or U4099 (N_4099,N_114,N_2359);
or U4100 (N_4100,N_2040,N_2109);
nor U4101 (N_4101,N_1086,N_136);
nor U4102 (N_4102,N_458,N_1480);
nand U4103 (N_4103,N_168,N_2323);
nand U4104 (N_4104,N_777,N_1617);
or U4105 (N_4105,N_202,N_2450);
nand U4106 (N_4106,N_1985,N_538);
nor U4107 (N_4107,N_994,N_628);
nand U4108 (N_4108,N_2197,N_905);
or U4109 (N_4109,N_1015,N_1141);
nor U4110 (N_4110,N_1197,N_377);
nor U4111 (N_4111,N_1170,N_1285);
nand U4112 (N_4112,N_1711,N_1705);
nand U4113 (N_4113,N_1937,N_1121);
or U4114 (N_4114,N_530,N_1473);
nand U4115 (N_4115,N_1185,N_1218);
nor U4116 (N_4116,N_2285,N_666);
nor U4117 (N_4117,N_1121,N_1977);
nor U4118 (N_4118,N_293,N_1502);
and U4119 (N_4119,N_2129,N_599);
xor U4120 (N_4120,N_2291,N_97);
or U4121 (N_4121,N_2354,N_1080);
and U4122 (N_4122,N_1635,N_1844);
and U4123 (N_4123,N_64,N_2292);
nor U4124 (N_4124,N_1706,N_1278);
or U4125 (N_4125,N_1326,N_1403);
nor U4126 (N_4126,N_2372,N_2497);
or U4127 (N_4127,N_1888,N_2159);
and U4128 (N_4128,N_2003,N_234);
nor U4129 (N_4129,N_1271,N_2467);
and U4130 (N_4130,N_1419,N_775);
or U4131 (N_4131,N_1180,N_2046);
and U4132 (N_4132,N_1283,N_977);
or U4133 (N_4133,N_1369,N_296);
and U4134 (N_4134,N_8,N_1945);
nand U4135 (N_4135,N_2271,N_61);
nor U4136 (N_4136,N_875,N_2496);
nand U4137 (N_4137,N_2151,N_2237);
or U4138 (N_4138,N_715,N_1020);
nor U4139 (N_4139,N_274,N_1975);
nand U4140 (N_4140,N_606,N_1361);
or U4141 (N_4141,N_1535,N_1779);
nor U4142 (N_4142,N_118,N_1298);
nor U4143 (N_4143,N_790,N_979);
and U4144 (N_4144,N_1089,N_725);
nor U4145 (N_4145,N_204,N_1756);
nand U4146 (N_4146,N_1579,N_373);
xor U4147 (N_4147,N_1066,N_1976);
or U4148 (N_4148,N_2459,N_1286);
and U4149 (N_4149,N_1111,N_2452);
or U4150 (N_4150,N_1890,N_2130);
or U4151 (N_4151,N_2076,N_2231);
nand U4152 (N_4152,N_2213,N_314);
nor U4153 (N_4153,N_1009,N_2219);
or U4154 (N_4154,N_677,N_312);
or U4155 (N_4155,N_2218,N_81);
and U4156 (N_4156,N_2102,N_412);
or U4157 (N_4157,N_1641,N_2258);
xnor U4158 (N_4158,N_639,N_850);
or U4159 (N_4159,N_273,N_411);
xnor U4160 (N_4160,N_560,N_2063);
and U4161 (N_4161,N_1144,N_1790);
or U4162 (N_4162,N_1395,N_2311);
or U4163 (N_4163,N_2111,N_1665);
and U4164 (N_4164,N_680,N_2489);
or U4165 (N_4165,N_791,N_1800);
nor U4166 (N_4166,N_2130,N_1180);
nand U4167 (N_4167,N_844,N_104);
nand U4168 (N_4168,N_2201,N_2485);
or U4169 (N_4169,N_685,N_2110);
nand U4170 (N_4170,N_1870,N_810);
and U4171 (N_4171,N_1900,N_1512);
nor U4172 (N_4172,N_9,N_2102);
nand U4173 (N_4173,N_2490,N_688);
nand U4174 (N_4174,N_386,N_1228);
nor U4175 (N_4175,N_818,N_1864);
and U4176 (N_4176,N_1103,N_2366);
nor U4177 (N_4177,N_818,N_1729);
and U4178 (N_4178,N_1178,N_1905);
or U4179 (N_4179,N_328,N_2242);
or U4180 (N_4180,N_1421,N_2442);
or U4181 (N_4181,N_1208,N_906);
nand U4182 (N_4182,N_2244,N_694);
and U4183 (N_4183,N_728,N_1135);
nand U4184 (N_4184,N_575,N_258);
nand U4185 (N_4185,N_2151,N_1231);
and U4186 (N_4186,N_451,N_1096);
or U4187 (N_4187,N_1302,N_1082);
or U4188 (N_4188,N_1541,N_2414);
nand U4189 (N_4189,N_2248,N_849);
and U4190 (N_4190,N_1668,N_673);
nor U4191 (N_4191,N_1075,N_988);
nor U4192 (N_4192,N_555,N_2144);
or U4193 (N_4193,N_255,N_1915);
and U4194 (N_4194,N_166,N_1246);
and U4195 (N_4195,N_629,N_2463);
nand U4196 (N_4196,N_1148,N_1317);
nor U4197 (N_4197,N_240,N_1408);
nor U4198 (N_4198,N_1611,N_305);
nor U4199 (N_4199,N_2100,N_916);
or U4200 (N_4200,N_568,N_2181);
nor U4201 (N_4201,N_548,N_521);
nor U4202 (N_4202,N_844,N_21);
nor U4203 (N_4203,N_769,N_1463);
and U4204 (N_4204,N_685,N_397);
or U4205 (N_4205,N_2301,N_951);
nand U4206 (N_4206,N_1212,N_1982);
and U4207 (N_4207,N_1052,N_2052);
nand U4208 (N_4208,N_2136,N_1775);
or U4209 (N_4209,N_1496,N_1739);
nand U4210 (N_4210,N_2000,N_143);
or U4211 (N_4211,N_2094,N_80);
nand U4212 (N_4212,N_1536,N_1068);
and U4213 (N_4213,N_104,N_1563);
nor U4214 (N_4214,N_1313,N_793);
nor U4215 (N_4215,N_433,N_91);
or U4216 (N_4216,N_1477,N_1091);
or U4217 (N_4217,N_1130,N_456);
or U4218 (N_4218,N_2253,N_1071);
or U4219 (N_4219,N_2472,N_1146);
nand U4220 (N_4220,N_1263,N_1044);
nor U4221 (N_4221,N_422,N_554);
or U4222 (N_4222,N_363,N_60);
and U4223 (N_4223,N_447,N_668);
nand U4224 (N_4224,N_1136,N_1983);
and U4225 (N_4225,N_2460,N_2024);
or U4226 (N_4226,N_1491,N_326);
nor U4227 (N_4227,N_1467,N_662);
nand U4228 (N_4228,N_1857,N_2109);
nor U4229 (N_4229,N_88,N_1651);
and U4230 (N_4230,N_1626,N_1860);
or U4231 (N_4231,N_725,N_288);
nor U4232 (N_4232,N_1829,N_1282);
or U4233 (N_4233,N_194,N_125);
nand U4234 (N_4234,N_933,N_502);
nor U4235 (N_4235,N_1944,N_2045);
nand U4236 (N_4236,N_1373,N_359);
nand U4237 (N_4237,N_1105,N_611);
or U4238 (N_4238,N_1250,N_256);
nand U4239 (N_4239,N_1868,N_2441);
nand U4240 (N_4240,N_1372,N_1585);
nor U4241 (N_4241,N_1327,N_1360);
nand U4242 (N_4242,N_1239,N_46);
or U4243 (N_4243,N_1662,N_1194);
or U4244 (N_4244,N_728,N_867);
nor U4245 (N_4245,N_2095,N_1338);
and U4246 (N_4246,N_606,N_797);
nand U4247 (N_4247,N_1187,N_931);
nand U4248 (N_4248,N_2090,N_1745);
nor U4249 (N_4249,N_1477,N_696);
nor U4250 (N_4250,N_868,N_56);
nand U4251 (N_4251,N_115,N_1344);
or U4252 (N_4252,N_143,N_2024);
and U4253 (N_4253,N_1480,N_869);
nand U4254 (N_4254,N_43,N_1156);
nand U4255 (N_4255,N_2042,N_131);
nand U4256 (N_4256,N_1342,N_1911);
nand U4257 (N_4257,N_39,N_213);
nand U4258 (N_4258,N_533,N_152);
nor U4259 (N_4259,N_1,N_1889);
nand U4260 (N_4260,N_2296,N_1933);
nor U4261 (N_4261,N_1689,N_1802);
xor U4262 (N_4262,N_1381,N_131);
or U4263 (N_4263,N_114,N_926);
and U4264 (N_4264,N_894,N_1189);
nor U4265 (N_4265,N_1081,N_133);
nand U4266 (N_4266,N_1958,N_249);
nor U4267 (N_4267,N_85,N_1949);
and U4268 (N_4268,N_1681,N_599);
or U4269 (N_4269,N_1789,N_804);
and U4270 (N_4270,N_2401,N_2400);
or U4271 (N_4271,N_1237,N_2470);
nor U4272 (N_4272,N_2443,N_1353);
nor U4273 (N_4273,N_2167,N_473);
and U4274 (N_4274,N_681,N_859);
nand U4275 (N_4275,N_2163,N_1122);
nand U4276 (N_4276,N_978,N_1225);
nor U4277 (N_4277,N_2193,N_1896);
or U4278 (N_4278,N_2171,N_1447);
or U4279 (N_4279,N_1428,N_1394);
nand U4280 (N_4280,N_1653,N_812);
nand U4281 (N_4281,N_340,N_1732);
and U4282 (N_4282,N_81,N_1287);
or U4283 (N_4283,N_1385,N_18);
nor U4284 (N_4284,N_627,N_1625);
or U4285 (N_4285,N_2318,N_448);
nor U4286 (N_4286,N_1679,N_913);
nand U4287 (N_4287,N_533,N_696);
and U4288 (N_4288,N_1741,N_216);
or U4289 (N_4289,N_570,N_1049);
and U4290 (N_4290,N_237,N_1457);
or U4291 (N_4291,N_648,N_2496);
and U4292 (N_4292,N_2343,N_1867);
nand U4293 (N_4293,N_1899,N_2420);
nor U4294 (N_4294,N_438,N_2470);
nor U4295 (N_4295,N_104,N_13);
or U4296 (N_4296,N_656,N_1595);
or U4297 (N_4297,N_1549,N_46);
or U4298 (N_4298,N_1812,N_490);
or U4299 (N_4299,N_1878,N_152);
and U4300 (N_4300,N_1254,N_1399);
nand U4301 (N_4301,N_545,N_1437);
or U4302 (N_4302,N_1452,N_412);
nor U4303 (N_4303,N_250,N_1963);
nand U4304 (N_4304,N_587,N_1717);
and U4305 (N_4305,N_1497,N_1380);
nand U4306 (N_4306,N_1293,N_419);
and U4307 (N_4307,N_959,N_413);
or U4308 (N_4308,N_1396,N_1410);
and U4309 (N_4309,N_594,N_1141);
or U4310 (N_4310,N_27,N_1327);
or U4311 (N_4311,N_1513,N_1108);
xor U4312 (N_4312,N_1639,N_1164);
or U4313 (N_4313,N_2094,N_2150);
nor U4314 (N_4314,N_23,N_701);
nand U4315 (N_4315,N_2306,N_1857);
nor U4316 (N_4316,N_1085,N_1972);
and U4317 (N_4317,N_2067,N_1435);
nor U4318 (N_4318,N_1983,N_131);
nand U4319 (N_4319,N_1611,N_1936);
and U4320 (N_4320,N_1946,N_948);
nand U4321 (N_4321,N_258,N_1185);
and U4322 (N_4322,N_1847,N_556);
xnor U4323 (N_4323,N_712,N_1685);
nand U4324 (N_4324,N_193,N_1124);
nor U4325 (N_4325,N_1830,N_1119);
nor U4326 (N_4326,N_830,N_232);
nand U4327 (N_4327,N_422,N_132);
nor U4328 (N_4328,N_1457,N_440);
and U4329 (N_4329,N_1076,N_1582);
nand U4330 (N_4330,N_2234,N_1417);
or U4331 (N_4331,N_1786,N_518);
nand U4332 (N_4332,N_2005,N_2343);
nand U4333 (N_4333,N_108,N_2030);
and U4334 (N_4334,N_657,N_2185);
and U4335 (N_4335,N_2075,N_1727);
and U4336 (N_4336,N_1428,N_1983);
nand U4337 (N_4337,N_1215,N_840);
and U4338 (N_4338,N_912,N_1940);
and U4339 (N_4339,N_2020,N_767);
or U4340 (N_4340,N_424,N_269);
nand U4341 (N_4341,N_2443,N_687);
nand U4342 (N_4342,N_1065,N_2424);
and U4343 (N_4343,N_2110,N_1271);
or U4344 (N_4344,N_1450,N_453);
nand U4345 (N_4345,N_368,N_482);
nand U4346 (N_4346,N_510,N_946);
nor U4347 (N_4347,N_867,N_1580);
or U4348 (N_4348,N_1675,N_2065);
nor U4349 (N_4349,N_1864,N_102);
nor U4350 (N_4350,N_1947,N_212);
nand U4351 (N_4351,N_517,N_1301);
nand U4352 (N_4352,N_2491,N_1858);
or U4353 (N_4353,N_518,N_1552);
and U4354 (N_4354,N_1677,N_2042);
nand U4355 (N_4355,N_1520,N_825);
and U4356 (N_4356,N_2443,N_2492);
nor U4357 (N_4357,N_92,N_1412);
and U4358 (N_4358,N_1806,N_587);
and U4359 (N_4359,N_2166,N_2361);
nand U4360 (N_4360,N_2226,N_1574);
or U4361 (N_4361,N_1913,N_1367);
nor U4362 (N_4362,N_37,N_1129);
nand U4363 (N_4363,N_505,N_1789);
or U4364 (N_4364,N_2305,N_57);
nor U4365 (N_4365,N_1291,N_2235);
and U4366 (N_4366,N_855,N_1325);
nor U4367 (N_4367,N_133,N_810);
nor U4368 (N_4368,N_1990,N_1554);
or U4369 (N_4369,N_1790,N_1813);
nor U4370 (N_4370,N_1390,N_490);
xor U4371 (N_4371,N_530,N_2494);
and U4372 (N_4372,N_1267,N_1675);
and U4373 (N_4373,N_2186,N_192);
or U4374 (N_4374,N_1608,N_2335);
and U4375 (N_4375,N_1998,N_1233);
and U4376 (N_4376,N_1752,N_1306);
and U4377 (N_4377,N_1558,N_1925);
and U4378 (N_4378,N_257,N_1158);
or U4379 (N_4379,N_286,N_1286);
nand U4380 (N_4380,N_1029,N_520);
nand U4381 (N_4381,N_1267,N_1336);
nor U4382 (N_4382,N_2026,N_671);
nor U4383 (N_4383,N_1916,N_497);
nand U4384 (N_4384,N_1099,N_2027);
or U4385 (N_4385,N_1055,N_716);
nand U4386 (N_4386,N_905,N_707);
and U4387 (N_4387,N_2432,N_1095);
and U4388 (N_4388,N_31,N_1246);
or U4389 (N_4389,N_1820,N_1529);
nor U4390 (N_4390,N_2287,N_1842);
and U4391 (N_4391,N_1221,N_1314);
nand U4392 (N_4392,N_694,N_2175);
nor U4393 (N_4393,N_647,N_2);
or U4394 (N_4394,N_1596,N_955);
and U4395 (N_4395,N_884,N_1481);
and U4396 (N_4396,N_1950,N_1133);
and U4397 (N_4397,N_315,N_1312);
and U4398 (N_4398,N_2459,N_1225);
or U4399 (N_4399,N_261,N_1310);
nand U4400 (N_4400,N_553,N_185);
and U4401 (N_4401,N_1570,N_1032);
nand U4402 (N_4402,N_1284,N_1022);
or U4403 (N_4403,N_2146,N_328);
nand U4404 (N_4404,N_1350,N_2200);
or U4405 (N_4405,N_758,N_1022);
and U4406 (N_4406,N_2153,N_653);
nand U4407 (N_4407,N_672,N_278);
and U4408 (N_4408,N_2421,N_1520);
and U4409 (N_4409,N_952,N_1165);
nor U4410 (N_4410,N_1156,N_1622);
nand U4411 (N_4411,N_1735,N_1958);
and U4412 (N_4412,N_1012,N_66);
nand U4413 (N_4413,N_1665,N_2227);
nor U4414 (N_4414,N_1957,N_730);
nor U4415 (N_4415,N_1665,N_1557);
or U4416 (N_4416,N_1790,N_126);
nand U4417 (N_4417,N_1970,N_1679);
nor U4418 (N_4418,N_2216,N_311);
nor U4419 (N_4419,N_2438,N_755);
nor U4420 (N_4420,N_837,N_159);
and U4421 (N_4421,N_623,N_567);
and U4422 (N_4422,N_730,N_791);
nand U4423 (N_4423,N_1992,N_251);
nand U4424 (N_4424,N_458,N_1427);
or U4425 (N_4425,N_1057,N_1761);
nor U4426 (N_4426,N_1967,N_1255);
and U4427 (N_4427,N_2467,N_243);
or U4428 (N_4428,N_112,N_606);
nor U4429 (N_4429,N_1003,N_2372);
or U4430 (N_4430,N_150,N_1829);
nor U4431 (N_4431,N_2496,N_1643);
or U4432 (N_4432,N_349,N_2494);
nand U4433 (N_4433,N_2484,N_1497);
or U4434 (N_4434,N_1171,N_473);
or U4435 (N_4435,N_793,N_829);
and U4436 (N_4436,N_196,N_2467);
and U4437 (N_4437,N_2265,N_341);
nand U4438 (N_4438,N_1254,N_1208);
or U4439 (N_4439,N_974,N_727);
and U4440 (N_4440,N_1695,N_225);
and U4441 (N_4441,N_17,N_1156);
nor U4442 (N_4442,N_1764,N_2093);
nor U4443 (N_4443,N_179,N_1170);
or U4444 (N_4444,N_1233,N_1753);
nor U4445 (N_4445,N_863,N_2254);
or U4446 (N_4446,N_328,N_2318);
nand U4447 (N_4447,N_2069,N_255);
and U4448 (N_4448,N_2169,N_2079);
or U4449 (N_4449,N_1185,N_1443);
nor U4450 (N_4450,N_1327,N_2132);
nor U4451 (N_4451,N_1461,N_808);
nor U4452 (N_4452,N_1434,N_2174);
nor U4453 (N_4453,N_220,N_630);
nor U4454 (N_4454,N_601,N_401);
nand U4455 (N_4455,N_82,N_1112);
nor U4456 (N_4456,N_2168,N_2326);
or U4457 (N_4457,N_406,N_2193);
and U4458 (N_4458,N_1195,N_2202);
nand U4459 (N_4459,N_2368,N_628);
nand U4460 (N_4460,N_200,N_65);
nor U4461 (N_4461,N_597,N_1740);
or U4462 (N_4462,N_1956,N_1748);
nand U4463 (N_4463,N_1472,N_1098);
xnor U4464 (N_4464,N_2233,N_1055);
nand U4465 (N_4465,N_1516,N_581);
and U4466 (N_4466,N_864,N_2065);
nand U4467 (N_4467,N_943,N_1671);
nand U4468 (N_4468,N_688,N_1355);
nand U4469 (N_4469,N_2410,N_238);
nand U4470 (N_4470,N_2324,N_2172);
nor U4471 (N_4471,N_555,N_2454);
xnor U4472 (N_4472,N_739,N_1516);
or U4473 (N_4473,N_846,N_1564);
or U4474 (N_4474,N_1393,N_110);
or U4475 (N_4475,N_2305,N_1075);
and U4476 (N_4476,N_1916,N_1673);
or U4477 (N_4477,N_1003,N_6);
nor U4478 (N_4478,N_1191,N_2364);
or U4479 (N_4479,N_2040,N_2285);
nor U4480 (N_4480,N_1034,N_2280);
and U4481 (N_4481,N_601,N_1166);
or U4482 (N_4482,N_2018,N_1347);
nor U4483 (N_4483,N_589,N_1576);
nand U4484 (N_4484,N_719,N_108);
or U4485 (N_4485,N_165,N_2149);
and U4486 (N_4486,N_1482,N_2022);
or U4487 (N_4487,N_1864,N_490);
nor U4488 (N_4488,N_406,N_1355);
and U4489 (N_4489,N_1755,N_273);
or U4490 (N_4490,N_1757,N_228);
nor U4491 (N_4491,N_375,N_1666);
and U4492 (N_4492,N_2323,N_1798);
or U4493 (N_4493,N_20,N_1863);
nand U4494 (N_4494,N_70,N_2261);
nor U4495 (N_4495,N_903,N_1055);
and U4496 (N_4496,N_2192,N_230);
nand U4497 (N_4497,N_147,N_26);
nor U4498 (N_4498,N_2030,N_2473);
or U4499 (N_4499,N_1370,N_373);
nand U4500 (N_4500,N_2312,N_1143);
or U4501 (N_4501,N_1135,N_1087);
nor U4502 (N_4502,N_1121,N_995);
and U4503 (N_4503,N_1859,N_2371);
and U4504 (N_4504,N_861,N_1436);
or U4505 (N_4505,N_1933,N_2379);
nor U4506 (N_4506,N_835,N_16);
or U4507 (N_4507,N_1793,N_370);
and U4508 (N_4508,N_384,N_225);
nand U4509 (N_4509,N_2344,N_1857);
nand U4510 (N_4510,N_2091,N_368);
or U4511 (N_4511,N_1332,N_777);
or U4512 (N_4512,N_1840,N_2218);
nor U4513 (N_4513,N_1707,N_1354);
nor U4514 (N_4514,N_452,N_1825);
nand U4515 (N_4515,N_1129,N_517);
or U4516 (N_4516,N_839,N_446);
or U4517 (N_4517,N_292,N_1794);
or U4518 (N_4518,N_1350,N_308);
nand U4519 (N_4519,N_486,N_224);
or U4520 (N_4520,N_2368,N_1011);
nand U4521 (N_4521,N_898,N_1643);
nand U4522 (N_4522,N_1669,N_1870);
or U4523 (N_4523,N_531,N_2412);
or U4524 (N_4524,N_498,N_1339);
and U4525 (N_4525,N_2371,N_1964);
or U4526 (N_4526,N_1418,N_319);
nand U4527 (N_4527,N_836,N_1092);
nand U4528 (N_4528,N_1306,N_47);
nor U4529 (N_4529,N_2192,N_383);
nor U4530 (N_4530,N_1238,N_258);
nor U4531 (N_4531,N_862,N_2498);
nor U4532 (N_4532,N_1991,N_855);
nand U4533 (N_4533,N_2173,N_2021);
nand U4534 (N_4534,N_2337,N_207);
and U4535 (N_4535,N_193,N_1693);
nand U4536 (N_4536,N_1472,N_873);
or U4537 (N_4537,N_458,N_2203);
and U4538 (N_4538,N_293,N_1777);
or U4539 (N_4539,N_229,N_1939);
nand U4540 (N_4540,N_2408,N_1561);
and U4541 (N_4541,N_1327,N_2275);
or U4542 (N_4542,N_1396,N_2118);
and U4543 (N_4543,N_619,N_1932);
and U4544 (N_4544,N_2304,N_1395);
or U4545 (N_4545,N_713,N_515);
and U4546 (N_4546,N_1224,N_1694);
nor U4547 (N_4547,N_1959,N_1673);
nand U4548 (N_4548,N_311,N_1899);
and U4549 (N_4549,N_1652,N_2273);
or U4550 (N_4550,N_1601,N_1155);
or U4551 (N_4551,N_2008,N_23);
xnor U4552 (N_4552,N_1615,N_2128);
nor U4553 (N_4553,N_1142,N_2328);
nand U4554 (N_4554,N_1555,N_1324);
nor U4555 (N_4555,N_992,N_1391);
nor U4556 (N_4556,N_2338,N_2079);
nand U4557 (N_4557,N_2112,N_1620);
or U4558 (N_4558,N_1448,N_495);
or U4559 (N_4559,N_2397,N_2073);
or U4560 (N_4560,N_2076,N_1481);
nor U4561 (N_4561,N_1882,N_1380);
and U4562 (N_4562,N_1646,N_23);
nand U4563 (N_4563,N_1982,N_132);
nor U4564 (N_4564,N_103,N_2106);
or U4565 (N_4565,N_434,N_247);
nand U4566 (N_4566,N_1416,N_2418);
nand U4567 (N_4567,N_2170,N_495);
or U4568 (N_4568,N_263,N_1927);
or U4569 (N_4569,N_1834,N_876);
nand U4570 (N_4570,N_296,N_120);
and U4571 (N_4571,N_1973,N_864);
nor U4572 (N_4572,N_1043,N_1249);
or U4573 (N_4573,N_1354,N_363);
or U4574 (N_4574,N_2058,N_1503);
nand U4575 (N_4575,N_740,N_1919);
or U4576 (N_4576,N_1178,N_517);
and U4577 (N_4577,N_1234,N_1730);
nor U4578 (N_4578,N_1933,N_2259);
nand U4579 (N_4579,N_2030,N_776);
and U4580 (N_4580,N_168,N_1111);
nor U4581 (N_4581,N_829,N_750);
and U4582 (N_4582,N_952,N_1416);
nor U4583 (N_4583,N_8,N_903);
nand U4584 (N_4584,N_1707,N_196);
or U4585 (N_4585,N_1444,N_572);
nand U4586 (N_4586,N_1481,N_930);
or U4587 (N_4587,N_1258,N_1010);
or U4588 (N_4588,N_2127,N_1417);
and U4589 (N_4589,N_2468,N_1212);
nand U4590 (N_4590,N_1775,N_574);
nand U4591 (N_4591,N_818,N_1549);
or U4592 (N_4592,N_2258,N_2455);
nand U4593 (N_4593,N_1198,N_1444);
and U4594 (N_4594,N_1957,N_999);
nand U4595 (N_4595,N_624,N_132);
and U4596 (N_4596,N_884,N_1757);
and U4597 (N_4597,N_793,N_1306);
nand U4598 (N_4598,N_200,N_2114);
and U4599 (N_4599,N_800,N_702);
or U4600 (N_4600,N_1780,N_1763);
or U4601 (N_4601,N_1334,N_2133);
or U4602 (N_4602,N_387,N_1457);
or U4603 (N_4603,N_1291,N_954);
nor U4604 (N_4604,N_1247,N_632);
or U4605 (N_4605,N_162,N_1857);
and U4606 (N_4606,N_1907,N_1356);
nand U4607 (N_4607,N_2290,N_1240);
nand U4608 (N_4608,N_1718,N_208);
or U4609 (N_4609,N_1584,N_2041);
or U4610 (N_4610,N_859,N_690);
nand U4611 (N_4611,N_299,N_2456);
nand U4612 (N_4612,N_829,N_603);
or U4613 (N_4613,N_753,N_800);
nand U4614 (N_4614,N_1406,N_1432);
and U4615 (N_4615,N_1089,N_1140);
or U4616 (N_4616,N_715,N_2329);
or U4617 (N_4617,N_1612,N_1736);
nor U4618 (N_4618,N_2195,N_253);
nor U4619 (N_4619,N_370,N_597);
or U4620 (N_4620,N_845,N_1376);
and U4621 (N_4621,N_1040,N_1367);
nand U4622 (N_4622,N_1049,N_1863);
and U4623 (N_4623,N_94,N_549);
nor U4624 (N_4624,N_391,N_1315);
nand U4625 (N_4625,N_673,N_1856);
nand U4626 (N_4626,N_2163,N_583);
and U4627 (N_4627,N_1513,N_1950);
and U4628 (N_4628,N_1727,N_2056);
nor U4629 (N_4629,N_641,N_127);
or U4630 (N_4630,N_2102,N_620);
nor U4631 (N_4631,N_792,N_578);
or U4632 (N_4632,N_1888,N_397);
and U4633 (N_4633,N_387,N_2147);
and U4634 (N_4634,N_1129,N_1217);
or U4635 (N_4635,N_2323,N_505);
nor U4636 (N_4636,N_1233,N_437);
nand U4637 (N_4637,N_1553,N_711);
or U4638 (N_4638,N_351,N_2148);
or U4639 (N_4639,N_622,N_1440);
nor U4640 (N_4640,N_1978,N_710);
nor U4641 (N_4641,N_462,N_1033);
nand U4642 (N_4642,N_1599,N_2312);
nor U4643 (N_4643,N_1424,N_2460);
nor U4644 (N_4644,N_866,N_1882);
and U4645 (N_4645,N_1549,N_2265);
or U4646 (N_4646,N_31,N_162);
nand U4647 (N_4647,N_132,N_878);
nand U4648 (N_4648,N_2121,N_1767);
or U4649 (N_4649,N_1133,N_1375);
nor U4650 (N_4650,N_2011,N_2250);
or U4651 (N_4651,N_212,N_119);
nand U4652 (N_4652,N_808,N_2447);
or U4653 (N_4653,N_751,N_1812);
nand U4654 (N_4654,N_114,N_1831);
and U4655 (N_4655,N_310,N_1840);
and U4656 (N_4656,N_2093,N_1797);
nor U4657 (N_4657,N_2133,N_2408);
nor U4658 (N_4658,N_2466,N_587);
and U4659 (N_4659,N_31,N_1298);
nor U4660 (N_4660,N_1798,N_230);
nor U4661 (N_4661,N_2119,N_705);
and U4662 (N_4662,N_783,N_899);
nor U4663 (N_4663,N_43,N_1595);
nand U4664 (N_4664,N_849,N_1939);
nor U4665 (N_4665,N_315,N_1763);
nor U4666 (N_4666,N_402,N_802);
and U4667 (N_4667,N_2455,N_827);
nand U4668 (N_4668,N_387,N_2350);
nor U4669 (N_4669,N_1415,N_1400);
or U4670 (N_4670,N_2142,N_1573);
or U4671 (N_4671,N_1687,N_760);
nor U4672 (N_4672,N_1795,N_1584);
or U4673 (N_4673,N_1503,N_1284);
nor U4674 (N_4674,N_641,N_2017);
and U4675 (N_4675,N_141,N_1978);
or U4676 (N_4676,N_2206,N_1549);
nor U4677 (N_4677,N_2074,N_6);
or U4678 (N_4678,N_1561,N_2036);
and U4679 (N_4679,N_1819,N_2294);
nand U4680 (N_4680,N_428,N_1082);
nand U4681 (N_4681,N_1674,N_1057);
nor U4682 (N_4682,N_799,N_958);
or U4683 (N_4683,N_1153,N_739);
nor U4684 (N_4684,N_1936,N_1984);
nor U4685 (N_4685,N_155,N_2457);
and U4686 (N_4686,N_2112,N_468);
nor U4687 (N_4687,N_1977,N_606);
or U4688 (N_4688,N_30,N_207);
or U4689 (N_4689,N_1514,N_808);
or U4690 (N_4690,N_828,N_1758);
nor U4691 (N_4691,N_443,N_784);
and U4692 (N_4692,N_1481,N_1460);
nand U4693 (N_4693,N_1916,N_600);
nand U4694 (N_4694,N_1372,N_943);
or U4695 (N_4695,N_1184,N_536);
nand U4696 (N_4696,N_1277,N_2119);
nand U4697 (N_4697,N_479,N_225);
nand U4698 (N_4698,N_2008,N_22);
or U4699 (N_4699,N_824,N_2274);
and U4700 (N_4700,N_1254,N_2276);
and U4701 (N_4701,N_800,N_1942);
nand U4702 (N_4702,N_1350,N_405);
nor U4703 (N_4703,N_802,N_1940);
nand U4704 (N_4704,N_1349,N_2098);
and U4705 (N_4705,N_160,N_663);
nand U4706 (N_4706,N_55,N_1300);
and U4707 (N_4707,N_962,N_1931);
xnor U4708 (N_4708,N_2104,N_2468);
nor U4709 (N_4709,N_1165,N_390);
nand U4710 (N_4710,N_1967,N_1957);
nand U4711 (N_4711,N_49,N_603);
nor U4712 (N_4712,N_2025,N_1077);
nor U4713 (N_4713,N_1243,N_408);
nor U4714 (N_4714,N_2337,N_1312);
or U4715 (N_4715,N_730,N_859);
xnor U4716 (N_4716,N_1619,N_1079);
nor U4717 (N_4717,N_1050,N_1868);
or U4718 (N_4718,N_1120,N_2082);
nand U4719 (N_4719,N_363,N_1971);
nor U4720 (N_4720,N_1988,N_917);
nor U4721 (N_4721,N_1328,N_1860);
and U4722 (N_4722,N_1082,N_1986);
nand U4723 (N_4723,N_1383,N_956);
nand U4724 (N_4724,N_240,N_2361);
or U4725 (N_4725,N_617,N_2222);
nand U4726 (N_4726,N_1221,N_2147);
and U4727 (N_4727,N_2347,N_2058);
nor U4728 (N_4728,N_619,N_641);
and U4729 (N_4729,N_709,N_2406);
or U4730 (N_4730,N_467,N_640);
or U4731 (N_4731,N_1522,N_1655);
and U4732 (N_4732,N_28,N_1453);
and U4733 (N_4733,N_375,N_792);
xnor U4734 (N_4734,N_1180,N_2196);
nor U4735 (N_4735,N_30,N_200);
and U4736 (N_4736,N_400,N_875);
nor U4737 (N_4737,N_2213,N_934);
nor U4738 (N_4738,N_2181,N_1013);
and U4739 (N_4739,N_65,N_76);
and U4740 (N_4740,N_2391,N_395);
or U4741 (N_4741,N_752,N_5);
nor U4742 (N_4742,N_1527,N_2226);
nand U4743 (N_4743,N_2078,N_939);
and U4744 (N_4744,N_1772,N_307);
and U4745 (N_4745,N_477,N_541);
and U4746 (N_4746,N_2090,N_977);
and U4747 (N_4747,N_1707,N_713);
nor U4748 (N_4748,N_2187,N_124);
and U4749 (N_4749,N_2387,N_1457);
nor U4750 (N_4750,N_2065,N_359);
or U4751 (N_4751,N_376,N_2288);
or U4752 (N_4752,N_2493,N_294);
and U4753 (N_4753,N_2188,N_705);
nand U4754 (N_4754,N_505,N_840);
and U4755 (N_4755,N_201,N_2083);
nand U4756 (N_4756,N_570,N_360);
and U4757 (N_4757,N_151,N_480);
and U4758 (N_4758,N_200,N_487);
nand U4759 (N_4759,N_1444,N_1015);
or U4760 (N_4760,N_2181,N_1288);
and U4761 (N_4761,N_1996,N_1768);
nor U4762 (N_4762,N_1064,N_797);
nor U4763 (N_4763,N_1678,N_7);
nor U4764 (N_4764,N_1830,N_2376);
or U4765 (N_4765,N_373,N_1582);
and U4766 (N_4766,N_1405,N_2420);
nand U4767 (N_4767,N_444,N_2069);
or U4768 (N_4768,N_2026,N_85);
or U4769 (N_4769,N_375,N_630);
and U4770 (N_4770,N_181,N_961);
and U4771 (N_4771,N_970,N_2157);
nor U4772 (N_4772,N_996,N_1312);
and U4773 (N_4773,N_793,N_2484);
and U4774 (N_4774,N_225,N_189);
or U4775 (N_4775,N_2332,N_1118);
or U4776 (N_4776,N_2230,N_225);
nand U4777 (N_4777,N_2454,N_379);
nand U4778 (N_4778,N_2361,N_335);
nor U4779 (N_4779,N_1198,N_863);
or U4780 (N_4780,N_2044,N_1996);
or U4781 (N_4781,N_1389,N_2351);
nand U4782 (N_4782,N_922,N_2269);
and U4783 (N_4783,N_906,N_1266);
nor U4784 (N_4784,N_1075,N_1934);
or U4785 (N_4785,N_3,N_1769);
and U4786 (N_4786,N_386,N_2238);
nand U4787 (N_4787,N_678,N_770);
nand U4788 (N_4788,N_506,N_2080);
nor U4789 (N_4789,N_1866,N_1023);
nor U4790 (N_4790,N_494,N_2188);
nand U4791 (N_4791,N_2452,N_2203);
and U4792 (N_4792,N_2200,N_1557);
or U4793 (N_4793,N_2101,N_860);
nor U4794 (N_4794,N_2146,N_1029);
nand U4795 (N_4795,N_815,N_1485);
nor U4796 (N_4796,N_1160,N_961);
or U4797 (N_4797,N_543,N_237);
nand U4798 (N_4798,N_1362,N_1520);
or U4799 (N_4799,N_109,N_1668);
nor U4800 (N_4800,N_1552,N_1357);
nand U4801 (N_4801,N_991,N_2273);
or U4802 (N_4802,N_643,N_1677);
and U4803 (N_4803,N_1554,N_1972);
or U4804 (N_4804,N_147,N_951);
nor U4805 (N_4805,N_475,N_263);
and U4806 (N_4806,N_1273,N_2490);
nand U4807 (N_4807,N_2019,N_2336);
nand U4808 (N_4808,N_996,N_2250);
nand U4809 (N_4809,N_1508,N_1450);
and U4810 (N_4810,N_1268,N_488);
and U4811 (N_4811,N_440,N_426);
nand U4812 (N_4812,N_826,N_2287);
nand U4813 (N_4813,N_226,N_1287);
nor U4814 (N_4814,N_1986,N_602);
and U4815 (N_4815,N_622,N_1990);
or U4816 (N_4816,N_538,N_24);
nor U4817 (N_4817,N_1734,N_2430);
or U4818 (N_4818,N_2012,N_626);
nand U4819 (N_4819,N_864,N_1879);
nand U4820 (N_4820,N_2330,N_348);
or U4821 (N_4821,N_2250,N_1506);
xor U4822 (N_4822,N_956,N_2366);
nand U4823 (N_4823,N_930,N_30);
or U4824 (N_4824,N_902,N_880);
nor U4825 (N_4825,N_872,N_19);
nor U4826 (N_4826,N_2132,N_1697);
or U4827 (N_4827,N_1871,N_2371);
and U4828 (N_4828,N_504,N_876);
nand U4829 (N_4829,N_1503,N_1472);
nor U4830 (N_4830,N_1089,N_1357);
and U4831 (N_4831,N_1695,N_461);
or U4832 (N_4832,N_2415,N_453);
or U4833 (N_4833,N_2026,N_1084);
nor U4834 (N_4834,N_2459,N_756);
and U4835 (N_4835,N_1540,N_819);
nand U4836 (N_4836,N_2397,N_1243);
nor U4837 (N_4837,N_278,N_238);
nor U4838 (N_4838,N_704,N_1557);
nor U4839 (N_4839,N_6,N_713);
nor U4840 (N_4840,N_540,N_1808);
and U4841 (N_4841,N_775,N_2148);
nand U4842 (N_4842,N_120,N_501);
nand U4843 (N_4843,N_811,N_1392);
xnor U4844 (N_4844,N_2299,N_1);
and U4845 (N_4845,N_1438,N_762);
xnor U4846 (N_4846,N_853,N_2479);
nor U4847 (N_4847,N_1364,N_1409);
nand U4848 (N_4848,N_1977,N_1623);
nor U4849 (N_4849,N_2178,N_894);
and U4850 (N_4850,N_2288,N_2121);
nor U4851 (N_4851,N_2257,N_1133);
nor U4852 (N_4852,N_106,N_1204);
xnor U4853 (N_4853,N_1653,N_449);
or U4854 (N_4854,N_1828,N_1027);
nand U4855 (N_4855,N_1490,N_34);
and U4856 (N_4856,N_1512,N_2391);
or U4857 (N_4857,N_76,N_945);
nand U4858 (N_4858,N_1719,N_1917);
and U4859 (N_4859,N_767,N_149);
nand U4860 (N_4860,N_418,N_1791);
nand U4861 (N_4861,N_595,N_601);
and U4862 (N_4862,N_1723,N_1438);
and U4863 (N_4863,N_2403,N_1421);
and U4864 (N_4864,N_672,N_1888);
and U4865 (N_4865,N_105,N_860);
or U4866 (N_4866,N_787,N_1537);
nand U4867 (N_4867,N_2247,N_1433);
and U4868 (N_4868,N_1287,N_386);
or U4869 (N_4869,N_1903,N_2166);
and U4870 (N_4870,N_1021,N_1016);
nor U4871 (N_4871,N_2419,N_2259);
and U4872 (N_4872,N_2168,N_469);
nor U4873 (N_4873,N_152,N_187);
nor U4874 (N_4874,N_191,N_1385);
nand U4875 (N_4875,N_2111,N_1185);
or U4876 (N_4876,N_1013,N_390);
and U4877 (N_4877,N_2367,N_528);
and U4878 (N_4878,N_1997,N_1592);
or U4879 (N_4879,N_232,N_790);
nand U4880 (N_4880,N_2426,N_1208);
and U4881 (N_4881,N_1758,N_1263);
nand U4882 (N_4882,N_1603,N_1521);
and U4883 (N_4883,N_234,N_2203);
nand U4884 (N_4884,N_542,N_1175);
nor U4885 (N_4885,N_1057,N_2188);
or U4886 (N_4886,N_1431,N_404);
or U4887 (N_4887,N_1206,N_1129);
nand U4888 (N_4888,N_1871,N_2380);
nand U4889 (N_4889,N_163,N_1642);
or U4890 (N_4890,N_1961,N_1966);
and U4891 (N_4891,N_954,N_111);
nor U4892 (N_4892,N_1855,N_642);
or U4893 (N_4893,N_233,N_1592);
nor U4894 (N_4894,N_1204,N_52);
nor U4895 (N_4895,N_1644,N_1002);
or U4896 (N_4896,N_813,N_468);
or U4897 (N_4897,N_850,N_2114);
nor U4898 (N_4898,N_439,N_696);
or U4899 (N_4899,N_53,N_102);
or U4900 (N_4900,N_2306,N_621);
nand U4901 (N_4901,N_2394,N_159);
nand U4902 (N_4902,N_1678,N_653);
and U4903 (N_4903,N_260,N_1492);
nand U4904 (N_4904,N_2150,N_2012);
or U4905 (N_4905,N_1765,N_1826);
nand U4906 (N_4906,N_1073,N_1009);
nand U4907 (N_4907,N_1675,N_700);
nand U4908 (N_4908,N_1335,N_796);
or U4909 (N_4909,N_2066,N_1831);
nor U4910 (N_4910,N_796,N_157);
nor U4911 (N_4911,N_139,N_260);
or U4912 (N_4912,N_191,N_1524);
or U4913 (N_4913,N_2055,N_1433);
or U4914 (N_4914,N_807,N_2323);
or U4915 (N_4915,N_583,N_625);
nor U4916 (N_4916,N_1790,N_93);
xnor U4917 (N_4917,N_1285,N_684);
nand U4918 (N_4918,N_2150,N_1178);
nand U4919 (N_4919,N_1523,N_1624);
nor U4920 (N_4920,N_1280,N_1039);
nand U4921 (N_4921,N_5,N_129);
or U4922 (N_4922,N_524,N_1041);
xor U4923 (N_4923,N_1157,N_1069);
or U4924 (N_4924,N_76,N_1414);
or U4925 (N_4925,N_974,N_2251);
or U4926 (N_4926,N_1175,N_1716);
nor U4927 (N_4927,N_1335,N_1714);
nand U4928 (N_4928,N_1775,N_1681);
or U4929 (N_4929,N_2118,N_2475);
nor U4930 (N_4930,N_2006,N_1642);
and U4931 (N_4931,N_656,N_285);
and U4932 (N_4932,N_1110,N_2018);
nand U4933 (N_4933,N_116,N_73);
and U4934 (N_4934,N_2104,N_1402);
nand U4935 (N_4935,N_631,N_93);
nor U4936 (N_4936,N_1213,N_2341);
nor U4937 (N_4937,N_994,N_1927);
or U4938 (N_4938,N_635,N_757);
nand U4939 (N_4939,N_556,N_1472);
or U4940 (N_4940,N_2116,N_2056);
nand U4941 (N_4941,N_2062,N_354);
and U4942 (N_4942,N_1820,N_1139);
and U4943 (N_4943,N_233,N_1265);
nor U4944 (N_4944,N_1429,N_462);
nand U4945 (N_4945,N_973,N_948);
nand U4946 (N_4946,N_1695,N_1760);
and U4947 (N_4947,N_1992,N_1525);
or U4948 (N_4948,N_1814,N_1763);
and U4949 (N_4949,N_1465,N_2297);
and U4950 (N_4950,N_2256,N_1780);
nor U4951 (N_4951,N_909,N_37);
nand U4952 (N_4952,N_1852,N_332);
nor U4953 (N_4953,N_1799,N_900);
nand U4954 (N_4954,N_2496,N_1277);
nor U4955 (N_4955,N_2408,N_1238);
and U4956 (N_4956,N_1958,N_140);
and U4957 (N_4957,N_858,N_414);
nor U4958 (N_4958,N_458,N_1933);
nor U4959 (N_4959,N_524,N_78);
or U4960 (N_4960,N_551,N_1382);
nor U4961 (N_4961,N_847,N_34);
or U4962 (N_4962,N_1255,N_848);
and U4963 (N_4963,N_1805,N_1221);
nand U4964 (N_4964,N_1094,N_264);
nor U4965 (N_4965,N_2293,N_1896);
and U4966 (N_4966,N_1669,N_2292);
nand U4967 (N_4967,N_1535,N_1846);
and U4968 (N_4968,N_57,N_1792);
xor U4969 (N_4969,N_384,N_1367);
nand U4970 (N_4970,N_265,N_388);
nor U4971 (N_4971,N_1105,N_455);
nand U4972 (N_4972,N_784,N_1819);
nor U4973 (N_4973,N_1315,N_483);
nor U4974 (N_4974,N_1459,N_1113);
or U4975 (N_4975,N_2061,N_1974);
nor U4976 (N_4976,N_639,N_12);
nor U4977 (N_4977,N_1191,N_2121);
nor U4978 (N_4978,N_2428,N_573);
nor U4979 (N_4979,N_2185,N_1870);
nand U4980 (N_4980,N_941,N_761);
nand U4981 (N_4981,N_908,N_1282);
nand U4982 (N_4982,N_896,N_531);
nand U4983 (N_4983,N_2096,N_1228);
and U4984 (N_4984,N_1669,N_418);
nand U4985 (N_4985,N_1105,N_65);
or U4986 (N_4986,N_2277,N_1203);
or U4987 (N_4987,N_1911,N_1758);
and U4988 (N_4988,N_1976,N_1623);
nand U4989 (N_4989,N_2482,N_2427);
nand U4990 (N_4990,N_947,N_2223);
and U4991 (N_4991,N_360,N_1054);
nand U4992 (N_4992,N_1682,N_1623);
or U4993 (N_4993,N_1153,N_2092);
nand U4994 (N_4994,N_128,N_2327);
or U4995 (N_4995,N_1544,N_1581);
and U4996 (N_4996,N_2184,N_2077);
nand U4997 (N_4997,N_2037,N_2290);
nand U4998 (N_4998,N_1376,N_656);
or U4999 (N_4999,N_697,N_1838);
nor UO_0 (O_0,N_4762,N_3213);
or UO_1 (O_1,N_2555,N_3752);
nand UO_2 (O_2,N_2592,N_3269);
xnor UO_3 (O_3,N_4331,N_2812);
nor UO_4 (O_4,N_4296,N_3224);
or UO_5 (O_5,N_4703,N_4832);
nand UO_6 (O_6,N_3415,N_4897);
nand UO_7 (O_7,N_3876,N_3483);
or UO_8 (O_8,N_3361,N_2605);
xnor UO_9 (O_9,N_4694,N_2781);
nor UO_10 (O_10,N_3428,N_3732);
or UO_11 (O_11,N_4979,N_4496);
nand UO_12 (O_12,N_2755,N_4308);
or UO_13 (O_13,N_2510,N_4605);
or UO_14 (O_14,N_3372,N_4285);
or UO_15 (O_15,N_4109,N_3206);
nand UO_16 (O_16,N_3639,N_4568);
or UO_17 (O_17,N_3823,N_3897);
nor UO_18 (O_18,N_4595,N_4314);
or UO_19 (O_19,N_3866,N_3848);
nor UO_20 (O_20,N_3416,N_3827);
nand UO_21 (O_21,N_4934,N_3649);
and UO_22 (O_22,N_4615,N_3507);
nor UO_23 (O_23,N_2545,N_2798);
or UO_24 (O_24,N_3395,N_3004);
and UO_25 (O_25,N_4561,N_3905);
and UO_26 (O_26,N_4952,N_3444);
or UO_27 (O_27,N_3700,N_4607);
or UO_28 (O_28,N_3977,N_2550);
nand UO_29 (O_29,N_4825,N_2949);
and UO_30 (O_30,N_4185,N_3646);
nand UO_31 (O_31,N_2867,N_4249);
and UO_32 (O_32,N_4685,N_2787);
nor UO_33 (O_33,N_2788,N_3344);
or UO_34 (O_34,N_4833,N_3571);
and UO_35 (O_35,N_4881,N_4333);
nand UO_36 (O_36,N_4553,N_2601);
and UO_37 (O_37,N_3185,N_4131);
nor UO_38 (O_38,N_4537,N_3329);
or UO_39 (O_39,N_4947,N_3653);
and UO_40 (O_40,N_3859,N_3586);
or UO_41 (O_41,N_4778,N_4542);
or UO_42 (O_42,N_3020,N_4978);
nand UO_43 (O_43,N_4468,N_4338);
nor UO_44 (O_44,N_4182,N_4323);
nand UO_45 (O_45,N_3760,N_3676);
or UO_46 (O_46,N_3898,N_3712);
and UO_47 (O_47,N_3660,N_2664);
nand UO_48 (O_48,N_3380,N_4573);
or UO_49 (O_49,N_2839,N_3478);
nand UO_50 (O_50,N_3750,N_3735);
nand UO_51 (O_51,N_4115,N_3006);
nor UO_52 (O_52,N_4655,N_4889);
nor UO_53 (O_53,N_3045,N_2843);
nand UO_54 (O_54,N_4016,N_3265);
nand UO_55 (O_55,N_3078,N_3641);
and UO_56 (O_56,N_3039,N_2985);
nor UO_57 (O_57,N_4558,N_4158);
nor UO_58 (O_58,N_2674,N_3999);
nand UO_59 (O_59,N_2777,N_3031);
nand UO_60 (O_60,N_3799,N_3057);
xnor UO_61 (O_61,N_3980,N_2847);
nor UO_62 (O_62,N_3715,N_2842);
nand UO_63 (O_63,N_3550,N_2871);
nor UO_64 (O_64,N_4671,N_3205);
nor UO_65 (O_65,N_3665,N_2604);
nand UO_66 (O_66,N_4309,N_4312);
nand UO_67 (O_67,N_2958,N_2786);
or UO_68 (O_68,N_3461,N_3446);
nor UO_69 (O_69,N_3535,N_2508);
and UO_70 (O_70,N_3277,N_4359);
and UO_71 (O_71,N_4099,N_4053);
or UO_72 (O_72,N_4820,N_4302);
nand UO_73 (O_73,N_3592,N_3734);
nor UO_74 (O_74,N_3605,N_3894);
or UO_75 (O_75,N_3606,N_4530);
or UO_76 (O_76,N_4996,N_4780);
or UO_77 (O_77,N_2589,N_3148);
nand UO_78 (O_78,N_3474,N_4365);
nor UO_79 (O_79,N_4596,N_2893);
nor UO_80 (O_80,N_3864,N_4394);
nor UO_81 (O_81,N_4387,N_3059);
or UO_82 (O_82,N_3456,N_2894);
nor UO_83 (O_83,N_4692,N_3939);
or UO_84 (O_84,N_2710,N_3194);
and UO_85 (O_85,N_4100,N_2935);
or UO_86 (O_86,N_4608,N_3947);
and UO_87 (O_87,N_4645,N_2502);
nand UO_88 (O_88,N_4725,N_4948);
or UO_89 (O_89,N_3383,N_4391);
nor UO_90 (O_90,N_3289,N_3011);
and UO_91 (O_91,N_4698,N_3617);
and UO_92 (O_92,N_4601,N_4098);
nand UO_93 (O_93,N_2831,N_2566);
and UO_94 (O_94,N_3008,N_3384);
nor UO_95 (O_95,N_3239,N_3637);
or UO_96 (O_96,N_2828,N_3249);
nand UO_97 (O_97,N_4386,N_2715);
and UO_98 (O_98,N_2908,N_3154);
nand UO_99 (O_99,N_4231,N_3235);
or UO_100 (O_100,N_3172,N_3303);
nor UO_101 (O_101,N_4423,N_3309);
nand UO_102 (O_102,N_4905,N_2793);
nor UO_103 (O_103,N_3187,N_3800);
or UO_104 (O_104,N_3447,N_2602);
or UO_105 (O_105,N_2688,N_4372);
or UO_106 (O_106,N_3498,N_4027);
nor UO_107 (O_107,N_2753,N_4173);
nand UO_108 (O_108,N_3690,N_3944);
or UO_109 (O_109,N_4872,N_4475);
or UO_110 (O_110,N_4926,N_4627);
and UO_111 (O_111,N_2872,N_2918);
nand UO_112 (O_112,N_3502,N_3257);
nand UO_113 (O_113,N_2695,N_4752);
nor UO_114 (O_114,N_3324,N_4519);
nand UO_115 (O_115,N_3557,N_4770);
nand UO_116 (O_116,N_3843,N_4495);
or UO_117 (O_117,N_3949,N_3515);
or UO_118 (O_118,N_4536,N_3293);
or UO_119 (O_119,N_4667,N_4265);
or UO_120 (O_120,N_4126,N_3563);
nand UO_121 (O_121,N_3354,N_3072);
or UO_122 (O_122,N_3844,N_3788);
or UO_123 (O_123,N_4712,N_3394);
nor UO_124 (O_124,N_3386,N_4317);
or UO_125 (O_125,N_3540,N_4807);
and UO_126 (O_126,N_2690,N_4543);
and UO_127 (O_127,N_2578,N_4818);
and UO_128 (O_128,N_4850,N_4447);
nor UO_129 (O_129,N_3625,N_2532);
nor UO_130 (O_130,N_4682,N_4942);
nand UO_131 (O_131,N_3382,N_3005);
and UO_132 (O_132,N_4117,N_3555);
xor UO_133 (O_133,N_2963,N_4229);
and UO_134 (O_134,N_2584,N_2683);
nor UO_135 (O_135,N_4188,N_4529);
or UO_136 (O_136,N_4389,N_4533);
and UO_137 (O_137,N_4963,N_3149);
or UO_138 (O_138,N_3623,N_3385);
or UO_139 (O_139,N_3163,N_4665);
or UO_140 (O_140,N_4041,N_4883);
nor UO_141 (O_141,N_3188,N_4194);
nand UO_142 (O_142,N_4436,N_4234);
nor UO_143 (O_143,N_4001,N_2892);
nor UO_144 (O_144,N_3445,N_3694);
and UO_145 (O_145,N_3778,N_3040);
or UO_146 (O_146,N_4499,N_2626);
or UO_147 (O_147,N_3353,N_3452);
nor UO_148 (O_148,N_3513,N_2512);
or UO_149 (O_149,N_3377,N_3680);
nand UO_150 (O_150,N_3400,N_4036);
xnor UO_151 (O_151,N_4798,N_3632);
and UO_152 (O_152,N_4767,N_3921);
xnor UO_153 (O_153,N_3294,N_3122);
nor UO_154 (O_154,N_4998,N_3202);
nand UO_155 (O_155,N_4823,N_3412);
nor UO_156 (O_156,N_4886,N_3655);
and UO_157 (O_157,N_4494,N_2511);
nand UO_158 (O_158,N_4754,N_4782);
nor UO_159 (O_159,N_3743,N_3465);
and UO_160 (O_160,N_3728,N_4364);
nand UO_161 (O_161,N_4751,N_2611);
nand UO_162 (O_162,N_2764,N_3260);
or UO_163 (O_163,N_3609,N_3169);
or UO_164 (O_164,N_4631,N_3270);
nor UO_165 (O_165,N_4708,N_4478);
nor UO_166 (O_166,N_2760,N_4498);
and UO_167 (O_167,N_3969,N_4300);
nand UO_168 (O_168,N_4461,N_4283);
nand UO_169 (O_169,N_3030,N_4409);
or UO_170 (O_170,N_3913,N_3583);
or UO_171 (O_171,N_4865,N_4813);
nand UO_172 (O_172,N_3620,N_4895);
or UO_173 (O_173,N_3339,N_4792);
xnor UO_174 (O_174,N_3076,N_2821);
or UO_175 (O_175,N_4235,N_4371);
nor UO_176 (O_176,N_4467,N_2616);
and UO_177 (O_177,N_2628,N_2932);
nand UO_178 (O_178,N_4735,N_3387);
nor UO_179 (O_179,N_4641,N_2906);
and UO_180 (O_180,N_2878,N_2917);
nor UO_181 (O_181,N_3526,N_4544);
or UO_182 (O_182,N_3741,N_3902);
nand UO_183 (O_183,N_4147,N_2704);
and UO_184 (O_184,N_4404,N_3120);
nand UO_185 (O_185,N_3796,N_4609);
or UO_186 (O_186,N_4878,N_4078);
nand UO_187 (O_187,N_3215,N_3577);
and UO_188 (O_188,N_3785,N_4839);
nor UO_189 (O_189,N_3692,N_3159);
or UO_190 (O_190,N_3895,N_4175);
nand UO_191 (O_191,N_4121,N_4012);
nor UO_192 (O_192,N_3325,N_4471);
and UO_193 (O_193,N_4280,N_3698);
nand UO_194 (O_194,N_2692,N_4955);
or UO_195 (O_195,N_2724,N_3765);
nand UO_196 (O_196,N_4857,N_2748);
nand UO_197 (O_197,N_4753,N_4428);
and UO_198 (O_198,N_2634,N_4965);
nand UO_199 (O_199,N_3141,N_4245);
nor UO_200 (O_200,N_4771,N_4431);
or UO_201 (O_201,N_4750,N_4438);
or UO_202 (O_202,N_3761,N_4023);
nor UO_203 (O_203,N_4258,N_2854);
and UO_204 (O_204,N_4113,N_3579);
or UO_205 (O_205,N_2557,N_4209);
and UO_206 (O_206,N_3705,N_4554);
or UO_207 (O_207,N_3495,N_4055);
nor UO_208 (O_208,N_4124,N_4246);
nand UO_209 (O_209,N_4637,N_2779);
nand UO_210 (O_210,N_3539,N_2808);
and UO_211 (O_211,N_2727,N_3287);
nand UO_212 (O_212,N_2513,N_4212);
or UO_213 (O_213,N_2740,N_2817);
nor UO_214 (O_214,N_4524,N_4384);
nand UO_215 (O_215,N_3246,N_4274);
or UO_216 (O_216,N_3909,N_4061);
or UO_217 (O_217,N_3716,N_4619);
and UO_218 (O_218,N_3389,N_4784);
nand UO_219 (O_219,N_2944,N_4731);
nor UO_220 (O_220,N_4038,N_4821);
or UO_221 (O_221,N_3168,N_4672);
nand UO_222 (O_222,N_4282,N_4487);
and UO_223 (O_223,N_4341,N_3390);
nand UO_224 (O_224,N_3589,N_4211);
nand UO_225 (O_225,N_4827,N_3580);
or UO_226 (O_226,N_4740,N_4340);
nor UO_227 (O_227,N_4303,N_4856);
nor UO_228 (O_228,N_2920,N_3553);
or UO_229 (O_229,N_4977,N_4935);
and UO_230 (O_230,N_4485,N_4128);
and UO_231 (O_231,N_4462,N_4638);
and UO_232 (O_232,N_3834,N_4974);
or UO_233 (O_233,N_2890,N_4982);
nand UO_234 (O_234,N_4921,N_3244);
or UO_235 (O_235,N_3401,N_4799);
or UO_236 (O_236,N_4819,N_4367);
nor UO_237 (O_237,N_4029,N_4097);
nor UO_238 (O_238,N_3467,N_4408);
nor UO_239 (O_239,N_4032,N_3178);
and UO_240 (O_240,N_2732,N_4149);
and UO_241 (O_241,N_4907,N_3508);
nor UO_242 (O_242,N_2758,N_3469);
nand UO_243 (O_243,N_4310,N_2687);
or UO_244 (O_244,N_3845,N_4973);
and UO_245 (O_245,N_4024,N_3892);
nor UO_246 (O_246,N_2883,N_4477);
nand UO_247 (O_247,N_3094,N_3127);
nor UO_248 (O_248,N_3731,N_4956);
nor UO_249 (O_249,N_4118,N_4442);
nor UO_250 (O_250,N_4186,N_4758);
or UO_251 (O_251,N_3745,N_4621);
and UO_252 (O_252,N_4505,N_3098);
nor UO_253 (O_253,N_4911,N_3096);
and UO_254 (O_254,N_4720,N_2603);
nand UO_255 (O_255,N_3802,N_3925);
or UO_256 (O_256,N_3114,N_3125);
and UO_257 (O_257,N_4060,N_2619);
nand UO_258 (O_258,N_4772,N_2708);
or UO_259 (O_259,N_2627,N_3597);
and UO_260 (O_260,N_2743,N_3422);
and UO_261 (O_261,N_2676,N_4575);
nor UO_262 (O_262,N_3146,N_3587);
nand UO_263 (O_263,N_3243,N_2823);
and UO_264 (O_264,N_2919,N_2610);
nand UO_265 (O_265,N_3774,N_4616);
or UO_266 (O_266,N_3408,N_4915);
or UO_267 (O_267,N_3972,N_4557);
nor UO_268 (O_268,N_4624,N_3704);
or UO_269 (O_269,N_4342,N_4794);
and UO_270 (O_270,N_2863,N_3493);
nor UO_271 (O_271,N_3248,N_3798);
xor UO_272 (O_272,N_4178,N_3320);
nand UO_273 (O_273,N_3861,N_4674);
and UO_274 (O_274,N_2803,N_3307);
nand UO_275 (O_275,N_4855,N_2929);
and UO_276 (O_276,N_4723,N_3170);
nand UO_277 (O_277,N_3863,N_4801);
or UO_278 (O_278,N_2606,N_3024);
nor UO_279 (O_279,N_3562,N_3811);
nor UO_280 (O_280,N_3706,N_3975);
and UO_281 (O_281,N_4961,N_4547);
or UO_282 (O_282,N_4125,N_2845);
and UO_283 (O_283,N_3564,N_3790);
nand UO_284 (O_284,N_3272,N_3840);
nor UO_285 (O_285,N_3105,N_4663);
and UO_286 (O_286,N_4183,N_3714);
nand UO_287 (O_287,N_4497,N_2543);
nand UO_288 (O_288,N_3573,N_4453);
nor UO_289 (O_289,N_3253,N_4717);
nand UO_290 (O_290,N_3523,N_3090);
or UO_291 (O_291,N_2940,N_3533);
nand UO_292 (O_292,N_2665,N_2765);
nand UO_293 (O_293,N_4888,N_4031);
nor UO_294 (O_294,N_3021,N_2588);
nor UO_295 (O_295,N_4220,N_4719);
and UO_296 (O_296,N_3060,N_4083);
nor UO_297 (O_297,N_2534,N_3251);
nand UO_298 (O_298,N_4373,N_3881);
nor UO_299 (O_299,N_2819,N_4744);
and UO_300 (O_300,N_2934,N_3266);
and UO_301 (O_301,N_4287,N_4702);
nor UO_302 (O_302,N_4757,N_3695);
nand UO_303 (O_303,N_3548,N_4434);
and UO_304 (O_304,N_3499,N_3711);
nand UO_305 (O_305,N_3849,N_3392);
and UO_306 (O_306,N_3262,N_4670);
and UO_307 (O_307,N_2542,N_3989);
nand UO_308 (O_308,N_3544,N_4347);
nor UO_309 (O_309,N_2910,N_3216);
or UO_310 (O_310,N_3247,N_4000);
and UO_311 (O_311,N_3914,N_3904);
nor UO_312 (O_312,N_4854,N_3922);
nor UO_313 (O_313,N_3979,N_4876);
and UO_314 (O_314,N_4983,N_4625);
nor UO_315 (O_315,N_3055,N_4361);
nor UO_316 (O_316,N_3846,N_3087);
nor UO_317 (O_317,N_3927,N_4874);
or UO_318 (O_318,N_3691,N_2586);
nand UO_319 (O_319,N_4301,N_3074);
and UO_320 (O_320,N_3803,N_3349);
and UO_321 (O_321,N_4228,N_3988);
xor UO_322 (O_322,N_2595,N_3402);
xnor UO_323 (O_323,N_4138,N_2804);
or UO_324 (O_324,N_4696,N_3662);
and UO_325 (O_325,N_2607,N_4205);
or UO_326 (O_326,N_2653,N_2694);
nor UO_327 (O_327,N_3874,N_4976);
or UO_328 (O_328,N_4577,N_3818);
nor UO_329 (O_329,N_3341,N_3987);
nand UO_330 (O_330,N_3650,N_3918);
and UO_331 (O_331,N_3953,N_4937);
and UO_332 (O_332,N_3865,N_3102);
or UO_333 (O_333,N_3733,N_4177);
and UO_334 (O_334,N_3162,N_4159);
nor UO_335 (O_335,N_4102,N_4680);
nand UO_336 (O_336,N_4425,N_2689);
and UO_337 (O_337,N_4986,N_4737);
and UO_338 (O_338,N_4120,N_4318);
and UO_339 (O_339,N_2815,N_3222);
and UO_340 (O_340,N_2716,N_4430);
nand UO_341 (O_341,N_4504,N_4091);
or UO_342 (O_342,N_2972,N_3857);
or UO_343 (O_343,N_3920,N_4829);
or UO_344 (O_344,N_4804,N_2852);
and UO_345 (O_345,N_4957,N_3186);
nor UO_346 (O_346,N_4635,N_3769);
or UO_347 (O_347,N_4932,N_2835);
nor UO_348 (O_348,N_4253,N_2832);
and UO_349 (O_349,N_3996,N_2982);
or UO_350 (O_350,N_3007,N_3306);
or UO_351 (O_351,N_3511,N_2914);
or UO_352 (O_352,N_4618,N_3976);
nand UO_353 (O_353,N_3722,N_3409);
and UO_354 (O_354,N_3358,N_3347);
or UO_355 (O_355,N_4210,N_3027);
nand UO_356 (O_356,N_4146,N_3019);
nor UO_357 (O_357,N_3286,N_3195);
or UO_358 (O_358,N_2703,N_3000);
or UO_359 (O_359,N_3932,N_4962);
or UO_360 (O_360,N_4755,N_2671);
and UO_361 (O_361,N_3175,N_4960);
nand UO_362 (O_362,N_2810,N_3123);
or UO_363 (O_363,N_2870,N_2826);
nand UO_364 (O_364,N_4925,N_4266);
or UO_365 (O_365,N_3438,N_3783);
and UO_366 (O_366,N_3296,N_2865);
nor UO_367 (O_367,N_3935,N_4441);
nor UO_368 (O_368,N_3193,N_4689);
nor UO_369 (O_369,N_3532,N_3440);
nand UO_370 (O_370,N_4069,N_3427);
and UO_371 (O_371,N_4612,N_4945);
and UO_372 (O_372,N_3686,N_3204);
nor UO_373 (O_373,N_3110,N_4134);
nor UO_374 (O_374,N_4336,N_2989);
nor UO_375 (O_375,N_3403,N_2561);
or UO_376 (O_376,N_3821,N_4020);
and UO_377 (O_377,N_4284,N_4695);
nand UO_378 (O_378,N_3492,N_3851);
or UO_379 (O_379,N_4292,N_3807);
nand UO_380 (O_380,N_4470,N_2936);
nand UO_381 (O_381,N_3381,N_4357);
nor UO_382 (O_382,N_4388,N_2912);
and UO_383 (O_383,N_4010,N_4510);
and UO_384 (O_384,N_4916,N_3992);
nor UO_385 (O_385,N_4920,N_4623);
nand UO_386 (O_386,N_4730,N_3313);
and UO_387 (O_387,N_3875,N_3472);
nand UO_388 (O_388,N_4643,N_4562);
nand UO_389 (O_389,N_2998,N_4259);
and UO_390 (O_390,N_2981,N_2580);
nor UO_391 (O_391,N_3893,N_4063);
nand UO_392 (O_392,N_4950,N_3673);
nor UO_393 (O_393,N_3219,N_2785);
xnor UO_394 (O_394,N_3940,N_4811);
nand UO_395 (O_395,N_2562,N_3411);
or UO_396 (O_396,N_2859,N_3104);
or UO_397 (O_397,N_3917,N_4075);
nand UO_398 (O_398,N_4705,N_3568);
and UO_399 (O_399,N_4406,N_3753);
and UO_400 (O_400,N_2736,N_3841);
nor UO_401 (O_401,N_2999,N_3288);
nor UO_402 (O_402,N_2806,N_3108);
nor UO_403 (O_403,N_3598,N_3737);
and UO_404 (O_404,N_3091,N_3762);
and UO_405 (O_405,N_2997,N_4805);
or UO_406 (O_406,N_3585,N_2898);
nor UO_407 (O_407,N_3870,N_4711);
nand UO_408 (O_408,N_3203,N_3873);
nor UO_409 (O_409,N_4437,N_3301);
and UO_410 (O_410,N_4473,N_4169);
nor UO_411 (O_411,N_2795,N_4217);
and UO_412 (O_412,N_3350,N_2563);
or UO_413 (O_413,N_4009,N_3558);
and UO_414 (O_414,N_3191,N_4927);
or UO_415 (O_415,N_3063,N_2801);
nor UO_416 (O_416,N_3238,N_3724);
and UO_417 (O_417,N_4144,N_3948);
and UO_418 (O_418,N_4329,N_2807);
nand UO_419 (O_419,N_3963,N_3782);
nand UO_420 (O_420,N_4765,N_3373);
xor UO_421 (O_421,N_4067,N_4786);
and UO_422 (O_422,N_4221,N_3407);
and UO_423 (O_423,N_4251,N_3425);
nand UO_424 (O_424,N_3142,N_3867);
and UO_425 (O_425,N_4260,N_4222);
and UO_426 (O_426,N_3847,N_3490);
nand UO_427 (O_427,N_3190,N_4398);
nor UO_428 (O_428,N_4511,N_4664);
nand UO_429 (O_429,N_4368,N_4729);
nand UO_430 (O_430,N_4539,N_4736);
nor UO_431 (O_431,N_4040,N_4401);
nor UO_432 (O_432,N_2726,N_3481);
or UO_433 (O_433,N_3164,N_3501);
nor UO_434 (O_434,N_2719,N_3479);
nand UO_435 (O_435,N_3484,N_4844);
or UO_436 (O_436,N_4656,N_3575);
nand UO_437 (O_437,N_4734,N_3696);
nor UO_438 (O_438,N_3310,N_4311);
or UO_439 (O_439,N_3693,N_4319);
nand UO_440 (O_440,N_4795,N_4899);
nor UO_441 (O_441,N_2952,N_3197);
nand UO_442 (O_442,N_2829,N_2539);
and UO_443 (O_443,N_2941,N_4417);
and UO_444 (O_444,N_4745,N_4742);
and UO_445 (O_445,N_3221,N_4747);
and UO_446 (O_446,N_2700,N_2691);
nor UO_447 (O_447,N_3058,N_3791);
nand UO_448 (O_448,N_3885,N_4959);
nor UO_449 (O_449,N_3107,N_3336);
nor UO_450 (O_450,N_4647,N_3421);
nor UO_451 (O_451,N_3025,N_2713);
nand UO_452 (O_452,N_4066,N_3509);
and UO_453 (O_453,N_2816,N_4861);
nor UO_454 (O_454,N_3174,N_4171);
or UO_455 (O_455,N_2881,N_3252);
and UO_456 (O_456,N_3946,N_2698);
nor UO_457 (O_457,N_3233,N_3572);
nand UO_458 (O_458,N_3448,N_3919);
or UO_459 (O_459,N_3362,N_4591);
and UO_460 (O_460,N_4039,N_3292);
and UO_461 (O_461,N_2874,N_2959);
or UO_462 (O_462,N_2684,N_3311);
nand UO_463 (O_463,N_2956,N_3830);
nor UO_464 (O_464,N_4405,N_4853);
nand UO_465 (O_465,N_3504,N_4917);
or UO_466 (O_466,N_4082,N_4545);
nand UO_467 (O_467,N_3209,N_4569);
or UO_468 (O_468,N_2811,N_3229);
and UO_469 (O_469,N_3962,N_2712);
nand UO_470 (O_470,N_4326,N_3832);
or UO_471 (O_471,N_4500,N_4451);
nor UO_472 (O_472,N_3593,N_4354);
nand UO_473 (O_473,N_4155,N_3835);
nor UO_474 (O_474,N_4137,N_4349);
or UO_475 (O_475,N_2617,N_3879);
or UO_476 (O_476,N_3167,N_3116);
nand UO_477 (O_477,N_3757,N_3633);
and UO_478 (O_478,N_3075,N_2685);
or UO_479 (O_479,N_2833,N_4741);
or UO_480 (O_480,N_4563,N_3519);
or UO_481 (O_481,N_2558,N_4184);
nand UO_482 (O_482,N_2506,N_2572);
and UO_483 (O_483,N_4914,N_3793);
nand UO_484 (O_484,N_4739,N_4532);
and UO_485 (O_485,N_3775,N_4227);
or UO_486 (O_486,N_4304,N_2911);
nor UO_487 (O_487,N_3340,N_3965);
or UO_488 (O_488,N_2913,N_2696);
nor UO_489 (O_489,N_3958,N_2967);
nand UO_490 (O_490,N_4426,N_3512);
or UO_491 (O_491,N_2618,N_4276);
and UO_492 (O_492,N_3143,N_4862);
nand UO_493 (O_493,N_2553,N_3139);
or UO_494 (O_494,N_4068,N_3601);
nand UO_495 (O_495,N_4059,N_2528);
nand UO_496 (O_496,N_3629,N_2693);
nand UO_497 (O_497,N_3323,N_4749);
or UO_498 (O_498,N_3855,N_3838);
and UO_499 (O_499,N_2525,N_4044);
and UO_500 (O_500,N_3453,N_3463);
and UO_501 (O_501,N_4035,N_3466);
nor UO_502 (O_502,N_3567,N_3819);
nand UO_503 (O_503,N_2520,N_4503);
or UO_504 (O_504,N_3984,N_4172);
nor UO_505 (O_505,N_2654,N_4777);
nor UO_506 (O_506,N_4981,N_4356);
or UO_507 (O_507,N_3437,N_3887);
nand UO_508 (O_508,N_2784,N_4868);
nand UO_509 (O_509,N_4610,N_3899);
nor UO_510 (O_510,N_4469,N_2769);
nand UO_511 (O_511,N_2650,N_4112);
or UO_512 (O_512,N_4293,N_4452);
and UO_513 (O_513,N_4328,N_3624);
and UO_514 (O_514,N_3321,N_3729);
or UO_515 (O_515,N_4062,N_4435);
and UO_516 (O_516,N_4081,N_2546);
and UO_517 (O_517,N_3126,N_3042);
nand UO_518 (O_518,N_3218,N_3388);
or UO_519 (O_519,N_2774,N_4571);
and UO_520 (O_520,N_3738,N_3547);
or UO_521 (O_521,N_3644,N_3237);
nand UO_522 (O_522,N_4199,N_3985);
or UO_523 (O_523,N_2675,N_3052);
or UO_524 (O_524,N_3817,N_4733);
or UO_525 (O_525,N_3065,N_4834);
nand UO_526 (O_526,N_4701,N_4225);
nand UO_527 (O_527,N_3332,N_3964);
nor UO_528 (O_528,N_2848,N_4116);
and UO_529 (O_529,N_2818,N_4800);
nor UO_530 (O_530,N_4521,N_2820);
or UO_531 (O_531,N_3664,N_3916);
and UO_532 (O_532,N_2517,N_4633);
nor UO_533 (O_533,N_2655,N_3363);
nand UO_534 (O_534,N_3454,N_4721);
or UO_535 (O_535,N_2635,N_4988);
and UO_536 (O_536,N_4779,N_4732);
nor UO_537 (O_537,N_4054,N_2614);
nand UO_538 (O_538,N_3978,N_3470);
nand UO_539 (O_539,N_4241,N_2916);
nand UO_540 (O_540,N_4922,N_4351);
and UO_541 (O_541,N_4585,N_2782);
and UO_542 (O_542,N_4570,N_4108);
nand UO_543 (O_543,N_4684,N_3781);
nor UO_544 (O_544,N_4243,N_3316);
nand UO_545 (O_545,N_4846,N_3574);
or UO_546 (O_546,N_4646,N_2789);
and UO_547 (O_547,N_4321,N_4017);
and UO_548 (O_548,N_4949,N_4968);
or UO_549 (O_549,N_3254,N_4572);
and UO_550 (O_550,N_3245,N_2772);
nor UO_551 (O_551,N_3643,N_4587);
nand UO_552 (O_552,N_3763,N_2599);
nand UO_553 (O_553,N_2960,N_2875);
or UO_554 (O_554,N_4176,N_4101);
or UO_555 (O_555,N_4273,N_2864);
nor UO_556 (O_556,N_4433,N_3654);
nor UO_557 (O_557,N_4377,N_4860);
or UO_558 (O_558,N_3322,N_4581);
nand UO_559 (O_559,N_3183,N_3717);
nor UO_560 (O_560,N_4161,N_4617);
nand UO_561 (O_561,N_3721,N_2629);
nor UO_562 (O_562,N_4913,N_3280);
or UO_563 (O_563,N_4796,N_2987);
and UO_564 (O_564,N_2905,N_4662);
and UO_565 (O_565,N_3071,N_3259);
and UO_566 (O_566,N_3442,N_2577);
nor UO_567 (O_567,N_3945,N_2637);
and UO_568 (O_568,N_3284,N_4879);
and UO_569 (O_569,N_4463,N_3177);
xor UO_570 (O_570,N_4127,N_2723);
nand UO_571 (O_571,N_4030,N_4488);
or UO_572 (O_572,N_4071,N_4939);
or UO_573 (O_573,N_2564,N_3619);
xnor UO_574 (O_574,N_4281,N_2896);
and UO_575 (O_575,N_4065,N_4869);
nand UO_576 (O_576,N_4890,N_4690);
nand UO_577 (O_577,N_3517,N_3957);
and UO_578 (O_578,N_2733,N_2659);
nand UO_579 (O_579,N_4901,N_4552);
nand UO_580 (O_580,N_3995,N_3675);
xnor UO_581 (O_581,N_3618,N_4015);
nand UO_582 (O_582,N_3462,N_4604);
and UO_583 (O_583,N_4693,N_4403);
nand UO_584 (O_584,N_2598,N_2873);
nand UO_585 (O_585,N_4337,N_4666);
and UO_586 (O_586,N_4327,N_3432);
nand UO_587 (O_587,N_4691,N_4482);
nand UO_588 (O_588,N_4592,N_3140);
nor UO_589 (O_589,N_3370,N_4444);
or UO_590 (O_590,N_4077,N_3748);
nor UO_591 (O_591,N_2527,N_4106);
and UO_592 (O_592,N_4845,N_4969);
or UO_593 (O_593,N_3404,N_4972);
nand UO_594 (O_594,N_2951,N_2868);
or UO_595 (O_595,N_2612,N_4516);
or UO_596 (O_596,N_4602,N_4880);
nand UO_597 (O_597,N_4507,N_2576);
nand UO_598 (O_598,N_3998,N_3549);
nand UO_599 (O_599,N_4993,N_4709);
nand UO_600 (O_600,N_4051,N_2945);
nand UO_601 (O_601,N_3697,N_2926);
or UO_602 (O_602,N_3707,N_3298);
nor UO_603 (O_603,N_3283,N_2682);
nand UO_604 (O_604,N_2625,N_4419);
xor UO_605 (O_605,N_4219,N_4679);
and UO_606 (O_606,N_3542,N_3825);
nor UO_607 (O_607,N_4538,N_3767);
or UO_608 (O_608,N_4474,N_2856);
nor UO_609 (O_609,N_3630,N_4597);
nand UO_610 (O_610,N_4250,N_3758);
nand UO_611 (O_611,N_3212,N_4218);
nor UO_612 (O_612,N_4279,N_3518);
nand UO_613 (O_613,N_4382,N_3529);
nand UO_614 (O_614,N_2879,N_4931);
and UO_615 (O_615,N_3566,N_4550);
nor UO_616 (O_616,N_2969,N_3491);
and UO_617 (O_617,N_4501,N_3133);
and UO_618 (O_618,N_2950,N_4906);
nor UO_619 (O_619,N_3460,N_4412);
nand UO_620 (O_620,N_3678,N_3672);
nand UO_621 (O_621,N_3088,N_4904);
nor UO_622 (O_622,N_4208,N_4070);
nor UO_623 (O_623,N_4306,N_2773);
nor UO_624 (O_624,N_4390,N_4714);
and UO_625 (O_625,N_3926,N_2924);
or UO_626 (O_626,N_4064,N_3375);
and UO_627 (O_627,N_3514,N_4202);
or UO_628 (O_628,N_3366,N_4847);
or UO_629 (O_629,N_2970,N_3966);
and UO_630 (O_630,N_2523,N_4204);
or UO_631 (O_631,N_4580,N_4985);
and UO_632 (O_632,N_4953,N_4513);
nand UO_633 (O_633,N_4187,N_4584);
nand UO_634 (O_634,N_2866,N_3431);
and UO_635 (O_635,N_4790,N_4145);
nand UO_636 (O_636,N_3941,N_4422);
and UO_637 (O_637,N_3688,N_3806);
or UO_638 (O_638,N_4630,N_4458);
and UO_639 (O_639,N_3525,N_3315);
and UO_640 (O_640,N_2946,N_3612);
or UO_641 (O_641,N_2988,N_4768);
and UO_642 (O_642,N_2927,N_3784);
and UO_643 (O_643,N_3570,N_4991);
or UO_644 (O_644,N_4658,N_4466);
nand UO_645 (O_645,N_4525,N_4089);
or UO_646 (O_646,N_4348,N_4191);
and UO_647 (O_647,N_3872,N_2830);
nor UO_648 (O_648,N_2587,N_3016);
nor UO_649 (O_649,N_3232,N_2533);
and UO_650 (O_650,N_4984,N_4887);
and UO_651 (O_651,N_4057,N_4810);
or UO_652 (O_652,N_4421,N_3364);
nor UO_653 (O_653,N_3584,N_2658);
and UO_654 (O_654,N_3291,N_3342);
nor UO_655 (O_655,N_2813,N_4167);
or UO_656 (O_656,N_4894,N_3766);
or UO_657 (O_657,N_3578,N_3070);
nor UO_658 (O_658,N_2656,N_4196);
nor UO_659 (O_659,N_2825,N_3417);
nor UO_660 (O_660,N_3158,N_4929);
and UO_661 (O_661,N_4838,N_2770);
nor UO_662 (O_662,N_4168,N_4822);
or UO_663 (O_663,N_3081,N_4727);
and UO_664 (O_664,N_4019,N_2591);
and UO_665 (O_665,N_3274,N_3089);
nand UO_666 (O_666,N_3755,N_4517);
and UO_667 (O_667,N_3115,N_4864);
or UO_668 (O_668,N_4541,N_4166);
and UO_669 (O_669,N_3982,N_3268);
and UO_670 (O_670,N_3877,N_4586);
and UO_671 (O_671,N_4885,N_4688);
or UO_672 (O_672,N_2541,N_4700);
and UO_673 (O_673,N_3330,N_4908);
nand UO_674 (O_674,N_3524,N_2746);
nor UO_675 (O_675,N_3494,N_2895);
and UO_676 (O_676,N_2780,N_3652);
nor UO_677 (O_677,N_2519,N_4206);
nor UO_678 (O_678,N_3062,N_2548);
or UO_679 (O_679,N_3777,N_4843);
and UO_680 (O_680,N_4527,N_4181);
and UO_681 (O_681,N_2968,N_3674);
and UO_682 (O_682,N_4898,N_2915);
and UO_683 (O_683,N_3770,N_3003);
or UO_684 (O_684,N_3527,N_4614);
and UO_685 (O_685,N_4157,N_4142);
or UO_686 (O_686,N_2609,N_4831);
and UO_687 (O_687,N_4613,N_2631);
nand UO_688 (O_688,N_3441,N_3787);
nor UO_689 (O_689,N_3670,N_3418);
xor UO_690 (O_690,N_3365,N_3230);
or UO_691 (O_691,N_3009,N_3896);
and UO_692 (O_692,N_4263,N_3901);
and UO_693 (O_693,N_3506,N_4400);
and UO_694 (O_694,N_3754,N_4657);
nand UO_695 (O_695,N_2802,N_4295);
or UO_696 (O_696,N_3683,N_4849);
nor UO_697 (O_697,N_3314,N_2500);
or UO_698 (O_698,N_4944,N_4086);
nor UO_699 (O_699,N_4756,N_4325);
nand UO_700 (O_700,N_4025,N_4224);
nand UO_701 (O_701,N_2702,N_4491);
and UO_702 (O_702,N_4835,N_4233);
or UO_703 (O_703,N_2666,N_3538);
and UO_704 (O_704,N_4546,N_4162);
and UO_705 (O_705,N_4649,N_4346);
nand UO_706 (O_706,N_4007,N_4746);
or UO_707 (O_707,N_3582,N_2840);
nor UO_708 (O_708,N_4535,N_3111);
and UO_709 (O_709,N_3742,N_3352);
or UO_710 (O_710,N_2762,N_3256);
or UO_711 (O_711,N_3086,N_2796);
nand UO_712 (O_712,N_3357,N_4514);
nand UO_713 (O_713,N_4903,N_3201);
nor UO_714 (O_714,N_3701,N_4345);
or UO_715 (O_715,N_4085,N_3682);
nand UO_716 (O_716,N_4034,N_4882);
or UO_717 (O_717,N_4668,N_3100);
and UO_718 (O_718,N_3510,N_4808);
or UO_719 (O_719,N_4710,N_4743);
and UO_720 (O_720,N_2678,N_3552);
or UO_721 (O_721,N_3374,N_4687);
and UO_722 (O_722,N_3130,N_4990);
nand UO_723 (O_723,N_2554,N_4305);
nand UO_724 (O_724,N_3497,N_3129);
and UO_725 (O_725,N_4579,N_3756);
and UO_726 (O_726,N_3092,N_3337);
or UO_727 (O_727,N_4440,N_3046);
nand UO_728 (O_728,N_3423,N_4699);
nor UO_729 (O_729,N_4193,N_4026);
nor UO_730 (O_730,N_3200,N_4678);
or UO_731 (O_731,N_4826,N_4122);
xor UO_732 (O_732,N_3180,N_4014);
or UO_733 (O_733,N_4629,N_3061);
nor UO_734 (O_734,N_3993,N_2742);
nand UO_735 (O_735,N_3505,N_4360);
nand UO_736 (O_736,N_3234,N_4013);
or UO_737 (O_737,N_3489,N_3559);
and UO_738 (O_738,N_3285,N_3276);
or UO_739 (O_739,N_3933,N_4343);
nand UO_740 (O_740,N_4397,N_3487);
and UO_741 (O_741,N_3636,N_2524);
nand UO_742 (O_742,N_3397,N_2585);
nor UO_743 (O_743,N_2961,N_3319);
nor UO_744 (O_744,N_2948,N_2721);
or UO_745 (O_745,N_3594,N_3271);
nand UO_746 (O_746,N_3581,N_2990);
or UO_747 (O_747,N_2544,N_3730);
nand UO_748 (O_748,N_2902,N_4093);
or UO_749 (O_749,N_4189,N_4718);
nor UO_750 (O_750,N_3137,N_3907);
or UO_751 (O_751,N_3603,N_3970);
nand UO_752 (O_752,N_3607,N_2992);
nor UO_753 (O_753,N_4938,N_3727);
nand UO_754 (O_754,N_4456,N_2582);
nand UO_755 (O_755,N_3273,N_3171);
and UO_756 (O_756,N_4045,N_4987);
and UO_757 (O_757,N_3049,N_4269);
and UO_758 (O_758,N_4074,N_3228);
or UO_759 (O_759,N_4139,N_4073);
nor UO_760 (O_760,N_4566,N_2504);
nor UO_761 (O_761,N_3398,N_2897);
nor UO_762 (O_762,N_3308,N_3250);
xnor UO_763 (O_763,N_3528,N_3371);
nor UO_764 (O_764,N_4958,N_3471);
nand UO_765 (O_765,N_4407,N_3196);
nand UO_766 (O_766,N_4160,N_3596);
nor UO_767 (O_767,N_3198,N_4576);
nand UO_768 (O_768,N_3882,N_4048);
nand UO_769 (O_769,N_4738,N_3815);
nand UO_770 (O_770,N_3101,N_3103);
nor UO_771 (O_771,N_3565,N_4776);
and UO_772 (O_772,N_3833,N_2759);
or UO_773 (O_773,N_2738,N_3145);
nand UO_774 (O_774,N_2624,N_3994);
nor UO_775 (O_775,N_4448,N_3659);
and UO_776 (O_776,N_4653,N_2790);
nor UO_777 (O_777,N_3546,N_4022);
nor UO_778 (O_778,N_2857,N_3355);
nand UO_779 (O_779,N_3600,N_4971);
nor UO_780 (O_780,N_3023,N_4748);
or UO_781 (O_781,N_4508,N_4460);
or UO_782 (O_782,N_2556,N_2657);
nand UO_783 (O_783,N_4951,N_4803);
or UO_784 (O_784,N_4815,N_4424);
nand UO_785 (O_785,N_3223,N_3602);
or UO_786 (O_786,N_4919,N_2547);
or UO_787 (O_787,N_2680,N_3771);
nand UO_788 (O_788,N_2549,N_3959);
nor UO_789 (O_789,N_3189,N_2581);
or UO_790 (O_790,N_3942,N_4216);
nor UO_791 (O_791,N_4104,N_2667);
and UO_792 (O_792,N_4628,N_3051);
nand UO_793 (O_793,N_2899,N_3588);
nand UO_794 (O_794,N_4634,N_2860);
or UO_795 (O_795,N_3056,N_3545);
or UO_796 (O_796,N_3900,N_4480);
nand UO_797 (O_797,N_4841,N_2876);
xnor UO_798 (O_798,N_3702,N_3326);
nor UO_799 (O_799,N_4277,N_4816);
nor UO_800 (O_800,N_3073,N_3012);
nand UO_801 (O_801,N_4639,N_3434);
or UO_802 (O_802,N_4726,N_2824);
or UO_803 (O_803,N_3192,N_3816);
nor UO_804 (O_804,N_3522,N_4379);
and UO_805 (O_805,N_4600,N_3069);
or UO_806 (O_806,N_4378,N_4320);
nand UO_807 (O_807,N_4363,N_4677);
nor UO_808 (O_808,N_2756,N_3638);
nor UO_809 (O_809,N_3599,N_3034);
nor UO_810 (O_810,N_4008,N_4759);
and UO_811 (O_811,N_4294,N_4203);
nor UO_812 (O_812,N_4449,N_2677);
xor UO_813 (O_813,N_2514,N_4851);
nor UO_814 (O_814,N_3343,N_3554);
nor UO_815 (O_815,N_4589,N_3220);
nand UO_816 (O_816,N_2516,N_4648);
or UO_817 (O_817,N_4715,N_3740);
and UO_818 (O_818,N_3663,N_4704);
or UO_819 (O_819,N_4418,N_3128);
nand UO_820 (O_820,N_2799,N_2537);
nand UO_821 (O_821,N_4606,N_3842);
and UO_822 (O_822,N_3138,N_2722);
or UO_823 (O_823,N_2538,N_4967);
and UO_824 (O_824,N_4090,N_4353);
nor UO_825 (O_825,N_4565,N_3473);
nor UO_826 (O_826,N_3531,N_4339);
nand UO_827 (O_827,N_2503,N_4154);
nor UO_828 (O_828,N_3211,N_4520);
and UO_829 (O_829,N_2996,N_3047);
nand UO_830 (O_830,N_4593,N_2639);
nor UO_831 (O_831,N_3983,N_4334);
nor UO_832 (O_832,N_4439,N_3068);
nand UO_833 (O_833,N_2709,N_2717);
and UO_834 (O_834,N_2767,N_3805);
and UO_835 (O_835,N_4564,N_2922);
nor UO_836 (O_836,N_4232,N_3616);
and UO_837 (O_837,N_4370,N_4170);
or UO_838 (O_838,N_4257,N_4797);
and UO_839 (O_839,N_3010,N_4195);
or UO_840 (O_840,N_3261,N_3669);
or UO_841 (O_841,N_3022,N_3150);
nor UO_842 (O_842,N_4848,N_4052);
nor UO_843 (O_843,N_3967,N_4111);
and UO_844 (O_844,N_2711,N_3496);
nand UO_845 (O_845,N_4350,N_2521);
and UO_846 (O_846,N_4242,N_4267);
or UO_847 (O_847,N_4033,N_2615);
or UO_848 (O_848,N_3093,N_2660);
nor UO_849 (O_849,N_3744,N_2930);
and UO_850 (O_850,N_4256,N_2531);
nor UO_851 (O_851,N_3954,N_2939);
and UO_852 (O_852,N_2535,N_3207);
nor UO_853 (O_853,N_3041,N_4239);
nand UO_854 (O_854,N_3938,N_4989);
or UO_855 (O_855,N_3723,N_3853);
or UO_856 (O_856,N_3153,N_2697);
and UO_857 (O_857,N_4943,N_3136);
or UO_858 (O_858,N_4414,N_4567);
nand UO_859 (O_859,N_3028,N_3736);
and UO_860 (O_860,N_3199,N_2735);
or UO_861 (O_861,N_3677,N_4923);
nand UO_862 (O_862,N_2891,N_3152);
xor UO_863 (O_863,N_2699,N_4084);
or UO_864 (O_864,N_4791,N_2593);
and UO_865 (O_865,N_3990,N_2552);
and UO_866 (O_866,N_2986,N_4774);
or UO_867 (O_867,N_3991,N_3956);
xor UO_868 (O_868,N_3242,N_4049);
nand UO_869 (O_869,N_3776,N_3812);
or UO_870 (O_870,N_3182,N_3053);
or UO_871 (O_871,N_3890,N_4393);
and UO_872 (O_872,N_4806,N_3952);
nand UO_873 (O_873,N_3225,N_3476);
or UO_874 (O_874,N_2745,N_2933);
nor UO_875 (O_875,N_4395,N_4683);
nand UO_876 (O_876,N_4896,N_4528);
nand UO_877 (O_877,N_4706,N_3208);
and UO_878 (O_878,N_3974,N_4760);
nor UO_879 (O_879,N_3176,N_4275);
and UO_880 (O_880,N_3396,N_3667);
nand UO_881 (O_881,N_2983,N_4215);
and UO_882 (O_882,N_3808,N_4556);
xnor UO_883 (O_883,N_3883,N_4396);
or UO_884 (O_884,N_2844,N_4450);
and UO_885 (O_885,N_4415,N_3451);
nor UO_886 (O_886,N_4954,N_2560);
or UO_887 (O_887,N_3429,N_4238);
nand UO_888 (O_888,N_2621,N_3590);
or UO_889 (O_889,N_4476,N_4999);
and UO_890 (O_890,N_4180,N_4909);
and UO_891 (O_891,N_2565,N_4966);
nand UO_892 (O_892,N_2739,N_4789);
and UO_893 (O_893,N_3475,N_3275);
nand UO_894 (O_894,N_4766,N_3084);
nand UO_895 (O_895,N_4830,N_3436);
nand UO_896 (O_896,N_4021,N_4910);
nand UO_897 (O_897,N_4046,N_2850);
nor UO_898 (O_898,N_4583,N_4763);
nand UO_899 (O_899,N_2978,N_3911);
or UO_900 (O_900,N_4559,N_2632);
nand UO_901 (O_901,N_3450,N_2955);
or UO_902 (O_902,N_3231,N_3378);
and UO_903 (O_903,N_3797,N_4299);
nand UO_904 (O_904,N_3135,N_4992);
nand UO_905 (O_905,N_4975,N_3279);
nand UO_906 (O_906,N_2880,N_3458);
nand UO_907 (O_907,N_4432,N_2526);
nand UO_908 (O_908,N_4413,N_3627);
and UO_909 (O_909,N_3267,N_3328);
nor UO_910 (O_910,N_4489,N_4355);
and UO_911 (O_911,N_2579,N_3015);
or UO_912 (O_912,N_4809,N_2904);
and UO_913 (O_913,N_2522,N_3376);
nand UO_914 (O_914,N_3837,N_2643);
nor UO_915 (O_915,N_3044,N_3335);
or UO_916 (O_916,N_4454,N_3109);
or UO_917 (O_917,N_4930,N_3854);
nor UO_918 (O_918,N_3955,N_4588);
nand UO_919 (O_919,N_3131,N_4787);
or UO_920 (O_920,N_2633,N_2771);
nor UO_921 (O_921,N_2600,N_4724);
nand UO_922 (O_922,N_3640,N_4207);
nand UO_923 (O_923,N_4248,N_3986);
nor UO_924 (O_924,N_4047,N_2530);
nor UO_925 (O_925,N_4769,N_4004);
or UO_926 (O_926,N_2775,N_3889);
or UO_927 (O_927,N_3943,N_4828);
nor UO_928 (O_928,N_4002,N_3657);
nand UO_929 (O_929,N_3348,N_4254);
or UO_930 (O_930,N_2792,N_3083);
nand UO_931 (O_931,N_2888,N_3820);
nor UO_932 (O_932,N_4190,N_2937);
nand UO_933 (O_933,N_2518,N_3809);
nand UO_934 (O_934,N_3713,N_2701);
nor UO_935 (O_935,N_3464,N_2652);
and UO_936 (O_936,N_2965,N_3503);
and UO_937 (O_937,N_4148,N_3631);
and UO_938 (O_938,N_3029,N_2729);
or UO_939 (O_939,N_3033,N_2623);
nand UO_940 (O_940,N_4551,N_4445);
and UO_941 (O_941,N_4096,N_2862);
nor UO_942 (O_942,N_4858,N_3227);
nor UO_943 (O_943,N_4344,N_3312);
and UO_944 (O_944,N_3318,N_3064);
nor UO_945 (O_945,N_2648,N_3792);
nor UO_946 (O_946,N_4291,N_2800);
and UO_947 (O_947,N_3910,N_4912);
nor UO_948 (O_948,N_2649,N_4270);
and UO_949 (O_949,N_3367,N_4050);
or UO_950 (O_950,N_3614,N_4366);
and UO_951 (O_951,N_2574,N_3561);
nor UO_952 (O_952,N_3718,N_4411);
and UO_953 (O_953,N_3356,N_3486);
nor UO_954 (O_954,N_2980,N_2670);
nand UO_955 (O_955,N_3391,N_4201);
nor UO_956 (O_956,N_3826,N_4472);
nor UO_957 (O_957,N_2661,N_4652);
or UO_958 (O_958,N_4374,N_3779);
or UO_959 (O_959,N_3118,N_4728);
nor UO_960 (O_960,N_4518,N_3828);
and UO_961 (O_961,N_3300,N_2507);
nand UO_962 (O_962,N_4200,N_3708);
and UO_963 (O_963,N_4673,N_4151);
nor UO_964 (O_964,N_2836,N_3181);
and UO_965 (O_965,N_3331,N_2928);
nand UO_966 (O_966,N_2734,N_4863);
or UO_967 (O_967,N_2877,N_4043);
and UO_968 (O_968,N_3699,N_2991);
nor UO_969 (O_969,N_4764,N_2731);
or UO_970 (O_970,N_3281,N_3405);
and UO_971 (O_971,N_4443,N_2822);
or UO_972 (O_972,N_4369,N_4540);
and UO_973 (O_973,N_2730,N_4226);
nand UO_974 (O_974,N_3345,N_2636);
nor UO_975 (O_975,N_3658,N_3856);
or UO_976 (O_976,N_4716,N_3858);
nand UO_977 (O_977,N_3165,N_4236);
or UO_978 (O_978,N_2540,N_3530);
or UO_979 (O_979,N_3468,N_3888);
and UO_980 (O_980,N_3604,N_4174);
and UO_981 (O_981,N_3666,N_3457);
and UO_982 (O_982,N_4940,N_4006);
or UO_983 (O_983,N_2672,N_2962);
and UO_984 (O_984,N_2622,N_2909);
and UO_985 (O_985,N_3687,N_4964);
or UO_986 (O_986,N_2640,N_3430);
nor UO_987 (O_987,N_4135,N_2995);
nand UO_988 (O_988,N_4003,N_3831);
and UO_989 (O_989,N_3648,N_4459);
and UO_990 (O_990,N_4644,N_3829);
and UO_991 (O_991,N_3013,N_3449);
and UO_992 (O_992,N_3217,N_4681);
nand UO_993 (O_993,N_3720,N_2993);
and UO_994 (O_994,N_4875,N_4058);
nor UO_995 (O_995,N_2957,N_3871);
nor UO_996 (O_996,N_4506,N_2741);
nand UO_997 (O_997,N_4526,N_3050);
nand UO_998 (O_998,N_4153,N_3608);
nor UO_999 (O_999,N_3161,N_3906);
endmodule