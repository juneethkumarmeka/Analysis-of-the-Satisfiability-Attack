module basic_500_3000_500_30_levels_5xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nor U0 (N_0,In_351,In_197);
xor U1 (N_1,In_433,In_283);
xnor U2 (N_2,In_342,In_336);
nor U3 (N_3,In_109,In_408);
and U4 (N_4,In_14,In_193);
nor U5 (N_5,In_353,In_117);
and U6 (N_6,In_455,In_365);
or U7 (N_7,In_491,In_40);
xor U8 (N_8,In_397,In_126);
nor U9 (N_9,In_371,In_121);
or U10 (N_10,In_84,In_360);
nor U11 (N_11,In_111,In_88);
or U12 (N_12,In_315,In_154);
or U13 (N_13,In_79,In_256);
nor U14 (N_14,In_431,In_392);
nor U15 (N_15,In_273,In_429);
xnor U16 (N_16,In_310,In_235);
nor U17 (N_17,In_391,In_161);
or U18 (N_18,In_114,In_214);
nand U19 (N_19,In_434,In_326);
and U20 (N_20,In_185,In_44);
nand U21 (N_21,In_382,In_258);
nor U22 (N_22,In_159,In_261);
or U23 (N_23,In_203,In_38);
nor U24 (N_24,In_291,In_296);
xor U25 (N_25,In_179,In_215);
nand U26 (N_26,In_267,In_401);
or U27 (N_27,In_212,In_217);
nor U28 (N_28,In_21,In_137);
nand U29 (N_29,In_37,In_142);
or U30 (N_30,In_430,In_294);
nor U31 (N_31,In_210,In_231);
nor U32 (N_32,In_356,In_373);
nand U33 (N_33,In_198,In_486);
nor U34 (N_34,In_441,In_64);
nor U35 (N_35,In_196,In_475);
and U36 (N_36,In_304,In_272);
and U37 (N_37,In_66,In_48);
or U38 (N_38,In_54,In_136);
nor U39 (N_39,In_411,In_262);
nor U40 (N_40,In_384,In_366);
or U41 (N_41,In_276,In_87);
nand U42 (N_42,In_421,In_15);
nand U43 (N_43,In_130,In_266);
nand U44 (N_44,In_308,In_181);
and U45 (N_45,In_333,In_167);
and U46 (N_46,In_337,In_419);
and U47 (N_47,In_359,In_160);
nor U48 (N_48,In_22,In_479);
or U49 (N_49,In_427,In_480);
and U50 (N_50,In_473,In_403);
nand U51 (N_51,In_76,In_13);
nand U52 (N_52,In_158,In_254);
and U53 (N_53,In_28,In_307);
or U54 (N_54,In_277,In_274);
nand U55 (N_55,In_335,In_106);
or U56 (N_56,In_334,In_200);
xor U57 (N_57,In_9,In_83);
nor U58 (N_58,In_318,In_343);
nor U59 (N_59,In_407,In_23);
or U60 (N_60,In_115,In_164);
nand U61 (N_61,In_497,In_388);
nor U62 (N_62,In_244,In_8);
or U63 (N_63,In_281,In_459);
or U64 (N_64,In_47,In_317);
xor U65 (N_65,In_338,In_144);
nand U66 (N_66,In_285,In_180);
nor U67 (N_67,In_102,In_119);
nand U68 (N_68,In_270,In_49);
xor U69 (N_69,In_293,In_331);
and U70 (N_70,In_127,In_29);
or U71 (N_71,In_349,In_344);
or U72 (N_72,In_11,In_314);
nor U73 (N_73,In_268,In_496);
xnor U74 (N_74,In_375,In_264);
and U75 (N_75,In_25,In_394);
nand U76 (N_76,In_406,In_70);
nor U77 (N_77,In_282,In_1);
and U78 (N_78,In_192,In_236);
and U79 (N_79,In_201,In_169);
and U80 (N_80,In_216,In_229);
nor U81 (N_81,In_374,In_279);
xnor U82 (N_82,In_494,In_362);
and U83 (N_83,In_461,In_489);
and U84 (N_84,In_250,In_146);
and U85 (N_85,In_2,In_467);
nor U86 (N_86,In_10,In_292);
and U87 (N_87,In_183,In_423);
and U88 (N_88,In_457,In_148);
and U89 (N_89,In_468,In_35);
nor U90 (N_90,In_470,In_389);
nand U91 (N_91,In_417,In_447);
nand U92 (N_92,In_445,In_393);
xor U93 (N_93,In_443,In_369);
or U94 (N_94,In_100,In_5);
nand U95 (N_95,In_298,In_206);
nand U96 (N_96,In_448,In_381);
nand U97 (N_97,In_499,In_379);
nand U98 (N_98,In_249,In_442);
xor U99 (N_99,In_347,In_73);
and U100 (N_100,In_402,In_472);
and U101 (N_101,In_484,In_6);
nand U102 (N_102,In_425,N_80);
nand U103 (N_103,In_46,In_147);
nand U104 (N_104,N_8,In_17);
nor U105 (N_105,In_124,In_450);
nor U106 (N_106,In_99,In_253);
nor U107 (N_107,In_350,N_87);
nand U108 (N_108,N_39,In_45);
nand U109 (N_109,In_354,In_116);
nand U110 (N_110,N_41,N_77);
nand U111 (N_111,In_151,N_93);
xnor U112 (N_112,N_44,In_20);
xor U113 (N_113,In_345,In_77);
nor U114 (N_114,N_12,In_0);
nor U115 (N_115,In_129,In_284);
or U116 (N_116,In_145,N_49);
nand U117 (N_117,N_15,N_35);
nand U118 (N_118,In_251,In_483);
and U119 (N_119,In_263,In_16);
or U120 (N_120,In_444,In_222);
nor U121 (N_121,N_85,In_439);
and U122 (N_122,In_81,In_172);
and U123 (N_123,In_39,In_245);
nor U124 (N_124,In_413,In_252);
and U125 (N_125,In_233,In_139);
or U126 (N_126,In_396,In_280);
and U127 (N_127,In_476,N_86);
xnor U128 (N_128,In_239,In_259);
xnor U129 (N_129,N_27,In_466);
and U130 (N_130,N_52,N_58);
nand U131 (N_131,In_61,N_32);
or U132 (N_132,In_395,In_24);
xnor U133 (N_133,In_68,In_464);
nor U134 (N_134,In_125,In_177);
and U135 (N_135,In_241,N_38);
nand U136 (N_136,N_59,In_4);
nor U137 (N_137,In_386,In_316);
nor U138 (N_138,N_17,In_12);
nor U139 (N_139,In_205,In_477);
and U140 (N_140,In_226,N_54);
or U141 (N_141,In_246,N_30);
and U142 (N_142,In_34,N_74);
xor U143 (N_143,In_238,In_438);
and U144 (N_144,N_22,In_352);
or U145 (N_145,In_120,N_29);
nand U146 (N_146,In_204,In_138);
or U147 (N_147,In_387,In_93);
or U148 (N_148,In_320,In_420);
xor U149 (N_149,N_28,In_287);
nand U150 (N_150,In_319,N_94);
and U151 (N_151,In_299,In_175);
nor U152 (N_152,N_51,In_78);
nor U153 (N_153,N_10,N_83);
nor U154 (N_154,N_14,In_474);
or U155 (N_155,In_110,In_227);
xor U156 (N_156,In_398,In_96);
nor U157 (N_157,N_67,In_437);
nor U158 (N_158,In_301,In_134);
and U159 (N_159,In_358,In_458);
nand U160 (N_160,N_61,In_415);
nor U161 (N_161,In_303,In_67);
nor U162 (N_162,N_60,In_103);
nor U163 (N_163,In_410,In_348);
nand U164 (N_164,In_242,In_456);
nor U165 (N_165,In_481,In_55);
nand U166 (N_166,In_323,In_27);
nor U167 (N_167,In_188,In_52);
or U168 (N_168,In_289,In_168);
nand U169 (N_169,In_328,N_46);
nor U170 (N_170,In_207,In_43);
nor U171 (N_171,In_327,N_42);
or U172 (N_172,N_1,N_40);
or U173 (N_173,N_36,In_133);
nor U174 (N_174,N_16,In_364);
and U175 (N_175,N_99,N_79);
and U176 (N_176,In_329,N_23);
nor U177 (N_177,In_313,N_73);
nor U178 (N_178,In_75,In_140);
or U179 (N_179,In_191,In_59);
nor U180 (N_180,In_141,In_19);
and U181 (N_181,In_53,N_50);
nor U182 (N_182,In_400,N_31);
nand U183 (N_183,In_265,In_302);
and U184 (N_184,In_156,N_37);
or U185 (N_185,In_454,In_367);
or U186 (N_186,In_300,N_11);
nand U187 (N_187,N_19,In_412);
and U188 (N_188,N_2,In_98);
nor U189 (N_189,N_57,N_84);
nor U190 (N_190,In_428,In_426);
and U191 (N_191,In_132,In_324);
or U192 (N_192,In_86,In_286);
xor U193 (N_193,In_385,In_153);
or U194 (N_194,In_432,In_460);
and U195 (N_195,In_436,N_82);
nand U196 (N_196,In_176,N_97);
and U197 (N_197,In_97,In_150);
nor U198 (N_198,In_162,In_165);
and U199 (N_199,In_213,In_449);
nor U200 (N_200,N_168,N_163);
and U201 (N_201,In_218,N_156);
and U202 (N_202,In_56,In_240);
or U203 (N_203,In_340,N_81);
nor U204 (N_204,In_311,N_110);
nor U205 (N_205,In_248,N_189);
xnor U206 (N_206,In_332,In_190);
nand U207 (N_207,N_145,In_143);
or U208 (N_208,In_199,N_68);
or U209 (N_209,In_361,In_257);
nand U210 (N_210,In_495,N_106);
nand U211 (N_211,In_424,In_186);
or U212 (N_212,In_187,In_422);
and U213 (N_213,In_123,In_390);
nor U214 (N_214,In_65,In_30);
and U215 (N_215,N_198,N_177);
nor U216 (N_216,N_65,N_88);
and U217 (N_217,N_185,In_306);
or U218 (N_218,In_219,In_74);
nand U219 (N_219,N_147,N_64);
nor U220 (N_220,N_132,N_193);
nand U221 (N_221,In_462,N_4);
nand U222 (N_222,In_26,N_9);
nand U223 (N_223,In_368,In_357);
or U224 (N_224,N_192,N_183);
or U225 (N_225,In_234,N_191);
or U226 (N_226,In_451,N_160);
xnor U227 (N_227,N_184,In_339);
or U228 (N_228,N_18,In_69);
nand U229 (N_229,In_269,In_91);
or U230 (N_230,N_96,N_111);
or U231 (N_231,N_91,In_108);
nor U232 (N_232,In_488,N_45);
and U233 (N_233,N_175,N_125);
or U234 (N_234,N_24,In_131);
and U235 (N_235,In_309,N_25);
nand U236 (N_236,N_56,N_78);
nor U237 (N_237,In_409,N_70);
nand U238 (N_238,N_104,N_171);
or U239 (N_239,In_405,In_290);
or U240 (N_240,N_63,In_255);
nand U241 (N_241,In_112,In_60);
nor U242 (N_242,In_418,N_119);
and U243 (N_243,N_149,N_0);
nor U244 (N_244,N_142,N_172);
nor U245 (N_245,In_225,In_72);
nor U246 (N_246,N_196,N_166);
and U247 (N_247,N_101,N_158);
or U248 (N_248,In_128,In_105);
nand U249 (N_249,N_116,In_446);
nand U250 (N_250,N_98,In_101);
or U251 (N_251,N_187,In_493);
and U252 (N_252,In_152,In_482);
or U253 (N_253,N_162,N_114);
and U254 (N_254,In_7,N_126);
xnor U255 (N_255,In_211,In_380);
nor U256 (N_256,In_195,N_71);
or U257 (N_257,N_33,N_130);
and U258 (N_258,N_20,In_247);
nor U259 (N_259,N_7,In_471);
and U260 (N_260,N_136,In_465);
nand U261 (N_261,In_295,N_143);
or U262 (N_262,N_154,N_146);
nor U263 (N_263,In_50,In_51);
nand U264 (N_264,In_485,In_122);
and U265 (N_265,In_104,In_82);
nand U266 (N_266,N_167,In_221);
xor U267 (N_267,N_108,N_161);
nand U268 (N_268,In_224,N_199);
xor U269 (N_269,N_95,In_487);
and U270 (N_270,In_492,In_92);
nand U271 (N_271,In_220,N_118);
nand U272 (N_272,In_32,N_186);
nor U273 (N_273,In_41,N_197);
or U274 (N_274,N_151,In_202);
or U275 (N_275,N_115,N_69);
nand U276 (N_276,N_34,In_3);
nand U277 (N_277,N_131,N_157);
nor U278 (N_278,N_159,N_140);
or U279 (N_279,N_5,In_208);
and U280 (N_280,In_404,In_435);
nand U281 (N_281,N_90,In_166);
nor U282 (N_282,N_195,N_122);
nor U283 (N_283,N_66,In_57);
nand U284 (N_284,N_165,In_33);
and U285 (N_285,N_141,N_48);
nand U286 (N_286,In_288,In_453);
nand U287 (N_287,In_377,In_271);
and U288 (N_288,In_376,In_414);
or U289 (N_289,In_230,In_341);
or U290 (N_290,N_181,In_62);
nor U291 (N_291,In_71,In_278);
nor U292 (N_292,N_107,In_440);
and U293 (N_293,In_149,N_62);
nor U294 (N_294,N_194,In_63);
nand U295 (N_295,In_95,In_243);
and U296 (N_296,In_42,In_498);
nor U297 (N_297,N_137,N_113);
nor U298 (N_298,In_330,In_194);
and U299 (N_299,N_173,In_469);
nor U300 (N_300,N_120,N_244);
and U301 (N_301,N_55,N_89);
nand U302 (N_302,N_260,N_286);
xor U303 (N_303,N_239,N_224);
or U304 (N_304,N_117,N_238);
nand U305 (N_305,N_208,N_263);
and U306 (N_306,N_225,N_294);
nand U307 (N_307,N_215,N_76);
and U308 (N_308,In_135,N_170);
and U309 (N_309,In_346,N_228);
nor U310 (N_310,N_169,N_237);
and U311 (N_311,N_258,In_452);
or U312 (N_312,N_284,N_297);
nor U313 (N_313,N_234,In_275);
or U314 (N_314,In_155,N_144);
nand U315 (N_315,In_170,N_291);
nor U316 (N_316,N_233,N_289);
xor U317 (N_317,In_383,N_152);
or U318 (N_318,N_75,N_47);
nor U319 (N_319,N_292,In_399);
xor U320 (N_320,N_112,In_228);
and U321 (N_321,N_241,N_226);
nand U322 (N_322,N_243,In_85);
nor U323 (N_323,N_264,N_21);
or U324 (N_324,N_188,N_26);
and U325 (N_325,In_378,N_133);
xor U326 (N_326,N_235,N_123);
nor U327 (N_327,N_281,N_43);
or U328 (N_328,N_287,In_163);
and U329 (N_329,N_295,N_210);
nor U330 (N_330,N_176,N_273);
nand U331 (N_331,N_53,N_13);
nand U332 (N_332,N_293,N_129);
or U333 (N_333,N_102,N_259);
nand U334 (N_334,N_275,N_298);
nor U335 (N_335,N_250,N_271);
nor U336 (N_336,N_203,In_321);
nor U337 (N_337,N_282,N_296);
nor U338 (N_338,N_214,In_209);
and U339 (N_339,N_249,N_229);
or U340 (N_340,N_201,In_113);
xnor U341 (N_341,N_211,N_262);
nor U342 (N_342,N_138,N_242);
nor U343 (N_343,In_232,In_18);
and U344 (N_344,N_231,In_322);
nor U345 (N_345,N_267,In_478);
xnor U346 (N_346,N_155,N_236);
or U347 (N_347,N_190,N_272);
or U348 (N_348,N_212,N_248);
and U349 (N_349,N_204,N_6);
nor U350 (N_350,In_312,N_3);
nor U351 (N_351,N_202,N_92);
xnor U352 (N_352,N_139,In_370);
or U353 (N_353,N_164,In_90);
and U354 (N_354,N_213,N_148);
nor U355 (N_355,N_180,In_325);
nor U356 (N_356,N_299,In_58);
or U357 (N_357,N_230,N_205);
and U358 (N_358,N_288,In_157);
or U359 (N_359,In_305,In_416);
nand U360 (N_360,N_251,In_490);
nor U361 (N_361,N_255,In_463);
nand U362 (N_362,N_207,N_252);
and U363 (N_363,In_178,N_240);
or U364 (N_364,N_153,N_109);
and U365 (N_365,N_206,N_223);
or U366 (N_366,In_363,N_216);
or U367 (N_367,N_269,N_105);
nand U368 (N_368,N_257,N_276);
or U369 (N_369,N_279,N_182);
nor U370 (N_370,In_118,N_134);
or U371 (N_371,N_103,N_179);
and U372 (N_372,N_72,N_174);
nand U373 (N_373,N_285,N_135);
nand U374 (N_374,N_217,N_222);
nor U375 (N_375,N_127,In_189);
or U376 (N_376,N_218,In_297);
xor U377 (N_377,In_237,In_372);
or U378 (N_378,N_278,N_178);
and U379 (N_379,N_247,In_171);
or U380 (N_380,In_107,N_254);
nand U381 (N_381,N_219,N_274);
nor U382 (N_382,N_227,In_173);
xnor U383 (N_383,N_150,N_220);
nand U384 (N_384,N_253,N_268);
nand U385 (N_385,N_221,N_209);
nor U386 (N_386,In_260,In_36);
xnor U387 (N_387,In_184,In_174);
nand U388 (N_388,N_232,N_270);
or U389 (N_389,N_128,N_256);
or U390 (N_390,N_283,In_355);
nor U391 (N_391,N_121,In_94);
nand U392 (N_392,N_246,In_89);
xnor U393 (N_393,N_290,N_277);
xnor U394 (N_394,In_182,N_265);
or U395 (N_395,In_31,N_200);
nor U396 (N_396,N_124,N_245);
or U397 (N_397,In_80,N_261);
and U398 (N_398,N_280,In_223);
or U399 (N_399,N_266,N_100);
nand U400 (N_400,N_333,N_360);
nand U401 (N_401,N_373,N_363);
and U402 (N_402,N_351,N_384);
nand U403 (N_403,N_327,N_346);
nand U404 (N_404,N_352,N_397);
or U405 (N_405,N_338,N_372);
or U406 (N_406,N_393,N_348);
nor U407 (N_407,N_362,N_356);
xor U408 (N_408,N_378,N_330);
and U409 (N_409,N_312,N_365);
xnor U410 (N_410,N_367,N_387);
or U411 (N_411,N_361,N_334);
nand U412 (N_412,N_305,N_308);
and U413 (N_413,N_355,N_339);
nor U414 (N_414,N_357,N_317);
nand U415 (N_415,N_336,N_370);
xor U416 (N_416,N_329,N_335);
and U417 (N_417,N_374,N_391);
or U418 (N_418,N_321,N_300);
nor U419 (N_419,N_381,N_396);
xor U420 (N_420,N_306,N_320);
and U421 (N_421,N_366,N_301);
or U422 (N_422,N_382,N_395);
nand U423 (N_423,N_328,N_394);
xor U424 (N_424,N_344,N_368);
nor U425 (N_425,N_340,N_302);
or U426 (N_426,N_303,N_324);
and U427 (N_427,N_322,N_380);
and U428 (N_428,N_375,N_377);
xnor U429 (N_429,N_392,N_314);
nor U430 (N_430,N_347,N_371);
xnor U431 (N_431,N_398,N_313);
and U432 (N_432,N_319,N_376);
nand U433 (N_433,N_354,N_316);
and U434 (N_434,N_399,N_311);
nand U435 (N_435,N_331,N_341);
nor U436 (N_436,N_304,N_358);
nor U437 (N_437,N_349,N_323);
and U438 (N_438,N_385,N_318);
or U439 (N_439,N_325,N_388);
nor U440 (N_440,N_309,N_326);
nand U441 (N_441,N_342,N_353);
and U442 (N_442,N_386,N_390);
or U443 (N_443,N_364,N_310);
nand U444 (N_444,N_345,N_337);
nor U445 (N_445,N_350,N_359);
nor U446 (N_446,N_343,N_307);
xnor U447 (N_447,N_379,N_369);
or U448 (N_448,N_332,N_389);
or U449 (N_449,N_383,N_315);
and U450 (N_450,N_309,N_393);
and U451 (N_451,N_300,N_370);
and U452 (N_452,N_393,N_383);
or U453 (N_453,N_312,N_324);
nand U454 (N_454,N_396,N_370);
and U455 (N_455,N_390,N_361);
and U456 (N_456,N_366,N_364);
xor U457 (N_457,N_336,N_386);
or U458 (N_458,N_374,N_370);
and U459 (N_459,N_336,N_345);
xor U460 (N_460,N_348,N_337);
nor U461 (N_461,N_310,N_377);
or U462 (N_462,N_342,N_335);
and U463 (N_463,N_339,N_316);
or U464 (N_464,N_302,N_385);
or U465 (N_465,N_312,N_300);
or U466 (N_466,N_389,N_398);
nor U467 (N_467,N_319,N_381);
and U468 (N_468,N_375,N_351);
nor U469 (N_469,N_389,N_363);
or U470 (N_470,N_327,N_369);
or U471 (N_471,N_306,N_343);
xnor U472 (N_472,N_384,N_318);
or U473 (N_473,N_357,N_316);
nand U474 (N_474,N_392,N_388);
nand U475 (N_475,N_387,N_369);
and U476 (N_476,N_381,N_391);
nand U477 (N_477,N_325,N_368);
nand U478 (N_478,N_363,N_337);
xor U479 (N_479,N_345,N_326);
nand U480 (N_480,N_362,N_305);
nor U481 (N_481,N_396,N_320);
and U482 (N_482,N_368,N_370);
and U483 (N_483,N_362,N_365);
or U484 (N_484,N_383,N_362);
nor U485 (N_485,N_390,N_307);
or U486 (N_486,N_327,N_337);
and U487 (N_487,N_321,N_343);
and U488 (N_488,N_314,N_322);
and U489 (N_489,N_311,N_312);
nor U490 (N_490,N_379,N_300);
nor U491 (N_491,N_397,N_338);
nor U492 (N_492,N_315,N_302);
nand U493 (N_493,N_381,N_345);
xor U494 (N_494,N_302,N_323);
nor U495 (N_495,N_385,N_340);
nor U496 (N_496,N_386,N_337);
nand U497 (N_497,N_303,N_322);
or U498 (N_498,N_362,N_325);
nor U499 (N_499,N_345,N_397);
or U500 (N_500,N_438,N_444);
nor U501 (N_501,N_414,N_485);
or U502 (N_502,N_497,N_455);
nor U503 (N_503,N_479,N_441);
or U504 (N_504,N_496,N_403);
or U505 (N_505,N_440,N_430);
or U506 (N_506,N_461,N_401);
xor U507 (N_507,N_437,N_458);
and U508 (N_508,N_415,N_431);
or U509 (N_509,N_498,N_474);
nor U510 (N_510,N_428,N_427);
xnor U511 (N_511,N_464,N_475);
nand U512 (N_512,N_468,N_484);
and U513 (N_513,N_400,N_499);
or U514 (N_514,N_442,N_443);
and U515 (N_515,N_466,N_448);
or U516 (N_516,N_404,N_463);
nor U517 (N_517,N_429,N_460);
or U518 (N_518,N_459,N_411);
or U519 (N_519,N_492,N_432);
nand U520 (N_520,N_446,N_433);
and U521 (N_521,N_476,N_491);
and U522 (N_522,N_451,N_453);
and U523 (N_523,N_471,N_421);
nand U524 (N_524,N_472,N_490);
nor U525 (N_525,N_450,N_405);
nor U526 (N_526,N_469,N_412);
and U527 (N_527,N_420,N_486);
or U528 (N_528,N_402,N_495);
and U529 (N_529,N_470,N_478);
nor U530 (N_530,N_473,N_447);
nand U531 (N_531,N_494,N_408);
nor U532 (N_532,N_423,N_409);
nor U533 (N_533,N_419,N_462);
nor U534 (N_534,N_467,N_482);
nor U535 (N_535,N_480,N_454);
nand U536 (N_536,N_416,N_445);
nor U537 (N_537,N_493,N_452);
nand U538 (N_538,N_483,N_426);
and U539 (N_539,N_456,N_457);
nand U540 (N_540,N_413,N_439);
or U541 (N_541,N_425,N_435);
nor U542 (N_542,N_418,N_449);
or U543 (N_543,N_488,N_424);
xor U544 (N_544,N_407,N_434);
or U545 (N_545,N_477,N_422);
or U546 (N_546,N_410,N_406);
nand U547 (N_547,N_417,N_436);
nand U548 (N_548,N_481,N_487);
and U549 (N_549,N_465,N_489);
xor U550 (N_550,N_428,N_479);
nor U551 (N_551,N_433,N_464);
or U552 (N_552,N_411,N_469);
and U553 (N_553,N_487,N_445);
and U554 (N_554,N_477,N_467);
nor U555 (N_555,N_497,N_474);
or U556 (N_556,N_431,N_465);
nand U557 (N_557,N_490,N_466);
xnor U558 (N_558,N_416,N_471);
and U559 (N_559,N_451,N_434);
or U560 (N_560,N_456,N_492);
nor U561 (N_561,N_405,N_465);
nand U562 (N_562,N_404,N_483);
nand U563 (N_563,N_466,N_474);
and U564 (N_564,N_442,N_485);
nand U565 (N_565,N_488,N_497);
and U566 (N_566,N_468,N_429);
or U567 (N_567,N_478,N_404);
nor U568 (N_568,N_494,N_485);
and U569 (N_569,N_482,N_472);
and U570 (N_570,N_433,N_441);
and U571 (N_571,N_425,N_484);
or U572 (N_572,N_456,N_477);
nand U573 (N_573,N_450,N_483);
nor U574 (N_574,N_405,N_423);
xnor U575 (N_575,N_456,N_452);
or U576 (N_576,N_487,N_484);
nor U577 (N_577,N_426,N_441);
nor U578 (N_578,N_469,N_401);
and U579 (N_579,N_418,N_487);
xor U580 (N_580,N_477,N_495);
nor U581 (N_581,N_426,N_488);
nor U582 (N_582,N_408,N_462);
and U583 (N_583,N_427,N_462);
xnor U584 (N_584,N_495,N_443);
nor U585 (N_585,N_414,N_408);
nor U586 (N_586,N_458,N_450);
nand U587 (N_587,N_435,N_430);
or U588 (N_588,N_473,N_492);
xnor U589 (N_589,N_422,N_456);
nor U590 (N_590,N_492,N_484);
or U591 (N_591,N_446,N_463);
and U592 (N_592,N_440,N_468);
xnor U593 (N_593,N_435,N_471);
and U594 (N_594,N_439,N_454);
or U595 (N_595,N_425,N_405);
nor U596 (N_596,N_465,N_475);
and U597 (N_597,N_492,N_443);
and U598 (N_598,N_484,N_419);
xnor U599 (N_599,N_405,N_490);
and U600 (N_600,N_553,N_560);
nor U601 (N_601,N_500,N_585);
or U602 (N_602,N_587,N_508);
and U603 (N_603,N_527,N_523);
or U604 (N_604,N_591,N_539);
and U605 (N_605,N_512,N_586);
and U606 (N_606,N_547,N_518);
xor U607 (N_607,N_558,N_574);
and U608 (N_608,N_532,N_505);
or U609 (N_609,N_564,N_517);
nand U610 (N_610,N_548,N_557);
nand U611 (N_611,N_502,N_521);
and U612 (N_612,N_542,N_573);
and U613 (N_613,N_568,N_597);
or U614 (N_614,N_504,N_596);
nor U615 (N_615,N_598,N_556);
nand U616 (N_616,N_524,N_584);
nand U617 (N_617,N_571,N_529);
and U618 (N_618,N_599,N_537);
and U619 (N_619,N_588,N_514);
nand U620 (N_620,N_575,N_538);
nand U621 (N_621,N_510,N_570);
or U622 (N_622,N_509,N_525);
or U623 (N_623,N_581,N_522);
or U624 (N_624,N_580,N_520);
nor U625 (N_625,N_530,N_569);
nor U626 (N_626,N_544,N_552);
nand U627 (N_627,N_565,N_540);
nand U628 (N_628,N_576,N_577);
or U629 (N_629,N_543,N_582);
nor U630 (N_630,N_583,N_506);
and U631 (N_631,N_516,N_562);
nor U632 (N_632,N_551,N_593);
nand U633 (N_633,N_541,N_566);
nand U634 (N_634,N_595,N_594);
nor U635 (N_635,N_536,N_579);
and U636 (N_636,N_507,N_572);
or U637 (N_637,N_526,N_563);
xor U638 (N_638,N_578,N_501);
nor U639 (N_639,N_519,N_513);
nor U640 (N_640,N_531,N_545);
or U641 (N_641,N_549,N_554);
nand U642 (N_642,N_546,N_534);
and U643 (N_643,N_528,N_535);
nand U644 (N_644,N_511,N_555);
nor U645 (N_645,N_503,N_533);
nand U646 (N_646,N_561,N_590);
nand U647 (N_647,N_559,N_550);
nor U648 (N_648,N_592,N_515);
nor U649 (N_649,N_567,N_589);
or U650 (N_650,N_517,N_553);
and U651 (N_651,N_595,N_557);
and U652 (N_652,N_517,N_597);
nand U653 (N_653,N_573,N_521);
nand U654 (N_654,N_554,N_537);
or U655 (N_655,N_590,N_547);
or U656 (N_656,N_505,N_556);
xnor U657 (N_657,N_565,N_570);
or U658 (N_658,N_544,N_523);
nor U659 (N_659,N_595,N_529);
or U660 (N_660,N_591,N_523);
nand U661 (N_661,N_573,N_586);
nor U662 (N_662,N_583,N_594);
or U663 (N_663,N_507,N_526);
nor U664 (N_664,N_516,N_542);
xor U665 (N_665,N_532,N_530);
or U666 (N_666,N_544,N_524);
nand U667 (N_667,N_537,N_589);
nand U668 (N_668,N_506,N_533);
xnor U669 (N_669,N_581,N_556);
nor U670 (N_670,N_553,N_556);
nand U671 (N_671,N_523,N_537);
nand U672 (N_672,N_514,N_516);
or U673 (N_673,N_591,N_548);
or U674 (N_674,N_526,N_559);
nor U675 (N_675,N_598,N_532);
or U676 (N_676,N_546,N_540);
or U677 (N_677,N_586,N_511);
and U678 (N_678,N_523,N_532);
nand U679 (N_679,N_596,N_531);
and U680 (N_680,N_539,N_500);
xor U681 (N_681,N_570,N_577);
nor U682 (N_682,N_547,N_504);
and U683 (N_683,N_534,N_564);
and U684 (N_684,N_551,N_574);
nand U685 (N_685,N_508,N_504);
or U686 (N_686,N_579,N_585);
or U687 (N_687,N_588,N_562);
or U688 (N_688,N_550,N_505);
nand U689 (N_689,N_504,N_595);
or U690 (N_690,N_508,N_585);
nand U691 (N_691,N_525,N_565);
or U692 (N_692,N_502,N_525);
nand U693 (N_693,N_565,N_538);
nor U694 (N_694,N_516,N_501);
xor U695 (N_695,N_556,N_559);
or U696 (N_696,N_541,N_535);
nor U697 (N_697,N_550,N_533);
nor U698 (N_698,N_513,N_507);
nand U699 (N_699,N_514,N_539);
xor U700 (N_700,N_618,N_612);
and U701 (N_701,N_688,N_646);
nor U702 (N_702,N_663,N_696);
or U703 (N_703,N_672,N_642);
and U704 (N_704,N_643,N_677);
nand U705 (N_705,N_621,N_640);
and U706 (N_706,N_699,N_611);
nor U707 (N_707,N_601,N_676);
and U708 (N_708,N_627,N_664);
or U709 (N_709,N_608,N_690);
nand U710 (N_710,N_683,N_686);
nor U711 (N_711,N_634,N_623);
or U712 (N_712,N_680,N_624);
or U713 (N_713,N_685,N_659);
nand U714 (N_714,N_671,N_668);
nand U715 (N_715,N_657,N_604);
or U716 (N_716,N_650,N_626);
nand U717 (N_717,N_691,N_630);
nand U718 (N_718,N_674,N_631);
nor U719 (N_719,N_605,N_665);
nor U720 (N_720,N_644,N_620);
or U721 (N_721,N_662,N_666);
xnor U722 (N_722,N_647,N_651);
or U723 (N_723,N_637,N_600);
and U724 (N_724,N_684,N_617);
nor U725 (N_725,N_682,N_609);
nand U726 (N_726,N_698,N_615);
and U727 (N_727,N_656,N_670);
nor U728 (N_728,N_629,N_675);
and U729 (N_729,N_669,N_689);
or U730 (N_730,N_697,N_693);
or U731 (N_731,N_614,N_692);
and U732 (N_732,N_649,N_622);
nand U733 (N_733,N_695,N_619);
xor U734 (N_734,N_658,N_628);
and U735 (N_735,N_679,N_606);
and U736 (N_736,N_638,N_613);
xor U737 (N_737,N_694,N_635);
nor U738 (N_738,N_654,N_616);
or U739 (N_739,N_687,N_602);
nor U740 (N_740,N_607,N_673);
and U741 (N_741,N_632,N_641);
and U742 (N_742,N_681,N_603);
and U743 (N_743,N_610,N_653);
or U744 (N_744,N_648,N_639);
nor U745 (N_745,N_660,N_645);
nand U746 (N_746,N_655,N_625);
and U747 (N_747,N_678,N_667);
and U748 (N_748,N_652,N_633);
nor U749 (N_749,N_661,N_636);
or U750 (N_750,N_655,N_689);
and U751 (N_751,N_692,N_643);
and U752 (N_752,N_636,N_600);
nand U753 (N_753,N_614,N_647);
and U754 (N_754,N_674,N_663);
or U755 (N_755,N_616,N_695);
or U756 (N_756,N_687,N_652);
or U757 (N_757,N_664,N_697);
nand U758 (N_758,N_657,N_667);
or U759 (N_759,N_618,N_619);
nand U760 (N_760,N_600,N_627);
xnor U761 (N_761,N_662,N_605);
nand U762 (N_762,N_685,N_617);
nand U763 (N_763,N_697,N_645);
xor U764 (N_764,N_650,N_617);
nand U765 (N_765,N_632,N_654);
and U766 (N_766,N_671,N_603);
nor U767 (N_767,N_613,N_653);
or U768 (N_768,N_693,N_652);
nand U769 (N_769,N_623,N_694);
xor U770 (N_770,N_645,N_608);
and U771 (N_771,N_696,N_623);
nor U772 (N_772,N_616,N_661);
or U773 (N_773,N_647,N_687);
or U774 (N_774,N_618,N_663);
nor U775 (N_775,N_600,N_611);
nor U776 (N_776,N_602,N_696);
nor U777 (N_777,N_659,N_681);
or U778 (N_778,N_601,N_652);
nor U779 (N_779,N_637,N_670);
and U780 (N_780,N_620,N_603);
nand U781 (N_781,N_654,N_653);
or U782 (N_782,N_675,N_698);
nand U783 (N_783,N_622,N_647);
nand U784 (N_784,N_672,N_635);
nor U785 (N_785,N_698,N_647);
and U786 (N_786,N_627,N_604);
nor U787 (N_787,N_633,N_670);
and U788 (N_788,N_661,N_697);
xnor U789 (N_789,N_676,N_662);
nand U790 (N_790,N_648,N_652);
or U791 (N_791,N_682,N_607);
or U792 (N_792,N_693,N_689);
nand U793 (N_793,N_686,N_608);
nor U794 (N_794,N_610,N_656);
nor U795 (N_795,N_676,N_648);
or U796 (N_796,N_640,N_600);
nor U797 (N_797,N_612,N_695);
nand U798 (N_798,N_615,N_636);
nor U799 (N_799,N_660,N_640);
nor U800 (N_800,N_744,N_730);
nor U801 (N_801,N_701,N_787);
xor U802 (N_802,N_781,N_716);
or U803 (N_803,N_767,N_705);
or U804 (N_804,N_712,N_735);
nor U805 (N_805,N_702,N_775);
or U806 (N_806,N_766,N_791);
nand U807 (N_807,N_727,N_770);
nor U808 (N_808,N_765,N_783);
nand U809 (N_809,N_714,N_725);
xnor U810 (N_810,N_737,N_792);
nor U811 (N_811,N_746,N_738);
or U812 (N_812,N_733,N_772);
xnor U813 (N_813,N_742,N_795);
xor U814 (N_814,N_711,N_752);
or U815 (N_815,N_762,N_718);
and U816 (N_816,N_754,N_773);
and U817 (N_817,N_768,N_736);
nor U818 (N_818,N_793,N_774);
nor U819 (N_819,N_782,N_786);
and U820 (N_820,N_759,N_731);
and U821 (N_821,N_704,N_753);
nand U822 (N_822,N_739,N_779);
or U823 (N_823,N_721,N_778);
or U824 (N_824,N_780,N_763);
nor U825 (N_825,N_761,N_700);
nor U826 (N_826,N_771,N_749);
or U827 (N_827,N_732,N_741);
nand U828 (N_828,N_799,N_729);
or U829 (N_829,N_709,N_788);
nand U830 (N_830,N_796,N_717);
nand U831 (N_831,N_745,N_760);
nand U832 (N_832,N_758,N_720);
and U833 (N_833,N_726,N_734);
and U834 (N_834,N_748,N_723);
and U835 (N_835,N_724,N_755);
or U836 (N_836,N_710,N_703);
and U837 (N_837,N_706,N_797);
nand U838 (N_838,N_751,N_708);
xnor U839 (N_839,N_713,N_776);
xnor U840 (N_840,N_719,N_707);
or U841 (N_841,N_757,N_740);
or U842 (N_842,N_747,N_784);
nor U843 (N_843,N_789,N_750);
nor U844 (N_844,N_769,N_777);
and U845 (N_845,N_785,N_743);
and U846 (N_846,N_790,N_794);
nand U847 (N_847,N_728,N_756);
and U848 (N_848,N_722,N_764);
nor U849 (N_849,N_715,N_798);
and U850 (N_850,N_737,N_779);
nor U851 (N_851,N_719,N_779);
or U852 (N_852,N_780,N_769);
nand U853 (N_853,N_789,N_719);
or U854 (N_854,N_763,N_757);
nor U855 (N_855,N_753,N_770);
or U856 (N_856,N_720,N_799);
and U857 (N_857,N_761,N_759);
or U858 (N_858,N_791,N_773);
nand U859 (N_859,N_756,N_755);
xor U860 (N_860,N_788,N_701);
xor U861 (N_861,N_743,N_779);
and U862 (N_862,N_763,N_770);
nand U863 (N_863,N_776,N_760);
and U864 (N_864,N_783,N_740);
or U865 (N_865,N_718,N_797);
nand U866 (N_866,N_717,N_727);
xnor U867 (N_867,N_754,N_786);
and U868 (N_868,N_736,N_748);
and U869 (N_869,N_713,N_774);
nand U870 (N_870,N_714,N_717);
and U871 (N_871,N_787,N_755);
and U872 (N_872,N_773,N_759);
and U873 (N_873,N_791,N_724);
nor U874 (N_874,N_766,N_735);
nand U875 (N_875,N_730,N_734);
nand U876 (N_876,N_703,N_745);
and U877 (N_877,N_763,N_708);
and U878 (N_878,N_735,N_739);
and U879 (N_879,N_779,N_776);
or U880 (N_880,N_731,N_741);
nor U881 (N_881,N_774,N_728);
or U882 (N_882,N_758,N_727);
and U883 (N_883,N_754,N_719);
or U884 (N_884,N_767,N_773);
nand U885 (N_885,N_793,N_787);
or U886 (N_886,N_772,N_713);
xnor U887 (N_887,N_796,N_707);
nand U888 (N_888,N_771,N_734);
nor U889 (N_889,N_771,N_784);
nand U890 (N_890,N_732,N_761);
and U891 (N_891,N_718,N_742);
nand U892 (N_892,N_750,N_704);
and U893 (N_893,N_705,N_756);
nor U894 (N_894,N_715,N_729);
nand U895 (N_895,N_755,N_727);
and U896 (N_896,N_742,N_788);
nand U897 (N_897,N_730,N_793);
nor U898 (N_898,N_761,N_747);
nor U899 (N_899,N_724,N_784);
and U900 (N_900,N_802,N_856);
or U901 (N_901,N_811,N_843);
or U902 (N_902,N_835,N_818);
xnor U903 (N_903,N_832,N_842);
xnor U904 (N_904,N_869,N_819);
nand U905 (N_905,N_801,N_836);
xnor U906 (N_906,N_866,N_851);
and U907 (N_907,N_810,N_840);
and U908 (N_908,N_897,N_875);
xor U909 (N_909,N_822,N_879);
nor U910 (N_910,N_839,N_855);
xor U911 (N_911,N_853,N_883);
nand U912 (N_912,N_884,N_820);
or U913 (N_913,N_837,N_824);
nand U914 (N_914,N_800,N_817);
nand U915 (N_915,N_878,N_877);
nand U916 (N_916,N_804,N_809);
nand U917 (N_917,N_889,N_826);
and U918 (N_918,N_895,N_821);
nand U919 (N_919,N_844,N_814);
or U920 (N_920,N_871,N_876);
and U921 (N_921,N_805,N_849);
and U922 (N_922,N_829,N_845);
nand U923 (N_923,N_860,N_854);
or U924 (N_924,N_813,N_899);
or U925 (N_925,N_867,N_887);
xor U926 (N_926,N_870,N_847);
or U927 (N_927,N_864,N_898);
nor U928 (N_928,N_896,N_865);
nor U929 (N_929,N_830,N_848);
or U930 (N_930,N_841,N_861);
and U931 (N_931,N_823,N_846);
nand U932 (N_932,N_868,N_880);
or U933 (N_933,N_850,N_833);
nor U934 (N_934,N_803,N_872);
nor U935 (N_935,N_807,N_891);
nor U936 (N_936,N_882,N_808);
and U937 (N_937,N_862,N_858);
or U938 (N_938,N_892,N_806);
and U939 (N_939,N_890,N_827);
and U940 (N_940,N_888,N_894);
nand U941 (N_941,N_834,N_893);
and U942 (N_942,N_838,N_825);
nand U943 (N_943,N_815,N_831);
or U944 (N_944,N_886,N_873);
nor U945 (N_945,N_812,N_859);
xnor U946 (N_946,N_874,N_828);
nand U947 (N_947,N_852,N_816);
nand U948 (N_948,N_863,N_857);
xnor U949 (N_949,N_885,N_881);
nor U950 (N_950,N_837,N_872);
nor U951 (N_951,N_899,N_821);
or U952 (N_952,N_819,N_879);
nand U953 (N_953,N_807,N_836);
nor U954 (N_954,N_818,N_814);
nor U955 (N_955,N_811,N_858);
and U956 (N_956,N_826,N_891);
or U957 (N_957,N_862,N_859);
and U958 (N_958,N_844,N_893);
nand U959 (N_959,N_854,N_818);
nor U960 (N_960,N_856,N_885);
or U961 (N_961,N_810,N_834);
and U962 (N_962,N_833,N_823);
or U963 (N_963,N_846,N_827);
nand U964 (N_964,N_849,N_813);
nand U965 (N_965,N_876,N_867);
or U966 (N_966,N_898,N_868);
or U967 (N_967,N_884,N_824);
nand U968 (N_968,N_856,N_811);
xnor U969 (N_969,N_894,N_835);
nand U970 (N_970,N_892,N_834);
nor U971 (N_971,N_849,N_821);
nor U972 (N_972,N_816,N_838);
nor U973 (N_973,N_868,N_859);
nand U974 (N_974,N_837,N_880);
nand U975 (N_975,N_801,N_825);
or U976 (N_976,N_806,N_818);
nand U977 (N_977,N_883,N_894);
or U978 (N_978,N_898,N_834);
nor U979 (N_979,N_887,N_884);
and U980 (N_980,N_836,N_859);
or U981 (N_981,N_884,N_885);
nor U982 (N_982,N_880,N_873);
xor U983 (N_983,N_895,N_899);
nor U984 (N_984,N_870,N_814);
and U985 (N_985,N_873,N_889);
nand U986 (N_986,N_807,N_804);
and U987 (N_987,N_874,N_875);
nand U988 (N_988,N_842,N_813);
nand U989 (N_989,N_887,N_817);
nor U990 (N_990,N_878,N_833);
nand U991 (N_991,N_808,N_872);
or U992 (N_992,N_841,N_877);
nand U993 (N_993,N_847,N_828);
nor U994 (N_994,N_820,N_861);
or U995 (N_995,N_860,N_835);
and U996 (N_996,N_817,N_854);
or U997 (N_997,N_865,N_863);
and U998 (N_998,N_832,N_860);
nand U999 (N_999,N_894,N_859);
or U1000 (N_1000,N_925,N_959);
xnor U1001 (N_1001,N_970,N_903);
or U1002 (N_1002,N_949,N_974);
and U1003 (N_1003,N_969,N_992);
and U1004 (N_1004,N_951,N_983);
nor U1005 (N_1005,N_968,N_953);
nand U1006 (N_1006,N_916,N_964);
nand U1007 (N_1007,N_991,N_962);
nor U1008 (N_1008,N_982,N_984);
or U1009 (N_1009,N_989,N_927);
nand U1010 (N_1010,N_977,N_996);
nand U1011 (N_1011,N_937,N_918);
and U1012 (N_1012,N_923,N_933);
nand U1013 (N_1013,N_935,N_911);
nand U1014 (N_1014,N_965,N_910);
nor U1015 (N_1015,N_913,N_939);
nor U1016 (N_1016,N_912,N_908);
nand U1017 (N_1017,N_955,N_952);
nor U1018 (N_1018,N_931,N_924);
and U1019 (N_1019,N_922,N_921);
and U1020 (N_1020,N_999,N_960);
nand U1021 (N_1021,N_920,N_917);
and U1022 (N_1022,N_915,N_919);
nor U1023 (N_1023,N_979,N_954);
or U1024 (N_1024,N_973,N_997);
xnor U1025 (N_1025,N_981,N_907);
nor U1026 (N_1026,N_987,N_948);
nor U1027 (N_1027,N_957,N_902);
nand U1028 (N_1028,N_958,N_944);
or U1029 (N_1029,N_929,N_928);
xnor U1030 (N_1030,N_942,N_995);
or U1031 (N_1031,N_978,N_909);
nor U1032 (N_1032,N_980,N_936);
xor U1033 (N_1033,N_967,N_994);
or U1034 (N_1034,N_945,N_963);
nand U1035 (N_1035,N_934,N_993);
or U1036 (N_1036,N_906,N_943);
and U1037 (N_1037,N_990,N_985);
or U1038 (N_1038,N_988,N_956);
and U1039 (N_1039,N_938,N_976);
xor U1040 (N_1040,N_901,N_914);
or U1041 (N_1041,N_947,N_966);
and U1042 (N_1042,N_904,N_930);
xor U1043 (N_1043,N_926,N_932);
nor U1044 (N_1044,N_961,N_940);
and U1045 (N_1045,N_986,N_905);
nand U1046 (N_1046,N_946,N_941);
nand U1047 (N_1047,N_998,N_972);
nand U1048 (N_1048,N_975,N_950);
nand U1049 (N_1049,N_971,N_900);
or U1050 (N_1050,N_990,N_982);
and U1051 (N_1051,N_937,N_997);
xnor U1052 (N_1052,N_954,N_912);
nor U1053 (N_1053,N_963,N_951);
nand U1054 (N_1054,N_972,N_944);
nor U1055 (N_1055,N_962,N_925);
nand U1056 (N_1056,N_950,N_900);
nor U1057 (N_1057,N_982,N_958);
or U1058 (N_1058,N_927,N_968);
or U1059 (N_1059,N_911,N_967);
nor U1060 (N_1060,N_924,N_921);
and U1061 (N_1061,N_908,N_943);
nand U1062 (N_1062,N_964,N_979);
and U1063 (N_1063,N_982,N_904);
nand U1064 (N_1064,N_907,N_913);
and U1065 (N_1065,N_921,N_986);
xor U1066 (N_1066,N_937,N_941);
nand U1067 (N_1067,N_939,N_968);
and U1068 (N_1068,N_940,N_959);
nor U1069 (N_1069,N_973,N_988);
and U1070 (N_1070,N_988,N_952);
and U1071 (N_1071,N_963,N_933);
xor U1072 (N_1072,N_937,N_982);
nor U1073 (N_1073,N_953,N_960);
or U1074 (N_1074,N_918,N_953);
or U1075 (N_1075,N_932,N_905);
and U1076 (N_1076,N_970,N_917);
or U1077 (N_1077,N_999,N_934);
nand U1078 (N_1078,N_981,N_919);
and U1079 (N_1079,N_937,N_987);
or U1080 (N_1080,N_920,N_951);
or U1081 (N_1081,N_950,N_998);
and U1082 (N_1082,N_906,N_921);
and U1083 (N_1083,N_971,N_933);
nand U1084 (N_1084,N_928,N_942);
xnor U1085 (N_1085,N_919,N_985);
or U1086 (N_1086,N_921,N_912);
nand U1087 (N_1087,N_937,N_957);
or U1088 (N_1088,N_944,N_947);
nand U1089 (N_1089,N_907,N_953);
or U1090 (N_1090,N_964,N_980);
or U1091 (N_1091,N_958,N_913);
and U1092 (N_1092,N_935,N_956);
xnor U1093 (N_1093,N_972,N_960);
and U1094 (N_1094,N_956,N_907);
nor U1095 (N_1095,N_917,N_950);
and U1096 (N_1096,N_916,N_918);
nand U1097 (N_1097,N_976,N_981);
nor U1098 (N_1098,N_989,N_985);
or U1099 (N_1099,N_930,N_987);
and U1100 (N_1100,N_1087,N_1099);
and U1101 (N_1101,N_1026,N_1004);
or U1102 (N_1102,N_1066,N_1031);
nor U1103 (N_1103,N_1092,N_1084);
nor U1104 (N_1104,N_1017,N_1063);
and U1105 (N_1105,N_1049,N_1057);
nand U1106 (N_1106,N_1091,N_1029);
nor U1107 (N_1107,N_1030,N_1023);
and U1108 (N_1108,N_1094,N_1032);
nor U1109 (N_1109,N_1076,N_1060);
and U1110 (N_1110,N_1075,N_1040);
and U1111 (N_1111,N_1007,N_1020);
nor U1112 (N_1112,N_1019,N_1078);
or U1113 (N_1113,N_1083,N_1041);
and U1114 (N_1114,N_1024,N_1038);
nor U1115 (N_1115,N_1003,N_1044);
or U1116 (N_1116,N_1055,N_1043);
nor U1117 (N_1117,N_1039,N_1065);
or U1118 (N_1118,N_1061,N_1018);
and U1119 (N_1119,N_1037,N_1001);
nor U1120 (N_1120,N_1062,N_1072);
or U1121 (N_1121,N_1077,N_1035);
or U1122 (N_1122,N_1027,N_1097);
nor U1123 (N_1123,N_1080,N_1006);
nand U1124 (N_1124,N_1089,N_1073);
or U1125 (N_1125,N_1047,N_1068);
nand U1126 (N_1126,N_1051,N_1033);
and U1127 (N_1127,N_1054,N_1088);
xor U1128 (N_1128,N_1013,N_1005);
xnor U1129 (N_1129,N_1015,N_1098);
nor U1130 (N_1130,N_1012,N_1000);
nor U1131 (N_1131,N_1002,N_1090);
or U1132 (N_1132,N_1011,N_1074);
or U1133 (N_1133,N_1095,N_1093);
nand U1134 (N_1134,N_1034,N_1079);
xnor U1135 (N_1135,N_1025,N_1064);
nor U1136 (N_1136,N_1045,N_1086);
xor U1137 (N_1137,N_1042,N_1067);
nand U1138 (N_1138,N_1016,N_1085);
nand U1139 (N_1139,N_1071,N_1096);
or U1140 (N_1140,N_1052,N_1008);
nor U1141 (N_1141,N_1010,N_1069);
nor U1142 (N_1142,N_1021,N_1070);
and U1143 (N_1143,N_1058,N_1050);
and U1144 (N_1144,N_1059,N_1036);
and U1145 (N_1145,N_1028,N_1014);
and U1146 (N_1146,N_1053,N_1046);
nand U1147 (N_1147,N_1009,N_1082);
or U1148 (N_1148,N_1022,N_1056);
nand U1149 (N_1149,N_1048,N_1081);
and U1150 (N_1150,N_1073,N_1054);
and U1151 (N_1151,N_1069,N_1072);
nand U1152 (N_1152,N_1047,N_1075);
and U1153 (N_1153,N_1072,N_1013);
and U1154 (N_1154,N_1002,N_1017);
and U1155 (N_1155,N_1092,N_1091);
nand U1156 (N_1156,N_1074,N_1090);
nor U1157 (N_1157,N_1000,N_1037);
nor U1158 (N_1158,N_1079,N_1001);
xnor U1159 (N_1159,N_1077,N_1061);
nand U1160 (N_1160,N_1091,N_1012);
or U1161 (N_1161,N_1080,N_1085);
and U1162 (N_1162,N_1062,N_1049);
and U1163 (N_1163,N_1021,N_1019);
nor U1164 (N_1164,N_1006,N_1082);
or U1165 (N_1165,N_1078,N_1044);
nor U1166 (N_1166,N_1053,N_1041);
or U1167 (N_1167,N_1042,N_1009);
and U1168 (N_1168,N_1078,N_1060);
and U1169 (N_1169,N_1024,N_1095);
and U1170 (N_1170,N_1031,N_1092);
nand U1171 (N_1171,N_1054,N_1049);
or U1172 (N_1172,N_1090,N_1022);
nand U1173 (N_1173,N_1049,N_1066);
nand U1174 (N_1174,N_1047,N_1043);
and U1175 (N_1175,N_1088,N_1055);
xor U1176 (N_1176,N_1088,N_1085);
or U1177 (N_1177,N_1068,N_1089);
xor U1178 (N_1178,N_1078,N_1038);
or U1179 (N_1179,N_1003,N_1081);
and U1180 (N_1180,N_1077,N_1016);
or U1181 (N_1181,N_1027,N_1089);
nand U1182 (N_1182,N_1099,N_1042);
xor U1183 (N_1183,N_1089,N_1082);
xnor U1184 (N_1184,N_1030,N_1042);
and U1185 (N_1185,N_1067,N_1014);
nand U1186 (N_1186,N_1008,N_1024);
nor U1187 (N_1187,N_1071,N_1006);
or U1188 (N_1188,N_1097,N_1076);
nor U1189 (N_1189,N_1062,N_1092);
or U1190 (N_1190,N_1093,N_1016);
xor U1191 (N_1191,N_1037,N_1068);
or U1192 (N_1192,N_1084,N_1001);
or U1193 (N_1193,N_1081,N_1086);
or U1194 (N_1194,N_1077,N_1033);
xnor U1195 (N_1195,N_1041,N_1004);
and U1196 (N_1196,N_1019,N_1000);
and U1197 (N_1197,N_1073,N_1099);
or U1198 (N_1198,N_1007,N_1013);
nor U1199 (N_1199,N_1012,N_1027);
and U1200 (N_1200,N_1111,N_1129);
or U1201 (N_1201,N_1149,N_1173);
nand U1202 (N_1202,N_1137,N_1164);
and U1203 (N_1203,N_1169,N_1153);
nor U1204 (N_1204,N_1194,N_1140);
nor U1205 (N_1205,N_1117,N_1132);
and U1206 (N_1206,N_1178,N_1109);
and U1207 (N_1207,N_1158,N_1185);
nand U1208 (N_1208,N_1191,N_1130);
nand U1209 (N_1209,N_1151,N_1126);
and U1210 (N_1210,N_1179,N_1182);
xnor U1211 (N_1211,N_1197,N_1120);
nand U1212 (N_1212,N_1199,N_1112);
or U1213 (N_1213,N_1105,N_1189);
nor U1214 (N_1214,N_1104,N_1174);
nand U1215 (N_1215,N_1113,N_1198);
or U1216 (N_1216,N_1157,N_1118);
nor U1217 (N_1217,N_1188,N_1196);
and U1218 (N_1218,N_1146,N_1102);
and U1219 (N_1219,N_1150,N_1119);
nor U1220 (N_1220,N_1123,N_1171);
and U1221 (N_1221,N_1186,N_1116);
or U1222 (N_1222,N_1177,N_1165);
or U1223 (N_1223,N_1124,N_1122);
xor U1224 (N_1224,N_1159,N_1160);
nand U1225 (N_1225,N_1175,N_1141);
or U1226 (N_1226,N_1145,N_1155);
nor U1227 (N_1227,N_1166,N_1156);
or U1228 (N_1228,N_1107,N_1110);
and U1229 (N_1229,N_1135,N_1192);
or U1230 (N_1230,N_1139,N_1187);
xor U1231 (N_1231,N_1163,N_1127);
nor U1232 (N_1232,N_1103,N_1154);
nand U1233 (N_1233,N_1134,N_1142);
or U1234 (N_1234,N_1193,N_1136);
and U1235 (N_1235,N_1101,N_1131);
nand U1236 (N_1236,N_1162,N_1133);
and U1237 (N_1237,N_1167,N_1195);
nand U1238 (N_1238,N_1125,N_1148);
nor U1239 (N_1239,N_1183,N_1114);
xnor U1240 (N_1240,N_1161,N_1128);
nor U1241 (N_1241,N_1143,N_1100);
nand U1242 (N_1242,N_1147,N_1108);
or U1243 (N_1243,N_1106,N_1180);
xnor U1244 (N_1244,N_1152,N_1181);
or U1245 (N_1245,N_1138,N_1115);
and U1246 (N_1246,N_1144,N_1170);
nand U1247 (N_1247,N_1190,N_1176);
and U1248 (N_1248,N_1184,N_1121);
and U1249 (N_1249,N_1168,N_1172);
or U1250 (N_1250,N_1128,N_1179);
nand U1251 (N_1251,N_1152,N_1117);
xnor U1252 (N_1252,N_1177,N_1196);
nand U1253 (N_1253,N_1176,N_1128);
nor U1254 (N_1254,N_1197,N_1185);
and U1255 (N_1255,N_1150,N_1133);
nand U1256 (N_1256,N_1118,N_1128);
nor U1257 (N_1257,N_1193,N_1154);
or U1258 (N_1258,N_1173,N_1131);
and U1259 (N_1259,N_1184,N_1190);
and U1260 (N_1260,N_1162,N_1157);
nor U1261 (N_1261,N_1153,N_1104);
or U1262 (N_1262,N_1113,N_1158);
and U1263 (N_1263,N_1102,N_1175);
nor U1264 (N_1264,N_1188,N_1157);
or U1265 (N_1265,N_1187,N_1178);
nor U1266 (N_1266,N_1166,N_1168);
or U1267 (N_1267,N_1179,N_1178);
and U1268 (N_1268,N_1192,N_1142);
nor U1269 (N_1269,N_1100,N_1189);
xnor U1270 (N_1270,N_1187,N_1121);
xnor U1271 (N_1271,N_1176,N_1116);
or U1272 (N_1272,N_1142,N_1199);
nand U1273 (N_1273,N_1182,N_1133);
nor U1274 (N_1274,N_1145,N_1148);
nor U1275 (N_1275,N_1111,N_1188);
nand U1276 (N_1276,N_1167,N_1128);
nor U1277 (N_1277,N_1151,N_1191);
nand U1278 (N_1278,N_1196,N_1180);
nand U1279 (N_1279,N_1168,N_1111);
and U1280 (N_1280,N_1116,N_1180);
or U1281 (N_1281,N_1173,N_1159);
nand U1282 (N_1282,N_1167,N_1106);
nor U1283 (N_1283,N_1120,N_1124);
and U1284 (N_1284,N_1122,N_1133);
nand U1285 (N_1285,N_1139,N_1171);
or U1286 (N_1286,N_1142,N_1126);
nand U1287 (N_1287,N_1179,N_1154);
and U1288 (N_1288,N_1196,N_1197);
and U1289 (N_1289,N_1109,N_1153);
nor U1290 (N_1290,N_1113,N_1135);
and U1291 (N_1291,N_1178,N_1111);
nor U1292 (N_1292,N_1151,N_1183);
nand U1293 (N_1293,N_1180,N_1186);
nor U1294 (N_1294,N_1141,N_1113);
nand U1295 (N_1295,N_1100,N_1162);
and U1296 (N_1296,N_1162,N_1134);
or U1297 (N_1297,N_1139,N_1191);
nor U1298 (N_1298,N_1176,N_1141);
nor U1299 (N_1299,N_1119,N_1106);
or U1300 (N_1300,N_1204,N_1207);
nand U1301 (N_1301,N_1298,N_1245);
nor U1302 (N_1302,N_1200,N_1213);
xnor U1303 (N_1303,N_1292,N_1224);
and U1304 (N_1304,N_1253,N_1265);
or U1305 (N_1305,N_1209,N_1285);
or U1306 (N_1306,N_1288,N_1262);
nor U1307 (N_1307,N_1293,N_1252);
or U1308 (N_1308,N_1210,N_1283);
and U1309 (N_1309,N_1244,N_1264);
and U1310 (N_1310,N_1220,N_1241);
and U1311 (N_1311,N_1231,N_1273);
nand U1312 (N_1312,N_1233,N_1257);
and U1313 (N_1313,N_1280,N_1259);
nand U1314 (N_1314,N_1297,N_1246);
or U1315 (N_1315,N_1277,N_1232);
nor U1316 (N_1316,N_1203,N_1261);
nor U1317 (N_1317,N_1222,N_1238);
xor U1318 (N_1318,N_1208,N_1291);
nor U1319 (N_1319,N_1254,N_1249);
and U1320 (N_1320,N_1202,N_1235);
nor U1321 (N_1321,N_1263,N_1230);
nand U1322 (N_1322,N_1279,N_1219);
nor U1323 (N_1323,N_1211,N_1229);
and U1324 (N_1324,N_1251,N_1296);
or U1325 (N_1325,N_1256,N_1276);
nand U1326 (N_1326,N_1278,N_1275);
nand U1327 (N_1327,N_1248,N_1289);
nor U1328 (N_1328,N_1295,N_1214);
nand U1329 (N_1329,N_1271,N_1247);
or U1330 (N_1330,N_1243,N_1221);
nor U1331 (N_1331,N_1223,N_1227);
or U1332 (N_1332,N_1242,N_1236);
nand U1333 (N_1333,N_1281,N_1260);
nand U1334 (N_1334,N_1216,N_1205);
or U1335 (N_1335,N_1299,N_1282);
or U1336 (N_1336,N_1274,N_1255);
and U1337 (N_1337,N_1284,N_1270);
nor U1338 (N_1338,N_1239,N_1206);
nor U1339 (N_1339,N_1225,N_1217);
nor U1340 (N_1340,N_1286,N_1294);
and U1341 (N_1341,N_1269,N_1228);
xor U1342 (N_1342,N_1201,N_1266);
or U1343 (N_1343,N_1258,N_1218);
or U1344 (N_1344,N_1240,N_1272);
nand U1345 (N_1345,N_1290,N_1287);
and U1346 (N_1346,N_1268,N_1237);
and U1347 (N_1347,N_1215,N_1226);
nand U1348 (N_1348,N_1267,N_1250);
or U1349 (N_1349,N_1212,N_1234);
nor U1350 (N_1350,N_1273,N_1291);
xor U1351 (N_1351,N_1220,N_1226);
and U1352 (N_1352,N_1266,N_1274);
nor U1353 (N_1353,N_1256,N_1233);
nand U1354 (N_1354,N_1214,N_1241);
nand U1355 (N_1355,N_1272,N_1201);
nor U1356 (N_1356,N_1216,N_1299);
or U1357 (N_1357,N_1285,N_1284);
nand U1358 (N_1358,N_1241,N_1244);
or U1359 (N_1359,N_1299,N_1220);
nand U1360 (N_1360,N_1270,N_1287);
nor U1361 (N_1361,N_1203,N_1229);
or U1362 (N_1362,N_1298,N_1239);
xor U1363 (N_1363,N_1273,N_1233);
nand U1364 (N_1364,N_1284,N_1298);
xnor U1365 (N_1365,N_1216,N_1239);
and U1366 (N_1366,N_1290,N_1271);
or U1367 (N_1367,N_1255,N_1269);
and U1368 (N_1368,N_1256,N_1241);
nand U1369 (N_1369,N_1275,N_1247);
and U1370 (N_1370,N_1272,N_1297);
or U1371 (N_1371,N_1286,N_1234);
or U1372 (N_1372,N_1262,N_1217);
or U1373 (N_1373,N_1225,N_1203);
xnor U1374 (N_1374,N_1212,N_1290);
nor U1375 (N_1375,N_1233,N_1293);
nand U1376 (N_1376,N_1208,N_1243);
nand U1377 (N_1377,N_1235,N_1274);
and U1378 (N_1378,N_1285,N_1216);
nand U1379 (N_1379,N_1254,N_1271);
and U1380 (N_1380,N_1200,N_1276);
and U1381 (N_1381,N_1254,N_1269);
nand U1382 (N_1382,N_1281,N_1289);
nor U1383 (N_1383,N_1211,N_1218);
nor U1384 (N_1384,N_1210,N_1239);
nand U1385 (N_1385,N_1230,N_1246);
or U1386 (N_1386,N_1284,N_1245);
xnor U1387 (N_1387,N_1277,N_1287);
nor U1388 (N_1388,N_1254,N_1244);
nor U1389 (N_1389,N_1205,N_1266);
or U1390 (N_1390,N_1299,N_1225);
nor U1391 (N_1391,N_1261,N_1297);
or U1392 (N_1392,N_1264,N_1271);
or U1393 (N_1393,N_1293,N_1284);
and U1394 (N_1394,N_1292,N_1288);
nand U1395 (N_1395,N_1248,N_1251);
nor U1396 (N_1396,N_1256,N_1205);
xor U1397 (N_1397,N_1282,N_1225);
or U1398 (N_1398,N_1284,N_1259);
or U1399 (N_1399,N_1244,N_1209);
and U1400 (N_1400,N_1309,N_1322);
nand U1401 (N_1401,N_1344,N_1383);
or U1402 (N_1402,N_1390,N_1382);
and U1403 (N_1403,N_1362,N_1371);
nand U1404 (N_1404,N_1300,N_1334);
and U1405 (N_1405,N_1324,N_1338);
nand U1406 (N_1406,N_1337,N_1384);
xnor U1407 (N_1407,N_1323,N_1319);
nor U1408 (N_1408,N_1389,N_1378);
and U1409 (N_1409,N_1341,N_1333);
nor U1410 (N_1410,N_1353,N_1398);
or U1411 (N_1411,N_1352,N_1381);
nor U1412 (N_1412,N_1386,N_1311);
nand U1413 (N_1413,N_1336,N_1376);
or U1414 (N_1414,N_1315,N_1327);
or U1415 (N_1415,N_1325,N_1303);
xnor U1416 (N_1416,N_1368,N_1346);
and U1417 (N_1417,N_1304,N_1366);
xnor U1418 (N_1418,N_1356,N_1365);
or U1419 (N_1419,N_1348,N_1375);
nor U1420 (N_1420,N_1354,N_1359);
or U1421 (N_1421,N_1310,N_1329);
or U1422 (N_1422,N_1330,N_1318);
and U1423 (N_1423,N_1392,N_1313);
nor U1424 (N_1424,N_1345,N_1360);
nor U1425 (N_1425,N_1340,N_1397);
or U1426 (N_1426,N_1363,N_1307);
or U1427 (N_1427,N_1373,N_1316);
or U1428 (N_1428,N_1342,N_1317);
or U1429 (N_1429,N_1374,N_1350);
xnor U1430 (N_1430,N_1347,N_1393);
nand U1431 (N_1431,N_1358,N_1391);
nor U1432 (N_1432,N_1305,N_1321);
and U1433 (N_1433,N_1332,N_1357);
and U1434 (N_1434,N_1361,N_1399);
nor U1435 (N_1435,N_1301,N_1302);
nor U1436 (N_1436,N_1388,N_1339);
xnor U1437 (N_1437,N_1380,N_1306);
nor U1438 (N_1438,N_1395,N_1370);
and U1439 (N_1439,N_1396,N_1343);
nand U1440 (N_1440,N_1326,N_1385);
and U1441 (N_1441,N_1367,N_1394);
and U1442 (N_1442,N_1308,N_1320);
or U1443 (N_1443,N_1335,N_1387);
or U1444 (N_1444,N_1349,N_1379);
and U1445 (N_1445,N_1377,N_1372);
and U1446 (N_1446,N_1351,N_1328);
and U1447 (N_1447,N_1314,N_1369);
xnor U1448 (N_1448,N_1364,N_1355);
or U1449 (N_1449,N_1312,N_1331);
or U1450 (N_1450,N_1349,N_1392);
or U1451 (N_1451,N_1398,N_1380);
nand U1452 (N_1452,N_1369,N_1364);
or U1453 (N_1453,N_1377,N_1332);
nor U1454 (N_1454,N_1331,N_1315);
nor U1455 (N_1455,N_1328,N_1325);
nand U1456 (N_1456,N_1355,N_1349);
and U1457 (N_1457,N_1389,N_1333);
xnor U1458 (N_1458,N_1359,N_1317);
xor U1459 (N_1459,N_1332,N_1380);
nor U1460 (N_1460,N_1349,N_1318);
nand U1461 (N_1461,N_1321,N_1369);
nor U1462 (N_1462,N_1317,N_1373);
xor U1463 (N_1463,N_1354,N_1360);
nand U1464 (N_1464,N_1327,N_1359);
nor U1465 (N_1465,N_1312,N_1303);
nor U1466 (N_1466,N_1333,N_1319);
and U1467 (N_1467,N_1333,N_1381);
nand U1468 (N_1468,N_1355,N_1334);
nand U1469 (N_1469,N_1330,N_1369);
or U1470 (N_1470,N_1324,N_1315);
or U1471 (N_1471,N_1393,N_1341);
nor U1472 (N_1472,N_1307,N_1395);
and U1473 (N_1473,N_1321,N_1312);
nand U1474 (N_1474,N_1312,N_1349);
nor U1475 (N_1475,N_1380,N_1316);
or U1476 (N_1476,N_1391,N_1347);
xor U1477 (N_1477,N_1358,N_1332);
nand U1478 (N_1478,N_1393,N_1370);
and U1479 (N_1479,N_1376,N_1384);
or U1480 (N_1480,N_1304,N_1332);
nand U1481 (N_1481,N_1326,N_1338);
or U1482 (N_1482,N_1332,N_1359);
xnor U1483 (N_1483,N_1347,N_1359);
xor U1484 (N_1484,N_1356,N_1377);
nor U1485 (N_1485,N_1367,N_1339);
or U1486 (N_1486,N_1388,N_1393);
nand U1487 (N_1487,N_1341,N_1331);
and U1488 (N_1488,N_1315,N_1349);
or U1489 (N_1489,N_1310,N_1313);
nand U1490 (N_1490,N_1385,N_1354);
or U1491 (N_1491,N_1319,N_1334);
and U1492 (N_1492,N_1361,N_1300);
or U1493 (N_1493,N_1379,N_1360);
and U1494 (N_1494,N_1358,N_1322);
xor U1495 (N_1495,N_1399,N_1382);
nor U1496 (N_1496,N_1324,N_1303);
nand U1497 (N_1497,N_1343,N_1384);
and U1498 (N_1498,N_1362,N_1396);
or U1499 (N_1499,N_1332,N_1390);
nor U1500 (N_1500,N_1446,N_1447);
nor U1501 (N_1501,N_1487,N_1445);
nand U1502 (N_1502,N_1474,N_1490);
or U1503 (N_1503,N_1460,N_1483);
xnor U1504 (N_1504,N_1481,N_1443);
or U1505 (N_1505,N_1444,N_1492);
and U1506 (N_1506,N_1424,N_1463);
or U1507 (N_1507,N_1478,N_1468);
nor U1508 (N_1508,N_1406,N_1488);
xor U1509 (N_1509,N_1485,N_1428);
or U1510 (N_1510,N_1470,N_1459);
or U1511 (N_1511,N_1491,N_1429);
nor U1512 (N_1512,N_1454,N_1438);
nand U1513 (N_1513,N_1453,N_1411);
nand U1514 (N_1514,N_1415,N_1426);
and U1515 (N_1515,N_1472,N_1482);
nand U1516 (N_1516,N_1440,N_1430);
nand U1517 (N_1517,N_1461,N_1419);
and U1518 (N_1518,N_1476,N_1402);
nor U1519 (N_1519,N_1442,N_1477);
and U1520 (N_1520,N_1400,N_1499);
and U1521 (N_1521,N_1416,N_1455);
or U1522 (N_1522,N_1464,N_1417);
nor U1523 (N_1523,N_1452,N_1433);
or U1524 (N_1524,N_1410,N_1404);
nor U1525 (N_1525,N_1493,N_1422);
nand U1526 (N_1526,N_1423,N_1401);
nand U1527 (N_1527,N_1449,N_1420);
nand U1528 (N_1528,N_1489,N_1418);
or U1529 (N_1529,N_1427,N_1412);
nand U1530 (N_1530,N_1467,N_1434);
or U1531 (N_1531,N_1462,N_1473);
and U1532 (N_1532,N_1479,N_1407);
or U1533 (N_1533,N_1439,N_1408);
and U1534 (N_1534,N_1436,N_1486);
nor U1535 (N_1535,N_1471,N_1495);
nand U1536 (N_1536,N_1457,N_1494);
and U1537 (N_1537,N_1437,N_1405);
nand U1538 (N_1538,N_1432,N_1435);
and U1539 (N_1539,N_1498,N_1409);
nand U1540 (N_1540,N_1484,N_1403);
nor U1541 (N_1541,N_1480,N_1475);
nand U1542 (N_1542,N_1450,N_1414);
or U1543 (N_1543,N_1431,N_1497);
or U1544 (N_1544,N_1458,N_1496);
and U1545 (N_1545,N_1421,N_1425);
nor U1546 (N_1546,N_1465,N_1456);
or U1547 (N_1547,N_1413,N_1469);
or U1548 (N_1548,N_1448,N_1466);
and U1549 (N_1549,N_1451,N_1441);
nor U1550 (N_1550,N_1435,N_1449);
nand U1551 (N_1551,N_1419,N_1423);
nor U1552 (N_1552,N_1404,N_1440);
or U1553 (N_1553,N_1430,N_1412);
nand U1554 (N_1554,N_1471,N_1427);
or U1555 (N_1555,N_1418,N_1475);
or U1556 (N_1556,N_1458,N_1468);
nor U1557 (N_1557,N_1425,N_1439);
or U1558 (N_1558,N_1458,N_1453);
nor U1559 (N_1559,N_1460,N_1406);
and U1560 (N_1560,N_1413,N_1470);
nand U1561 (N_1561,N_1417,N_1445);
or U1562 (N_1562,N_1491,N_1413);
and U1563 (N_1563,N_1413,N_1439);
or U1564 (N_1564,N_1429,N_1464);
or U1565 (N_1565,N_1453,N_1419);
nand U1566 (N_1566,N_1406,N_1444);
or U1567 (N_1567,N_1434,N_1446);
or U1568 (N_1568,N_1412,N_1417);
nor U1569 (N_1569,N_1462,N_1489);
nand U1570 (N_1570,N_1431,N_1465);
nor U1571 (N_1571,N_1451,N_1490);
or U1572 (N_1572,N_1454,N_1486);
nor U1573 (N_1573,N_1465,N_1421);
xnor U1574 (N_1574,N_1409,N_1418);
or U1575 (N_1575,N_1415,N_1441);
nor U1576 (N_1576,N_1410,N_1487);
xnor U1577 (N_1577,N_1468,N_1467);
nand U1578 (N_1578,N_1445,N_1497);
nand U1579 (N_1579,N_1401,N_1477);
xor U1580 (N_1580,N_1482,N_1498);
xor U1581 (N_1581,N_1495,N_1474);
xnor U1582 (N_1582,N_1439,N_1433);
or U1583 (N_1583,N_1433,N_1445);
nor U1584 (N_1584,N_1428,N_1417);
xor U1585 (N_1585,N_1458,N_1406);
and U1586 (N_1586,N_1426,N_1461);
or U1587 (N_1587,N_1472,N_1416);
and U1588 (N_1588,N_1450,N_1497);
and U1589 (N_1589,N_1479,N_1493);
or U1590 (N_1590,N_1494,N_1450);
or U1591 (N_1591,N_1437,N_1465);
and U1592 (N_1592,N_1407,N_1440);
or U1593 (N_1593,N_1400,N_1411);
xnor U1594 (N_1594,N_1423,N_1411);
and U1595 (N_1595,N_1454,N_1418);
nand U1596 (N_1596,N_1423,N_1409);
xnor U1597 (N_1597,N_1490,N_1466);
or U1598 (N_1598,N_1455,N_1436);
or U1599 (N_1599,N_1474,N_1457);
and U1600 (N_1600,N_1523,N_1596);
or U1601 (N_1601,N_1546,N_1576);
nand U1602 (N_1602,N_1510,N_1530);
or U1603 (N_1603,N_1502,N_1504);
nand U1604 (N_1604,N_1593,N_1532);
nand U1605 (N_1605,N_1515,N_1568);
nor U1606 (N_1606,N_1558,N_1579);
or U1607 (N_1607,N_1524,N_1506);
and U1608 (N_1608,N_1552,N_1551);
or U1609 (N_1609,N_1525,N_1560);
nand U1610 (N_1610,N_1538,N_1561);
or U1611 (N_1611,N_1567,N_1574);
nor U1612 (N_1612,N_1597,N_1543);
and U1613 (N_1613,N_1501,N_1583);
nand U1614 (N_1614,N_1549,N_1589);
xnor U1615 (N_1615,N_1586,N_1598);
nand U1616 (N_1616,N_1587,N_1557);
or U1617 (N_1617,N_1585,N_1595);
and U1618 (N_1618,N_1513,N_1518);
xnor U1619 (N_1619,N_1516,N_1545);
and U1620 (N_1620,N_1580,N_1590);
nor U1621 (N_1621,N_1533,N_1522);
and U1622 (N_1622,N_1584,N_1521);
and U1623 (N_1623,N_1550,N_1534);
or U1624 (N_1624,N_1503,N_1535);
or U1625 (N_1625,N_1527,N_1565);
or U1626 (N_1626,N_1573,N_1582);
nor U1627 (N_1627,N_1547,N_1517);
or U1628 (N_1628,N_1508,N_1520);
nand U1629 (N_1629,N_1581,N_1507);
nand U1630 (N_1630,N_1539,N_1536);
xnor U1631 (N_1631,N_1559,N_1572);
or U1632 (N_1632,N_1514,N_1511);
nand U1633 (N_1633,N_1528,N_1519);
nor U1634 (N_1634,N_1540,N_1591);
and U1635 (N_1635,N_1505,N_1577);
and U1636 (N_1636,N_1556,N_1575);
nor U1637 (N_1637,N_1541,N_1578);
xor U1638 (N_1638,N_1555,N_1544);
nand U1639 (N_1639,N_1594,N_1571);
or U1640 (N_1640,N_1553,N_1531);
and U1641 (N_1641,N_1512,N_1569);
nand U1642 (N_1642,N_1563,N_1548);
nand U1643 (N_1643,N_1588,N_1562);
nor U1644 (N_1644,N_1554,N_1500);
nand U1645 (N_1645,N_1526,N_1529);
or U1646 (N_1646,N_1564,N_1542);
or U1647 (N_1647,N_1566,N_1570);
or U1648 (N_1648,N_1537,N_1592);
and U1649 (N_1649,N_1599,N_1509);
nor U1650 (N_1650,N_1556,N_1574);
nor U1651 (N_1651,N_1556,N_1562);
or U1652 (N_1652,N_1527,N_1513);
nor U1653 (N_1653,N_1509,N_1536);
or U1654 (N_1654,N_1549,N_1551);
and U1655 (N_1655,N_1545,N_1513);
and U1656 (N_1656,N_1599,N_1507);
or U1657 (N_1657,N_1577,N_1578);
xor U1658 (N_1658,N_1581,N_1552);
and U1659 (N_1659,N_1553,N_1591);
and U1660 (N_1660,N_1579,N_1555);
and U1661 (N_1661,N_1578,N_1525);
nand U1662 (N_1662,N_1531,N_1512);
or U1663 (N_1663,N_1591,N_1527);
or U1664 (N_1664,N_1579,N_1544);
nor U1665 (N_1665,N_1502,N_1569);
or U1666 (N_1666,N_1530,N_1587);
nand U1667 (N_1667,N_1546,N_1536);
nor U1668 (N_1668,N_1566,N_1580);
nand U1669 (N_1669,N_1517,N_1546);
and U1670 (N_1670,N_1577,N_1529);
nand U1671 (N_1671,N_1521,N_1505);
nand U1672 (N_1672,N_1509,N_1579);
or U1673 (N_1673,N_1504,N_1561);
nor U1674 (N_1674,N_1588,N_1591);
and U1675 (N_1675,N_1512,N_1575);
or U1676 (N_1676,N_1582,N_1515);
or U1677 (N_1677,N_1541,N_1588);
or U1678 (N_1678,N_1559,N_1579);
and U1679 (N_1679,N_1595,N_1513);
nand U1680 (N_1680,N_1546,N_1574);
nand U1681 (N_1681,N_1587,N_1507);
nand U1682 (N_1682,N_1543,N_1552);
xnor U1683 (N_1683,N_1517,N_1566);
or U1684 (N_1684,N_1558,N_1574);
and U1685 (N_1685,N_1553,N_1543);
nor U1686 (N_1686,N_1531,N_1501);
nand U1687 (N_1687,N_1555,N_1521);
nand U1688 (N_1688,N_1565,N_1564);
nand U1689 (N_1689,N_1576,N_1571);
xor U1690 (N_1690,N_1505,N_1550);
and U1691 (N_1691,N_1579,N_1560);
and U1692 (N_1692,N_1581,N_1596);
nor U1693 (N_1693,N_1572,N_1552);
nor U1694 (N_1694,N_1592,N_1531);
or U1695 (N_1695,N_1569,N_1561);
nand U1696 (N_1696,N_1519,N_1540);
nor U1697 (N_1697,N_1516,N_1543);
nor U1698 (N_1698,N_1512,N_1570);
and U1699 (N_1699,N_1505,N_1595);
and U1700 (N_1700,N_1637,N_1613);
and U1701 (N_1701,N_1691,N_1622);
or U1702 (N_1702,N_1635,N_1620);
nor U1703 (N_1703,N_1669,N_1663);
xnor U1704 (N_1704,N_1658,N_1606);
nor U1705 (N_1705,N_1661,N_1608);
and U1706 (N_1706,N_1642,N_1654);
and U1707 (N_1707,N_1660,N_1629);
xor U1708 (N_1708,N_1632,N_1670);
nor U1709 (N_1709,N_1696,N_1648);
and U1710 (N_1710,N_1664,N_1610);
or U1711 (N_1711,N_1619,N_1655);
nor U1712 (N_1712,N_1600,N_1602);
xnor U1713 (N_1713,N_1607,N_1690);
nor U1714 (N_1714,N_1639,N_1653);
xor U1715 (N_1715,N_1671,N_1640);
and U1716 (N_1716,N_1621,N_1684);
nand U1717 (N_1717,N_1689,N_1627);
or U1718 (N_1718,N_1611,N_1644);
or U1719 (N_1719,N_1617,N_1666);
nor U1720 (N_1720,N_1659,N_1626);
or U1721 (N_1721,N_1618,N_1657);
and U1722 (N_1722,N_1677,N_1628);
and U1723 (N_1723,N_1634,N_1630);
nand U1724 (N_1724,N_1652,N_1674);
and U1725 (N_1725,N_1638,N_1609);
or U1726 (N_1726,N_1636,N_1625);
nor U1727 (N_1727,N_1631,N_1603);
or U1728 (N_1728,N_1675,N_1699);
and U1729 (N_1729,N_1698,N_1643);
and U1730 (N_1730,N_1679,N_1656);
or U1731 (N_1731,N_1678,N_1641);
nor U1732 (N_1732,N_1649,N_1685);
and U1733 (N_1733,N_1605,N_1697);
nand U1734 (N_1734,N_1647,N_1633);
and U1735 (N_1735,N_1680,N_1604);
xor U1736 (N_1736,N_1645,N_1612);
or U1737 (N_1737,N_1695,N_1624);
nor U1738 (N_1738,N_1694,N_1667);
nand U1739 (N_1739,N_1615,N_1651);
and U1740 (N_1740,N_1688,N_1683);
nor U1741 (N_1741,N_1692,N_1601);
and U1742 (N_1742,N_1646,N_1672);
and U1743 (N_1743,N_1681,N_1650);
and U1744 (N_1744,N_1662,N_1676);
xnor U1745 (N_1745,N_1614,N_1673);
nand U1746 (N_1746,N_1686,N_1693);
nor U1747 (N_1747,N_1623,N_1616);
xor U1748 (N_1748,N_1687,N_1665);
nor U1749 (N_1749,N_1682,N_1668);
nand U1750 (N_1750,N_1625,N_1641);
or U1751 (N_1751,N_1601,N_1691);
nor U1752 (N_1752,N_1608,N_1648);
nand U1753 (N_1753,N_1640,N_1605);
nor U1754 (N_1754,N_1627,N_1633);
nand U1755 (N_1755,N_1661,N_1619);
xnor U1756 (N_1756,N_1605,N_1637);
nand U1757 (N_1757,N_1600,N_1691);
and U1758 (N_1758,N_1656,N_1689);
and U1759 (N_1759,N_1604,N_1602);
nand U1760 (N_1760,N_1614,N_1643);
nor U1761 (N_1761,N_1657,N_1621);
or U1762 (N_1762,N_1658,N_1660);
and U1763 (N_1763,N_1625,N_1694);
and U1764 (N_1764,N_1621,N_1615);
nand U1765 (N_1765,N_1696,N_1606);
nor U1766 (N_1766,N_1680,N_1646);
and U1767 (N_1767,N_1626,N_1635);
xnor U1768 (N_1768,N_1622,N_1633);
and U1769 (N_1769,N_1602,N_1662);
and U1770 (N_1770,N_1637,N_1679);
and U1771 (N_1771,N_1614,N_1679);
nor U1772 (N_1772,N_1677,N_1690);
or U1773 (N_1773,N_1643,N_1692);
and U1774 (N_1774,N_1671,N_1638);
nand U1775 (N_1775,N_1687,N_1681);
or U1776 (N_1776,N_1666,N_1630);
nor U1777 (N_1777,N_1678,N_1601);
or U1778 (N_1778,N_1668,N_1674);
or U1779 (N_1779,N_1670,N_1644);
nor U1780 (N_1780,N_1610,N_1634);
and U1781 (N_1781,N_1679,N_1674);
nand U1782 (N_1782,N_1675,N_1680);
nor U1783 (N_1783,N_1629,N_1678);
and U1784 (N_1784,N_1651,N_1693);
and U1785 (N_1785,N_1698,N_1640);
nand U1786 (N_1786,N_1652,N_1660);
or U1787 (N_1787,N_1632,N_1661);
and U1788 (N_1788,N_1675,N_1640);
or U1789 (N_1789,N_1633,N_1691);
or U1790 (N_1790,N_1654,N_1660);
nand U1791 (N_1791,N_1619,N_1674);
xor U1792 (N_1792,N_1642,N_1664);
xor U1793 (N_1793,N_1602,N_1696);
and U1794 (N_1794,N_1666,N_1628);
nand U1795 (N_1795,N_1657,N_1697);
and U1796 (N_1796,N_1666,N_1602);
nor U1797 (N_1797,N_1653,N_1641);
and U1798 (N_1798,N_1626,N_1647);
nand U1799 (N_1799,N_1602,N_1663);
xnor U1800 (N_1800,N_1761,N_1720);
and U1801 (N_1801,N_1746,N_1732);
xnor U1802 (N_1802,N_1780,N_1769);
nor U1803 (N_1803,N_1730,N_1735);
nor U1804 (N_1804,N_1794,N_1710);
nor U1805 (N_1805,N_1701,N_1791);
nor U1806 (N_1806,N_1742,N_1762);
nand U1807 (N_1807,N_1733,N_1727);
or U1808 (N_1808,N_1707,N_1764);
xnor U1809 (N_1809,N_1771,N_1752);
nand U1810 (N_1810,N_1795,N_1728);
and U1811 (N_1811,N_1777,N_1750);
or U1812 (N_1812,N_1779,N_1766);
nand U1813 (N_1813,N_1745,N_1773);
nand U1814 (N_1814,N_1747,N_1703);
or U1815 (N_1815,N_1711,N_1799);
or U1816 (N_1816,N_1724,N_1778);
and U1817 (N_1817,N_1751,N_1709);
xnor U1818 (N_1818,N_1772,N_1700);
nand U1819 (N_1819,N_1785,N_1726);
nand U1820 (N_1820,N_1706,N_1797);
nand U1821 (N_1821,N_1790,N_1757);
xnor U1822 (N_1822,N_1725,N_1789);
or U1823 (N_1823,N_1774,N_1756);
or U1824 (N_1824,N_1718,N_1731);
xnor U1825 (N_1825,N_1719,N_1739);
nand U1826 (N_1826,N_1763,N_1759);
or U1827 (N_1827,N_1776,N_1737);
or U1828 (N_1828,N_1743,N_1741);
xor U1829 (N_1829,N_1765,N_1786);
nand U1830 (N_1830,N_1770,N_1715);
nand U1831 (N_1831,N_1721,N_1760);
and U1832 (N_1832,N_1784,N_1734);
and U1833 (N_1833,N_1792,N_1783);
nand U1834 (N_1834,N_1702,N_1708);
xor U1835 (N_1835,N_1753,N_1714);
nand U1836 (N_1836,N_1788,N_1781);
nor U1837 (N_1837,N_1767,N_1793);
and U1838 (N_1838,N_1740,N_1717);
and U1839 (N_1839,N_1744,N_1713);
and U1840 (N_1840,N_1705,N_1782);
nor U1841 (N_1841,N_1755,N_1736);
and U1842 (N_1842,N_1787,N_1754);
nand U1843 (N_1843,N_1729,N_1749);
nor U1844 (N_1844,N_1738,N_1704);
or U1845 (N_1845,N_1775,N_1716);
and U1846 (N_1846,N_1748,N_1768);
and U1847 (N_1847,N_1722,N_1758);
nand U1848 (N_1848,N_1723,N_1796);
nor U1849 (N_1849,N_1712,N_1798);
or U1850 (N_1850,N_1723,N_1746);
nand U1851 (N_1851,N_1795,N_1787);
and U1852 (N_1852,N_1781,N_1755);
xnor U1853 (N_1853,N_1722,N_1739);
nor U1854 (N_1854,N_1774,N_1734);
nor U1855 (N_1855,N_1770,N_1797);
nand U1856 (N_1856,N_1741,N_1764);
nor U1857 (N_1857,N_1702,N_1713);
or U1858 (N_1858,N_1706,N_1748);
nand U1859 (N_1859,N_1783,N_1746);
or U1860 (N_1860,N_1793,N_1730);
nor U1861 (N_1861,N_1730,N_1792);
nor U1862 (N_1862,N_1731,N_1711);
nor U1863 (N_1863,N_1741,N_1780);
nand U1864 (N_1864,N_1759,N_1798);
xor U1865 (N_1865,N_1717,N_1738);
xnor U1866 (N_1866,N_1733,N_1781);
or U1867 (N_1867,N_1713,N_1720);
nor U1868 (N_1868,N_1731,N_1759);
nand U1869 (N_1869,N_1789,N_1751);
nor U1870 (N_1870,N_1708,N_1780);
or U1871 (N_1871,N_1796,N_1774);
or U1872 (N_1872,N_1725,N_1780);
and U1873 (N_1873,N_1783,N_1748);
xnor U1874 (N_1874,N_1784,N_1742);
nand U1875 (N_1875,N_1776,N_1760);
or U1876 (N_1876,N_1727,N_1772);
nand U1877 (N_1877,N_1711,N_1741);
or U1878 (N_1878,N_1720,N_1702);
nor U1879 (N_1879,N_1741,N_1733);
nor U1880 (N_1880,N_1794,N_1759);
and U1881 (N_1881,N_1752,N_1732);
xor U1882 (N_1882,N_1747,N_1791);
nand U1883 (N_1883,N_1755,N_1775);
nand U1884 (N_1884,N_1780,N_1706);
nor U1885 (N_1885,N_1768,N_1744);
nand U1886 (N_1886,N_1751,N_1705);
nand U1887 (N_1887,N_1777,N_1795);
nand U1888 (N_1888,N_1745,N_1780);
and U1889 (N_1889,N_1761,N_1734);
or U1890 (N_1890,N_1777,N_1763);
or U1891 (N_1891,N_1757,N_1767);
nor U1892 (N_1892,N_1741,N_1726);
nand U1893 (N_1893,N_1784,N_1717);
xor U1894 (N_1894,N_1752,N_1764);
or U1895 (N_1895,N_1784,N_1704);
and U1896 (N_1896,N_1753,N_1794);
and U1897 (N_1897,N_1724,N_1719);
and U1898 (N_1898,N_1721,N_1782);
and U1899 (N_1899,N_1739,N_1703);
and U1900 (N_1900,N_1880,N_1855);
and U1901 (N_1901,N_1803,N_1846);
xnor U1902 (N_1902,N_1887,N_1856);
and U1903 (N_1903,N_1868,N_1832);
and U1904 (N_1904,N_1802,N_1892);
nor U1905 (N_1905,N_1828,N_1879);
or U1906 (N_1906,N_1869,N_1801);
nand U1907 (N_1907,N_1821,N_1889);
or U1908 (N_1908,N_1848,N_1805);
or U1909 (N_1909,N_1815,N_1891);
or U1910 (N_1910,N_1885,N_1837);
nor U1911 (N_1911,N_1864,N_1840);
or U1912 (N_1912,N_1820,N_1863);
and U1913 (N_1913,N_1852,N_1886);
and U1914 (N_1914,N_1861,N_1881);
nand U1915 (N_1915,N_1822,N_1862);
nand U1916 (N_1916,N_1808,N_1850);
nand U1917 (N_1917,N_1882,N_1829);
and U1918 (N_1918,N_1810,N_1831);
or U1919 (N_1919,N_1812,N_1898);
and U1920 (N_1920,N_1811,N_1841);
xnor U1921 (N_1921,N_1873,N_1899);
nand U1922 (N_1922,N_1858,N_1893);
and U1923 (N_1923,N_1872,N_1878);
nor U1924 (N_1924,N_1826,N_1884);
nor U1925 (N_1925,N_1895,N_1897);
or U1926 (N_1926,N_1871,N_1816);
nand U1927 (N_1927,N_1813,N_1827);
and U1928 (N_1928,N_1807,N_1875);
or U1929 (N_1929,N_1890,N_1835);
nor U1930 (N_1930,N_1847,N_1844);
nand U1931 (N_1931,N_1853,N_1870);
or U1932 (N_1932,N_1845,N_1888);
xnor U1933 (N_1933,N_1833,N_1883);
nand U1934 (N_1934,N_1854,N_1867);
or U1935 (N_1935,N_1896,N_1836);
xor U1936 (N_1936,N_1823,N_1834);
or U1937 (N_1937,N_1877,N_1843);
or U1938 (N_1938,N_1824,N_1866);
nand U1939 (N_1939,N_1849,N_1839);
nor U1940 (N_1940,N_1830,N_1819);
xor U1941 (N_1941,N_1814,N_1851);
nand U1942 (N_1942,N_1894,N_1876);
nand U1943 (N_1943,N_1838,N_1859);
nor U1944 (N_1944,N_1818,N_1857);
nand U1945 (N_1945,N_1874,N_1800);
nand U1946 (N_1946,N_1806,N_1825);
nand U1947 (N_1947,N_1842,N_1809);
or U1948 (N_1948,N_1865,N_1804);
nor U1949 (N_1949,N_1860,N_1817);
nand U1950 (N_1950,N_1836,N_1875);
or U1951 (N_1951,N_1868,N_1888);
and U1952 (N_1952,N_1817,N_1816);
nand U1953 (N_1953,N_1801,N_1896);
nand U1954 (N_1954,N_1883,N_1859);
nand U1955 (N_1955,N_1845,N_1819);
and U1956 (N_1956,N_1810,N_1863);
nor U1957 (N_1957,N_1839,N_1889);
nor U1958 (N_1958,N_1853,N_1896);
xnor U1959 (N_1959,N_1876,N_1810);
nor U1960 (N_1960,N_1893,N_1857);
and U1961 (N_1961,N_1815,N_1835);
and U1962 (N_1962,N_1885,N_1839);
xor U1963 (N_1963,N_1884,N_1831);
xnor U1964 (N_1964,N_1872,N_1846);
or U1965 (N_1965,N_1860,N_1825);
or U1966 (N_1966,N_1814,N_1805);
xnor U1967 (N_1967,N_1841,N_1839);
or U1968 (N_1968,N_1852,N_1833);
and U1969 (N_1969,N_1807,N_1833);
nand U1970 (N_1970,N_1811,N_1873);
nand U1971 (N_1971,N_1898,N_1892);
nor U1972 (N_1972,N_1828,N_1808);
nand U1973 (N_1973,N_1884,N_1804);
and U1974 (N_1974,N_1829,N_1861);
nor U1975 (N_1975,N_1827,N_1800);
and U1976 (N_1976,N_1894,N_1845);
and U1977 (N_1977,N_1870,N_1892);
nor U1978 (N_1978,N_1823,N_1847);
and U1979 (N_1979,N_1865,N_1809);
xor U1980 (N_1980,N_1892,N_1835);
nand U1981 (N_1981,N_1876,N_1889);
nor U1982 (N_1982,N_1848,N_1897);
nor U1983 (N_1983,N_1886,N_1885);
nand U1984 (N_1984,N_1859,N_1827);
nor U1985 (N_1985,N_1836,N_1881);
nand U1986 (N_1986,N_1884,N_1872);
and U1987 (N_1987,N_1851,N_1816);
nor U1988 (N_1988,N_1874,N_1883);
nor U1989 (N_1989,N_1851,N_1807);
or U1990 (N_1990,N_1842,N_1818);
and U1991 (N_1991,N_1846,N_1894);
or U1992 (N_1992,N_1857,N_1883);
and U1993 (N_1993,N_1835,N_1805);
or U1994 (N_1994,N_1888,N_1803);
nor U1995 (N_1995,N_1848,N_1803);
and U1996 (N_1996,N_1869,N_1867);
or U1997 (N_1997,N_1871,N_1886);
nand U1998 (N_1998,N_1878,N_1890);
or U1999 (N_1999,N_1889,N_1823);
nor U2000 (N_2000,N_1951,N_1989);
nand U2001 (N_2001,N_1983,N_1941);
nor U2002 (N_2002,N_1969,N_1986);
or U2003 (N_2003,N_1990,N_1996);
and U2004 (N_2004,N_1916,N_1909);
nor U2005 (N_2005,N_1977,N_1925);
xnor U2006 (N_2006,N_1964,N_1905);
xnor U2007 (N_2007,N_1952,N_1939);
nor U2008 (N_2008,N_1912,N_1999);
and U2009 (N_2009,N_1953,N_1934);
and U2010 (N_2010,N_1904,N_1943);
and U2011 (N_2011,N_1937,N_1921);
and U2012 (N_2012,N_1947,N_1928);
nor U2013 (N_2013,N_1998,N_1900);
xor U2014 (N_2014,N_1915,N_1973);
or U2015 (N_2015,N_1957,N_1902);
nor U2016 (N_2016,N_1945,N_1994);
nor U2017 (N_2017,N_1995,N_1929);
and U2018 (N_2018,N_1955,N_1931);
nor U2019 (N_2019,N_1903,N_1917);
xnor U2020 (N_2020,N_1993,N_1984);
xor U2021 (N_2021,N_1906,N_1944);
xor U2022 (N_2022,N_1997,N_1948);
or U2023 (N_2023,N_1914,N_1949);
nand U2024 (N_2024,N_1918,N_1959);
and U2025 (N_2025,N_1936,N_1942);
or U2026 (N_2026,N_1910,N_1975);
and U2027 (N_2027,N_1930,N_1935);
nor U2028 (N_2028,N_1981,N_1967);
and U2029 (N_2029,N_1924,N_1954);
nand U2030 (N_2030,N_1991,N_1985);
xor U2031 (N_2031,N_1923,N_1926);
or U2032 (N_2032,N_1982,N_1960);
nor U2033 (N_2033,N_1956,N_1938);
nand U2034 (N_2034,N_1976,N_1922);
nor U2035 (N_2035,N_1979,N_1911);
nor U2036 (N_2036,N_1919,N_1907);
xor U2037 (N_2037,N_1940,N_1988);
or U2038 (N_2038,N_1974,N_1978);
and U2039 (N_2039,N_1972,N_1913);
nand U2040 (N_2040,N_1950,N_1927);
nor U2041 (N_2041,N_1962,N_1933);
nor U2042 (N_2042,N_1992,N_1963);
nand U2043 (N_2043,N_1920,N_1980);
nand U2044 (N_2044,N_1965,N_1946);
nor U2045 (N_2045,N_1961,N_1932);
or U2046 (N_2046,N_1987,N_1901);
xor U2047 (N_2047,N_1971,N_1958);
xnor U2048 (N_2048,N_1908,N_1970);
or U2049 (N_2049,N_1966,N_1968);
nor U2050 (N_2050,N_1913,N_1944);
nand U2051 (N_2051,N_1950,N_1980);
or U2052 (N_2052,N_1975,N_1983);
nand U2053 (N_2053,N_1912,N_1976);
nand U2054 (N_2054,N_1929,N_1972);
and U2055 (N_2055,N_1903,N_1966);
and U2056 (N_2056,N_1980,N_1938);
or U2057 (N_2057,N_1944,N_1908);
or U2058 (N_2058,N_1971,N_1924);
and U2059 (N_2059,N_1904,N_1914);
xnor U2060 (N_2060,N_1997,N_1989);
nand U2061 (N_2061,N_1937,N_1994);
nand U2062 (N_2062,N_1931,N_1924);
and U2063 (N_2063,N_1947,N_1985);
or U2064 (N_2064,N_1991,N_1905);
or U2065 (N_2065,N_1984,N_1936);
nor U2066 (N_2066,N_1954,N_1996);
xnor U2067 (N_2067,N_1990,N_1910);
or U2068 (N_2068,N_1962,N_1945);
xor U2069 (N_2069,N_1994,N_1974);
or U2070 (N_2070,N_1996,N_1904);
and U2071 (N_2071,N_1963,N_1987);
and U2072 (N_2072,N_1952,N_1933);
nand U2073 (N_2073,N_1912,N_1980);
nand U2074 (N_2074,N_1990,N_1909);
nor U2075 (N_2075,N_1968,N_1915);
nor U2076 (N_2076,N_1987,N_1973);
and U2077 (N_2077,N_1932,N_1918);
xor U2078 (N_2078,N_1991,N_1938);
nor U2079 (N_2079,N_1933,N_1965);
nor U2080 (N_2080,N_1971,N_1964);
and U2081 (N_2081,N_1951,N_1907);
xor U2082 (N_2082,N_1942,N_1915);
nand U2083 (N_2083,N_1960,N_1902);
nand U2084 (N_2084,N_1996,N_1913);
or U2085 (N_2085,N_1917,N_1999);
and U2086 (N_2086,N_1940,N_1961);
and U2087 (N_2087,N_1905,N_1963);
xnor U2088 (N_2088,N_1970,N_1969);
xor U2089 (N_2089,N_1974,N_1933);
and U2090 (N_2090,N_1913,N_1993);
nor U2091 (N_2091,N_1947,N_1970);
and U2092 (N_2092,N_1976,N_1953);
or U2093 (N_2093,N_1975,N_1915);
or U2094 (N_2094,N_1946,N_1978);
or U2095 (N_2095,N_1983,N_1968);
nand U2096 (N_2096,N_1992,N_1951);
nor U2097 (N_2097,N_1983,N_1955);
nor U2098 (N_2098,N_1992,N_1944);
nand U2099 (N_2099,N_1992,N_1998);
nor U2100 (N_2100,N_2002,N_2005);
nand U2101 (N_2101,N_2073,N_2044);
nand U2102 (N_2102,N_2042,N_2035);
nand U2103 (N_2103,N_2037,N_2095);
and U2104 (N_2104,N_2015,N_2043);
or U2105 (N_2105,N_2077,N_2008);
nor U2106 (N_2106,N_2034,N_2093);
nand U2107 (N_2107,N_2084,N_2061);
nor U2108 (N_2108,N_2091,N_2089);
or U2109 (N_2109,N_2051,N_2083);
nand U2110 (N_2110,N_2020,N_2071);
nor U2111 (N_2111,N_2063,N_2070);
nor U2112 (N_2112,N_2009,N_2076);
xor U2113 (N_2113,N_2014,N_2012);
xor U2114 (N_2114,N_2048,N_2081);
xor U2115 (N_2115,N_2041,N_2033);
or U2116 (N_2116,N_2017,N_2056);
xor U2117 (N_2117,N_2052,N_2053);
nor U2118 (N_2118,N_2036,N_2040);
nand U2119 (N_2119,N_2062,N_2059);
nand U2120 (N_2120,N_2087,N_2075);
nand U2121 (N_2121,N_2025,N_2060);
nand U2122 (N_2122,N_2004,N_2039);
nand U2123 (N_2123,N_2047,N_2066);
or U2124 (N_2124,N_2068,N_2079);
and U2125 (N_2125,N_2003,N_2046);
and U2126 (N_2126,N_2023,N_2085);
nor U2127 (N_2127,N_2064,N_2054);
nand U2128 (N_2128,N_2080,N_2099);
nor U2129 (N_2129,N_2049,N_2058);
nor U2130 (N_2130,N_2018,N_2074);
nand U2131 (N_2131,N_2078,N_2098);
nand U2132 (N_2132,N_2072,N_2090);
and U2133 (N_2133,N_2045,N_2096);
nand U2134 (N_2134,N_2050,N_2057);
nor U2135 (N_2135,N_2097,N_2026);
or U2136 (N_2136,N_2030,N_2019);
nor U2137 (N_2137,N_2001,N_2088);
or U2138 (N_2138,N_2067,N_2055);
nand U2139 (N_2139,N_2094,N_2082);
or U2140 (N_2140,N_2086,N_2011);
and U2141 (N_2141,N_2069,N_2029);
or U2142 (N_2142,N_2027,N_2024);
and U2143 (N_2143,N_2092,N_2065);
nor U2144 (N_2144,N_2031,N_2010);
and U2145 (N_2145,N_2038,N_2006);
or U2146 (N_2146,N_2000,N_2016);
and U2147 (N_2147,N_2021,N_2032);
and U2148 (N_2148,N_2022,N_2013);
nor U2149 (N_2149,N_2028,N_2007);
nor U2150 (N_2150,N_2067,N_2014);
nor U2151 (N_2151,N_2052,N_2094);
nor U2152 (N_2152,N_2052,N_2050);
nand U2153 (N_2153,N_2072,N_2085);
nor U2154 (N_2154,N_2069,N_2021);
xor U2155 (N_2155,N_2016,N_2083);
and U2156 (N_2156,N_2050,N_2017);
xnor U2157 (N_2157,N_2085,N_2028);
nand U2158 (N_2158,N_2020,N_2067);
nor U2159 (N_2159,N_2083,N_2097);
or U2160 (N_2160,N_2016,N_2066);
and U2161 (N_2161,N_2057,N_2047);
nand U2162 (N_2162,N_2047,N_2076);
nor U2163 (N_2163,N_2045,N_2092);
or U2164 (N_2164,N_2041,N_2008);
and U2165 (N_2165,N_2019,N_2037);
nor U2166 (N_2166,N_2034,N_2081);
nand U2167 (N_2167,N_2060,N_2089);
and U2168 (N_2168,N_2003,N_2014);
or U2169 (N_2169,N_2090,N_2065);
and U2170 (N_2170,N_2087,N_2095);
nand U2171 (N_2171,N_2033,N_2066);
or U2172 (N_2172,N_2059,N_2003);
xnor U2173 (N_2173,N_2045,N_2084);
or U2174 (N_2174,N_2092,N_2095);
or U2175 (N_2175,N_2006,N_2024);
or U2176 (N_2176,N_2090,N_2084);
xnor U2177 (N_2177,N_2055,N_2097);
nor U2178 (N_2178,N_2090,N_2097);
nand U2179 (N_2179,N_2088,N_2011);
nand U2180 (N_2180,N_2030,N_2060);
nand U2181 (N_2181,N_2095,N_2051);
nor U2182 (N_2182,N_2058,N_2022);
nand U2183 (N_2183,N_2099,N_2009);
and U2184 (N_2184,N_2008,N_2063);
and U2185 (N_2185,N_2077,N_2097);
nor U2186 (N_2186,N_2002,N_2066);
or U2187 (N_2187,N_2034,N_2051);
nor U2188 (N_2188,N_2024,N_2017);
or U2189 (N_2189,N_2033,N_2024);
and U2190 (N_2190,N_2021,N_2006);
nor U2191 (N_2191,N_2080,N_2090);
or U2192 (N_2192,N_2058,N_2088);
nand U2193 (N_2193,N_2042,N_2068);
nand U2194 (N_2194,N_2012,N_2020);
and U2195 (N_2195,N_2011,N_2016);
nand U2196 (N_2196,N_2004,N_2040);
or U2197 (N_2197,N_2039,N_2094);
xor U2198 (N_2198,N_2086,N_2010);
nand U2199 (N_2199,N_2011,N_2079);
and U2200 (N_2200,N_2113,N_2195);
xor U2201 (N_2201,N_2128,N_2112);
xnor U2202 (N_2202,N_2147,N_2118);
nand U2203 (N_2203,N_2102,N_2188);
or U2204 (N_2204,N_2160,N_2194);
nor U2205 (N_2205,N_2121,N_2138);
nor U2206 (N_2206,N_2199,N_2175);
nand U2207 (N_2207,N_2124,N_2184);
nor U2208 (N_2208,N_2137,N_2198);
or U2209 (N_2209,N_2153,N_2176);
nor U2210 (N_2210,N_2130,N_2109);
and U2211 (N_2211,N_2142,N_2185);
and U2212 (N_2212,N_2151,N_2174);
and U2213 (N_2213,N_2107,N_2190);
and U2214 (N_2214,N_2155,N_2144);
nand U2215 (N_2215,N_2132,N_2187);
xnor U2216 (N_2216,N_2189,N_2161);
nand U2217 (N_2217,N_2149,N_2143);
or U2218 (N_2218,N_2179,N_2163);
nor U2219 (N_2219,N_2100,N_2114);
and U2220 (N_2220,N_2182,N_2191);
nand U2221 (N_2221,N_2192,N_2172);
nor U2222 (N_2222,N_2120,N_2145);
nor U2223 (N_2223,N_2186,N_2181);
nor U2224 (N_2224,N_2171,N_2125);
nand U2225 (N_2225,N_2183,N_2152);
and U2226 (N_2226,N_2111,N_2156);
or U2227 (N_2227,N_2164,N_2173);
nor U2228 (N_2228,N_2115,N_2140);
nand U2229 (N_2229,N_2178,N_2158);
and U2230 (N_2230,N_2131,N_2166);
and U2231 (N_2231,N_2197,N_2154);
nor U2232 (N_2232,N_2146,N_2134);
xnor U2233 (N_2233,N_2135,N_2127);
nand U2234 (N_2234,N_2157,N_2104);
nor U2235 (N_2235,N_2165,N_2169);
nor U2236 (N_2236,N_2148,N_2177);
xor U2237 (N_2237,N_2141,N_2116);
nor U2238 (N_2238,N_2136,N_2110);
nand U2239 (N_2239,N_2103,N_2193);
xnor U2240 (N_2240,N_2122,N_2126);
nand U2241 (N_2241,N_2108,N_2117);
nor U2242 (N_2242,N_2159,N_2119);
xnor U2243 (N_2243,N_2168,N_2106);
and U2244 (N_2244,N_2139,N_2105);
or U2245 (N_2245,N_2123,N_2167);
nor U2246 (N_2246,N_2101,N_2180);
xor U2247 (N_2247,N_2196,N_2133);
and U2248 (N_2248,N_2129,N_2150);
xnor U2249 (N_2249,N_2162,N_2170);
and U2250 (N_2250,N_2171,N_2139);
nor U2251 (N_2251,N_2182,N_2170);
nor U2252 (N_2252,N_2164,N_2195);
nor U2253 (N_2253,N_2105,N_2103);
nand U2254 (N_2254,N_2197,N_2106);
nor U2255 (N_2255,N_2185,N_2100);
or U2256 (N_2256,N_2193,N_2172);
or U2257 (N_2257,N_2119,N_2154);
nand U2258 (N_2258,N_2192,N_2114);
and U2259 (N_2259,N_2120,N_2130);
nor U2260 (N_2260,N_2155,N_2141);
or U2261 (N_2261,N_2152,N_2139);
and U2262 (N_2262,N_2173,N_2157);
xor U2263 (N_2263,N_2182,N_2143);
nor U2264 (N_2264,N_2174,N_2167);
nor U2265 (N_2265,N_2125,N_2193);
and U2266 (N_2266,N_2150,N_2187);
and U2267 (N_2267,N_2104,N_2166);
or U2268 (N_2268,N_2193,N_2154);
or U2269 (N_2269,N_2103,N_2107);
nor U2270 (N_2270,N_2107,N_2133);
or U2271 (N_2271,N_2165,N_2122);
or U2272 (N_2272,N_2141,N_2158);
xor U2273 (N_2273,N_2130,N_2104);
nand U2274 (N_2274,N_2172,N_2148);
or U2275 (N_2275,N_2158,N_2143);
and U2276 (N_2276,N_2131,N_2160);
or U2277 (N_2277,N_2197,N_2160);
nor U2278 (N_2278,N_2169,N_2124);
nand U2279 (N_2279,N_2195,N_2170);
nor U2280 (N_2280,N_2175,N_2124);
nor U2281 (N_2281,N_2107,N_2165);
nor U2282 (N_2282,N_2110,N_2188);
nand U2283 (N_2283,N_2164,N_2117);
nor U2284 (N_2284,N_2128,N_2115);
and U2285 (N_2285,N_2135,N_2122);
nand U2286 (N_2286,N_2191,N_2139);
nand U2287 (N_2287,N_2123,N_2194);
xnor U2288 (N_2288,N_2179,N_2132);
xnor U2289 (N_2289,N_2151,N_2117);
nor U2290 (N_2290,N_2175,N_2176);
nand U2291 (N_2291,N_2195,N_2160);
and U2292 (N_2292,N_2168,N_2185);
or U2293 (N_2293,N_2108,N_2184);
and U2294 (N_2294,N_2111,N_2113);
xnor U2295 (N_2295,N_2133,N_2174);
nor U2296 (N_2296,N_2121,N_2189);
and U2297 (N_2297,N_2128,N_2132);
nand U2298 (N_2298,N_2149,N_2102);
nand U2299 (N_2299,N_2187,N_2159);
or U2300 (N_2300,N_2299,N_2230);
nand U2301 (N_2301,N_2298,N_2284);
and U2302 (N_2302,N_2257,N_2244);
nand U2303 (N_2303,N_2231,N_2218);
xor U2304 (N_2304,N_2253,N_2229);
xnor U2305 (N_2305,N_2248,N_2208);
xnor U2306 (N_2306,N_2236,N_2201);
xnor U2307 (N_2307,N_2237,N_2245);
nor U2308 (N_2308,N_2275,N_2295);
nor U2309 (N_2309,N_2225,N_2289);
or U2310 (N_2310,N_2293,N_2222);
or U2311 (N_2311,N_2297,N_2249);
and U2312 (N_2312,N_2277,N_2261);
and U2313 (N_2313,N_2272,N_2203);
nand U2314 (N_2314,N_2264,N_2281);
or U2315 (N_2315,N_2221,N_2217);
and U2316 (N_2316,N_2287,N_2292);
and U2317 (N_2317,N_2274,N_2256);
or U2318 (N_2318,N_2279,N_2267);
and U2319 (N_2319,N_2210,N_2226);
nand U2320 (N_2320,N_2270,N_2276);
nand U2321 (N_2321,N_2202,N_2212);
nand U2322 (N_2322,N_2215,N_2265);
nand U2323 (N_2323,N_2250,N_2234);
or U2324 (N_2324,N_2241,N_2294);
and U2325 (N_2325,N_2204,N_2269);
or U2326 (N_2326,N_2296,N_2252);
and U2327 (N_2327,N_2238,N_2278);
nand U2328 (N_2328,N_2228,N_2227);
or U2329 (N_2329,N_2273,N_2235);
or U2330 (N_2330,N_2255,N_2239);
or U2331 (N_2331,N_2213,N_2266);
nand U2332 (N_2332,N_2219,N_2200);
or U2333 (N_2333,N_2286,N_2263);
nand U2334 (N_2334,N_2282,N_2209);
nor U2335 (N_2335,N_2268,N_2216);
and U2336 (N_2336,N_2240,N_2224);
nand U2337 (N_2337,N_2232,N_2211);
and U2338 (N_2338,N_2283,N_2280);
or U2339 (N_2339,N_2260,N_2243);
and U2340 (N_2340,N_2258,N_2291);
nand U2341 (N_2341,N_2290,N_2271);
or U2342 (N_2342,N_2262,N_2223);
nand U2343 (N_2343,N_2288,N_2242);
or U2344 (N_2344,N_2205,N_2251);
nand U2345 (N_2345,N_2247,N_2206);
nand U2346 (N_2346,N_2220,N_2214);
and U2347 (N_2347,N_2285,N_2207);
xnor U2348 (N_2348,N_2233,N_2259);
nand U2349 (N_2349,N_2246,N_2254);
and U2350 (N_2350,N_2227,N_2220);
or U2351 (N_2351,N_2249,N_2296);
nand U2352 (N_2352,N_2249,N_2232);
or U2353 (N_2353,N_2240,N_2277);
xnor U2354 (N_2354,N_2203,N_2200);
nand U2355 (N_2355,N_2271,N_2237);
or U2356 (N_2356,N_2216,N_2283);
and U2357 (N_2357,N_2284,N_2230);
and U2358 (N_2358,N_2217,N_2234);
or U2359 (N_2359,N_2256,N_2276);
or U2360 (N_2360,N_2252,N_2248);
or U2361 (N_2361,N_2285,N_2264);
nand U2362 (N_2362,N_2222,N_2294);
and U2363 (N_2363,N_2250,N_2210);
and U2364 (N_2364,N_2215,N_2263);
nand U2365 (N_2365,N_2270,N_2256);
nor U2366 (N_2366,N_2292,N_2247);
nor U2367 (N_2367,N_2232,N_2288);
or U2368 (N_2368,N_2229,N_2267);
nand U2369 (N_2369,N_2241,N_2209);
nand U2370 (N_2370,N_2272,N_2245);
nor U2371 (N_2371,N_2252,N_2257);
and U2372 (N_2372,N_2282,N_2215);
and U2373 (N_2373,N_2213,N_2222);
or U2374 (N_2374,N_2267,N_2231);
or U2375 (N_2375,N_2298,N_2236);
nand U2376 (N_2376,N_2288,N_2220);
nand U2377 (N_2377,N_2278,N_2204);
nand U2378 (N_2378,N_2256,N_2294);
nand U2379 (N_2379,N_2298,N_2215);
nor U2380 (N_2380,N_2238,N_2217);
nor U2381 (N_2381,N_2251,N_2203);
nor U2382 (N_2382,N_2270,N_2206);
or U2383 (N_2383,N_2231,N_2251);
and U2384 (N_2384,N_2225,N_2271);
xor U2385 (N_2385,N_2277,N_2283);
nand U2386 (N_2386,N_2233,N_2214);
nand U2387 (N_2387,N_2245,N_2273);
or U2388 (N_2388,N_2211,N_2203);
and U2389 (N_2389,N_2228,N_2209);
nand U2390 (N_2390,N_2281,N_2279);
nand U2391 (N_2391,N_2272,N_2220);
and U2392 (N_2392,N_2258,N_2261);
or U2393 (N_2393,N_2248,N_2280);
xnor U2394 (N_2394,N_2225,N_2209);
nand U2395 (N_2395,N_2221,N_2273);
nand U2396 (N_2396,N_2216,N_2262);
nand U2397 (N_2397,N_2230,N_2206);
or U2398 (N_2398,N_2208,N_2288);
nand U2399 (N_2399,N_2202,N_2278);
or U2400 (N_2400,N_2357,N_2330);
nor U2401 (N_2401,N_2395,N_2303);
nor U2402 (N_2402,N_2362,N_2387);
nor U2403 (N_2403,N_2397,N_2339);
nor U2404 (N_2404,N_2353,N_2358);
or U2405 (N_2405,N_2315,N_2342);
and U2406 (N_2406,N_2329,N_2371);
nand U2407 (N_2407,N_2327,N_2369);
or U2408 (N_2408,N_2352,N_2302);
and U2409 (N_2409,N_2365,N_2321);
and U2410 (N_2410,N_2335,N_2318);
nand U2411 (N_2411,N_2322,N_2364);
and U2412 (N_2412,N_2394,N_2307);
and U2413 (N_2413,N_2382,N_2319);
and U2414 (N_2414,N_2366,N_2381);
or U2415 (N_2415,N_2347,N_2363);
or U2416 (N_2416,N_2309,N_2323);
and U2417 (N_2417,N_2338,N_2390);
or U2418 (N_2418,N_2380,N_2379);
or U2419 (N_2419,N_2310,N_2348);
and U2420 (N_2420,N_2367,N_2350);
nand U2421 (N_2421,N_2372,N_2361);
and U2422 (N_2422,N_2317,N_2328);
and U2423 (N_2423,N_2332,N_2378);
and U2424 (N_2424,N_2393,N_2313);
xnor U2425 (N_2425,N_2396,N_2311);
xnor U2426 (N_2426,N_2391,N_2370);
nor U2427 (N_2427,N_2392,N_2354);
or U2428 (N_2428,N_2334,N_2373);
or U2429 (N_2429,N_2356,N_2388);
or U2430 (N_2430,N_2337,N_2377);
or U2431 (N_2431,N_2341,N_2320);
nor U2432 (N_2432,N_2389,N_2340);
and U2433 (N_2433,N_2344,N_2312);
xnor U2434 (N_2434,N_2305,N_2324);
nand U2435 (N_2435,N_2336,N_2306);
or U2436 (N_2436,N_2374,N_2301);
and U2437 (N_2437,N_2349,N_2304);
nand U2438 (N_2438,N_2314,N_2375);
or U2439 (N_2439,N_2331,N_2351);
nor U2440 (N_2440,N_2360,N_2399);
and U2441 (N_2441,N_2326,N_2343);
xnor U2442 (N_2442,N_2368,N_2355);
or U2443 (N_2443,N_2385,N_2300);
and U2444 (N_2444,N_2398,N_2316);
nand U2445 (N_2445,N_2383,N_2376);
nor U2446 (N_2446,N_2346,N_2386);
or U2447 (N_2447,N_2345,N_2333);
or U2448 (N_2448,N_2384,N_2308);
and U2449 (N_2449,N_2359,N_2325);
or U2450 (N_2450,N_2314,N_2368);
xnor U2451 (N_2451,N_2373,N_2332);
nand U2452 (N_2452,N_2365,N_2389);
nor U2453 (N_2453,N_2395,N_2381);
nor U2454 (N_2454,N_2391,N_2392);
nor U2455 (N_2455,N_2364,N_2341);
or U2456 (N_2456,N_2329,N_2309);
and U2457 (N_2457,N_2326,N_2350);
nor U2458 (N_2458,N_2359,N_2389);
nor U2459 (N_2459,N_2372,N_2340);
and U2460 (N_2460,N_2327,N_2356);
and U2461 (N_2461,N_2344,N_2366);
nand U2462 (N_2462,N_2367,N_2338);
nor U2463 (N_2463,N_2353,N_2374);
nand U2464 (N_2464,N_2307,N_2315);
nand U2465 (N_2465,N_2327,N_2357);
or U2466 (N_2466,N_2369,N_2356);
or U2467 (N_2467,N_2324,N_2343);
or U2468 (N_2468,N_2301,N_2366);
xor U2469 (N_2469,N_2351,N_2396);
and U2470 (N_2470,N_2357,N_2335);
nor U2471 (N_2471,N_2337,N_2378);
xnor U2472 (N_2472,N_2303,N_2341);
and U2473 (N_2473,N_2367,N_2377);
xnor U2474 (N_2474,N_2359,N_2353);
nor U2475 (N_2475,N_2336,N_2370);
or U2476 (N_2476,N_2383,N_2357);
and U2477 (N_2477,N_2392,N_2311);
and U2478 (N_2478,N_2335,N_2302);
nand U2479 (N_2479,N_2363,N_2384);
and U2480 (N_2480,N_2331,N_2339);
and U2481 (N_2481,N_2390,N_2381);
nor U2482 (N_2482,N_2386,N_2371);
and U2483 (N_2483,N_2391,N_2372);
nor U2484 (N_2484,N_2319,N_2368);
or U2485 (N_2485,N_2329,N_2393);
nand U2486 (N_2486,N_2306,N_2366);
xor U2487 (N_2487,N_2322,N_2392);
nand U2488 (N_2488,N_2377,N_2386);
and U2489 (N_2489,N_2332,N_2390);
or U2490 (N_2490,N_2323,N_2327);
nor U2491 (N_2491,N_2338,N_2391);
nor U2492 (N_2492,N_2325,N_2386);
xnor U2493 (N_2493,N_2360,N_2304);
and U2494 (N_2494,N_2369,N_2324);
nor U2495 (N_2495,N_2322,N_2344);
nor U2496 (N_2496,N_2397,N_2379);
nand U2497 (N_2497,N_2327,N_2350);
or U2498 (N_2498,N_2343,N_2304);
xor U2499 (N_2499,N_2393,N_2368);
nor U2500 (N_2500,N_2451,N_2435);
or U2501 (N_2501,N_2460,N_2446);
and U2502 (N_2502,N_2401,N_2470);
and U2503 (N_2503,N_2466,N_2491);
xnor U2504 (N_2504,N_2452,N_2437);
and U2505 (N_2505,N_2480,N_2440);
nor U2506 (N_2506,N_2422,N_2476);
nand U2507 (N_2507,N_2405,N_2485);
or U2508 (N_2508,N_2434,N_2493);
and U2509 (N_2509,N_2431,N_2445);
and U2510 (N_2510,N_2455,N_2478);
and U2511 (N_2511,N_2436,N_2459);
and U2512 (N_2512,N_2461,N_2468);
nor U2513 (N_2513,N_2462,N_2419);
or U2514 (N_2514,N_2417,N_2463);
or U2515 (N_2515,N_2499,N_2426);
and U2516 (N_2516,N_2424,N_2494);
and U2517 (N_2517,N_2406,N_2409);
and U2518 (N_2518,N_2475,N_2400);
nand U2519 (N_2519,N_2448,N_2486);
xor U2520 (N_2520,N_2418,N_2489);
nand U2521 (N_2521,N_2414,N_2439);
and U2522 (N_2522,N_2428,N_2433);
or U2523 (N_2523,N_2427,N_2420);
xnor U2524 (N_2524,N_2444,N_2438);
or U2525 (N_2525,N_2410,N_2496);
nand U2526 (N_2526,N_2487,N_2492);
nand U2527 (N_2527,N_2425,N_2472);
or U2528 (N_2528,N_2495,N_2477);
and U2529 (N_2529,N_2423,N_2415);
and U2530 (N_2530,N_2408,N_2416);
or U2531 (N_2531,N_2484,N_2488);
nand U2532 (N_2532,N_2442,N_2411);
nor U2533 (N_2533,N_2421,N_2490);
xor U2534 (N_2534,N_2407,N_2402);
nor U2535 (N_2535,N_2412,N_2447);
and U2536 (N_2536,N_2498,N_2429);
nand U2537 (N_2537,N_2473,N_2474);
or U2538 (N_2538,N_2441,N_2449);
nand U2539 (N_2539,N_2457,N_2456);
and U2540 (N_2540,N_2481,N_2482);
or U2541 (N_2541,N_2479,N_2465);
and U2542 (N_2542,N_2467,N_2469);
nand U2543 (N_2543,N_2432,N_2413);
and U2544 (N_2544,N_2404,N_2430);
nand U2545 (N_2545,N_2464,N_2443);
nand U2546 (N_2546,N_2483,N_2471);
nor U2547 (N_2547,N_2497,N_2403);
or U2548 (N_2548,N_2454,N_2458);
nand U2549 (N_2549,N_2450,N_2453);
or U2550 (N_2550,N_2414,N_2464);
and U2551 (N_2551,N_2459,N_2458);
nand U2552 (N_2552,N_2432,N_2423);
nor U2553 (N_2553,N_2420,N_2459);
nor U2554 (N_2554,N_2419,N_2471);
nor U2555 (N_2555,N_2480,N_2402);
nor U2556 (N_2556,N_2434,N_2400);
and U2557 (N_2557,N_2473,N_2416);
or U2558 (N_2558,N_2483,N_2430);
nor U2559 (N_2559,N_2494,N_2432);
or U2560 (N_2560,N_2435,N_2486);
nand U2561 (N_2561,N_2494,N_2473);
or U2562 (N_2562,N_2473,N_2450);
and U2563 (N_2563,N_2470,N_2463);
nor U2564 (N_2564,N_2467,N_2476);
nor U2565 (N_2565,N_2439,N_2406);
xnor U2566 (N_2566,N_2487,N_2402);
nor U2567 (N_2567,N_2484,N_2416);
and U2568 (N_2568,N_2425,N_2446);
xnor U2569 (N_2569,N_2414,N_2460);
and U2570 (N_2570,N_2451,N_2409);
nand U2571 (N_2571,N_2415,N_2458);
nand U2572 (N_2572,N_2408,N_2437);
or U2573 (N_2573,N_2400,N_2401);
or U2574 (N_2574,N_2431,N_2402);
nand U2575 (N_2575,N_2419,N_2444);
nand U2576 (N_2576,N_2432,N_2417);
or U2577 (N_2577,N_2413,N_2464);
or U2578 (N_2578,N_2483,N_2490);
nand U2579 (N_2579,N_2423,N_2442);
or U2580 (N_2580,N_2484,N_2475);
nor U2581 (N_2581,N_2419,N_2412);
nor U2582 (N_2582,N_2419,N_2448);
xor U2583 (N_2583,N_2473,N_2481);
and U2584 (N_2584,N_2421,N_2477);
or U2585 (N_2585,N_2421,N_2485);
nor U2586 (N_2586,N_2417,N_2409);
or U2587 (N_2587,N_2432,N_2478);
or U2588 (N_2588,N_2484,N_2470);
xnor U2589 (N_2589,N_2489,N_2425);
nand U2590 (N_2590,N_2445,N_2402);
and U2591 (N_2591,N_2450,N_2482);
nand U2592 (N_2592,N_2401,N_2476);
nand U2593 (N_2593,N_2428,N_2458);
nand U2594 (N_2594,N_2426,N_2427);
and U2595 (N_2595,N_2419,N_2498);
nand U2596 (N_2596,N_2443,N_2403);
nor U2597 (N_2597,N_2447,N_2489);
and U2598 (N_2598,N_2444,N_2439);
nand U2599 (N_2599,N_2425,N_2427);
xor U2600 (N_2600,N_2583,N_2565);
nand U2601 (N_2601,N_2586,N_2574);
nand U2602 (N_2602,N_2510,N_2503);
xnor U2603 (N_2603,N_2525,N_2555);
nand U2604 (N_2604,N_2560,N_2504);
nand U2605 (N_2605,N_2506,N_2522);
and U2606 (N_2606,N_2571,N_2532);
nor U2607 (N_2607,N_2584,N_2569);
nor U2608 (N_2608,N_2592,N_2597);
nor U2609 (N_2609,N_2577,N_2579);
and U2610 (N_2610,N_2502,N_2538);
nand U2611 (N_2611,N_2553,N_2527);
nand U2612 (N_2612,N_2582,N_2549);
and U2613 (N_2613,N_2585,N_2546);
xnor U2614 (N_2614,N_2562,N_2517);
nor U2615 (N_2615,N_2540,N_2543);
nor U2616 (N_2616,N_2594,N_2590);
or U2617 (N_2617,N_2530,N_2593);
or U2618 (N_2618,N_2533,N_2535);
and U2619 (N_2619,N_2598,N_2575);
and U2620 (N_2620,N_2531,N_2580);
nand U2621 (N_2621,N_2544,N_2509);
and U2622 (N_2622,N_2542,N_2558);
nand U2623 (N_2623,N_2550,N_2576);
nor U2624 (N_2624,N_2591,N_2514);
nand U2625 (N_2625,N_2568,N_2528);
or U2626 (N_2626,N_2578,N_2547);
and U2627 (N_2627,N_2519,N_2552);
and U2628 (N_2628,N_2507,N_2539);
nor U2629 (N_2629,N_2567,N_2520);
and U2630 (N_2630,N_2511,N_2566);
nor U2631 (N_2631,N_2554,N_2518);
nand U2632 (N_2632,N_2524,N_2572);
nor U2633 (N_2633,N_2573,N_2599);
or U2634 (N_2634,N_2563,N_2537);
or U2635 (N_2635,N_2551,N_2541);
nor U2636 (N_2636,N_2512,N_2501);
and U2637 (N_2637,N_2534,N_2523);
or U2638 (N_2638,N_2513,N_2559);
nor U2639 (N_2639,N_2589,N_2545);
or U2640 (N_2640,N_2596,N_2595);
nor U2641 (N_2641,N_2548,N_2526);
nand U2642 (N_2642,N_2515,N_2564);
xnor U2643 (N_2643,N_2508,N_2588);
and U2644 (N_2644,N_2536,N_2557);
nor U2645 (N_2645,N_2570,N_2556);
or U2646 (N_2646,N_2561,N_2500);
and U2647 (N_2647,N_2529,N_2505);
nand U2648 (N_2648,N_2587,N_2521);
and U2649 (N_2649,N_2581,N_2516);
or U2650 (N_2650,N_2507,N_2531);
and U2651 (N_2651,N_2547,N_2585);
nand U2652 (N_2652,N_2566,N_2544);
or U2653 (N_2653,N_2542,N_2535);
nand U2654 (N_2654,N_2502,N_2504);
and U2655 (N_2655,N_2591,N_2573);
nor U2656 (N_2656,N_2505,N_2526);
nand U2657 (N_2657,N_2550,N_2528);
nand U2658 (N_2658,N_2580,N_2514);
and U2659 (N_2659,N_2552,N_2503);
and U2660 (N_2660,N_2563,N_2551);
nand U2661 (N_2661,N_2505,N_2558);
nor U2662 (N_2662,N_2540,N_2592);
xor U2663 (N_2663,N_2559,N_2587);
nor U2664 (N_2664,N_2559,N_2500);
nand U2665 (N_2665,N_2527,N_2575);
nand U2666 (N_2666,N_2598,N_2549);
nand U2667 (N_2667,N_2503,N_2590);
nand U2668 (N_2668,N_2560,N_2558);
nor U2669 (N_2669,N_2582,N_2599);
nand U2670 (N_2670,N_2529,N_2546);
and U2671 (N_2671,N_2506,N_2570);
nand U2672 (N_2672,N_2528,N_2595);
nand U2673 (N_2673,N_2538,N_2532);
and U2674 (N_2674,N_2555,N_2577);
xor U2675 (N_2675,N_2553,N_2562);
and U2676 (N_2676,N_2502,N_2560);
nand U2677 (N_2677,N_2551,N_2522);
nor U2678 (N_2678,N_2557,N_2527);
or U2679 (N_2679,N_2592,N_2583);
and U2680 (N_2680,N_2577,N_2521);
or U2681 (N_2681,N_2520,N_2575);
and U2682 (N_2682,N_2514,N_2572);
nor U2683 (N_2683,N_2548,N_2554);
or U2684 (N_2684,N_2547,N_2500);
or U2685 (N_2685,N_2526,N_2509);
nand U2686 (N_2686,N_2569,N_2587);
nor U2687 (N_2687,N_2515,N_2581);
nand U2688 (N_2688,N_2502,N_2527);
and U2689 (N_2689,N_2574,N_2513);
xor U2690 (N_2690,N_2569,N_2533);
and U2691 (N_2691,N_2560,N_2585);
nand U2692 (N_2692,N_2524,N_2542);
and U2693 (N_2693,N_2576,N_2501);
nand U2694 (N_2694,N_2557,N_2517);
and U2695 (N_2695,N_2537,N_2524);
nor U2696 (N_2696,N_2555,N_2543);
or U2697 (N_2697,N_2507,N_2526);
nor U2698 (N_2698,N_2539,N_2544);
and U2699 (N_2699,N_2534,N_2579);
or U2700 (N_2700,N_2605,N_2692);
nor U2701 (N_2701,N_2667,N_2656);
nor U2702 (N_2702,N_2653,N_2641);
and U2703 (N_2703,N_2625,N_2633);
xor U2704 (N_2704,N_2612,N_2621);
and U2705 (N_2705,N_2699,N_2663);
or U2706 (N_2706,N_2690,N_2662);
and U2707 (N_2707,N_2639,N_2674);
xnor U2708 (N_2708,N_2647,N_2638);
or U2709 (N_2709,N_2617,N_2623);
or U2710 (N_2710,N_2697,N_2686);
and U2711 (N_2711,N_2644,N_2635);
nor U2712 (N_2712,N_2630,N_2670);
or U2713 (N_2713,N_2637,N_2676);
xor U2714 (N_2714,N_2618,N_2616);
nand U2715 (N_2715,N_2679,N_2643);
nor U2716 (N_2716,N_2603,N_2626);
or U2717 (N_2717,N_2660,N_2677);
and U2718 (N_2718,N_2684,N_2610);
nor U2719 (N_2719,N_2646,N_2600);
nor U2720 (N_2720,N_2666,N_2675);
or U2721 (N_2721,N_2614,N_2624);
nand U2722 (N_2722,N_2659,N_2628);
and U2723 (N_2723,N_2608,N_2652);
nor U2724 (N_2724,N_2678,N_2627);
nand U2725 (N_2725,N_2665,N_2622);
nor U2726 (N_2726,N_2604,N_2658);
nor U2727 (N_2727,N_2668,N_2629);
and U2728 (N_2728,N_2654,N_2619);
or U2729 (N_2729,N_2671,N_2680);
or U2730 (N_2730,N_2689,N_2613);
or U2731 (N_2731,N_2645,N_2601);
nand U2732 (N_2732,N_2682,N_2651);
or U2733 (N_2733,N_2606,N_2669);
and U2734 (N_2734,N_2640,N_2681);
nor U2735 (N_2735,N_2602,N_2649);
xor U2736 (N_2736,N_2650,N_2688);
and U2737 (N_2737,N_2636,N_2632);
nand U2738 (N_2738,N_2696,N_2611);
or U2739 (N_2739,N_2655,N_2693);
xor U2740 (N_2740,N_2620,N_2631);
or U2741 (N_2741,N_2673,N_2685);
and U2742 (N_2742,N_2664,N_2694);
nor U2743 (N_2743,N_2648,N_2698);
nand U2744 (N_2744,N_2642,N_2661);
or U2745 (N_2745,N_2615,N_2695);
xnor U2746 (N_2746,N_2657,N_2687);
nor U2747 (N_2747,N_2607,N_2672);
and U2748 (N_2748,N_2683,N_2634);
or U2749 (N_2749,N_2691,N_2609);
and U2750 (N_2750,N_2618,N_2655);
and U2751 (N_2751,N_2656,N_2686);
xnor U2752 (N_2752,N_2650,N_2685);
nand U2753 (N_2753,N_2646,N_2640);
nand U2754 (N_2754,N_2654,N_2652);
and U2755 (N_2755,N_2624,N_2673);
nor U2756 (N_2756,N_2613,N_2635);
or U2757 (N_2757,N_2678,N_2697);
or U2758 (N_2758,N_2655,N_2620);
or U2759 (N_2759,N_2685,N_2617);
nor U2760 (N_2760,N_2666,N_2649);
and U2761 (N_2761,N_2658,N_2654);
or U2762 (N_2762,N_2648,N_2604);
nor U2763 (N_2763,N_2625,N_2664);
nor U2764 (N_2764,N_2644,N_2684);
nand U2765 (N_2765,N_2681,N_2680);
or U2766 (N_2766,N_2672,N_2601);
nand U2767 (N_2767,N_2633,N_2631);
nor U2768 (N_2768,N_2610,N_2642);
xnor U2769 (N_2769,N_2665,N_2647);
nor U2770 (N_2770,N_2655,N_2650);
xnor U2771 (N_2771,N_2625,N_2618);
or U2772 (N_2772,N_2610,N_2694);
xor U2773 (N_2773,N_2656,N_2685);
and U2774 (N_2774,N_2673,N_2691);
and U2775 (N_2775,N_2618,N_2658);
and U2776 (N_2776,N_2630,N_2616);
nand U2777 (N_2777,N_2695,N_2652);
nor U2778 (N_2778,N_2630,N_2680);
nor U2779 (N_2779,N_2630,N_2626);
and U2780 (N_2780,N_2665,N_2693);
nand U2781 (N_2781,N_2684,N_2681);
nor U2782 (N_2782,N_2635,N_2657);
or U2783 (N_2783,N_2606,N_2661);
nor U2784 (N_2784,N_2693,N_2634);
xor U2785 (N_2785,N_2694,N_2619);
nand U2786 (N_2786,N_2651,N_2655);
nor U2787 (N_2787,N_2699,N_2683);
nand U2788 (N_2788,N_2682,N_2698);
and U2789 (N_2789,N_2627,N_2658);
or U2790 (N_2790,N_2633,N_2673);
or U2791 (N_2791,N_2630,N_2696);
nand U2792 (N_2792,N_2660,N_2639);
nor U2793 (N_2793,N_2637,N_2647);
nand U2794 (N_2794,N_2673,N_2605);
nand U2795 (N_2795,N_2664,N_2693);
or U2796 (N_2796,N_2655,N_2601);
or U2797 (N_2797,N_2646,N_2656);
nor U2798 (N_2798,N_2638,N_2601);
nand U2799 (N_2799,N_2699,N_2635);
nor U2800 (N_2800,N_2728,N_2735);
nor U2801 (N_2801,N_2727,N_2712);
nor U2802 (N_2802,N_2781,N_2782);
and U2803 (N_2803,N_2787,N_2799);
and U2804 (N_2804,N_2706,N_2731);
and U2805 (N_2805,N_2790,N_2736);
xor U2806 (N_2806,N_2777,N_2778);
or U2807 (N_2807,N_2761,N_2769);
or U2808 (N_2808,N_2793,N_2776);
nor U2809 (N_2809,N_2708,N_2742);
nor U2810 (N_2810,N_2700,N_2709);
nor U2811 (N_2811,N_2744,N_2798);
and U2812 (N_2812,N_2738,N_2713);
nand U2813 (N_2813,N_2703,N_2704);
and U2814 (N_2814,N_2737,N_2760);
nor U2815 (N_2815,N_2711,N_2755);
or U2816 (N_2816,N_2789,N_2734);
nor U2817 (N_2817,N_2741,N_2785);
nor U2818 (N_2818,N_2774,N_2796);
nor U2819 (N_2819,N_2717,N_2795);
and U2820 (N_2820,N_2783,N_2743);
nand U2821 (N_2821,N_2716,N_2752);
nand U2822 (N_2822,N_2748,N_2718);
nand U2823 (N_2823,N_2722,N_2732);
nor U2824 (N_2824,N_2715,N_2773);
and U2825 (N_2825,N_2719,N_2756);
nor U2826 (N_2826,N_2775,N_2750);
nor U2827 (N_2827,N_2771,N_2786);
nand U2828 (N_2828,N_2725,N_2762);
nor U2829 (N_2829,N_2733,N_2747);
or U2830 (N_2830,N_2739,N_2751);
and U2831 (N_2831,N_2740,N_2745);
nor U2832 (N_2832,N_2792,N_2726);
and U2833 (N_2833,N_2705,N_2720);
nand U2834 (N_2834,N_2758,N_2721);
and U2835 (N_2835,N_2757,N_2754);
nor U2836 (N_2836,N_2763,N_2730);
or U2837 (N_2837,N_2765,N_2780);
and U2838 (N_2838,N_2788,N_2707);
xor U2839 (N_2839,N_2701,N_2723);
or U2840 (N_2840,N_2710,N_2729);
xor U2841 (N_2841,N_2772,N_2784);
and U2842 (N_2842,N_2779,N_2797);
xnor U2843 (N_2843,N_2764,N_2767);
and U2844 (N_2844,N_2759,N_2702);
or U2845 (N_2845,N_2714,N_2768);
and U2846 (N_2846,N_2753,N_2749);
nand U2847 (N_2847,N_2724,N_2794);
or U2848 (N_2848,N_2770,N_2746);
nor U2849 (N_2849,N_2766,N_2791);
nand U2850 (N_2850,N_2746,N_2742);
or U2851 (N_2851,N_2786,N_2779);
nor U2852 (N_2852,N_2713,N_2782);
nand U2853 (N_2853,N_2721,N_2772);
and U2854 (N_2854,N_2768,N_2755);
nand U2855 (N_2855,N_2779,N_2790);
nor U2856 (N_2856,N_2707,N_2757);
and U2857 (N_2857,N_2739,N_2723);
and U2858 (N_2858,N_2785,N_2758);
or U2859 (N_2859,N_2759,N_2732);
or U2860 (N_2860,N_2734,N_2750);
nand U2861 (N_2861,N_2772,N_2780);
nand U2862 (N_2862,N_2751,N_2723);
nor U2863 (N_2863,N_2727,N_2771);
and U2864 (N_2864,N_2710,N_2786);
or U2865 (N_2865,N_2792,N_2782);
nor U2866 (N_2866,N_2779,N_2787);
nor U2867 (N_2867,N_2771,N_2762);
nand U2868 (N_2868,N_2770,N_2786);
nor U2869 (N_2869,N_2744,N_2706);
nor U2870 (N_2870,N_2712,N_2789);
or U2871 (N_2871,N_2773,N_2792);
nor U2872 (N_2872,N_2722,N_2712);
xor U2873 (N_2873,N_2722,N_2713);
nand U2874 (N_2874,N_2779,N_2702);
or U2875 (N_2875,N_2789,N_2792);
and U2876 (N_2876,N_2725,N_2731);
nor U2877 (N_2877,N_2709,N_2799);
nand U2878 (N_2878,N_2762,N_2734);
and U2879 (N_2879,N_2796,N_2799);
xor U2880 (N_2880,N_2762,N_2727);
nand U2881 (N_2881,N_2759,N_2735);
or U2882 (N_2882,N_2793,N_2722);
and U2883 (N_2883,N_2744,N_2762);
nand U2884 (N_2884,N_2763,N_2720);
or U2885 (N_2885,N_2711,N_2745);
and U2886 (N_2886,N_2769,N_2765);
or U2887 (N_2887,N_2785,N_2781);
nor U2888 (N_2888,N_2775,N_2741);
or U2889 (N_2889,N_2748,N_2787);
or U2890 (N_2890,N_2750,N_2727);
and U2891 (N_2891,N_2733,N_2777);
nor U2892 (N_2892,N_2761,N_2764);
or U2893 (N_2893,N_2799,N_2757);
nand U2894 (N_2894,N_2771,N_2767);
or U2895 (N_2895,N_2743,N_2714);
nand U2896 (N_2896,N_2765,N_2753);
and U2897 (N_2897,N_2726,N_2738);
nor U2898 (N_2898,N_2747,N_2741);
nor U2899 (N_2899,N_2787,N_2766);
or U2900 (N_2900,N_2841,N_2893);
or U2901 (N_2901,N_2828,N_2805);
and U2902 (N_2902,N_2819,N_2861);
or U2903 (N_2903,N_2800,N_2886);
nand U2904 (N_2904,N_2826,N_2847);
nor U2905 (N_2905,N_2843,N_2870);
and U2906 (N_2906,N_2834,N_2890);
and U2907 (N_2907,N_2860,N_2806);
or U2908 (N_2908,N_2888,N_2863);
nand U2909 (N_2909,N_2894,N_2885);
and U2910 (N_2910,N_2812,N_2840);
nor U2911 (N_2911,N_2884,N_2831);
nand U2912 (N_2912,N_2803,N_2830);
or U2913 (N_2913,N_2877,N_2839);
or U2914 (N_2914,N_2876,N_2898);
and U2915 (N_2915,N_2856,N_2801);
nand U2916 (N_2916,N_2899,N_2837);
nand U2917 (N_2917,N_2807,N_2857);
nand U2918 (N_2918,N_2848,N_2845);
or U2919 (N_2919,N_2859,N_2862);
nor U2920 (N_2920,N_2833,N_2846);
nand U2921 (N_2921,N_2897,N_2891);
nand U2922 (N_2922,N_2866,N_2882);
nor U2923 (N_2923,N_2896,N_2864);
and U2924 (N_2924,N_2869,N_2850);
nand U2925 (N_2925,N_2842,N_2849);
xnor U2926 (N_2926,N_2851,N_2804);
nand U2927 (N_2927,N_2810,N_2871);
nand U2928 (N_2928,N_2817,N_2844);
or U2929 (N_2929,N_2824,N_2821);
nor U2930 (N_2930,N_2820,N_2808);
or U2931 (N_2931,N_2818,N_2878);
or U2932 (N_2932,N_2868,N_2892);
and U2933 (N_2933,N_2813,N_2865);
or U2934 (N_2934,N_2838,N_2874);
and U2935 (N_2935,N_2836,N_2809);
and U2936 (N_2936,N_2811,N_2822);
nor U2937 (N_2937,N_2835,N_2875);
and U2938 (N_2938,N_2852,N_2802);
nand U2939 (N_2939,N_2895,N_2887);
and U2940 (N_2940,N_2816,N_2815);
or U2941 (N_2941,N_2829,N_2855);
and U2942 (N_2942,N_2832,N_2879);
and U2943 (N_2943,N_2854,N_2823);
nor U2944 (N_2944,N_2889,N_2872);
nand U2945 (N_2945,N_2883,N_2881);
nand U2946 (N_2946,N_2853,N_2858);
and U2947 (N_2947,N_2825,N_2814);
nand U2948 (N_2948,N_2827,N_2873);
nand U2949 (N_2949,N_2867,N_2880);
xor U2950 (N_2950,N_2845,N_2830);
and U2951 (N_2951,N_2877,N_2872);
nand U2952 (N_2952,N_2866,N_2861);
and U2953 (N_2953,N_2889,N_2830);
nor U2954 (N_2954,N_2858,N_2872);
xor U2955 (N_2955,N_2849,N_2854);
or U2956 (N_2956,N_2859,N_2876);
nor U2957 (N_2957,N_2853,N_2841);
nor U2958 (N_2958,N_2837,N_2867);
nand U2959 (N_2959,N_2841,N_2846);
and U2960 (N_2960,N_2838,N_2855);
nor U2961 (N_2961,N_2877,N_2833);
and U2962 (N_2962,N_2892,N_2898);
nor U2963 (N_2963,N_2855,N_2851);
or U2964 (N_2964,N_2876,N_2852);
nor U2965 (N_2965,N_2820,N_2803);
nand U2966 (N_2966,N_2802,N_2899);
nand U2967 (N_2967,N_2839,N_2830);
nand U2968 (N_2968,N_2839,N_2814);
nor U2969 (N_2969,N_2824,N_2814);
and U2970 (N_2970,N_2876,N_2805);
or U2971 (N_2971,N_2820,N_2836);
or U2972 (N_2972,N_2850,N_2886);
xnor U2973 (N_2973,N_2837,N_2818);
nor U2974 (N_2974,N_2808,N_2836);
nand U2975 (N_2975,N_2899,N_2832);
nor U2976 (N_2976,N_2881,N_2890);
and U2977 (N_2977,N_2812,N_2826);
nor U2978 (N_2978,N_2894,N_2850);
nand U2979 (N_2979,N_2803,N_2839);
nor U2980 (N_2980,N_2844,N_2870);
nand U2981 (N_2981,N_2825,N_2831);
nor U2982 (N_2982,N_2873,N_2886);
xor U2983 (N_2983,N_2813,N_2803);
or U2984 (N_2984,N_2870,N_2853);
and U2985 (N_2985,N_2847,N_2855);
nand U2986 (N_2986,N_2883,N_2816);
and U2987 (N_2987,N_2802,N_2820);
nor U2988 (N_2988,N_2894,N_2832);
and U2989 (N_2989,N_2804,N_2839);
or U2990 (N_2990,N_2845,N_2891);
nor U2991 (N_2991,N_2862,N_2895);
and U2992 (N_2992,N_2809,N_2831);
nand U2993 (N_2993,N_2818,N_2835);
and U2994 (N_2994,N_2880,N_2831);
nor U2995 (N_2995,N_2833,N_2815);
nor U2996 (N_2996,N_2830,N_2882);
nor U2997 (N_2997,N_2826,N_2831);
nor U2998 (N_2998,N_2804,N_2873);
and U2999 (N_2999,N_2806,N_2816);
nand UO_0 (O_0,N_2934,N_2948);
or UO_1 (O_1,N_2905,N_2936);
nand UO_2 (O_2,N_2950,N_2938);
nor UO_3 (O_3,N_2977,N_2990);
nor UO_4 (O_4,N_2961,N_2949);
nand UO_5 (O_5,N_2988,N_2903);
and UO_6 (O_6,N_2970,N_2942);
nand UO_7 (O_7,N_2935,N_2901);
or UO_8 (O_8,N_2967,N_2929);
nor UO_9 (O_9,N_2939,N_2925);
nor UO_10 (O_10,N_2907,N_2960);
nor UO_11 (O_11,N_2911,N_2943);
and UO_12 (O_12,N_2941,N_2912);
nor UO_13 (O_13,N_2926,N_2946);
or UO_14 (O_14,N_2974,N_2962);
nand UO_15 (O_15,N_2906,N_2932);
xor UO_16 (O_16,N_2922,N_2947);
or UO_17 (O_17,N_2921,N_2965);
and UO_18 (O_18,N_2957,N_2933);
nor UO_19 (O_19,N_2958,N_2973);
xor UO_20 (O_20,N_2963,N_2964);
nor UO_21 (O_21,N_2952,N_2914);
nand UO_22 (O_22,N_2953,N_2993);
and UO_23 (O_23,N_2919,N_2920);
nor UO_24 (O_24,N_2916,N_2937);
nand UO_25 (O_25,N_2986,N_2992);
nand UO_26 (O_26,N_2910,N_2902);
and UO_27 (O_27,N_2904,N_2931);
nor UO_28 (O_28,N_2984,N_2940);
or UO_29 (O_29,N_2956,N_2918);
nor UO_30 (O_30,N_2930,N_2989);
or UO_31 (O_31,N_2976,N_2966);
and UO_32 (O_32,N_2980,N_2915);
and UO_33 (O_33,N_2987,N_2900);
nor UO_34 (O_34,N_2944,N_2951);
or UO_35 (O_35,N_2923,N_2998);
nor UO_36 (O_36,N_2997,N_2995);
nor UO_37 (O_37,N_2969,N_2972);
xnor UO_38 (O_38,N_2983,N_2985);
nand UO_39 (O_39,N_2955,N_2927);
nor UO_40 (O_40,N_2975,N_2917);
nor UO_41 (O_41,N_2996,N_2978);
nor UO_42 (O_42,N_2982,N_2994);
nor UO_43 (O_43,N_2924,N_2971);
and UO_44 (O_44,N_2909,N_2991);
or UO_45 (O_45,N_2908,N_2979);
or UO_46 (O_46,N_2981,N_2954);
nand UO_47 (O_47,N_2928,N_2913);
or UO_48 (O_48,N_2959,N_2945);
nand UO_49 (O_49,N_2968,N_2999);
nor UO_50 (O_50,N_2963,N_2982);
nand UO_51 (O_51,N_2956,N_2932);
nor UO_52 (O_52,N_2993,N_2958);
nand UO_53 (O_53,N_2926,N_2924);
or UO_54 (O_54,N_2903,N_2934);
nor UO_55 (O_55,N_2940,N_2904);
nor UO_56 (O_56,N_2972,N_2983);
or UO_57 (O_57,N_2970,N_2951);
xnor UO_58 (O_58,N_2923,N_2976);
or UO_59 (O_59,N_2993,N_2918);
and UO_60 (O_60,N_2912,N_2980);
and UO_61 (O_61,N_2988,N_2916);
or UO_62 (O_62,N_2926,N_2909);
nor UO_63 (O_63,N_2931,N_2922);
and UO_64 (O_64,N_2976,N_2924);
nand UO_65 (O_65,N_2997,N_2910);
nand UO_66 (O_66,N_2977,N_2969);
or UO_67 (O_67,N_2919,N_2971);
and UO_68 (O_68,N_2982,N_2996);
nand UO_69 (O_69,N_2995,N_2913);
nand UO_70 (O_70,N_2941,N_2948);
xnor UO_71 (O_71,N_2934,N_2920);
nand UO_72 (O_72,N_2957,N_2960);
or UO_73 (O_73,N_2933,N_2993);
nor UO_74 (O_74,N_2961,N_2935);
nor UO_75 (O_75,N_2975,N_2939);
nand UO_76 (O_76,N_2995,N_2908);
nor UO_77 (O_77,N_2994,N_2905);
nor UO_78 (O_78,N_2908,N_2943);
and UO_79 (O_79,N_2984,N_2944);
nor UO_80 (O_80,N_2915,N_2974);
nor UO_81 (O_81,N_2932,N_2970);
and UO_82 (O_82,N_2983,N_2969);
and UO_83 (O_83,N_2918,N_2941);
and UO_84 (O_84,N_2994,N_2948);
nand UO_85 (O_85,N_2930,N_2900);
or UO_86 (O_86,N_2946,N_2981);
nor UO_87 (O_87,N_2958,N_2900);
nand UO_88 (O_88,N_2948,N_2912);
or UO_89 (O_89,N_2938,N_2934);
and UO_90 (O_90,N_2995,N_2994);
and UO_91 (O_91,N_2937,N_2950);
xnor UO_92 (O_92,N_2910,N_2941);
or UO_93 (O_93,N_2932,N_2903);
xor UO_94 (O_94,N_2901,N_2977);
nand UO_95 (O_95,N_2986,N_2994);
nand UO_96 (O_96,N_2905,N_2900);
or UO_97 (O_97,N_2959,N_2968);
and UO_98 (O_98,N_2961,N_2998);
nand UO_99 (O_99,N_2953,N_2981);
nor UO_100 (O_100,N_2978,N_2919);
nand UO_101 (O_101,N_2926,N_2996);
nand UO_102 (O_102,N_2931,N_2999);
nor UO_103 (O_103,N_2959,N_2930);
nor UO_104 (O_104,N_2965,N_2975);
nand UO_105 (O_105,N_2927,N_2989);
nor UO_106 (O_106,N_2939,N_2977);
nand UO_107 (O_107,N_2909,N_2939);
and UO_108 (O_108,N_2946,N_2957);
nand UO_109 (O_109,N_2903,N_2941);
and UO_110 (O_110,N_2995,N_2990);
or UO_111 (O_111,N_2926,N_2929);
or UO_112 (O_112,N_2943,N_2988);
and UO_113 (O_113,N_2968,N_2907);
and UO_114 (O_114,N_2993,N_2974);
nor UO_115 (O_115,N_2977,N_2929);
xnor UO_116 (O_116,N_2929,N_2920);
or UO_117 (O_117,N_2930,N_2990);
or UO_118 (O_118,N_2989,N_2904);
and UO_119 (O_119,N_2962,N_2949);
nor UO_120 (O_120,N_2971,N_2955);
and UO_121 (O_121,N_2987,N_2929);
and UO_122 (O_122,N_2901,N_2998);
and UO_123 (O_123,N_2954,N_2933);
and UO_124 (O_124,N_2902,N_2975);
nor UO_125 (O_125,N_2964,N_2946);
or UO_126 (O_126,N_2938,N_2932);
nor UO_127 (O_127,N_2964,N_2918);
nand UO_128 (O_128,N_2905,N_2967);
nand UO_129 (O_129,N_2978,N_2916);
or UO_130 (O_130,N_2926,N_2943);
and UO_131 (O_131,N_2958,N_2941);
nor UO_132 (O_132,N_2909,N_2998);
xor UO_133 (O_133,N_2934,N_2926);
or UO_134 (O_134,N_2976,N_2931);
and UO_135 (O_135,N_2903,N_2929);
nand UO_136 (O_136,N_2930,N_2998);
nor UO_137 (O_137,N_2963,N_2978);
nand UO_138 (O_138,N_2934,N_2918);
or UO_139 (O_139,N_2967,N_2934);
nand UO_140 (O_140,N_2908,N_2927);
xnor UO_141 (O_141,N_2990,N_2974);
and UO_142 (O_142,N_2917,N_2997);
or UO_143 (O_143,N_2991,N_2941);
or UO_144 (O_144,N_2929,N_2950);
nor UO_145 (O_145,N_2982,N_2972);
xor UO_146 (O_146,N_2904,N_2922);
nand UO_147 (O_147,N_2983,N_2961);
xor UO_148 (O_148,N_2938,N_2952);
or UO_149 (O_149,N_2968,N_2935);
and UO_150 (O_150,N_2968,N_2994);
or UO_151 (O_151,N_2948,N_2983);
nand UO_152 (O_152,N_2987,N_2931);
nand UO_153 (O_153,N_2934,N_2906);
nand UO_154 (O_154,N_2986,N_2998);
or UO_155 (O_155,N_2993,N_2952);
nor UO_156 (O_156,N_2934,N_2921);
and UO_157 (O_157,N_2999,N_2967);
or UO_158 (O_158,N_2909,N_2947);
nand UO_159 (O_159,N_2990,N_2944);
or UO_160 (O_160,N_2904,N_2953);
and UO_161 (O_161,N_2904,N_2977);
and UO_162 (O_162,N_2964,N_2903);
or UO_163 (O_163,N_2923,N_2914);
and UO_164 (O_164,N_2923,N_2910);
nor UO_165 (O_165,N_2936,N_2963);
xnor UO_166 (O_166,N_2927,N_2994);
nor UO_167 (O_167,N_2932,N_2936);
xor UO_168 (O_168,N_2987,N_2908);
or UO_169 (O_169,N_2945,N_2925);
or UO_170 (O_170,N_2968,N_2938);
nand UO_171 (O_171,N_2935,N_2929);
nand UO_172 (O_172,N_2950,N_2997);
and UO_173 (O_173,N_2935,N_2942);
xor UO_174 (O_174,N_2990,N_2905);
or UO_175 (O_175,N_2903,N_2973);
and UO_176 (O_176,N_2998,N_2957);
nand UO_177 (O_177,N_2968,N_2915);
or UO_178 (O_178,N_2950,N_2933);
and UO_179 (O_179,N_2934,N_2990);
nor UO_180 (O_180,N_2952,N_2964);
nor UO_181 (O_181,N_2907,N_2902);
nand UO_182 (O_182,N_2914,N_2947);
nand UO_183 (O_183,N_2941,N_2929);
and UO_184 (O_184,N_2963,N_2903);
nor UO_185 (O_185,N_2942,N_2968);
nor UO_186 (O_186,N_2910,N_2982);
nor UO_187 (O_187,N_2998,N_2985);
or UO_188 (O_188,N_2919,N_2951);
or UO_189 (O_189,N_2929,N_2932);
nor UO_190 (O_190,N_2906,N_2974);
or UO_191 (O_191,N_2965,N_2901);
nand UO_192 (O_192,N_2990,N_2949);
and UO_193 (O_193,N_2942,N_2937);
xnor UO_194 (O_194,N_2984,N_2982);
and UO_195 (O_195,N_2906,N_2918);
or UO_196 (O_196,N_2913,N_2911);
nor UO_197 (O_197,N_2994,N_2904);
nand UO_198 (O_198,N_2954,N_2988);
nor UO_199 (O_199,N_2961,N_2952);
nor UO_200 (O_200,N_2910,N_2948);
nor UO_201 (O_201,N_2908,N_2981);
and UO_202 (O_202,N_2945,N_2926);
nor UO_203 (O_203,N_2979,N_2932);
or UO_204 (O_204,N_2975,N_2954);
or UO_205 (O_205,N_2971,N_2907);
nor UO_206 (O_206,N_2911,N_2945);
or UO_207 (O_207,N_2954,N_2999);
nor UO_208 (O_208,N_2974,N_2943);
or UO_209 (O_209,N_2939,N_2949);
nand UO_210 (O_210,N_2954,N_2979);
and UO_211 (O_211,N_2956,N_2919);
nand UO_212 (O_212,N_2976,N_2961);
and UO_213 (O_213,N_2950,N_2954);
or UO_214 (O_214,N_2904,N_2998);
or UO_215 (O_215,N_2938,N_2969);
and UO_216 (O_216,N_2959,N_2934);
xor UO_217 (O_217,N_2970,N_2957);
and UO_218 (O_218,N_2968,N_2922);
nor UO_219 (O_219,N_2933,N_2931);
and UO_220 (O_220,N_2939,N_2929);
nor UO_221 (O_221,N_2983,N_2939);
or UO_222 (O_222,N_2961,N_2970);
nand UO_223 (O_223,N_2941,N_2998);
nor UO_224 (O_224,N_2905,N_2955);
nor UO_225 (O_225,N_2937,N_2994);
nand UO_226 (O_226,N_2954,N_2992);
or UO_227 (O_227,N_2962,N_2948);
nor UO_228 (O_228,N_2925,N_2907);
or UO_229 (O_229,N_2990,N_2954);
and UO_230 (O_230,N_2969,N_2961);
nand UO_231 (O_231,N_2997,N_2938);
and UO_232 (O_232,N_2943,N_2977);
and UO_233 (O_233,N_2942,N_2905);
nand UO_234 (O_234,N_2919,N_2915);
nor UO_235 (O_235,N_2961,N_2957);
nor UO_236 (O_236,N_2973,N_2938);
nand UO_237 (O_237,N_2987,N_2927);
nand UO_238 (O_238,N_2907,N_2959);
nand UO_239 (O_239,N_2943,N_2928);
nand UO_240 (O_240,N_2933,N_2995);
or UO_241 (O_241,N_2919,N_2946);
or UO_242 (O_242,N_2932,N_2991);
nand UO_243 (O_243,N_2994,N_2984);
nor UO_244 (O_244,N_2939,N_2933);
xor UO_245 (O_245,N_2936,N_2907);
nor UO_246 (O_246,N_2983,N_2953);
or UO_247 (O_247,N_2942,N_2992);
nor UO_248 (O_248,N_2956,N_2922);
nor UO_249 (O_249,N_2946,N_2969);
or UO_250 (O_250,N_2919,N_2959);
nand UO_251 (O_251,N_2929,N_2964);
xnor UO_252 (O_252,N_2926,N_2965);
nor UO_253 (O_253,N_2986,N_2901);
xor UO_254 (O_254,N_2914,N_2924);
nor UO_255 (O_255,N_2993,N_2937);
or UO_256 (O_256,N_2969,N_2955);
and UO_257 (O_257,N_2956,N_2945);
nand UO_258 (O_258,N_2916,N_2902);
nor UO_259 (O_259,N_2981,N_2915);
nor UO_260 (O_260,N_2925,N_2968);
or UO_261 (O_261,N_2977,N_2935);
nand UO_262 (O_262,N_2900,N_2942);
nand UO_263 (O_263,N_2971,N_2991);
nand UO_264 (O_264,N_2933,N_2978);
and UO_265 (O_265,N_2928,N_2967);
xor UO_266 (O_266,N_2940,N_2990);
nor UO_267 (O_267,N_2998,N_2964);
or UO_268 (O_268,N_2996,N_2925);
nor UO_269 (O_269,N_2905,N_2923);
xnor UO_270 (O_270,N_2950,N_2904);
nor UO_271 (O_271,N_2912,N_2916);
nor UO_272 (O_272,N_2975,N_2919);
and UO_273 (O_273,N_2921,N_2913);
and UO_274 (O_274,N_2923,N_2992);
and UO_275 (O_275,N_2940,N_2972);
or UO_276 (O_276,N_2986,N_2937);
nand UO_277 (O_277,N_2902,N_2955);
nand UO_278 (O_278,N_2926,N_2987);
or UO_279 (O_279,N_2939,N_2971);
xor UO_280 (O_280,N_2940,N_2927);
or UO_281 (O_281,N_2912,N_2943);
or UO_282 (O_282,N_2983,N_2912);
nand UO_283 (O_283,N_2914,N_2959);
nor UO_284 (O_284,N_2920,N_2989);
nor UO_285 (O_285,N_2983,N_2966);
and UO_286 (O_286,N_2929,N_2993);
nand UO_287 (O_287,N_2916,N_2996);
and UO_288 (O_288,N_2994,N_2953);
or UO_289 (O_289,N_2995,N_2931);
or UO_290 (O_290,N_2982,N_2993);
xnor UO_291 (O_291,N_2958,N_2989);
nor UO_292 (O_292,N_2918,N_2974);
or UO_293 (O_293,N_2944,N_2928);
nor UO_294 (O_294,N_2947,N_2984);
and UO_295 (O_295,N_2960,N_2985);
or UO_296 (O_296,N_2939,N_2967);
nor UO_297 (O_297,N_2971,N_2990);
or UO_298 (O_298,N_2923,N_2966);
or UO_299 (O_299,N_2998,N_2967);
nand UO_300 (O_300,N_2963,N_2904);
xnor UO_301 (O_301,N_2977,N_2928);
or UO_302 (O_302,N_2953,N_2901);
or UO_303 (O_303,N_2901,N_2980);
and UO_304 (O_304,N_2907,N_2955);
nand UO_305 (O_305,N_2959,N_2901);
and UO_306 (O_306,N_2924,N_2939);
or UO_307 (O_307,N_2955,N_2943);
nand UO_308 (O_308,N_2901,N_2976);
and UO_309 (O_309,N_2978,N_2942);
and UO_310 (O_310,N_2903,N_2995);
nand UO_311 (O_311,N_2983,N_2903);
nand UO_312 (O_312,N_2946,N_2928);
nand UO_313 (O_313,N_2951,N_2910);
nand UO_314 (O_314,N_2927,N_2952);
nand UO_315 (O_315,N_2901,N_2934);
or UO_316 (O_316,N_2916,N_2943);
xor UO_317 (O_317,N_2915,N_2905);
or UO_318 (O_318,N_2978,N_2954);
and UO_319 (O_319,N_2994,N_2916);
or UO_320 (O_320,N_2945,N_2957);
nor UO_321 (O_321,N_2919,N_2964);
or UO_322 (O_322,N_2928,N_2966);
and UO_323 (O_323,N_2986,N_2964);
nand UO_324 (O_324,N_2994,N_2966);
nand UO_325 (O_325,N_2933,N_2952);
xnor UO_326 (O_326,N_2948,N_2938);
or UO_327 (O_327,N_2972,N_2930);
and UO_328 (O_328,N_2943,N_2957);
nor UO_329 (O_329,N_2983,N_2915);
or UO_330 (O_330,N_2927,N_2965);
and UO_331 (O_331,N_2911,N_2908);
xnor UO_332 (O_332,N_2903,N_2901);
or UO_333 (O_333,N_2900,N_2907);
nor UO_334 (O_334,N_2919,N_2988);
nor UO_335 (O_335,N_2989,N_2910);
nand UO_336 (O_336,N_2910,N_2953);
and UO_337 (O_337,N_2964,N_2920);
or UO_338 (O_338,N_2949,N_2951);
and UO_339 (O_339,N_2932,N_2993);
xor UO_340 (O_340,N_2995,N_2999);
nand UO_341 (O_341,N_2915,N_2920);
nand UO_342 (O_342,N_2996,N_2975);
and UO_343 (O_343,N_2931,N_2972);
nand UO_344 (O_344,N_2913,N_2939);
nand UO_345 (O_345,N_2904,N_2900);
nor UO_346 (O_346,N_2907,N_2940);
nand UO_347 (O_347,N_2995,N_2977);
nand UO_348 (O_348,N_2918,N_2994);
and UO_349 (O_349,N_2987,N_2992);
or UO_350 (O_350,N_2922,N_2944);
nor UO_351 (O_351,N_2995,N_2938);
or UO_352 (O_352,N_2968,N_2904);
nor UO_353 (O_353,N_2936,N_2990);
nor UO_354 (O_354,N_2958,N_2940);
xnor UO_355 (O_355,N_2995,N_2979);
nor UO_356 (O_356,N_2955,N_2928);
xor UO_357 (O_357,N_2978,N_2900);
nor UO_358 (O_358,N_2941,N_2913);
or UO_359 (O_359,N_2980,N_2928);
nor UO_360 (O_360,N_2978,N_2961);
and UO_361 (O_361,N_2902,N_2923);
nand UO_362 (O_362,N_2995,N_2936);
nand UO_363 (O_363,N_2973,N_2996);
and UO_364 (O_364,N_2936,N_2928);
and UO_365 (O_365,N_2993,N_2927);
nor UO_366 (O_366,N_2953,N_2928);
nand UO_367 (O_367,N_2907,N_2903);
or UO_368 (O_368,N_2917,N_2977);
nand UO_369 (O_369,N_2969,N_2912);
or UO_370 (O_370,N_2939,N_2955);
or UO_371 (O_371,N_2999,N_2918);
nand UO_372 (O_372,N_2918,N_2926);
or UO_373 (O_373,N_2937,N_2923);
nor UO_374 (O_374,N_2994,N_2933);
nor UO_375 (O_375,N_2926,N_2938);
and UO_376 (O_376,N_2948,N_2915);
xor UO_377 (O_377,N_2985,N_2976);
nand UO_378 (O_378,N_2922,N_2938);
or UO_379 (O_379,N_2967,N_2922);
nand UO_380 (O_380,N_2983,N_2908);
nand UO_381 (O_381,N_2923,N_2918);
or UO_382 (O_382,N_2975,N_2972);
and UO_383 (O_383,N_2933,N_2992);
or UO_384 (O_384,N_2953,N_2908);
nand UO_385 (O_385,N_2942,N_2985);
nor UO_386 (O_386,N_2907,N_2941);
or UO_387 (O_387,N_2907,N_2932);
or UO_388 (O_388,N_2981,N_2921);
or UO_389 (O_389,N_2901,N_2927);
nor UO_390 (O_390,N_2985,N_2969);
and UO_391 (O_391,N_2903,N_2999);
nor UO_392 (O_392,N_2910,N_2958);
and UO_393 (O_393,N_2931,N_2917);
nand UO_394 (O_394,N_2927,N_2954);
or UO_395 (O_395,N_2938,N_2942);
or UO_396 (O_396,N_2923,N_2951);
nor UO_397 (O_397,N_2954,N_2951);
xnor UO_398 (O_398,N_2938,N_2990);
nand UO_399 (O_399,N_2929,N_2907);
and UO_400 (O_400,N_2917,N_2949);
nor UO_401 (O_401,N_2932,N_2982);
nor UO_402 (O_402,N_2900,N_2997);
nand UO_403 (O_403,N_2973,N_2901);
xor UO_404 (O_404,N_2923,N_2946);
nor UO_405 (O_405,N_2977,N_2915);
and UO_406 (O_406,N_2957,N_2944);
and UO_407 (O_407,N_2925,N_2931);
or UO_408 (O_408,N_2917,N_2930);
or UO_409 (O_409,N_2948,N_2961);
and UO_410 (O_410,N_2967,N_2937);
and UO_411 (O_411,N_2965,N_2950);
nor UO_412 (O_412,N_2928,N_2945);
nor UO_413 (O_413,N_2927,N_2998);
nor UO_414 (O_414,N_2976,N_2959);
and UO_415 (O_415,N_2918,N_2936);
or UO_416 (O_416,N_2974,N_2964);
nand UO_417 (O_417,N_2932,N_2950);
and UO_418 (O_418,N_2997,N_2944);
or UO_419 (O_419,N_2931,N_2990);
xor UO_420 (O_420,N_2973,N_2902);
nand UO_421 (O_421,N_2956,N_2985);
nor UO_422 (O_422,N_2914,N_2935);
xnor UO_423 (O_423,N_2966,N_2992);
nand UO_424 (O_424,N_2981,N_2914);
and UO_425 (O_425,N_2917,N_2971);
and UO_426 (O_426,N_2959,N_2944);
or UO_427 (O_427,N_2926,N_2956);
nor UO_428 (O_428,N_2909,N_2944);
nor UO_429 (O_429,N_2963,N_2913);
or UO_430 (O_430,N_2971,N_2946);
or UO_431 (O_431,N_2954,N_2974);
nor UO_432 (O_432,N_2924,N_2951);
and UO_433 (O_433,N_2955,N_2960);
or UO_434 (O_434,N_2984,N_2985);
or UO_435 (O_435,N_2917,N_2961);
nand UO_436 (O_436,N_2980,N_2951);
nor UO_437 (O_437,N_2973,N_2912);
and UO_438 (O_438,N_2915,N_2914);
nand UO_439 (O_439,N_2935,N_2952);
and UO_440 (O_440,N_2935,N_2920);
nand UO_441 (O_441,N_2932,N_2958);
nor UO_442 (O_442,N_2918,N_2916);
nor UO_443 (O_443,N_2996,N_2909);
and UO_444 (O_444,N_2901,N_2966);
xnor UO_445 (O_445,N_2926,N_2964);
nor UO_446 (O_446,N_2985,N_2946);
or UO_447 (O_447,N_2993,N_2924);
or UO_448 (O_448,N_2988,N_2995);
nand UO_449 (O_449,N_2979,N_2944);
and UO_450 (O_450,N_2911,N_2912);
nand UO_451 (O_451,N_2940,N_2969);
and UO_452 (O_452,N_2990,N_2914);
or UO_453 (O_453,N_2987,N_2997);
nor UO_454 (O_454,N_2961,N_2909);
or UO_455 (O_455,N_2949,N_2958);
or UO_456 (O_456,N_2904,N_2919);
or UO_457 (O_457,N_2944,N_2975);
nand UO_458 (O_458,N_2986,N_2947);
and UO_459 (O_459,N_2974,N_2979);
nor UO_460 (O_460,N_2913,N_2972);
or UO_461 (O_461,N_2987,N_2916);
nor UO_462 (O_462,N_2976,N_2960);
or UO_463 (O_463,N_2926,N_2970);
nor UO_464 (O_464,N_2957,N_2967);
nand UO_465 (O_465,N_2920,N_2965);
or UO_466 (O_466,N_2970,N_2997);
and UO_467 (O_467,N_2938,N_2987);
nor UO_468 (O_468,N_2925,N_2960);
and UO_469 (O_469,N_2946,N_2940);
and UO_470 (O_470,N_2916,N_2958);
and UO_471 (O_471,N_2975,N_2977);
and UO_472 (O_472,N_2954,N_2928);
or UO_473 (O_473,N_2947,N_2977);
or UO_474 (O_474,N_2974,N_2930);
nand UO_475 (O_475,N_2946,N_2955);
nand UO_476 (O_476,N_2923,N_2900);
or UO_477 (O_477,N_2967,N_2952);
or UO_478 (O_478,N_2998,N_2988);
and UO_479 (O_479,N_2998,N_2979);
nand UO_480 (O_480,N_2986,N_2975);
or UO_481 (O_481,N_2987,N_2915);
and UO_482 (O_482,N_2928,N_2900);
and UO_483 (O_483,N_2979,N_2992);
nor UO_484 (O_484,N_2936,N_2914);
or UO_485 (O_485,N_2995,N_2925);
nor UO_486 (O_486,N_2974,N_2966);
nor UO_487 (O_487,N_2972,N_2978);
and UO_488 (O_488,N_2941,N_2905);
xnor UO_489 (O_489,N_2965,N_2959);
or UO_490 (O_490,N_2943,N_2981);
and UO_491 (O_491,N_2909,N_2974);
and UO_492 (O_492,N_2936,N_2981);
or UO_493 (O_493,N_2901,N_2944);
nand UO_494 (O_494,N_2941,N_2920);
or UO_495 (O_495,N_2917,N_2932);
or UO_496 (O_496,N_2913,N_2931);
or UO_497 (O_497,N_2936,N_2917);
or UO_498 (O_498,N_2997,N_2935);
and UO_499 (O_499,N_2954,N_2914);
endmodule