module basic_3000_30000_3500_6_levels_10xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
or U0 (N_0,In_1315,In_1951);
or U1 (N_1,In_2124,In_1869);
and U2 (N_2,In_2424,In_1108);
nand U3 (N_3,In_2133,In_34);
nor U4 (N_4,In_867,In_1449);
or U5 (N_5,In_726,In_2453);
nand U6 (N_6,In_2159,In_404);
and U7 (N_7,In_1807,In_599);
nor U8 (N_8,In_2041,In_1554);
nor U9 (N_9,In_2832,In_2307);
xor U10 (N_10,In_865,In_1387);
or U11 (N_11,In_1700,In_2071);
nor U12 (N_12,In_703,In_2875);
xor U13 (N_13,In_1144,In_1656);
nand U14 (N_14,In_1321,In_229);
xor U15 (N_15,In_1585,In_1228);
or U16 (N_16,In_879,In_2940);
or U17 (N_17,In_1252,In_138);
xnor U18 (N_18,In_2695,In_1767);
nor U19 (N_19,In_365,In_2949);
nand U20 (N_20,In_1533,In_2951);
and U21 (N_21,In_1134,In_979);
or U22 (N_22,In_1051,In_479);
nor U23 (N_23,In_1495,In_935);
or U24 (N_24,In_2791,In_2002);
or U25 (N_25,In_840,In_2272);
xnor U26 (N_26,In_716,In_1422);
nand U27 (N_27,In_1112,In_1780);
nor U28 (N_28,In_561,In_1589);
nor U29 (N_29,In_2254,In_2256);
nor U30 (N_30,In_427,In_2952);
nor U31 (N_31,In_2584,In_2934);
xnor U32 (N_32,In_1674,In_1600);
or U33 (N_33,In_806,In_2652);
xor U34 (N_34,In_1011,In_745);
xor U35 (N_35,In_1372,In_1615);
nor U36 (N_36,In_725,In_2800);
nor U37 (N_37,In_2570,In_2937);
xnor U38 (N_38,In_507,In_1128);
and U39 (N_39,In_1703,In_2001);
nand U40 (N_40,In_1403,In_2233);
and U41 (N_41,In_2946,In_2004);
or U42 (N_42,In_2162,In_272);
nand U43 (N_43,In_1029,In_2242);
nand U44 (N_44,In_2099,In_2623);
and U45 (N_45,In_1695,In_554);
nor U46 (N_46,In_2724,In_338);
nand U47 (N_47,In_2353,In_2586);
nor U48 (N_48,In_931,In_2948);
or U49 (N_49,In_199,In_89);
or U50 (N_50,In_2838,In_2651);
nor U51 (N_51,In_735,In_2578);
nor U52 (N_52,In_1133,In_523);
nand U53 (N_53,In_406,In_1844);
nor U54 (N_54,In_1084,In_283);
or U55 (N_55,In_2332,In_2715);
xor U56 (N_56,In_2964,In_1804);
nor U57 (N_57,In_496,In_36);
or U58 (N_58,In_2348,In_1588);
and U59 (N_59,In_2249,In_2330);
or U60 (N_60,In_1294,In_25);
nand U61 (N_61,In_2521,In_2788);
and U62 (N_62,In_2011,In_2169);
xnor U63 (N_63,In_746,In_2881);
or U64 (N_64,In_2527,In_817);
nor U65 (N_65,In_1361,In_1826);
nand U66 (N_66,In_1789,In_331);
xnor U67 (N_67,In_339,In_620);
xor U68 (N_68,In_2892,In_2554);
xor U69 (N_69,In_2545,In_2112);
xor U70 (N_70,In_922,In_1408);
xor U71 (N_71,In_2693,In_531);
and U72 (N_72,In_891,In_1611);
nor U73 (N_73,In_580,In_1979);
xnor U74 (N_74,In_1904,In_1945);
or U75 (N_75,In_2761,In_2670);
nor U76 (N_76,In_141,In_170);
or U77 (N_77,In_150,In_1500);
xnor U78 (N_78,In_1671,In_2437);
xor U79 (N_79,In_307,In_1790);
or U80 (N_80,In_1241,In_103);
nand U81 (N_81,In_1707,In_133);
xor U82 (N_82,In_933,In_1073);
and U83 (N_83,In_2624,In_69);
nand U84 (N_84,In_2529,In_1149);
and U85 (N_85,In_2536,In_1302);
or U86 (N_86,In_648,In_828);
and U87 (N_87,In_1210,In_1960);
or U88 (N_88,In_1092,In_1222);
nor U89 (N_89,In_1863,In_1924);
or U90 (N_90,In_752,In_796);
nor U91 (N_91,In_1362,In_1182);
nand U92 (N_92,In_2565,In_2503);
nor U93 (N_93,In_2901,In_1511);
nand U94 (N_94,In_2762,In_913);
nand U95 (N_95,In_1028,In_2969);
xnor U96 (N_96,In_348,In_642);
or U97 (N_97,In_2911,In_2583);
or U98 (N_98,In_2198,In_1308);
nand U99 (N_99,In_1666,In_2597);
or U100 (N_100,In_1351,In_2375);
xor U101 (N_101,In_2380,In_2073);
or U102 (N_102,In_1292,In_619);
or U103 (N_103,In_1360,In_2590);
and U104 (N_104,In_1591,In_1451);
or U105 (N_105,In_2379,In_1584);
nor U106 (N_106,In_2417,In_704);
or U107 (N_107,In_246,In_2833);
xor U108 (N_108,In_929,In_139);
nand U109 (N_109,In_2500,In_2081);
nor U110 (N_110,In_904,In_1270);
nor U111 (N_111,In_183,In_2701);
nor U112 (N_112,In_37,In_2768);
nor U113 (N_113,In_1848,In_2033);
xor U114 (N_114,In_649,In_189);
or U115 (N_115,In_1738,In_854);
nor U116 (N_116,In_1535,In_2939);
and U117 (N_117,In_739,In_1755);
xnor U118 (N_118,In_938,In_563);
nor U119 (N_119,In_2100,In_15);
xor U120 (N_120,In_2372,In_1670);
or U121 (N_121,In_2920,In_368);
xor U122 (N_122,In_2735,In_117);
nand U123 (N_123,In_187,In_2271);
or U124 (N_124,In_2136,In_968);
nor U125 (N_125,In_361,In_795);
xor U126 (N_126,In_2406,In_537);
nor U127 (N_127,In_1400,In_2672);
nand U128 (N_128,In_737,In_255);
and U129 (N_129,In_1499,In_1934);
or U130 (N_130,In_831,In_1528);
and U131 (N_131,In_2741,In_1344);
or U132 (N_132,In_2535,In_993);
nor U133 (N_133,In_1933,In_306);
or U134 (N_134,In_1353,In_991);
nand U135 (N_135,In_878,In_1727);
and U136 (N_136,In_44,In_462);
and U137 (N_137,In_329,In_2727);
nor U138 (N_138,In_1405,In_1768);
nand U139 (N_139,In_1218,In_851);
and U140 (N_140,In_2110,In_2804);
and U141 (N_141,In_1527,In_345);
xor U142 (N_142,In_2258,In_829);
nor U143 (N_143,In_946,In_151);
nor U144 (N_144,In_321,In_1635);
and U145 (N_145,In_1053,In_812);
nand U146 (N_146,In_1660,In_2058);
nand U147 (N_147,In_2607,In_2582);
nor U148 (N_148,In_2903,In_274);
xor U149 (N_149,In_2154,In_2251);
nand U150 (N_150,In_822,In_2671);
xnor U151 (N_151,In_2673,In_1483);
or U152 (N_152,In_808,In_502);
xor U153 (N_153,In_2856,In_1783);
xor U154 (N_154,In_1506,In_457);
nand U155 (N_155,In_1090,In_1607);
xnor U156 (N_156,In_299,In_1438);
and U157 (N_157,In_2636,In_2177);
nand U158 (N_158,In_676,In_2322);
xnor U159 (N_159,In_1349,In_2354);
nor U160 (N_160,In_2132,In_1243);
nor U161 (N_161,In_1096,In_1632);
xnor U162 (N_162,In_39,In_130);
xnor U163 (N_163,In_2926,In_143);
and U164 (N_164,In_1881,In_1900);
nor U165 (N_165,In_2622,In_2560);
nor U166 (N_166,In_1159,In_257);
or U167 (N_167,In_750,In_2070);
xor U168 (N_168,In_1048,In_1452);
nand U169 (N_169,In_392,In_1192);
nor U170 (N_170,In_1818,In_2489);
and U171 (N_171,In_2596,In_2274);
nor U172 (N_172,In_790,In_1289);
or U173 (N_173,In_2135,In_2577);
nor U174 (N_174,In_572,In_72);
and U175 (N_175,In_1828,In_2748);
xor U176 (N_176,In_1056,In_131);
or U177 (N_177,In_2302,In_679);
and U178 (N_178,In_358,In_625);
nor U179 (N_179,In_2462,In_22);
or U180 (N_180,In_733,In_1079);
or U181 (N_181,In_695,In_2614);
xnor U182 (N_182,In_2241,In_2792);
nor U183 (N_183,In_2435,In_270);
nand U184 (N_184,In_1411,In_90);
or U185 (N_185,In_1023,In_2495);
nand U186 (N_186,In_2669,In_2632);
nand U187 (N_187,In_1166,In_2490);
or U188 (N_188,In_1212,In_2359);
nand U189 (N_189,In_2405,In_107);
or U190 (N_190,In_2660,In_2763);
and U191 (N_191,In_1074,In_1570);
and U192 (N_192,In_1184,In_2456);
and U193 (N_193,In_1172,In_2820);
nor U194 (N_194,In_74,In_1278);
nor U195 (N_195,In_495,In_2181);
and U196 (N_196,In_460,In_1718);
nor U197 (N_197,In_363,In_954);
nand U198 (N_198,In_2769,In_426);
xor U199 (N_199,In_2817,In_1474);
and U200 (N_200,In_1312,In_2824);
or U201 (N_201,In_237,In_2396);
nor U202 (N_202,In_2218,In_1713);
xor U203 (N_203,In_1138,In_2979);
xor U204 (N_204,In_2822,In_273);
xnor U205 (N_205,In_45,In_227);
nor U206 (N_206,In_254,In_2690);
or U207 (N_207,In_10,In_798);
nand U208 (N_208,In_503,In_1675);
nand U209 (N_209,In_962,In_2191);
nor U210 (N_210,In_2047,In_815);
nand U211 (N_211,In_1823,In_1970);
or U212 (N_212,In_2857,In_197);
xor U213 (N_213,In_2953,In_435);
xnor U214 (N_214,In_93,In_1062);
or U215 (N_215,In_2096,In_2784);
xnor U216 (N_216,In_1299,In_1432);
xor U217 (N_217,In_97,In_2329);
nor U218 (N_218,In_1513,In_288);
and U219 (N_219,In_2814,In_2328);
xnor U220 (N_220,In_26,In_1923);
and U221 (N_221,In_1910,In_1442);
nor U222 (N_222,In_1476,In_585);
xor U223 (N_223,In_2340,In_494);
or U224 (N_224,In_1851,In_659);
or U225 (N_225,In_2259,In_223);
nand U226 (N_226,In_2131,In_1874);
or U227 (N_227,In_1634,In_2883);
xor U228 (N_228,In_2163,In_477);
xnor U229 (N_229,In_1428,In_1541);
nor U230 (N_230,In_830,In_1811);
nor U231 (N_231,In_2643,In_264);
xor U232 (N_232,In_190,In_686);
xor U233 (N_233,In_2831,In_767);
and U234 (N_234,In_1803,In_1944);
and U235 (N_235,In_1809,In_1275);
or U236 (N_236,In_2179,In_82);
nor U237 (N_237,In_2567,In_756);
xnor U238 (N_238,In_2368,In_5);
nand U239 (N_239,In_838,In_2611);
and U240 (N_240,In_2757,In_527);
nand U241 (N_241,In_2336,In_2556);
nor U242 (N_242,In_536,In_973);
and U243 (N_243,In_2114,In_284);
and U244 (N_244,In_1510,In_1371);
or U245 (N_245,In_33,In_779);
nand U246 (N_246,In_2884,In_1211);
xor U247 (N_247,In_2166,In_458);
nand U248 (N_248,In_2882,In_66);
nand U249 (N_249,In_2127,In_1751);
xor U250 (N_250,In_970,In_244);
or U251 (N_251,In_1505,In_2014);
nor U252 (N_252,In_2350,In_1490);
or U253 (N_253,In_378,In_755);
nor U254 (N_254,In_2157,In_1447);
or U255 (N_255,In_1203,In_2247);
or U256 (N_256,In_2472,In_129);
xnor U257 (N_257,In_2513,In_1880);
and U258 (N_258,In_628,In_1586);
or U259 (N_259,In_1991,In_2551);
nand U260 (N_260,In_2160,In_2463);
nand U261 (N_261,In_1524,In_1825);
or U262 (N_262,In_2877,In_1471);
nand U263 (N_263,In_720,In_2518);
xor U264 (N_264,In_940,In_2487);
nor U265 (N_265,In_101,In_296);
or U266 (N_266,In_397,In_2726);
nand U267 (N_267,In_1161,In_1123);
nor U268 (N_268,In_2559,In_586);
and U269 (N_269,In_896,In_2180);
or U270 (N_270,In_860,In_1151);
or U271 (N_271,In_401,In_2694);
nand U272 (N_272,In_159,In_1287);
xnor U273 (N_273,In_2494,In_881);
or U274 (N_274,In_1852,In_1042);
and U275 (N_275,In_1415,In_1193);
nand U276 (N_276,In_2716,In_2801);
nor U277 (N_277,In_2092,In_1325);
nand U278 (N_278,In_239,In_1052);
and U279 (N_279,In_781,In_609);
nor U280 (N_280,In_1046,In_2917);
or U281 (N_281,In_2326,In_529);
nor U282 (N_282,In_224,In_76);
and U283 (N_283,In_431,In_952);
nand U284 (N_284,In_1639,In_1988);
or U285 (N_285,In_1550,In_2268);
or U286 (N_286,In_2187,In_196);
nor U287 (N_287,In_783,In_2305);
xnor U288 (N_288,In_2021,In_1534);
xnor U289 (N_289,In_1508,In_2993);
or U290 (N_290,In_682,In_1257);
nand U291 (N_291,In_1005,In_2199);
xnor U292 (N_292,In_2044,In_846);
xor U293 (N_293,In_2200,In_380);
xor U294 (N_294,In_2931,In_32);
or U295 (N_295,In_1076,In_1322);
xor U296 (N_296,In_1304,In_622);
nand U297 (N_297,In_2129,In_1838);
or U298 (N_298,In_489,In_579);
and U299 (N_299,In_2366,In_1791);
or U300 (N_300,In_1016,In_1446);
xor U301 (N_301,In_629,In_1463);
or U302 (N_302,In_1364,In_2645);
nand U303 (N_303,In_80,In_2444);
nor U304 (N_304,In_897,In_2928);
xnor U305 (N_305,In_900,In_2138);
nor U306 (N_306,In_2246,In_589);
nand U307 (N_307,In_1375,In_16);
nor U308 (N_308,In_2561,In_576);
or U309 (N_309,In_2059,In_2525);
nor U310 (N_310,In_1840,In_1756);
xnor U311 (N_311,In_774,In_1641);
or U312 (N_312,In_2467,In_376);
or U313 (N_313,In_2470,In_1676);
or U314 (N_314,In_2052,In_1793);
and U315 (N_315,In_1894,In_1081);
or U316 (N_316,In_2563,In_1575);
and U317 (N_317,In_108,In_2369);
or U318 (N_318,In_930,In_455);
xnor U319 (N_319,In_1231,In_1114);
xor U320 (N_320,In_486,In_438);
xnor U321 (N_321,In_1014,In_2035);
xor U322 (N_322,In_127,In_213);
and U323 (N_323,In_2304,In_1317);
xor U324 (N_324,In_1942,In_882);
nand U325 (N_325,In_594,In_985);
nor U326 (N_326,In_81,In_1063);
xnor U327 (N_327,In_560,In_2466);
nand U328 (N_328,In_1905,In_1984);
nand U329 (N_329,In_461,In_1858);
or U330 (N_330,In_1097,In_2790);
nand U331 (N_331,In_2313,In_2501);
nor U332 (N_332,In_18,In_2203);
and U333 (N_333,In_969,In_419);
nand U334 (N_334,In_2238,In_1009);
nand U335 (N_335,In_1843,In_2922);
nor U336 (N_336,In_1552,In_872);
xnor U337 (N_337,In_472,In_2981);
xor U338 (N_338,In_1737,In_1902);
nand U339 (N_339,In_2223,In_195);
or U340 (N_340,In_506,In_688);
or U341 (N_341,In_2730,In_782);
or U342 (N_342,In_1847,In_2987);
xor U343 (N_343,In_1819,In_293);
or U344 (N_344,In_2502,In_2849);
nor U345 (N_345,In_1850,In_210);
xnor U346 (N_346,In_2867,In_1204);
xnor U347 (N_347,In_2534,In_1341);
or U348 (N_348,In_2595,In_324);
xnor U349 (N_349,In_2683,In_1329);
nand U350 (N_350,In_2451,In_1785);
nand U351 (N_351,In_1024,In_2147);
xor U352 (N_352,In_9,In_422);
nor U353 (N_353,In_1070,In_2030);
nand U354 (N_354,In_2758,In_1339);
nor U355 (N_355,In_1548,In_673);
and U356 (N_356,In_2686,In_2300);
nand U357 (N_357,In_2327,In_1565);
xor U358 (N_358,In_2550,In_1072);
or U359 (N_359,In_1217,In_759);
nor U360 (N_360,In_2255,In_1017);
or U361 (N_361,In_1004,In_1055);
or U362 (N_362,In_2260,In_1202);
or U363 (N_363,In_2775,In_2844);
and U364 (N_364,In_1260,In_276);
nand U365 (N_365,In_1669,In_584);
or U366 (N_366,In_861,In_96);
nor U367 (N_367,In_1687,In_853);
and U368 (N_368,In_2571,In_1020);
nor U369 (N_369,In_1116,In_1340);
nor U370 (N_370,In_1295,In_2539);
or U371 (N_371,In_2383,In_2141);
xnor U372 (N_372,In_723,In_841);
nand U373 (N_373,In_41,In_298);
and U374 (N_374,In_568,In_1741);
or U375 (N_375,In_1201,In_1493);
and U376 (N_376,In_2712,In_2034);
and U377 (N_377,In_2668,In_1736);
nand U378 (N_378,In_2921,In_1121);
nor U379 (N_379,In_1514,In_874);
or U380 (N_380,In_595,In_2699);
nand U381 (N_381,In_520,In_999);
xnor U382 (N_382,In_2342,In_2056);
nor U383 (N_383,In_2943,In_308);
nand U384 (N_384,In_627,In_1194);
xnor U385 (N_385,In_248,In_2760);
nand U386 (N_386,In_1925,In_1244);
nor U387 (N_387,In_1069,In_487);
nand U388 (N_388,In_2175,In_2066);
or U389 (N_389,In_948,In_1698);
nand U390 (N_390,In_656,In_2789);
nand U391 (N_391,In_2457,In_2171);
nand U392 (N_392,In_1410,In_1781);
nor U393 (N_393,In_168,In_2063);
and U394 (N_394,In_2213,In_504);
or U395 (N_395,In_678,In_943);
nor U396 (N_396,In_754,In_2235);
nand U397 (N_397,In_1367,In_364);
nand U398 (N_398,In_1547,In_1000);
nand U399 (N_399,In_2656,In_1553);
xor U400 (N_400,In_1597,In_1147);
nand U401 (N_401,In_730,In_945);
nor U402 (N_402,In_1283,In_2961);
and U403 (N_403,In_309,In_233);
xnor U404 (N_404,In_1383,In_2122);
xnor U405 (N_405,In_888,In_1378);
or U406 (N_406,In_593,In_1143);
nor U407 (N_407,In_2493,In_1573);
and U408 (N_408,In_884,In_245);
and U409 (N_409,In_2054,In_2086);
and U410 (N_410,In_1154,In_1911);
and U411 (N_411,In_1494,In_1022);
nand U412 (N_412,In_1593,In_102);
and U413 (N_413,In_2709,In_1488);
nand U414 (N_414,In_1163,In_371);
and U415 (N_415,In_714,In_1636);
or U416 (N_416,In_105,In_161);
xnor U417 (N_417,In_1532,In_996);
xor U418 (N_418,In_417,In_1327);
nand U419 (N_419,In_2403,In_1814);
nand U420 (N_420,In_344,In_2438);
nor U421 (N_421,In_2729,In_2192);
nand U422 (N_422,In_1131,In_230);
xor U423 (N_423,In_2853,In_243);
nand U424 (N_424,In_2479,In_2025);
nand U425 (N_425,In_1155,In_1730);
xor U426 (N_426,In_1256,In_1877);
nand U427 (N_427,In_1436,In_624);
and U428 (N_428,In_350,In_2777);
and U429 (N_429,In_2331,In_43);
and U430 (N_430,In_2226,In_2074);
xnor U431 (N_431,In_1221,In_2812);
xnor U432 (N_432,In_2846,In_1457);
nand U433 (N_433,In_2930,In_1999);
xnor U434 (N_434,In_1871,In_2638);
and U435 (N_435,In_2772,In_690);
and U436 (N_436,In_2834,In_663);
or U437 (N_437,In_2447,In_2958);
nor U438 (N_438,In_124,In_2776);
and U439 (N_439,In_1758,In_1509);
or U440 (N_440,In_1647,In_2983);
nor U441 (N_441,In_2514,In_1622);
or U442 (N_442,In_645,In_1605);
nor U443 (N_443,In_2286,In_2659);
nor U444 (N_444,In_464,In_2400);
and U445 (N_445,In_2057,In_1664);
nand U446 (N_446,In_1778,In_286);
nand U447 (N_447,In_1916,In_640);
nand U448 (N_448,In_1075,In_2810);
nor U449 (N_449,In_1036,In_149);
or U450 (N_450,In_982,In_2899);
nand U451 (N_451,In_1437,In_1355);
nand U452 (N_452,In_864,In_956);
nor U453 (N_453,In_2579,In_2333);
xor U454 (N_454,In_2870,In_1728);
or U455 (N_455,In_100,In_349);
nor U456 (N_456,In_4,In_497);
nor U457 (N_457,In_1898,In_1420);
nand U458 (N_458,In_801,In_1536);
nand U459 (N_459,In_2989,In_1067);
or U460 (N_460,In_2334,In_615);
nor U461 (N_461,In_153,In_939);
nor U462 (N_462,In_971,In_180);
xor U463 (N_463,In_2619,In_1642);
and U464 (N_464,In_1724,In_2997);
and U465 (N_465,In_616,In_1571);
xnor U466 (N_466,In_509,In_175);
nor U467 (N_467,In_2277,In_116);
or U468 (N_468,In_1873,In_1380);
nand U469 (N_469,In_1199,In_297);
and U470 (N_470,In_2207,In_1441);
or U471 (N_471,In_2868,In_875);
and U472 (N_472,In_858,In_708);
nor U473 (N_473,In_657,In_2984);
nand U474 (N_474,In_498,In_1196);
or U475 (N_475,In_2782,In_1566);
nand U476 (N_476,In_1136,In_2010);
nand U477 (N_477,In_2767,In_277);
nor U478 (N_478,In_1258,In_1467);
or U479 (N_479,In_2480,In_613);
xor U480 (N_480,In_2031,In_1444);
or U481 (N_481,In_2278,In_388);
and U482 (N_482,In_1901,In_611);
nand U483 (N_483,In_2257,In_605);
xnor U484 (N_484,In_972,In_1579);
nor U485 (N_485,In_2013,In_1526);
nor U486 (N_486,In_1595,In_1205);
xnor U487 (N_487,In_148,In_2914);
and U488 (N_488,In_2751,In_1557);
nand U489 (N_489,In_538,In_184);
and U490 (N_490,In_758,In_570);
or U491 (N_491,In_1358,In_2053);
and U492 (N_492,In_386,In_2684);
nor U493 (N_493,In_1649,In_1139);
xnor U494 (N_494,In_451,In_2471);
xor U495 (N_495,In_2971,In_905);
and U496 (N_496,In_1104,In_2364);
or U497 (N_497,In_707,In_2204);
nor U498 (N_498,In_268,In_2287);
and U499 (N_499,In_1188,In_1065);
xnor U500 (N_500,In_1592,In_1033);
or U501 (N_501,In_169,In_2509);
nand U502 (N_502,In_42,In_855);
nor U503 (N_503,In_2675,In_55);
xnor U504 (N_504,In_1862,In_2641);
nor U505 (N_505,In_1684,In_2318);
nand U506 (N_506,In_399,In_1148);
or U507 (N_507,In_771,In_528);
nand U508 (N_508,In_2009,In_313);
nand U509 (N_509,In_849,In_1972);
and U510 (N_510,In_2866,In_1187);
or U511 (N_511,In_2404,In_967);
nor U512 (N_512,In_1849,In_1884);
and U513 (N_513,In_1821,In_453);
and U514 (N_514,In_748,In_1518);
or U515 (N_515,In_2900,In_2786);
and U516 (N_516,In_886,In_1854);
and U517 (N_517,In_792,In_1832);
and U518 (N_518,In_221,In_512);
or U519 (N_519,In_1460,In_1426);
nor U520 (N_520,In_119,In_1389);
xnor U521 (N_521,In_488,In_2077);
nor U522 (N_522,In_2061,In_145);
xor U523 (N_523,In_1215,In_2345);
nand U524 (N_524,In_957,In_1558);
nor U525 (N_525,In_1425,In_2944);
and U526 (N_526,In_2793,In_2523);
xor U527 (N_527,In_1305,In_2826);
and U528 (N_528,In_1887,In_2125);
or U529 (N_529,In_1961,In_58);
and U530 (N_530,In_330,In_1926);
nor U531 (N_531,In_1157,In_661);
and U532 (N_532,In_2923,In_1745);
nand U533 (N_533,In_2072,In_48);
and U534 (N_534,In_850,In_1797);
nor U535 (N_535,In_721,In_816);
or U536 (N_536,In_430,In_396);
nand U537 (N_537,In_2553,In_2173);
and U538 (N_538,In_2108,In_852);
and U539 (N_539,In_393,In_2309);
nor U540 (N_540,In_1087,In_3);
xnor U541 (N_541,In_677,In_62);
xor U542 (N_542,In_1485,In_1227);
nand U543 (N_543,In_2387,In_2893);
nand U544 (N_544,In_30,In_377);
or U545 (N_545,In_1333,In_549);
nor U546 (N_546,In_207,In_786);
or U547 (N_547,In_1773,In_1058);
or U548 (N_548,In_670,In_135);
xnor U549 (N_549,In_919,In_610);
nor U550 (N_550,In_2575,In_302);
and U551 (N_551,In_542,In_1454);
nor U552 (N_552,In_471,In_2802);
nor U553 (N_553,In_2732,In_2687);
or U554 (N_554,In_2774,In_2644);
nand U555 (N_555,In_2977,In_718);
nor U556 (N_556,In_1958,In_87);
nand U557 (N_557,In_1842,In_1010);
and U558 (N_558,In_1846,In_1171);
and U559 (N_559,In_409,In_1279);
nor U560 (N_560,In_2739,In_1829);
xor U561 (N_561,In_2408,In_2880);
or U562 (N_562,In_2592,In_2864);
nor U563 (N_563,In_2418,In_1354);
or U564 (N_564,In_1234,In_734);
or U565 (N_565,In_2894,In_581);
nand U566 (N_566,In_2394,In_1559);
and U567 (N_567,In_2411,In_2121);
xor U568 (N_568,In_1127,In_2787);
xor U569 (N_569,In_1678,In_1419);
or U570 (N_570,In_1750,In_1150);
and U571 (N_571,In_711,In_1975);
nor U572 (N_572,In_1608,In_2308);
nand U573 (N_573,In_1130,In_1384);
and U574 (N_574,In_2642,In_1612);
nand U575 (N_575,In_1692,In_741);
nor U576 (N_576,In_2458,In_499);
or U577 (N_577,In_425,In_94);
and U578 (N_578,In_78,In_155);
nor U579 (N_579,In_1041,In_1968);
or U580 (N_580,In_1930,In_2341);
xnor U581 (N_581,In_1263,In_1037);
xnor U582 (N_582,In_1817,In_2219);
nor U583 (N_583,In_7,In_446);
xnor U584 (N_584,In_2616,In_343);
xnor U585 (N_585,In_1782,In_1752);
or U586 (N_586,In_2012,In_2423);
or U587 (N_587,In_179,In_433);
or U588 (N_588,In_1313,In_2499);
nand U589 (N_589,In_2778,In_2442);
or U590 (N_590,In_1233,In_1481);
and U591 (N_591,In_2850,In_2610);
nand U592 (N_592,In_1857,In_1050);
and U593 (N_593,In_304,In_1099);
and U594 (N_594,In_1907,In_421);
or U595 (N_595,In_2320,In_2401);
nand U596 (N_596,In_327,In_1619);
nand U597 (N_597,In_1953,In_500);
xnor U598 (N_598,In_804,In_2816);
and U599 (N_599,In_2798,In_1583);
nor U600 (N_600,In_1480,In_1717);
xor U601 (N_601,In_226,In_1342);
and U602 (N_602,In_1722,In_398);
xor U603 (N_603,In_2183,In_1316);
nor U604 (N_604,In_2541,In_1516);
nand U605 (N_605,In_191,In_2796);
xor U606 (N_606,In_1347,In_990);
or U607 (N_607,In_2842,In_1543);
or U608 (N_608,In_1685,In_1563);
and U609 (N_609,In_2865,In_1195);
nand U610 (N_610,In_963,In_2427);
nor U611 (N_611,In_1274,In_1679);
nand U612 (N_612,In_2734,In_1820);
and U613 (N_613,In_1981,In_2708);
and U614 (N_614,In_391,In_1653);
xnor U615 (N_615,In_1061,In_552);
or U616 (N_616,In_305,In_2311);
nor U617 (N_617,In_1802,In_1191);
and U618 (N_618,In_2743,In_2087);
nor U619 (N_619,In_1609,In_2091);
xnor U620 (N_620,In_709,In_1078);
or U621 (N_621,In_285,In_2915);
xor U622 (N_622,In_1235,In_578);
and U623 (N_623,In_193,In_2615);
nor U624 (N_624,In_1969,In_2297);
nor U625 (N_625,In_2655,In_1667);
nand U626 (N_626,In_1937,In_442);
and U627 (N_627,In_429,In_1486);
and U628 (N_628,In_2722,In_2587);
xor U629 (N_629,In_869,In_983);
nor U630 (N_630,In_701,In_1875);
nor U631 (N_631,In_2212,In_174);
and U632 (N_632,In_2508,In_1531);
nand U633 (N_633,In_2208,In_181);
xor U634 (N_634,In_1,In_2312);
and U635 (N_635,In_1654,In_2210);
or U636 (N_636,In_188,In_1002);
xnor U637 (N_637,In_478,In_1677);
or U638 (N_638,In_2895,In_2750);
nor U639 (N_639,In_2860,In_1711);
nand U640 (N_640,In_1324,In_71);
or U641 (N_641,In_1537,In_778);
and U642 (N_642,In_590,In_19);
xor U643 (N_643,In_793,In_799);
and U644 (N_644,In_2317,In_715);
or U645 (N_645,In_743,In_1165);
or U646 (N_646,In_541,In_1796);
nand U647 (N_647,In_1186,In_447);
or U648 (N_648,In_1038,In_2891);
and U649 (N_649,In_1435,In_524);
nor U650 (N_650,In_1868,In_1920);
xor U651 (N_651,In_232,In_2443);
nand U652 (N_652,In_998,In_2542);
nor U653 (N_653,In_518,In_1393);
nor U654 (N_654,In_1974,In_253);
nor U655 (N_655,In_641,In_23);
and U656 (N_656,In_2469,In_1746);
or U657 (N_657,In_2588,In_1792);
xor U658 (N_658,In_1469,In_47);
and U659 (N_659,In_1117,In_2771);
or U660 (N_660,In_1652,In_218);
nor U661 (N_661,In_328,In_1060);
nand U662 (N_662,In_764,In_997);
nand U663 (N_663,In_2460,In_986);
nand U664 (N_664,In_2859,In_2229);
xor U665 (N_665,In_1245,In_2970);
and U666 (N_666,In_68,In_1427);
or U667 (N_667,In_209,In_2089);
xnor U668 (N_668,In_1976,In_2555);
and U669 (N_669,In_1963,In_222);
nand U670 (N_670,In_2773,In_1491);
or U671 (N_671,In_918,In_2468);
or U672 (N_672,In_310,In_2950);
or U673 (N_673,In_2538,In_2351);
or U674 (N_674,In_1098,In_2925);
or U675 (N_675,In_612,In_1836);
and U676 (N_676,In_1008,In_763);
or U677 (N_677,In_1306,In_1334);
or U678 (N_678,In_157,In_2123);
xor U679 (N_679,In_1236,In_443);
nor U680 (N_680,In_566,In_738);
and U681 (N_681,In_247,In_1226);
nand U682 (N_682,In_978,In_753);
and U683 (N_683,In_2060,In_1917);
nand U684 (N_684,In_2105,In_165);
nor U685 (N_685,In_178,In_2196);
and U686 (N_686,In_826,In_2301);
xor U687 (N_687,In_2710,In_287);
and U688 (N_688,In_942,In_1190);
xnor U689 (N_689,In_2080,In_2050);
nand U690 (N_690,In_1105,In_216);
xor U691 (N_691,In_2506,In_1777);
or U692 (N_692,In_876,In_424);
and U693 (N_693,In_2688,In_1498);
xor U694 (N_694,In_1977,In_164);
and U695 (N_695,In_1691,In_450);
nor U696 (N_696,In_548,In_652);
and U697 (N_697,In_2885,In_49);
nand U698 (N_698,In_1995,In_1044);
and U699 (N_699,In_2803,In_981);
nand U700 (N_700,In_749,In_1160);
xnor U701 (N_701,In_702,In_1335);
nand U702 (N_702,In_1921,In_1626);
nor U703 (N_703,In_2098,In_2662);
xnor U704 (N_704,In_1122,In_1896);
nand U705 (N_705,In_2391,In_2474);
nor U706 (N_706,In_698,In_1280);
nor U707 (N_707,In_211,In_2558);
nor U708 (N_708,In_2049,In_1662);
nor U709 (N_709,In_2190,In_2705);
xor U710 (N_710,In_1035,In_448);
nor U711 (N_711,In_2497,In_2473);
nand U712 (N_712,In_693,In_1238);
xnor U713 (N_713,In_2431,In_2533);
nor U714 (N_714,In_2663,In_2573);
xnor U715 (N_715,In_2231,In_1464);
nor U716 (N_716,In_2809,In_768);
xnor U717 (N_717,In_2830,In_2855);
xnor U718 (N_718,In_104,In_2164);
nand U719 (N_719,In_1068,In_1398);
nand U720 (N_720,In_2422,In_699);
or U721 (N_721,In_740,In_2352);
xor U722 (N_722,In_2085,In_2167);
nor U723 (N_723,In_2998,In_1546);
or U724 (N_724,In_2023,In_2315);
xnor U725 (N_725,In_926,In_924);
or U726 (N_726,In_1462,In_2745);
and U727 (N_727,In_1748,In_2837);
or U728 (N_728,In_2685,In_200);
or U729 (N_729,In_354,In_2753);
xnor U730 (N_730,In_1088,In_468);
xnor U731 (N_731,In_2346,In_1232);
and U732 (N_732,In_228,In_587);
nor U733 (N_733,In_2498,In_1477);
or U734 (N_734,In_1725,In_522);
nor U735 (N_735,In_2243,In_12);
and U736 (N_736,In_1919,In_2065);
nand U737 (N_737,In_8,In_1156);
nor U738 (N_738,In_797,In_2886);
nor U739 (N_739,In_201,In_353);
xor U740 (N_740,In_1686,In_2261);
or U741 (N_741,In_1599,In_1409);
nor U742 (N_742,In_1225,In_118);
and U743 (N_743,In_2955,In_1286);
and U744 (N_744,In_1715,In_83);
nor U745 (N_745,In_251,In_705);
nor U746 (N_746,In_144,In_2647);
and U747 (N_747,In_2252,In_1683);
xor U748 (N_748,In_562,In_2137);
xnor U749 (N_749,In_1374,In_833);
or U750 (N_750,In_2381,In_2933);
or U751 (N_751,In_2232,In_2839);
nor U752 (N_752,In_2674,In_1859);
nand U753 (N_753,In_2285,In_2504);
or U754 (N_754,In_825,In_588);
nor U755 (N_755,In_132,In_2612);
nand U756 (N_756,In_2544,In_182);
nand U757 (N_757,In_2496,In_1475);
nand U758 (N_758,In_67,In_653);
or U759 (N_759,In_519,In_807);
nor U760 (N_760,In_1251,In_2805);
nor U761 (N_761,In_1983,In_2202);
xnor U762 (N_762,In_2725,In_732);
nor U763 (N_763,In_2426,In_2419);
or U764 (N_764,In_1946,In_2520);
nor U765 (N_765,In_21,In_1771);
nor U766 (N_766,In_1967,In_2161);
nand U767 (N_767,In_1610,In_323);
and U768 (N_768,In_1965,In_1545);
or U769 (N_769,In_1616,In_539);
xnor U770 (N_770,In_2082,In_2120);
nand U771 (N_771,In_1542,In_2747);
nor U772 (N_772,In_1443,In_6);
nor U773 (N_773,In_2430,In_1015);
and U774 (N_774,In_1529,In_1177);
and U775 (N_775,In_2314,In_2631);
or U776 (N_776,In_1086,In_1310);
nand U777 (N_777,In_989,In_1638);
xnor U778 (N_778,In_2702,In_2323);
nand U779 (N_779,In_1947,In_803);
nand U780 (N_780,In_2835,In_582);
or U781 (N_781,In_2292,In_1929);
and U782 (N_782,In_202,In_1107);
or U783 (N_783,In_236,In_2042);
nand U784 (N_784,In_2532,In_1922);
nand U785 (N_785,In_2151,In_2393);
and U786 (N_786,In_1867,In_1300);
and U787 (N_787,In_681,In_242);
xnor U788 (N_788,In_1694,In_2390);
or U789 (N_789,In_2008,In_2564);
and U790 (N_790,In_1385,In_761);
or U791 (N_791,In_1888,In_2095);
and U792 (N_792,In_1996,In_1479);
xnor U793 (N_793,In_614,In_2963);
nor U794 (N_794,In_2851,In_2967);
nor U795 (N_795,In_2707,In_2759);
nand U796 (N_796,In_1576,In_2719);
and U797 (N_797,In_2905,In_280);
nor U798 (N_798,In_791,In_1285);
and U799 (N_799,In_592,In_2020);
nand U800 (N_800,In_974,In_959);
or U801 (N_801,In_1689,In_632);
nand U802 (N_802,In_2858,In_1962);
and U803 (N_803,In_1080,In_2711);
nor U804 (N_804,In_1472,In_1623);
xor U805 (N_805,In_2609,In_2413);
or U806 (N_806,In_1892,In_2339);
nand U807 (N_807,In_2382,In_31);
nand U808 (N_808,In_2755,In_2143);
and U809 (N_809,In_256,In_1111);
or U810 (N_810,In_1326,In_788);
nor U811 (N_811,In_664,In_1242);
nand U812 (N_812,In_1198,In_2216);
or U813 (N_813,In_2384,In_845);
nor U814 (N_814,In_262,In_1954);
xnor U815 (N_815,In_965,In_2661);
xor U816 (N_816,In_665,In_1101);
xnor U817 (N_817,In_814,In_2103);
xnor U818 (N_818,In_2441,In_909);
or U819 (N_819,In_2626,In_1406);
nand U820 (N_820,In_2876,In_1578);
nor U821 (N_821,In_2941,In_1401);
or U822 (N_822,In_630,In_1214);
xnor U823 (N_823,In_1824,In_921);
and U824 (N_824,In_2144,In_1672);
nand U825 (N_825,In_2428,In_2825);
or U826 (N_826,In_894,In_583);
nor U827 (N_827,In_987,In_719);
and U828 (N_828,In_1175,In_1830);
nand U829 (N_829,In_2621,In_2581);
xor U830 (N_830,In_950,In_271);
xnor U831 (N_831,In_29,In_2079);
nand U832 (N_832,In_265,In_1365);
nand U833 (N_833,In_467,In_1624);
nor U834 (N_834,In_385,In_2016);
or U835 (N_835,In_311,In_2276);
xnor U836 (N_836,In_818,In_1739);
and U837 (N_837,In_1174,In_389);
xnor U838 (N_838,In_413,In_215);
nor U839 (N_839,In_1397,In_2806);
xnor U840 (N_840,In_1185,In_1769);
nand U841 (N_841,In_1866,In_646);
and U842 (N_842,In_1761,In_526);
and U843 (N_843,In_1501,In_1208);
and U844 (N_844,In_98,In_2646);
or U845 (N_845,In_1273,In_1453);
and U846 (N_846,In_2517,In_1992);
nand U847 (N_847,In_1598,In_219);
nand U848 (N_848,In_1357,In_2037);
or U849 (N_849,In_2236,In_1320);
nor U850 (N_850,In_2158,In_2338);
xor U851 (N_851,In_2902,In_760);
or U852 (N_852,In_357,In_2111);
nor U853 (N_853,In_322,In_1282);
xnor U854 (N_854,In_463,In_1264);
xor U855 (N_855,In_2043,In_2324);
and U856 (N_856,In_2385,In_459);
nand U857 (N_857,In_449,In_2543);
nand U858 (N_858,In_469,In_2075);
xnor U859 (N_859,In_2205,In_2959);
nor U860 (N_860,In_2148,In_2454);
xor U861 (N_861,In_608,In_1680);
xor U862 (N_862,In_2618,In_1350);
xnor U863 (N_863,In_79,In_2819);
xor U864 (N_864,In_490,In_1189);
nor U865 (N_865,In_2706,In_1288);
nor U866 (N_866,In_2908,In_1448);
or U867 (N_867,In_2358,In_485);
nand U868 (N_868,In_573,In_1729);
xor U869 (N_869,In_259,In_2913);
and U870 (N_870,In_1941,In_2440);
nor U871 (N_871,In_2975,In_1897);
nand U872 (N_872,In_2594,In_880);
nand U873 (N_873,In_231,In_631);
xnor U874 (N_874,In_334,In_1132);
and U875 (N_875,In_2863,In_1071);
xor U876 (N_876,In_2740,In_1927);
nand U877 (N_877,In_217,In_2119);
xnor U878 (N_878,In_152,In_729);
nand U879 (N_879,In_134,In_1754);
or U880 (N_880,In_2634,In_400);
xor U881 (N_881,In_671,In_809);
nor U882 (N_882,In_441,In_1001);
nor U883 (N_883,In_2653,In_372);
or U884 (N_884,In_728,In_367);
or U885 (N_885,In_176,In_381);
xor U886 (N_886,In_20,In_2185);
xnor U887 (N_887,In_84,In_694);
and U888 (N_888,In_544,In_267);
and U889 (N_889,In_1412,In_712);
and U890 (N_890,In_1265,In_235);
nor U891 (N_891,In_885,In_412);
nand U892 (N_892,In_2389,In_731);
nand U893 (N_893,In_2357,In_2116);
or U894 (N_894,In_2240,In_2515);
nand U895 (N_895,In_2680,In_115);
or U896 (N_896,In_2585,In_1699);
xnor U897 (N_897,In_185,In_1461);
nor U898 (N_898,In_1539,In_1618);
nand U899 (N_899,In_1665,In_1109);
and U900 (N_900,In_240,In_2475);
and U901 (N_901,In_2228,In_2942);
xor U902 (N_902,In_2370,In_899);
nand U903 (N_903,In_2409,In_416);
xor U904 (N_904,In_1369,In_491);
nand U905 (N_905,In_2029,In_1503);
nand U906 (N_906,In_2386,In_2781);
and U907 (N_907,In_2230,In_2106);
or U908 (N_908,In_88,In_557);
nand U909 (N_909,In_1606,In_250);
or U910 (N_910,In_2754,In_269);
nor U911 (N_911,In_2797,In_2999);
nand U912 (N_912,In_1414,In_466);
and U913 (N_913,In_454,In_445);
or U914 (N_914,In_1742,In_832);
xor U915 (N_915,In_789,In_2874);
nand U916 (N_916,In_2465,In_301);
and U917 (N_917,In_1045,In_1580);
or U918 (N_918,In_2220,In_976);
xor U919 (N_919,In_1955,In_2349);
or U920 (N_920,In_1805,In_525);
nand U921 (N_921,In_1220,In_140);
or U922 (N_922,In_1994,In_1893);
or U923 (N_923,In_2084,In_390);
and U924 (N_924,In_1141,In_2604);
xor U925 (N_925,In_2270,In_532);
xnor U926 (N_926,In_505,In_925);
or U927 (N_927,In_2294,In_1512);
and U928 (N_928,In_1561,In_1319);
and U929 (N_929,In_314,In_1140);
xor U930 (N_930,In_966,In_1267);
and U931 (N_931,In_2507,In_56);
or U932 (N_932,In_2854,In_1827);
xor U933 (N_933,In_2484,In_638);
and U934 (N_934,In_85,In_2799);
and U935 (N_935,In_890,In_411);
or U936 (N_936,In_666,In_1839);
nor U937 (N_937,In_1522,In_2954);
nor U938 (N_938,In_2039,In_1644);
nand U939 (N_939,In_1837,In_437);
or U940 (N_940,In_2083,In_2174);
xor U941 (N_941,In_1314,In_2003);
or U942 (N_942,In_2682,In_1482);
and U943 (N_943,In_493,In_1816);
or U944 (N_944,In_1456,In_290);
and U945 (N_945,In_1417,In_2239);
or U946 (N_946,In_2519,In_1883);
or U947 (N_947,In_167,In_303);
nor U948 (N_948,In_2696,In_1352);
and U949 (N_949,In_915,In_1255);
nand U950 (N_950,In_351,In_916);
xor U951 (N_951,In_2919,In_2361);
and U952 (N_952,In_546,In_903);
and U953 (N_953,In_1604,In_2101);
nand U954 (N_954,In_2549,In_1966);
xor U955 (N_955,In_2746,In_2599);
nand U956 (N_956,In_2343,In_1856);
xor U957 (N_957,In_1562,In_1468);
nand U958 (N_958,In_995,In_1237);
or U959 (N_959,In_1569,In_2172);
xnor U960 (N_960,In_1082,In_555);
xor U961 (N_961,In_2843,In_1085);
and U962 (N_962,In_2960,In_2733);
xnor U963 (N_963,In_501,In_2436);
and U964 (N_964,In_2482,In_514);
and U965 (N_965,In_2929,In_46);
and U966 (N_966,In_2818,In_2697);
nand U967 (N_967,In_550,In_238);
nand U968 (N_968,In_1458,In_2211);
or U969 (N_969,In_266,In_2093);
nand U970 (N_970,In_516,In_1770);
xnor U971 (N_971,In_1261,In_1744);
nand U972 (N_972,In_559,In_1271);
nand U973 (N_973,In_439,In_1034);
nor U974 (N_974,In_1870,In_598);
or U975 (N_975,In_1590,In_2363);
nand U976 (N_976,In_2598,In_2224);
or U977 (N_977,In_2036,In_2721);
nor U978 (N_978,In_2155,In_691);
or U979 (N_979,In_2186,In_319);
or U980 (N_980,In_2439,In_1716);
and U981 (N_981,In_1366,In_944);
nand U982 (N_982,In_1169,In_1094);
nor U983 (N_983,In_2847,In_172);
and U984 (N_984,In_2227,In_1120);
nor U985 (N_985,In_1651,In_2310);
and U986 (N_986,In_936,In_1413);
xnor U987 (N_987,In_1704,In_1115);
or U988 (N_988,In_1872,In_1795);
and U989 (N_989,In_2995,In_2511);
or U990 (N_990,In_1822,In_1433);
nor U991 (N_991,In_958,In_1799);
or U992 (N_992,In_2275,In_1331);
or U993 (N_993,In_2813,In_2126);
or U994 (N_994,In_2737,In_379);
and U995 (N_995,In_1370,In_2827);
or U996 (N_996,In_1392,In_220);
xnor U997 (N_997,In_1450,In_1307);
and U998 (N_998,In_510,In_2303);
nand U999 (N_999,In_38,In_545);
xnor U1000 (N_1000,In_820,In_2878);
xor U1001 (N_1001,In_2402,In_1640);
xor U1002 (N_1002,In_1899,In_1224);
xnor U1003 (N_1003,In_2766,In_2990);
nor U1004 (N_1004,In_1808,In_1776);
nand U1005 (N_1005,In_1434,In_1841);
and U1006 (N_1006,In_2910,In_1784);
nand U1007 (N_1007,In_2546,In_1249);
or U1008 (N_1008,In_326,In_2676);
or U1009 (N_1009,In_2704,In_1054);
xnor U1010 (N_1010,In_300,In_408);
and U1011 (N_1011,In_407,In_214);
and U1012 (N_1012,In_1835,In_2522);
or U1013 (N_1013,In_112,In_434);
and U1014 (N_1014,In_2362,In_772);
xnor U1015 (N_1015,In_51,In_1332);
nand U1016 (N_1016,In_1284,In_1146);
xor U1017 (N_1017,In_1336,In_403);
nor U1018 (N_1018,In_777,In_547);
xnor U1019 (N_1019,In_54,In_2836);
nand U1020 (N_1020,In_1077,In_859);
xnor U1021 (N_1021,In_1772,In_1620);
or U1022 (N_1022,In_1497,In_984);
nor U1023 (N_1023,In_57,In_675);
xnor U1024 (N_1024,In_898,In_700);
or U1025 (N_1025,In_375,In_607);
or U1026 (N_1026,In_173,In_2356);
and U1027 (N_1027,In_1702,In_1197);
and U1028 (N_1028,In_1723,In_2399);
or U1029 (N_1029,In_2295,In_1939);
or U1030 (N_1030,In_384,In_1732);
nor U1031 (N_1031,In_2665,In_1577);
xor U1032 (N_1032,In_2115,In_1423);
and U1033 (N_1033,In_1952,In_1269);
or U1034 (N_1034,In_263,In_2640);
and U1035 (N_1035,In_569,In_2994);
nand U1036 (N_1036,In_1812,In_1291);
or U1037 (N_1037,In_1059,In_1391);
nor U1038 (N_1038,In_2102,In_1178);
and U1039 (N_1039,In_2140,In_2459);
nor U1040 (N_1040,In_1864,In_618);
nand U1041 (N_1041,In_1200,In_1124);
nand U1042 (N_1042,In_2068,In_2319);
nand U1043 (N_1043,In_1731,In_1540);
nor U1044 (N_1044,In_1368,In_1137);
nand U1045 (N_1045,In_1708,In_685);
xnor U1046 (N_1046,In_410,In_1216);
and U1047 (N_1047,In_692,In_465);
xnor U1048 (N_1048,In_2046,In_2094);
nor U1049 (N_1049,In_680,In_40);
nor U1050 (N_1050,In_2608,In_444);
nand U1051 (N_1051,In_689,In_1712);
nor U1052 (N_1052,In_1879,In_920);
nand U1053 (N_1053,In_2510,In_2449);
nand U1054 (N_1054,In_395,In_2445);
xor U1055 (N_1055,In_1889,In_2603);
nand U1056 (N_1056,In_2378,In_52);
and U1057 (N_1057,In_192,In_2265);
or U1058 (N_1058,In_2635,In_2250);
nor U1059 (N_1059,In_2117,In_654);
nand U1060 (N_1060,In_1657,In_1834);
nor U1061 (N_1061,In_1668,In_163);
nand U1062 (N_1062,In_961,In_2450);
xnor U1063 (N_1063,In_1895,In_1645);
xnor U1064 (N_1064,In_889,In_1396);
or U1065 (N_1065,In_2823,In_1223);
and U1066 (N_1066,In_805,In_205);
nor U1067 (N_1067,In_1735,In_362);
nand U1068 (N_1068,In_77,In_60);
nand U1069 (N_1069,In_383,In_643);
xor U1070 (N_1070,In_848,In_206);
or U1071 (N_1071,In_1431,In_2214);
and U1072 (N_1072,In_2176,In_1328);
and U1073 (N_1073,In_1459,In_2407);
xnor U1074 (N_1074,In_147,In_1621);
nor U1075 (N_1075,In_1602,In_2015);
or U1076 (N_1076,In_713,In_2421);
xnor U1077 (N_1077,In_1574,In_2909);
or U1078 (N_1078,In_558,In_1572);
xnor U1079 (N_1079,In_1630,In_114);
nor U1080 (N_1080,In_511,In_2692);
nor U1081 (N_1081,In_346,In_2476);
or U1082 (N_1082,In_279,In_1100);
nor U1083 (N_1083,In_660,In_394);
and U1084 (N_1084,In_2637,In_1359);
and U1085 (N_1085,In_2526,In_414);
and U1086 (N_1086,In_1276,In_1709);
xnor U1087 (N_1087,In_260,In_1309);
and U1088 (N_1088,In_856,In_1890);
or U1089 (N_1089,In_1661,In_658);
or U1090 (N_1090,In_870,In_24);
or U1091 (N_1091,In_317,In_2221);
xor U1092 (N_1092,In_717,In_480);
or U1093 (N_1093,In_53,In_684);
xnor U1094 (N_1094,In_1007,In_1909);
nor U1095 (N_1095,In_2848,In_1629);
nor U1096 (N_1096,In_203,In_2628);
and U1097 (N_1097,In_2606,In_2195);
nand U1098 (N_1098,In_1179,In_1455);
nand U1099 (N_1099,In_360,In_617);
or U1100 (N_1100,In_2262,In_234);
nor U1101 (N_1101,In_843,In_2593);
nor U1102 (N_1102,In_1928,In_373);
nand U1103 (N_1103,In_2749,In_171);
or U1104 (N_1104,In_1544,In_1487);
or U1105 (N_1105,In_2873,In_1394);
nand U1106 (N_1106,In_1787,In_281);
or U1107 (N_1107,In_2182,In_2552);
or U1108 (N_1108,In_877,In_2689);
xor U1109 (N_1109,In_2040,In_2879);
and U1110 (N_1110,In_883,In_2904);
nor U1111 (N_1111,In_1125,In_2524);
nand U1112 (N_1112,In_337,In_2764);
nand U1113 (N_1113,In_2986,In_1266);
and U1114 (N_1114,In_2374,In_2783);
nand U1115 (N_1115,In_356,In_1990);
nand U1116 (N_1116,In_2245,In_927);
nor U1117 (N_1117,In_1521,In_655);
nand U1118 (N_1118,In_811,In_1648);
xnor U1119 (N_1119,In_2678,In_1126);
or U1120 (N_1120,In_1948,In_436);
and U1121 (N_1121,In_2957,In_2872);
nor U1122 (N_1122,In_1345,In_1658);
xor U1123 (N_1123,In_186,In_2293);
or U1124 (N_1124,In_1701,In_1774);
xnor U1125 (N_1125,In_2976,In_2486);
or U1126 (N_1126,In_591,In_415);
xnor U1127 (N_1127,In_2681,In_483);
nand U1128 (N_1128,In_420,In_2973);
nand U1129 (N_1129,In_1388,In_1882);
or U1130 (N_1130,In_1766,In_955);
nand U1131 (N_1131,In_1129,In_2620);
and U1132 (N_1132,In_2828,In_2184);
xnor U1133 (N_1133,In_1027,In_1031);
and U1134 (N_1134,In_2022,In_2206);
xor U1135 (N_1135,In_2464,In_1323);
xor U1136 (N_1136,In_1402,In_2371);
and U1137 (N_1137,In_785,In_2728);
nand U1138 (N_1138,In_473,In_1318);
nor U1139 (N_1139,In_1049,In_2547);
xnor U1140 (N_1140,In_873,In_1145);
or U1141 (N_1141,In_2630,In_1914);
nor U1142 (N_1142,In_564,In_2296);
xor U1143 (N_1143,In_1903,In_1213);
nand U1144 (N_1144,In_2365,In_1418);
xor U1145 (N_1145,In_667,In_1183);
xor U1146 (N_1146,In_1985,In_1560);
xor U1147 (N_1147,In_1594,In_2209);
and U1148 (N_1148,In_1083,In_1230);
and U1149 (N_1149,In_336,In_934);
nor U1150 (N_1150,In_751,In_2978);
and U1151 (N_1151,In_776,In_1473);
and U1152 (N_1152,In_2720,In_1346);
xor U1153 (N_1153,In_198,In_423);
xnor U1154 (N_1154,In_1993,In_359);
or U1155 (N_1155,In_2189,In_2530);
or U1156 (N_1156,In_937,In_1989);
nor U1157 (N_1157,In_727,In_2512);
or U1158 (N_1158,In_2898,In_2064);
xor U1159 (N_1159,In_1064,In_61);
nor U1160 (N_1160,In_2279,In_1026);
xor U1161 (N_1161,In_1330,In_2264);
or U1162 (N_1162,In_1628,In_2974);
and U1163 (N_1163,In_2217,In_2736);
or U1164 (N_1164,In_1831,In_1779);
nand U1165 (N_1165,In_1338,In_2713);
nand U1166 (N_1166,In_1614,In_2845);
xnor U1167 (N_1167,In_2045,In_1176);
or U1168 (N_1168,In_1886,In_1018);
xnor U1169 (N_1169,In_1936,In_2067);
and U1170 (N_1170,In_2531,In_2097);
and U1171 (N_1171,In_902,In_530);
nor U1172 (N_1172,In_1706,In_2807);
xnor U1173 (N_1173,In_225,In_1959);
xor U1174 (N_1174,In_2027,In_603);
nor U1175 (N_1175,In_2291,In_1551);
nand U1176 (N_1176,In_813,In_2889);
nor U1177 (N_1177,In_824,In_794);
nand U1178 (N_1178,In_2625,In_2237);
or U1179 (N_1179,In_325,In_1039);
nand U1180 (N_1180,In_1416,In_2657);
nor U1181 (N_1181,In_27,In_1379);
xor U1182 (N_1182,In_1798,In_1643);
nand U1183 (N_1183,In_1613,In_2455);
xnor U1184 (N_1184,In_571,In_63);
and U1185 (N_1185,In_2966,In_428);
nor U1186 (N_1186,In_2633,In_1047);
nand U1187 (N_1187,In_352,In_2574);
nand U1188 (N_1188,In_2703,In_2118);
and U1189 (N_1189,In_2718,In_1173);
and U1190 (N_1190,In_120,In_374);
xor U1191 (N_1191,In_2691,In_742);
and U1192 (N_1192,In_2924,In_2907);
or U1193 (N_1193,In_2028,In_2048);
or U1194 (N_1194,In_2916,In_2617);
nand U1195 (N_1195,In_142,In_156);
or U1196 (N_1196,In_1568,In_906);
nor U1197 (N_1197,In_294,In_1801);
and U1198 (N_1198,In_95,In_1259);
and U1199 (N_1199,In_600,In_1209);
nor U1200 (N_1200,In_1705,In_2723);
xor U1201 (N_1201,In_1021,In_2156);
nand U1202 (N_1202,In_1404,In_1253);
or U1203 (N_1203,In_551,In_2654);
xor U1204 (N_1204,In_1915,In_1356);
nand U1205 (N_1205,In_1517,In_1733);
nand U1206 (N_1206,In_482,In_1429);
and U1207 (N_1207,In_1301,In_2968);
nor U1208 (N_1208,In_1110,In_355);
nor U1209 (N_1209,In_1158,In_901);
xor U1210 (N_1210,In_1876,In_744);
xnor U1211 (N_1211,In_1885,In_1119);
nor U1212 (N_1212,In_964,In_2483);
and U1213 (N_1213,In_914,In_1421);
nor U1214 (N_1214,In_1012,In_2282);
xor U1215 (N_1215,In_912,In_2780);
or U1216 (N_1216,In_1587,In_1978);
and U1217 (N_1217,In_2602,In_2090);
nand U1218 (N_1218,In_1650,In_1019);
nand U1219 (N_1219,In_839,In_1757);
nor U1220 (N_1220,In_2811,In_2325);
or U1221 (N_1221,In_1582,In_1721);
and U1222 (N_1222,In_2700,In_2152);
nor U1223 (N_1223,In_863,In_1681);
or U1224 (N_1224,In_644,In_2677);
xor U1225 (N_1225,In_1949,In_2432);
nand U1226 (N_1226,In_2537,In_1726);
nand U1227 (N_1227,In_382,In_1564);
or U1228 (N_1228,In_2113,In_1439);
nand U1229 (N_1229,In_1337,In_669);
nor U1230 (N_1230,In_2938,In_1855);
or U1231 (N_1231,In_2569,In_1030);
xnor U1232 (N_1232,In_535,In_2991);
nand U1233 (N_1233,In_2269,In_635);
nor U1234 (N_1234,In_1095,In_1693);
nor U1235 (N_1235,In_291,In_2808);
nor U1236 (N_1236,In_1032,In_577);
or U1237 (N_1237,In_2145,In_1833);
nand U1238 (N_1238,In_2613,In_1555);
and U1239 (N_1239,In_1180,In_1363);
and U1240 (N_1240,In_650,In_1290);
nor U1241 (N_1241,In_602,In_2481);
and U1242 (N_1242,In_784,In_835);
nand U1243 (N_1243,In_887,In_2153);
or U1244 (N_1244,In_2142,In_765);
nor U1245 (N_1245,In_1986,In_2605);
nand U1246 (N_1246,In_1719,In_475);
or U1247 (N_1247,In_1373,In_626);
nand U1248 (N_1248,In_35,In_1878);
xnor U1249 (N_1249,In_1250,In_1740);
nand U1250 (N_1250,In_1765,In_1135);
and U1251 (N_1251,In_474,In_2316);
xnor U1252 (N_1252,In_2717,In_1943);
and U1253 (N_1253,In_2335,In_1860);
xor U1254 (N_1254,In_2398,In_892);
nand U1255 (N_1255,In_2918,In_1971);
nand U1256 (N_1256,In_917,In_533);
and U1257 (N_1257,In_1935,In_1813);
nand U1258 (N_1258,In_941,In_601);
nor U1259 (N_1259,In_634,In_335);
and U1260 (N_1260,In_2996,In_1390);
nor U1261 (N_1261,In_369,In_318);
xnor U1262 (N_1262,In_2415,In_1998);
nor U1263 (N_1263,In_2267,In_2107);
nor U1264 (N_1264,In_86,In_1815);
or U1265 (N_1265,In_1646,In_1168);
and U1266 (N_1266,In_64,In_295);
and U1267 (N_1267,In_633,In_2648);
nand U1268 (N_1268,In_2869,In_2666);
xnor U1269 (N_1269,In_639,In_2698);
or U1270 (N_1270,In_1747,In_1006);
and U1271 (N_1271,In_810,In_2794);
nand U1272 (N_1272,In_2170,In_2360);
nand U1273 (N_1273,In_111,In_821);
nand U1274 (N_1274,In_476,In_1956);
or U1275 (N_1275,In_1673,In_2377);
or U1276 (N_1276,In_1800,In_844);
nand U1277 (N_1277,In_780,In_1386);
xnor U1278 (N_1278,In_1381,In_312);
nand U1279 (N_1279,In_2744,In_2639);
nor U1280 (N_1280,In_137,In_160);
nand U1281 (N_1281,In_2234,In_672);
nand U1282 (N_1282,In_1982,In_2516);
nor U1283 (N_1283,In_1601,In_2492);
nand U1284 (N_1284,In_847,In_2139);
and U1285 (N_1285,In_1407,In_1753);
nand U1286 (N_1286,In_606,In_50);
nand U1287 (N_1287,In_2829,In_2299);
xnor U1288 (N_1288,In_92,In_484);
or U1289 (N_1289,In_910,In_370);
nand U1290 (N_1290,In_2795,In_1040);
nand U1291 (N_1291,In_2446,In_2785);
or U1292 (N_1292,In_866,In_2714);
nor U1293 (N_1293,In_2841,In_1440);
nand U1294 (N_1294,In_2572,In_28);
and U1295 (N_1295,In_2896,In_1891);
xor U1296 (N_1296,In_432,In_1973);
and U1297 (N_1297,In_258,In_515);
xnor U1298 (N_1298,In_1298,In_2852);
or U1299 (N_1299,In_1950,In_1348);
xnor U1300 (N_1300,In_2266,In_683);
nand U1301 (N_1301,In_1303,In_1142);
nand U1302 (N_1302,In_2935,In_762);
or U1303 (N_1303,In_1515,In_1720);
and U1304 (N_1304,In_2491,In_2505);
xnor U1305 (N_1305,In_1603,In_2627);
or U1306 (N_1306,In_2006,In_687);
nand U1307 (N_1307,In_2298,In_1164);
or U1308 (N_1308,In_2344,In_1206);
nand U1309 (N_1309,In_75,In_1240);
nor U1310 (N_1310,In_1219,In_2667);
xor U1311 (N_1311,In_2128,In_1103);
nor U1312 (N_1312,In_1631,In_1810);
nand U1313 (N_1313,In_2017,In_316);
xor U1314 (N_1314,In_2972,In_1617);
nor U1315 (N_1315,In_2283,In_492);
xnor U1316 (N_1316,In_2280,In_2038);
nor U1317 (N_1317,In_1519,In_1794);
and U1318 (N_1318,In_2580,In_2871);
and U1319 (N_1319,In_1382,In_2134);
nor U1320 (N_1320,In_604,In_1931);
xor U1321 (N_1321,In_366,In_597);
or U1322 (N_1322,In_1760,In_1538);
nor U1323 (N_1323,In_2397,In_636);
and U1324 (N_1324,In_842,In_521);
nand U1325 (N_1325,In_2932,In_2945);
and U1326 (N_1326,In_1659,In_1764);
and U1327 (N_1327,In_2731,In_252);
or U1328 (N_1328,In_773,In_2273);
and U1329 (N_1329,In_2936,In_2576);
xor U1330 (N_1330,In_932,In_14);
and U1331 (N_1331,In_121,In_2051);
xnor U1332 (N_1332,In_623,In_2290);
and U1333 (N_1333,In_1093,In_166);
nand U1334 (N_1334,In_1520,In_109);
or U1335 (N_1335,In_278,In_162);
or U1336 (N_1336,In_2650,In_567);
xor U1337 (N_1337,In_2253,In_2373);
nor U1338 (N_1338,In_2321,In_975);
or U1339 (N_1339,In_1987,In_1908);
and U1340 (N_1340,In_2388,In_1343);
nand U1341 (N_1341,In_836,In_907);
xor U1342 (N_1342,In_1167,In_2410);
and U1343 (N_1343,In_770,In_819);
xor U1344 (N_1344,In_1690,In_953);
nor U1345 (N_1345,In_2104,In_802);
or U1346 (N_1346,In_2244,In_1806);
and U1347 (N_1347,In_1466,In_123);
xor U1348 (N_1348,In_2562,In_1484);
nor U1349 (N_1349,In_99,In_1938);
or U1350 (N_1350,In_2815,In_2347);
nor U1351 (N_1351,In_1025,In_1913);
nand U1352 (N_1352,In_1395,In_1492);
xor U1353 (N_1353,In_1940,In_1470);
xor U1354 (N_1354,In_1523,In_868);
and U1355 (N_1355,In_827,In_1980);
or U1356 (N_1356,In_440,In_1763);
xnor U1357 (N_1357,In_960,In_2912);
and U1358 (N_1358,In_1865,In_146);
nand U1359 (N_1359,In_405,In_1853);
and U1360 (N_1360,In_862,In_2861);
or U1361 (N_1361,In_647,In_106);
and U1362 (N_1362,In_1106,In_992);
or U1363 (N_1363,In_1997,In_2664);
or U1364 (N_1364,In_1162,In_1637);
xor U1365 (N_1365,In_320,In_204);
nor U1366 (N_1366,In_342,In_1399);
and U1367 (N_1367,In_2649,In_315);
and U1368 (N_1368,In_2485,In_747);
nor U1369 (N_1369,In_2601,In_2988);
and U1370 (N_1370,In_575,In_1478);
xnor U1371 (N_1371,In_1688,In_1153);
and U1372 (N_1372,In_2281,In_282);
nor U1373 (N_1373,In_1246,In_2429);
and U1374 (N_1374,In_2448,In_697);
and U1375 (N_1375,In_2146,In_565);
nand U1376 (N_1376,In_757,In_0);
xor U1377 (N_1377,In_1247,In_1272);
and U1378 (N_1378,In_787,In_2005);
or U1379 (N_1379,In_2756,In_1496);
xnor U1380 (N_1380,In_637,In_2215);
nand U1381 (N_1381,In_2738,In_2178);
nor U1382 (N_1382,In_1229,In_2188);
nor U1383 (N_1383,In_724,In_1170);
nand U1384 (N_1384,In_470,In_994);
or U1385 (N_1385,In_1091,In_2018);
or U1386 (N_1386,In_1633,In_110);
nand U1387 (N_1387,In_402,In_1567);
xnor U1388 (N_1388,In_73,In_2752);
nand U1389 (N_1389,In_1430,In_1239);
xnor U1390 (N_1390,In_2225,In_508);
xor U1391 (N_1391,In_800,In_1655);
nor U1392 (N_1392,In_517,In_1297);
nand U1393 (N_1393,In_2024,In_775);
nand U1394 (N_1394,In_1465,In_1502);
xor U1395 (N_1395,In_2927,In_2461);
or U1396 (N_1396,In_241,In_158);
nor U1397 (N_1397,In_2965,In_1043);
and U1398 (N_1398,In_2956,In_2589);
nor U1399 (N_1399,In_2629,In_2062);
nand U1400 (N_1400,In_2600,In_2540);
nor U1401 (N_1401,In_2376,In_1248);
nor U1402 (N_1402,In_2888,In_2367);
and U1403 (N_1403,In_208,In_1556);
nor U1404 (N_1404,In_1549,In_2078);
nor U1405 (N_1405,In_1445,In_1296);
nor U1406 (N_1406,In_2109,In_2088);
nor U1407 (N_1407,In_347,In_2263);
nand U1408 (N_1408,In_2477,In_1376);
nor U1409 (N_1409,In_977,In_2032);
xor U1410 (N_1410,In_1759,In_2149);
nand U1411 (N_1411,In_2069,In_668);
nand U1412 (N_1412,In_249,In_1207);
or U1413 (N_1413,In_1596,In_2821);
nand U1414 (N_1414,In_2980,In_1845);
xor U1415 (N_1415,In_2306,In_857);
nand U1416 (N_1416,In_1262,In_1089);
and U1417 (N_1417,In_2452,In_2862);
nor U1418 (N_1418,In_2355,In_2679);
nand U1419 (N_1419,In_154,In_988);
or U1420 (N_1420,In_2425,In_387);
or U1421 (N_1421,In_333,In_194);
nand U1422 (N_1422,In_928,In_456);
xor U1423 (N_1423,In_452,In_332);
nand U1424 (N_1424,In_2150,In_1504);
xor U1425 (N_1425,In_2779,In_1786);
or U1426 (N_1426,In_1932,In_1957);
nand U1427 (N_1427,In_1749,In_2000);
nand U1428 (N_1428,In_128,In_769);
nor U1429 (N_1429,In_1696,In_126);
and U1430 (N_1430,In_722,In_1762);
and U1431 (N_1431,In_1530,In_1268);
nand U1432 (N_1432,In_2433,In_2026);
xor U1433 (N_1433,In_540,In_212);
nand U1434 (N_1434,In_2201,In_1710);
or U1435 (N_1435,In_1102,In_951);
or U1436 (N_1436,In_1277,In_11);
and U1437 (N_1437,In_834,In_113);
nand U1438 (N_1438,In_823,In_2168);
xnor U1439 (N_1439,In_2,In_1964);
or U1440 (N_1440,In_1775,In_136);
and U1441 (N_1441,In_1377,In_2193);
xor U1442 (N_1442,In_871,In_1152);
and U1443 (N_1443,In_2897,In_1118);
nor U1444 (N_1444,In_2568,In_1254);
xor U1445 (N_1445,In_2248,In_13);
xnor U1446 (N_1446,In_2288,In_949);
nor U1447 (N_1447,In_1057,In_923);
nor U1448 (N_1448,In_1663,In_1912);
nand U1449 (N_1449,In_2130,In_2488);
nand U1450 (N_1450,In_292,In_2770);
and U1451 (N_1451,In_706,In_125);
nand U1452 (N_1452,In_2566,In_2887);
xor U1453 (N_1453,In_2992,In_1424);
nand U1454 (N_1454,In_1714,In_1311);
and U1455 (N_1455,In_543,In_91);
and U1456 (N_1456,In_908,In_1113);
and U1457 (N_1457,In_2982,In_696);
nor U1458 (N_1458,In_2284,In_2222);
nand U1459 (N_1459,In_481,In_553);
xor U1460 (N_1460,In_513,In_2165);
and U1461 (N_1461,In_2765,In_1906);
xnor U1462 (N_1462,In_893,In_662);
or U1463 (N_1463,In_122,In_596);
xnor U1464 (N_1464,In_1003,In_1581);
nand U1465 (N_1465,In_2414,In_1525);
nor U1466 (N_1466,In_177,In_2890);
and U1467 (N_1467,In_2906,In_1861);
or U1468 (N_1468,In_1743,In_2194);
and U1469 (N_1469,In_2947,In_2197);
and U1470 (N_1470,In_2420,In_418);
or U1471 (N_1471,In_1627,In_1181);
xor U1472 (N_1472,In_2055,In_2337);
xor U1473 (N_1473,In_275,In_556);
nor U1474 (N_1474,In_2840,In_1013);
and U1475 (N_1475,In_2019,In_980);
nor U1476 (N_1476,In_2416,In_1281);
xor U1477 (N_1477,In_947,In_2289);
nand U1478 (N_1478,In_2962,In_1788);
or U1479 (N_1479,In_1066,In_2076);
nand U1480 (N_1480,In_837,In_574);
or U1481 (N_1481,In_895,In_59);
and U1482 (N_1482,In_710,In_534);
nand U1483 (N_1483,In_261,In_2395);
or U1484 (N_1484,In_674,In_1507);
xnor U1485 (N_1485,In_1918,In_911);
xnor U1486 (N_1486,In_289,In_2412);
nor U1487 (N_1487,In_70,In_651);
nor U1488 (N_1488,In_341,In_1734);
or U1489 (N_1489,In_340,In_2985);
and U1490 (N_1490,In_736,In_1625);
or U1491 (N_1491,In_2742,In_1682);
and U1492 (N_1492,In_2434,In_2658);
and U1493 (N_1493,In_1697,In_621);
and U1494 (N_1494,In_1293,In_65);
xnor U1495 (N_1495,In_2478,In_1489);
xnor U1496 (N_1496,In_2557,In_766);
or U1497 (N_1497,In_2392,In_2528);
nand U1498 (N_1498,In_17,In_2548);
nand U1499 (N_1499,In_2007,In_2591);
and U1500 (N_1500,In_982,In_2738);
nand U1501 (N_1501,In_151,In_2215);
or U1502 (N_1502,In_2908,In_1395);
xor U1503 (N_1503,In_1600,In_718);
or U1504 (N_1504,In_2213,In_1763);
and U1505 (N_1505,In_2443,In_2167);
nor U1506 (N_1506,In_795,In_2715);
and U1507 (N_1507,In_1170,In_1595);
or U1508 (N_1508,In_1062,In_1060);
and U1509 (N_1509,In_1859,In_1556);
nor U1510 (N_1510,In_2365,In_2341);
and U1511 (N_1511,In_899,In_1788);
nand U1512 (N_1512,In_1093,In_972);
xor U1513 (N_1513,In_652,In_1255);
and U1514 (N_1514,In_1895,In_2033);
or U1515 (N_1515,In_2131,In_535);
and U1516 (N_1516,In_295,In_1413);
and U1517 (N_1517,In_1218,In_2265);
and U1518 (N_1518,In_511,In_2708);
nand U1519 (N_1519,In_2739,In_1444);
nand U1520 (N_1520,In_1963,In_2690);
nor U1521 (N_1521,In_101,In_2412);
and U1522 (N_1522,In_1221,In_2648);
nor U1523 (N_1523,In_1761,In_284);
nor U1524 (N_1524,In_1705,In_1772);
xor U1525 (N_1525,In_2756,In_1240);
xnor U1526 (N_1526,In_2728,In_1815);
or U1527 (N_1527,In_1468,In_2849);
and U1528 (N_1528,In_640,In_948);
or U1529 (N_1529,In_198,In_2900);
nor U1530 (N_1530,In_710,In_293);
or U1531 (N_1531,In_1312,In_2456);
xnor U1532 (N_1532,In_1429,In_2092);
xor U1533 (N_1533,In_2639,In_2207);
nor U1534 (N_1534,In_916,In_550);
or U1535 (N_1535,In_1257,In_2162);
and U1536 (N_1536,In_2328,In_1069);
and U1537 (N_1537,In_2839,In_756);
nand U1538 (N_1538,In_2080,In_2612);
or U1539 (N_1539,In_2912,In_404);
nand U1540 (N_1540,In_1362,In_311);
nor U1541 (N_1541,In_488,In_1117);
and U1542 (N_1542,In_406,In_629);
or U1543 (N_1543,In_2790,In_1300);
xor U1544 (N_1544,In_790,In_712);
xor U1545 (N_1545,In_1095,In_1493);
nand U1546 (N_1546,In_94,In_1206);
nand U1547 (N_1547,In_2286,In_705);
nor U1548 (N_1548,In_886,In_1196);
nor U1549 (N_1549,In_2467,In_1312);
and U1550 (N_1550,In_1426,In_46);
xnor U1551 (N_1551,In_1283,In_2771);
nor U1552 (N_1552,In_1926,In_2130);
or U1553 (N_1553,In_1762,In_1162);
or U1554 (N_1554,In_1624,In_1772);
xor U1555 (N_1555,In_2530,In_2239);
and U1556 (N_1556,In_248,In_1337);
nor U1557 (N_1557,In_1283,In_843);
or U1558 (N_1558,In_161,In_2674);
and U1559 (N_1559,In_2939,In_1484);
nor U1560 (N_1560,In_1733,In_2257);
or U1561 (N_1561,In_2848,In_645);
and U1562 (N_1562,In_233,In_1912);
xnor U1563 (N_1563,In_2095,In_2651);
nand U1564 (N_1564,In_598,In_460);
and U1565 (N_1565,In_218,In_869);
xor U1566 (N_1566,In_1332,In_143);
nand U1567 (N_1567,In_2643,In_2247);
nand U1568 (N_1568,In_617,In_404);
or U1569 (N_1569,In_773,In_2721);
and U1570 (N_1570,In_2360,In_559);
nor U1571 (N_1571,In_2913,In_2740);
xnor U1572 (N_1572,In_2175,In_460);
nor U1573 (N_1573,In_1429,In_389);
or U1574 (N_1574,In_2353,In_1830);
and U1575 (N_1575,In_2894,In_60);
and U1576 (N_1576,In_2790,In_1412);
or U1577 (N_1577,In_1725,In_1795);
and U1578 (N_1578,In_2512,In_2344);
or U1579 (N_1579,In_1450,In_708);
or U1580 (N_1580,In_2936,In_356);
nand U1581 (N_1581,In_2659,In_2880);
nand U1582 (N_1582,In_433,In_1920);
nand U1583 (N_1583,In_2191,In_1425);
nor U1584 (N_1584,In_85,In_1121);
nand U1585 (N_1585,In_2991,In_352);
nor U1586 (N_1586,In_1455,In_420);
or U1587 (N_1587,In_2011,In_1267);
xnor U1588 (N_1588,In_540,In_2930);
and U1589 (N_1589,In_2088,In_635);
and U1590 (N_1590,In_904,In_961);
and U1591 (N_1591,In_2878,In_2853);
nand U1592 (N_1592,In_317,In_417);
xor U1593 (N_1593,In_2604,In_2287);
nand U1594 (N_1594,In_652,In_1734);
or U1595 (N_1595,In_277,In_647);
or U1596 (N_1596,In_606,In_275);
and U1597 (N_1597,In_2534,In_260);
xnor U1598 (N_1598,In_2561,In_1553);
nor U1599 (N_1599,In_1440,In_2951);
xnor U1600 (N_1600,In_290,In_296);
nand U1601 (N_1601,In_1986,In_2412);
or U1602 (N_1602,In_2257,In_683);
or U1603 (N_1603,In_740,In_2229);
xor U1604 (N_1604,In_1532,In_2236);
nor U1605 (N_1605,In_2501,In_1378);
and U1606 (N_1606,In_640,In_1283);
nor U1607 (N_1607,In_1206,In_1822);
nor U1608 (N_1608,In_715,In_507);
or U1609 (N_1609,In_2516,In_2758);
xor U1610 (N_1610,In_2211,In_2142);
nor U1611 (N_1611,In_509,In_282);
nand U1612 (N_1612,In_2399,In_796);
nor U1613 (N_1613,In_2397,In_1134);
nand U1614 (N_1614,In_1257,In_2103);
or U1615 (N_1615,In_1307,In_1091);
xnor U1616 (N_1616,In_826,In_2467);
or U1617 (N_1617,In_1525,In_1676);
and U1618 (N_1618,In_1703,In_1843);
xnor U1619 (N_1619,In_376,In_802);
and U1620 (N_1620,In_274,In_1639);
nand U1621 (N_1621,In_140,In_1785);
or U1622 (N_1622,In_2175,In_455);
and U1623 (N_1623,In_1073,In_1557);
or U1624 (N_1624,In_513,In_2091);
nand U1625 (N_1625,In_2032,In_1915);
nor U1626 (N_1626,In_2172,In_391);
or U1627 (N_1627,In_1838,In_2323);
and U1628 (N_1628,In_2162,In_1097);
xnor U1629 (N_1629,In_235,In_1030);
xor U1630 (N_1630,In_2786,In_1473);
or U1631 (N_1631,In_673,In_2946);
and U1632 (N_1632,In_133,In_1161);
nand U1633 (N_1633,In_1021,In_438);
or U1634 (N_1634,In_2331,In_2679);
xor U1635 (N_1635,In_1590,In_1602);
or U1636 (N_1636,In_2721,In_159);
nand U1637 (N_1637,In_1529,In_1094);
nand U1638 (N_1638,In_1393,In_1945);
nor U1639 (N_1639,In_847,In_2425);
nand U1640 (N_1640,In_42,In_473);
nand U1641 (N_1641,In_2072,In_1037);
nor U1642 (N_1642,In_2729,In_820);
xor U1643 (N_1643,In_2485,In_1707);
nand U1644 (N_1644,In_308,In_1892);
nand U1645 (N_1645,In_869,In_856);
or U1646 (N_1646,In_971,In_1743);
nand U1647 (N_1647,In_1232,In_2257);
and U1648 (N_1648,In_1505,In_469);
nor U1649 (N_1649,In_1095,In_2736);
xor U1650 (N_1650,In_235,In_1126);
and U1651 (N_1651,In_2290,In_1703);
nor U1652 (N_1652,In_933,In_2258);
or U1653 (N_1653,In_2524,In_2024);
xnor U1654 (N_1654,In_350,In_1403);
xnor U1655 (N_1655,In_541,In_1322);
and U1656 (N_1656,In_722,In_2720);
or U1657 (N_1657,In_1077,In_567);
xnor U1658 (N_1658,In_2674,In_1304);
nor U1659 (N_1659,In_1261,In_1254);
or U1660 (N_1660,In_2925,In_533);
nor U1661 (N_1661,In_856,In_2465);
nand U1662 (N_1662,In_448,In_614);
or U1663 (N_1663,In_2177,In_1096);
nor U1664 (N_1664,In_396,In_1570);
nor U1665 (N_1665,In_1309,In_1996);
nand U1666 (N_1666,In_1477,In_1084);
and U1667 (N_1667,In_1495,In_765);
and U1668 (N_1668,In_2124,In_1802);
and U1669 (N_1669,In_262,In_1913);
or U1670 (N_1670,In_258,In_1893);
or U1671 (N_1671,In_2890,In_2344);
or U1672 (N_1672,In_1805,In_2386);
xor U1673 (N_1673,In_891,In_1498);
or U1674 (N_1674,In_400,In_2325);
and U1675 (N_1675,In_47,In_1582);
or U1676 (N_1676,In_1746,In_2103);
and U1677 (N_1677,In_1896,In_2216);
xnor U1678 (N_1678,In_1011,In_1335);
and U1679 (N_1679,In_2850,In_1888);
or U1680 (N_1680,In_1943,In_1115);
nor U1681 (N_1681,In_898,In_611);
xor U1682 (N_1682,In_1658,In_1606);
and U1683 (N_1683,In_479,In_1456);
or U1684 (N_1684,In_620,In_1335);
nand U1685 (N_1685,In_2119,In_336);
nand U1686 (N_1686,In_1746,In_2794);
and U1687 (N_1687,In_896,In_971);
xnor U1688 (N_1688,In_2680,In_85);
xnor U1689 (N_1689,In_1138,In_2933);
xor U1690 (N_1690,In_1301,In_1911);
and U1691 (N_1691,In_1869,In_80);
or U1692 (N_1692,In_2869,In_2823);
nand U1693 (N_1693,In_1108,In_692);
xor U1694 (N_1694,In_33,In_375);
and U1695 (N_1695,In_599,In_86);
or U1696 (N_1696,In_2429,In_1203);
xnor U1697 (N_1697,In_2144,In_1892);
or U1698 (N_1698,In_1703,In_2141);
or U1699 (N_1699,In_1598,In_281);
or U1700 (N_1700,In_950,In_652);
xnor U1701 (N_1701,In_1,In_2402);
or U1702 (N_1702,In_1346,In_234);
and U1703 (N_1703,In_795,In_593);
or U1704 (N_1704,In_2068,In_281);
or U1705 (N_1705,In_2556,In_2061);
nor U1706 (N_1706,In_1719,In_215);
xnor U1707 (N_1707,In_1274,In_1179);
xor U1708 (N_1708,In_2730,In_480);
and U1709 (N_1709,In_519,In_1515);
or U1710 (N_1710,In_1356,In_1711);
nor U1711 (N_1711,In_1877,In_2627);
xor U1712 (N_1712,In_934,In_1178);
nand U1713 (N_1713,In_2947,In_530);
nand U1714 (N_1714,In_760,In_798);
nor U1715 (N_1715,In_1198,In_1207);
nor U1716 (N_1716,In_2625,In_389);
and U1717 (N_1717,In_1273,In_2726);
xnor U1718 (N_1718,In_2430,In_2361);
nand U1719 (N_1719,In_862,In_2186);
nor U1720 (N_1720,In_327,In_1008);
nand U1721 (N_1721,In_1958,In_133);
xor U1722 (N_1722,In_1577,In_542);
or U1723 (N_1723,In_635,In_2880);
xor U1724 (N_1724,In_1572,In_1039);
nor U1725 (N_1725,In_2363,In_740);
or U1726 (N_1726,In_1924,In_2690);
xor U1727 (N_1727,In_1651,In_1347);
nand U1728 (N_1728,In_1643,In_2054);
nor U1729 (N_1729,In_698,In_1578);
or U1730 (N_1730,In_2124,In_1112);
nand U1731 (N_1731,In_1174,In_1068);
and U1732 (N_1732,In_1080,In_898);
nand U1733 (N_1733,In_2535,In_1279);
nand U1734 (N_1734,In_1647,In_830);
and U1735 (N_1735,In_1616,In_2860);
xnor U1736 (N_1736,In_1739,In_1992);
nor U1737 (N_1737,In_2590,In_539);
and U1738 (N_1738,In_212,In_237);
xor U1739 (N_1739,In_1139,In_1365);
nand U1740 (N_1740,In_933,In_985);
nor U1741 (N_1741,In_2795,In_205);
and U1742 (N_1742,In_1949,In_974);
nor U1743 (N_1743,In_1631,In_915);
and U1744 (N_1744,In_114,In_2197);
or U1745 (N_1745,In_61,In_373);
or U1746 (N_1746,In_2490,In_1742);
nor U1747 (N_1747,In_2521,In_2112);
nand U1748 (N_1748,In_1451,In_145);
nand U1749 (N_1749,In_1821,In_1175);
and U1750 (N_1750,In_2716,In_2081);
xor U1751 (N_1751,In_2861,In_594);
nor U1752 (N_1752,In_1706,In_2112);
xor U1753 (N_1753,In_506,In_913);
nor U1754 (N_1754,In_1743,In_451);
or U1755 (N_1755,In_2913,In_2020);
xor U1756 (N_1756,In_942,In_225);
or U1757 (N_1757,In_1514,In_1598);
or U1758 (N_1758,In_296,In_2832);
and U1759 (N_1759,In_2417,In_973);
nand U1760 (N_1760,In_2836,In_229);
nand U1761 (N_1761,In_1761,In_2199);
nor U1762 (N_1762,In_887,In_1085);
or U1763 (N_1763,In_2723,In_760);
nor U1764 (N_1764,In_1620,In_447);
or U1765 (N_1765,In_2005,In_2531);
nand U1766 (N_1766,In_719,In_738);
nor U1767 (N_1767,In_339,In_1960);
xor U1768 (N_1768,In_2578,In_438);
nand U1769 (N_1769,In_1096,In_1638);
xor U1770 (N_1770,In_997,In_1297);
and U1771 (N_1771,In_492,In_573);
or U1772 (N_1772,In_957,In_2853);
and U1773 (N_1773,In_2885,In_1574);
xnor U1774 (N_1774,In_745,In_1598);
and U1775 (N_1775,In_703,In_485);
xor U1776 (N_1776,In_973,In_1546);
and U1777 (N_1777,In_1163,In_2550);
and U1778 (N_1778,In_427,In_1467);
or U1779 (N_1779,In_241,In_2007);
or U1780 (N_1780,In_639,In_30);
nor U1781 (N_1781,In_820,In_700);
xor U1782 (N_1782,In_734,In_812);
or U1783 (N_1783,In_707,In_2520);
nand U1784 (N_1784,In_1403,In_887);
and U1785 (N_1785,In_2224,In_266);
and U1786 (N_1786,In_481,In_1625);
or U1787 (N_1787,In_2145,In_2579);
nor U1788 (N_1788,In_2022,In_1487);
nor U1789 (N_1789,In_543,In_2653);
or U1790 (N_1790,In_2930,In_2476);
nor U1791 (N_1791,In_839,In_2405);
nor U1792 (N_1792,In_2424,In_1924);
or U1793 (N_1793,In_439,In_2843);
or U1794 (N_1794,In_2704,In_979);
nand U1795 (N_1795,In_1305,In_1233);
or U1796 (N_1796,In_2231,In_635);
nor U1797 (N_1797,In_656,In_2418);
xnor U1798 (N_1798,In_2659,In_1042);
nor U1799 (N_1799,In_1957,In_850);
and U1800 (N_1800,In_723,In_2197);
nand U1801 (N_1801,In_209,In_2682);
nor U1802 (N_1802,In_207,In_1012);
nand U1803 (N_1803,In_692,In_943);
and U1804 (N_1804,In_254,In_2793);
nor U1805 (N_1805,In_430,In_1443);
nand U1806 (N_1806,In_1048,In_1580);
or U1807 (N_1807,In_2538,In_426);
or U1808 (N_1808,In_2300,In_1409);
nor U1809 (N_1809,In_434,In_1416);
nor U1810 (N_1810,In_2464,In_2143);
nand U1811 (N_1811,In_1268,In_1469);
nand U1812 (N_1812,In_701,In_2441);
and U1813 (N_1813,In_2948,In_590);
nor U1814 (N_1814,In_246,In_381);
or U1815 (N_1815,In_596,In_762);
xnor U1816 (N_1816,In_1866,In_1162);
and U1817 (N_1817,In_1735,In_1217);
nand U1818 (N_1818,In_152,In_2975);
xor U1819 (N_1819,In_1023,In_2769);
or U1820 (N_1820,In_2486,In_2851);
nor U1821 (N_1821,In_804,In_1300);
xor U1822 (N_1822,In_2428,In_673);
or U1823 (N_1823,In_1991,In_1980);
nand U1824 (N_1824,In_1545,In_940);
xnor U1825 (N_1825,In_1857,In_1336);
xor U1826 (N_1826,In_917,In_1571);
nor U1827 (N_1827,In_79,In_38);
or U1828 (N_1828,In_1080,In_2479);
nor U1829 (N_1829,In_742,In_1706);
nor U1830 (N_1830,In_2022,In_1653);
or U1831 (N_1831,In_2150,In_216);
xor U1832 (N_1832,In_2849,In_871);
or U1833 (N_1833,In_945,In_429);
and U1834 (N_1834,In_1649,In_1238);
xnor U1835 (N_1835,In_2394,In_827);
and U1836 (N_1836,In_530,In_969);
nor U1837 (N_1837,In_1118,In_438);
nand U1838 (N_1838,In_2658,In_732);
nand U1839 (N_1839,In_2769,In_2948);
and U1840 (N_1840,In_26,In_2779);
and U1841 (N_1841,In_977,In_322);
or U1842 (N_1842,In_2446,In_558);
nor U1843 (N_1843,In_766,In_906);
nand U1844 (N_1844,In_743,In_1688);
or U1845 (N_1845,In_1235,In_1045);
or U1846 (N_1846,In_1155,In_6);
nand U1847 (N_1847,In_109,In_125);
nand U1848 (N_1848,In_1688,In_1832);
nand U1849 (N_1849,In_1665,In_2764);
nand U1850 (N_1850,In_491,In_2853);
nand U1851 (N_1851,In_1519,In_1363);
nand U1852 (N_1852,In_389,In_491);
nor U1853 (N_1853,In_132,In_1018);
or U1854 (N_1854,In_2422,In_830);
nand U1855 (N_1855,In_2267,In_1259);
xor U1856 (N_1856,In_2975,In_400);
nor U1857 (N_1857,In_294,In_527);
nor U1858 (N_1858,In_2572,In_2597);
nor U1859 (N_1859,In_1893,In_154);
nand U1860 (N_1860,In_1329,In_733);
xnor U1861 (N_1861,In_2239,In_2801);
or U1862 (N_1862,In_1319,In_578);
nor U1863 (N_1863,In_2855,In_2927);
or U1864 (N_1864,In_1503,In_1310);
nor U1865 (N_1865,In_1168,In_1998);
nor U1866 (N_1866,In_2707,In_1120);
nand U1867 (N_1867,In_955,In_2786);
nand U1868 (N_1868,In_808,In_2028);
and U1869 (N_1869,In_2145,In_1985);
xor U1870 (N_1870,In_1214,In_194);
nand U1871 (N_1871,In_411,In_922);
nand U1872 (N_1872,In_2888,In_323);
nor U1873 (N_1873,In_1412,In_131);
xnor U1874 (N_1874,In_1071,In_2880);
nand U1875 (N_1875,In_2606,In_1918);
nor U1876 (N_1876,In_2882,In_2438);
nand U1877 (N_1877,In_1157,In_1091);
nand U1878 (N_1878,In_1569,In_1294);
nand U1879 (N_1879,In_2278,In_187);
xor U1880 (N_1880,In_1207,In_1586);
nand U1881 (N_1881,In_2210,In_980);
nor U1882 (N_1882,In_1090,In_1502);
nand U1883 (N_1883,In_454,In_1147);
nor U1884 (N_1884,In_2305,In_2428);
and U1885 (N_1885,In_1239,In_1753);
and U1886 (N_1886,In_938,In_1268);
nand U1887 (N_1887,In_2517,In_673);
nor U1888 (N_1888,In_1129,In_2285);
or U1889 (N_1889,In_2014,In_2015);
nand U1890 (N_1890,In_2834,In_2915);
and U1891 (N_1891,In_295,In_2036);
and U1892 (N_1892,In_419,In_76);
nand U1893 (N_1893,In_1094,In_195);
xnor U1894 (N_1894,In_817,In_2880);
nor U1895 (N_1895,In_99,In_2895);
or U1896 (N_1896,In_26,In_619);
xnor U1897 (N_1897,In_1891,In_1215);
xor U1898 (N_1898,In_37,In_97);
xor U1899 (N_1899,In_311,In_485);
nor U1900 (N_1900,In_1080,In_2788);
nor U1901 (N_1901,In_771,In_557);
nand U1902 (N_1902,In_1158,In_382);
nand U1903 (N_1903,In_1373,In_1208);
or U1904 (N_1904,In_2581,In_948);
and U1905 (N_1905,In_1848,In_2068);
xor U1906 (N_1906,In_2093,In_1514);
and U1907 (N_1907,In_1316,In_935);
nor U1908 (N_1908,In_758,In_1700);
and U1909 (N_1909,In_1911,In_1901);
nand U1910 (N_1910,In_2042,In_212);
or U1911 (N_1911,In_2581,In_1536);
nand U1912 (N_1912,In_1861,In_1268);
and U1913 (N_1913,In_1100,In_2567);
nand U1914 (N_1914,In_352,In_1148);
xor U1915 (N_1915,In_1036,In_2886);
and U1916 (N_1916,In_2658,In_2870);
nor U1917 (N_1917,In_174,In_1086);
nand U1918 (N_1918,In_2687,In_83);
and U1919 (N_1919,In_2549,In_1838);
nand U1920 (N_1920,In_569,In_2531);
and U1921 (N_1921,In_2962,In_2632);
xor U1922 (N_1922,In_763,In_1984);
and U1923 (N_1923,In_1829,In_2660);
nor U1924 (N_1924,In_2516,In_1694);
xnor U1925 (N_1925,In_970,In_371);
or U1926 (N_1926,In_1919,In_365);
nand U1927 (N_1927,In_2994,In_1509);
xor U1928 (N_1928,In_2187,In_203);
or U1929 (N_1929,In_1283,In_2897);
and U1930 (N_1930,In_2860,In_510);
nor U1931 (N_1931,In_2838,In_1868);
nor U1932 (N_1932,In_2503,In_1757);
xor U1933 (N_1933,In_299,In_393);
or U1934 (N_1934,In_1050,In_2933);
xnor U1935 (N_1935,In_2078,In_138);
and U1936 (N_1936,In_2394,In_2336);
nand U1937 (N_1937,In_1356,In_872);
or U1938 (N_1938,In_2600,In_950);
nor U1939 (N_1939,In_668,In_1307);
nor U1940 (N_1940,In_287,In_665);
nor U1941 (N_1941,In_635,In_1085);
nor U1942 (N_1942,In_1786,In_589);
nor U1943 (N_1943,In_2762,In_2781);
xnor U1944 (N_1944,In_1100,In_2438);
nor U1945 (N_1945,In_80,In_2545);
or U1946 (N_1946,In_2959,In_1387);
and U1947 (N_1947,In_471,In_2731);
xnor U1948 (N_1948,In_2440,In_2576);
or U1949 (N_1949,In_2619,In_147);
and U1950 (N_1950,In_2013,In_780);
and U1951 (N_1951,In_1006,In_939);
or U1952 (N_1952,In_2497,In_1831);
or U1953 (N_1953,In_1450,In_2475);
xnor U1954 (N_1954,In_1149,In_648);
xor U1955 (N_1955,In_2350,In_1496);
xnor U1956 (N_1956,In_577,In_2232);
and U1957 (N_1957,In_1649,In_1582);
nor U1958 (N_1958,In_1918,In_82);
nor U1959 (N_1959,In_2009,In_2228);
nor U1960 (N_1960,In_404,In_512);
and U1961 (N_1961,In_2900,In_837);
and U1962 (N_1962,In_2947,In_1039);
or U1963 (N_1963,In_1621,In_1375);
and U1964 (N_1964,In_1737,In_1121);
nand U1965 (N_1965,In_2590,In_1356);
and U1966 (N_1966,In_311,In_1370);
nand U1967 (N_1967,In_90,In_2225);
nand U1968 (N_1968,In_2386,In_2208);
and U1969 (N_1969,In_2213,In_2302);
xor U1970 (N_1970,In_700,In_2552);
nand U1971 (N_1971,In_2704,In_573);
xor U1972 (N_1972,In_2754,In_108);
nand U1973 (N_1973,In_2443,In_1099);
or U1974 (N_1974,In_950,In_2105);
nor U1975 (N_1975,In_1510,In_1560);
xnor U1976 (N_1976,In_2107,In_643);
nand U1977 (N_1977,In_1933,In_2627);
and U1978 (N_1978,In_150,In_2563);
and U1979 (N_1979,In_530,In_878);
nand U1980 (N_1980,In_1779,In_1802);
nand U1981 (N_1981,In_406,In_1799);
nor U1982 (N_1982,In_583,In_2682);
or U1983 (N_1983,In_1349,In_1359);
nor U1984 (N_1984,In_1164,In_2668);
and U1985 (N_1985,In_895,In_3);
nand U1986 (N_1986,In_1541,In_2156);
and U1987 (N_1987,In_1630,In_2205);
nor U1988 (N_1988,In_2708,In_553);
nand U1989 (N_1989,In_2329,In_2012);
or U1990 (N_1990,In_2445,In_1962);
or U1991 (N_1991,In_1115,In_1786);
nor U1992 (N_1992,In_2021,In_1619);
xnor U1993 (N_1993,In_615,In_1876);
and U1994 (N_1994,In_2574,In_1336);
nand U1995 (N_1995,In_1295,In_726);
and U1996 (N_1996,In_2759,In_1520);
and U1997 (N_1997,In_2982,In_1893);
xor U1998 (N_1998,In_2811,In_154);
xor U1999 (N_1999,In_2188,In_2903);
nand U2000 (N_2000,In_2673,In_480);
nand U2001 (N_2001,In_2242,In_452);
and U2002 (N_2002,In_2232,In_2427);
nand U2003 (N_2003,In_2872,In_2411);
nor U2004 (N_2004,In_1881,In_130);
and U2005 (N_2005,In_988,In_1267);
xnor U2006 (N_2006,In_2565,In_2050);
and U2007 (N_2007,In_557,In_2541);
and U2008 (N_2008,In_2654,In_1329);
nor U2009 (N_2009,In_859,In_1154);
or U2010 (N_2010,In_1106,In_102);
nor U2011 (N_2011,In_926,In_2203);
or U2012 (N_2012,In_1833,In_1687);
nand U2013 (N_2013,In_527,In_171);
or U2014 (N_2014,In_2923,In_1140);
or U2015 (N_2015,In_2001,In_2918);
or U2016 (N_2016,In_1425,In_101);
xnor U2017 (N_2017,In_2104,In_2581);
or U2018 (N_2018,In_726,In_1967);
or U2019 (N_2019,In_1450,In_1380);
and U2020 (N_2020,In_380,In_2106);
xnor U2021 (N_2021,In_2498,In_1177);
and U2022 (N_2022,In_755,In_753);
nand U2023 (N_2023,In_2749,In_2417);
nor U2024 (N_2024,In_2563,In_2543);
and U2025 (N_2025,In_2765,In_744);
nand U2026 (N_2026,In_1572,In_457);
nor U2027 (N_2027,In_1364,In_328);
xnor U2028 (N_2028,In_1902,In_2085);
xor U2029 (N_2029,In_1382,In_2440);
xnor U2030 (N_2030,In_1121,In_2384);
nand U2031 (N_2031,In_434,In_351);
nand U2032 (N_2032,In_1435,In_2424);
nand U2033 (N_2033,In_1816,In_800);
nand U2034 (N_2034,In_1387,In_32);
or U2035 (N_2035,In_442,In_1944);
nand U2036 (N_2036,In_1547,In_1631);
nand U2037 (N_2037,In_737,In_1779);
xor U2038 (N_2038,In_1550,In_2593);
and U2039 (N_2039,In_1868,In_2140);
xor U2040 (N_2040,In_1778,In_2323);
or U2041 (N_2041,In_674,In_703);
xnor U2042 (N_2042,In_396,In_2279);
xnor U2043 (N_2043,In_2984,In_1578);
or U2044 (N_2044,In_328,In_1341);
xnor U2045 (N_2045,In_1072,In_461);
nand U2046 (N_2046,In_2141,In_231);
and U2047 (N_2047,In_2439,In_678);
or U2048 (N_2048,In_612,In_2580);
nand U2049 (N_2049,In_1872,In_1879);
nand U2050 (N_2050,In_1671,In_735);
xnor U2051 (N_2051,In_1355,In_2464);
nand U2052 (N_2052,In_56,In_2391);
or U2053 (N_2053,In_2275,In_2829);
nor U2054 (N_2054,In_236,In_66);
nand U2055 (N_2055,In_1661,In_175);
nor U2056 (N_2056,In_1276,In_1423);
nand U2057 (N_2057,In_2397,In_2819);
nand U2058 (N_2058,In_389,In_1554);
or U2059 (N_2059,In_657,In_142);
and U2060 (N_2060,In_931,In_2518);
nand U2061 (N_2061,In_799,In_1607);
nand U2062 (N_2062,In_1347,In_2848);
or U2063 (N_2063,In_2113,In_1816);
or U2064 (N_2064,In_564,In_68);
and U2065 (N_2065,In_1585,In_2391);
or U2066 (N_2066,In_2429,In_550);
or U2067 (N_2067,In_1547,In_2494);
or U2068 (N_2068,In_375,In_589);
or U2069 (N_2069,In_98,In_1845);
or U2070 (N_2070,In_2908,In_2573);
or U2071 (N_2071,In_2179,In_2651);
or U2072 (N_2072,In_751,In_2773);
nand U2073 (N_2073,In_1448,In_2604);
nor U2074 (N_2074,In_1154,In_1186);
or U2075 (N_2075,In_325,In_1371);
xor U2076 (N_2076,In_698,In_2578);
and U2077 (N_2077,In_450,In_1756);
or U2078 (N_2078,In_636,In_2888);
or U2079 (N_2079,In_2373,In_2091);
or U2080 (N_2080,In_662,In_117);
or U2081 (N_2081,In_2427,In_474);
nor U2082 (N_2082,In_1432,In_150);
xnor U2083 (N_2083,In_762,In_2642);
nand U2084 (N_2084,In_2036,In_2926);
xor U2085 (N_2085,In_1064,In_382);
and U2086 (N_2086,In_1527,In_980);
xor U2087 (N_2087,In_2763,In_779);
xnor U2088 (N_2088,In_173,In_359);
nand U2089 (N_2089,In_1742,In_583);
nor U2090 (N_2090,In_2686,In_1986);
or U2091 (N_2091,In_2863,In_1072);
nor U2092 (N_2092,In_2659,In_1457);
xnor U2093 (N_2093,In_1573,In_1758);
xnor U2094 (N_2094,In_2727,In_194);
xor U2095 (N_2095,In_2063,In_351);
or U2096 (N_2096,In_489,In_2456);
nand U2097 (N_2097,In_1147,In_1958);
or U2098 (N_2098,In_2408,In_1208);
and U2099 (N_2099,In_2054,In_1622);
or U2100 (N_2100,In_1786,In_1438);
or U2101 (N_2101,In_2384,In_985);
and U2102 (N_2102,In_1945,In_2023);
nor U2103 (N_2103,In_149,In_2871);
nand U2104 (N_2104,In_1818,In_630);
xor U2105 (N_2105,In_1348,In_2618);
xor U2106 (N_2106,In_543,In_2614);
xnor U2107 (N_2107,In_2358,In_1601);
and U2108 (N_2108,In_1873,In_2905);
xor U2109 (N_2109,In_922,In_2484);
or U2110 (N_2110,In_2963,In_1102);
nor U2111 (N_2111,In_639,In_1425);
or U2112 (N_2112,In_2599,In_1025);
xor U2113 (N_2113,In_1854,In_178);
nand U2114 (N_2114,In_1978,In_63);
nor U2115 (N_2115,In_2040,In_1454);
and U2116 (N_2116,In_1150,In_754);
nand U2117 (N_2117,In_1411,In_1596);
and U2118 (N_2118,In_2352,In_1499);
xor U2119 (N_2119,In_835,In_1422);
nand U2120 (N_2120,In_903,In_302);
and U2121 (N_2121,In_1998,In_1792);
xor U2122 (N_2122,In_1076,In_2872);
or U2123 (N_2123,In_999,In_555);
nor U2124 (N_2124,In_2093,In_2396);
xor U2125 (N_2125,In_608,In_941);
or U2126 (N_2126,In_696,In_169);
or U2127 (N_2127,In_1212,In_1651);
nand U2128 (N_2128,In_2770,In_49);
nand U2129 (N_2129,In_531,In_263);
and U2130 (N_2130,In_1030,In_1325);
xor U2131 (N_2131,In_1893,In_2626);
nand U2132 (N_2132,In_144,In_2531);
xor U2133 (N_2133,In_1410,In_192);
or U2134 (N_2134,In_659,In_969);
and U2135 (N_2135,In_389,In_1519);
and U2136 (N_2136,In_2711,In_2915);
or U2137 (N_2137,In_2657,In_1360);
nand U2138 (N_2138,In_235,In_730);
and U2139 (N_2139,In_1451,In_1844);
xnor U2140 (N_2140,In_648,In_1296);
nand U2141 (N_2141,In_1861,In_2619);
nor U2142 (N_2142,In_1488,In_2834);
nand U2143 (N_2143,In_2532,In_2386);
or U2144 (N_2144,In_590,In_2088);
nor U2145 (N_2145,In_2764,In_2474);
and U2146 (N_2146,In_1908,In_2406);
nand U2147 (N_2147,In_2563,In_1094);
nand U2148 (N_2148,In_1030,In_1244);
nand U2149 (N_2149,In_2872,In_2976);
and U2150 (N_2150,In_567,In_2538);
xor U2151 (N_2151,In_2278,In_896);
nor U2152 (N_2152,In_1432,In_1804);
or U2153 (N_2153,In_234,In_1641);
xnor U2154 (N_2154,In_1368,In_1355);
nor U2155 (N_2155,In_982,In_906);
nor U2156 (N_2156,In_989,In_1119);
xnor U2157 (N_2157,In_1784,In_1603);
nor U2158 (N_2158,In_2074,In_1818);
xnor U2159 (N_2159,In_2667,In_566);
xor U2160 (N_2160,In_2952,In_596);
nand U2161 (N_2161,In_370,In_570);
nand U2162 (N_2162,In_1720,In_2655);
or U2163 (N_2163,In_27,In_672);
or U2164 (N_2164,In_1957,In_2817);
nand U2165 (N_2165,In_2703,In_692);
nand U2166 (N_2166,In_57,In_1272);
nor U2167 (N_2167,In_954,In_816);
or U2168 (N_2168,In_2511,In_350);
or U2169 (N_2169,In_699,In_734);
or U2170 (N_2170,In_2359,In_235);
xnor U2171 (N_2171,In_2340,In_2004);
and U2172 (N_2172,In_210,In_1839);
xnor U2173 (N_2173,In_436,In_2345);
nor U2174 (N_2174,In_2045,In_452);
nand U2175 (N_2175,In_2338,In_1772);
nand U2176 (N_2176,In_1005,In_2140);
xnor U2177 (N_2177,In_1201,In_326);
xor U2178 (N_2178,In_1580,In_1617);
and U2179 (N_2179,In_235,In_1021);
nor U2180 (N_2180,In_1090,In_1666);
and U2181 (N_2181,In_54,In_641);
and U2182 (N_2182,In_90,In_834);
xor U2183 (N_2183,In_1285,In_956);
nor U2184 (N_2184,In_1972,In_1856);
nand U2185 (N_2185,In_1978,In_305);
and U2186 (N_2186,In_1100,In_1060);
nand U2187 (N_2187,In_704,In_898);
and U2188 (N_2188,In_1828,In_1044);
and U2189 (N_2189,In_802,In_1015);
nor U2190 (N_2190,In_1229,In_356);
or U2191 (N_2191,In_1906,In_2227);
nor U2192 (N_2192,In_1569,In_2478);
xor U2193 (N_2193,In_663,In_2548);
xor U2194 (N_2194,In_1392,In_1456);
nor U2195 (N_2195,In_653,In_1010);
and U2196 (N_2196,In_2455,In_1597);
nand U2197 (N_2197,In_1745,In_1604);
nand U2198 (N_2198,In_352,In_1835);
nor U2199 (N_2199,In_422,In_1932);
or U2200 (N_2200,In_905,In_2923);
or U2201 (N_2201,In_870,In_1770);
or U2202 (N_2202,In_946,In_327);
xor U2203 (N_2203,In_278,In_1698);
nand U2204 (N_2204,In_109,In_1177);
or U2205 (N_2205,In_113,In_539);
xor U2206 (N_2206,In_770,In_1618);
and U2207 (N_2207,In_1775,In_123);
nor U2208 (N_2208,In_4,In_1448);
xor U2209 (N_2209,In_664,In_1383);
nor U2210 (N_2210,In_2908,In_1333);
nor U2211 (N_2211,In_963,In_801);
or U2212 (N_2212,In_976,In_1913);
xor U2213 (N_2213,In_91,In_27);
nor U2214 (N_2214,In_2091,In_1016);
nand U2215 (N_2215,In_2065,In_2707);
or U2216 (N_2216,In_1361,In_1302);
or U2217 (N_2217,In_1816,In_834);
nor U2218 (N_2218,In_601,In_1588);
and U2219 (N_2219,In_2506,In_2201);
nor U2220 (N_2220,In_607,In_2314);
or U2221 (N_2221,In_1554,In_2080);
nand U2222 (N_2222,In_708,In_855);
nand U2223 (N_2223,In_79,In_2810);
and U2224 (N_2224,In_116,In_2860);
nand U2225 (N_2225,In_2083,In_93);
and U2226 (N_2226,In_2480,In_1140);
and U2227 (N_2227,In_1394,In_1047);
xnor U2228 (N_2228,In_2869,In_186);
nor U2229 (N_2229,In_779,In_2139);
nor U2230 (N_2230,In_1549,In_982);
nor U2231 (N_2231,In_2538,In_2714);
nor U2232 (N_2232,In_1840,In_2609);
nor U2233 (N_2233,In_20,In_1215);
nand U2234 (N_2234,In_1045,In_438);
xnor U2235 (N_2235,In_2029,In_1817);
or U2236 (N_2236,In_1508,In_1480);
nor U2237 (N_2237,In_1946,In_190);
and U2238 (N_2238,In_2744,In_1601);
nand U2239 (N_2239,In_1100,In_2839);
nor U2240 (N_2240,In_2350,In_108);
nand U2241 (N_2241,In_1456,In_96);
xor U2242 (N_2242,In_1085,In_337);
nand U2243 (N_2243,In_517,In_2302);
nand U2244 (N_2244,In_1915,In_303);
and U2245 (N_2245,In_1134,In_1378);
and U2246 (N_2246,In_2271,In_2990);
and U2247 (N_2247,In_890,In_1646);
xnor U2248 (N_2248,In_778,In_1869);
nor U2249 (N_2249,In_104,In_1243);
or U2250 (N_2250,In_1262,In_2728);
or U2251 (N_2251,In_1083,In_693);
xnor U2252 (N_2252,In_1549,In_1822);
nand U2253 (N_2253,In_1682,In_1753);
nand U2254 (N_2254,In_2531,In_408);
nand U2255 (N_2255,In_304,In_1094);
nor U2256 (N_2256,In_2560,In_2820);
nand U2257 (N_2257,In_890,In_1335);
nor U2258 (N_2258,In_612,In_291);
nand U2259 (N_2259,In_591,In_911);
and U2260 (N_2260,In_2674,In_1766);
or U2261 (N_2261,In_2105,In_451);
nand U2262 (N_2262,In_1305,In_1285);
or U2263 (N_2263,In_2099,In_204);
nor U2264 (N_2264,In_651,In_2125);
xor U2265 (N_2265,In_509,In_1510);
xor U2266 (N_2266,In_1041,In_869);
nor U2267 (N_2267,In_2457,In_541);
and U2268 (N_2268,In_1586,In_2858);
nand U2269 (N_2269,In_1668,In_950);
nand U2270 (N_2270,In_1243,In_1254);
or U2271 (N_2271,In_610,In_754);
or U2272 (N_2272,In_2814,In_2733);
or U2273 (N_2273,In_1830,In_1459);
or U2274 (N_2274,In_2640,In_2277);
and U2275 (N_2275,In_1780,In_2001);
xnor U2276 (N_2276,In_2507,In_1410);
or U2277 (N_2277,In_2081,In_472);
and U2278 (N_2278,In_2249,In_2069);
and U2279 (N_2279,In_1964,In_2151);
or U2280 (N_2280,In_2864,In_578);
or U2281 (N_2281,In_676,In_2272);
nor U2282 (N_2282,In_741,In_831);
nor U2283 (N_2283,In_2840,In_1567);
nor U2284 (N_2284,In_389,In_1136);
and U2285 (N_2285,In_553,In_2640);
nand U2286 (N_2286,In_120,In_1968);
nor U2287 (N_2287,In_1908,In_2329);
nand U2288 (N_2288,In_347,In_581);
and U2289 (N_2289,In_581,In_1903);
xnor U2290 (N_2290,In_517,In_791);
nor U2291 (N_2291,In_793,In_1505);
nand U2292 (N_2292,In_2982,In_278);
nor U2293 (N_2293,In_2986,In_1926);
nor U2294 (N_2294,In_1999,In_516);
nor U2295 (N_2295,In_2474,In_1007);
or U2296 (N_2296,In_2942,In_422);
or U2297 (N_2297,In_2021,In_1715);
nand U2298 (N_2298,In_2656,In_1);
xor U2299 (N_2299,In_2937,In_894);
nor U2300 (N_2300,In_1712,In_2221);
and U2301 (N_2301,In_773,In_2289);
or U2302 (N_2302,In_604,In_1459);
and U2303 (N_2303,In_1755,In_148);
nand U2304 (N_2304,In_369,In_1408);
xnor U2305 (N_2305,In_372,In_2071);
nor U2306 (N_2306,In_1719,In_265);
and U2307 (N_2307,In_1005,In_877);
nand U2308 (N_2308,In_590,In_514);
or U2309 (N_2309,In_995,In_2132);
nor U2310 (N_2310,In_1049,In_1955);
xnor U2311 (N_2311,In_2977,In_780);
and U2312 (N_2312,In_2740,In_2620);
xor U2313 (N_2313,In_2974,In_478);
nor U2314 (N_2314,In_496,In_2063);
xor U2315 (N_2315,In_1858,In_1393);
nand U2316 (N_2316,In_932,In_818);
nand U2317 (N_2317,In_2421,In_1173);
nor U2318 (N_2318,In_1534,In_1808);
xnor U2319 (N_2319,In_53,In_671);
or U2320 (N_2320,In_2728,In_1786);
nor U2321 (N_2321,In_2947,In_2613);
and U2322 (N_2322,In_2702,In_1261);
nand U2323 (N_2323,In_2325,In_1787);
and U2324 (N_2324,In_441,In_2194);
nor U2325 (N_2325,In_1486,In_2806);
nand U2326 (N_2326,In_1395,In_1929);
and U2327 (N_2327,In_2376,In_190);
xor U2328 (N_2328,In_1518,In_1547);
nand U2329 (N_2329,In_1994,In_1872);
nor U2330 (N_2330,In_1765,In_688);
or U2331 (N_2331,In_39,In_750);
nor U2332 (N_2332,In_60,In_835);
nand U2333 (N_2333,In_1565,In_405);
nor U2334 (N_2334,In_2868,In_174);
nand U2335 (N_2335,In_2667,In_2509);
nor U2336 (N_2336,In_979,In_431);
nor U2337 (N_2337,In_795,In_2093);
and U2338 (N_2338,In_490,In_922);
or U2339 (N_2339,In_1422,In_1111);
xnor U2340 (N_2340,In_495,In_2163);
xnor U2341 (N_2341,In_1854,In_382);
or U2342 (N_2342,In_2605,In_698);
and U2343 (N_2343,In_2409,In_585);
and U2344 (N_2344,In_1535,In_2097);
and U2345 (N_2345,In_2112,In_2581);
xor U2346 (N_2346,In_1664,In_2272);
nor U2347 (N_2347,In_2777,In_2011);
xnor U2348 (N_2348,In_1607,In_1943);
nor U2349 (N_2349,In_2952,In_108);
nand U2350 (N_2350,In_1579,In_488);
or U2351 (N_2351,In_512,In_212);
xor U2352 (N_2352,In_2389,In_885);
nand U2353 (N_2353,In_2635,In_1893);
nor U2354 (N_2354,In_1924,In_2783);
xnor U2355 (N_2355,In_25,In_1731);
nand U2356 (N_2356,In_86,In_2040);
xnor U2357 (N_2357,In_889,In_238);
nor U2358 (N_2358,In_1240,In_1849);
xnor U2359 (N_2359,In_2540,In_2709);
xor U2360 (N_2360,In_918,In_732);
and U2361 (N_2361,In_846,In_1443);
and U2362 (N_2362,In_1339,In_157);
nor U2363 (N_2363,In_2552,In_1330);
and U2364 (N_2364,In_1325,In_1126);
xor U2365 (N_2365,In_310,In_2181);
and U2366 (N_2366,In_153,In_492);
xnor U2367 (N_2367,In_1833,In_2774);
nand U2368 (N_2368,In_1054,In_642);
xnor U2369 (N_2369,In_857,In_1015);
and U2370 (N_2370,In_186,In_84);
and U2371 (N_2371,In_2764,In_6);
nor U2372 (N_2372,In_1016,In_1613);
nor U2373 (N_2373,In_529,In_1415);
or U2374 (N_2374,In_1073,In_2057);
nand U2375 (N_2375,In_1062,In_588);
nand U2376 (N_2376,In_2296,In_2630);
and U2377 (N_2377,In_2987,In_1235);
nor U2378 (N_2378,In_2098,In_2261);
and U2379 (N_2379,In_1021,In_2012);
and U2380 (N_2380,In_1908,In_712);
or U2381 (N_2381,In_1296,In_1683);
xor U2382 (N_2382,In_2491,In_1797);
or U2383 (N_2383,In_2721,In_1571);
nand U2384 (N_2384,In_2020,In_1177);
and U2385 (N_2385,In_328,In_1304);
nor U2386 (N_2386,In_1718,In_2703);
xnor U2387 (N_2387,In_2421,In_1547);
nor U2388 (N_2388,In_2380,In_746);
nor U2389 (N_2389,In_1416,In_2624);
and U2390 (N_2390,In_1611,In_1025);
xor U2391 (N_2391,In_1302,In_400);
and U2392 (N_2392,In_284,In_2501);
or U2393 (N_2393,In_1873,In_2794);
nand U2394 (N_2394,In_2009,In_2339);
or U2395 (N_2395,In_1858,In_2109);
and U2396 (N_2396,In_1984,In_2394);
xor U2397 (N_2397,In_2130,In_1401);
nor U2398 (N_2398,In_1459,In_1007);
or U2399 (N_2399,In_2840,In_1729);
and U2400 (N_2400,In_176,In_2463);
nor U2401 (N_2401,In_1754,In_2883);
nor U2402 (N_2402,In_951,In_319);
or U2403 (N_2403,In_751,In_620);
xor U2404 (N_2404,In_427,In_22);
or U2405 (N_2405,In_2457,In_1958);
and U2406 (N_2406,In_493,In_324);
nand U2407 (N_2407,In_306,In_2707);
or U2408 (N_2408,In_1161,In_2582);
or U2409 (N_2409,In_942,In_1721);
or U2410 (N_2410,In_579,In_2881);
nand U2411 (N_2411,In_1578,In_900);
or U2412 (N_2412,In_707,In_2876);
and U2413 (N_2413,In_1799,In_1582);
nor U2414 (N_2414,In_948,In_519);
nand U2415 (N_2415,In_515,In_2619);
nand U2416 (N_2416,In_2182,In_2169);
and U2417 (N_2417,In_2351,In_809);
nor U2418 (N_2418,In_128,In_2408);
or U2419 (N_2419,In_1436,In_721);
xor U2420 (N_2420,In_2008,In_1516);
nand U2421 (N_2421,In_2640,In_438);
nand U2422 (N_2422,In_2469,In_1436);
xnor U2423 (N_2423,In_2407,In_2073);
xnor U2424 (N_2424,In_722,In_627);
nor U2425 (N_2425,In_1655,In_191);
and U2426 (N_2426,In_2064,In_2893);
and U2427 (N_2427,In_499,In_2329);
nand U2428 (N_2428,In_1373,In_788);
and U2429 (N_2429,In_1275,In_2090);
or U2430 (N_2430,In_390,In_2733);
xor U2431 (N_2431,In_530,In_1559);
and U2432 (N_2432,In_48,In_2349);
xor U2433 (N_2433,In_152,In_1534);
nand U2434 (N_2434,In_2028,In_2596);
nand U2435 (N_2435,In_511,In_1866);
nand U2436 (N_2436,In_2822,In_1225);
and U2437 (N_2437,In_1234,In_2470);
or U2438 (N_2438,In_2423,In_1691);
and U2439 (N_2439,In_1480,In_2282);
xnor U2440 (N_2440,In_2558,In_1649);
or U2441 (N_2441,In_23,In_251);
and U2442 (N_2442,In_2843,In_507);
and U2443 (N_2443,In_1316,In_1404);
and U2444 (N_2444,In_2862,In_89);
nand U2445 (N_2445,In_1252,In_2046);
nand U2446 (N_2446,In_1884,In_1836);
nor U2447 (N_2447,In_1943,In_892);
nor U2448 (N_2448,In_107,In_1134);
and U2449 (N_2449,In_2751,In_1695);
and U2450 (N_2450,In_1673,In_341);
nand U2451 (N_2451,In_2298,In_645);
nand U2452 (N_2452,In_629,In_2660);
and U2453 (N_2453,In_1362,In_1767);
and U2454 (N_2454,In_2429,In_2727);
xor U2455 (N_2455,In_1750,In_1728);
nand U2456 (N_2456,In_1824,In_2270);
nor U2457 (N_2457,In_1793,In_1000);
and U2458 (N_2458,In_2052,In_1904);
nor U2459 (N_2459,In_706,In_1593);
nor U2460 (N_2460,In_959,In_2150);
nand U2461 (N_2461,In_1655,In_196);
and U2462 (N_2462,In_1897,In_1971);
nor U2463 (N_2463,In_200,In_1918);
xor U2464 (N_2464,In_1851,In_2574);
or U2465 (N_2465,In_1656,In_503);
nor U2466 (N_2466,In_186,In_1369);
xor U2467 (N_2467,In_226,In_2128);
nor U2468 (N_2468,In_2667,In_182);
or U2469 (N_2469,In_1157,In_1308);
and U2470 (N_2470,In_1655,In_1454);
or U2471 (N_2471,In_2773,In_419);
and U2472 (N_2472,In_633,In_2797);
and U2473 (N_2473,In_122,In_2309);
and U2474 (N_2474,In_1395,In_358);
or U2475 (N_2475,In_940,In_2683);
and U2476 (N_2476,In_1161,In_1872);
nand U2477 (N_2477,In_1470,In_2915);
or U2478 (N_2478,In_1552,In_1897);
xor U2479 (N_2479,In_1908,In_1162);
nor U2480 (N_2480,In_2022,In_236);
nor U2481 (N_2481,In_1764,In_1476);
and U2482 (N_2482,In_780,In_1324);
nor U2483 (N_2483,In_85,In_2897);
and U2484 (N_2484,In_49,In_1805);
nor U2485 (N_2485,In_2397,In_282);
nor U2486 (N_2486,In_2505,In_2697);
xnor U2487 (N_2487,In_2256,In_2050);
nand U2488 (N_2488,In_1293,In_49);
xnor U2489 (N_2489,In_2413,In_2951);
or U2490 (N_2490,In_740,In_343);
xor U2491 (N_2491,In_2467,In_2361);
nor U2492 (N_2492,In_1786,In_1891);
and U2493 (N_2493,In_1951,In_2289);
nor U2494 (N_2494,In_593,In_18);
nand U2495 (N_2495,In_634,In_138);
xor U2496 (N_2496,In_446,In_1301);
nand U2497 (N_2497,In_1707,In_1537);
nor U2498 (N_2498,In_1701,In_1827);
and U2499 (N_2499,In_1459,In_1329);
or U2500 (N_2500,In_2596,In_1604);
nand U2501 (N_2501,In_13,In_1864);
nand U2502 (N_2502,In_393,In_1854);
nor U2503 (N_2503,In_257,In_1989);
nand U2504 (N_2504,In_1492,In_1833);
and U2505 (N_2505,In_2451,In_1171);
and U2506 (N_2506,In_1575,In_429);
nand U2507 (N_2507,In_2049,In_1948);
nor U2508 (N_2508,In_2990,In_1537);
nand U2509 (N_2509,In_2039,In_1201);
or U2510 (N_2510,In_1554,In_963);
nor U2511 (N_2511,In_1861,In_656);
xnor U2512 (N_2512,In_1202,In_2100);
xor U2513 (N_2513,In_2584,In_1478);
and U2514 (N_2514,In_1512,In_161);
or U2515 (N_2515,In_1441,In_751);
or U2516 (N_2516,In_322,In_230);
nor U2517 (N_2517,In_785,In_1026);
xnor U2518 (N_2518,In_2802,In_309);
and U2519 (N_2519,In_207,In_1331);
or U2520 (N_2520,In_2794,In_153);
nor U2521 (N_2521,In_887,In_1503);
and U2522 (N_2522,In_1188,In_617);
xor U2523 (N_2523,In_2242,In_1953);
nand U2524 (N_2524,In_1306,In_1189);
nand U2525 (N_2525,In_2874,In_448);
nand U2526 (N_2526,In_1530,In_1273);
and U2527 (N_2527,In_2271,In_1022);
and U2528 (N_2528,In_1575,In_2821);
xnor U2529 (N_2529,In_1280,In_552);
nand U2530 (N_2530,In_1340,In_2324);
nand U2531 (N_2531,In_1000,In_412);
nand U2532 (N_2532,In_1002,In_2673);
and U2533 (N_2533,In_681,In_1499);
xor U2534 (N_2534,In_1747,In_1801);
nand U2535 (N_2535,In_597,In_719);
xnor U2536 (N_2536,In_646,In_2715);
xnor U2537 (N_2537,In_1921,In_2897);
xnor U2538 (N_2538,In_2850,In_1092);
and U2539 (N_2539,In_1083,In_1027);
nor U2540 (N_2540,In_399,In_2935);
or U2541 (N_2541,In_2328,In_2322);
and U2542 (N_2542,In_544,In_1035);
and U2543 (N_2543,In_623,In_1287);
or U2544 (N_2544,In_1578,In_2521);
xor U2545 (N_2545,In_391,In_607);
or U2546 (N_2546,In_956,In_2068);
nor U2547 (N_2547,In_33,In_1872);
nor U2548 (N_2548,In_2630,In_2996);
nand U2549 (N_2549,In_2589,In_2918);
or U2550 (N_2550,In_2232,In_1923);
xnor U2551 (N_2551,In_633,In_483);
xor U2552 (N_2552,In_2583,In_780);
xnor U2553 (N_2553,In_125,In_1780);
or U2554 (N_2554,In_2729,In_1965);
xnor U2555 (N_2555,In_1568,In_546);
or U2556 (N_2556,In_1667,In_2161);
xor U2557 (N_2557,In_631,In_422);
nor U2558 (N_2558,In_2732,In_2956);
nor U2559 (N_2559,In_2743,In_1660);
xor U2560 (N_2560,In_2292,In_513);
nand U2561 (N_2561,In_740,In_1949);
and U2562 (N_2562,In_1877,In_2888);
or U2563 (N_2563,In_2067,In_1216);
xnor U2564 (N_2564,In_961,In_1969);
or U2565 (N_2565,In_1522,In_1067);
nand U2566 (N_2566,In_393,In_761);
nand U2567 (N_2567,In_332,In_1620);
and U2568 (N_2568,In_47,In_1526);
xor U2569 (N_2569,In_2404,In_940);
and U2570 (N_2570,In_2029,In_345);
and U2571 (N_2571,In_1617,In_2764);
or U2572 (N_2572,In_1910,In_761);
nand U2573 (N_2573,In_26,In_1692);
or U2574 (N_2574,In_1082,In_1563);
xnor U2575 (N_2575,In_1799,In_354);
xor U2576 (N_2576,In_2402,In_1823);
xnor U2577 (N_2577,In_876,In_1894);
nand U2578 (N_2578,In_266,In_125);
or U2579 (N_2579,In_1519,In_2534);
or U2580 (N_2580,In_1160,In_2607);
xnor U2581 (N_2581,In_2902,In_424);
nand U2582 (N_2582,In_1808,In_585);
nand U2583 (N_2583,In_1344,In_2457);
or U2584 (N_2584,In_2159,In_1207);
or U2585 (N_2585,In_2022,In_339);
xnor U2586 (N_2586,In_2270,In_1257);
xnor U2587 (N_2587,In_2601,In_783);
or U2588 (N_2588,In_2904,In_2485);
xnor U2589 (N_2589,In_1049,In_1820);
nand U2590 (N_2590,In_1759,In_1602);
and U2591 (N_2591,In_431,In_1737);
nand U2592 (N_2592,In_2039,In_1152);
and U2593 (N_2593,In_1063,In_2556);
or U2594 (N_2594,In_963,In_2806);
or U2595 (N_2595,In_1528,In_1905);
and U2596 (N_2596,In_212,In_1808);
nand U2597 (N_2597,In_637,In_1728);
and U2598 (N_2598,In_1146,In_2752);
or U2599 (N_2599,In_629,In_647);
xnor U2600 (N_2600,In_88,In_2586);
or U2601 (N_2601,In_412,In_2675);
nor U2602 (N_2602,In_1217,In_1309);
or U2603 (N_2603,In_1007,In_908);
xnor U2604 (N_2604,In_30,In_1451);
and U2605 (N_2605,In_101,In_2089);
nand U2606 (N_2606,In_181,In_2867);
nor U2607 (N_2607,In_1984,In_1720);
nand U2608 (N_2608,In_1493,In_282);
or U2609 (N_2609,In_1624,In_2546);
nor U2610 (N_2610,In_730,In_2672);
or U2611 (N_2611,In_2520,In_395);
xnor U2612 (N_2612,In_2390,In_2745);
xor U2613 (N_2613,In_475,In_2502);
nand U2614 (N_2614,In_44,In_1945);
nor U2615 (N_2615,In_263,In_2382);
xor U2616 (N_2616,In_2883,In_529);
nor U2617 (N_2617,In_641,In_1833);
nor U2618 (N_2618,In_1925,In_1825);
nand U2619 (N_2619,In_2549,In_2328);
nand U2620 (N_2620,In_2093,In_2136);
xnor U2621 (N_2621,In_706,In_788);
nor U2622 (N_2622,In_1502,In_2535);
nor U2623 (N_2623,In_2509,In_2315);
or U2624 (N_2624,In_2289,In_319);
nand U2625 (N_2625,In_1849,In_405);
and U2626 (N_2626,In_308,In_1478);
nor U2627 (N_2627,In_2134,In_2718);
nand U2628 (N_2628,In_2008,In_2994);
nor U2629 (N_2629,In_439,In_1522);
nand U2630 (N_2630,In_2594,In_1831);
xnor U2631 (N_2631,In_158,In_1977);
nor U2632 (N_2632,In_1050,In_1798);
or U2633 (N_2633,In_922,In_2961);
or U2634 (N_2634,In_2912,In_1754);
and U2635 (N_2635,In_1573,In_300);
or U2636 (N_2636,In_2984,In_2268);
xor U2637 (N_2637,In_197,In_365);
and U2638 (N_2638,In_2631,In_1640);
nor U2639 (N_2639,In_1104,In_1847);
or U2640 (N_2640,In_864,In_1492);
or U2641 (N_2641,In_1591,In_1579);
or U2642 (N_2642,In_1635,In_2733);
nor U2643 (N_2643,In_195,In_2746);
or U2644 (N_2644,In_393,In_368);
xor U2645 (N_2645,In_1038,In_2056);
xor U2646 (N_2646,In_261,In_488);
or U2647 (N_2647,In_617,In_76);
or U2648 (N_2648,In_695,In_618);
and U2649 (N_2649,In_2589,In_2167);
or U2650 (N_2650,In_120,In_2025);
and U2651 (N_2651,In_694,In_2856);
or U2652 (N_2652,In_1645,In_1956);
or U2653 (N_2653,In_2510,In_2753);
and U2654 (N_2654,In_1616,In_1288);
or U2655 (N_2655,In_1996,In_1825);
xor U2656 (N_2656,In_1230,In_2682);
nor U2657 (N_2657,In_46,In_2136);
or U2658 (N_2658,In_442,In_1576);
and U2659 (N_2659,In_1249,In_1200);
or U2660 (N_2660,In_2111,In_715);
nor U2661 (N_2661,In_943,In_2658);
nor U2662 (N_2662,In_2170,In_2753);
nand U2663 (N_2663,In_2725,In_774);
and U2664 (N_2664,In_2087,In_1904);
and U2665 (N_2665,In_968,In_2941);
or U2666 (N_2666,In_1108,In_690);
nand U2667 (N_2667,In_1172,In_106);
xor U2668 (N_2668,In_2166,In_2322);
and U2669 (N_2669,In_1277,In_1901);
xnor U2670 (N_2670,In_2992,In_1349);
xor U2671 (N_2671,In_440,In_723);
or U2672 (N_2672,In_258,In_2585);
and U2673 (N_2673,In_519,In_1388);
and U2674 (N_2674,In_73,In_339);
xnor U2675 (N_2675,In_385,In_1931);
nor U2676 (N_2676,In_632,In_2002);
xnor U2677 (N_2677,In_1010,In_337);
nand U2678 (N_2678,In_1589,In_514);
xnor U2679 (N_2679,In_1206,In_134);
nor U2680 (N_2680,In_581,In_1986);
nand U2681 (N_2681,In_2327,In_618);
and U2682 (N_2682,In_2746,In_2336);
xor U2683 (N_2683,In_2663,In_720);
nor U2684 (N_2684,In_1483,In_2712);
nand U2685 (N_2685,In_1226,In_1436);
and U2686 (N_2686,In_618,In_2508);
nor U2687 (N_2687,In_1177,In_155);
and U2688 (N_2688,In_1720,In_2706);
or U2689 (N_2689,In_2746,In_221);
or U2690 (N_2690,In_2329,In_2815);
xor U2691 (N_2691,In_1953,In_405);
xor U2692 (N_2692,In_382,In_1436);
nand U2693 (N_2693,In_51,In_1863);
and U2694 (N_2694,In_5,In_665);
nor U2695 (N_2695,In_419,In_367);
nand U2696 (N_2696,In_1310,In_316);
and U2697 (N_2697,In_1951,In_1523);
or U2698 (N_2698,In_900,In_1691);
or U2699 (N_2699,In_493,In_2223);
or U2700 (N_2700,In_2225,In_387);
xnor U2701 (N_2701,In_2643,In_1126);
and U2702 (N_2702,In_943,In_1729);
or U2703 (N_2703,In_1116,In_521);
or U2704 (N_2704,In_1795,In_2006);
and U2705 (N_2705,In_160,In_2830);
and U2706 (N_2706,In_1659,In_589);
and U2707 (N_2707,In_153,In_2246);
xnor U2708 (N_2708,In_2862,In_2608);
nand U2709 (N_2709,In_1467,In_377);
xnor U2710 (N_2710,In_109,In_1220);
nor U2711 (N_2711,In_1093,In_2475);
xnor U2712 (N_2712,In_692,In_1521);
or U2713 (N_2713,In_2970,In_1864);
nor U2714 (N_2714,In_2217,In_860);
xnor U2715 (N_2715,In_749,In_2030);
xor U2716 (N_2716,In_2856,In_2738);
nor U2717 (N_2717,In_2971,In_68);
or U2718 (N_2718,In_1529,In_1536);
nand U2719 (N_2719,In_1228,In_2349);
nand U2720 (N_2720,In_2803,In_1440);
xnor U2721 (N_2721,In_1127,In_1223);
and U2722 (N_2722,In_1718,In_1074);
xnor U2723 (N_2723,In_206,In_262);
and U2724 (N_2724,In_2149,In_2683);
and U2725 (N_2725,In_385,In_1002);
nor U2726 (N_2726,In_507,In_2892);
nor U2727 (N_2727,In_972,In_2812);
nor U2728 (N_2728,In_1718,In_2140);
or U2729 (N_2729,In_1022,In_2519);
and U2730 (N_2730,In_1456,In_1233);
xnor U2731 (N_2731,In_2985,In_482);
nor U2732 (N_2732,In_2653,In_2165);
and U2733 (N_2733,In_156,In_1970);
or U2734 (N_2734,In_1013,In_2157);
xnor U2735 (N_2735,In_2790,In_2519);
xnor U2736 (N_2736,In_1993,In_414);
or U2737 (N_2737,In_281,In_1951);
and U2738 (N_2738,In_925,In_1367);
nor U2739 (N_2739,In_935,In_514);
nand U2740 (N_2740,In_1524,In_2581);
and U2741 (N_2741,In_534,In_1227);
and U2742 (N_2742,In_2300,In_2011);
and U2743 (N_2743,In_2167,In_965);
and U2744 (N_2744,In_1137,In_2941);
or U2745 (N_2745,In_2006,In_2835);
xnor U2746 (N_2746,In_1442,In_2587);
and U2747 (N_2747,In_2070,In_546);
nor U2748 (N_2748,In_203,In_2876);
nand U2749 (N_2749,In_326,In_2961);
nand U2750 (N_2750,In_2496,In_1571);
nand U2751 (N_2751,In_1353,In_1819);
and U2752 (N_2752,In_2571,In_949);
or U2753 (N_2753,In_2255,In_1374);
nand U2754 (N_2754,In_2257,In_231);
xnor U2755 (N_2755,In_2248,In_2994);
nor U2756 (N_2756,In_2021,In_2115);
nor U2757 (N_2757,In_2345,In_1947);
nor U2758 (N_2758,In_2580,In_690);
and U2759 (N_2759,In_785,In_156);
or U2760 (N_2760,In_2408,In_818);
xor U2761 (N_2761,In_620,In_2398);
xnor U2762 (N_2762,In_1698,In_2964);
and U2763 (N_2763,In_1116,In_1390);
or U2764 (N_2764,In_2706,In_1918);
and U2765 (N_2765,In_2268,In_135);
and U2766 (N_2766,In_2567,In_103);
and U2767 (N_2767,In_2485,In_546);
nor U2768 (N_2768,In_241,In_2675);
or U2769 (N_2769,In_2737,In_1689);
nand U2770 (N_2770,In_180,In_59);
or U2771 (N_2771,In_616,In_1943);
and U2772 (N_2772,In_202,In_1094);
nand U2773 (N_2773,In_1230,In_2807);
nor U2774 (N_2774,In_772,In_2839);
nor U2775 (N_2775,In_2209,In_612);
or U2776 (N_2776,In_83,In_110);
xnor U2777 (N_2777,In_2394,In_1172);
nor U2778 (N_2778,In_2128,In_438);
nor U2779 (N_2779,In_574,In_312);
xnor U2780 (N_2780,In_961,In_307);
and U2781 (N_2781,In_48,In_122);
nand U2782 (N_2782,In_155,In_2300);
nand U2783 (N_2783,In_235,In_2699);
nand U2784 (N_2784,In_1303,In_1363);
xnor U2785 (N_2785,In_2875,In_1740);
xnor U2786 (N_2786,In_291,In_2003);
nor U2787 (N_2787,In_1480,In_733);
or U2788 (N_2788,In_2877,In_1962);
xor U2789 (N_2789,In_680,In_243);
nor U2790 (N_2790,In_2049,In_2112);
nand U2791 (N_2791,In_862,In_424);
nand U2792 (N_2792,In_2195,In_911);
nand U2793 (N_2793,In_857,In_2883);
or U2794 (N_2794,In_2025,In_675);
and U2795 (N_2795,In_1218,In_2158);
nor U2796 (N_2796,In_413,In_2663);
or U2797 (N_2797,In_624,In_404);
and U2798 (N_2798,In_1075,In_702);
xnor U2799 (N_2799,In_21,In_1260);
nand U2800 (N_2800,In_2,In_1210);
or U2801 (N_2801,In_2199,In_1845);
xnor U2802 (N_2802,In_2501,In_2372);
nor U2803 (N_2803,In_2577,In_488);
and U2804 (N_2804,In_561,In_230);
nor U2805 (N_2805,In_1253,In_1401);
or U2806 (N_2806,In_527,In_919);
nand U2807 (N_2807,In_2919,In_2475);
or U2808 (N_2808,In_2025,In_698);
and U2809 (N_2809,In_1473,In_1424);
and U2810 (N_2810,In_2847,In_808);
xor U2811 (N_2811,In_1328,In_815);
and U2812 (N_2812,In_391,In_667);
or U2813 (N_2813,In_1574,In_1967);
nor U2814 (N_2814,In_1963,In_2681);
and U2815 (N_2815,In_1489,In_2633);
nand U2816 (N_2816,In_2647,In_2807);
xnor U2817 (N_2817,In_1028,In_1086);
and U2818 (N_2818,In_2220,In_1327);
and U2819 (N_2819,In_1243,In_718);
nor U2820 (N_2820,In_1102,In_165);
xnor U2821 (N_2821,In_2736,In_1288);
nor U2822 (N_2822,In_1924,In_1185);
or U2823 (N_2823,In_574,In_1851);
nor U2824 (N_2824,In_606,In_270);
and U2825 (N_2825,In_1980,In_2003);
and U2826 (N_2826,In_1207,In_829);
nor U2827 (N_2827,In_417,In_1714);
xnor U2828 (N_2828,In_746,In_1388);
nand U2829 (N_2829,In_1992,In_1236);
nor U2830 (N_2830,In_2126,In_2380);
and U2831 (N_2831,In_1922,In_2065);
xnor U2832 (N_2832,In_2609,In_2366);
xor U2833 (N_2833,In_2723,In_710);
and U2834 (N_2834,In_2797,In_308);
xnor U2835 (N_2835,In_1842,In_752);
or U2836 (N_2836,In_579,In_417);
nor U2837 (N_2837,In_1711,In_2192);
or U2838 (N_2838,In_531,In_1559);
nor U2839 (N_2839,In_2448,In_716);
nand U2840 (N_2840,In_1240,In_111);
or U2841 (N_2841,In_1558,In_1152);
xor U2842 (N_2842,In_2077,In_1312);
and U2843 (N_2843,In_348,In_2786);
xor U2844 (N_2844,In_2576,In_1991);
and U2845 (N_2845,In_2,In_1763);
nand U2846 (N_2846,In_2036,In_858);
and U2847 (N_2847,In_2654,In_1380);
xor U2848 (N_2848,In_2414,In_2535);
nor U2849 (N_2849,In_1273,In_2541);
and U2850 (N_2850,In_1723,In_149);
xnor U2851 (N_2851,In_2799,In_458);
and U2852 (N_2852,In_2814,In_988);
nand U2853 (N_2853,In_2988,In_692);
nor U2854 (N_2854,In_1128,In_2261);
xor U2855 (N_2855,In_650,In_300);
or U2856 (N_2856,In_308,In_2653);
or U2857 (N_2857,In_2919,In_1466);
nor U2858 (N_2858,In_2509,In_46);
or U2859 (N_2859,In_345,In_2436);
nor U2860 (N_2860,In_2185,In_2546);
or U2861 (N_2861,In_2366,In_38);
nor U2862 (N_2862,In_2949,In_1755);
and U2863 (N_2863,In_1093,In_2582);
xnor U2864 (N_2864,In_938,In_2536);
or U2865 (N_2865,In_2021,In_2788);
and U2866 (N_2866,In_2473,In_1325);
and U2867 (N_2867,In_2128,In_2389);
nor U2868 (N_2868,In_66,In_302);
xnor U2869 (N_2869,In_30,In_2818);
nor U2870 (N_2870,In_104,In_1551);
xor U2871 (N_2871,In_1667,In_2759);
and U2872 (N_2872,In_856,In_2585);
and U2873 (N_2873,In_2697,In_2747);
or U2874 (N_2874,In_134,In_2949);
xnor U2875 (N_2875,In_2191,In_802);
or U2876 (N_2876,In_2546,In_165);
nor U2877 (N_2877,In_618,In_1591);
and U2878 (N_2878,In_1946,In_327);
nor U2879 (N_2879,In_1706,In_451);
and U2880 (N_2880,In_948,In_1992);
nand U2881 (N_2881,In_575,In_2704);
and U2882 (N_2882,In_2878,In_2909);
and U2883 (N_2883,In_2614,In_1136);
nor U2884 (N_2884,In_2916,In_2099);
nand U2885 (N_2885,In_1241,In_224);
and U2886 (N_2886,In_2798,In_1870);
or U2887 (N_2887,In_2964,In_1083);
nand U2888 (N_2888,In_2423,In_836);
xnor U2889 (N_2889,In_2947,In_2004);
nand U2890 (N_2890,In_944,In_2572);
nor U2891 (N_2891,In_554,In_778);
nand U2892 (N_2892,In_2630,In_770);
nor U2893 (N_2893,In_1692,In_1134);
nand U2894 (N_2894,In_2783,In_858);
nor U2895 (N_2895,In_2117,In_559);
or U2896 (N_2896,In_2728,In_1275);
nand U2897 (N_2897,In_2937,In_2864);
xnor U2898 (N_2898,In_151,In_2146);
xnor U2899 (N_2899,In_308,In_852);
and U2900 (N_2900,In_2990,In_2468);
xor U2901 (N_2901,In_1226,In_962);
nand U2902 (N_2902,In_1418,In_1629);
nand U2903 (N_2903,In_10,In_820);
xor U2904 (N_2904,In_851,In_944);
nor U2905 (N_2905,In_1573,In_2365);
nand U2906 (N_2906,In_2684,In_2088);
and U2907 (N_2907,In_1776,In_782);
nand U2908 (N_2908,In_1790,In_101);
nand U2909 (N_2909,In_1879,In_2260);
nand U2910 (N_2910,In_901,In_2533);
nor U2911 (N_2911,In_983,In_2887);
xnor U2912 (N_2912,In_788,In_2570);
or U2913 (N_2913,In_135,In_2045);
and U2914 (N_2914,In_752,In_206);
xnor U2915 (N_2915,In_1678,In_2764);
xor U2916 (N_2916,In_2575,In_1602);
or U2917 (N_2917,In_2116,In_1830);
or U2918 (N_2918,In_893,In_801);
nor U2919 (N_2919,In_354,In_1562);
nand U2920 (N_2920,In_1523,In_2865);
xor U2921 (N_2921,In_1216,In_1828);
or U2922 (N_2922,In_1132,In_2009);
nor U2923 (N_2923,In_1781,In_734);
nor U2924 (N_2924,In_2043,In_2384);
and U2925 (N_2925,In_1767,In_2785);
nand U2926 (N_2926,In_1341,In_2446);
nand U2927 (N_2927,In_2495,In_2135);
nand U2928 (N_2928,In_2685,In_2768);
or U2929 (N_2929,In_1545,In_1944);
or U2930 (N_2930,In_1747,In_669);
xnor U2931 (N_2931,In_2882,In_2433);
and U2932 (N_2932,In_170,In_2785);
nor U2933 (N_2933,In_722,In_662);
nand U2934 (N_2934,In_816,In_2436);
and U2935 (N_2935,In_1376,In_109);
or U2936 (N_2936,In_2396,In_2276);
xor U2937 (N_2937,In_2618,In_1036);
and U2938 (N_2938,In_2557,In_2250);
nand U2939 (N_2939,In_2068,In_2522);
or U2940 (N_2940,In_591,In_380);
nand U2941 (N_2941,In_819,In_2198);
or U2942 (N_2942,In_2661,In_2304);
or U2943 (N_2943,In_2137,In_1347);
and U2944 (N_2944,In_772,In_281);
and U2945 (N_2945,In_974,In_705);
and U2946 (N_2946,In_676,In_1063);
or U2947 (N_2947,In_2323,In_2619);
xor U2948 (N_2948,In_1350,In_2432);
or U2949 (N_2949,In_2203,In_2109);
xnor U2950 (N_2950,In_2825,In_764);
and U2951 (N_2951,In_2173,In_2989);
nand U2952 (N_2952,In_806,In_1603);
nor U2953 (N_2953,In_1763,In_2223);
and U2954 (N_2954,In_1137,In_2808);
or U2955 (N_2955,In_2947,In_1410);
or U2956 (N_2956,In_1145,In_2912);
xnor U2957 (N_2957,In_1321,In_751);
or U2958 (N_2958,In_1231,In_222);
nand U2959 (N_2959,In_2938,In_2473);
or U2960 (N_2960,In_2617,In_2834);
xnor U2961 (N_2961,In_524,In_1252);
nand U2962 (N_2962,In_1443,In_2613);
and U2963 (N_2963,In_301,In_2678);
xor U2964 (N_2964,In_1101,In_1605);
nor U2965 (N_2965,In_2987,In_110);
xor U2966 (N_2966,In_2532,In_2801);
and U2967 (N_2967,In_839,In_727);
nand U2968 (N_2968,In_985,In_996);
nand U2969 (N_2969,In_2006,In_929);
nand U2970 (N_2970,In_2715,In_2890);
xor U2971 (N_2971,In_2848,In_750);
nor U2972 (N_2972,In_828,In_2143);
or U2973 (N_2973,In_1739,In_2567);
xor U2974 (N_2974,In_1650,In_207);
or U2975 (N_2975,In_861,In_2864);
or U2976 (N_2976,In_377,In_2134);
and U2977 (N_2977,In_1302,In_1547);
nor U2978 (N_2978,In_832,In_1929);
nor U2979 (N_2979,In_276,In_2533);
or U2980 (N_2980,In_2970,In_1049);
nand U2981 (N_2981,In_2180,In_2752);
nor U2982 (N_2982,In_1615,In_1000);
nand U2983 (N_2983,In_2526,In_776);
xnor U2984 (N_2984,In_1609,In_2978);
nor U2985 (N_2985,In_1190,In_1538);
and U2986 (N_2986,In_2940,In_473);
xor U2987 (N_2987,In_2599,In_2411);
nor U2988 (N_2988,In_1784,In_1256);
xor U2989 (N_2989,In_1594,In_72);
xnor U2990 (N_2990,In_595,In_1680);
nor U2991 (N_2991,In_504,In_2782);
and U2992 (N_2992,In_548,In_929);
nor U2993 (N_2993,In_1157,In_1451);
or U2994 (N_2994,In_2093,In_1728);
xnor U2995 (N_2995,In_1893,In_1235);
or U2996 (N_2996,In_495,In_1459);
or U2997 (N_2997,In_2994,In_1958);
or U2998 (N_2998,In_2816,In_605);
nand U2999 (N_2999,In_1601,In_880);
or U3000 (N_3000,In_1733,In_1164);
nand U3001 (N_3001,In_2781,In_423);
nand U3002 (N_3002,In_1475,In_638);
nor U3003 (N_3003,In_113,In_277);
or U3004 (N_3004,In_522,In_1386);
nor U3005 (N_3005,In_591,In_1408);
xor U3006 (N_3006,In_2277,In_1766);
nand U3007 (N_3007,In_1792,In_176);
and U3008 (N_3008,In_87,In_95);
xnor U3009 (N_3009,In_659,In_2618);
and U3010 (N_3010,In_1722,In_1482);
nor U3011 (N_3011,In_1566,In_435);
xnor U3012 (N_3012,In_2576,In_2994);
or U3013 (N_3013,In_1088,In_1812);
xnor U3014 (N_3014,In_2176,In_2795);
or U3015 (N_3015,In_2308,In_362);
or U3016 (N_3016,In_0,In_737);
xor U3017 (N_3017,In_640,In_2659);
xor U3018 (N_3018,In_443,In_712);
xnor U3019 (N_3019,In_2858,In_1063);
or U3020 (N_3020,In_979,In_639);
nand U3021 (N_3021,In_1418,In_598);
xor U3022 (N_3022,In_270,In_393);
and U3023 (N_3023,In_2251,In_295);
or U3024 (N_3024,In_2729,In_937);
xnor U3025 (N_3025,In_1009,In_1347);
and U3026 (N_3026,In_2654,In_1654);
or U3027 (N_3027,In_2454,In_2432);
nand U3028 (N_3028,In_2161,In_1501);
nor U3029 (N_3029,In_2665,In_1915);
and U3030 (N_3030,In_425,In_891);
and U3031 (N_3031,In_2564,In_1301);
nor U3032 (N_3032,In_2075,In_520);
nand U3033 (N_3033,In_2156,In_50);
and U3034 (N_3034,In_2623,In_400);
nand U3035 (N_3035,In_2286,In_2145);
and U3036 (N_3036,In_1033,In_948);
xor U3037 (N_3037,In_49,In_1637);
nand U3038 (N_3038,In_720,In_1002);
nand U3039 (N_3039,In_2410,In_803);
nand U3040 (N_3040,In_859,In_255);
and U3041 (N_3041,In_2684,In_1049);
nor U3042 (N_3042,In_516,In_2419);
nor U3043 (N_3043,In_2162,In_1166);
xor U3044 (N_3044,In_297,In_2937);
nor U3045 (N_3045,In_2160,In_1002);
nor U3046 (N_3046,In_1993,In_2538);
nand U3047 (N_3047,In_1815,In_1282);
xor U3048 (N_3048,In_503,In_1454);
nor U3049 (N_3049,In_2540,In_687);
xor U3050 (N_3050,In_2301,In_2176);
or U3051 (N_3051,In_1269,In_2764);
and U3052 (N_3052,In_2311,In_1821);
or U3053 (N_3053,In_262,In_450);
nand U3054 (N_3054,In_19,In_2966);
or U3055 (N_3055,In_354,In_1807);
and U3056 (N_3056,In_1437,In_171);
and U3057 (N_3057,In_1324,In_2181);
xor U3058 (N_3058,In_1659,In_1037);
or U3059 (N_3059,In_2745,In_2213);
nand U3060 (N_3060,In_2436,In_49);
nor U3061 (N_3061,In_86,In_2590);
xor U3062 (N_3062,In_2975,In_2323);
nand U3063 (N_3063,In_2974,In_2450);
nand U3064 (N_3064,In_2585,In_1788);
nor U3065 (N_3065,In_1421,In_2494);
or U3066 (N_3066,In_2567,In_168);
nand U3067 (N_3067,In_783,In_2377);
nor U3068 (N_3068,In_2781,In_2903);
nand U3069 (N_3069,In_450,In_1427);
xor U3070 (N_3070,In_1834,In_2145);
or U3071 (N_3071,In_1991,In_1936);
nor U3072 (N_3072,In_1519,In_1638);
nand U3073 (N_3073,In_709,In_341);
and U3074 (N_3074,In_254,In_1218);
xor U3075 (N_3075,In_935,In_476);
nor U3076 (N_3076,In_338,In_1795);
nor U3077 (N_3077,In_239,In_2673);
nand U3078 (N_3078,In_775,In_1418);
nor U3079 (N_3079,In_1968,In_1789);
and U3080 (N_3080,In_671,In_2323);
xor U3081 (N_3081,In_2762,In_457);
nor U3082 (N_3082,In_880,In_2383);
nor U3083 (N_3083,In_288,In_2864);
or U3084 (N_3084,In_2377,In_2733);
or U3085 (N_3085,In_540,In_1653);
nand U3086 (N_3086,In_395,In_2719);
or U3087 (N_3087,In_1872,In_2920);
xnor U3088 (N_3088,In_1722,In_2870);
nor U3089 (N_3089,In_271,In_1563);
nand U3090 (N_3090,In_669,In_2622);
nor U3091 (N_3091,In_280,In_992);
nor U3092 (N_3092,In_184,In_1130);
or U3093 (N_3093,In_2150,In_902);
nor U3094 (N_3094,In_2323,In_268);
and U3095 (N_3095,In_1134,In_1590);
or U3096 (N_3096,In_2537,In_356);
nand U3097 (N_3097,In_2838,In_668);
nand U3098 (N_3098,In_2248,In_2923);
or U3099 (N_3099,In_938,In_332);
or U3100 (N_3100,In_1097,In_2969);
and U3101 (N_3101,In_783,In_1192);
xor U3102 (N_3102,In_542,In_1442);
nor U3103 (N_3103,In_2920,In_2222);
nand U3104 (N_3104,In_170,In_1328);
and U3105 (N_3105,In_1150,In_447);
or U3106 (N_3106,In_1897,In_265);
or U3107 (N_3107,In_1118,In_1698);
or U3108 (N_3108,In_606,In_127);
or U3109 (N_3109,In_2967,In_2566);
xor U3110 (N_3110,In_1948,In_877);
nand U3111 (N_3111,In_1861,In_2499);
xnor U3112 (N_3112,In_180,In_2251);
or U3113 (N_3113,In_1926,In_791);
or U3114 (N_3114,In_2774,In_2633);
nand U3115 (N_3115,In_267,In_1416);
nand U3116 (N_3116,In_1080,In_977);
or U3117 (N_3117,In_2275,In_592);
nand U3118 (N_3118,In_2240,In_1492);
nand U3119 (N_3119,In_1118,In_1586);
nor U3120 (N_3120,In_2406,In_2258);
nor U3121 (N_3121,In_1445,In_2925);
or U3122 (N_3122,In_1165,In_85);
or U3123 (N_3123,In_2050,In_2966);
nand U3124 (N_3124,In_174,In_2314);
or U3125 (N_3125,In_1913,In_311);
nor U3126 (N_3126,In_1324,In_2729);
xor U3127 (N_3127,In_2159,In_2678);
xor U3128 (N_3128,In_2737,In_1908);
or U3129 (N_3129,In_1111,In_2574);
or U3130 (N_3130,In_778,In_218);
nand U3131 (N_3131,In_2502,In_2222);
nor U3132 (N_3132,In_583,In_1792);
nor U3133 (N_3133,In_1731,In_9);
nand U3134 (N_3134,In_337,In_1011);
or U3135 (N_3135,In_1211,In_2616);
xor U3136 (N_3136,In_2665,In_667);
and U3137 (N_3137,In_1363,In_2313);
xnor U3138 (N_3138,In_267,In_1857);
nor U3139 (N_3139,In_814,In_130);
nand U3140 (N_3140,In_720,In_2565);
and U3141 (N_3141,In_751,In_1001);
xor U3142 (N_3142,In_2787,In_2489);
and U3143 (N_3143,In_2137,In_1922);
nor U3144 (N_3144,In_1525,In_879);
or U3145 (N_3145,In_2733,In_17);
nand U3146 (N_3146,In_1364,In_1967);
and U3147 (N_3147,In_392,In_489);
nand U3148 (N_3148,In_2079,In_2365);
and U3149 (N_3149,In_1407,In_2979);
xor U3150 (N_3150,In_1977,In_794);
nand U3151 (N_3151,In_1900,In_2743);
xnor U3152 (N_3152,In_2864,In_1892);
or U3153 (N_3153,In_1622,In_1792);
nor U3154 (N_3154,In_1332,In_1580);
nand U3155 (N_3155,In_1408,In_187);
nor U3156 (N_3156,In_805,In_2471);
or U3157 (N_3157,In_2266,In_868);
nor U3158 (N_3158,In_2281,In_916);
and U3159 (N_3159,In_937,In_1834);
nor U3160 (N_3160,In_2563,In_2765);
nand U3161 (N_3161,In_309,In_1433);
nor U3162 (N_3162,In_944,In_1433);
nor U3163 (N_3163,In_2167,In_1354);
xor U3164 (N_3164,In_2451,In_2326);
xor U3165 (N_3165,In_1726,In_751);
or U3166 (N_3166,In_1575,In_1735);
nand U3167 (N_3167,In_726,In_847);
xor U3168 (N_3168,In_2840,In_916);
nand U3169 (N_3169,In_462,In_787);
or U3170 (N_3170,In_2596,In_621);
or U3171 (N_3171,In_2152,In_595);
and U3172 (N_3172,In_1994,In_668);
and U3173 (N_3173,In_1926,In_978);
nand U3174 (N_3174,In_2540,In_249);
or U3175 (N_3175,In_1962,In_118);
or U3176 (N_3176,In_750,In_923);
nand U3177 (N_3177,In_2117,In_1024);
nor U3178 (N_3178,In_2554,In_729);
nor U3179 (N_3179,In_81,In_261);
xor U3180 (N_3180,In_2844,In_2674);
xor U3181 (N_3181,In_2796,In_1882);
or U3182 (N_3182,In_1800,In_455);
nor U3183 (N_3183,In_2749,In_716);
nor U3184 (N_3184,In_99,In_116);
and U3185 (N_3185,In_499,In_39);
and U3186 (N_3186,In_2977,In_697);
nor U3187 (N_3187,In_2038,In_2159);
nor U3188 (N_3188,In_875,In_1363);
and U3189 (N_3189,In_1569,In_1339);
or U3190 (N_3190,In_652,In_529);
and U3191 (N_3191,In_319,In_19);
xor U3192 (N_3192,In_481,In_650);
xor U3193 (N_3193,In_2920,In_140);
xor U3194 (N_3194,In_894,In_1000);
nand U3195 (N_3195,In_286,In_1440);
or U3196 (N_3196,In_125,In_2223);
xnor U3197 (N_3197,In_1970,In_2585);
nand U3198 (N_3198,In_2812,In_1840);
nand U3199 (N_3199,In_547,In_2451);
nand U3200 (N_3200,In_1562,In_1227);
xnor U3201 (N_3201,In_2367,In_296);
nor U3202 (N_3202,In_2417,In_852);
and U3203 (N_3203,In_2176,In_268);
xor U3204 (N_3204,In_800,In_1719);
nand U3205 (N_3205,In_1748,In_313);
and U3206 (N_3206,In_2081,In_1225);
xnor U3207 (N_3207,In_2041,In_2699);
xor U3208 (N_3208,In_396,In_2324);
and U3209 (N_3209,In_2455,In_1670);
nor U3210 (N_3210,In_2804,In_2901);
and U3211 (N_3211,In_1408,In_2105);
or U3212 (N_3212,In_2551,In_2708);
nor U3213 (N_3213,In_1369,In_2478);
and U3214 (N_3214,In_1807,In_173);
and U3215 (N_3215,In_2700,In_2751);
nand U3216 (N_3216,In_1829,In_1863);
nand U3217 (N_3217,In_1416,In_1494);
or U3218 (N_3218,In_1212,In_1149);
nor U3219 (N_3219,In_2893,In_1452);
and U3220 (N_3220,In_304,In_130);
nand U3221 (N_3221,In_1584,In_381);
and U3222 (N_3222,In_2750,In_1600);
or U3223 (N_3223,In_2378,In_693);
nand U3224 (N_3224,In_615,In_1999);
nand U3225 (N_3225,In_2016,In_2813);
nor U3226 (N_3226,In_2691,In_1331);
and U3227 (N_3227,In_2854,In_1652);
xor U3228 (N_3228,In_2387,In_868);
xor U3229 (N_3229,In_360,In_211);
nand U3230 (N_3230,In_2918,In_2801);
xnor U3231 (N_3231,In_1562,In_677);
nand U3232 (N_3232,In_1443,In_2194);
nor U3233 (N_3233,In_1560,In_2362);
and U3234 (N_3234,In_2191,In_1105);
xnor U3235 (N_3235,In_1354,In_2260);
xnor U3236 (N_3236,In_1327,In_332);
nor U3237 (N_3237,In_310,In_749);
xnor U3238 (N_3238,In_884,In_1290);
nand U3239 (N_3239,In_2919,In_2643);
xor U3240 (N_3240,In_1086,In_2763);
and U3241 (N_3241,In_266,In_1382);
xor U3242 (N_3242,In_1732,In_2930);
nor U3243 (N_3243,In_2179,In_386);
or U3244 (N_3244,In_155,In_1952);
nand U3245 (N_3245,In_1721,In_590);
xor U3246 (N_3246,In_732,In_2813);
or U3247 (N_3247,In_2978,In_536);
nor U3248 (N_3248,In_2311,In_1849);
nand U3249 (N_3249,In_2774,In_1850);
nand U3250 (N_3250,In_1375,In_2602);
or U3251 (N_3251,In_1644,In_1326);
nand U3252 (N_3252,In_2173,In_1494);
nand U3253 (N_3253,In_57,In_1232);
nor U3254 (N_3254,In_1676,In_1544);
nor U3255 (N_3255,In_172,In_2918);
nor U3256 (N_3256,In_2195,In_2525);
or U3257 (N_3257,In_546,In_1471);
or U3258 (N_3258,In_1625,In_2425);
nor U3259 (N_3259,In_304,In_256);
nand U3260 (N_3260,In_1098,In_2811);
xnor U3261 (N_3261,In_1154,In_2369);
or U3262 (N_3262,In_1497,In_2185);
and U3263 (N_3263,In_2755,In_801);
xor U3264 (N_3264,In_1311,In_1864);
nor U3265 (N_3265,In_1082,In_1915);
or U3266 (N_3266,In_2749,In_636);
xnor U3267 (N_3267,In_906,In_36);
or U3268 (N_3268,In_170,In_2596);
or U3269 (N_3269,In_2409,In_2492);
and U3270 (N_3270,In_2619,In_885);
xnor U3271 (N_3271,In_2305,In_2786);
nand U3272 (N_3272,In_2373,In_2042);
and U3273 (N_3273,In_2062,In_636);
xor U3274 (N_3274,In_42,In_2881);
or U3275 (N_3275,In_143,In_2624);
xnor U3276 (N_3276,In_1398,In_2668);
xor U3277 (N_3277,In_2527,In_1779);
and U3278 (N_3278,In_1453,In_2840);
nor U3279 (N_3279,In_938,In_2970);
nor U3280 (N_3280,In_1016,In_874);
nor U3281 (N_3281,In_1595,In_1157);
and U3282 (N_3282,In_2477,In_102);
nand U3283 (N_3283,In_1734,In_1559);
nor U3284 (N_3284,In_1651,In_2677);
xnor U3285 (N_3285,In_159,In_2990);
nand U3286 (N_3286,In_2050,In_1451);
xnor U3287 (N_3287,In_305,In_1680);
or U3288 (N_3288,In_2847,In_1076);
and U3289 (N_3289,In_1856,In_464);
and U3290 (N_3290,In_2707,In_1736);
or U3291 (N_3291,In_1635,In_655);
xnor U3292 (N_3292,In_1653,In_1777);
nand U3293 (N_3293,In_1215,In_2474);
nand U3294 (N_3294,In_1529,In_1936);
nand U3295 (N_3295,In_1501,In_1012);
nand U3296 (N_3296,In_736,In_1170);
nand U3297 (N_3297,In_2917,In_2337);
nand U3298 (N_3298,In_1349,In_2496);
or U3299 (N_3299,In_1218,In_2013);
or U3300 (N_3300,In_2715,In_170);
and U3301 (N_3301,In_652,In_2240);
or U3302 (N_3302,In_2797,In_2718);
xnor U3303 (N_3303,In_1112,In_194);
nor U3304 (N_3304,In_526,In_84);
or U3305 (N_3305,In_2245,In_2713);
or U3306 (N_3306,In_1545,In_2502);
or U3307 (N_3307,In_1653,In_2718);
or U3308 (N_3308,In_2773,In_890);
nor U3309 (N_3309,In_105,In_350);
or U3310 (N_3310,In_2312,In_681);
and U3311 (N_3311,In_349,In_536);
xor U3312 (N_3312,In_2549,In_302);
nand U3313 (N_3313,In_2827,In_1696);
xor U3314 (N_3314,In_1205,In_2037);
and U3315 (N_3315,In_1531,In_1663);
nand U3316 (N_3316,In_1579,In_1404);
or U3317 (N_3317,In_694,In_2434);
and U3318 (N_3318,In_1606,In_887);
or U3319 (N_3319,In_2488,In_2693);
nor U3320 (N_3320,In_2206,In_1081);
or U3321 (N_3321,In_2208,In_2986);
xnor U3322 (N_3322,In_1547,In_1027);
xor U3323 (N_3323,In_961,In_709);
nand U3324 (N_3324,In_2850,In_2515);
xor U3325 (N_3325,In_402,In_1304);
or U3326 (N_3326,In_2742,In_546);
nor U3327 (N_3327,In_2714,In_71);
nand U3328 (N_3328,In_2320,In_54);
and U3329 (N_3329,In_2981,In_2957);
xor U3330 (N_3330,In_2708,In_2902);
and U3331 (N_3331,In_2285,In_2137);
nor U3332 (N_3332,In_637,In_883);
or U3333 (N_3333,In_2302,In_2301);
nor U3334 (N_3334,In_146,In_2854);
or U3335 (N_3335,In_2139,In_825);
nand U3336 (N_3336,In_1368,In_388);
and U3337 (N_3337,In_1332,In_2927);
or U3338 (N_3338,In_617,In_2880);
xor U3339 (N_3339,In_335,In_2505);
and U3340 (N_3340,In_815,In_67);
and U3341 (N_3341,In_1561,In_2271);
and U3342 (N_3342,In_762,In_2162);
nor U3343 (N_3343,In_330,In_10);
xor U3344 (N_3344,In_991,In_197);
and U3345 (N_3345,In_1530,In_1676);
xor U3346 (N_3346,In_2967,In_709);
or U3347 (N_3347,In_178,In_1125);
and U3348 (N_3348,In_2583,In_460);
and U3349 (N_3349,In_2794,In_881);
nor U3350 (N_3350,In_1292,In_1603);
nand U3351 (N_3351,In_2987,In_627);
and U3352 (N_3352,In_2162,In_933);
nand U3353 (N_3353,In_2610,In_964);
nor U3354 (N_3354,In_1461,In_67);
or U3355 (N_3355,In_1007,In_959);
nand U3356 (N_3356,In_2460,In_870);
or U3357 (N_3357,In_1311,In_521);
nand U3358 (N_3358,In_983,In_1865);
nor U3359 (N_3359,In_273,In_1588);
xnor U3360 (N_3360,In_507,In_156);
xor U3361 (N_3361,In_1599,In_975);
or U3362 (N_3362,In_1672,In_1509);
xnor U3363 (N_3363,In_1701,In_2368);
nor U3364 (N_3364,In_2067,In_2064);
nor U3365 (N_3365,In_1088,In_2119);
xor U3366 (N_3366,In_797,In_1180);
nand U3367 (N_3367,In_2205,In_1830);
or U3368 (N_3368,In_960,In_1913);
nor U3369 (N_3369,In_1808,In_1587);
nor U3370 (N_3370,In_156,In_755);
xnor U3371 (N_3371,In_45,In_914);
xnor U3372 (N_3372,In_1893,In_2246);
or U3373 (N_3373,In_1907,In_2818);
nand U3374 (N_3374,In_1478,In_1387);
xor U3375 (N_3375,In_754,In_1840);
xnor U3376 (N_3376,In_803,In_1888);
nor U3377 (N_3377,In_428,In_2736);
nand U3378 (N_3378,In_944,In_2195);
xnor U3379 (N_3379,In_2559,In_2785);
nor U3380 (N_3380,In_2210,In_2415);
nand U3381 (N_3381,In_2470,In_1878);
or U3382 (N_3382,In_507,In_2978);
nor U3383 (N_3383,In_2355,In_2979);
and U3384 (N_3384,In_2289,In_1278);
xor U3385 (N_3385,In_2938,In_1601);
or U3386 (N_3386,In_1600,In_2740);
nor U3387 (N_3387,In_1797,In_1375);
nor U3388 (N_3388,In_967,In_1806);
and U3389 (N_3389,In_468,In_826);
and U3390 (N_3390,In_799,In_442);
nor U3391 (N_3391,In_1520,In_1285);
nand U3392 (N_3392,In_775,In_1566);
or U3393 (N_3393,In_1611,In_1744);
and U3394 (N_3394,In_197,In_1350);
nand U3395 (N_3395,In_2817,In_387);
xnor U3396 (N_3396,In_2842,In_2491);
nor U3397 (N_3397,In_533,In_1144);
or U3398 (N_3398,In_1300,In_131);
or U3399 (N_3399,In_2116,In_2840);
nor U3400 (N_3400,In_1599,In_27);
xnor U3401 (N_3401,In_2401,In_2791);
xnor U3402 (N_3402,In_1798,In_2015);
nand U3403 (N_3403,In_103,In_88);
xor U3404 (N_3404,In_288,In_663);
and U3405 (N_3405,In_95,In_791);
or U3406 (N_3406,In_2499,In_2387);
nand U3407 (N_3407,In_2506,In_2385);
nor U3408 (N_3408,In_401,In_633);
and U3409 (N_3409,In_535,In_1362);
and U3410 (N_3410,In_1741,In_1935);
xnor U3411 (N_3411,In_2441,In_925);
nand U3412 (N_3412,In_1513,In_2132);
nor U3413 (N_3413,In_2237,In_2896);
xnor U3414 (N_3414,In_334,In_2647);
and U3415 (N_3415,In_2980,In_2709);
and U3416 (N_3416,In_2210,In_2678);
nor U3417 (N_3417,In_522,In_870);
or U3418 (N_3418,In_1794,In_19);
xnor U3419 (N_3419,In_698,In_1022);
xor U3420 (N_3420,In_2583,In_2032);
xnor U3421 (N_3421,In_2842,In_434);
and U3422 (N_3422,In_579,In_773);
nand U3423 (N_3423,In_164,In_1868);
and U3424 (N_3424,In_1779,In_2415);
nand U3425 (N_3425,In_1740,In_1770);
xnor U3426 (N_3426,In_1095,In_2491);
xor U3427 (N_3427,In_1815,In_419);
nand U3428 (N_3428,In_2588,In_30);
or U3429 (N_3429,In_533,In_1972);
and U3430 (N_3430,In_1164,In_2744);
nand U3431 (N_3431,In_237,In_696);
or U3432 (N_3432,In_2122,In_2508);
or U3433 (N_3433,In_38,In_185);
and U3434 (N_3434,In_2894,In_1776);
xnor U3435 (N_3435,In_1379,In_534);
nor U3436 (N_3436,In_2516,In_1069);
nand U3437 (N_3437,In_1623,In_1232);
xnor U3438 (N_3438,In_355,In_2115);
nor U3439 (N_3439,In_1821,In_2067);
nor U3440 (N_3440,In_2947,In_178);
nand U3441 (N_3441,In_1607,In_5);
nand U3442 (N_3442,In_2607,In_70);
nor U3443 (N_3443,In_473,In_1903);
nand U3444 (N_3444,In_1427,In_35);
and U3445 (N_3445,In_1809,In_2357);
or U3446 (N_3446,In_1355,In_849);
nor U3447 (N_3447,In_87,In_2095);
nand U3448 (N_3448,In_1314,In_1943);
xnor U3449 (N_3449,In_2110,In_2470);
nor U3450 (N_3450,In_2563,In_1327);
xor U3451 (N_3451,In_1187,In_1776);
and U3452 (N_3452,In_1249,In_1013);
and U3453 (N_3453,In_603,In_2580);
and U3454 (N_3454,In_460,In_2168);
nor U3455 (N_3455,In_367,In_2595);
or U3456 (N_3456,In_1803,In_2008);
and U3457 (N_3457,In_1478,In_1965);
or U3458 (N_3458,In_2726,In_2412);
xor U3459 (N_3459,In_2871,In_2622);
xnor U3460 (N_3460,In_2167,In_2484);
nand U3461 (N_3461,In_1542,In_910);
xor U3462 (N_3462,In_2487,In_51);
and U3463 (N_3463,In_2802,In_1962);
and U3464 (N_3464,In_2843,In_936);
and U3465 (N_3465,In_282,In_2155);
nand U3466 (N_3466,In_1761,In_606);
nand U3467 (N_3467,In_1520,In_232);
and U3468 (N_3468,In_1643,In_962);
and U3469 (N_3469,In_2930,In_568);
or U3470 (N_3470,In_1051,In_1744);
or U3471 (N_3471,In_775,In_1289);
nor U3472 (N_3472,In_1912,In_482);
and U3473 (N_3473,In_393,In_387);
nor U3474 (N_3474,In_1309,In_1513);
nor U3475 (N_3475,In_2114,In_1318);
xor U3476 (N_3476,In_1755,In_2803);
nand U3477 (N_3477,In_806,In_1767);
and U3478 (N_3478,In_38,In_979);
xnor U3479 (N_3479,In_1079,In_2163);
xnor U3480 (N_3480,In_589,In_1012);
or U3481 (N_3481,In_2710,In_1466);
nand U3482 (N_3482,In_1970,In_2583);
nand U3483 (N_3483,In_465,In_896);
nand U3484 (N_3484,In_2061,In_1872);
nor U3485 (N_3485,In_725,In_1964);
and U3486 (N_3486,In_905,In_2919);
and U3487 (N_3487,In_2078,In_2450);
xnor U3488 (N_3488,In_2613,In_1874);
or U3489 (N_3489,In_1914,In_2281);
and U3490 (N_3490,In_1302,In_18);
or U3491 (N_3491,In_2045,In_1416);
and U3492 (N_3492,In_2450,In_1978);
or U3493 (N_3493,In_687,In_608);
nor U3494 (N_3494,In_512,In_2052);
and U3495 (N_3495,In_362,In_2086);
and U3496 (N_3496,In_567,In_1504);
or U3497 (N_3497,In_2142,In_2811);
nand U3498 (N_3498,In_2193,In_1783);
nor U3499 (N_3499,In_2717,In_31);
nor U3500 (N_3500,In_1480,In_1656);
or U3501 (N_3501,In_2932,In_2212);
or U3502 (N_3502,In_769,In_842);
and U3503 (N_3503,In_1505,In_832);
nand U3504 (N_3504,In_795,In_2682);
or U3505 (N_3505,In_912,In_676);
nand U3506 (N_3506,In_1722,In_1597);
nor U3507 (N_3507,In_251,In_2736);
nand U3508 (N_3508,In_2366,In_1229);
nand U3509 (N_3509,In_65,In_367);
and U3510 (N_3510,In_1350,In_2995);
nand U3511 (N_3511,In_2519,In_232);
nand U3512 (N_3512,In_267,In_869);
nor U3513 (N_3513,In_2098,In_792);
or U3514 (N_3514,In_2066,In_490);
nor U3515 (N_3515,In_422,In_2853);
xor U3516 (N_3516,In_2635,In_2647);
nand U3517 (N_3517,In_2500,In_226);
and U3518 (N_3518,In_2204,In_2541);
and U3519 (N_3519,In_282,In_2919);
and U3520 (N_3520,In_266,In_763);
nor U3521 (N_3521,In_500,In_2093);
nor U3522 (N_3522,In_1222,In_2041);
or U3523 (N_3523,In_2935,In_1510);
or U3524 (N_3524,In_2858,In_944);
and U3525 (N_3525,In_701,In_2226);
and U3526 (N_3526,In_2221,In_1494);
nor U3527 (N_3527,In_2264,In_2236);
nor U3528 (N_3528,In_326,In_2049);
or U3529 (N_3529,In_2676,In_1691);
or U3530 (N_3530,In_279,In_1586);
nand U3531 (N_3531,In_1474,In_1829);
nor U3532 (N_3532,In_975,In_2930);
and U3533 (N_3533,In_348,In_1540);
or U3534 (N_3534,In_988,In_1022);
nand U3535 (N_3535,In_1029,In_2264);
and U3536 (N_3536,In_566,In_867);
xnor U3537 (N_3537,In_2744,In_214);
or U3538 (N_3538,In_1781,In_992);
xnor U3539 (N_3539,In_1471,In_2395);
nand U3540 (N_3540,In_3,In_2568);
nor U3541 (N_3541,In_2527,In_93);
xnor U3542 (N_3542,In_2441,In_1860);
and U3543 (N_3543,In_1008,In_847);
and U3544 (N_3544,In_642,In_1687);
or U3545 (N_3545,In_345,In_578);
or U3546 (N_3546,In_831,In_62);
nor U3547 (N_3547,In_730,In_2398);
nor U3548 (N_3548,In_2531,In_403);
nor U3549 (N_3549,In_2716,In_475);
nor U3550 (N_3550,In_1560,In_1092);
nor U3551 (N_3551,In_2919,In_2890);
nor U3552 (N_3552,In_1757,In_1773);
xor U3553 (N_3553,In_1650,In_2834);
nand U3554 (N_3554,In_1472,In_661);
or U3555 (N_3555,In_1136,In_1164);
nor U3556 (N_3556,In_1869,In_2822);
nor U3557 (N_3557,In_18,In_1903);
nand U3558 (N_3558,In_2027,In_2071);
nand U3559 (N_3559,In_994,In_267);
and U3560 (N_3560,In_1914,In_486);
nand U3561 (N_3561,In_2137,In_566);
nand U3562 (N_3562,In_540,In_19);
xnor U3563 (N_3563,In_593,In_2352);
and U3564 (N_3564,In_607,In_2568);
and U3565 (N_3565,In_2746,In_1414);
xor U3566 (N_3566,In_124,In_1595);
or U3567 (N_3567,In_854,In_967);
nand U3568 (N_3568,In_1507,In_2108);
nand U3569 (N_3569,In_1887,In_1100);
and U3570 (N_3570,In_2920,In_1862);
or U3571 (N_3571,In_873,In_372);
nor U3572 (N_3572,In_2950,In_2788);
or U3573 (N_3573,In_946,In_2259);
nor U3574 (N_3574,In_849,In_2868);
xnor U3575 (N_3575,In_501,In_331);
xnor U3576 (N_3576,In_1021,In_701);
or U3577 (N_3577,In_2116,In_76);
nand U3578 (N_3578,In_719,In_7);
nor U3579 (N_3579,In_990,In_678);
or U3580 (N_3580,In_1447,In_1323);
or U3581 (N_3581,In_947,In_993);
or U3582 (N_3582,In_1093,In_2871);
and U3583 (N_3583,In_1942,In_1634);
nor U3584 (N_3584,In_259,In_1668);
or U3585 (N_3585,In_1644,In_803);
xnor U3586 (N_3586,In_926,In_899);
and U3587 (N_3587,In_1740,In_2482);
nand U3588 (N_3588,In_471,In_217);
and U3589 (N_3589,In_2218,In_300);
nand U3590 (N_3590,In_300,In_2132);
nor U3591 (N_3591,In_1966,In_1408);
and U3592 (N_3592,In_1437,In_804);
or U3593 (N_3593,In_2285,In_247);
nor U3594 (N_3594,In_1451,In_2765);
nor U3595 (N_3595,In_2837,In_608);
or U3596 (N_3596,In_1163,In_2731);
and U3597 (N_3597,In_1427,In_1842);
nand U3598 (N_3598,In_787,In_2247);
nand U3599 (N_3599,In_1446,In_2640);
xor U3600 (N_3600,In_1603,In_471);
or U3601 (N_3601,In_132,In_1139);
and U3602 (N_3602,In_897,In_732);
xnor U3603 (N_3603,In_122,In_1467);
xor U3604 (N_3604,In_1683,In_938);
nor U3605 (N_3605,In_1362,In_1575);
or U3606 (N_3606,In_379,In_484);
or U3607 (N_3607,In_2880,In_505);
and U3608 (N_3608,In_2668,In_1022);
nor U3609 (N_3609,In_1590,In_2533);
nor U3610 (N_3610,In_294,In_444);
nor U3611 (N_3611,In_1583,In_585);
xor U3612 (N_3612,In_1549,In_1340);
xor U3613 (N_3613,In_423,In_237);
nor U3614 (N_3614,In_1692,In_1658);
or U3615 (N_3615,In_707,In_1059);
nand U3616 (N_3616,In_2714,In_93);
xor U3617 (N_3617,In_1972,In_1228);
and U3618 (N_3618,In_1009,In_2968);
xnor U3619 (N_3619,In_1585,In_712);
and U3620 (N_3620,In_489,In_2265);
or U3621 (N_3621,In_2715,In_2125);
nand U3622 (N_3622,In_116,In_1248);
nand U3623 (N_3623,In_1275,In_2847);
or U3624 (N_3624,In_2362,In_2439);
xnor U3625 (N_3625,In_768,In_1382);
and U3626 (N_3626,In_2018,In_2861);
xor U3627 (N_3627,In_2549,In_2384);
xnor U3628 (N_3628,In_1852,In_2159);
or U3629 (N_3629,In_481,In_374);
or U3630 (N_3630,In_2549,In_352);
and U3631 (N_3631,In_1173,In_1597);
and U3632 (N_3632,In_2435,In_1202);
and U3633 (N_3633,In_531,In_412);
xnor U3634 (N_3634,In_166,In_2146);
nand U3635 (N_3635,In_1266,In_249);
nand U3636 (N_3636,In_1402,In_183);
nand U3637 (N_3637,In_1056,In_1337);
and U3638 (N_3638,In_905,In_791);
nand U3639 (N_3639,In_1124,In_1458);
xor U3640 (N_3640,In_227,In_601);
xor U3641 (N_3641,In_1751,In_2089);
xnor U3642 (N_3642,In_231,In_2839);
nand U3643 (N_3643,In_1664,In_2274);
xnor U3644 (N_3644,In_1235,In_2560);
or U3645 (N_3645,In_2815,In_1633);
nor U3646 (N_3646,In_914,In_276);
or U3647 (N_3647,In_2548,In_28);
nor U3648 (N_3648,In_2753,In_2552);
xor U3649 (N_3649,In_1270,In_1454);
nand U3650 (N_3650,In_1928,In_958);
or U3651 (N_3651,In_245,In_65);
or U3652 (N_3652,In_897,In_1782);
xnor U3653 (N_3653,In_241,In_1869);
or U3654 (N_3654,In_2025,In_2892);
nor U3655 (N_3655,In_446,In_28);
nor U3656 (N_3656,In_192,In_966);
or U3657 (N_3657,In_565,In_1026);
or U3658 (N_3658,In_2766,In_1265);
or U3659 (N_3659,In_355,In_2667);
and U3660 (N_3660,In_1067,In_129);
or U3661 (N_3661,In_1118,In_2388);
nand U3662 (N_3662,In_940,In_2401);
or U3663 (N_3663,In_2303,In_2902);
or U3664 (N_3664,In_309,In_2313);
nand U3665 (N_3665,In_2303,In_2715);
or U3666 (N_3666,In_2291,In_465);
and U3667 (N_3667,In_366,In_996);
xor U3668 (N_3668,In_2911,In_1510);
nor U3669 (N_3669,In_517,In_2744);
nand U3670 (N_3670,In_1677,In_1926);
or U3671 (N_3671,In_938,In_919);
xor U3672 (N_3672,In_11,In_379);
or U3673 (N_3673,In_217,In_2627);
nor U3674 (N_3674,In_1933,In_1172);
and U3675 (N_3675,In_372,In_424);
nor U3676 (N_3676,In_1670,In_988);
xor U3677 (N_3677,In_452,In_545);
nand U3678 (N_3678,In_181,In_1825);
xor U3679 (N_3679,In_1536,In_2222);
nand U3680 (N_3680,In_152,In_2928);
nand U3681 (N_3681,In_738,In_684);
nor U3682 (N_3682,In_1717,In_1791);
nand U3683 (N_3683,In_523,In_2182);
xor U3684 (N_3684,In_214,In_1042);
or U3685 (N_3685,In_576,In_337);
and U3686 (N_3686,In_2513,In_2190);
xnor U3687 (N_3687,In_1800,In_1514);
nand U3688 (N_3688,In_2661,In_1340);
and U3689 (N_3689,In_2720,In_1247);
or U3690 (N_3690,In_1616,In_1387);
nand U3691 (N_3691,In_2490,In_2713);
or U3692 (N_3692,In_1404,In_77);
xnor U3693 (N_3693,In_553,In_1870);
xor U3694 (N_3694,In_1627,In_2723);
or U3695 (N_3695,In_2693,In_1936);
and U3696 (N_3696,In_802,In_2217);
or U3697 (N_3697,In_401,In_2960);
nor U3698 (N_3698,In_2684,In_1628);
xor U3699 (N_3699,In_223,In_751);
xnor U3700 (N_3700,In_2209,In_707);
nor U3701 (N_3701,In_292,In_1810);
or U3702 (N_3702,In_1970,In_487);
xnor U3703 (N_3703,In_1011,In_191);
or U3704 (N_3704,In_1820,In_780);
nor U3705 (N_3705,In_2684,In_1797);
xor U3706 (N_3706,In_1205,In_1424);
and U3707 (N_3707,In_2245,In_1933);
or U3708 (N_3708,In_428,In_2274);
nor U3709 (N_3709,In_2829,In_2485);
or U3710 (N_3710,In_1077,In_1528);
or U3711 (N_3711,In_895,In_1599);
nor U3712 (N_3712,In_395,In_1167);
or U3713 (N_3713,In_672,In_1022);
nand U3714 (N_3714,In_1304,In_1415);
xnor U3715 (N_3715,In_2708,In_120);
nor U3716 (N_3716,In_1815,In_695);
nand U3717 (N_3717,In_1464,In_1566);
and U3718 (N_3718,In_723,In_653);
nand U3719 (N_3719,In_2701,In_2892);
nand U3720 (N_3720,In_2324,In_2565);
nor U3721 (N_3721,In_1481,In_2548);
or U3722 (N_3722,In_1945,In_1496);
and U3723 (N_3723,In_1068,In_605);
nor U3724 (N_3724,In_774,In_2074);
or U3725 (N_3725,In_2592,In_1202);
nor U3726 (N_3726,In_1272,In_355);
nor U3727 (N_3727,In_1917,In_514);
or U3728 (N_3728,In_337,In_526);
and U3729 (N_3729,In_1302,In_1464);
and U3730 (N_3730,In_2563,In_427);
nor U3731 (N_3731,In_591,In_77);
nand U3732 (N_3732,In_2818,In_2189);
nand U3733 (N_3733,In_1089,In_730);
nand U3734 (N_3734,In_2773,In_2554);
xor U3735 (N_3735,In_393,In_873);
xor U3736 (N_3736,In_973,In_1802);
and U3737 (N_3737,In_2633,In_1148);
nor U3738 (N_3738,In_1298,In_1097);
and U3739 (N_3739,In_1725,In_2687);
xor U3740 (N_3740,In_1557,In_1603);
or U3741 (N_3741,In_2608,In_1881);
and U3742 (N_3742,In_1306,In_1795);
xnor U3743 (N_3743,In_304,In_346);
xnor U3744 (N_3744,In_1569,In_784);
and U3745 (N_3745,In_1637,In_262);
nand U3746 (N_3746,In_488,In_1498);
or U3747 (N_3747,In_2544,In_1566);
xnor U3748 (N_3748,In_974,In_1079);
or U3749 (N_3749,In_52,In_1191);
or U3750 (N_3750,In_2837,In_1507);
nor U3751 (N_3751,In_2978,In_1880);
xor U3752 (N_3752,In_1123,In_2329);
nor U3753 (N_3753,In_1861,In_1878);
and U3754 (N_3754,In_2657,In_794);
xnor U3755 (N_3755,In_2995,In_2060);
nand U3756 (N_3756,In_716,In_2281);
or U3757 (N_3757,In_2640,In_1185);
nor U3758 (N_3758,In_1278,In_2667);
xor U3759 (N_3759,In_2165,In_772);
nor U3760 (N_3760,In_1596,In_25);
and U3761 (N_3761,In_6,In_812);
nand U3762 (N_3762,In_220,In_2099);
nand U3763 (N_3763,In_2922,In_1906);
or U3764 (N_3764,In_753,In_907);
and U3765 (N_3765,In_1071,In_1173);
nor U3766 (N_3766,In_2147,In_2173);
or U3767 (N_3767,In_2027,In_1461);
nor U3768 (N_3768,In_1723,In_2548);
xor U3769 (N_3769,In_1464,In_280);
nand U3770 (N_3770,In_774,In_917);
or U3771 (N_3771,In_104,In_408);
and U3772 (N_3772,In_885,In_2862);
nand U3773 (N_3773,In_748,In_1563);
nor U3774 (N_3774,In_732,In_2358);
xor U3775 (N_3775,In_1669,In_1635);
or U3776 (N_3776,In_1113,In_243);
xnor U3777 (N_3777,In_2888,In_2473);
nor U3778 (N_3778,In_785,In_2984);
nor U3779 (N_3779,In_2777,In_698);
and U3780 (N_3780,In_2137,In_1598);
and U3781 (N_3781,In_2301,In_525);
nand U3782 (N_3782,In_1527,In_933);
nor U3783 (N_3783,In_366,In_887);
nand U3784 (N_3784,In_1716,In_509);
xor U3785 (N_3785,In_239,In_146);
or U3786 (N_3786,In_175,In_1728);
or U3787 (N_3787,In_1865,In_195);
and U3788 (N_3788,In_2694,In_2807);
nor U3789 (N_3789,In_1103,In_747);
nor U3790 (N_3790,In_2708,In_662);
and U3791 (N_3791,In_1785,In_1688);
nor U3792 (N_3792,In_710,In_1732);
and U3793 (N_3793,In_1205,In_1312);
nor U3794 (N_3794,In_1402,In_447);
xor U3795 (N_3795,In_81,In_442);
and U3796 (N_3796,In_260,In_312);
and U3797 (N_3797,In_1838,In_100);
xor U3798 (N_3798,In_2652,In_2510);
nor U3799 (N_3799,In_2941,In_2095);
xnor U3800 (N_3800,In_2899,In_2955);
nand U3801 (N_3801,In_2018,In_2929);
nand U3802 (N_3802,In_2795,In_1504);
nand U3803 (N_3803,In_764,In_1638);
xor U3804 (N_3804,In_52,In_696);
nor U3805 (N_3805,In_1988,In_1928);
and U3806 (N_3806,In_1739,In_3);
nand U3807 (N_3807,In_2615,In_1056);
nand U3808 (N_3808,In_493,In_442);
xor U3809 (N_3809,In_2055,In_1016);
or U3810 (N_3810,In_709,In_1350);
xnor U3811 (N_3811,In_444,In_2885);
and U3812 (N_3812,In_2226,In_1429);
and U3813 (N_3813,In_1502,In_763);
nor U3814 (N_3814,In_460,In_776);
or U3815 (N_3815,In_664,In_888);
or U3816 (N_3816,In_2945,In_2486);
xor U3817 (N_3817,In_1569,In_1378);
and U3818 (N_3818,In_2960,In_1068);
and U3819 (N_3819,In_2715,In_907);
nor U3820 (N_3820,In_125,In_2979);
nand U3821 (N_3821,In_2594,In_124);
nand U3822 (N_3822,In_810,In_1943);
nand U3823 (N_3823,In_830,In_2951);
nor U3824 (N_3824,In_444,In_1303);
and U3825 (N_3825,In_2430,In_319);
xnor U3826 (N_3826,In_567,In_316);
xor U3827 (N_3827,In_1495,In_436);
nand U3828 (N_3828,In_913,In_2400);
xnor U3829 (N_3829,In_983,In_1348);
and U3830 (N_3830,In_1067,In_979);
nor U3831 (N_3831,In_300,In_2339);
and U3832 (N_3832,In_2968,In_1043);
nor U3833 (N_3833,In_211,In_640);
and U3834 (N_3834,In_1485,In_2244);
and U3835 (N_3835,In_2848,In_844);
or U3836 (N_3836,In_718,In_2939);
and U3837 (N_3837,In_2505,In_2217);
nand U3838 (N_3838,In_286,In_603);
nand U3839 (N_3839,In_2438,In_2991);
nor U3840 (N_3840,In_913,In_1082);
and U3841 (N_3841,In_170,In_1109);
and U3842 (N_3842,In_1763,In_2455);
nor U3843 (N_3843,In_2530,In_1392);
nand U3844 (N_3844,In_2469,In_1035);
nand U3845 (N_3845,In_917,In_2372);
or U3846 (N_3846,In_1215,In_1873);
nor U3847 (N_3847,In_2652,In_781);
xor U3848 (N_3848,In_481,In_928);
xor U3849 (N_3849,In_823,In_110);
or U3850 (N_3850,In_2680,In_190);
nor U3851 (N_3851,In_711,In_1720);
or U3852 (N_3852,In_441,In_2200);
and U3853 (N_3853,In_1279,In_1463);
nor U3854 (N_3854,In_825,In_96);
and U3855 (N_3855,In_2933,In_640);
and U3856 (N_3856,In_2758,In_2742);
nand U3857 (N_3857,In_2134,In_2463);
and U3858 (N_3858,In_2483,In_2344);
and U3859 (N_3859,In_975,In_585);
and U3860 (N_3860,In_1518,In_1828);
and U3861 (N_3861,In_1485,In_2012);
and U3862 (N_3862,In_1684,In_732);
xor U3863 (N_3863,In_1152,In_2357);
nor U3864 (N_3864,In_942,In_611);
xnor U3865 (N_3865,In_2752,In_423);
nand U3866 (N_3866,In_1956,In_2806);
nor U3867 (N_3867,In_2036,In_193);
or U3868 (N_3868,In_2541,In_1113);
or U3869 (N_3869,In_2067,In_1749);
or U3870 (N_3870,In_851,In_2049);
nand U3871 (N_3871,In_620,In_288);
xor U3872 (N_3872,In_309,In_2438);
xor U3873 (N_3873,In_451,In_1909);
nand U3874 (N_3874,In_1323,In_504);
and U3875 (N_3875,In_359,In_1358);
nor U3876 (N_3876,In_824,In_1942);
nand U3877 (N_3877,In_701,In_2653);
nor U3878 (N_3878,In_1500,In_1833);
and U3879 (N_3879,In_1615,In_2189);
and U3880 (N_3880,In_1940,In_2368);
nand U3881 (N_3881,In_1029,In_563);
nand U3882 (N_3882,In_2383,In_551);
nand U3883 (N_3883,In_832,In_1599);
or U3884 (N_3884,In_846,In_1169);
nand U3885 (N_3885,In_576,In_2493);
and U3886 (N_3886,In_1229,In_46);
or U3887 (N_3887,In_186,In_493);
and U3888 (N_3888,In_2220,In_1128);
or U3889 (N_3889,In_1386,In_1882);
xor U3890 (N_3890,In_984,In_1097);
and U3891 (N_3891,In_2911,In_232);
nor U3892 (N_3892,In_2664,In_358);
and U3893 (N_3893,In_3,In_455);
nor U3894 (N_3894,In_2935,In_1079);
nor U3895 (N_3895,In_1698,In_1015);
nor U3896 (N_3896,In_155,In_2925);
and U3897 (N_3897,In_246,In_322);
and U3898 (N_3898,In_2558,In_26);
or U3899 (N_3899,In_860,In_663);
nor U3900 (N_3900,In_2455,In_821);
xnor U3901 (N_3901,In_904,In_1341);
and U3902 (N_3902,In_500,In_1488);
and U3903 (N_3903,In_482,In_1451);
and U3904 (N_3904,In_560,In_83);
and U3905 (N_3905,In_2534,In_2338);
nor U3906 (N_3906,In_2616,In_1415);
nor U3907 (N_3907,In_2718,In_1110);
xnor U3908 (N_3908,In_2834,In_1033);
and U3909 (N_3909,In_158,In_1652);
nor U3910 (N_3910,In_285,In_2379);
nand U3911 (N_3911,In_122,In_2243);
and U3912 (N_3912,In_1795,In_600);
and U3913 (N_3913,In_2511,In_1508);
nor U3914 (N_3914,In_2773,In_544);
nand U3915 (N_3915,In_884,In_1902);
or U3916 (N_3916,In_1904,In_2402);
and U3917 (N_3917,In_1216,In_2895);
or U3918 (N_3918,In_2671,In_1562);
xnor U3919 (N_3919,In_365,In_1393);
nand U3920 (N_3920,In_2370,In_1561);
and U3921 (N_3921,In_785,In_2103);
or U3922 (N_3922,In_381,In_1724);
nand U3923 (N_3923,In_378,In_2964);
xor U3924 (N_3924,In_2737,In_170);
and U3925 (N_3925,In_2181,In_233);
or U3926 (N_3926,In_868,In_786);
and U3927 (N_3927,In_2405,In_601);
or U3928 (N_3928,In_643,In_1476);
nor U3929 (N_3929,In_109,In_234);
xor U3930 (N_3930,In_798,In_576);
and U3931 (N_3931,In_1703,In_1970);
xnor U3932 (N_3932,In_1421,In_768);
xnor U3933 (N_3933,In_2821,In_1678);
xnor U3934 (N_3934,In_1559,In_1628);
xnor U3935 (N_3935,In_2885,In_401);
nor U3936 (N_3936,In_1291,In_2308);
nor U3937 (N_3937,In_2105,In_553);
nand U3938 (N_3938,In_741,In_2981);
and U3939 (N_3939,In_824,In_711);
nand U3940 (N_3940,In_1684,In_2293);
xnor U3941 (N_3941,In_1459,In_2576);
or U3942 (N_3942,In_883,In_2365);
or U3943 (N_3943,In_2458,In_782);
xnor U3944 (N_3944,In_2084,In_2737);
nor U3945 (N_3945,In_2166,In_2675);
or U3946 (N_3946,In_1380,In_362);
nand U3947 (N_3947,In_717,In_177);
nor U3948 (N_3948,In_264,In_2705);
xnor U3949 (N_3949,In_2173,In_1658);
nor U3950 (N_3950,In_1760,In_2401);
nor U3951 (N_3951,In_2223,In_805);
and U3952 (N_3952,In_825,In_902);
nor U3953 (N_3953,In_1598,In_2188);
nor U3954 (N_3954,In_2192,In_1609);
nor U3955 (N_3955,In_2878,In_2868);
and U3956 (N_3956,In_1353,In_1556);
or U3957 (N_3957,In_1696,In_694);
xor U3958 (N_3958,In_825,In_1989);
xor U3959 (N_3959,In_2820,In_2341);
and U3960 (N_3960,In_2964,In_2796);
and U3961 (N_3961,In_1704,In_571);
xnor U3962 (N_3962,In_2172,In_1986);
xnor U3963 (N_3963,In_353,In_190);
and U3964 (N_3964,In_2439,In_2635);
xor U3965 (N_3965,In_2584,In_1303);
nand U3966 (N_3966,In_1075,In_2945);
and U3967 (N_3967,In_1198,In_985);
nor U3968 (N_3968,In_2359,In_2991);
xnor U3969 (N_3969,In_2016,In_429);
nor U3970 (N_3970,In_1839,In_912);
nor U3971 (N_3971,In_31,In_1280);
nor U3972 (N_3972,In_1865,In_793);
and U3973 (N_3973,In_685,In_1825);
and U3974 (N_3974,In_1148,In_1941);
nand U3975 (N_3975,In_1226,In_739);
nor U3976 (N_3976,In_969,In_616);
or U3977 (N_3977,In_2521,In_771);
nand U3978 (N_3978,In_1720,In_773);
or U3979 (N_3979,In_1377,In_2997);
nor U3980 (N_3980,In_2603,In_83);
xnor U3981 (N_3981,In_2488,In_2468);
nor U3982 (N_3982,In_82,In_2159);
and U3983 (N_3983,In_772,In_605);
nor U3984 (N_3984,In_454,In_2295);
nor U3985 (N_3985,In_1390,In_2641);
or U3986 (N_3986,In_1903,In_2883);
nor U3987 (N_3987,In_2629,In_680);
nand U3988 (N_3988,In_2196,In_1875);
or U3989 (N_3989,In_1098,In_2199);
or U3990 (N_3990,In_2853,In_115);
and U3991 (N_3991,In_2181,In_1576);
xnor U3992 (N_3992,In_1688,In_715);
nand U3993 (N_3993,In_582,In_2706);
xor U3994 (N_3994,In_2389,In_2702);
xor U3995 (N_3995,In_2384,In_928);
and U3996 (N_3996,In_759,In_2418);
nand U3997 (N_3997,In_1221,In_1817);
xor U3998 (N_3998,In_1494,In_1062);
nand U3999 (N_3999,In_1088,In_278);
xor U4000 (N_4000,In_2290,In_2298);
xnor U4001 (N_4001,In_2756,In_1752);
xnor U4002 (N_4002,In_2518,In_1101);
nand U4003 (N_4003,In_610,In_2309);
nor U4004 (N_4004,In_2822,In_754);
and U4005 (N_4005,In_1113,In_2123);
and U4006 (N_4006,In_813,In_1924);
nand U4007 (N_4007,In_141,In_2690);
and U4008 (N_4008,In_683,In_1298);
nor U4009 (N_4009,In_789,In_435);
nor U4010 (N_4010,In_46,In_2408);
xor U4011 (N_4011,In_904,In_1982);
nand U4012 (N_4012,In_1380,In_2400);
and U4013 (N_4013,In_1868,In_356);
or U4014 (N_4014,In_2783,In_373);
and U4015 (N_4015,In_2336,In_261);
nand U4016 (N_4016,In_335,In_236);
xnor U4017 (N_4017,In_1659,In_1117);
xnor U4018 (N_4018,In_2921,In_801);
or U4019 (N_4019,In_1204,In_2817);
nor U4020 (N_4020,In_2104,In_2189);
nor U4021 (N_4021,In_80,In_1979);
nor U4022 (N_4022,In_2204,In_1293);
xor U4023 (N_4023,In_1157,In_759);
nand U4024 (N_4024,In_1670,In_1957);
nor U4025 (N_4025,In_2916,In_2746);
nand U4026 (N_4026,In_1504,In_2960);
nor U4027 (N_4027,In_451,In_1614);
nand U4028 (N_4028,In_2242,In_2865);
xor U4029 (N_4029,In_738,In_2);
or U4030 (N_4030,In_729,In_913);
or U4031 (N_4031,In_452,In_2852);
nor U4032 (N_4032,In_765,In_77);
nor U4033 (N_4033,In_294,In_1557);
nor U4034 (N_4034,In_132,In_214);
or U4035 (N_4035,In_2104,In_1658);
xor U4036 (N_4036,In_2777,In_19);
nor U4037 (N_4037,In_1249,In_883);
or U4038 (N_4038,In_2805,In_733);
or U4039 (N_4039,In_2569,In_698);
nor U4040 (N_4040,In_2060,In_1329);
or U4041 (N_4041,In_431,In_1307);
xnor U4042 (N_4042,In_1792,In_2562);
nor U4043 (N_4043,In_1172,In_1735);
and U4044 (N_4044,In_1196,In_2768);
and U4045 (N_4045,In_1927,In_2294);
nand U4046 (N_4046,In_2227,In_1511);
and U4047 (N_4047,In_2908,In_1211);
xnor U4048 (N_4048,In_1268,In_2800);
and U4049 (N_4049,In_528,In_457);
nand U4050 (N_4050,In_1609,In_1698);
nand U4051 (N_4051,In_2535,In_69);
nand U4052 (N_4052,In_553,In_2754);
and U4053 (N_4053,In_1733,In_2154);
and U4054 (N_4054,In_2071,In_1497);
xor U4055 (N_4055,In_1743,In_2250);
or U4056 (N_4056,In_973,In_1383);
nand U4057 (N_4057,In_50,In_543);
and U4058 (N_4058,In_669,In_2558);
or U4059 (N_4059,In_1458,In_2681);
or U4060 (N_4060,In_740,In_580);
xor U4061 (N_4061,In_2039,In_2208);
or U4062 (N_4062,In_2375,In_874);
or U4063 (N_4063,In_768,In_2602);
and U4064 (N_4064,In_2993,In_1665);
nor U4065 (N_4065,In_1380,In_1926);
or U4066 (N_4066,In_2244,In_1760);
nor U4067 (N_4067,In_2636,In_2297);
or U4068 (N_4068,In_1511,In_277);
and U4069 (N_4069,In_1563,In_2466);
nor U4070 (N_4070,In_397,In_2172);
nand U4071 (N_4071,In_1603,In_2361);
or U4072 (N_4072,In_1805,In_2703);
nor U4073 (N_4073,In_171,In_2725);
and U4074 (N_4074,In_261,In_932);
and U4075 (N_4075,In_2622,In_1590);
xor U4076 (N_4076,In_2259,In_521);
nand U4077 (N_4077,In_2507,In_1120);
and U4078 (N_4078,In_963,In_1609);
or U4079 (N_4079,In_849,In_1431);
nor U4080 (N_4080,In_356,In_861);
and U4081 (N_4081,In_2971,In_1622);
nand U4082 (N_4082,In_2402,In_2137);
xor U4083 (N_4083,In_1511,In_2925);
xnor U4084 (N_4084,In_100,In_874);
and U4085 (N_4085,In_1006,In_1197);
or U4086 (N_4086,In_2402,In_1540);
and U4087 (N_4087,In_423,In_1048);
and U4088 (N_4088,In_2759,In_2797);
nor U4089 (N_4089,In_701,In_2027);
xnor U4090 (N_4090,In_1992,In_2492);
or U4091 (N_4091,In_495,In_2020);
nor U4092 (N_4092,In_2902,In_1994);
xor U4093 (N_4093,In_2872,In_2190);
or U4094 (N_4094,In_2516,In_293);
or U4095 (N_4095,In_2360,In_332);
or U4096 (N_4096,In_2767,In_2397);
xor U4097 (N_4097,In_371,In_1318);
nand U4098 (N_4098,In_2625,In_178);
nand U4099 (N_4099,In_85,In_2456);
xor U4100 (N_4100,In_1158,In_2318);
or U4101 (N_4101,In_1058,In_201);
nor U4102 (N_4102,In_2988,In_2084);
nand U4103 (N_4103,In_2089,In_647);
nor U4104 (N_4104,In_477,In_1372);
xor U4105 (N_4105,In_951,In_995);
or U4106 (N_4106,In_74,In_152);
and U4107 (N_4107,In_317,In_2664);
nor U4108 (N_4108,In_2884,In_828);
nor U4109 (N_4109,In_756,In_1187);
nor U4110 (N_4110,In_1283,In_1837);
xor U4111 (N_4111,In_704,In_1189);
and U4112 (N_4112,In_1012,In_2338);
nor U4113 (N_4113,In_974,In_907);
and U4114 (N_4114,In_805,In_43);
or U4115 (N_4115,In_493,In_1998);
xnor U4116 (N_4116,In_2583,In_2483);
or U4117 (N_4117,In_1177,In_2261);
xor U4118 (N_4118,In_2853,In_2191);
and U4119 (N_4119,In_179,In_896);
or U4120 (N_4120,In_423,In_2341);
xor U4121 (N_4121,In_778,In_756);
or U4122 (N_4122,In_2374,In_1421);
and U4123 (N_4123,In_2559,In_876);
nor U4124 (N_4124,In_578,In_929);
xor U4125 (N_4125,In_1844,In_41);
and U4126 (N_4126,In_87,In_501);
or U4127 (N_4127,In_1649,In_2488);
and U4128 (N_4128,In_126,In_1958);
and U4129 (N_4129,In_823,In_2042);
and U4130 (N_4130,In_1714,In_1305);
and U4131 (N_4131,In_1055,In_1917);
nand U4132 (N_4132,In_2154,In_2238);
nor U4133 (N_4133,In_943,In_2049);
or U4134 (N_4134,In_2004,In_2895);
xor U4135 (N_4135,In_560,In_1565);
nor U4136 (N_4136,In_1850,In_2868);
nor U4137 (N_4137,In_2750,In_2277);
nand U4138 (N_4138,In_1157,In_1988);
and U4139 (N_4139,In_1644,In_2150);
or U4140 (N_4140,In_973,In_621);
xor U4141 (N_4141,In_766,In_913);
xor U4142 (N_4142,In_22,In_1149);
nand U4143 (N_4143,In_1717,In_1319);
nor U4144 (N_4144,In_1821,In_1437);
and U4145 (N_4145,In_1424,In_2251);
xnor U4146 (N_4146,In_384,In_1635);
nor U4147 (N_4147,In_914,In_442);
xnor U4148 (N_4148,In_189,In_1268);
nand U4149 (N_4149,In_1402,In_2855);
nor U4150 (N_4150,In_2687,In_2074);
nor U4151 (N_4151,In_1939,In_1853);
xor U4152 (N_4152,In_2400,In_533);
nor U4153 (N_4153,In_28,In_1465);
nand U4154 (N_4154,In_1886,In_1144);
and U4155 (N_4155,In_1138,In_1751);
nor U4156 (N_4156,In_1500,In_2606);
xor U4157 (N_4157,In_1432,In_535);
nor U4158 (N_4158,In_2963,In_781);
and U4159 (N_4159,In_375,In_1628);
nand U4160 (N_4160,In_2850,In_1231);
or U4161 (N_4161,In_2316,In_544);
or U4162 (N_4162,In_1304,In_1138);
nor U4163 (N_4163,In_1333,In_467);
or U4164 (N_4164,In_173,In_2135);
nand U4165 (N_4165,In_42,In_1937);
nor U4166 (N_4166,In_719,In_202);
or U4167 (N_4167,In_2908,In_668);
nand U4168 (N_4168,In_1096,In_1620);
and U4169 (N_4169,In_1674,In_502);
and U4170 (N_4170,In_1396,In_2114);
nor U4171 (N_4171,In_906,In_293);
or U4172 (N_4172,In_1283,In_2188);
nand U4173 (N_4173,In_1107,In_2184);
and U4174 (N_4174,In_108,In_2015);
and U4175 (N_4175,In_2014,In_2357);
xnor U4176 (N_4176,In_2002,In_34);
nor U4177 (N_4177,In_635,In_1814);
xnor U4178 (N_4178,In_1784,In_604);
xnor U4179 (N_4179,In_1312,In_960);
or U4180 (N_4180,In_1590,In_1939);
and U4181 (N_4181,In_1968,In_2667);
and U4182 (N_4182,In_2129,In_2266);
nand U4183 (N_4183,In_731,In_2787);
nand U4184 (N_4184,In_2964,In_2378);
nor U4185 (N_4185,In_309,In_2437);
xnor U4186 (N_4186,In_555,In_1429);
nand U4187 (N_4187,In_2918,In_2126);
or U4188 (N_4188,In_1280,In_2909);
and U4189 (N_4189,In_1304,In_211);
or U4190 (N_4190,In_1023,In_2585);
nand U4191 (N_4191,In_2881,In_1460);
xor U4192 (N_4192,In_884,In_1042);
nor U4193 (N_4193,In_847,In_1306);
and U4194 (N_4194,In_1327,In_1030);
and U4195 (N_4195,In_1214,In_267);
and U4196 (N_4196,In_583,In_362);
or U4197 (N_4197,In_1458,In_2050);
and U4198 (N_4198,In_1148,In_1380);
nand U4199 (N_4199,In_896,In_1763);
and U4200 (N_4200,In_288,In_1200);
xnor U4201 (N_4201,In_2690,In_2688);
and U4202 (N_4202,In_2750,In_346);
nor U4203 (N_4203,In_2013,In_2101);
xnor U4204 (N_4204,In_1254,In_2318);
xnor U4205 (N_4205,In_2053,In_1921);
xor U4206 (N_4206,In_2612,In_140);
nand U4207 (N_4207,In_2604,In_1497);
nand U4208 (N_4208,In_1191,In_260);
xor U4209 (N_4209,In_20,In_1952);
nor U4210 (N_4210,In_1579,In_1654);
xor U4211 (N_4211,In_2676,In_887);
and U4212 (N_4212,In_1220,In_1042);
or U4213 (N_4213,In_1231,In_786);
xnor U4214 (N_4214,In_1437,In_221);
nand U4215 (N_4215,In_2089,In_2558);
and U4216 (N_4216,In_399,In_1395);
nor U4217 (N_4217,In_2906,In_7);
nand U4218 (N_4218,In_607,In_379);
and U4219 (N_4219,In_265,In_1463);
nor U4220 (N_4220,In_2729,In_1297);
xor U4221 (N_4221,In_307,In_1663);
or U4222 (N_4222,In_51,In_1259);
or U4223 (N_4223,In_938,In_102);
nand U4224 (N_4224,In_1499,In_1338);
and U4225 (N_4225,In_520,In_1713);
xor U4226 (N_4226,In_199,In_2289);
xor U4227 (N_4227,In_2545,In_77);
xor U4228 (N_4228,In_1444,In_2882);
nor U4229 (N_4229,In_2087,In_308);
nand U4230 (N_4230,In_327,In_1957);
or U4231 (N_4231,In_1088,In_1543);
xor U4232 (N_4232,In_1497,In_1366);
xor U4233 (N_4233,In_1513,In_2068);
and U4234 (N_4234,In_1460,In_492);
xor U4235 (N_4235,In_708,In_1735);
or U4236 (N_4236,In_701,In_88);
and U4237 (N_4237,In_1087,In_477);
nor U4238 (N_4238,In_2531,In_50);
or U4239 (N_4239,In_1902,In_2141);
or U4240 (N_4240,In_362,In_38);
nand U4241 (N_4241,In_222,In_2052);
nand U4242 (N_4242,In_1511,In_2505);
and U4243 (N_4243,In_20,In_360);
nand U4244 (N_4244,In_299,In_1385);
nand U4245 (N_4245,In_2233,In_2213);
nand U4246 (N_4246,In_318,In_1160);
or U4247 (N_4247,In_2727,In_2062);
and U4248 (N_4248,In_2239,In_2946);
xnor U4249 (N_4249,In_750,In_684);
nand U4250 (N_4250,In_2169,In_2638);
xor U4251 (N_4251,In_100,In_2027);
nand U4252 (N_4252,In_614,In_1347);
nor U4253 (N_4253,In_2397,In_2892);
xnor U4254 (N_4254,In_1337,In_2803);
or U4255 (N_4255,In_2736,In_2590);
or U4256 (N_4256,In_608,In_1891);
nand U4257 (N_4257,In_889,In_377);
or U4258 (N_4258,In_53,In_2827);
and U4259 (N_4259,In_253,In_812);
or U4260 (N_4260,In_722,In_2000);
nand U4261 (N_4261,In_1720,In_2336);
or U4262 (N_4262,In_1528,In_1617);
xor U4263 (N_4263,In_1807,In_1250);
nor U4264 (N_4264,In_207,In_2402);
or U4265 (N_4265,In_1712,In_1918);
nor U4266 (N_4266,In_2867,In_1365);
nor U4267 (N_4267,In_1123,In_2070);
or U4268 (N_4268,In_2794,In_2129);
nand U4269 (N_4269,In_2383,In_2976);
nand U4270 (N_4270,In_2622,In_1019);
nor U4271 (N_4271,In_2313,In_2806);
nor U4272 (N_4272,In_2731,In_1048);
nand U4273 (N_4273,In_2421,In_2067);
nor U4274 (N_4274,In_2032,In_1179);
xor U4275 (N_4275,In_2841,In_2536);
nand U4276 (N_4276,In_1950,In_842);
nor U4277 (N_4277,In_174,In_1880);
and U4278 (N_4278,In_2962,In_87);
nand U4279 (N_4279,In_1909,In_2910);
or U4280 (N_4280,In_2666,In_514);
and U4281 (N_4281,In_416,In_940);
and U4282 (N_4282,In_1206,In_577);
nand U4283 (N_4283,In_660,In_1728);
nor U4284 (N_4284,In_2164,In_1837);
or U4285 (N_4285,In_1022,In_453);
xnor U4286 (N_4286,In_1587,In_2703);
or U4287 (N_4287,In_2625,In_2238);
xor U4288 (N_4288,In_693,In_2688);
xnor U4289 (N_4289,In_130,In_1714);
nor U4290 (N_4290,In_1917,In_1355);
nor U4291 (N_4291,In_2401,In_460);
xor U4292 (N_4292,In_2848,In_2982);
xnor U4293 (N_4293,In_765,In_1806);
or U4294 (N_4294,In_769,In_2809);
nor U4295 (N_4295,In_2788,In_2619);
xnor U4296 (N_4296,In_1436,In_893);
xnor U4297 (N_4297,In_321,In_302);
nor U4298 (N_4298,In_2889,In_194);
nor U4299 (N_4299,In_332,In_1626);
or U4300 (N_4300,In_2522,In_1241);
xnor U4301 (N_4301,In_1670,In_930);
xor U4302 (N_4302,In_1176,In_1049);
xnor U4303 (N_4303,In_871,In_210);
and U4304 (N_4304,In_1960,In_139);
or U4305 (N_4305,In_1155,In_891);
and U4306 (N_4306,In_700,In_595);
or U4307 (N_4307,In_1619,In_2659);
and U4308 (N_4308,In_2299,In_1490);
or U4309 (N_4309,In_2579,In_1551);
nor U4310 (N_4310,In_711,In_295);
and U4311 (N_4311,In_1685,In_2432);
xnor U4312 (N_4312,In_2591,In_10);
nor U4313 (N_4313,In_434,In_212);
xor U4314 (N_4314,In_2816,In_626);
or U4315 (N_4315,In_1372,In_1695);
nor U4316 (N_4316,In_1159,In_268);
and U4317 (N_4317,In_2889,In_1174);
nor U4318 (N_4318,In_358,In_1462);
and U4319 (N_4319,In_1689,In_661);
and U4320 (N_4320,In_587,In_2632);
or U4321 (N_4321,In_246,In_2220);
nor U4322 (N_4322,In_789,In_207);
and U4323 (N_4323,In_2005,In_2815);
nand U4324 (N_4324,In_1086,In_2499);
nand U4325 (N_4325,In_679,In_1407);
nor U4326 (N_4326,In_1060,In_269);
and U4327 (N_4327,In_1205,In_2750);
xor U4328 (N_4328,In_340,In_2276);
and U4329 (N_4329,In_1544,In_750);
or U4330 (N_4330,In_542,In_740);
and U4331 (N_4331,In_1219,In_371);
nor U4332 (N_4332,In_88,In_349);
and U4333 (N_4333,In_1836,In_1139);
and U4334 (N_4334,In_641,In_2079);
nand U4335 (N_4335,In_822,In_801);
nor U4336 (N_4336,In_308,In_150);
and U4337 (N_4337,In_381,In_1766);
or U4338 (N_4338,In_1945,In_1711);
and U4339 (N_4339,In_2508,In_1736);
and U4340 (N_4340,In_698,In_2476);
and U4341 (N_4341,In_2337,In_394);
or U4342 (N_4342,In_2081,In_1446);
and U4343 (N_4343,In_2150,In_2541);
nand U4344 (N_4344,In_460,In_1192);
and U4345 (N_4345,In_2749,In_280);
or U4346 (N_4346,In_725,In_39);
and U4347 (N_4347,In_1595,In_620);
nor U4348 (N_4348,In_799,In_1412);
xor U4349 (N_4349,In_2552,In_147);
or U4350 (N_4350,In_908,In_628);
nand U4351 (N_4351,In_2784,In_738);
nand U4352 (N_4352,In_816,In_1259);
or U4353 (N_4353,In_601,In_248);
xnor U4354 (N_4354,In_2505,In_2280);
or U4355 (N_4355,In_2364,In_2950);
nor U4356 (N_4356,In_1021,In_2575);
or U4357 (N_4357,In_1652,In_2462);
and U4358 (N_4358,In_660,In_411);
xnor U4359 (N_4359,In_2247,In_2564);
nor U4360 (N_4360,In_234,In_2493);
nand U4361 (N_4361,In_790,In_1659);
nor U4362 (N_4362,In_111,In_842);
nand U4363 (N_4363,In_2253,In_1509);
nor U4364 (N_4364,In_562,In_1473);
or U4365 (N_4365,In_2214,In_835);
or U4366 (N_4366,In_663,In_1884);
xnor U4367 (N_4367,In_1122,In_1417);
nor U4368 (N_4368,In_2864,In_2997);
nand U4369 (N_4369,In_919,In_848);
or U4370 (N_4370,In_218,In_2570);
or U4371 (N_4371,In_2219,In_2239);
and U4372 (N_4372,In_1781,In_1797);
nor U4373 (N_4373,In_996,In_31);
or U4374 (N_4374,In_2930,In_2514);
xor U4375 (N_4375,In_1068,In_2328);
xnor U4376 (N_4376,In_1812,In_1617);
xor U4377 (N_4377,In_1451,In_1791);
or U4378 (N_4378,In_644,In_1224);
nand U4379 (N_4379,In_293,In_1430);
and U4380 (N_4380,In_2633,In_1759);
or U4381 (N_4381,In_305,In_2845);
and U4382 (N_4382,In_1577,In_2287);
and U4383 (N_4383,In_2799,In_2257);
xnor U4384 (N_4384,In_2089,In_1249);
nand U4385 (N_4385,In_2017,In_640);
xnor U4386 (N_4386,In_552,In_1547);
nand U4387 (N_4387,In_1399,In_2975);
nor U4388 (N_4388,In_2027,In_781);
xor U4389 (N_4389,In_1040,In_1617);
nand U4390 (N_4390,In_1128,In_1293);
or U4391 (N_4391,In_2462,In_2418);
or U4392 (N_4392,In_425,In_2682);
xnor U4393 (N_4393,In_654,In_58);
and U4394 (N_4394,In_2507,In_2554);
and U4395 (N_4395,In_1617,In_769);
and U4396 (N_4396,In_49,In_2857);
and U4397 (N_4397,In_341,In_51);
nand U4398 (N_4398,In_679,In_2253);
and U4399 (N_4399,In_1679,In_2394);
nand U4400 (N_4400,In_36,In_2799);
and U4401 (N_4401,In_47,In_2776);
or U4402 (N_4402,In_2894,In_1726);
and U4403 (N_4403,In_2777,In_1455);
or U4404 (N_4404,In_2354,In_490);
and U4405 (N_4405,In_2104,In_1000);
xnor U4406 (N_4406,In_1353,In_722);
nand U4407 (N_4407,In_810,In_1357);
xnor U4408 (N_4408,In_2656,In_2015);
nand U4409 (N_4409,In_405,In_1733);
nor U4410 (N_4410,In_335,In_243);
xor U4411 (N_4411,In_1385,In_468);
nand U4412 (N_4412,In_198,In_2096);
nand U4413 (N_4413,In_2175,In_1628);
nand U4414 (N_4414,In_266,In_1751);
nand U4415 (N_4415,In_2661,In_356);
nor U4416 (N_4416,In_1177,In_1255);
and U4417 (N_4417,In_790,In_2460);
or U4418 (N_4418,In_917,In_2309);
xor U4419 (N_4419,In_560,In_2762);
nor U4420 (N_4420,In_2138,In_1275);
and U4421 (N_4421,In_1763,In_1459);
nand U4422 (N_4422,In_287,In_2589);
xnor U4423 (N_4423,In_1018,In_2958);
nor U4424 (N_4424,In_295,In_1060);
xnor U4425 (N_4425,In_2098,In_1728);
nor U4426 (N_4426,In_1091,In_1437);
and U4427 (N_4427,In_344,In_276);
xor U4428 (N_4428,In_406,In_376);
nand U4429 (N_4429,In_1070,In_2147);
and U4430 (N_4430,In_1911,In_2253);
xnor U4431 (N_4431,In_64,In_1592);
xnor U4432 (N_4432,In_890,In_151);
xnor U4433 (N_4433,In_402,In_2769);
or U4434 (N_4434,In_1217,In_1833);
xor U4435 (N_4435,In_2872,In_141);
and U4436 (N_4436,In_910,In_774);
nor U4437 (N_4437,In_1,In_920);
or U4438 (N_4438,In_1477,In_1267);
xor U4439 (N_4439,In_1486,In_261);
nor U4440 (N_4440,In_2858,In_2028);
nand U4441 (N_4441,In_2644,In_1294);
nand U4442 (N_4442,In_2120,In_74);
xnor U4443 (N_4443,In_2367,In_2647);
nand U4444 (N_4444,In_478,In_343);
nand U4445 (N_4445,In_2854,In_500);
nand U4446 (N_4446,In_1927,In_1438);
nand U4447 (N_4447,In_1492,In_587);
nor U4448 (N_4448,In_1454,In_2527);
xor U4449 (N_4449,In_166,In_1669);
xnor U4450 (N_4450,In_2874,In_2072);
or U4451 (N_4451,In_280,In_1266);
and U4452 (N_4452,In_2960,In_2295);
nand U4453 (N_4453,In_330,In_2262);
and U4454 (N_4454,In_2129,In_2123);
and U4455 (N_4455,In_2680,In_1060);
nand U4456 (N_4456,In_2030,In_1103);
nor U4457 (N_4457,In_1128,In_1960);
nor U4458 (N_4458,In_855,In_2759);
and U4459 (N_4459,In_2730,In_2360);
nor U4460 (N_4460,In_2730,In_1028);
or U4461 (N_4461,In_181,In_2281);
nor U4462 (N_4462,In_2323,In_2438);
xor U4463 (N_4463,In_2574,In_1478);
nand U4464 (N_4464,In_2178,In_2421);
and U4465 (N_4465,In_1497,In_2154);
nand U4466 (N_4466,In_1363,In_2848);
nand U4467 (N_4467,In_813,In_2172);
nor U4468 (N_4468,In_680,In_928);
or U4469 (N_4469,In_203,In_807);
or U4470 (N_4470,In_482,In_61);
nor U4471 (N_4471,In_1188,In_933);
xnor U4472 (N_4472,In_1230,In_444);
or U4473 (N_4473,In_2501,In_207);
nor U4474 (N_4474,In_1326,In_2176);
and U4475 (N_4475,In_854,In_843);
xnor U4476 (N_4476,In_2453,In_2580);
nand U4477 (N_4477,In_1332,In_550);
or U4478 (N_4478,In_593,In_2866);
nand U4479 (N_4479,In_2858,In_2645);
and U4480 (N_4480,In_2841,In_14);
and U4481 (N_4481,In_2945,In_2542);
nor U4482 (N_4482,In_2359,In_2238);
nand U4483 (N_4483,In_2650,In_2235);
nor U4484 (N_4484,In_2124,In_33);
xor U4485 (N_4485,In_460,In_2574);
or U4486 (N_4486,In_945,In_1261);
nor U4487 (N_4487,In_1829,In_773);
xnor U4488 (N_4488,In_2440,In_1737);
xor U4489 (N_4489,In_1613,In_2501);
nor U4490 (N_4490,In_54,In_1387);
or U4491 (N_4491,In_518,In_2383);
and U4492 (N_4492,In_119,In_1339);
and U4493 (N_4493,In_1849,In_1209);
nand U4494 (N_4494,In_1280,In_1661);
and U4495 (N_4495,In_391,In_2641);
nor U4496 (N_4496,In_1380,In_959);
or U4497 (N_4497,In_2570,In_1309);
or U4498 (N_4498,In_1306,In_1143);
or U4499 (N_4499,In_2744,In_312);
or U4500 (N_4500,In_966,In_420);
and U4501 (N_4501,In_703,In_923);
and U4502 (N_4502,In_2801,In_1903);
and U4503 (N_4503,In_1626,In_1390);
and U4504 (N_4504,In_2158,In_2256);
nand U4505 (N_4505,In_1110,In_1395);
xnor U4506 (N_4506,In_1539,In_2361);
nand U4507 (N_4507,In_2600,In_1743);
or U4508 (N_4508,In_80,In_2077);
xor U4509 (N_4509,In_1191,In_1549);
and U4510 (N_4510,In_1073,In_1926);
xor U4511 (N_4511,In_232,In_1028);
and U4512 (N_4512,In_2387,In_1390);
nand U4513 (N_4513,In_303,In_1379);
nor U4514 (N_4514,In_1647,In_2798);
nor U4515 (N_4515,In_1239,In_1609);
nor U4516 (N_4516,In_1190,In_414);
nor U4517 (N_4517,In_358,In_858);
xor U4518 (N_4518,In_222,In_1096);
xor U4519 (N_4519,In_2511,In_608);
and U4520 (N_4520,In_1169,In_2751);
or U4521 (N_4521,In_1517,In_892);
or U4522 (N_4522,In_1043,In_2120);
nor U4523 (N_4523,In_772,In_2646);
and U4524 (N_4524,In_2219,In_1843);
or U4525 (N_4525,In_1446,In_2633);
and U4526 (N_4526,In_2888,In_2168);
xnor U4527 (N_4527,In_527,In_1117);
and U4528 (N_4528,In_1907,In_320);
nand U4529 (N_4529,In_547,In_1124);
xor U4530 (N_4530,In_1090,In_1855);
nor U4531 (N_4531,In_1415,In_1457);
xnor U4532 (N_4532,In_2183,In_991);
nand U4533 (N_4533,In_2905,In_1355);
and U4534 (N_4534,In_1097,In_1631);
and U4535 (N_4535,In_2071,In_2938);
and U4536 (N_4536,In_962,In_994);
nor U4537 (N_4537,In_2270,In_488);
or U4538 (N_4538,In_1616,In_504);
xnor U4539 (N_4539,In_247,In_2577);
or U4540 (N_4540,In_1289,In_2746);
and U4541 (N_4541,In_1866,In_1404);
or U4542 (N_4542,In_130,In_2688);
or U4543 (N_4543,In_1716,In_1453);
or U4544 (N_4544,In_1298,In_1116);
xnor U4545 (N_4545,In_1805,In_491);
or U4546 (N_4546,In_475,In_851);
nor U4547 (N_4547,In_2631,In_408);
nor U4548 (N_4548,In_1565,In_1581);
and U4549 (N_4549,In_2965,In_1765);
xor U4550 (N_4550,In_2619,In_1858);
and U4551 (N_4551,In_1632,In_2052);
nand U4552 (N_4552,In_2456,In_1136);
nand U4553 (N_4553,In_2165,In_2213);
or U4554 (N_4554,In_2425,In_2628);
xor U4555 (N_4555,In_2059,In_2650);
nor U4556 (N_4556,In_2102,In_57);
or U4557 (N_4557,In_1107,In_2996);
xnor U4558 (N_4558,In_1645,In_2635);
nand U4559 (N_4559,In_1622,In_538);
and U4560 (N_4560,In_643,In_2894);
xnor U4561 (N_4561,In_935,In_1368);
nor U4562 (N_4562,In_468,In_2116);
or U4563 (N_4563,In_293,In_1943);
xnor U4564 (N_4564,In_1549,In_1568);
nor U4565 (N_4565,In_2384,In_2768);
nor U4566 (N_4566,In_144,In_1231);
and U4567 (N_4567,In_2683,In_2841);
and U4568 (N_4568,In_493,In_1898);
and U4569 (N_4569,In_1070,In_232);
or U4570 (N_4570,In_1367,In_1213);
nor U4571 (N_4571,In_2554,In_50);
nor U4572 (N_4572,In_18,In_2978);
or U4573 (N_4573,In_2895,In_984);
xor U4574 (N_4574,In_1658,In_2163);
and U4575 (N_4575,In_2584,In_1959);
and U4576 (N_4576,In_2872,In_705);
nor U4577 (N_4577,In_1241,In_2288);
or U4578 (N_4578,In_66,In_2923);
nand U4579 (N_4579,In_2685,In_2294);
nand U4580 (N_4580,In_2766,In_1164);
and U4581 (N_4581,In_2532,In_1275);
or U4582 (N_4582,In_2398,In_1317);
xor U4583 (N_4583,In_1647,In_2052);
and U4584 (N_4584,In_1094,In_1604);
xor U4585 (N_4585,In_712,In_1303);
and U4586 (N_4586,In_177,In_1394);
nor U4587 (N_4587,In_2350,In_418);
or U4588 (N_4588,In_888,In_111);
and U4589 (N_4589,In_31,In_1725);
or U4590 (N_4590,In_174,In_1677);
xor U4591 (N_4591,In_421,In_2801);
or U4592 (N_4592,In_153,In_1270);
or U4593 (N_4593,In_1121,In_1396);
xor U4594 (N_4594,In_1219,In_1125);
nor U4595 (N_4595,In_1859,In_253);
xor U4596 (N_4596,In_554,In_263);
or U4597 (N_4597,In_611,In_2704);
nor U4598 (N_4598,In_2817,In_2392);
nand U4599 (N_4599,In_370,In_710);
or U4600 (N_4600,In_2924,In_315);
and U4601 (N_4601,In_2469,In_432);
nand U4602 (N_4602,In_709,In_1737);
and U4603 (N_4603,In_1281,In_2436);
nand U4604 (N_4604,In_976,In_500);
nor U4605 (N_4605,In_42,In_2241);
nor U4606 (N_4606,In_1120,In_2807);
xor U4607 (N_4607,In_841,In_2713);
nor U4608 (N_4608,In_2093,In_2830);
nor U4609 (N_4609,In_2622,In_2999);
or U4610 (N_4610,In_1189,In_1877);
xnor U4611 (N_4611,In_1063,In_1008);
xnor U4612 (N_4612,In_717,In_1544);
nor U4613 (N_4613,In_180,In_2003);
nor U4614 (N_4614,In_1120,In_2647);
nand U4615 (N_4615,In_2803,In_2594);
nor U4616 (N_4616,In_2523,In_1111);
xnor U4617 (N_4617,In_2355,In_1624);
xnor U4618 (N_4618,In_1591,In_2735);
and U4619 (N_4619,In_543,In_76);
nand U4620 (N_4620,In_1209,In_956);
xnor U4621 (N_4621,In_1532,In_2809);
and U4622 (N_4622,In_502,In_1514);
and U4623 (N_4623,In_1742,In_2423);
or U4624 (N_4624,In_2883,In_202);
nand U4625 (N_4625,In_468,In_110);
and U4626 (N_4626,In_2595,In_1956);
or U4627 (N_4627,In_1163,In_698);
nor U4628 (N_4628,In_230,In_1167);
xor U4629 (N_4629,In_508,In_1505);
xor U4630 (N_4630,In_333,In_1363);
nand U4631 (N_4631,In_118,In_955);
xor U4632 (N_4632,In_295,In_688);
and U4633 (N_4633,In_1163,In_2427);
or U4634 (N_4634,In_505,In_622);
or U4635 (N_4635,In_2036,In_1252);
or U4636 (N_4636,In_2746,In_1775);
xor U4637 (N_4637,In_1015,In_137);
or U4638 (N_4638,In_429,In_1341);
xor U4639 (N_4639,In_2504,In_2396);
nand U4640 (N_4640,In_784,In_145);
nand U4641 (N_4641,In_2169,In_1672);
xnor U4642 (N_4642,In_872,In_661);
nor U4643 (N_4643,In_750,In_1922);
nor U4644 (N_4644,In_268,In_2087);
and U4645 (N_4645,In_2452,In_883);
nor U4646 (N_4646,In_1919,In_429);
xnor U4647 (N_4647,In_1141,In_828);
and U4648 (N_4648,In_484,In_2293);
or U4649 (N_4649,In_1321,In_1087);
xnor U4650 (N_4650,In_2761,In_176);
and U4651 (N_4651,In_1859,In_2315);
or U4652 (N_4652,In_2280,In_2063);
or U4653 (N_4653,In_21,In_1302);
xnor U4654 (N_4654,In_2647,In_2424);
xnor U4655 (N_4655,In_1503,In_1826);
nor U4656 (N_4656,In_699,In_2086);
nand U4657 (N_4657,In_513,In_1566);
or U4658 (N_4658,In_1832,In_1173);
nor U4659 (N_4659,In_1009,In_125);
nand U4660 (N_4660,In_2243,In_588);
nand U4661 (N_4661,In_2201,In_406);
nand U4662 (N_4662,In_2990,In_28);
xnor U4663 (N_4663,In_1175,In_881);
and U4664 (N_4664,In_1243,In_1814);
and U4665 (N_4665,In_786,In_1939);
nand U4666 (N_4666,In_1303,In_1481);
xnor U4667 (N_4667,In_2880,In_2090);
nand U4668 (N_4668,In_1196,In_2034);
or U4669 (N_4669,In_819,In_764);
xnor U4670 (N_4670,In_2865,In_107);
nor U4671 (N_4671,In_818,In_1649);
nand U4672 (N_4672,In_2419,In_996);
or U4673 (N_4673,In_1560,In_2000);
or U4674 (N_4674,In_177,In_1023);
nor U4675 (N_4675,In_2562,In_2320);
xnor U4676 (N_4676,In_1159,In_2974);
and U4677 (N_4677,In_2721,In_2875);
nand U4678 (N_4678,In_1379,In_2776);
nand U4679 (N_4679,In_344,In_819);
nor U4680 (N_4680,In_2849,In_2563);
xor U4681 (N_4681,In_927,In_2498);
nor U4682 (N_4682,In_1448,In_2687);
nor U4683 (N_4683,In_1998,In_2901);
xor U4684 (N_4684,In_2228,In_1723);
and U4685 (N_4685,In_2500,In_2036);
xnor U4686 (N_4686,In_1201,In_990);
or U4687 (N_4687,In_2446,In_744);
and U4688 (N_4688,In_1441,In_2330);
nand U4689 (N_4689,In_298,In_1678);
or U4690 (N_4690,In_2717,In_1300);
and U4691 (N_4691,In_2311,In_1900);
and U4692 (N_4692,In_322,In_834);
and U4693 (N_4693,In_2679,In_1019);
nand U4694 (N_4694,In_2397,In_2612);
or U4695 (N_4695,In_1450,In_2722);
nor U4696 (N_4696,In_2045,In_2755);
xnor U4697 (N_4697,In_107,In_1579);
xnor U4698 (N_4698,In_2554,In_1832);
xnor U4699 (N_4699,In_2781,In_2063);
or U4700 (N_4700,In_1253,In_2682);
nor U4701 (N_4701,In_932,In_1330);
xor U4702 (N_4702,In_57,In_11);
nor U4703 (N_4703,In_2420,In_1665);
or U4704 (N_4704,In_1946,In_1832);
xor U4705 (N_4705,In_2742,In_2357);
nand U4706 (N_4706,In_1712,In_1573);
nand U4707 (N_4707,In_1449,In_2696);
or U4708 (N_4708,In_656,In_647);
nor U4709 (N_4709,In_360,In_2586);
xor U4710 (N_4710,In_1334,In_619);
xnor U4711 (N_4711,In_323,In_832);
or U4712 (N_4712,In_744,In_2140);
xnor U4713 (N_4713,In_1573,In_1283);
nor U4714 (N_4714,In_2257,In_877);
xnor U4715 (N_4715,In_1536,In_905);
xor U4716 (N_4716,In_767,In_2293);
nand U4717 (N_4717,In_1828,In_1055);
xor U4718 (N_4718,In_761,In_2655);
or U4719 (N_4719,In_980,In_93);
or U4720 (N_4720,In_1092,In_328);
and U4721 (N_4721,In_2221,In_292);
xor U4722 (N_4722,In_1083,In_2099);
nand U4723 (N_4723,In_617,In_270);
xnor U4724 (N_4724,In_1058,In_813);
or U4725 (N_4725,In_2930,In_1915);
nor U4726 (N_4726,In_838,In_517);
and U4727 (N_4727,In_755,In_831);
xor U4728 (N_4728,In_1868,In_84);
and U4729 (N_4729,In_2924,In_922);
or U4730 (N_4730,In_1475,In_722);
nand U4731 (N_4731,In_98,In_1753);
nor U4732 (N_4732,In_2300,In_2250);
or U4733 (N_4733,In_1757,In_230);
nor U4734 (N_4734,In_1675,In_995);
nor U4735 (N_4735,In_2631,In_295);
and U4736 (N_4736,In_265,In_2033);
nand U4737 (N_4737,In_456,In_1765);
xnor U4738 (N_4738,In_1346,In_284);
nor U4739 (N_4739,In_2874,In_2070);
nor U4740 (N_4740,In_232,In_1864);
xor U4741 (N_4741,In_2923,In_1381);
xnor U4742 (N_4742,In_2744,In_2965);
and U4743 (N_4743,In_1706,In_2579);
xnor U4744 (N_4744,In_586,In_2351);
or U4745 (N_4745,In_313,In_146);
and U4746 (N_4746,In_538,In_1561);
and U4747 (N_4747,In_489,In_210);
nand U4748 (N_4748,In_2857,In_1353);
xor U4749 (N_4749,In_578,In_2964);
and U4750 (N_4750,In_640,In_721);
and U4751 (N_4751,In_1214,In_1357);
nand U4752 (N_4752,In_1954,In_2996);
or U4753 (N_4753,In_11,In_2220);
nor U4754 (N_4754,In_273,In_2696);
or U4755 (N_4755,In_1613,In_109);
nor U4756 (N_4756,In_2541,In_2657);
nor U4757 (N_4757,In_2315,In_150);
nor U4758 (N_4758,In_376,In_2861);
nand U4759 (N_4759,In_52,In_1891);
nand U4760 (N_4760,In_1508,In_224);
nor U4761 (N_4761,In_771,In_523);
nand U4762 (N_4762,In_1165,In_654);
nand U4763 (N_4763,In_1386,In_2624);
nand U4764 (N_4764,In_2962,In_1128);
xnor U4765 (N_4765,In_1290,In_887);
xnor U4766 (N_4766,In_1109,In_2022);
and U4767 (N_4767,In_967,In_385);
or U4768 (N_4768,In_1258,In_1446);
and U4769 (N_4769,In_1074,In_2364);
and U4770 (N_4770,In_184,In_384);
or U4771 (N_4771,In_2327,In_239);
or U4772 (N_4772,In_646,In_254);
and U4773 (N_4773,In_284,In_1981);
and U4774 (N_4774,In_2366,In_840);
nor U4775 (N_4775,In_271,In_807);
or U4776 (N_4776,In_2093,In_2735);
or U4777 (N_4777,In_1270,In_1575);
or U4778 (N_4778,In_1333,In_1163);
and U4779 (N_4779,In_1593,In_2509);
nand U4780 (N_4780,In_2506,In_2613);
nand U4781 (N_4781,In_2598,In_1922);
nand U4782 (N_4782,In_1495,In_1133);
nand U4783 (N_4783,In_1564,In_1901);
xor U4784 (N_4784,In_475,In_2576);
nand U4785 (N_4785,In_2938,In_2943);
nor U4786 (N_4786,In_1207,In_2522);
or U4787 (N_4787,In_2397,In_701);
nand U4788 (N_4788,In_802,In_2669);
nor U4789 (N_4789,In_2497,In_234);
xnor U4790 (N_4790,In_1488,In_1070);
nand U4791 (N_4791,In_1850,In_2465);
xnor U4792 (N_4792,In_2909,In_2151);
and U4793 (N_4793,In_1660,In_2092);
nor U4794 (N_4794,In_1523,In_2);
nor U4795 (N_4795,In_1944,In_324);
nand U4796 (N_4796,In_2675,In_1311);
nand U4797 (N_4797,In_79,In_1294);
nor U4798 (N_4798,In_2149,In_2448);
xor U4799 (N_4799,In_506,In_862);
nand U4800 (N_4800,In_2743,In_1569);
nand U4801 (N_4801,In_728,In_1657);
xor U4802 (N_4802,In_1133,In_2095);
nor U4803 (N_4803,In_2166,In_1833);
nor U4804 (N_4804,In_470,In_2876);
nor U4805 (N_4805,In_553,In_1731);
xnor U4806 (N_4806,In_2927,In_159);
or U4807 (N_4807,In_88,In_2547);
nor U4808 (N_4808,In_1943,In_910);
nor U4809 (N_4809,In_1550,In_926);
or U4810 (N_4810,In_2602,In_1570);
or U4811 (N_4811,In_1005,In_2578);
or U4812 (N_4812,In_2920,In_153);
xor U4813 (N_4813,In_1050,In_2043);
nor U4814 (N_4814,In_1401,In_1544);
nand U4815 (N_4815,In_670,In_421);
xor U4816 (N_4816,In_928,In_329);
or U4817 (N_4817,In_1720,In_639);
xnor U4818 (N_4818,In_619,In_2296);
nand U4819 (N_4819,In_1360,In_477);
nand U4820 (N_4820,In_2122,In_1582);
nand U4821 (N_4821,In_2803,In_2163);
xor U4822 (N_4822,In_1464,In_2027);
xor U4823 (N_4823,In_2834,In_1160);
nand U4824 (N_4824,In_1442,In_2399);
nor U4825 (N_4825,In_2344,In_465);
or U4826 (N_4826,In_530,In_702);
nor U4827 (N_4827,In_2613,In_747);
nand U4828 (N_4828,In_929,In_1292);
and U4829 (N_4829,In_753,In_1672);
and U4830 (N_4830,In_2684,In_182);
and U4831 (N_4831,In_2736,In_417);
or U4832 (N_4832,In_2298,In_859);
or U4833 (N_4833,In_1492,In_1371);
or U4834 (N_4834,In_1139,In_231);
xnor U4835 (N_4835,In_1038,In_1275);
or U4836 (N_4836,In_1169,In_1223);
and U4837 (N_4837,In_2256,In_2539);
and U4838 (N_4838,In_1021,In_2436);
or U4839 (N_4839,In_1629,In_1152);
and U4840 (N_4840,In_1530,In_1036);
or U4841 (N_4841,In_231,In_726);
xor U4842 (N_4842,In_1520,In_2829);
and U4843 (N_4843,In_390,In_1972);
xnor U4844 (N_4844,In_65,In_2285);
nor U4845 (N_4845,In_165,In_1124);
nor U4846 (N_4846,In_2981,In_2313);
nor U4847 (N_4847,In_703,In_2670);
xnor U4848 (N_4848,In_25,In_475);
nand U4849 (N_4849,In_2784,In_238);
or U4850 (N_4850,In_1998,In_290);
nand U4851 (N_4851,In_179,In_2491);
and U4852 (N_4852,In_2779,In_2744);
or U4853 (N_4853,In_1098,In_326);
and U4854 (N_4854,In_1797,In_539);
and U4855 (N_4855,In_2734,In_1145);
or U4856 (N_4856,In_8,In_1210);
xor U4857 (N_4857,In_1282,In_793);
nand U4858 (N_4858,In_755,In_2025);
nor U4859 (N_4859,In_1493,In_1318);
xor U4860 (N_4860,In_2301,In_2426);
or U4861 (N_4861,In_2301,In_2478);
nand U4862 (N_4862,In_2357,In_939);
xnor U4863 (N_4863,In_2352,In_2448);
nor U4864 (N_4864,In_1088,In_2525);
nand U4865 (N_4865,In_2134,In_2832);
or U4866 (N_4866,In_503,In_2992);
and U4867 (N_4867,In_1306,In_2344);
and U4868 (N_4868,In_151,In_717);
nor U4869 (N_4869,In_638,In_377);
or U4870 (N_4870,In_2842,In_42);
or U4871 (N_4871,In_224,In_1257);
nand U4872 (N_4872,In_501,In_2359);
nand U4873 (N_4873,In_2194,In_1206);
nor U4874 (N_4874,In_874,In_1842);
nor U4875 (N_4875,In_2378,In_1293);
and U4876 (N_4876,In_2205,In_755);
and U4877 (N_4877,In_1725,In_2338);
and U4878 (N_4878,In_1626,In_2705);
nand U4879 (N_4879,In_2502,In_2727);
or U4880 (N_4880,In_2370,In_2131);
nand U4881 (N_4881,In_411,In_2344);
or U4882 (N_4882,In_17,In_1953);
nor U4883 (N_4883,In_1041,In_279);
nand U4884 (N_4884,In_2232,In_980);
nor U4885 (N_4885,In_2006,In_557);
nor U4886 (N_4886,In_738,In_2211);
xor U4887 (N_4887,In_354,In_971);
xnor U4888 (N_4888,In_1044,In_2320);
xnor U4889 (N_4889,In_2644,In_265);
nand U4890 (N_4890,In_837,In_588);
nor U4891 (N_4891,In_2959,In_1298);
nand U4892 (N_4892,In_971,In_2968);
or U4893 (N_4893,In_1741,In_2202);
and U4894 (N_4894,In_227,In_1541);
or U4895 (N_4895,In_841,In_2545);
and U4896 (N_4896,In_1462,In_1945);
nor U4897 (N_4897,In_418,In_1495);
xor U4898 (N_4898,In_361,In_1298);
nand U4899 (N_4899,In_2951,In_1485);
or U4900 (N_4900,In_1170,In_1669);
or U4901 (N_4901,In_828,In_206);
xnor U4902 (N_4902,In_572,In_971);
nor U4903 (N_4903,In_2130,In_2149);
and U4904 (N_4904,In_724,In_315);
and U4905 (N_4905,In_706,In_2791);
nand U4906 (N_4906,In_756,In_135);
nor U4907 (N_4907,In_2350,In_2281);
nand U4908 (N_4908,In_2731,In_600);
nor U4909 (N_4909,In_246,In_2543);
or U4910 (N_4910,In_1941,In_987);
and U4911 (N_4911,In_2630,In_2671);
and U4912 (N_4912,In_1563,In_2235);
and U4913 (N_4913,In_1188,In_2253);
and U4914 (N_4914,In_2490,In_1526);
nand U4915 (N_4915,In_626,In_1939);
nor U4916 (N_4916,In_51,In_2029);
xnor U4917 (N_4917,In_1703,In_2420);
nor U4918 (N_4918,In_1738,In_688);
nand U4919 (N_4919,In_2647,In_986);
or U4920 (N_4920,In_2358,In_741);
nand U4921 (N_4921,In_1147,In_659);
xnor U4922 (N_4922,In_2674,In_1908);
nor U4923 (N_4923,In_1713,In_1342);
nand U4924 (N_4924,In_222,In_2137);
or U4925 (N_4925,In_2455,In_1940);
or U4926 (N_4926,In_2533,In_1947);
xor U4927 (N_4927,In_78,In_2619);
xnor U4928 (N_4928,In_1953,In_479);
and U4929 (N_4929,In_1681,In_2950);
and U4930 (N_4930,In_522,In_1108);
nand U4931 (N_4931,In_265,In_209);
and U4932 (N_4932,In_92,In_2128);
nor U4933 (N_4933,In_2119,In_412);
nor U4934 (N_4934,In_2157,In_528);
nand U4935 (N_4935,In_1335,In_2291);
nand U4936 (N_4936,In_1061,In_1878);
nor U4937 (N_4937,In_1207,In_2676);
or U4938 (N_4938,In_621,In_1277);
or U4939 (N_4939,In_64,In_1326);
nor U4940 (N_4940,In_162,In_574);
nand U4941 (N_4941,In_1754,In_2101);
nor U4942 (N_4942,In_1907,In_2988);
and U4943 (N_4943,In_2638,In_1631);
xnor U4944 (N_4944,In_2798,In_644);
xor U4945 (N_4945,In_2348,In_1082);
xnor U4946 (N_4946,In_266,In_1922);
or U4947 (N_4947,In_2346,In_910);
and U4948 (N_4948,In_311,In_500);
nor U4949 (N_4949,In_2612,In_789);
nor U4950 (N_4950,In_2618,In_1555);
and U4951 (N_4951,In_266,In_1483);
and U4952 (N_4952,In_1221,In_2284);
nor U4953 (N_4953,In_158,In_214);
and U4954 (N_4954,In_1702,In_2881);
and U4955 (N_4955,In_1691,In_2938);
xnor U4956 (N_4956,In_2353,In_2421);
or U4957 (N_4957,In_1915,In_2627);
and U4958 (N_4958,In_2522,In_2169);
nor U4959 (N_4959,In_2887,In_850);
nor U4960 (N_4960,In_1389,In_2219);
and U4961 (N_4961,In_2414,In_90);
or U4962 (N_4962,In_2049,In_1547);
and U4963 (N_4963,In_2012,In_2358);
xor U4964 (N_4964,In_1670,In_2909);
nand U4965 (N_4965,In_1258,In_689);
nand U4966 (N_4966,In_395,In_513);
xnor U4967 (N_4967,In_1203,In_2120);
nor U4968 (N_4968,In_557,In_2874);
or U4969 (N_4969,In_347,In_2267);
or U4970 (N_4970,In_1940,In_1194);
and U4971 (N_4971,In_2725,In_2605);
or U4972 (N_4972,In_1281,In_934);
nor U4973 (N_4973,In_419,In_2319);
xor U4974 (N_4974,In_1481,In_1036);
or U4975 (N_4975,In_1074,In_437);
nand U4976 (N_4976,In_1754,In_1074);
or U4977 (N_4977,In_2231,In_261);
nor U4978 (N_4978,In_2225,In_382);
nor U4979 (N_4979,In_2683,In_1286);
nor U4980 (N_4980,In_575,In_2317);
nor U4981 (N_4981,In_1044,In_451);
xor U4982 (N_4982,In_2140,In_1181);
or U4983 (N_4983,In_212,In_68);
nand U4984 (N_4984,In_1787,In_339);
nor U4985 (N_4985,In_1011,In_2015);
and U4986 (N_4986,In_781,In_2269);
or U4987 (N_4987,In_2129,In_650);
nand U4988 (N_4988,In_140,In_612);
nand U4989 (N_4989,In_414,In_1812);
xor U4990 (N_4990,In_274,In_906);
or U4991 (N_4991,In_470,In_913);
and U4992 (N_4992,In_842,In_2971);
xnor U4993 (N_4993,In_2002,In_156);
nor U4994 (N_4994,In_622,In_494);
and U4995 (N_4995,In_1311,In_1913);
and U4996 (N_4996,In_2463,In_1709);
nand U4997 (N_4997,In_2838,In_840);
nor U4998 (N_4998,In_31,In_1211);
nor U4999 (N_4999,In_2311,In_1771);
or U5000 (N_5000,N_4022,N_2250);
nand U5001 (N_5001,N_3706,N_3310);
and U5002 (N_5002,N_3365,N_1874);
nand U5003 (N_5003,N_587,N_3152);
and U5004 (N_5004,N_3574,N_942);
and U5005 (N_5005,N_205,N_2781);
xnor U5006 (N_5006,N_559,N_3969);
or U5007 (N_5007,N_1862,N_3539);
nand U5008 (N_5008,N_3733,N_3331);
or U5009 (N_5009,N_2759,N_451);
nor U5010 (N_5010,N_2367,N_506);
xor U5011 (N_5011,N_831,N_4799);
nor U5012 (N_5012,N_4178,N_2703);
nand U5013 (N_5013,N_2033,N_3529);
xnor U5014 (N_5014,N_784,N_4423);
nor U5015 (N_5015,N_4099,N_4051);
xor U5016 (N_5016,N_1484,N_3983);
nand U5017 (N_5017,N_420,N_2305);
xnor U5018 (N_5018,N_9,N_1181);
or U5019 (N_5019,N_310,N_4764);
nand U5020 (N_5020,N_2137,N_766);
xor U5021 (N_5021,N_1787,N_2417);
and U5022 (N_5022,N_3831,N_296);
nand U5023 (N_5023,N_3345,N_3013);
xor U5024 (N_5024,N_3887,N_1518);
xor U5025 (N_5025,N_2784,N_1587);
xor U5026 (N_5026,N_2618,N_1118);
nand U5027 (N_5027,N_3396,N_343);
nand U5028 (N_5028,N_2511,N_413);
and U5029 (N_5029,N_4006,N_2867);
nand U5030 (N_5030,N_351,N_3725);
nand U5031 (N_5031,N_100,N_525);
nand U5032 (N_5032,N_2188,N_3827);
or U5033 (N_5033,N_3193,N_4445);
xor U5034 (N_5034,N_3896,N_3314);
nand U5035 (N_5035,N_2197,N_2036);
nor U5036 (N_5036,N_3726,N_2174);
nand U5037 (N_5037,N_17,N_1114);
nand U5038 (N_5038,N_797,N_249);
or U5039 (N_5039,N_4595,N_1322);
nand U5040 (N_5040,N_1071,N_4730);
xor U5041 (N_5041,N_3940,N_4430);
or U5042 (N_5042,N_148,N_1182);
nor U5043 (N_5043,N_3260,N_4377);
and U5044 (N_5044,N_241,N_1526);
or U5045 (N_5045,N_1213,N_271);
xnor U5046 (N_5046,N_3103,N_2030);
and U5047 (N_5047,N_3992,N_3342);
nand U5048 (N_5048,N_652,N_4875);
and U5049 (N_5049,N_1104,N_666);
or U5050 (N_5050,N_2870,N_907);
and U5051 (N_5051,N_4405,N_1632);
xnor U5052 (N_5052,N_558,N_2278);
or U5053 (N_5053,N_626,N_4741);
nand U5054 (N_5054,N_2873,N_1225);
nor U5055 (N_5055,N_605,N_2000);
xnor U5056 (N_5056,N_1726,N_439);
nor U5057 (N_5057,N_2762,N_1817);
and U5058 (N_5058,N_4695,N_263);
xor U5059 (N_5059,N_1597,N_260);
or U5060 (N_5060,N_1543,N_863);
and U5061 (N_5061,N_4633,N_4743);
nand U5062 (N_5062,N_2946,N_162);
or U5063 (N_5063,N_2459,N_2653);
nor U5064 (N_5064,N_870,N_673);
xor U5065 (N_5065,N_865,N_2735);
xor U5066 (N_5066,N_4355,N_2347);
nand U5067 (N_5067,N_679,N_4637);
nor U5068 (N_5068,N_2930,N_767);
xor U5069 (N_5069,N_920,N_3130);
and U5070 (N_5070,N_1220,N_3366);
xor U5071 (N_5071,N_3868,N_1955);
nor U5072 (N_5072,N_4837,N_1900);
or U5073 (N_5073,N_2374,N_3120);
nand U5074 (N_5074,N_1873,N_4465);
xor U5075 (N_5075,N_2026,N_3466);
nand U5076 (N_5076,N_1139,N_3339);
nand U5077 (N_5077,N_1984,N_3836);
xor U5078 (N_5078,N_408,N_1174);
xor U5079 (N_5079,N_4946,N_4979);
nand U5080 (N_5080,N_3079,N_2106);
nor U5081 (N_5081,N_3343,N_2832);
nor U5082 (N_5082,N_4783,N_4719);
xor U5083 (N_5083,N_2922,N_1903);
and U5084 (N_5084,N_4521,N_3904);
or U5085 (N_5085,N_1827,N_1801);
or U5086 (N_5086,N_3768,N_4203);
xor U5087 (N_5087,N_1615,N_3481);
and U5088 (N_5088,N_2678,N_3008);
xnor U5089 (N_5089,N_4847,N_3709);
and U5090 (N_5090,N_435,N_1081);
or U5091 (N_5091,N_2982,N_3026);
and U5092 (N_5092,N_2632,N_2894);
nor U5093 (N_5093,N_1574,N_4326);
nor U5094 (N_5094,N_4149,N_3112);
or U5095 (N_5095,N_991,N_4863);
and U5096 (N_5096,N_30,N_2071);
xnor U5097 (N_5097,N_540,N_1812);
nor U5098 (N_5098,N_1284,N_1309);
nand U5099 (N_5099,N_892,N_3338);
nand U5100 (N_5100,N_2447,N_1033);
and U5101 (N_5101,N_3304,N_1111);
or U5102 (N_5102,N_951,N_2985);
xnor U5103 (N_5103,N_2998,N_1208);
or U5104 (N_5104,N_4693,N_2782);
nor U5105 (N_5105,N_820,N_819);
nand U5106 (N_5106,N_2282,N_4190);
nor U5107 (N_5107,N_2048,N_636);
xnor U5108 (N_5108,N_4587,N_1375);
nand U5109 (N_5109,N_2908,N_3843);
nor U5110 (N_5110,N_1261,N_4933);
or U5111 (N_5111,N_3235,N_1944);
nor U5112 (N_5112,N_749,N_2205);
and U5113 (N_5113,N_4842,N_2390);
or U5114 (N_5114,N_599,N_459);
nand U5115 (N_5115,N_3218,N_4329);
xnor U5116 (N_5116,N_3275,N_1476);
and U5117 (N_5117,N_1557,N_4852);
or U5118 (N_5118,N_1937,N_1363);
nor U5119 (N_5119,N_4116,N_4);
or U5120 (N_5120,N_3579,N_3611);
and U5121 (N_5121,N_1788,N_3938);
xnor U5122 (N_5122,N_2542,N_4573);
nor U5123 (N_5123,N_3866,N_3067);
and U5124 (N_5124,N_826,N_614);
nor U5125 (N_5125,N_1214,N_2302);
or U5126 (N_5126,N_2338,N_2151);
xnor U5127 (N_5127,N_4610,N_3771);
or U5128 (N_5128,N_3714,N_2012);
xor U5129 (N_5129,N_2220,N_4762);
xor U5130 (N_5130,N_1443,N_4824);
and U5131 (N_5131,N_4567,N_2830);
xnor U5132 (N_5132,N_2791,N_4963);
nand U5133 (N_5133,N_3181,N_2163);
nand U5134 (N_5134,N_2105,N_438);
xnor U5135 (N_5135,N_2642,N_4958);
and U5136 (N_5136,N_989,N_1028);
and U5137 (N_5137,N_2715,N_1973);
xnor U5138 (N_5138,N_616,N_837);
and U5139 (N_5139,N_4474,N_2175);
nand U5140 (N_5140,N_2740,N_4578);
nor U5141 (N_5141,N_4155,N_3608);
xnor U5142 (N_5142,N_2724,N_1527);
nand U5143 (N_5143,N_2441,N_3662);
nor U5144 (N_5144,N_3212,N_3609);
and U5145 (N_5145,N_732,N_4194);
nand U5146 (N_5146,N_3948,N_4471);
nand U5147 (N_5147,N_1292,N_1079);
xor U5148 (N_5148,N_3164,N_3773);
or U5149 (N_5149,N_4612,N_4057);
xor U5150 (N_5150,N_2321,N_3142);
nand U5151 (N_5151,N_1659,N_1537);
nand U5152 (N_5152,N_3431,N_3162);
or U5153 (N_5153,N_2817,N_456);
or U5154 (N_5154,N_3257,N_4965);
and U5155 (N_5155,N_3533,N_2749);
nand U5156 (N_5156,N_1538,N_2610);
and U5157 (N_5157,N_403,N_3941);
or U5158 (N_5158,N_1343,N_3173);
xnor U5159 (N_5159,N_3823,N_846);
nor U5160 (N_5160,N_1512,N_4228);
nor U5161 (N_5161,N_3177,N_522);
or U5162 (N_5162,N_3435,N_428);
nor U5163 (N_5163,N_4440,N_4053);
nor U5164 (N_5164,N_1455,N_2869);
and U5165 (N_5165,N_1120,N_1599);
or U5166 (N_5166,N_1896,N_2159);
xor U5167 (N_5167,N_746,N_1137);
and U5168 (N_5168,N_3264,N_1656);
and U5169 (N_5169,N_1525,N_3408);
and U5170 (N_5170,N_4561,N_27);
nor U5171 (N_5171,N_3293,N_3790);
xnor U5172 (N_5172,N_579,N_4596);
or U5173 (N_5173,N_4859,N_2629);
nand U5174 (N_5174,N_2187,N_4473);
and U5175 (N_5175,N_4131,N_3096);
xnor U5176 (N_5176,N_1127,N_4461);
or U5177 (N_5177,N_142,N_3950);
nor U5178 (N_5178,N_346,N_3295);
nand U5179 (N_5179,N_359,N_4655);
xor U5180 (N_5180,N_580,N_4247);
xnor U5181 (N_5181,N_4124,N_1766);
nand U5182 (N_5182,N_4248,N_3349);
nor U5183 (N_5183,N_1218,N_2694);
nor U5184 (N_5184,N_3614,N_4046);
or U5185 (N_5185,N_4255,N_2586);
and U5186 (N_5186,N_2277,N_2172);
and U5187 (N_5187,N_3475,N_2168);
nor U5188 (N_5188,N_1915,N_4011);
xor U5189 (N_5189,N_3740,N_352);
or U5190 (N_5190,N_467,N_3406);
or U5191 (N_5191,N_2325,N_3317);
xor U5192 (N_5192,N_3751,N_3037);
xnor U5193 (N_5193,N_4721,N_458);
nand U5194 (N_5194,N_1135,N_1027);
xor U5195 (N_5195,N_2630,N_3901);
nand U5196 (N_5196,N_606,N_4460);
nand U5197 (N_5197,N_1505,N_2720);
nor U5198 (N_5198,N_2640,N_193);
and U5199 (N_5199,N_4780,N_1831);
nand U5200 (N_5200,N_2206,N_4093);
nand U5201 (N_5201,N_3968,N_2937);
nor U5202 (N_5202,N_4603,N_2446);
and U5203 (N_5203,N_1275,N_3984);
and U5204 (N_5204,N_3498,N_3015);
and U5205 (N_5205,N_388,N_4642);
and U5206 (N_5206,N_3862,N_280);
nor U5207 (N_5207,N_1049,N_4819);
or U5208 (N_5208,N_3384,N_2001);
and U5209 (N_5209,N_3514,N_4292);
nor U5210 (N_5210,N_3374,N_4197);
nor U5211 (N_5211,N_3057,N_3963);
xor U5212 (N_5212,N_2017,N_3214);
nor U5213 (N_5213,N_410,N_382);
nor U5214 (N_5214,N_3245,N_1160);
or U5215 (N_5215,N_4160,N_3501);
xor U5216 (N_5216,N_2409,N_3936);
and U5217 (N_5217,N_4411,N_2283);
xor U5218 (N_5218,N_1629,N_2761);
nor U5219 (N_5219,N_1100,N_1157);
nor U5220 (N_5220,N_4260,N_1841);
nor U5221 (N_5221,N_686,N_3551);
nand U5222 (N_5222,N_3750,N_1916);
or U5223 (N_5223,N_194,N_4572);
nor U5224 (N_5224,N_2522,N_3176);
xor U5225 (N_5225,N_608,N_804);
nor U5226 (N_5226,N_3929,N_1792);
nor U5227 (N_5227,N_161,N_345);
or U5228 (N_5228,N_3379,N_734);
nor U5229 (N_5229,N_584,N_3849);
nor U5230 (N_5230,N_1192,N_3283);
xor U5231 (N_5231,N_937,N_2684);
xor U5232 (N_5232,N_2200,N_1405);
and U5233 (N_5233,N_4645,N_2676);
nor U5234 (N_5234,N_709,N_4607);
or U5235 (N_5235,N_3532,N_4315);
nor U5236 (N_5236,N_1005,N_3538);
xnor U5237 (N_5237,N_1972,N_2580);
and U5238 (N_5238,N_3794,N_3454);
and U5239 (N_5239,N_1878,N_2774);
nor U5240 (N_5240,N_665,N_3035);
nand U5241 (N_5241,N_3604,N_1573);
or U5242 (N_5242,N_1159,N_4480);
and U5243 (N_5243,N_548,N_371);
or U5244 (N_5244,N_1130,N_2796);
or U5245 (N_5245,N_2686,N_1230);
nor U5246 (N_5246,N_2103,N_2445);
and U5247 (N_5247,N_3660,N_3912);
nand U5248 (N_5248,N_967,N_1450);
nor U5249 (N_5249,N_3806,N_4122);
and U5250 (N_5250,N_3847,N_1523);
xor U5251 (N_5251,N_3934,N_678);
nor U5252 (N_5252,N_79,N_1064);
xnor U5253 (N_5253,N_4786,N_214);
or U5254 (N_5254,N_1408,N_4841);
xnor U5255 (N_5255,N_943,N_2350);
nand U5256 (N_5256,N_4280,N_1063);
xor U5257 (N_5257,N_3548,N_2330);
nand U5258 (N_5258,N_4969,N_3016);
xor U5259 (N_5259,N_1634,N_823);
nor U5260 (N_5260,N_2666,N_396);
nand U5261 (N_5261,N_22,N_230);
xor U5262 (N_5262,N_1928,N_3420);
nor U5263 (N_5263,N_886,N_1035);
nand U5264 (N_5264,N_4271,N_1459);
xor U5265 (N_5265,N_1103,N_672);
and U5266 (N_5266,N_4731,N_4167);
xnor U5267 (N_5267,N_2695,N_1191);
nor U5268 (N_5268,N_925,N_240);
or U5269 (N_5269,N_2790,N_4798);
nor U5270 (N_5270,N_3736,N_2429);
nor U5271 (N_5271,N_1889,N_2153);
nand U5272 (N_5272,N_1199,N_3743);
xor U5273 (N_5273,N_234,N_3588);
nand U5274 (N_5274,N_3975,N_2015);
nor U5275 (N_5275,N_1395,N_2186);
nor U5276 (N_5276,N_3920,N_1215);
or U5277 (N_5277,N_2387,N_1383);
or U5278 (N_5278,N_2889,N_2956);
nor U5279 (N_5279,N_1332,N_3596);
nand U5280 (N_5280,N_2534,N_4787);
or U5281 (N_5281,N_1777,N_4697);
and U5282 (N_5282,N_3411,N_2107);
nand U5283 (N_5283,N_332,N_1641);
and U5284 (N_5284,N_3553,N_4481);
nand U5285 (N_5285,N_2764,N_1410);
or U5286 (N_5286,N_349,N_1549);
nand U5287 (N_5287,N_4904,N_3213);
and U5288 (N_5288,N_2497,N_4150);
nor U5289 (N_5289,N_2371,N_1194);
nand U5290 (N_5290,N_3643,N_4078);
nand U5291 (N_5291,N_3119,N_798);
or U5292 (N_5292,N_4188,N_4590);
nand U5293 (N_5293,N_3344,N_4365);
nand U5294 (N_5294,N_1779,N_589);
nor U5295 (N_5295,N_2932,N_3597);
nor U5296 (N_5296,N_91,N_2198);
nor U5297 (N_5297,N_4112,N_776);
or U5298 (N_5298,N_1361,N_4414);
or U5299 (N_5299,N_3185,N_3677);
xor U5300 (N_5300,N_3032,N_64);
nor U5301 (N_5301,N_3762,N_3517);
nor U5302 (N_5302,N_3415,N_143);
and U5303 (N_5303,N_4953,N_3271);
nor U5304 (N_5304,N_1935,N_3889);
and U5305 (N_5305,N_935,N_3873);
and U5306 (N_5306,N_575,N_1314);
xnor U5307 (N_5307,N_3097,N_3888);
nor U5308 (N_5308,N_1286,N_191);
xor U5309 (N_5309,N_2814,N_622);
nor U5310 (N_5310,N_527,N_631);
nor U5311 (N_5311,N_4483,N_3278);
xor U5312 (N_5312,N_4737,N_3133);
nand U5313 (N_5313,N_1280,N_4264);
or U5314 (N_5314,N_1113,N_4692);
nor U5315 (N_5315,N_3520,N_4477);
and U5316 (N_5316,N_4240,N_3606);
or U5317 (N_5317,N_2977,N_1430);
nor U5318 (N_5318,N_288,N_4109);
nand U5319 (N_5319,N_2303,N_2756);
and U5320 (N_5320,N_4984,N_598);
or U5321 (N_5321,N_594,N_2418);
xor U5322 (N_5322,N_335,N_4808);
xor U5323 (N_5323,N_3956,N_4304);
or U5324 (N_5324,N_867,N_3179);
nand U5325 (N_5325,N_1051,N_2847);
nor U5326 (N_5326,N_2507,N_4113);
nor U5327 (N_5327,N_1942,N_2816);
and U5328 (N_5328,N_2649,N_2955);
or U5329 (N_5329,N_730,N_1201);
and U5330 (N_5330,N_4129,N_2969);
nand U5331 (N_5331,N_3616,N_3369);
nand U5332 (N_5332,N_2261,N_566);
nand U5333 (N_5333,N_379,N_3252);
or U5334 (N_5334,N_4681,N_4845);
nor U5335 (N_5335,N_1729,N_2785);
and U5336 (N_5336,N_4991,N_648);
and U5337 (N_5337,N_2248,N_509);
and U5338 (N_5338,N_524,N_2748);
nor U5339 (N_5339,N_4284,N_1211);
or U5340 (N_5340,N_1461,N_1252);
xnor U5341 (N_5341,N_4742,N_1773);
and U5342 (N_5342,N_2727,N_3014);
xnor U5343 (N_5343,N_4043,N_4147);
or U5344 (N_5344,N_2288,N_1463);
or U5345 (N_5345,N_4059,N_911);
xnor U5346 (N_5346,N_482,N_4135);
or U5347 (N_5347,N_90,N_3870);
nor U5348 (N_5348,N_315,N_4382);
or U5349 (N_5349,N_226,N_2963);
and U5350 (N_5350,N_4183,N_3897);
or U5351 (N_5351,N_4784,N_511);
xnor U5352 (N_5352,N_3042,N_4544);
or U5353 (N_5353,N_3977,N_838);
or U5354 (N_5354,N_3957,N_4911);
nand U5355 (N_5355,N_3728,N_4955);
or U5356 (N_5356,N_3687,N_712);
or U5357 (N_5357,N_3263,N_1657);
nand U5358 (N_5358,N_2845,N_1339);
nor U5359 (N_5359,N_4106,N_146);
nand U5360 (N_5360,N_1301,N_1384);
or U5361 (N_5361,N_1188,N_2259);
or U5362 (N_5362,N_3226,N_701);
xnor U5363 (N_5363,N_414,N_2664);
or U5364 (N_5364,N_3443,N_4281);
xor U5365 (N_5365,N_742,N_1588);
xor U5366 (N_5366,N_2055,N_2608);
xnor U5367 (N_5367,N_2673,N_933);
xor U5368 (N_5368,N_1303,N_2972);
or U5369 (N_5369,N_2611,N_4138);
or U5370 (N_5370,N_3699,N_1699);
and U5371 (N_5371,N_2861,N_1091);
xor U5372 (N_5372,N_4234,N_1800);
xor U5373 (N_5373,N_3744,N_4728);
and U5374 (N_5374,N_860,N_180);
nor U5375 (N_5375,N_1711,N_334);
xnor U5376 (N_5376,N_2425,N_4425);
or U5377 (N_5377,N_708,N_1452);
or U5378 (N_5378,N_2912,N_1094);
nor U5379 (N_5379,N_2403,N_3166);
or U5380 (N_5380,N_3385,N_4105);
xnor U5381 (N_5381,N_400,N_3188);
nand U5382 (N_5382,N_33,N_4899);
nand U5383 (N_5383,N_3364,N_319);
nor U5384 (N_5384,N_4273,N_3457);
or U5385 (N_5385,N_3913,N_2269);
nor U5386 (N_5386,N_630,N_430);
nand U5387 (N_5387,N_3253,N_3433);
xnor U5388 (N_5388,N_3544,N_3468);
xnor U5389 (N_5389,N_4039,N_790);
xor U5390 (N_5390,N_1373,N_3495);
nor U5391 (N_5391,N_4988,N_115);
nand U5392 (N_5392,N_1241,N_3426);
or U5393 (N_5393,N_2381,N_1962);
nand U5394 (N_5394,N_3640,N_3703);
nor U5395 (N_5395,N_2892,N_3020);
or U5396 (N_5396,N_1429,N_731);
or U5397 (N_5397,N_402,N_1036);
and U5398 (N_5398,N_107,N_1555);
or U5399 (N_5399,N_1631,N_2014);
nand U5400 (N_5400,N_2344,N_3315);
and U5401 (N_5401,N_131,N_4755);
nor U5402 (N_5402,N_2800,N_4027);
nand U5403 (N_5403,N_3361,N_2512);
and U5404 (N_5404,N_3600,N_1835);
or U5405 (N_5405,N_3895,N_1423);
or U5406 (N_5406,N_2115,N_2718);
nor U5407 (N_5407,N_390,N_1364);
or U5408 (N_5408,N_3880,N_917);
nand U5409 (N_5409,N_3954,N_29);
and U5410 (N_5410,N_4221,N_781);
and U5411 (N_5411,N_2906,N_2383);
xor U5412 (N_5412,N_2506,N_1017);
nand U5413 (N_5413,N_1226,N_2059);
nand U5414 (N_5414,N_761,N_1012);
nand U5415 (N_5415,N_1697,N_3146);
and U5416 (N_5416,N_4996,N_615);
xnor U5417 (N_5417,N_2566,N_3926);
or U5418 (N_5418,N_1872,N_2472);
or U5419 (N_5419,N_4372,N_4490);
nor U5420 (N_5420,N_1400,N_4371);
xor U5421 (N_5421,N_801,N_374);
nor U5422 (N_5422,N_3741,N_4727);
xor U5423 (N_5423,N_657,N_2672);
and U5424 (N_5424,N_3769,N_1347);
or U5425 (N_5425,N_3294,N_3650);
or U5426 (N_5426,N_2165,N_2890);
nor U5427 (N_5427,N_3464,N_4530);
or U5428 (N_5428,N_4517,N_329);
and U5429 (N_5429,N_4564,N_3324);
nand U5430 (N_5430,N_223,N_2599);
or U5431 (N_5431,N_1238,N_1565);
or U5432 (N_5432,N_195,N_4045);
and U5433 (N_5433,N_4734,N_4606);
and U5434 (N_5434,N_2891,N_1427);
xnor U5435 (N_5435,N_4455,N_4957);
and U5436 (N_5436,N_1184,N_1290);
xor U5437 (N_5437,N_4503,N_2980);
or U5438 (N_5438,N_3370,N_3565);
xnor U5439 (N_5439,N_775,N_1170);
nor U5440 (N_5440,N_4522,N_45);
xnor U5441 (N_5441,N_2505,N_1311);
and U5442 (N_5442,N_2359,N_406);
nand U5443 (N_5443,N_897,N_92);
or U5444 (N_5444,N_3507,N_2757);
or U5445 (N_5445,N_4512,N_4349);
nand U5446 (N_5446,N_4615,N_1070);
or U5447 (N_5447,N_825,N_874);
and U5448 (N_5448,N_4774,N_499);
xnor U5449 (N_5449,N_416,N_956);
and U5450 (N_5450,N_4800,N_1377);
xnor U5451 (N_5451,N_4206,N_1611);
and U5452 (N_5452,N_1289,N_2380);
nand U5453 (N_5453,N_2404,N_3357);
or U5454 (N_5454,N_4827,N_2602);
nor U5455 (N_5455,N_1863,N_85);
nor U5456 (N_5456,N_2934,N_2355);
nor U5457 (N_5457,N_2366,N_2714);
nor U5458 (N_5458,N_2293,N_1501);
or U5459 (N_5459,N_3208,N_256);
and U5460 (N_5460,N_2682,N_1195);
xnor U5461 (N_5461,N_2529,N_472);
and U5462 (N_5462,N_116,N_1269);
and U5463 (N_5463,N_2591,N_695);
nand U5464 (N_5464,N_2287,N_1456);
and U5465 (N_5465,N_2074,N_2595);
xor U5466 (N_5466,N_4752,N_4286);
or U5467 (N_5467,N_4019,N_560);
xor U5468 (N_5468,N_3101,N_1076);
and U5469 (N_5469,N_4708,N_818);
and U5470 (N_5470,N_1689,N_3612);
and U5471 (N_5471,N_412,N_4350);
and U5472 (N_5472,N_4758,N_1851);
or U5473 (N_5473,N_3389,N_1316);
xor U5474 (N_5474,N_2289,N_2848);
nand U5475 (N_5475,N_370,N_903);
nor U5476 (N_5476,N_3046,N_2585);
nor U5477 (N_5477,N_4209,N_3022);
nand U5478 (N_5478,N_3256,N_1407);
nor U5479 (N_5479,N_433,N_504);
or U5480 (N_5480,N_3159,N_3512);
or U5481 (N_5481,N_3853,N_3107);
xnor U5482 (N_5482,N_2473,N_4501);
or U5483 (N_5483,N_4432,N_2964);
nor U5484 (N_5484,N_1710,N_2812);
xnor U5485 (N_5485,N_3203,N_893);
nor U5486 (N_5486,N_13,N_3777);
nand U5487 (N_5487,N_550,N_2307);
nor U5488 (N_5488,N_1999,N_4532);
and U5489 (N_5489,N_23,N_354);
and U5490 (N_5490,N_4328,N_3094);
nor U5491 (N_5491,N_4220,N_171);
xnor U5492 (N_5492,N_4981,N_2923);
and U5493 (N_5493,N_3391,N_568);
nor U5494 (N_5494,N_126,N_4058);
or U5495 (N_5495,N_94,N_4975);
and U5496 (N_5496,N_970,N_3919);
nand U5497 (N_5497,N_1894,N_3224);
and U5498 (N_5498,N_2438,N_4182);
xnor U5499 (N_5499,N_3590,N_2528);
and U5500 (N_5500,N_3137,N_2851);
xor U5501 (N_5501,N_2143,N_2603);
nand U5502 (N_5502,N_496,N_977);
nor U5503 (N_5503,N_4811,N_1925);
xnor U5504 (N_5504,N_1023,N_724);
and U5505 (N_5505,N_2138,N_1494);
and U5506 (N_5506,N_4041,N_1379);
xor U5507 (N_5507,N_4851,N_1265);
xor U5508 (N_5508,N_4066,N_4128);
xor U5509 (N_5509,N_4210,N_1980);
nor U5510 (N_5510,N_1664,N_2571);
nand U5511 (N_5511,N_1059,N_3816);
xnor U5512 (N_5512,N_172,N_1818);
or U5513 (N_5513,N_4623,N_3326);
xor U5514 (N_5514,N_1946,N_4756);
and U5515 (N_5515,N_340,N_1575);
nor U5516 (N_5516,N_1598,N_3078);
and U5517 (N_5517,N_4060,N_4224);
xor U5518 (N_5518,N_2635,N_4137);
nor U5519 (N_5519,N_4789,N_3865);
nor U5520 (N_5520,N_3136,N_2950);
and U5521 (N_5521,N_3795,N_1979);
xor U5522 (N_5522,N_4962,N_880);
and U5523 (N_5523,N_2146,N_857);
nand U5524 (N_5524,N_1852,N_2876);
xnor U5525 (N_5525,N_2141,N_1969);
nor U5526 (N_5526,N_3858,N_1352);
nor U5527 (N_5527,N_294,N_1510);
nor U5528 (N_5528,N_3585,N_768);
nor U5529 (N_5529,N_4239,N_780);
nor U5530 (N_5530,N_3439,N_258);
xor U5531 (N_5531,N_623,N_2336);
nand U5532 (N_5532,N_2444,N_2214);
nor U5533 (N_5533,N_305,N_2877);
xnor U5534 (N_5534,N_4960,N_2706);
nand U5535 (N_5535,N_4404,N_2885);
and U5536 (N_5536,N_4861,N_4064);
or U5537 (N_5537,N_624,N_245);
and U5538 (N_5538,N_2967,N_4608);
or U5539 (N_5539,N_581,N_2886);
xor U5540 (N_5540,N_3153,N_206);
and U5541 (N_5541,N_1660,N_3194);
and U5542 (N_5542,N_1209,N_2940);
nand U5543 (N_5543,N_531,N_607);
nand U5544 (N_5544,N_3698,N_3070);
and U5545 (N_5545,N_760,N_4308);
or U5546 (N_5546,N_170,N_4486);
xnor U5547 (N_5547,N_3639,N_2519);
nand U5548 (N_5548,N_974,N_4511);
and U5549 (N_5549,N_851,N_660);
xnor U5550 (N_5550,N_4339,N_2559);
or U5551 (N_5551,N_3802,N_2597);
or U5552 (N_5552,N_1471,N_2554);
and U5553 (N_5553,N_87,N_3407);
nor U5554 (N_5554,N_4747,N_3392);
and U5555 (N_5555,N_3727,N_2266);
nand U5556 (N_5556,N_3440,N_3198);
nand U5557 (N_5557,N_2834,N_1278);
and U5558 (N_5558,N_2925,N_3692);
or U5559 (N_5559,N_2826,N_461);
or U5560 (N_5560,N_2063,N_3222);
xnor U5561 (N_5561,N_3098,N_931);
or U5562 (N_5562,N_4997,N_4466);
nor U5563 (N_5563,N_4256,N_1553);
nand U5564 (N_5564,N_1257,N_610);
xor U5565 (N_5565,N_3363,N_74);
nand U5566 (N_5566,N_1654,N_398);
nor U5567 (N_5567,N_997,N_2652);
nor U5568 (N_5568,N_4044,N_3223);
nor U5569 (N_5569,N_1623,N_4246);
xnor U5570 (N_5570,N_188,N_2797);
xor U5571 (N_5571,N_1092,N_1391);
nand U5572 (N_5572,N_2846,N_3000);
xor U5573 (N_5573,N_132,N_2155);
nand U5574 (N_5574,N_1758,N_4146);
nand U5575 (N_5575,N_2057,N_4008);
nand U5576 (N_5576,N_2045,N_3864);
and U5577 (N_5577,N_3810,N_308);
xnor U5578 (N_5578,N_4162,N_2637);
nor U5579 (N_5579,N_1534,N_3309);
or U5580 (N_5580,N_3601,N_3958);
nand U5581 (N_5581,N_1328,N_145);
and U5582 (N_5582,N_3300,N_1105);
and U5583 (N_5583,N_4433,N_4844);
or U5584 (N_5584,N_2741,N_521);
xnor U5585 (N_5585,N_1374,N_2058);
nand U5586 (N_5586,N_462,N_4971);
xnor U5587 (N_5587,N_4472,N_387);
or U5588 (N_5588,N_4661,N_4175);
nor U5589 (N_5589,N_1843,N_592);
nor U5590 (N_5590,N_4482,N_676);
or U5591 (N_5591,N_4860,N_4306);
nand U5592 (N_5592,N_3908,N_3441);
nand U5593 (N_5593,N_3267,N_2803);
or U5594 (N_5594,N_1437,N_4435);
and U5595 (N_5595,N_813,N_2421);
nand U5596 (N_5596,N_2859,N_3997);
or U5597 (N_5597,N_3019,N_1780);
nor U5598 (N_5598,N_1725,N_4848);
nor U5599 (N_5599,N_3716,N_67);
xnor U5600 (N_5600,N_1670,N_399);
nand U5601 (N_5601,N_4682,N_395);
xor U5602 (N_5602,N_975,N_3132);
xnor U5603 (N_5603,N_1021,N_418);
and U5604 (N_5604,N_3262,N_3400);
nor U5605 (N_5605,N_1073,N_4812);
nand U5606 (N_5606,N_4999,N_644);
nor U5607 (N_5607,N_4071,N_3233);
nand U5608 (N_5608,N_2495,N_4513);
nand U5609 (N_5609,N_1321,N_1431);
and U5610 (N_5610,N_1834,N_1740);
nand U5611 (N_5611,N_135,N_2075);
or U5612 (N_5612,N_2818,N_291);
nor U5613 (N_5613,N_1169,N_1771);
nor U5614 (N_5614,N_889,N_4913);
or U5615 (N_5615,N_4395,N_77);
xor U5616 (N_5616,N_1585,N_2291);
xnor U5617 (N_5617,N_4985,N_1614);
xnor U5618 (N_5618,N_755,N_4267);
or U5619 (N_5619,N_3319,N_481);
nand U5620 (N_5620,N_208,N_2110);
and U5621 (N_5621,N_3760,N_4526);
xnor U5622 (N_5622,N_179,N_2679);
nand U5623 (N_5623,N_4676,N_4002);
and U5624 (N_5624,N_2084,N_3735);
nand U5625 (N_5625,N_4588,N_2032);
nand U5626 (N_5626,N_357,N_246);
xnor U5627 (N_5627,N_4342,N_3713);
or U5628 (N_5628,N_1223,N_3474);
nor U5629 (N_5629,N_3819,N_3249);
or U5630 (N_5630,N_3061,N_3684);
or U5631 (N_5631,N_949,N_4417);
and U5632 (N_5632,N_276,N_2907);
and U5633 (N_5633,N_3519,N_4939);
and U5634 (N_5634,N_3279,N_4278);
and U5635 (N_5635,N_3757,N_1376);
nand U5636 (N_5636,N_1306,N_3054);
xnor U5637 (N_5637,N_2641,N_4456);
xor U5638 (N_5638,N_2651,N_2726);
nand U5639 (N_5639,N_2911,N_2843);
nor U5640 (N_5640,N_1187,N_1607);
xor U5641 (N_5641,N_122,N_3982);
and U5642 (N_5642,N_128,N_235);
xor U5643 (N_5643,N_1068,N_3602);
nor U5644 (N_5644,N_1462,N_1602);
nand U5645 (N_5645,N_4098,N_1262);
xnor U5646 (N_5646,N_2126,N_3050);
xor U5647 (N_5647,N_544,N_4452);
nor U5648 (N_5648,N_1380,N_3781);
xnor U5649 (N_5649,N_1006,N_2807);
xor U5650 (N_5650,N_2431,N_4566);
nor U5651 (N_5651,N_3155,N_4302);
xnor U5652 (N_5652,N_2267,N_3033);
nor U5653 (N_5653,N_4702,N_268);
nor U5654 (N_5654,N_3526,N_2477);
nand U5655 (N_5655,N_2463,N_2677);
and U5656 (N_5656,N_4592,N_1719);
or U5657 (N_5657,N_3290,N_1433);
or U5658 (N_5658,N_3485,N_3093);
nand U5659 (N_5659,N_1963,N_4186);
nor U5660 (N_5660,N_564,N_3924);
and U5661 (N_5661,N_1090,N_3946);
nor U5662 (N_5662,N_2025,N_4386);
nand U5663 (N_5663,N_839,N_266);
or U5664 (N_5664,N_1887,N_740);
nor U5665 (N_5665,N_2406,N_510);
and U5666 (N_5666,N_4518,N_3649);
nor U5667 (N_5667,N_585,N_1752);
nor U5668 (N_5668,N_212,N_3486);
and U5669 (N_5669,N_487,N_1869);
xnor U5670 (N_5670,N_3644,N_2135);
or U5671 (N_5671,N_2361,N_1502);
xnor U5672 (N_5672,N_209,N_1504);
nand U5673 (N_5673,N_1814,N_3782);
nand U5674 (N_5674,N_4401,N_3998);
xor U5675 (N_5675,N_4901,N_4403);
xor U5676 (N_5676,N_1520,N_2222);
nor U5677 (N_5677,N_1388,N_707);
nor U5678 (N_5678,N_697,N_4717);
or U5679 (N_5679,N_1865,N_1082);
or U5680 (N_5680,N_4858,N_1691);
xnor U5681 (N_5681,N_1990,N_841);
or U5682 (N_5682,N_3993,N_2745);
xnor U5683 (N_5683,N_2013,N_793);
nand U5684 (N_5684,N_3797,N_899);
xor U5685 (N_5685,N_3282,N_2824);
nor U5686 (N_5686,N_3560,N_2631);
and U5687 (N_5687,N_4354,N_4886);
nor U5688 (N_5688,N_4193,N_3321);
nor U5689 (N_5689,N_2548,N_1948);
nor U5690 (N_5690,N_2272,N_2578);
xnor U5691 (N_5691,N_2503,N_1369);
or U5692 (N_5692,N_3482,N_233);
nand U5693 (N_5693,N_532,N_603);
nor U5694 (N_5694,N_1351,N_4749);
nand U5695 (N_5695,N_4882,N_73);
or U5696 (N_5696,N_2962,N_1348);
or U5697 (N_5697,N_3272,N_103);
xnor U5698 (N_5698,N_4601,N_3659);
and U5699 (N_5699,N_3671,N_1007);
nand U5700 (N_5700,N_2621,N_1465);
and U5701 (N_5701,N_4289,N_4156);
nand U5702 (N_5702,N_2113,N_2193);
nor U5703 (N_5703,N_2550,N_3978);
and U5704 (N_5704,N_2878,N_2356);
or U5705 (N_5705,N_4973,N_4555);
xnor U5706 (N_5706,N_1675,N_426);
and U5707 (N_5707,N_3437,N_407);
and U5708 (N_5708,N_2401,N_3428);
and U5709 (N_5709,N_432,N_4683);
xor U5710 (N_5710,N_512,N_4930);
or U5711 (N_5711,N_4200,N_2368);
nor U5712 (N_5712,N_2656,N_1349);
or U5713 (N_5713,N_4318,N_2958);
and U5714 (N_5714,N_4976,N_4543);
nand U5715 (N_5715,N_2620,N_2661);
xnor U5716 (N_5716,N_1734,N_2732);
nand U5717 (N_5717,N_1325,N_2688);
and U5718 (N_5718,N_1608,N_3678);
or U5719 (N_5719,N_1338,N_2199);
or U5720 (N_5720,N_4856,N_284);
xnor U5721 (N_5721,N_12,N_1406);
nor U5722 (N_5722,N_2420,N_2536);
nor U5723 (N_5723,N_2100,N_2211);
xor U5724 (N_5724,N_2052,N_1883);
xnor U5725 (N_5725,N_2194,N_3058);
nand U5726 (N_5726,N_4463,N_2150);
or U5727 (N_5727,N_2540,N_1676);
nor U5728 (N_5728,N_4000,N_2879);
nand U5729 (N_5729,N_494,N_983);
or U5730 (N_5730,N_3742,N_269);
or U5731 (N_5731,N_2701,N_1330);
nand U5732 (N_5732,N_692,N_990);
nor U5733 (N_5733,N_3108,N_1983);
or U5734 (N_5734,N_2095,N_4716);
xor U5735 (N_5735,N_1989,N_4136);
or U5736 (N_5736,N_1336,N_4871);
xnor U5737 (N_5737,N_2166,N_2315);
or U5738 (N_5738,N_1360,N_2183);
nand U5739 (N_5739,N_3308,N_1245);
nor U5740 (N_5740,N_4179,N_4750);
xor U5741 (N_5741,N_836,N_4118);
and U5742 (N_5742,N_2898,N_1649);
nor U5743 (N_5743,N_4635,N_3336);
or U5744 (N_5744,N_2481,N_3658);
or U5745 (N_5745,N_4529,N_1626);
nand U5746 (N_5746,N_4275,N_3442);
nand U5747 (N_5747,N_1819,N_2713);
xor U5748 (N_5748,N_4408,N_1454);
or U5749 (N_5749,N_2866,N_4163);
nand U5750 (N_5750,N_3,N_300);
nor U5751 (N_5751,N_200,N_2128);
xor U5752 (N_5752,N_2062,N_3818);
xnor U5753 (N_5753,N_4688,N_908);
nor U5754 (N_5754,N_1850,N_3259);
xor U5755 (N_5755,N_373,N_337);
nand U5756 (N_5756,N_939,N_2167);
xnor U5757 (N_5757,N_2488,N_1627);
and U5758 (N_5758,N_4317,N_323);
nor U5759 (N_5759,N_1778,N_2842);
nor U5760 (N_5760,N_4902,N_3547);
or U5761 (N_5761,N_201,N_3573);
and U5762 (N_5762,N_2462,N_1732);
and U5763 (N_5763,N_4549,N_4542);
xor U5764 (N_5764,N_3562,N_3511);
nor U5765 (N_5765,N_3691,N_4020);
or U5766 (N_5766,N_2479,N_1517);
nor U5767 (N_5767,N_1366,N_3053);
nand U5768 (N_5768,N_1272,N_4468);
or U5769 (N_5769,N_3550,N_3068);
or U5770 (N_5770,N_3065,N_417);
xor U5771 (N_5771,N_4785,N_2489);
nand U5772 (N_5772,N_4888,N_577);
and U5773 (N_5773,N_1624,N_1524);
nand U5774 (N_5774,N_984,N_3930);
and U5775 (N_5775,N_2709,N_324);
or U5776 (N_5776,N_4944,N_613);
and U5777 (N_5777,N_227,N_3200);
xnor U5778 (N_5778,N_4890,N_1848);
nor U5779 (N_5779,N_2270,N_491);
nor U5780 (N_5780,N_2320,N_1222);
xnor U5781 (N_5781,N_259,N_155);
or U5782 (N_5782,N_32,N_224);
and U5783 (N_5783,N_3557,N_3884);
nor U5784 (N_5784,N_4660,N_3911);
nor U5785 (N_5785,N_111,N_2788);
and U5786 (N_5786,N_653,N_3580);
nand U5787 (N_5787,N_4092,N_1702);
or U5788 (N_5788,N_2051,N_1274);
or U5789 (N_5789,N_2567,N_1253);
or U5790 (N_5790,N_2587,N_3527);
and U5791 (N_5791,N_3933,N_1596);
xnor U5792 (N_5792,N_4180,N_1612);
nand U5793 (N_5793,N_4829,N_869);
and U5794 (N_5794,N_3524,N_650);
nand U5795 (N_5795,N_1256,N_2098);
and U5796 (N_5796,N_4583,N_1922);
and U5797 (N_5797,N_4450,N_1583);
nor U5798 (N_5798,N_2304,N_167);
nor U5799 (N_5799,N_3006,N_2377);
nor U5800 (N_5800,N_513,N_721);
and U5801 (N_5801,N_484,N_2612);
nor U5802 (N_5802,N_2273,N_3109);
nor U5803 (N_5803,N_2451,N_4753);
or U5804 (N_5804,N_4216,N_39);
and U5805 (N_5805,N_4476,N_3592);
nor U5806 (N_5806,N_4791,N_542);
and U5807 (N_5807,N_4770,N_3756);
nor U5808 (N_5808,N_1912,N_2773);
nor U5809 (N_5809,N_2991,N_1426);
nand U5810 (N_5810,N_4236,N_1647);
or U5811 (N_5811,N_1926,N_4145);
nor U5812 (N_5812,N_2047,N_4624);
xnor U5813 (N_5813,N_4983,N_2657);
and U5814 (N_5814,N_4434,N_3491);
xor U5815 (N_5815,N_3480,N_3071);
or U5816 (N_5816,N_1001,N_4504);
nor U5817 (N_5817,N_2201,N_4320);
or U5818 (N_5818,N_363,N_1938);
xor U5819 (N_5819,N_4067,N_3123);
nand U5820 (N_5820,N_2504,N_2655);
xnor U5821 (N_5821,N_4394,N_18);
or U5822 (N_5822,N_2929,N_668);
and U5823 (N_5823,N_4712,N_4534);
and U5824 (N_5824,N_4571,N_876);
and U5825 (N_5825,N_979,N_3629);
nor U5826 (N_5826,N_2813,N_204);
or U5827 (N_5827,N_728,N_4288);
and U5828 (N_5828,N_3241,N_2258);
nand U5829 (N_5829,N_1993,N_164);
nor U5830 (N_5830,N_1554,N_4843);
xnor U5831 (N_5831,N_1992,N_654);
and U5832 (N_5832,N_3455,N_3341);
or U5833 (N_5833,N_3617,N_518);
xor U5834 (N_5834,N_1205,N_198);
nor U5835 (N_5835,N_127,N_2968);
and U5836 (N_5836,N_1809,N_3673);
or U5837 (N_5837,N_3619,N_1957);
or U5838 (N_5838,N_4012,N_2888);
nor U5839 (N_5839,N_328,N_1981);
and U5840 (N_5840,N_316,N_4126);
and U5841 (N_5841,N_1345,N_279);
nand U5842 (N_5842,N_4368,N_2875);
or U5843 (N_5843,N_2485,N_553);
nand U5844 (N_5844,N_913,N_556);
nand U5845 (N_5845,N_1134,N_4667);
nand U5846 (N_5846,N_4413,N_3383);
and U5847 (N_5847,N_2260,N_3377);
nand U5848 (N_5848,N_2190,N_4914);
nor U5849 (N_5849,N_110,N_1741);
nor U5850 (N_5850,N_1633,N_1885);
xnor U5851 (N_5851,N_1389,N_434);
or U5852 (N_5852,N_250,N_2124);
nor U5853 (N_5853,N_555,N_3325);
nor U5854 (N_5854,N_2264,N_4940);
nand U5855 (N_5855,N_546,N_3100);
nand U5856 (N_5856,N_4191,N_2265);
or U5857 (N_5857,N_1891,N_4235);
or U5858 (N_5858,N_1350,N_1976);
nor U5859 (N_5859,N_1684,N_2499);
nand U5860 (N_5860,N_4084,N_1491);
or U5861 (N_5861,N_4277,N_3126);
and U5862 (N_5862,N_4334,N_4835);
xor U5863 (N_5863,N_3871,N_2461);
xor U5864 (N_5864,N_1606,N_2563);
nor U5865 (N_5865,N_3029,N_3572);
xnor U5866 (N_5866,N_415,N_4775);
xor U5867 (N_5867,N_4585,N_2811);
or U5868 (N_5868,N_1305,N_2037);
xor U5869 (N_5869,N_1368,N_4912);
nor U5870 (N_5870,N_1415,N_4035);
xnor U5871 (N_5871,N_4420,N_3221);
and U5872 (N_5872,N_24,N_4628);
and U5873 (N_5873,N_3723,N_4076);
xor U5874 (N_5874,N_4510,N_2921);
nand U5875 (N_5875,N_3073,N_4771);
xor U5876 (N_5876,N_1069,N_3250);
xor U5877 (N_5877,N_4698,N_4778);
nor U5878 (N_5878,N_273,N_1297);
nor U5879 (N_5879,N_1582,N_1581);
xnor U5880 (N_5880,N_4563,N_2647);
and U5881 (N_5881,N_4241,N_4714);
and U5882 (N_5882,N_1717,N_2767);
nor U5883 (N_5883,N_3693,N_3002);
or U5884 (N_5884,N_4516,N_627);
nand U5885 (N_5885,N_1846,N_3332);
nor U5886 (N_5886,N_2897,N_4484);
or U5887 (N_5887,N_4325,N_3603);
nor U5888 (N_5888,N_3623,N_1712);
xnor U5889 (N_5889,N_4640,N_2884);
nor U5890 (N_5890,N_868,N_3266);
nor U5891 (N_5891,N_1178,N_3285);
nor U5892 (N_5892,N_2496,N_1066);
nor U5893 (N_5893,N_3064,N_2035);
and U5894 (N_5894,N_1445,N_1709);
and U5895 (N_5895,N_1716,N_4507);
and U5896 (N_5896,N_2232,N_154);
nor U5897 (N_5897,N_4884,N_56);
xnor U5898 (N_5898,N_4497,N_2823);
nor U5899 (N_5899,N_1414,N_3360);
or U5900 (N_5900,N_4554,N_4091);
nand U5901 (N_5901,N_2665,N_437);
nor U5902 (N_5902,N_3251,N_3207);
nor U5903 (N_5903,N_1567,N_1044);
nand U5904 (N_5904,N_123,N_1138);
nor U5905 (N_5905,N_93,N_2557);
and U5906 (N_5906,N_1378,N_2170);
xor U5907 (N_5907,N_2806,N_1556);
and U5908 (N_5908,N_2195,N_4222);
nor U5909 (N_5909,N_3092,N_2698);
xnor U5910 (N_5910,N_1307,N_3798);
and U5911 (N_5911,N_3780,N_479);
or U5912 (N_5912,N_3313,N_26);
nand U5913 (N_5913,N_3932,N_2142);
xor U5914 (N_5914,N_261,N_1665);
nand U5915 (N_5915,N_552,N_685);
and U5916 (N_5916,N_4978,N_878);
or U5917 (N_5917,N_3255,N_4231);
xnor U5918 (N_5918,N_166,N_176);
xnor U5919 (N_5919,N_4015,N_864);
xnor U5920 (N_5920,N_2960,N_1830);
nand U5921 (N_5921,N_1988,N_457);
nor U5922 (N_5922,N_3114,N_2178);
nand U5923 (N_5923,N_4772,N_1409);
xnor U5924 (N_5924,N_83,N_1796);
or U5925 (N_5925,N_2249,N_796);
and U5926 (N_5926,N_1866,N_1288);
nand U5927 (N_5927,N_3598,N_4905);
or U5928 (N_5928,N_392,N_3530);
xnor U5929 (N_5929,N_2041,N_2339);
and U5930 (N_5930,N_1467,N_3299);
nand U5931 (N_5931,N_855,N_2434);
xor U5932 (N_5932,N_778,N_2681);
and U5933 (N_5933,N_4704,N_4629);
nor U5934 (N_5934,N_3710,N_1768);
and U5935 (N_5935,N_3239,N_2601);
or U5936 (N_5936,N_762,N_700);
and U5937 (N_5937,N_549,N_1358);
nor U5938 (N_5938,N_1331,N_4010);
xnor U5939 (N_5939,N_2801,N_4117);
and U5940 (N_5940,N_1031,N_314);
xnor U5941 (N_5941,N_4272,N_2936);
and U5942 (N_5942,N_1826,N_4736);
nor U5943 (N_5943,N_1613,N_1832);
nor U5944 (N_5944,N_3838,N_2935);
nand U5945 (N_5945,N_3219,N_3082);
or U5946 (N_5946,N_2643,N_4796);
and U5947 (N_5947,N_2872,N_3348);
and U5948 (N_5948,N_1640,N_1497);
nand U5949 (N_5949,N_2516,N_1151);
nand U5950 (N_5950,N_362,N_4907);
nor U5951 (N_5951,N_2326,N_2023);
or U5952 (N_5952,N_1786,N_4568);
and U5953 (N_5953,N_4687,N_3834);
and U5954 (N_5954,N_1892,N_3306);
nor U5955 (N_5955,N_2369,N_4710);
nand U5956 (N_5956,N_3080,N_130);
or U5957 (N_5957,N_2004,N_1176);
or U5958 (N_5958,N_3555,N_3149);
or U5959 (N_5959,N_4725,N_4565);
xor U5960 (N_5960,N_3497,N_1216);
nor U5961 (N_5961,N_641,N_1533);
or U5962 (N_5962,N_480,N_1447);
nand U5963 (N_5963,N_265,N_3833);
nor U5964 (N_5964,N_2469,N_3388);
and U5965 (N_5965,N_1075,N_3236);
nor U5966 (N_5966,N_2831,N_3238);
nor U5967 (N_5967,N_4056,N_4016);
or U5968 (N_5968,N_2122,N_3509);
and U5969 (N_5969,N_139,N_218);
nor U5970 (N_5970,N_2156,N_1888);
and U5971 (N_5971,N_1698,N_42);
nand U5972 (N_5972,N_1793,N_3298);
nor U5973 (N_5973,N_4311,N_4846);
xnor U5974 (N_5974,N_4214,N_3863);
nand U5975 (N_5975,N_2614,N_2308);
or U5976 (N_5976,N_1340,N_4024);
xor U5977 (N_5977,N_3656,N_3031);
xnor U5978 (N_5978,N_3661,N_3183);
and U5979 (N_5979,N_3625,N_4332);
nand U5980 (N_5980,N_3610,N_3228);
and U5981 (N_5981,N_4369,N_4968);
xnor U5982 (N_5982,N_1546,N_722);
nand U5983 (N_5983,N_3883,N_726);
and U5984 (N_5984,N_3001,N_507);
xor U5985 (N_5985,N_1475,N_69);
xnor U5986 (N_5986,N_488,N_348);
xor U5987 (N_5987,N_44,N_1966);
nor U5988 (N_5988,N_1838,N_262);
nand U5989 (N_5989,N_4143,N_3124);
xor U5990 (N_5990,N_609,N_2317);
nand U5991 (N_5991,N_1868,N_601);
nand U5992 (N_5992,N_1353,N_2021);
nor U5993 (N_5993,N_894,N_3971);
or U5994 (N_5994,N_4047,N_236);
xnor U5995 (N_5995,N_3416,N_4815);
and U5996 (N_5996,N_4972,N_4094);
nand U5997 (N_5997,N_744,N_1956);
and U5998 (N_5998,N_4296,N_4679);
and U5999 (N_5999,N_2680,N_2101);
nor U6000 (N_6000,N_651,N_4873);
nand U6001 (N_6001,N_4213,N_2092);
and U6002 (N_6002,N_638,N_914);
nor U6003 (N_6003,N_4877,N_1011);
nor U6004 (N_6004,N_1478,N_3824);
or U6005 (N_6005,N_1087,N_149);
or U6006 (N_6006,N_1965,N_2453);
nor U6007 (N_6007,N_3765,N_3730);
nor U6008 (N_6008,N_4779,N_1337);
and U6009 (N_6009,N_965,N_1251);
nand U6010 (N_6010,N_916,N_4366);
nand U6011 (N_6011,N_3478,N_2396);
or U6012 (N_6012,N_1749,N_1917);
nand U6013 (N_6013,N_3593,N_2213);
and U6014 (N_6014,N_3607,N_1171);
and U6015 (N_6015,N_2835,N_347);
nor U6016 (N_6016,N_3296,N_4120);
nor U6017 (N_6017,N_3937,N_999);
xor U6018 (N_6018,N_634,N_62);
nand U6019 (N_6019,N_3900,N_4082);
or U6020 (N_6020,N_736,N_1971);
or U6021 (N_6021,N_2645,N_1065);
nor U6022 (N_6022,N_909,N_1735);
and U6023 (N_6023,N_702,N_3320);
and U6024 (N_6024,N_4204,N_2501);
nor U6025 (N_6025,N_492,N_3903);
or U6026 (N_6026,N_682,N_4918);
and U6027 (N_6027,N_4706,N_1849);
nand U6028 (N_6028,N_221,N_4760);
xnor U6029 (N_6029,N_3959,N_3423);
or U6030 (N_6030,N_2408,N_4164);
and U6031 (N_6031,N_1738,N_112);
or U6032 (N_6032,N_4880,N_3409);
xnor U6033 (N_6033,N_476,N_3039);
and U6034 (N_6034,N_4527,N_2079);
nor U6035 (N_6035,N_738,N_2589);
nand U6036 (N_6036,N_2568,N_1242);
xor U6037 (N_6037,N_966,N_2605);
or U6038 (N_6038,N_1239,N_215);
or U6039 (N_6039,N_4108,N_3459);
and U6040 (N_6040,N_4838,N_108);
and U6041 (N_6041,N_747,N_691);
nand U6042 (N_6042,N_792,N_232);
and U6043 (N_6043,N_1837,N_2050);
nand U6044 (N_6044,N_2648,N_331);
nand U6045 (N_6045,N_4424,N_1183);
and U6046 (N_6046,N_2760,N_1248);
or U6047 (N_6047,N_2060,N_995);
nand U6048 (N_6048,N_1899,N_765);
xor U6049 (N_6049,N_3525,N_4205);
or U6050 (N_6050,N_1279,N_4026);
xnor U6051 (N_6051,N_1692,N_8);
or U6052 (N_6052,N_1528,N_384);
or U6053 (N_6053,N_489,N_572);
nor U6054 (N_6054,N_4307,N_3196);
xnor U6055 (N_6055,N_783,N_1008);
nor U6056 (N_6056,N_698,N_4040);
xnor U6057 (N_6057,N_3269,N_4680);
nand U6058 (N_6058,N_503,N_3499);
or U6059 (N_6059,N_3793,N_1934);
xor U6060 (N_6060,N_3496,N_495);
and U6061 (N_6061,N_3734,N_794);
or U6062 (N_6062,N_2212,N_1671);
xor U6063 (N_6063,N_2737,N_1947);
and U6064 (N_6064,N_96,N_1560);
xnor U6065 (N_6065,N_2391,N_3542);
and U6066 (N_6066,N_3566,N_3131);
nand U6067 (N_6067,N_3534,N_443);
nand U6068 (N_6068,N_1568,N_578);
nand U6069 (N_6069,N_659,N_4356);
nor U6070 (N_6070,N_2573,N_3568);
or U6071 (N_6071,N_4065,N_2254);
and U6072 (N_6072,N_1398,N_2384);
and U6073 (N_6073,N_3558,N_2335);
nor U6074 (N_6074,N_4127,N_1532);
xnor U6075 (N_6075,N_3168,N_2600);
and U6076 (N_6076,N_2179,N_1442);
or U6077 (N_6077,N_4133,N_677);
nand U6078 (N_6078,N_313,N_808);
and U6079 (N_6079,N_1397,N_385);
nand U6080 (N_6080,N_535,N_1329);
nor U6081 (N_6081,N_1039,N_4282);
or U6082 (N_6082,N_3301,N_3747);
or U6083 (N_6083,N_2324,N_1203);
and U6084 (N_6084,N_4557,N_3048);
or U6085 (N_6085,N_486,N_2471);
and U6086 (N_6086,N_4735,N_4809);
nand U6087 (N_6087,N_4396,N_2360);
and U6088 (N_6088,N_1775,N_3909);
nor U6089 (N_6089,N_1206,N_3234);
and U6090 (N_6090,N_1959,N_3516);
nor U6091 (N_6091,N_2954,N_3445);
xnor U6092 (N_6092,N_687,N_4438);
nor U6093 (N_6093,N_140,N_4807);
or U6094 (N_6094,N_1055,N_2357);
nor U6095 (N_6095,N_3062,N_4936);
nand U6096 (N_6096,N_4375,N_3907);
xnor U6097 (N_6097,N_1385,N_1403);
nand U6098 (N_6098,N_2458,N_1718);
nor U6099 (N_6099,N_4358,N_4684);
nand U6100 (N_6100,N_1616,N_4322);
xor U6101 (N_6101,N_3630,N_1133);
nand U6102 (N_6102,N_1755,N_1106);
and U6103 (N_6103,N_1890,N_3697);
or U6104 (N_6104,N_2435,N_3796);
and U6105 (N_6105,N_941,N_3775);
xnor U6106 (N_6106,N_4169,N_1895);
and U6107 (N_6107,N_4367,N_4062);
nor U6108 (N_6108,N_4469,N_4699);
nor U6109 (N_6109,N_3567,N_16);
and U6110 (N_6110,N_3128,N_2638);
nor U6111 (N_6111,N_2109,N_3990);
and U6112 (N_6112,N_4101,N_1277);
nand U6113 (N_6113,N_1285,N_4351);
nor U6114 (N_6114,N_2999,N_1240);
or U6115 (N_6115,N_3003,N_1593);
nand U6116 (N_6116,N_4345,N_4048);
or U6117 (N_6117,N_4990,N_3302);
nor U6118 (N_6118,N_3962,N_3376);
nand U6119 (N_6119,N_1590,N_2087);
xor U6120 (N_6120,N_2944,N_3945);
nor U6121 (N_6121,N_2755,N_78);
nor U6122 (N_6122,N_1085,N_4379);
or U6123 (N_6123,N_1295,N_1970);
xor U6124 (N_6124,N_1308,N_4389);
or U6125 (N_6125,N_3394,N_2711);
nor U6126 (N_6126,N_4908,N_2294);
xnor U6127 (N_6127,N_2622,N_576);
nor U6128 (N_6128,N_378,N_4253);
xnor U6129 (N_6129,N_1842,N_1041);
nor U6130 (N_6130,N_4499,N_1453);
xor U6131 (N_6131,N_2633,N_928);
xnor U6132 (N_6132,N_2158,N_4547);
nor U6133 (N_6133,N_3886,N_3582);
nor U6134 (N_6134,N_4009,N_2370);
or U6135 (N_6135,N_2844,N_366);
nor U6136 (N_6136,N_1164,N_1141);
xnor U6137 (N_6137,N_3951,N_2674);
or U6138 (N_6138,N_4616,N_468);
nand U6139 (N_6139,N_3452,N_2426);
xor U6140 (N_6140,N_4740,N_3641);
nand U6141 (N_6141,N_1056,N_986);
nand U6142 (N_6142,N_4919,N_1667);
or U6143 (N_6143,N_1168,N_3334);
or U6144 (N_6144,N_4104,N_1098);
nand U6145 (N_6145,N_2414,N_4855);
nor U6146 (N_6146,N_4872,N_1355);
nor U6147 (N_6147,N_1714,N_1644);
or U6148 (N_6148,N_4090,N_244);
or U6149 (N_6149,N_3811,N_2837);
nor U6150 (N_6150,N_3135,N_2532);
xor U6151 (N_6151,N_88,N_1481);
xor U6152 (N_6152,N_3012,N_3701);
or U6153 (N_6153,N_3861,N_3809);
xor U6154 (N_6154,N_2464,N_3021);
xor U6155 (N_6155,N_3125,N_930);
nor U6156 (N_6156,N_4768,N_1236);
nor U6157 (N_6157,N_7,N_4745);
and U6158 (N_6158,N_4023,N_3085);
nor U6159 (N_6159,N_2691,N_807);
xnor U6160 (N_6160,N_3448,N_1513);
and U6161 (N_6161,N_3817,N_3571);
or U6162 (N_6162,N_3960,N_1165);
xnor U6163 (N_6163,N_1618,N_1186);
xnor U6164 (N_6164,N_2223,N_424);
and U6165 (N_6165,N_1950,N_3987);
nor U6166 (N_6166,N_153,N_1561);
xor U6167 (N_6167,N_455,N_4052);
xnor U6168 (N_6168,N_4038,N_47);
xnor U6169 (N_6169,N_2624,N_4100);
nor U6170 (N_6170,N_670,N_2604);
or U6171 (N_6171,N_1499,N_2518);
nand U6172 (N_6172,N_929,N_1259);
nor U6173 (N_6173,N_3353,N_4036);
and U6174 (N_6174,N_3633,N_640);
xnor U6175 (N_6175,N_538,N_2575);
and U6176 (N_6176,N_1084,N_4722);
and U6177 (N_6177,N_3632,N_2096);
and U6178 (N_6178,N_3187,N_2793);
and U6179 (N_6179,N_4553,N_1739);
nand U6180 (N_6180,N_475,N_1703);
or U6181 (N_6181,N_2524,N_2538);
and U6182 (N_6182,N_2349,N_3129);
or U6183 (N_6183,N_2234,N_3479);
nor U6184 (N_6184,N_985,N_1125);
xor U6185 (N_6185,N_1229,N_1189);
nor U6186 (N_6186,N_2729,N_2139);
or U6187 (N_6187,N_1529,N_473);
xnor U6188 (N_6188,N_2570,N_3402);
nor U6189 (N_6189,N_4834,N_1);
nand U6190 (N_6190,N_4903,N_2839);
and U6191 (N_6191,N_4158,N_625);
nand U6192 (N_6192,N_3351,N_3143);
nand U6193 (N_6193,N_1977,N_1172);
xnor U6194 (N_6194,N_4007,N_2077);
nand U6195 (N_6195,N_940,N_3502);
nand U6196 (N_6196,N_3004,N_2588);
xnor U6197 (N_6197,N_2225,N_3683);
nor U6198 (N_6198,N_1260,N_2564);
nand U6199 (N_6199,N_764,N_2692);
nand U6200 (N_6200,N_448,N_3925);
or U6201 (N_6201,N_219,N_2852);
and U6202 (N_6202,N_565,N_2989);
nand U6203 (N_6203,N_1822,N_4492);
xor U6204 (N_6204,N_2494,N_2002);
nand U6205 (N_6205,N_1669,N_921);
nor U6206 (N_6206,N_1335,N_737);
or U6207 (N_6207,N_4291,N_4925);
and U6208 (N_6208,N_3820,N_2850);
or U6209 (N_6209,N_2066,N_1217);
nor U6210 (N_6210,N_1500,N_2176);
nor U6211 (N_6211,N_2393,N_228);
xnor U6212 (N_6212,N_2993,N_3453);
nor U6213 (N_6213,N_3410,N_3680);
nor U6214 (N_6214,N_3776,N_2836);
and U6215 (N_6215,N_4701,N_4641);
or U6216 (N_6216,N_1761,N_2904);
xor U6217 (N_6217,N_3916,N_978);
xnor U6218 (N_6218,N_3654,N_4514);
or U6219 (N_6219,N_4935,N_3965);
nor U6220 (N_6220,N_1270,N_231);
nor U6221 (N_6221,N_4669,N_3034);
nor U6222 (N_6222,N_4887,N_177);
xnor U6223 (N_6223,N_3878,N_4943);
xor U6224 (N_6224,N_3882,N_1402);
or U6225 (N_6225,N_4528,N_4069);
xor U6226 (N_6226,N_1677,N_3460);
or U6227 (N_6227,N_1424,N_649);
and U6228 (N_6228,N_3724,N_1688);
and U6229 (N_6229,N_4451,N_3594);
or U6230 (N_6230,N_405,N_992);
xnor U6231 (N_6231,N_699,N_1276);
or U6232 (N_6232,N_973,N_788);
xnor U6233 (N_6233,N_3545,N_3312);
and U6234 (N_6234,N_4192,N_216);
xnor U6235 (N_6235,N_1781,N_2274);
nor U6236 (N_6236,N_2508,N_3867);
and U6237 (N_6237,N_4464,N_2617);
nor U6238 (N_6238,N_2162,N_1024);
xnor U6239 (N_6239,N_4258,N_2228);
and U6240 (N_6240,N_3876,N_4448);
xor U6241 (N_6241,N_4013,N_1435);
or U6242 (N_6242,N_3541,N_3307);
or U6243 (N_6243,N_1179,N_3028);
and U6244 (N_6244,N_611,N_4980);
and U6245 (N_6245,N_303,N_4226);
and U6246 (N_6246,N_104,N_2316);
nor U6247 (N_6247,N_463,N_2117);
nor U6248 (N_6248,N_4244,N_2208);
and U6249 (N_6249,N_1422,N_2752);
xnor U6250 (N_6250,N_2314,N_4268);
or U6251 (N_6251,N_1449,N_1666);
nor U6252 (N_6252,N_1721,N_4626);
xor U6253 (N_6253,N_680,N_1795);
and U6254 (N_6254,N_1967,N_3705);
and U6255 (N_6255,N_633,N_136);
nor U6256 (N_6256,N_302,N_1019);
or U6257 (N_6257,N_3801,N_3059);
or U6258 (N_6258,N_3881,N_3515);
nor U6259 (N_6259,N_1974,N_1762);
or U6260 (N_6260,N_3537,N_275);
xor U6261 (N_6261,N_3209,N_812);
or U6262 (N_6262,N_3041,N_2941);
or U6263 (N_6263,N_2626,N_1458);
nand U6264 (N_6264,N_49,N_2144);
nor U6265 (N_6265,N_4491,N_2916);
nand U6266 (N_6266,N_4347,N_3169);
and U6267 (N_6267,N_1680,N_2029);
xnor U6268 (N_6268,N_1110,N_1495);
nand U6269 (N_6269,N_1794,N_3803);
or U6270 (N_6270,N_1161,N_1296);
xnor U6271 (N_6271,N_3084,N_4195);
nor U6272 (N_6272,N_1961,N_2569);
or U6273 (N_6273,N_213,N_715);
xnor U6274 (N_6274,N_2331,N_3425);
nand U6275 (N_6275,N_4948,N_3017);
or U6276 (N_6276,N_4088,N_4276);
nor U6277 (N_6277,N_2354,N_4416);
nand U6278 (N_6278,N_1951,N_3007);
nand U6279 (N_6279,N_3647,N_3484);
xnor U6280 (N_6280,N_2992,N_1050);
xnor U6281 (N_6281,N_3825,N_2702);
and U6282 (N_6282,N_1493,N_547);
and U6283 (N_6283,N_3869,N_2901);
xnor U6284 (N_6284,N_3745,N_1678);
xnor U6285 (N_6285,N_184,N_2312);
nor U6286 (N_6286,N_2204,N_4085);
xor U6287 (N_6287,N_4673,N_2399);
nand U6288 (N_6288,N_3712,N_508);
or U6289 (N_6289,N_3670,N_2947);
nor U6290 (N_6290,N_902,N_4211);
xnor U6291 (N_6291,N_1404,N_1515);
and U6292 (N_6292,N_661,N_174);
or U6293 (N_6293,N_1115,N_4144);
nand U6294 (N_6294,N_4233,N_2207);
nand U6295 (N_6295,N_645,N_822);
nor U6296 (N_6296,N_1143,N_4243);
xnor U6297 (N_6297,N_252,N_2280);
nor U6298 (N_6298,N_4814,N_53);
nor U6299 (N_6299,N_4898,N_34);
or U6300 (N_6300,N_1700,N_25);
xor U6301 (N_6301,N_3855,N_113);
xor U6302 (N_6302,N_3346,N_2085);
nand U6303 (N_6303,N_723,N_1857);
nand U6304 (N_6304,N_2218,N_4054);
and U6305 (N_6305,N_4788,N_2644);
nand U6306 (N_6306,N_782,N_4249);
xnor U6307 (N_6307,N_4648,N_1362);
and U6308 (N_6308,N_2776,N_4335);
nor U6309 (N_6309,N_1359,N_3556);
and U6310 (N_6310,N_646,N_1025);
or U6311 (N_6311,N_1508,N_705);
nor U6312 (N_6312,N_1897,N_2215);
and U6313 (N_6313,N_4994,N_2543);
nand U6314 (N_6314,N_3779,N_4966);
or U6315 (N_6315,N_1009,N_2576);
and U6316 (N_6316,N_1592,N_1029);
nand U6317 (N_6317,N_2281,N_4142);
xor U6318 (N_6318,N_1998,N_4559);
xnor U6319 (N_6319,N_6,N_4773);
xnor U6320 (N_6320,N_3195,N_756);
nor U6321 (N_6321,N_4376,N_444);
nand U6322 (N_6322,N_770,N_4533);
nor U6323 (N_6323,N_2763,N_3167);
and U6324 (N_6324,N_4079,N_1914);
nor U6325 (N_6325,N_368,N_376);
or U6326 (N_6326,N_2572,N_1509);
nand U6327 (N_6327,N_919,N_1022);
nand U6328 (N_6328,N_1466,N_694);
nor U6329 (N_6329,N_1235,N_1145);
nor U6330 (N_6330,N_2310,N_541);
xor U6331 (N_6331,N_4373,N_1078);
nor U6332 (N_6332,N_3086,N_4618);
or U6333 (N_6333,N_2840,N_1298);
nand U6334 (N_6334,N_4739,N_1061);
nand U6335 (N_6335,N_3115,N_1727);
xor U6336 (N_6336,N_635,N_393);
nor U6337 (N_6337,N_3738,N_905);
or U6338 (N_6338,N_1342,N_186);
xnor U6339 (N_6339,N_454,N_2231);
and U6340 (N_6340,N_3211,N_1708);
xnor U6341 (N_6341,N_2487,N_4312);
nor U6342 (N_6342,N_4581,N_1921);
and U6343 (N_6343,N_1715,N_4001);
and U6344 (N_6344,N_1776,N_152);
and U6345 (N_6345,N_1326,N_4801);
nand U6346 (N_6346,N_3184,N_4072);
or U6347 (N_6347,N_1909,N_4397);
nor U6348 (N_6348,N_1060,N_2042);
nand U6349 (N_6349,N_106,N_2020);
or U6350 (N_6350,N_3340,N_1271);
or U6351 (N_6351,N_4300,N_830);
or U6352 (N_6352,N_4672,N_3421);
nor U6353 (N_6353,N_168,N_318);
xor U6354 (N_6354,N_70,N_211);
nor U6355 (N_6355,N_3696,N_1871);
nor U6356 (N_6356,N_1399,N_844);
nor U6357 (N_6357,N_4720,N_537);
and U6358 (N_6358,N_3850,N_3281);
and U6359 (N_6359,N_3044,N_4074);
nor U6360 (N_6360,N_4823,N_1232);
nand U6361 (N_6361,N_2243,N_2022);
nor U6362 (N_6362,N_1420,N_4560);
and U6363 (N_6363,N_2577,N_1101);
nor U6364 (N_6364,N_3899,N_1756);
nor U6365 (N_6365,N_4654,N_4970);
xnor U6366 (N_6366,N_1088,N_4285);
nor U6367 (N_6367,N_719,N_944);
and U6368 (N_6368,N_2038,N_4121);
nand U6369 (N_6369,N_3174,N_2476);
or U6370 (N_6370,N_1722,N_1536);
or U6371 (N_6371,N_203,N_2675);
and U6372 (N_6372,N_4398,N_690);
xor U6373 (N_6373,N_460,N_3893);
or U6374 (N_6374,N_3979,N_3690);
xor U6375 (N_6375,N_1030,N_4632);
xnor U6376 (N_6376,N_3800,N_4298);
and U6377 (N_6377,N_2509,N_2027);
nand U6378 (N_6378,N_3513,N_2995);
nand U6379 (N_6379,N_3988,N_1881);
nor U6380 (N_6380,N_1119,N_1291);
xor U6381 (N_6381,N_4508,N_4353);
xor U6382 (N_6382,N_2716,N_2952);
xnor U6383 (N_6383,N_2475,N_2104);
nor U6384 (N_6384,N_1185,N_3589);
nor U6385 (N_6385,N_1346,N_2899);
nand U6386 (N_6386,N_2539,N_3401);
or U6387 (N_6387,N_4767,N_3704);
and U6388 (N_6388,N_3231,N_3935);
or U6389 (N_6389,N_517,N_4757);
and U6390 (N_6390,N_3718,N_3761);
or U6391 (N_6391,N_3113,N_1591);
and U6392 (N_6392,N_3500,N_3754);
and U6393 (N_6393,N_2221,N_2130);
and U6394 (N_6394,N_4374,N_254);
and U6395 (N_6395,N_3679,N_3875);
or U6396 (N_6396,N_4402,N_1146);
or U6397 (N_6397,N_3075,N_1784);
or U6398 (N_6398,N_237,N_355);
nor U6399 (N_6399,N_3637,N_1020);
nand U6400 (N_6400,N_4409,N_3642);
nor U6401 (N_6401,N_2236,N_2491);
nand U6402 (N_6402,N_600,N_4593);
nor U6403 (N_6403,N_1907,N_554);
or U6404 (N_6404,N_1913,N_2994);
and U6405 (N_6405,N_2871,N_2699);
or U6406 (N_6406,N_1425,N_4713);
nor U6407 (N_6407,N_3122,N_3731);
or U6408 (N_6408,N_2181,N_1393);
nor U6409 (N_6409,N_4262,N_1898);
xor U6410 (N_6410,N_3615,N_2108);
nand U6411 (N_6411,N_2068,N_2808);
and U6412 (N_6412,N_516,N_3456);
xor U6413 (N_6413,N_1886,N_3413);
nor U6414 (N_6414,N_10,N_1018);
nand U6415 (N_6415,N_3318,N_2820);
and U6416 (N_6416,N_4157,N_4894);
nor U6417 (N_6417,N_4805,N_3561);
xnor U6418 (N_6418,N_1150,N_465);
nor U6419 (N_6419,N_2120,N_1002);
nor U6420 (N_6420,N_1707,N_2140);
nor U6421 (N_6421,N_4937,N_4207);
and U6422 (N_6422,N_689,N_4998);
nand U6423 (N_6423,N_3292,N_2743);
or U6424 (N_6424,N_2739,N_1652);
nand U6425 (N_6425,N_953,N_3577);
or U6426 (N_6426,N_4862,N_4830);
xnor U6427 (N_6427,N_745,N_3056);
and U6428 (N_6428,N_3199,N_4853);
xnor U6429 (N_6429,N_2668,N_4649);
xnor U6430 (N_6430,N_948,N_2016);
or U6431 (N_6431,N_1994,N_3578);
or U6432 (N_6432,N_827,N_2210);
or U6433 (N_6433,N_1124,N_514);
nor U6434 (N_6434,N_4506,N_4259);
and U6435 (N_6435,N_2114,N_637);
xnor U6436 (N_6436,N_885,N_1829);
nand U6437 (N_6437,N_1244,N_639);
nand U6438 (N_6438,N_409,N_1177);
nand U6439 (N_6439,N_1129,N_3877);
nand U6440 (N_6440,N_1097,N_2700);
nor U6441 (N_6441,N_257,N_1390);
nand U6442 (N_6442,N_1713,N_3225);
and U6443 (N_6443,N_1765,N_2245);
and U6444 (N_6444,N_1760,N_1790);
xnor U6445 (N_6445,N_4348,N_1317);
xor U6446 (N_6446,N_1570,N_4691);
and U6447 (N_6447,N_1109,N_267);
nand U6448 (N_6448,N_2933,N_1958);
xor U6449 (N_6449,N_1931,N_4227);
or U6450 (N_6450,N_4917,N_2152);
nor U6451 (N_6451,N_4850,N_2959);
nor U6452 (N_6452,N_2246,N_1267);
and U6453 (N_6453,N_274,N_3081);
and U6454 (N_6454,N_1638,N_2402);
nand U6455 (N_6455,N_771,N_3190);
nand U6456 (N_6456,N_3419,N_3047);
nand U6457 (N_6457,N_573,N_1604);
xor U6458 (N_6458,N_4776,N_4487);
and U6459 (N_6459,N_4964,N_173);
nor U6460 (N_6460,N_1263,N_4604);
xnor U6461 (N_6461,N_3689,N_4864);
xor U6462 (N_6462,N_3371,N_4575);
nor U6463 (N_6463,N_1949,N_474);
or U6464 (N_6464,N_3077,N_3189);
or U6465 (N_6465,N_4949,N_3635);
or U6466 (N_6466,N_3227,N_1531);
nand U6467 (N_6467,N_3117,N_4301);
xnor U6468 (N_6468,N_341,N_4134);
or U6469 (N_6469,N_497,N_2009);
nand U6470 (N_6470,N_54,N_2411);
nand U6471 (N_6471,N_4674,N_502);
or U6472 (N_6472,N_4609,N_2961);
or U6473 (N_6473,N_2520,N_629);
nor U6474 (N_6474,N_1884,N_1154);
or U6475 (N_6475,N_4795,N_19);
nor U6476 (N_6476,N_278,N_4653);
and U6477 (N_6477,N_2747,N_714);
or U6478 (N_6478,N_4087,N_4478);
nand U6479 (N_6479,N_1535,N_2457);
nor U6480 (N_6480,N_3620,N_2541);
nand U6481 (N_6481,N_1745,N_3613);
nand U6482 (N_6482,N_3655,N_4475);
xnor U6483 (N_6483,N_1731,N_3845);
or U6484 (N_6484,N_2299,N_1418);
or U6485 (N_6485,N_383,N_1662);
or U6486 (N_6486,N_647,N_3676);
nor U6487 (N_6487,N_2229,N_501);
or U6488 (N_6488,N_4878,N_4644);
nand U6489 (N_6489,N_2768,N_196);
xnor U6490 (N_6490,N_3424,N_1828);
and U6491 (N_6491,N_2828,N_4343);
or U6492 (N_6492,N_3872,N_847);
nor U6493 (N_6493,N_2298,N_4383);
and U6494 (N_6494,N_4580,N_2771);
xnor U6495 (N_6495,N_2549,N_2593);
and U6496 (N_6496,N_4381,N_3807);
or U6497 (N_6497,N_464,N_2433);
nand U6498 (N_6498,N_2775,N_2351);
nand U6499 (N_6499,N_377,N_918);
nor U6500 (N_6500,N_2772,N_3273);
xor U6501 (N_6501,N_3778,N_1757);
xor U6502 (N_6502,N_1464,N_286);
xnor U6503 (N_6503,N_2561,N_20);
nand U6504 (N_6504,N_2240,N_207);
and U6505 (N_6505,N_3812,N_58);
xnor U6506 (N_6506,N_105,N_1686);
xnor U6507 (N_6507,N_2685,N_2662);
nor U6508 (N_6508,N_834,N_4790);
or U6509 (N_6509,N_2758,N_1586);
xnor U6510 (N_6510,N_2285,N_2705);
nor U6511 (N_6511,N_4305,N_1619);
and U6512 (N_6512,N_500,N_3191);
xnor U6513 (N_6513,N_2669,N_2650);
or U6514 (N_6514,N_1566,N_1382);
nor U6515 (N_6515,N_1083,N_1724);
or U6516 (N_6516,N_4390,N_3905);
xor U6517 (N_6517,N_843,N_297);
xnor U6518 (N_6518,N_4357,N_5);
or U6519 (N_6519,N_1304,N_1747);
nand U6520 (N_6520,N_2751,N_2719);
and U6521 (N_6521,N_2574,N_3722);
and U6522 (N_6522,N_2428,N_4361);
nand U6523 (N_6523,N_4942,N_3458);
and U6524 (N_6524,N_4840,N_436);
and U6525 (N_6525,N_1572,N_1880);
or U6526 (N_6526,N_2046,N_4921);
nand U6527 (N_6527,N_1918,N_1387);
and U6528 (N_6528,N_1601,N_36);
or U6529 (N_6529,N_3914,N_3631);
or U6530 (N_6530,N_3994,N_3427);
nor U6531 (N_6531,N_4168,N_1312);
nor U6532 (N_6532,N_1486,N_1836);
xor U6533 (N_6533,N_1936,N_2531);
xor U6534 (N_6534,N_2607,N_394);
xor U6535 (N_6535,N_1750,N_3327);
and U6536 (N_6536,N_1744,N_2582);
xnor U6537 (N_6537,N_1121,N_2552);
xor U6538 (N_6538,N_4232,N_389);
nor U6539 (N_6539,N_187,N_299);
and U6540 (N_6540,N_3618,N_2432);
or U6541 (N_6541,N_3390,N_2192);
or U6542 (N_6542,N_2909,N_4196);
or U6543 (N_6543,N_4836,N_4531);
or U6544 (N_6544,N_1266,N_2667);
or U6545 (N_6545,N_2483,N_1043);
nor U6546 (N_6546,N_3763,N_1893);
xnor U6547 (N_6547,N_3316,N_3083);
nand U6548 (N_6548,N_895,N_2343);
xor U6549 (N_6549,N_4453,N_4229);
or U6550 (N_6550,N_4337,N_2424);
nor U6551 (N_6551,N_4399,N_632);
or U6552 (N_6552,N_994,N_1249);
xor U6553 (N_6553,N_4494,N_960);
and U6554 (N_6554,N_3280,N_4891);
nor U6555 (N_6555,N_3178,N_4867);
nor U6556 (N_6556,N_1428,N_1635);
nand U6557 (N_6557,N_2802,N_593);
xnor U6558 (N_6558,N_4173,N_1577);
and U6559 (N_6559,N_4658,N_4089);
nor U6560 (N_6560,N_3595,N_1472);
nand U6561 (N_6561,N_2920,N_4989);
nor U6562 (N_6562,N_4111,N_2226);
nand U6563 (N_6563,N_65,N_2598);
nand U6564 (N_6564,N_4159,N_1545);
xnor U6565 (N_6565,N_4266,N_3138);
nor U6566 (N_6566,N_1559,N_1576);
or U6567 (N_6567,N_2448,N_2660);
nand U6568 (N_6568,N_4584,N_4831);
xor U6569 (N_6569,N_4489,N_3784);
nand U6570 (N_6570,N_3104,N_2392);
and U6571 (N_6571,N_3980,N_4031);
xnor U6572 (N_6572,N_1323,N_753);
or U6573 (N_6573,N_595,N_4340);
and U6574 (N_6574,N_344,N_3989);
nor U6575 (N_6575,N_82,N_4832);
nand U6576 (N_6576,N_3333,N_656);
or U6577 (N_6577,N_1853,N_2118);
or U6578 (N_6578,N_3540,N_4077);
or U6579 (N_6579,N_1876,N_4257);
and U6580 (N_6580,N_1571,N_618);
or U6581 (N_6581,N_551,N_4651);
xor U6582 (N_6582,N_888,N_1370);
and U6583 (N_6583,N_4050,N_1605);
and U6584 (N_6584,N_3669,N_4362);
or U6585 (N_6585,N_669,N_3788);
xnor U6586 (N_6586,N_4187,N_1620);
and U6587 (N_6587,N_2945,N_2537);
nor U6588 (N_6588,N_4171,N_117);
xor U6589 (N_6589,N_3489,N_1810);
xor U6590 (N_6590,N_3986,N_2082);
nor U6591 (N_6591,N_2525,N_4909);
xor U6592 (N_6592,N_539,N_4746);
xnor U6593 (N_6593,N_3774,N_75);
or U6594 (N_6594,N_1128,N_453);
or U6595 (N_6595,N_2951,N_3121);
nand U6596 (N_6596,N_3362,N_4184);
xor U6597 (N_6597,N_3395,N_1730);
xnor U6598 (N_6598,N_3646,N_3922);
xnor U6599 (N_6599,N_4927,N_441);
or U6600 (N_6600,N_4309,N_4230);
xor U6601 (N_6601,N_2121,N_4619);
and U6602 (N_6602,N_2914,N_3412);
xor U6603 (N_6603,N_2227,N_3894);
or U6604 (N_6604,N_2822,N_4732);
nand U6605 (N_6605,N_4818,N_202);
nand U6606 (N_6606,N_2990,N_4443);
or U6607 (N_6607,N_1293,N_2492);
or U6608 (N_6608,N_4086,N_4004);
nand U6609 (N_6609,N_55,N_3622);
nor U6610 (N_6610,N_1483,N_3549);
nand U6611 (N_6611,N_2295,N_3210);
or U6612 (N_6612,N_1167,N_1228);
and U6613 (N_6613,N_1643,N_2099);
or U6614 (N_6614,N_1639,N_320);
xor U6615 (N_6615,N_693,N_1799);
xnor U6616 (N_6616,N_2949,N_3543);
and U6617 (N_6617,N_3171,N_298);
nor U6618 (N_6618,N_2882,N_2112);
or U6619 (N_6619,N_4931,N_3721);
and U6620 (N_6620,N_789,N_1439);
or U6621 (N_6621,N_84,N_1166);
or U6622 (N_6622,N_671,N_1820);
and U6623 (N_6623,N_4421,N_1600);
nor U6624 (N_6624,N_1960,N_4447);
nor U6625 (N_6625,N_2639,N_2853);
xor U6626 (N_6626,N_1743,N_452);
nand U6627 (N_6627,N_3928,N_1763);
xnor U6628 (N_6628,N_2407,N_1807);
xnor U6629 (N_6629,N_3848,N_2147);
nand U6630 (N_6630,N_121,N_4110);
nor U6631 (N_6631,N_3063,N_2498);
or U6632 (N_6632,N_4705,N_4338);
or U6633 (N_6633,N_1058,N_3386);
or U6634 (N_6634,N_4444,N_2365);
xor U6635 (N_6635,N_543,N_3240);
xnor U6636 (N_6636,N_2819,N_220);
or U6637 (N_6637,N_862,N_1053);
nor U6638 (N_6638,N_972,N_4295);
nand U6639 (N_6639,N_4552,N_2722);
nor U6640 (N_6640,N_2443,N_3328);
nor U6641 (N_6641,N_2129,N_3563);
nand U6642 (N_6642,N_367,N_959);
xnor U6643 (N_6643,N_875,N_2388);
nand U6644 (N_6644,N_1864,N_1197);
and U6645 (N_6645,N_1584,N_3087);
xnor U6646 (N_6646,N_3664,N_1908);
and U6647 (N_6647,N_446,N_2696);
and U6648 (N_6648,N_2185,N_336);
xor U6649 (N_6649,N_741,N_3018);
nor U6650 (N_6650,N_1451,N_3570);
or U6651 (N_6651,N_4154,N_3380);
or U6652 (N_6652,N_1281,N_3805);
and U6653 (N_6653,N_4319,N_773);
xnor U6654 (N_6654,N_4333,N_2405);
and U6655 (N_6655,N_1401,N_1808);
xnor U6656 (N_6656,N_4647,N_1642);
nand U6657 (N_6657,N_381,N_3156);
or U6658 (N_6658,N_996,N_816);
xor U6659 (N_6659,N_534,N_1077);
and U6660 (N_6660,N_2300,N_4165);
and U6661 (N_6661,N_4765,N_1816);
and U6662 (N_6662,N_1294,N_569);
nand U6663 (N_6663,N_59,N_1016);
xor U6664 (N_6664,N_3552,N_2341);
and U6665 (N_6665,N_4869,N_2348);
or U6666 (N_6666,N_2276,N_3844);
and U6667 (N_6667,N_1485,N_1333);
nor U6668 (N_6668,N_2423,N_2474);
xor U6669 (N_6669,N_3559,N_3856);
and U6670 (N_6670,N_1748,N_3748);
and U6671 (N_6671,N_1978,N_2379);
or U6672 (N_6672,N_774,N_3832);
nand U6673 (N_6673,N_957,N_4650);
or U6674 (N_6674,N_3467,N_4754);
or U6675 (N_6675,N_968,N_4003);
xor U6676 (N_6676,N_1655,N_197);
or U6677 (N_6677,N_4151,N_1037);
and U6678 (N_6678,N_3702,N_3072);
nor U6679 (N_6679,N_4777,N_3732);
nand U6680 (N_6680,N_1701,N_4330);
or U6681 (N_6681,N_2731,N_1099);
and U6682 (N_6682,N_2988,N_4141);
nor U6683 (N_6683,N_4073,N_1492);
nor U6684 (N_6684,N_4493,N_2358);
or U6685 (N_6685,N_1365,N_3160);
xor U6686 (N_6686,N_806,N_915);
nand U6687 (N_6687,N_3030,N_4923);
xor U6688 (N_6688,N_4428,N_282);
and U6689 (N_6689,N_3974,N_1180);
or U6690 (N_6690,N_2855,N_3991);
and U6691 (N_6691,N_1341,N_2323);
and U6692 (N_6692,N_2239,N_2887);
and U6693 (N_6693,N_664,N_3837);
nor U6694 (N_6694,N_1156,N_3981);
nand U6695 (N_6695,N_1685,N_3393);
nor U6696 (N_6696,N_4509,N_3289);
nand U6697 (N_6697,N_1558,N_3605);
xor U6698 (N_6698,N_2119,N_3229);
nand U6699 (N_6699,N_1219,N_2131);
xor U6700 (N_6700,N_3359,N_264);
or U6701 (N_6701,N_2943,N_3675);
and U6702 (N_6702,N_4049,N_628);
nand U6703 (N_6703,N_3488,N_4945);
nor U6704 (N_6704,N_4562,N_4636);
or U6705 (N_6705,N_1093,N_1324);
xnor U6706 (N_6706,N_292,N_800);
nor U6707 (N_6707,N_1457,N_4442);
nand U6708 (N_6708,N_4299,N_4429);
or U6709 (N_6709,N_4627,N_1367);
and U6710 (N_6710,N_440,N_4540);
nand U6711 (N_6711,N_4810,N_2551);
nand U6712 (N_6712,N_1589,N_2203);
nand U6713 (N_6713,N_2526,N_3147);
nand U6714 (N_6714,N_3851,N_99);
nor U6715 (N_6715,N_824,N_124);
nand U6716 (N_6716,N_2318,N_490);
and U6717 (N_6717,N_2530,N_4485);
and U6718 (N_6718,N_1578,N_3069);
or U6719 (N_6719,N_466,N_4951);
and U6720 (N_6720,N_4630,N_290);
nand U6721 (N_6721,N_2734,N_4910);
and U6722 (N_6722,N_2257,N_1153);
and U6723 (N_6723,N_1318,N_4537);
and U6724 (N_6724,N_3638,N_2825);
xor U6725 (N_6725,N_1507,N_222);
xor U6726 (N_6726,N_4663,N_1237);
nand U6727 (N_6727,N_4678,N_1854);
or U6728 (N_6728,N_3011,N_1833);
nor U6729 (N_6729,N_138,N_1516);
nand U6730 (N_6730,N_1200,N_3432);
nor U6731 (N_6731,N_3583,N_4254);
nor U6732 (N_6732,N_3668,N_4242);
nor U6733 (N_6733,N_619,N_4556);
and U6734 (N_6734,N_1774,N_1396);
xor U6735 (N_6735,N_2484,N_4324);
and U6736 (N_6736,N_3444,N_1840);
nor U6737 (N_6737,N_4668,N_4005);
xnor U6738 (N_6738,N_2896,N_1964);
nand U6739 (N_6739,N_2340,N_4068);
nand U6740 (N_6740,N_4458,N_1986);
nor U6741 (N_6741,N_4294,N_4218);
xor U6742 (N_6742,N_1802,N_1823);
and U6743 (N_6743,N_1519,N_4336);
nor U6744 (N_6744,N_2149,N_225);
xnor U6745 (N_6745,N_4378,N_2500);
xnor U6746 (N_6746,N_3355,N_2275);
and U6747 (N_6747,N_3254,N_2704);
or U6748 (N_6748,N_2924,N_4419);
or U6749 (N_6749,N_620,N_2262);
xor U6750 (N_6750,N_31,N_4751);
or U6751 (N_6751,N_2415,N_1996);
xor U6752 (N_6752,N_3813,N_1636);
and U6753 (N_6753,N_3584,N_1539);
or U6754 (N_6754,N_842,N_3175);
or U6755 (N_6755,N_4290,N_3186);
and U6756 (N_6756,N_4614,N_2590);
or U6757 (N_6757,N_1299,N_987);
or U6758 (N_6758,N_4359,N_927);
or U6759 (N_6759,N_881,N_48);
xnor U6760 (N_6760,N_2809,N_4763);
and U6761 (N_6761,N_3438,N_2917);
nor U6762 (N_6762,N_2627,N_2003);
xor U6763 (N_6763,N_365,N_2502);
nor U6764 (N_6764,N_2088,N_4929);
xnor U6765 (N_6765,N_786,N_2);
xor U6766 (N_6766,N_2478,N_4075);
nand U6767 (N_6767,N_189,N_4422);
xor U6768 (N_6768,N_2233,N_803);
and U6769 (N_6769,N_1767,N_2219);
nand U6770 (N_6770,N_4961,N_2043);
or U6771 (N_6771,N_3461,N_427);
and U6772 (N_6772,N_1327,N_3051);
nor U6773 (N_6773,N_4114,N_969);
and U6774 (N_6774,N_1126,N_2754);
nor U6775 (N_6775,N_4535,N_4310);
xnor U6776 (N_6776,N_3469,N_156);
xnor U6777 (N_6777,N_1985,N_2125);
nor U6778 (N_6778,N_3422,N_2770);
or U6779 (N_6779,N_829,N_2976);
or U6780 (N_6780,N_1250,N_3973);
xor U6781 (N_6781,N_4652,N_4153);
nor U6782 (N_6782,N_2804,N_2810);
xnor U6783 (N_6783,N_2081,N_3322);
or U6784 (N_6784,N_2978,N_3764);
nand U6785 (N_6785,N_3627,N_4675);
nand U6786 (N_6786,N_2053,N_3621);
and U6787 (N_6787,N_2169,N_3839);
nand U6788 (N_6788,N_1693,N_952);
and U6789 (N_6789,N_642,N_3323);
nor U6790 (N_6790,N_4889,N_2658);
xor U6791 (N_6791,N_4657,N_4959);
and U6792 (N_6792,N_528,N_2854);
or U6793 (N_6793,N_4659,N_1158);
and U6794 (N_6794,N_2689,N_1754);
xor U6795 (N_6795,N_2581,N_2373);
xor U6796 (N_6796,N_3522,N_157);
or U6797 (N_6797,N_621,N_309);
nand U6798 (N_6798,N_325,N_1438);
and U6799 (N_6799,N_3737,N_4238);
nor U6800 (N_6800,N_243,N_1770);
or U6801 (N_6801,N_3902,N_2049);
or U6802 (N_6802,N_4130,N_2926);
xnor U6803 (N_6803,N_4096,N_3399);
xnor U6804 (N_6804,N_2161,N_2857);
nor U6805 (N_6805,N_2753,N_4388);
and U6806 (N_6806,N_1906,N_3854);
xor U6807 (N_6807,N_11,N_799);
nor U6808 (N_6808,N_3358,N_2948);
nand U6809 (N_6809,N_3587,N_3791);
xnor U6810 (N_6810,N_3554,N_4977);
or U6811 (N_6811,N_4671,N_2815);
nand U6812 (N_6812,N_3436,N_704);
nand U6813 (N_6813,N_4502,N_2363);
nor U6814 (N_6814,N_2780,N_591);
xor U6815 (N_6815,N_57,N_3024);
nand U6816 (N_6816,N_2712,N_1672);
nor U6817 (N_6817,N_3258,N_3505);
or U6818 (N_6818,N_4665,N_981);
or U6819 (N_6819,N_133,N_4664);
or U6820 (N_6820,N_2010,N_924);
or U6821 (N_6821,N_891,N_2779);
or U6822 (N_6822,N_681,N_2750);
and U6823 (N_6823,N_934,N_483);
xor U6824 (N_6824,N_1421,N_2253);
xor U6825 (N_6825,N_879,N_1595);
and U6826 (N_6826,N_545,N_4274);
xor U6827 (N_6827,N_4639,N_1014);
nand U6828 (N_6828,N_3404,N_3674);
nor U6829 (N_6829,N_4270,N_1791);
nor U6830 (N_6830,N_530,N_1470);
or U6831 (N_6831,N_3665,N_2279);
nor U6832 (N_6832,N_242,N_2584);
or U6833 (N_6833,N_2736,N_4995);
nand U6834 (N_6834,N_3720,N_1026);
nor U6835 (N_6835,N_3217,N_1224);
nor U6836 (N_6836,N_1193,N_4457);
nor U6837 (N_6837,N_4103,N_4385);
and U6838 (N_6838,N_852,N_353);
nand U6839 (N_6839,N_3446,N_1930);
xor U6840 (N_6840,N_1038,N_4686);
xnor U6841 (N_6841,N_1048,N_1003);
or U6842 (N_6842,N_2069,N_3277);
nor U6843 (N_6843,N_2895,N_3657);
or U6844 (N_6844,N_4868,N_4321);
nor U6845 (N_6845,N_643,N_2659);
nand U6846 (N_6846,N_4709,N_3891);
nor U6847 (N_6847,N_3398,N_3487);
nand U6848 (N_6848,N_3145,N_1975);
and U6849 (N_6849,N_1855,N_2342);
nor U6850 (N_6850,N_4208,N_4782);
nor U6851 (N_6851,N_1844,N_1661);
xor U6852 (N_6852,N_2397,N_4454);
and U6853 (N_6853,N_4412,N_1434);
xnor U6854 (N_6854,N_2778,N_217);
and U6855 (N_6855,N_2191,N_1542);
and U6856 (N_6856,N_4406,N_1046);
nand U6857 (N_6857,N_3447,N_4794);
nand U6858 (N_6858,N_119,N_163);
or U6859 (N_6859,N_3711,N_1436);
or U6860 (N_6860,N_2083,N_3118);
and U6861 (N_6861,N_2583,N_1769);
nand U6862 (N_6862,N_815,N_1648);
xnor U6863 (N_6863,N_1901,N_1797);
and U6864 (N_6864,N_2849,N_663);
nor U6865 (N_6865,N_2625,N_4724);
xor U6866 (N_6866,N_4617,N_1190);
nor U6867 (N_6867,N_41,N_169);
nand U6868 (N_6868,N_350,N_2693);
nand U6869 (N_6869,N_2419,N_1706);
xnor U6870 (N_6870,N_3247,N_4820);
xor U6871 (N_6871,N_2296,N_4014);
nor U6872 (N_6872,N_809,N_358);
nand U6873 (N_6873,N_3783,N_4170);
or U6874 (N_6874,N_2974,N_1514);
and U6875 (N_6875,N_2067,N_2019);
xnor U6876 (N_6876,N_301,N_1845);
and U6877 (N_6877,N_2334,N_4550);
and U6878 (N_6878,N_4488,N_4441);
nand U6879 (N_6879,N_421,N_596);
xor U6880 (N_6880,N_317,N_2616);
nor U6881 (N_6881,N_287,N_3237);
or U6882 (N_6882,N_4759,N_3074);
and U6883 (N_6883,N_3636,N_1733);
xnor U6884 (N_6884,N_4915,N_4941);
nand U6885 (N_6885,N_4600,N_4125);
nand U6886 (N_6886,N_4594,N_2510);
or U6887 (N_6887,N_1487,N_1441);
xor U6888 (N_6888,N_3879,N_3287);
nand U6889 (N_6889,N_971,N_3230);
and U6890 (N_6890,N_4427,N_1112);
nand U6891 (N_6891,N_471,N_1695);
or U6892 (N_6892,N_750,N_751);
xnor U6893 (N_6893,N_3815,N_0);
xnor U6894 (N_6894,N_4536,N_144);
nor U6895 (N_6895,N_2646,N_2076);
nand U6896 (N_6896,N_248,N_583);
or U6897 (N_6897,N_2093,N_945);
or U6898 (N_6898,N_3106,N_327);
xor U6899 (N_6899,N_1444,N_1910);
and U6900 (N_6900,N_3375,N_1720);
nor U6901 (N_6901,N_2717,N_1751);
nor U6902 (N_6902,N_4545,N_3564);
nand U6903 (N_6903,N_81,N_76);
nand U6904 (N_6904,N_2263,N_1870);
and U6905 (N_6905,N_35,N_2996);
nor U6906 (N_6906,N_1746,N_2097);
and U6907 (N_6907,N_3397,N_4519);
xor U6908 (N_6908,N_1067,N_520);
xor U6909 (N_6909,N_2527,N_4500);
or U6910 (N_6910,N_1927,N_3036);
and U6911 (N_6911,N_3786,N_3232);
nand U6912 (N_6912,N_3330,N_3708);
nand U6913 (N_6913,N_306,N_3161);
xor U6914 (N_6914,N_4462,N_21);
nand U6915 (N_6915,N_1929,N_3274);
nor U6916 (N_6916,N_2544,N_1506);
xor U6917 (N_6917,N_2634,N_1663);
or U6918 (N_6918,N_923,N_14);
xnor U6919 (N_6919,N_1432,N_1386);
xor U6920 (N_6920,N_2322,N_2792);
or U6921 (N_6921,N_2437,N_4314);
or U6922 (N_6922,N_743,N_2619);
and U6923 (N_6923,N_2394,N_1924);
and U6924 (N_6924,N_4893,N_1490);
nor U6925 (N_6925,N_2514,N_3040);
and U6926 (N_6926,N_4579,N_3591);
or U6927 (N_6927,N_1313,N_674);
nor U6928 (N_6928,N_912,N_4954);
or U6929 (N_6929,N_2697,N_356);
or U6930 (N_6930,N_2382,N_2111);
or U6931 (N_6931,N_3943,N_2154);
nor U6932 (N_6932,N_4792,N_2410);
nor U6933 (N_6933,N_588,N_3476);
xor U6934 (N_6934,N_4467,N_1175);
xor U6935 (N_6935,N_4928,N_304);
nor U6936 (N_6936,N_2467,N_3985);
and U6937 (N_6937,N_2786,N_338);
and U6938 (N_6938,N_958,N_1875);
and U6939 (N_6939,N_3009,N_2011);
nand U6940 (N_6940,N_1080,N_4881);
xor U6941 (N_6941,N_2217,N_1879);
nand U6942 (N_6942,N_3352,N_675);
nor U6943 (N_6943,N_4479,N_4631);
nand U6944 (N_6944,N_859,N_1645);
nand U6945 (N_6945,N_1923,N_2821);
xnor U6946 (N_6946,N_1482,N_4392);
xnor U6947 (N_6947,N_3528,N_3503);
nand U6948 (N_6948,N_4316,N_2306);
nor U6949 (N_6949,N_1860,N_380);
xor U6950 (N_6950,N_567,N_2981);
and U6951 (N_6951,N_3297,N_604);
nand U6952 (N_6952,N_1859,N_4802);
or U6953 (N_6953,N_3695,N_4283);
nand U6954 (N_6954,N_832,N_2251);
and U6955 (N_6955,N_4744,N_4986);
nor U6956 (N_6956,N_80,N_3027);
nor U6957 (N_6957,N_3648,N_2078);
xnor U6958 (N_6958,N_515,N_4870);
and U6959 (N_6959,N_3964,N_2241);
nor U6960 (N_6960,N_2268,N_1610);
and U6961 (N_6961,N_833,N_4201);
or U6962 (N_6962,N_2413,N_4352);
and U6963 (N_6963,N_1696,N_147);
and U6964 (N_6964,N_3005,N_2385);
nor U6965 (N_6965,N_4161,N_72);
xnor U6966 (N_6966,N_3835,N_1856);
nor U6967 (N_6967,N_98,N_2482);
nor U6968 (N_6968,N_1540,N_3785);
nor U6969 (N_6969,N_2327,N_2910);
nor U6970 (N_6970,N_4217,N_523);
nand U6971 (N_6971,N_947,N_1658);
nor U6972 (N_6972,N_617,N_2332);
xnor U6973 (N_6973,N_3215,N_61);
and U6974 (N_6974,N_2533,N_1394);
nor U6975 (N_6975,N_850,N_1052);
nor U6976 (N_6976,N_2915,N_2547);
and U6977 (N_6977,N_3531,N_1904);
or U6978 (N_6978,N_4344,N_3102);
and U6979 (N_6979,N_3645,N_1131);
nand U6980 (N_6980,N_3368,N_277);
xor U6981 (N_6981,N_898,N_1142);
xor U6982 (N_6982,N_2196,N_3045);
and U6983 (N_6983,N_710,N_2663);
or U6984 (N_6984,N_4574,N_1651);
or U6985 (N_6985,N_4694,N_3088);
or U6986 (N_6986,N_4874,N_1521);
and U6987 (N_6987,N_716,N_4042);
nor U6988 (N_6988,N_1646,N_4723);
nand U6989 (N_6989,N_1468,N_4198);
and U6990 (N_6990,N_1102,N_533);
nor U6991 (N_6991,N_101,N_160);
xor U6992 (N_6992,N_2352,N_2065);
xor U6993 (N_6993,N_1045,N_1212);
and U6994 (N_6994,N_2535,N_3490);
and U6995 (N_6995,N_1117,N_4729);
and U6996 (N_6996,N_1144,N_2319);
and U6997 (N_6997,N_1440,N_199);
nor U6998 (N_6998,N_1013,N_293);
nand U6999 (N_6999,N_729,N_150);
nor U7000 (N_7000,N_109,N_3841);
nor U7001 (N_7001,N_3719,N_4761);
or U7002 (N_7002,N_2609,N_4993);
nor U7003 (N_7003,N_3694,N_3151);
xnor U7004 (N_7004,N_1987,N_2671);
nand U7005 (N_7005,N_1268,N_4538);
or U7006 (N_7006,N_3329,N_1074);
xor U7007 (N_7007,N_3898,N_2795);
nor U7008 (N_7008,N_4323,N_2794);
nor U7009 (N_7009,N_3403,N_2942);
nand U7010 (N_7010,N_2452,N_835);
nand U7011 (N_7011,N_4327,N_1805);
nor U7012 (N_7012,N_1653,N_360);
or U7013 (N_7013,N_2031,N_1198);
xor U7014 (N_7014,N_4341,N_4269);
or U7015 (N_7015,N_95,N_2255);
xor U7016 (N_7016,N_2903,N_4696);
xor U7017 (N_7017,N_2439,N_2970);
or U7018 (N_7018,N_4690,N_470);
and U7019 (N_7019,N_4215,N_2375);
xnor U7020 (N_7020,N_2189,N_922);
nor U7021 (N_7021,N_3449,N_2252);
nor U7022 (N_7022,N_703,N_442);
xor U7023 (N_7023,N_3842,N_4748);
nand U7024 (N_7024,N_3192,N_2513);
nor U7025 (N_7025,N_3634,N_2386);
nand U7026 (N_7026,N_4387,N_2145);
or U7027 (N_7027,N_4621,N_1932);
or U7028 (N_7028,N_1302,N_326);
and U7029 (N_7029,N_3772,N_718);
nand U7030 (N_7030,N_1148,N_856);
or U7031 (N_7031,N_2018,N_890);
and U7032 (N_7032,N_2292,N_720);
nand U7033 (N_7033,N_1086,N_3418);
xnor U7034 (N_7034,N_1736,N_3220);
xor U7035 (N_7035,N_4646,N_3216);
or U7036 (N_7036,N_3154,N_2064);
xor U7037 (N_7037,N_3158,N_3038);
and U7038 (N_7038,N_3892,N_1480);
or U7039 (N_7039,N_3939,N_2721);
or U7040 (N_7040,N_904,N_4662);
or U7041 (N_7041,N_3688,N_3451);
xor U7042 (N_7042,N_3700,N_375);
nor U7043 (N_7043,N_2690,N_817);
xor U7044 (N_7044,N_3518,N_4987);
nand U7045 (N_7045,N_3163,N_2938);
nand U7046 (N_7046,N_571,N_2436);
and U7047 (N_7047,N_2024,N_574);
xor U7048 (N_7048,N_159,N_419);
nor U7049 (N_7049,N_1287,N_2858);
and U7050 (N_7050,N_1095,N_2238);
or U7051 (N_7051,N_3860,N_882);
xnor U7052 (N_7052,N_562,N_877);
nand U7053 (N_7053,N_2372,N_4602);
xnor U7054 (N_7054,N_1723,N_711);
or U7055 (N_7055,N_60,N_4225);
and U7056 (N_7056,N_3089,N_2039);
nor U7057 (N_7057,N_713,N_795);
or U7058 (N_7058,N_1580,N_185);
nand U7059 (N_7059,N_1995,N_469);
and U7060 (N_7060,N_4176,N_3890);
or U7061 (N_7061,N_2346,N_582);
nor U7062 (N_7062,N_2523,N_1204);
nor U7063 (N_7063,N_2290,N_3382);
xor U7064 (N_7064,N_3955,N_2244);
and U7065 (N_7065,N_561,N_4541);
nand U7066 (N_7066,N_4523,N_3354);
nor U7067 (N_7067,N_563,N_3066);
xnor U7068 (N_7068,N_4384,N_281);
nor U7069 (N_7069,N_2313,N_4879);
nand U7070 (N_7070,N_3356,N_4967);
nand U7071 (N_7071,N_3242,N_3822);
nor U7072 (N_7072,N_954,N_4495);
xor U7073 (N_7073,N_364,N_4279);
xnor U7074 (N_7074,N_2116,N_4080);
and U7075 (N_7075,N_4245,N_125);
nor U7076 (N_7076,N_1821,N_3311);
xnor U7077 (N_7077,N_4897,N_866);
or U7078 (N_7078,N_4766,N_3244);
or U7079 (N_7079,N_1522,N_2864);
nand U7080 (N_7080,N_597,N_2881);
or U7081 (N_7081,N_1550,N_2133);
nor U7082 (N_7082,N_4505,N_4806);
xnor U7083 (N_7083,N_71,N_2056);
nand U7084 (N_7084,N_4083,N_3303);
nor U7085 (N_7085,N_2971,N_1136);
or U7086 (N_7086,N_1704,N_4816);
xnor U7087 (N_7087,N_536,N_752);
xnor U7088 (N_7088,N_386,N_1062);
nor U7089 (N_7089,N_3821,N_1381);
xnor U7090 (N_7090,N_1954,N_3134);
nor U7091 (N_7091,N_3405,N_2271);
or U7092 (N_7092,N_1300,N_3291);
nor U7093 (N_7093,N_900,N_3999);
and U7094 (N_7094,N_289,N_2061);
xor U7095 (N_7095,N_50,N_3381);
nand U7096 (N_7096,N_1196,N_4821);
nor U7097 (N_7097,N_955,N_2957);
nand U7098 (N_7098,N_2579,N_51);
and U7099 (N_7099,N_2546,N_4813);
nor U7100 (N_7100,N_3378,N_1674);
or U7101 (N_7101,N_2148,N_37);
nor U7102 (N_7102,N_684,N_3052);
and U7103 (N_7103,N_4436,N_477);
xnor U7104 (N_7104,N_450,N_4885);
or U7105 (N_7105,N_887,N_4866);
and U7106 (N_7106,N_3504,N_3828);
nand U7107 (N_7107,N_3799,N_1825);
nand U7108 (N_7108,N_4061,N_4817);
nand U7109 (N_7109,N_4711,N_1552);
and U7110 (N_7110,N_3477,N_3023);
or U7111 (N_7111,N_1227,N_2919);
and U7112 (N_7112,N_2230,N_1132);
or U7113 (N_7113,N_4293,N_2256);
nor U7114 (N_7114,N_1411,N_1530);
and U7115 (N_7115,N_2893,N_4906);
nor U7116 (N_7116,N_2827,N_1392);
or U7117 (N_7117,N_748,N_2628);
nand U7118 (N_7118,N_3367,N_1356);
nor U7119 (N_7119,N_993,N_1473);
nor U7120 (N_7120,N_3749,N_1803);
and U7121 (N_7121,N_2400,N_1258);
and U7122 (N_7122,N_1905,N_1940);
and U7123 (N_7123,N_3417,N_4029);
nand U7124 (N_7124,N_769,N_1933);
and U7125 (N_7125,N_3927,N_3746);
or U7126 (N_7126,N_1681,N_871);
or U7127 (N_7127,N_449,N_759);
and U7128 (N_7128,N_1089,N_2007);
or U7129 (N_7129,N_4287,N_3373);
nand U7130 (N_7130,N_4597,N_1344);
or U7131 (N_7131,N_4992,N_1705);
nor U7132 (N_7132,N_3450,N_739);
xnor U7133 (N_7133,N_4331,N_4947);
nor U7134 (N_7134,N_1815,N_4822);
nor U7135 (N_7135,N_2789,N_3286);
xnor U7136 (N_7136,N_2798,N_178);
or U7137 (N_7137,N_1254,N_422);
or U7138 (N_7138,N_2345,N_3885);
and U7139 (N_7139,N_2470,N_586);
or U7140 (N_7140,N_3996,N_1357);
and U7141 (N_7141,N_1417,N_802);
nor U7142 (N_7142,N_3091,N_3127);
nor U7143 (N_7143,N_2442,N_2738);
nand U7144 (N_7144,N_429,N_3921);
and U7145 (N_7145,N_3165,N_2983);
and U7146 (N_7146,N_2515,N_1544);
xor U7147 (N_7147,N_4033,N_1173);
nand U7148 (N_7148,N_3961,N_2733);
and U7149 (N_7149,N_2769,N_285);
nor U7150 (N_7150,N_2517,N_1798);
or U7151 (N_7151,N_3110,N_1953);
and U7152 (N_7152,N_1867,N_4177);
nand U7153 (N_7153,N_247,N_1858);
and U7154 (N_7154,N_4119,N_1122);
or U7155 (N_7155,N_936,N_2766);
or U7156 (N_7156,N_1162,N_1412);
xor U7157 (N_7157,N_1764,N_2710);
or U7158 (N_7158,N_4689,N_754);
xor U7159 (N_7159,N_330,N_2073);
and U7160 (N_7160,N_849,N_1630);
nor U7161 (N_7161,N_4139,N_2725);
xor U7162 (N_7162,N_1811,N_1919);
and U7163 (N_7163,N_2430,N_2683);
nor U7164 (N_7164,N_4922,N_2913);
xor U7165 (N_7165,N_3483,N_311);
or U7166 (N_7166,N_2480,N_845);
nand U7167 (N_7167,N_3663,N_3715);
xnor U7168 (N_7168,N_342,N_3508);
nand U7169 (N_7169,N_1282,N_4063);
xnor U7170 (N_7170,N_4926,N_2008);
nor U7171 (N_7171,N_1372,N_425);
nand U7172 (N_7172,N_785,N_2863);
xor U7173 (N_7173,N_40,N_980);
and U7174 (N_7174,N_1460,N_4202);
xnor U7175 (N_7175,N_3826,N_1477);
nand U7176 (N_7176,N_1489,N_270);
and U7177 (N_7177,N_4643,N_3170);
xnor U7178 (N_7178,N_165,N_4199);
and U7179 (N_7179,N_175,N_404);
and U7180 (N_7180,N_910,N_3536);
and U7181 (N_7181,N_3753,N_1040);
and U7182 (N_7182,N_1563,N_1123);
nor U7183 (N_7183,N_3025,N_4081);
xor U7184 (N_7184,N_2856,N_4437);
or U7185 (N_7185,N_2931,N_4174);
nand U7186 (N_7186,N_3043,N_1107);
nor U7187 (N_7187,N_4380,N_3535);
and U7188 (N_7188,N_4097,N_229);
and U7189 (N_7189,N_3172,N_2838);
nor U7190 (N_7190,N_4223,N_1694);
xor U7191 (N_7191,N_2615,N_3510);
and U7192 (N_7192,N_43,N_4426);
nor U7193 (N_7193,N_2416,N_3430);
and U7194 (N_7194,N_4733,N_3804);
or U7195 (N_7195,N_1541,N_2449);
xor U7196 (N_7196,N_4876,N_3141);
xor U7197 (N_7197,N_2594,N_2927);
and U7198 (N_7198,N_478,N_2799);
and U7199 (N_7199,N_3434,N_445);
nor U7200 (N_7200,N_1882,N_4895);
or U7201 (N_7201,N_2123,N_2094);
nand U7202 (N_7202,N_2833,N_2040);
nor U7203 (N_7203,N_3667,N_4055);
nand U7204 (N_7204,N_3350,N_4037);
xor U7205 (N_7205,N_2173,N_4446);
xnor U7206 (N_7206,N_283,N_4952);
nand U7207 (N_7207,N_2209,N_3284);
xor U7208 (N_7208,N_2805,N_4263);
nand U7209 (N_7209,N_3918,N_1945);
nor U7210 (N_7210,N_667,N_1806);
and U7211 (N_7211,N_1474,N_4854);
nor U7212 (N_7212,N_4297,N_2455);
xor U7213 (N_7213,N_3492,N_1140);
and U7214 (N_7214,N_1789,N_251);
or U7215 (N_7215,N_2164,N_3288);
nand U7216 (N_7216,N_4449,N_1354);
xor U7217 (N_7217,N_2160,N_2329);
or U7218 (N_7218,N_411,N_4018);
xnor U7219 (N_7219,N_1628,N_1772);
nand U7220 (N_7220,N_1861,N_3261);
or U7221 (N_7221,N_1562,N_772);
or U7222 (N_7222,N_1968,N_3976);
xor U7223 (N_7223,N_3276,N_1785);
xnor U7224 (N_7224,N_2466,N_3569);
nor U7225 (N_7225,N_3852,N_2286);
and U7226 (N_7226,N_1247,N_391);
nand U7227 (N_7227,N_3859,N_2783);
and U7228 (N_7228,N_725,N_1503);
or U7229 (N_7229,N_1034,N_3910);
xor U7230 (N_7230,N_570,N_295);
and U7231 (N_7231,N_2224,N_4551);
and U7232 (N_7232,N_2654,N_4707);
and U7233 (N_7233,N_1728,N_901);
nand U7234 (N_7234,N_4496,N_3792);
nand U7235 (N_7235,N_151,N_4123);
or U7236 (N_7236,N_4950,N_3090);
or U7237 (N_7237,N_3372,N_4439);
and U7238 (N_7238,N_4102,N_3829);
xnor U7239 (N_7239,N_811,N_2553);
xnor U7240 (N_7240,N_4956,N_1687);
nor U7241 (N_7241,N_3681,N_1683);
nand U7242 (N_7242,N_1233,N_1690);
and U7243 (N_7243,N_3840,N_322);
nor U7244 (N_7244,N_3672,N_655);
and U7245 (N_7245,N_805,N_2328);
and U7246 (N_7246,N_1015,N_52);
and U7247 (N_7247,N_3830,N_120);
or U7248 (N_7248,N_3915,N_102);
xnor U7249 (N_7249,N_3337,N_3471);
nor U7250 (N_7250,N_2309,N_4132);
or U7251 (N_7251,N_1511,N_1551);
nand U7252 (N_7252,N_3099,N_3305);
and U7253 (N_7253,N_4252,N_1991);
and U7254 (N_7254,N_1004,N_3814);
nor U7255 (N_7255,N_1047,N_3707);
and U7256 (N_7256,N_2829,N_2521);
or U7257 (N_7257,N_962,N_2490);
or U7258 (N_7258,N_1479,N_15);
and U7259 (N_7259,N_1149,N_118);
nand U7260 (N_7260,N_431,N_1609);
or U7261 (N_7261,N_2596,N_2297);
nor U7262 (N_7262,N_253,N_3201);
xnor U7263 (N_7263,N_2427,N_423);
nor U7264 (N_7264,N_1152,N_114);
or U7265 (N_7265,N_4974,N_2364);
or U7266 (N_7266,N_4524,N_2687);
nor U7267 (N_7267,N_2493,N_883);
and U7268 (N_7268,N_4515,N_791);
xnor U7269 (N_7269,N_89,N_1742);
nor U7270 (N_7270,N_4715,N_3931);
or U7271 (N_7271,N_1032,N_3917);
nand U7272 (N_7272,N_2311,N_1594);
nand U7273 (N_7273,N_3717,N_814);
nor U7274 (N_7274,N_998,N_2235);
nand U7275 (N_7275,N_2606,N_141);
or U7276 (N_7276,N_3767,N_97);
nand U7277 (N_7277,N_2939,N_66);
or U7278 (N_7278,N_2918,N_2965);
nand U7279 (N_7279,N_4828,N_4793);
nand U7280 (N_7280,N_3651,N_3265);
nand U7281 (N_7281,N_3755,N_976);
nand U7282 (N_7282,N_557,N_2005);
xor U7283 (N_7283,N_2460,N_2558);
nand U7284 (N_7284,N_1783,N_4219);
nand U7285 (N_7285,N_321,N_2613);
nand U7286 (N_7286,N_1679,N_4520);
nor U7287 (N_7287,N_1782,N_4577);
nor U7288 (N_7288,N_2862,N_926);
or U7289 (N_7289,N_2742,N_3139);
nor U7290 (N_7290,N_4804,N_3182);
nand U7291 (N_7291,N_372,N_1813);
xnor U7292 (N_7292,N_821,N_2072);
xor U7293 (N_7293,N_2440,N_2623);
nand U7294 (N_7294,N_2707,N_2247);
or U7295 (N_7295,N_63,N_688);
xor U7296 (N_7296,N_4857,N_4569);
nand U7297 (N_7297,N_1413,N_1163);
nand U7298 (N_7298,N_727,N_590);
nand U7299 (N_7299,N_447,N_1824);
nand U7300 (N_7300,N_854,N_1847);
and U7301 (N_7301,N_4261,N_3966);
or U7302 (N_7302,N_4634,N_4415);
nand U7303 (N_7303,N_4148,N_68);
xnor U7304 (N_7304,N_2730,N_3506);
xor U7305 (N_7305,N_828,N_3846);
nand U7306 (N_7306,N_3414,N_401);
or U7307 (N_7307,N_2184,N_4459);
xnor U7308 (N_7308,N_4189,N_86);
nand U7309 (N_7309,N_2333,N_3653);
or U7310 (N_7310,N_2841,N_2202);
xor U7311 (N_7311,N_963,N_3060);
or U7312 (N_7312,N_872,N_3148);
nor U7313 (N_7313,N_4251,N_3970);
nor U7314 (N_7314,N_884,N_1753);
or U7315 (N_7315,N_1057,N_787);
or U7316 (N_7316,N_1207,N_777);
xor U7317 (N_7317,N_1419,N_982);
or U7318 (N_7318,N_3599,N_3523);
xor U7319 (N_7319,N_1547,N_2636);
nor U7320 (N_7320,N_2284,N_3586);
and U7321 (N_7321,N_2902,N_2242);
and U7322 (N_7322,N_190,N_2454);
and U7323 (N_7323,N_4407,N_4032);
or U7324 (N_7324,N_1319,N_3686);
or U7325 (N_7325,N_2080,N_2180);
and U7326 (N_7326,N_602,N_238);
or U7327 (N_7327,N_3944,N_3472);
nor U7328 (N_7328,N_3874,N_1902);
nor U7329 (N_7329,N_2070,N_4670);
xor U7330 (N_7330,N_735,N_2171);
xnor U7331 (N_7331,N_3759,N_3463);
nor U7332 (N_7332,N_4916,N_4400);
or U7333 (N_7333,N_1283,N_129);
nor U7334 (N_7334,N_46,N_4685);
nand U7335 (N_7335,N_1637,N_3076);
and U7336 (N_7336,N_1569,N_3010);
and U7337 (N_7337,N_662,N_2102);
xor U7338 (N_7338,N_1943,N_1320);
or U7339 (N_7339,N_1315,N_4017);
or U7340 (N_7340,N_1072,N_4303);
nor U7341 (N_7341,N_3546,N_2865);
nand U7342 (N_7342,N_1920,N_4826);
xor U7343 (N_7343,N_2744,N_2975);
and U7344 (N_7344,N_2979,N_1488);
and U7345 (N_7345,N_3243,N_1000);
nor U7346 (N_7346,N_2723,N_2565);
and U7347 (N_7347,N_2398,N_896);
xor U7348 (N_7348,N_3581,N_4611);
nor U7349 (N_7349,N_3248,N_3947);
or U7350 (N_7350,N_4034,N_3575);
or U7351 (N_7351,N_3268,N_3347);
and U7352 (N_7352,N_3429,N_858);
nor U7353 (N_7353,N_4677,N_1982);
and U7354 (N_7354,N_2986,N_2997);
nor U7355 (N_7355,N_3682,N_4028);
xor U7356 (N_7356,N_2216,N_3144);
and U7357 (N_7357,N_2987,N_3493);
and U7358 (N_7358,N_2422,N_4638);
nand U7359 (N_7359,N_38,N_4726);
or U7360 (N_7360,N_4582,N_182);
or U7361 (N_7361,N_339,N_4625);
or U7362 (N_7362,N_4265,N_938);
and U7363 (N_7363,N_1202,N_3857);
nor U7364 (N_7364,N_733,N_2412);
or U7365 (N_7365,N_1548,N_4938);
nor U7366 (N_7366,N_2765,N_2237);
nand U7367 (N_7367,N_4140,N_1579);
nor U7368 (N_7368,N_1682,N_2353);
xnor U7369 (N_7369,N_1621,N_2560);
and U7370 (N_7370,N_840,N_2389);
or U7371 (N_7371,N_2132,N_3758);
xnor U7372 (N_7372,N_361,N_3685);
nor U7373 (N_7373,N_4558,N_4865);
nand U7374 (N_7374,N_4803,N_1310);
or U7375 (N_7375,N_1673,N_4431);
nand U7376 (N_7376,N_1010,N_4025);
nor U7377 (N_7377,N_2337,N_3206);
and U7378 (N_7378,N_1155,N_333);
nand U7379 (N_7379,N_2044,N_3335);
and U7380 (N_7380,N_4839,N_3906);
nor U7381 (N_7381,N_4470,N_4586);
or U7382 (N_7382,N_1498,N_158);
or U7383 (N_7383,N_2450,N_4070);
or U7384 (N_7384,N_873,N_3150);
xor U7385 (N_7385,N_3205,N_3949);
nand U7386 (N_7386,N_3180,N_2136);
xnor U7387 (N_7387,N_4883,N_4920);
and U7388 (N_7388,N_3049,N_4982);
nor U7389 (N_7389,N_1210,N_4718);
nor U7390 (N_7390,N_183,N_4900);
nand U7391 (N_7391,N_4892,N_4107);
or U7392 (N_7392,N_1446,N_2028);
nor U7393 (N_7393,N_3789,N_3652);
nor U7394 (N_7394,N_1939,N_3739);
nor U7395 (N_7395,N_1804,N_2456);
nor U7396 (N_7396,N_696,N_3055);
nand U7397 (N_7397,N_529,N_4181);
nor U7398 (N_7398,N_3202,N_4591);
nand U7399 (N_7399,N_3140,N_3995);
xnor U7400 (N_7400,N_3462,N_1334);
nor U7401 (N_7401,N_2091,N_1231);
xnor U7402 (N_7402,N_397,N_4924);
xnor U7403 (N_7403,N_2670,N_706);
and U7404 (N_7404,N_4548,N_210);
or U7405 (N_7405,N_683,N_2868);
or U7406 (N_7406,N_4021,N_906);
nor U7407 (N_7407,N_1243,N_2486);
or U7408 (N_7408,N_4363,N_1617);
and U7409 (N_7409,N_4115,N_1448);
nand U7410 (N_7410,N_3752,N_1273);
xor U7411 (N_7411,N_4656,N_612);
xor U7412 (N_7412,N_4934,N_2556);
or U7413 (N_7413,N_2376,N_4364);
nor U7414 (N_7414,N_3521,N_255);
or U7415 (N_7415,N_519,N_4360);
xnor U7416 (N_7416,N_3470,N_1246);
or U7417 (N_7417,N_2545,N_3246);
and U7418 (N_7418,N_4237,N_2787);
or U7419 (N_7419,N_988,N_946);
xor U7420 (N_7420,N_1147,N_134);
or U7421 (N_7421,N_853,N_4598);
or U7422 (N_7422,N_4576,N_239);
and U7423 (N_7423,N_4738,N_810);
xnor U7424 (N_7424,N_4212,N_4370);
or U7425 (N_7425,N_493,N_1737);
or U7426 (N_7426,N_964,N_3157);
xnor U7427 (N_7427,N_1952,N_4620);
xnor U7428 (N_7428,N_1997,N_4605);
and U7429 (N_7429,N_3465,N_4825);
xor U7430 (N_7430,N_4391,N_4152);
nand U7431 (N_7431,N_763,N_2555);
nand U7432 (N_7432,N_1759,N_3116);
or U7433 (N_7433,N_1603,N_3808);
nand U7434 (N_7434,N_4346,N_4781);
nand U7435 (N_7435,N_4539,N_4700);
nand U7436 (N_7436,N_4393,N_1221);
and U7437 (N_7437,N_312,N_1255);
nor U7438 (N_7438,N_2134,N_779);
nand U7439 (N_7439,N_2973,N_2182);
and U7440 (N_7440,N_4410,N_2006);
and U7441 (N_7441,N_3628,N_3624);
nand U7442 (N_7442,N_2465,N_4589);
and U7443 (N_7443,N_1371,N_1622);
and U7444 (N_7444,N_2984,N_28);
nor U7445 (N_7445,N_3729,N_2746);
or U7446 (N_7446,N_505,N_2860);
and U7447 (N_7447,N_4185,N_1668);
nor U7448 (N_7448,N_3787,N_1877);
xnor U7449 (N_7449,N_950,N_3972);
or U7450 (N_7450,N_3942,N_3111);
nand U7451 (N_7451,N_369,N_2127);
nor U7452 (N_7452,N_1054,N_4666);
xor U7453 (N_7453,N_758,N_1234);
and U7454 (N_7454,N_2378,N_2874);
nand U7455 (N_7455,N_4030,N_848);
xor U7456 (N_7456,N_2905,N_4599);
nand U7457 (N_7457,N_4769,N_4095);
or U7458 (N_7458,N_4797,N_3095);
nand U7459 (N_7459,N_4622,N_1108);
and U7460 (N_7460,N_4525,N_4833);
and U7461 (N_7461,N_526,N_4703);
nand U7462 (N_7462,N_272,N_2966);
nor U7463 (N_7463,N_3770,N_2708);
and U7464 (N_7464,N_1839,N_2928);
xnor U7465 (N_7465,N_1264,N_757);
or U7466 (N_7466,N_192,N_2090);
or U7467 (N_7467,N_2562,N_1116);
or U7468 (N_7468,N_2395,N_181);
nand U7469 (N_7469,N_2086,N_717);
nand U7470 (N_7470,N_4932,N_3967);
nor U7471 (N_7471,N_137,N_1469);
nor U7472 (N_7472,N_2728,N_3473);
nand U7473 (N_7473,N_4896,N_4313);
or U7474 (N_7474,N_3270,N_3666);
nor U7475 (N_7475,N_2034,N_2953);
or U7476 (N_7476,N_498,N_4570);
and U7477 (N_7477,N_3387,N_2468);
and U7478 (N_7478,N_2900,N_307);
xor U7479 (N_7479,N_2362,N_1650);
xnor U7480 (N_7480,N_3204,N_3626);
or U7481 (N_7481,N_3766,N_4546);
and U7482 (N_7482,N_2301,N_3953);
or U7483 (N_7483,N_2089,N_2777);
nor U7484 (N_7484,N_3576,N_1096);
or U7485 (N_7485,N_3923,N_3197);
xor U7486 (N_7486,N_961,N_932);
nand U7487 (N_7487,N_1042,N_4498);
and U7488 (N_7488,N_485,N_2177);
or U7489 (N_7489,N_3105,N_2883);
or U7490 (N_7490,N_861,N_4613);
nor U7491 (N_7491,N_1496,N_2054);
xor U7492 (N_7492,N_2157,N_2592);
or U7493 (N_7493,N_4849,N_3952);
and U7494 (N_7494,N_1941,N_1416);
nor U7495 (N_7495,N_3494,N_1564);
and U7496 (N_7496,N_658,N_2880);
nand U7497 (N_7497,N_1911,N_4172);
nand U7498 (N_7498,N_4250,N_4418);
xor U7499 (N_7499,N_4166,N_1625);
nor U7500 (N_7500,N_1713,N_586);
xor U7501 (N_7501,N_2348,N_1326);
or U7502 (N_7502,N_330,N_720);
nor U7503 (N_7503,N_1841,N_4064);
nor U7504 (N_7504,N_4360,N_478);
or U7505 (N_7505,N_2761,N_3835);
xor U7506 (N_7506,N_2254,N_2890);
xnor U7507 (N_7507,N_62,N_390);
or U7508 (N_7508,N_2494,N_4643);
and U7509 (N_7509,N_425,N_661);
and U7510 (N_7510,N_937,N_4873);
and U7511 (N_7511,N_428,N_1619);
xnor U7512 (N_7512,N_3672,N_1396);
or U7513 (N_7513,N_1946,N_3217);
and U7514 (N_7514,N_4358,N_2632);
nand U7515 (N_7515,N_2476,N_2960);
and U7516 (N_7516,N_4334,N_3478);
nand U7517 (N_7517,N_4524,N_3384);
or U7518 (N_7518,N_4378,N_3899);
nor U7519 (N_7519,N_4487,N_4159);
xor U7520 (N_7520,N_191,N_4351);
or U7521 (N_7521,N_567,N_1872);
nor U7522 (N_7522,N_1014,N_2018);
nand U7523 (N_7523,N_1517,N_781);
or U7524 (N_7524,N_1540,N_3240);
or U7525 (N_7525,N_1577,N_271);
and U7526 (N_7526,N_1772,N_2605);
xor U7527 (N_7527,N_2118,N_4229);
or U7528 (N_7528,N_2198,N_2952);
and U7529 (N_7529,N_4573,N_1271);
and U7530 (N_7530,N_2773,N_490);
xor U7531 (N_7531,N_2854,N_2627);
xor U7532 (N_7532,N_450,N_1820);
or U7533 (N_7533,N_4315,N_2480);
and U7534 (N_7534,N_4460,N_4323);
xnor U7535 (N_7535,N_2709,N_1216);
and U7536 (N_7536,N_2475,N_632);
xnor U7537 (N_7537,N_4994,N_4223);
xor U7538 (N_7538,N_4228,N_578);
nor U7539 (N_7539,N_1262,N_4738);
nor U7540 (N_7540,N_2953,N_3833);
nor U7541 (N_7541,N_1063,N_3961);
and U7542 (N_7542,N_699,N_3609);
xor U7543 (N_7543,N_590,N_4146);
nor U7544 (N_7544,N_3941,N_354);
xnor U7545 (N_7545,N_1673,N_1939);
nor U7546 (N_7546,N_3027,N_3758);
nor U7547 (N_7547,N_2842,N_3156);
nand U7548 (N_7548,N_1322,N_1838);
xor U7549 (N_7549,N_2299,N_1667);
and U7550 (N_7550,N_3748,N_3289);
or U7551 (N_7551,N_3275,N_1514);
nand U7552 (N_7552,N_2478,N_4001);
and U7553 (N_7553,N_3281,N_2706);
and U7554 (N_7554,N_4047,N_2675);
nand U7555 (N_7555,N_3394,N_3410);
nand U7556 (N_7556,N_2483,N_2702);
nand U7557 (N_7557,N_4643,N_3516);
xnor U7558 (N_7558,N_3327,N_326);
nand U7559 (N_7559,N_4291,N_1059);
nand U7560 (N_7560,N_29,N_4254);
nor U7561 (N_7561,N_2441,N_4797);
or U7562 (N_7562,N_732,N_2453);
xnor U7563 (N_7563,N_162,N_4121);
or U7564 (N_7564,N_1840,N_1935);
xor U7565 (N_7565,N_4498,N_1075);
or U7566 (N_7566,N_2907,N_1897);
and U7567 (N_7567,N_4086,N_4686);
or U7568 (N_7568,N_1646,N_3226);
and U7569 (N_7569,N_4138,N_3520);
or U7570 (N_7570,N_2082,N_3382);
or U7571 (N_7571,N_2594,N_1845);
nor U7572 (N_7572,N_1616,N_3611);
nand U7573 (N_7573,N_1614,N_2070);
xor U7574 (N_7574,N_1960,N_754);
nand U7575 (N_7575,N_2402,N_2972);
nor U7576 (N_7576,N_525,N_1037);
xor U7577 (N_7577,N_1414,N_253);
and U7578 (N_7578,N_3263,N_1834);
or U7579 (N_7579,N_2106,N_229);
or U7580 (N_7580,N_4581,N_85);
xor U7581 (N_7581,N_3173,N_1163);
nand U7582 (N_7582,N_4755,N_1288);
nor U7583 (N_7583,N_1803,N_852);
nand U7584 (N_7584,N_2077,N_1039);
nor U7585 (N_7585,N_1264,N_644);
or U7586 (N_7586,N_3396,N_969);
nand U7587 (N_7587,N_3880,N_336);
and U7588 (N_7588,N_2597,N_312);
or U7589 (N_7589,N_2435,N_4124);
or U7590 (N_7590,N_439,N_3691);
and U7591 (N_7591,N_155,N_1466);
or U7592 (N_7592,N_917,N_349);
nor U7593 (N_7593,N_1221,N_1618);
or U7594 (N_7594,N_3386,N_1972);
nand U7595 (N_7595,N_260,N_332);
nor U7596 (N_7596,N_3131,N_13);
xor U7597 (N_7597,N_3144,N_1329);
or U7598 (N_7598,N_834,N_3851);
nand U7599 (N_7599,N_4894,N_4416);
or U7600 (N_7600,N_1338,N_2856);
xor U7601 (N_7601,N_1578,N_3978);
or U7602 (N_7602,N_95,N_1267);
or U7603 (N_7603,N_550,N_4251);
nor U7604 (N_7604,N_1226,N_2197);
and U7605 (N_7605,N_24,N_1919);
nand U7606 (N_7606,N_4966,N_2302);
xor U7607 (N_7607,N_173,N_969);
or U7608 (N_7608,N_16,N_3546);
nor U7609 (N_7609,N_4515,N_3711);
nand U7610 (N_7610,N_4448,N_3489);
and U7611 (N_7611,N_3588,N_4077);
or U7612 (N_7612,N_3803,N_786);
nor U7613 (N_7613,N_3995,N_152);
nand U7614 (N_7614,N_3553,N_1576);
nor U7615 (N_7615,N_491,N_4349);
or U7616 (N_7616,N_3709,N_738);
nand U7617 (N_7617,N_3475,N_277);
nand U7618 (N_7618,N_4788,N_2509);
xor U7619 (N_7619,N_2315,N_2342);
and U7620 (N_7620,N_2575,N_2040);
and U7621 (N_7621,N_1289,N_4554);
nor U7622 (N_7622,N_2359,N_2444);
xnor U7623 (N_7623,N_2927,N_2922);
nor U7624 (N_7624,N_3417,N_4344);
nor U7625 (N_7625,N_2978,N_1775);
nor U7626 (N_7626,N_4218,N_4127);
nand U7627 (N_7627,N_2043,N_968);
or U7628 (N_7628,N_2129,N_2436);
nor U7629 (N_7629,N_4444,N_2114);
xnor U7630 (N_7630,N_607,N_324);
or U7631 (N_7631,N_4946,N_4669);
or U7632 (N_7632,N_1066,N_2430);
or U7633 (N_7633,N_1442,N_591);
and U7634 (N_7634,N_3618,N_31);
and U7635 (N_7635,N_640,N_3466);
and U7636 (N_7636,N_134,N_102);
nor U7637 (N_7637,N_4952,N_4294);
or U7638 (N_7638,N_1684,N_1359);
nand U7639 (N_7639,N_3880,N_1179);
or U7640 (N_7640,N_4295,N_4895);
nor U7641 (N_7641,N_3375,N_1433);
and U7642 (N_7642,N_586,N_4259);
nor U7643 (N_7643,N_1982,N_3586);
and U7644 (N_7644,N_4367,N_1389);
nand U7645 (N_7645,N_4004,N_620);
nand U7646 (N_7646,N_3225,N_2127);
or U7647 (N_7647,N_4224,N_1866);
nand U7648 (N_7648,N_2858,N_4198);
or U7649 (N_7649,N_1380,N_3281);
nand U7650 (N_7650,N_951,N_1298);
and U7651 (N_7651,N_3421,N_3561);
nor U7652 (N_7652,N_2751,N_2017);
or U7653 (N_7653,N_152,N_2377);
nor U7654 (N_7654,N_3041,N_423);
xor U7655 (N_7655,N_189,N_3122);
and U7656 (N_7656,N_1467,N_4180);
nor U7657 (N_7657,N_4542,N_315);
nand U7658 (N_7658,N_95,N_4076);
nor U7659 (N_7659,N_368,N_778);
nand U7660 (N_7660,N_2507,N_1515);
and U7661 (N_7661,N_1641,N_508);
nor U7662 (N_7662,N_1125,N_4395);
nor U7663 (N_7663,N_2330,N_1200);
or U7664 (N_7664,N_2502,N_3886);
xnor U7665 (N_7665,N_4089,N_96);
nand U7666 (N_7666,N_1615,N_4043);
nor U7667 (N_7667,N_2363,N_1460);
xor U7668 (N_7668,N_1262,N_1012);
nor U7669 (N_7669,N_3942,N_4445);
xor U7670 (N_7670,N_3228,N_1311);
nor U7671 (N_7671,N_2182,N_4391);
nand U7672 (N_7672,N_2131,N_478);
nand U7673 (N_7673,N_2728,N_2882);
nor U7674 (N_7674,N_3706,N_213);
or U7675 (N_7675,N_2490,N_2229);
nand U7676 (N_7676,N_680,N_2092);
nand U7677 (N_7677,N_3357,N_4436);
and U7678 (N_7678,N_3650,N_4983);
and U7679 (N_7679,N_4332,N_2974);
nand U7680 (N_7680,N_912,N_2965);
and U7681 (N_7681,N_3381,N_3827);
nor U7682 (N_7682,N_3949,N_3889);
or U7683 (N_7683,N_2954,N_3317);
nand U7684 (N_7684,N_1555,N_2175);
xnor U7685 (N_7685,N_1951,N_2221);
and U7686 (N_7686,N_1128,N_1166);
nand U7687 (N_7687,N_1896,N_4505);
nor U7688 (N_7688,N_3746,N_2622);
and U7689 (N_7689,N_706,N_4023);
or U7690 (N_7690,N_1078,N_3946);
xnor U7691 (N_7691,N_4403,N_4022);
xnor U7692 (N_7692,N_3775,N_4821);
nor U7693 (N_7693,N_817,N_222);
nor U7694 (N_7694,N_4335,N_144);
nor U7695 (N_7695,N_1057,N_4);
xnor U7696 (N_7696,N_3520,N_4847);
nand U7697 (N_7697,N_1556,N_1541);
nand U7698 (N_7698,N_4392,N_940);
or U7699 (N_7699,N_1539,N_4884);
xnor U7700 (N_7700,N_3530,N_2908);
or U7701 (N_7701,N_620,N_1970);
nor U7702 (N_7702,N_2598,N_918);
nand U7703 (N_7703,N_1740,N_4424);
xor U7704 (N_7704,N_1940,N_1774);
xor U7705 (N_7705,N_3902,N_465);
or U7706 (N_7706,N_2962,N_3564);
nor U7707 (N_7707,N_2813,N_4044);
nand U7708 (N_7708,N_46,N_4484);
and U7709 (N_7709,N_1196,N_743);
nand U7710 (N_7710,N_355,N_230);
or U7711 (N_7711,N_959,N_794);
nor U7712 (N_7712,N_693,N_150);
nand U7713 (N_7713,N_4238,N_1661);
xnor U7714 (N_7714,N_4308,N_3098);
xnor U7715 (N_7715,N_3714,N_588);
or U7716 (N_7716,N_4274,N_996);
nand U7717 (N_7717,N_4332,N_2752);
nor U7718 (N_7718,N_4924,N_354);
nand U7719 (N_7719,N_1462,N_1091);
nor U7720 (N_7720,N_1040,N_2639);
or U7721 (N_7721,N_1126,N_2530);
nand U7722 (N_7722,N_1680,N_1642);
nor U7723 (N_7723,N_449,N_3003);
and U7724 (N_7724,N_96,N_3891);
nand U7725 (N_7725,N_4336,N_4169);
and U7726 (N_7726,N_999,N_1538);
nor U7727 (N_7727,N_2378,N_829);
nand U7728 (N_7728,N_2994,N_3307);
or U7729 (N_7729,N_513,N_4912);
nor U7730 (N_7730,N_4389,N_566);
and U7731 (N_7731,N_4138,N_3921);
nand U7732 (N_7732,N_4682,N_2624);
and U7733 (N_7733,N_406,N_2373);
nand U7734 (N_7734,N_1171,N_3957);
nand U7735 (N_7735,N_1981,N_1474);
nand U7736 (N_7736,N_4224,N_1128);
nor U7737 (N_7737,N_1909,N_4282);
and U7738 (N_7738,N_4200,N_2588);
xnor U7739 (N_7739,N_3059,N_4402);
and U7740 (N_7740,N_2639,N_4507);
or U7741 (N_7741,N_4172,N_175);
xor U7742 (N_7742,N_2628,N_4408);
and U7743 (N_7743,N_3950,N_1897);
and U7744 (N_7744,N_1366,N_3479);
xor U7745 (N_7745,N_3147,N_2555);
and U7746 (N_7746,N_4193,N_3916);
and U7747 (N_7747,N_2813,N_982);
xor U7748 (N_7748,N_121,N_798);
and U7749 (N_7749,N_3813,N_4864);
nor U7750 (N_7750,N_36,N_765);
and U7751 (N_7751,N_4419,N_222);
or U7752 (N_7752,N_833,N_4683);
nor U7753 (N_7753,N_1466,N_3009);
and U7754 (N_7754,N_2894,N_4030);
nor U7755 (N_7755,N_435,N_669);
xor U7756 (N_7756,N_4115,N_2856);
and U7757 (N_7757,N_452,N_483);
nand U7758 (N_7758,N_3445,N_3031);
nor U7759 (N_7759,N_1452,N_1275);
and U7760 (N_7760,N_3925,N_1861);
nand U7761 (N_7761,N_3953,N_3310);
nand U7762 (N_7762,N_4639,N_4932);
nand U7763 (N_7763,N_2516,N_215);
and U7764 (N_7764,N_3014,N_4819);
nand U7765 (N_7765,N_3086,N_3066);
nand U7766 (N_7766,N_1303,N_339);
nand U7767 (N_7767,N_3347,N_4624);
xnor U7768 (N_7768,N_4143,N_4456);
nand U7769 (N_7769,N_3526,N_362);
nor U7770 (N_7770,N_796,N_1051);
and U7771 (N_7771,N_4286,N_1181);
and U7772 (N_7772,N_4699,N_4673);
nand U7773 (N_7773,N_1748,N_4095);
nand U7774 (N_7774,N_2000,N_3103);
and U7775 (N_7775,N_2482,N_3328);
and U7776 (N_7776,N_3738,N_3600);
xnor U7777 (N_7777,N_2204,N_508);
and U7778 (N_7778,N_39,N_2476);
nand U7779 (N_7779,N_3162,N_3343);
and U7780 (N_7780,N_1931,N_2548);
and U7781 (N_7781,N_20,N_2715);
xnor U7782 (N_7782,N_193,N_4003);
nand U7783 (N_7783,N_1343,N_726);
nand U7784 (N_7784,N_3131,N_4993);
or U7785 (N_7785,N_1397,N_1442);
nor U7786 (N_7786,N_2028,N_3243);
and U7787 (N_7787,N_858,N_1056);
or U7788 (N_7788,N_1447,N_1561);
or U7789 (N_7789,N_3159,N_1767);
or U7790 (N_7790,N_3301,N_1481);
and U7791 (N_7791,N_3354,N_1767);
nand U7792 (N_7792,N_4931,N_4131);
and U7793 (N_7793,N_1605,N_225);
nand U7794 (N_7794,N_2906,N_464);
nand U7795 (N_7795,N_799,N_4486);
nand U7796 (N_7796,N_3547,N_973);
or U7797 (N_7797,N_4270,N_4949);
nand U7798 (N_7798,N_2120,N_4287);
and U7799 (N_7799,N_683,N_2796);
or U7800 (N_7800,N_3866,N_855);
xnor U7801 (N_7801,N_2960,N_1026);
or U7802 (N_7802,N_2501,N_1060);
and U7803 (N_7803,N_293,N_1156);
or U7804 (N_7804,N_3300,N_2425);
nand U7805 (N_7805,N_3398,N_2681);
xnor U7806 (N_7806,N_1116,N_2457);
nor U7807 (N_7807,N_631,N_3239);
and U7808 (N_7808,N_4601,N_3541);
or U7809 (N_7809,N_4163,N_3857);
nor U7810 (N_7810,N_715,N_133);
and U7811 (N_7811,N_3376,N_2684);
nor U7812 (N_7812,N_4189,N_4048);
nor U7813 (N_7813,N_4824,N_3644);
or U7814 (N_7814,N_3366,N_3478);
xor U7815 (N_7815,N_2167,N_3789);
nand U7816 (N_7816,N_2133,N_71);
nor U7817 (N_7817,N_4786,N_349);
nor U7818 (N_7818,N_1964,N_1745);
xnor U7819 (N_7819,N_1116,N_2666);
nor U7820 (N_7820,N_3572,N_557);
and U7821 (N_7821,N_417,N_561);
or U7822 (N_7822,N_1343,N_3962);
nand U7823 (N_7823,N_549,N_1311);
nor U7824 (N_7824,N_209,N_3116);
xor U7825 (N_7825,N_730,N_3767);
or U7826 (N_7826,N_4261,N_4768);
xnor U7827 (N_7827,N_1172,N_2588);
nand U7828 (N_7828,N_2738,N_3338);
nor U7829 (N_7829,N_3643,N_3957);
or U7830 (N_7830,N_2482,N_1255);
or U7831 (N_7831,N_2444,N_1330);
nor U7832 (N_7832,N_2287,N_4635);
nand U7833 (N_7833,N_652,N_537);
xor U7834 (N_7834,N_2333,N_153);
nand U7835 (N_7835,N_4347,N_1);
nor U7836 (N_7836,N_4741,N_2820);
nor U7837 (N_7837,N_1765,N_4138);
or U7838 (N_7838,N_1797,N_322);
and U7839 (N_7839,N_2185,N_556);
xor U7840 (N_7840,N_40,N_2724);
and U7841 (N_7841,N_2809,N_2634);
nor U7842 (N_7842,N_4259,N_705);
and U7843 (N_7843,N_4108,N_1615);
and U7844 (N_7844,N_877,N_533);
nor U7845 (N_7845,N_2072,N_1112);
xor U7846 (N_7846,N_3329,N_3853);
and U7847 (N_7847,N_268,N_4035);
or U7848 (N_7848,N_298,N_1493);
or U7849 (N_7849,N_2148,N_1390);
nor U7850 (N_7850,N_1295,N_2699);
or U7851 (N_7851,N_57,N_3791);
nand U7852 (N_7852,N_1619,N_1552);
nor U7853 (N_7853,N_412,N_3994);
and U7854 (N_7854,N_4391,N_4182);
xor U7855 (N_7855,N_4280,N_137);
xnor U7856 (N_7856,N_2855,N_4611);
nand U7857 (N_7857,N_1254,N_4968);
xnor U7858 (N_7858,N_865,N_3579);
or U7859 (N_7859,N_4276,N_2226);
and U7860 (N_7860,N_4580,N_4142);
nor U7861 (N_7861,N_2772,N_337);
xnor U7862 (N_7862,N_3381,N_4648);
or U7863 (N_7863,N_1012,N_3355);
nor U7864 (N_7864,N_724,N_1361);
and U7865 (N_7865,N_4465,N_1664);
xor U7866 (N_7866,N_4606,N_2104);
or U7867 (N_7867,N_3969,N_3619);
and U7868 (N_7868,N_4248,N_4689);
nor U7869 (N_7869,N_1138,N_817);
xnor U7870 (N_7870,N_2544,N_4397);
and U7871 (N_7871,N_2160,N_4067);
nand U7872 (N_7872,N_838,N_108);
nor U7873 (N_7873,N_1753,N_1934);
and U7874 (N_7874,N_2244,N_2691);
xnor U7875 (N_7875,N_1463,N_3577);
and U7876 (N_7876,N_671,N_0);
nand U7877 (N_7877,N_3513,N_4599);
nand U7878 (N_7878,N_4919,N_2439);
or U7879 (N_7879,N_597,N_1356);
and U7880 (N_7880,N_3119,N_616);
xnor U7881 (N_7881,N_4133,N_4786);
and U7882 (N_7882,N_586,N_4593);
nand U7883 (N_7883,N_3335,N_3025);
nor U7884 (N_7884,N_3128,N_4451);
xor U7885 (N_7885,N_3017,N_1464);
nor U7886 (N_7886,N_447,N_4507);
and U7887 (N_7887,N_533,N_3570);
or U7888 (N_7888,N_3506,N_3443);
nor U7889 (N_7889,N_4041,N_4575);
and U7890 (N_7890,N_2670,N_1355);
and U7891 (N_7891,N_2456,N_1506);
xnor U7892 (N_7892,N_4778,N_1407);
nand U7893 (N_7893,N_4889,N_2307);
and U7894 (N_7894,N_3361,N_666);
nor U7895 (N_7895,N_4906,N_1897);
or U7896 (N_7896,N_4629,N_3235);
or U7897 (N_7897,N_1449,N_1040);
and U7898 (N_7898,N_288,N_2706);
nor U7899 (N_7899,N_3939,N_3444);
and U7900 (N_7900,N_719,N_4081);
nand U7901 (N_7901,N_1403,N_3977);
nand U7902 (N_7902,N_1759,N_1784);
xor U7903 (N_7903,N_1216,N_4735);
nor U7904 (N_7904,N_1970,N_4586);
nand U7905 (N_7905,N_564,N_3820);
or U7906 (N_7906,N_3396,N_2544);
xnor U7907 (N_7907,N_3411,N_4356);
or U7908 (N_7908,N_3323,N_2655);
or U7909 (N_7909,N_3352,N_4517);
nor U7910 (N_7910,N_3236,N_459);
or U7911 (N_7911,N_3363,N_3128);
xnor U7912 (N_7912,N_3970,N_4583);
xor U7913 (N_7913,N_4641,N_705);
nand U7914 (N_7914,N_417,N_1859);
nor U7915 (N_7915,N_1048,N_1648);
nor U7916 (N_7916,N_4885,N_2735);
xnor U7917 (N_7917,N_1461,N_4722);
and U7918 (N_7918,N_4857,N_153);
nor U7919 (N_7919,N_2801,N_4222);
nor U7920 (N_7920,N_3191,N_4252);
nor U7921 (N_7921,N_1833,N_2076);
nor U7922 (N_7922,N_3470,N_25);
and U7923 (N_7923,N_567,N_3673);
nand U7924 (N_7924,N_3344,N_3707);
or U7925 (N_7925,N_1490,N_933);
nand U7926 (N_7926,N_1281,N_2200);
or U7927 (N_7927,N_3789,N_251);
nand U7928 (N_7928,N_1657,N_2764);
nand U7929 (N_7929,N_3208,N_866);
xor U7930 (N_7930,N_3853,N_4084);
nand U7931 (N_7931,N_45,N_1657);
xor U7932 (N_7932,N_1831,N_4569);
nand U7933 (N_7933,N_3359,N_733);
and U7934 (N_7934,N_2900,N_4522);
nor U7935 (N_7935,N_2891,N_3217);
xnor U7936 (N_7936,N_1969,N_4030);
or U7937 (N_7937,N_3944,N_2074);
nand U7938 (N_7938,N_1920,N_1279);
xor U7939 (N_7939,N_232,N_4337);
nor U7940 (N_7940,N_1477,N_3990);
nand U7941 (N_7941,N_2311,N_1545);
nand U7942 (N_7942,N_575,N_532);
or U7943 (N_7943,N_2423,N_2039);
and U7944 (N_7944,N_1029,N_2149);
nand U7945 (N_7945,N_390,N_1807);
xnor U7946 (N_7946,N_2322,N_2419);
or U7947 (N_7947,N_996,N_2656);
xor U7948 (N_7948,N_678,N_1564);
nor U7949 (N_7949,N_459,N_4608);
and U7950 (N_7950,N_2743,N_1189);
and U7951 (N_7951,N_782,N_2969);
and U7952 (N_7952,N_2068,N_2035);
and U7953 (N_7953,N_4246,N_106);
or U7954 (N_7954,N_3,N_3578);
xor U7955 (N_7955,N_3278,N_4807);
or U7956 (N_7956,N_69,N_850);
or U7957 (N_7957,N_479,N_4899);
and U7958 (N_7958,N_1877,N_1990);
xor U7959 (N_7959,N_2750,N_943);
and U7960 (N_7960,N_3574,N_4715);
or U7961 (N_7961,N_2574,N_4572);
nor U7962 (N_7962,N_1702,N_4513);
nand U7963 (N_7963,N_4045,N_1310);
or U7964 (N_7964,N_3209,N_663);
nand U7965 (N_7965,N_4424,N_3203);
and U7966 (N_7966,N_3135,N_3383);
nand U7967 (N_7967,N_961,N_1989);
nor U7968 (N_7968,N_3070,N_1392);
nor U7969 (N_7969,N_3300,N_3619);
or U7970 (N_7970,N_1727,N_1406);
nand U7971 (N_7971,N_3912,N_2950);
nor U7972 (N_7972,N_3454,N_4802);
or U7973 (N_7973,N_1296,N_1346);
nand U7974 (N_7974,N_3975,N_4053);
nor U7975 (N_7975,N_143,N_1303);
nor U7976 (N_7976,N_145,N_1712);
or U7977 (N_7977,N_2837,N_983);
or U7978 (N_7978,N_1015,N_3319);
xnor U7979 (N_7979,N_3999,N_4526);
nand U7980 (N_7980,N_534,N_2803);
nor U7981 (N_7981,N_608,N_2876);
xnor U7982 (N_7982,N_4442,N_3433);
and U7983 (N_7983,N_2993,N_1792);
nor U7984 (N_7984,N_3227,N_3869);
xor U7985 (N_7985,N_637,N_4929);
nor U7986 (N_7986,N_445,N_929);
and U7987 (N_7987,N_800,N_1514);
xnor U7988 (N_7988,N_2442,N_4934);
and U7989 (N_7989,N_1861,N_1538);
or U7990 (N_7990,N_1271,N_1641);
and U7991 (N_7991,N_1944,N_3928);
or U7992 (N_7992,N_2739,N_4632);
nor U7993 (N_7993,N_1836,N_2854);
nand U7994 (N_7994,N_252,N_4397);
nor U7995 (N_7995,N_4837,N_2823);
and U7996 (N_7996,N_1412,N_1181);
or U7997 (N_7997,N_1252,N_1478);
and U7998 (N_7998,N_555,N_863);
or U7999 (N_7999,N_1479,N_2092);
nand U8000 (N_8000,N_2947,N_2415);
xnor U8001 (N_8001,N_4295,N_3106);
nor U8002 (N_8002,N_2128,N_881);
or U8003 (N_8003,N_2568,N_652);
or U8004 (N_8004,N_2254,N_1459);
xnor U8005 (N_8005,N_2641,N_4640);
or U8006 (N_8006,N_4229,N_2678);
nand U8007 (N_8007,N_4897,N_3614);
and U8008 (N_8008,N_1940,N_334);
nand U8009 (N_8009,N_3425,N_2227);
nand U8010 (N_8010,N_3122,N_1720);
nand U8011 (N_8011,N_3662,N_2303);
nand U8012 (N_8012,N_2019,N_3964);
xnor U8013 (N_8013,N_4606,N_2867);
or U8014 (N_8014,N_1594,N_4166);
or U8015 (N_8015,N_3904,N_3646);
nor U8016 (N_8016,N_4155,N_2180);
xor U8017 (N_8017,N_1069,N_3770);
and U8018 (N_8018,N_2745,N_2262);
nand U8019 (N_8019,N_805,N_133);
or U8020 (N_8020,N_3393,N_4967);
nand U8021 (N_8021,N_3953,N_4063);
nand U8022 (N_8022,N_3050,N_3063);
xor U8023 (N_8023,N_1378,N_2758);
or U8024 (N_8024,N_2654,N_4414);
xor U8025 (N_8025,N_4635,N_3344);
xnor U8026 (N_8026,N_3835,N_1789);
or U8027 (N_8027,N_1141,N_148);
nand U8028 (N_8028,N_4634,N_833);
xor U8029 (N_8029,N_3213,N_3663);
xnor U8030 (N_8030,N_4558,N_4920);
xnor U8031 (N_8031,N_3426,N_469);
or U8032 (N_8032,N_571,N_2739);
or U8033 (N_8033,N_323,N_3116);
nor U8034 (N_8034,N_4150,N_573);
or U8035 (N_8035,N_2325,N_29);
nand U8036 (N_8036,N_4833,N_3985);
nand U8037 (N_8037,N_4257,N_4858);
nor U8038 (N_8038,N_815,N_2061);
nand U8039 (N_8039,N_3949,N_2914);
nand U8040 (N_8040,N_918,N_4729);
nor U8041 (N_8041,N_2237,N_4824);
nand U8042 (N_8042,N_1224,N_2331);
or U8043 (N_8043,N_2915,N_1853);
or U8044 (N_8044,N_4838,N_3166);
nor U8045 (N_8045,N_3557,N_3742);
or U8046 (N_8046,N_1850,N_3987);
nor U8047 (N_8047,N_4558,N_2883);
nor U8048 (N_8048,N_2317,N_2750);
and U8049 (N_8049,N_1839,N_3444);
nor U8050 (N_8050,N_1301,N_3200);
nor U8051 (N_8051,N_1153,N_2402);
and U8052 (N_8052,N_689,N_2279);
nor U8053 (N_8053,N_4357,N_1731);
xnor U8054 (N_8054,N_295,N_3132);
or U8055 (N_8055,N_4462,N_1338);
nand U8056 (N_8056,N_2161,N_2380);
nand U8057 (N_8057,N_2708,N_2609);
or U8058 (N_8058,N_300,N_1506);
xor U8059 (N_8059,N_1810,N_2379);
and U8060 (N_8060,N_2002,N_3850);
and U8061 (N_8061,N_4933,N_939);
or U8062 (N_8062,N_4862,N_1125);
or U8063 (N_8063,N_921,N_1199);
nand U8064 (N_8064,N_2195,N_222);
nor U8065 (N_8065,N_4322,N_1942);
xnor U8066 (N_8066,N_4558,N_1431);
nand U8067 (N_8067,N_1208,N_3872);
nand U8068 (N_8068,N_2282,N_276);
or U8069 (N_8069,N_204,N_3449);
nor U8070 (N_8070,N_203,N_3664);
or U8071 (N_8071,N_423,N_2459);
xnor U8072 (N_8072,N_1202,N_224);
nor U8073 (N_8073,N_2800,N_1320);
and U8074 (N_8074,N_2199,N_408);
or U8075 (N_8075,N_452,N_3344);
xnor U8076 (N_8076,N_2266,N_105);
nand U8077 (N_8077,N_2985,N_4987);
nor U8078 (N_8078,N_500,N_1088);
xor U8079 (N_8079,N_3298,N_4161);
xor U8080 (N_8080,N_4789,N_2494);
and U8081 (N_8081,N_3352,N_2730);
or U8082 (N_8082,N_4998,N_4825);
xnor U8083 (N_8083,N_1587,N_4897);
nor U8084 (N_8084,N_619,N_3571);
and U8085 (N_8085,N_3882,N_4892);
xor U8086 (N_8086,N_4798,N_1499);
nand U8087 (N_8087,N_491,N_508);
nor U8088 (N_8088,N_1021,N_4289);
nor U8089 (N_8089,N_4988,N_562);
or U8090 (N_8090,N_4478,N_1376);
nand U8091 (N_8091,N_1234,N_3553);
xnor U8092 (N_8092,N_3499,N_1833);
and U8093 (N_8093,N_3828,N_3215);
and U8094 (N_8094,N_1391,N_1639);
nor U8095 (N_8095,N_3503,N_4042);
nand U8096 (N_8096,N_2204,N_4086);
nor U8097 (N_8097,N_4179,N_2208);
xor U8098 (N_8098,N_321,N_208);
xor U8099 (N_8099,N_2536,N_1775);
xnor U8100 (N_8100,N_3359,N_3099);
xnor U8101 (N_8101,N_220,N_2100);
and U8102 (N_8102,N_3423,N_3342);
and U8103 (N_8103,N_781,N_4252);
xor U8104 (N_8104,N_4240,N_3242);
and U8105 (N_8105,N_1466,N_34);
xnor U8106 (N_8106,N_4123,N_4078);
nand U8107 (N_8107,N_969,N_2525);
nand U8108 (N_8108,N_3229,N_2358);
nand U8109 (N_8109,N_2372,N_1067);
and U8110 (N_8110,N_858,N_939);
or U8111 (N_8111,N_3735,N_4496);
nand U8112 (N_8112,N_4203,N_4270);
or U8113 (N_8113,N_1597,N_3370);
nor U8114 (N_8114,N_1626,N_4717);
xor U8115 (N_8115,N_2827,N_428);
and U8116 (N_8116,N_4665,N_2068);
xnor U8117 (N_8117,N_1105,N_1629);
and U8118 (N_8118,N_2359,N_3983);
or U8119 (N_8119,N_3714,N_3530);
or U8120 (N_8120,N_1849,N_3720);
xor U8121 (N_8121,N_3710,N_752);
xnor U8122 (N_8122,N_2746,N_3433);
or U8123 (N_8123,N_4274,N_4986);
and U8124 (N_8124,N_4663,N_287);
nand U8125 (N_8125,N_4148,N_2509);
and U8126 (N_8126,N_2388,N_571);
or U8127 (N_8127,N_108,N_4368);
and U8128 (N_8128,N_215,N_2590);
and U8129 (N_8129,N_1604,N_690);
or U8130 (N_8130,N_3406,N_4863);
and U8131 (N_8131,N_2558,N_37);
nor U8132 (N_8132,N_303,N_1540);
or U8133 (N_8133,N_2895,N_1114);
or U8134 (N_8134,N_1968,N_1224);
xor U8135 (N_8135,N_4306,N_3351);
and U8136 (N_8136,N_4950,N_4655);
or U8137 (N_8137,N_2856,N_4540);
or U8138 (N_8138,N_1199,N_3677);
nand U8139 (N_8139,N_1102,N_1758);
nand U8140 (N_8140,N_3151,N_1675);
and U8141 (N_8141,N_3573,N_2700);
xor U8142 (N_8142,N_4335,N_1501);
and U8143 (N_8143,N_2596,N_1137);
and U8144 (N_8144,N_2322,N_3009);
or U8145 (N_8145,N_3023,N_1158);
xor U8146 (N_8146,N_2681,N_178);
nand U8147 (N_8147,N_4876,N_1071);
xnor U8148 (N_8148,N_4595,N_4752);
nand U8149 (N_8149,N_71,N_372);
nand U8150 (N_8150,N_2364,N_1827);
and U8151 (N_8151,N_3115,N_2270);
or U8152 (N_8152,N_4336,N_3105);
xor U8153 (N_8153,N_2327,N_2498);
nand U8154 (N_8154,N_2228,N_2634);
nand U8155 (N_8155,N_4361,N_2135);
nor U8156 (N_8156,N_2731,N_4806);
nand U8157 (N_8157,N_1392,N_3135);
xor U8158 (N_8158,N_2761,N_3508);
nand U8159 (N_8159,N_3477,N_2826);
xnor U8160 (N_8160,N_3408,N_4328);
and U8161 (N_8161,N_4378,N_4059);
nor U8162 (N_8162,N_3618,N_3532);
and U8163 (N_8163,N_4953,N_1897);
nand U8164 (N_8164,N_2651,N_38);
xnor U8165 (N_8165,N_2186,N_2666);
nand U8166 (N_8166,N_4758,N_4627);
xnor U8167 (N_8167,N_879,N_1860);
or U8168 (N_8168,N_3725,N_52);
nor U8169 (N_8169,N_1918,N_1592);
nor U8170 (N_8170,N_4273,N_623);
and U8171 (N_8171,N_2660,N_553);
or U8172 (N_8172,N_1371,N_2804);
and U8173 (N_8173,N_1537,N_964);
or U8174 (N_8174,N_518,N_1541);
nand U8175 (N_8175,N_1700,N_2914);
xnor U8176 (N_8176,N_1806,N_685);
nor U8177 (N_8177,N_3890,N_2548);
nor U8178 (N_8178,N_2741,N_611);
or U8179 (N_8179,N_3429,N_4276);
or U8180 (N_8180,N_3937,N_864);
or U8181 (N_8181,N_2796,N_4856);
nor U8182 (N_8182,N_4700,N_3136);
or U8183 (N_8183,N_2021,N_831);
nand U8184 (N_8184,N_2213,N_4380);
nor U8185 (N_8185,N_3718,N_361);
nor U8186 (N_8186,N_1074,N_227);
and U8187 (N_8187,N_297,N_4323);
or U8188 (N_8188,N_4337,N_1071);
nor U8189 (N_8189,N_2579,N_4435);
or U8190 (N_8190,N_3195,N_925);
and U8191 (N_8191,N_2998,N_3980);
xnor U8192 (N_8192,N_2520,N_1157);
or U8193 (N_8193,N_803,N_2611);
nor U8194 (N_8194,N_1059,N_4411);
nand U8195 (N_8195,N_3209,N_270);
or U8196 (N_8196,N_3689,N_253);
nand U8197 (N_8197,N_2303,N_1193);
xor U8198 (N_8198,N_2136,N_1079);
or U8199 (N_8199,N_3184,N_525);
nand U8200 (N_8200,N_253,N_2742);
nor U8201 (N_8201,N_4343,N_4465);
and U8202 (N_8202,N_4741,N_1922);
and U8203 (N_8203,N_1516,N_3483);
nand U8204 (N_8204,N_4949,N_19);
nor U8205 (N_8205,N_1743,N_3309);
and U8206 (N_8206,N_329,N_631);
or U8207 (N_8207,N_4544,N_3777);
xor U8208 (N_8208,N_607,N_512);
xor U8209 (N_8209,N_4290,N_9);
nand U8210 (N_8210,N_3451,N_941);
and U8211 (N_8211,N_955,N_3896);
nand U8212 (N_8212,N_1088,N_4918);
or U8213 (N_8213,N_3389,N_4059);
nor U8214 (N_8214,N_1245,N_3717);
nand U8215 (N_8215,N_2177,N_2350);
nand U8216 (N_8216,N_1215,N_4956);
or U8217 (N_8217,N_4254,N_4405);
nand U8218 (N_8218,N_4906,N_353);
nor U8219 (N_8219,N_3873,N_2324);
nor U8220 (N_8220,N_2923,N_1534);
or U8221 (N_8221,N_820,N_2467);
or U8222 (N_8222,N_3290,N_1453);
or U8223 (N_8223,N_4442,N_4054);
xnor U8224 (N_8224,N_3364,N_1568);
nor U8225 (N_8225,N_999,N_3443);
and U8226 (N_8226,N_2531,N_3606);
nand U8227 (N_8227,N_211,N_2410);
and U8228 (N_8228,N_1010,N_4867);
or U8229 (N_8229,N_1449,N_3177);
and U8230 (N_8230,N_2458,N_1565);
xnor U8231 (N_8231,N_1926,N_1149);
and U8232 (N_8232,N_1057,N_3668);
nor U8233 (N_8233,N_818,N_1676);
nor U8234 (N_8234,N_4352,N_1735);
xnor U8235 (N_8235,N_155,N_4769);
or U8236 (N_8236,N_4925,N_4550);
and U8237 (N_8237,N_3648,N_2721);
or U8238 (N_8238,N_446,N_4950);
nand U8239 (N_8239,N_978,N_1811);
nor U8240 (N_8240,N_2361,N_3978);
xor U8241 (N_8241,N_509,N_4169);
or U8242 (N_8242,N_4430,N_1324);
and U8243 (N_8243,N_465,N_3873);
xor U8244 (N_8244,N_2603,N_2604);
or U8245 (N_8245,N_392,N_791);
nor U8246 (N_8246,N_1660,N_631);
nor U8247 (N_8247,N_4045,N_4462);
or U8248 (N_8248,N_2448,N_3937);
or U8249 (N_8249,N_4608,N_377);
xnor U8250 (N_8250,N_4326,N_4403);
nor U8251 (N_8251,N_3457,N_43);
or U8252 (N_8252,N_565,N_632);
or U8253 (N_8253,N_2826,N_748);
xor U8254 (N_8254,N_4022,N_2491);
nand U8255 (N_8255,N_3466,N_3209);
xnor U8256 (N_8256,N_3964,N_1180);
xnor U8257 (N_8257,N_216,N_3492);
xnor U8258 (N_8258,N_2154,N_393);
nor U8259 (N_8259,N_3138,N_494);
nand U8260 (N_8260,N_656,N_185);
nand U8261 (N_8261,N_809,N_2730);
nor U8262 (N_8262,N_3282,N_2715);
xor U8263 (N_8263,N_1376,N_868);
and U8264 (N_8264,N_1702,N_4471);
or U8265 (N_8265,N_3776,N_2107);
xor U8266 (N_8266,N_4251,N_1752);
or U8267 (N_8267,N_3671,N_1942);
or U8268 (N_8268,N_1476,N_380);
nand U8269 (N_8269,N_2984,N_1802);
xor U8270 (N_8270,N_4805,N_4984);
nand U8271 (N_8271,N_4156,N_4032);
nor U8272 (N_8272,N_560,N_831);
nand U8273 (N_8273,N_2162,N_1765);
and U8274 (N_8274,N_4883,N_3622);
or U8275 (N_8275,N_3223,N_1651);
xnor U8276 (N_8276,N_4492,N_3409);
and U8277 (N_8277,N_1145,N_4966);
xnor U8278 (N_8278,N_66,N_1925);
or U8279 (N_8279,N_2856,N_4074);
or U8280 (N_8280,N_589,N_4456);
and U8281 (N_8281,N_676,N_912);
and U8282 (N_8282,N_2166,N_2528);
nor U8283 (N_8283,N_1372,N_1153);
nor U8284 (N_8284,N_4831,N_1021);
or U8285 (N_8285,N_2214,N_3608);
xnor U8286 (N_8286,N_2827,N_2098);
nor U8287 (N_8287,N_202,N_1185);
nand U8288 (N_8288,N_3255,N_1304);
and U8289 (N_8289,N_2453,N_4886);
nor U8290 (N_8290,N_3568,N_942);
xnor U8291 (N_8291,N_2607,N_2231);
or U8292 (N_8292,N_2475,N_3245);
xor U8293 (N_8293,N_3735,N_2083);
or U8294 (N_8294,N_2161,N_2088);
nand U8295 (N_8295,N_3992,N_3530);
nand U8296 (N_8296,N_3469,N_2228);
nand U8297 (N_8297,N_3074,N_2996);
or U8298 (N_8298,N_4134,N_678);
and U8299 (N_8299,N_3348,N_373);
or U8300 (N_8300,N_3707,N_628);
nand U8301 (N_8301,N_3262,N_3735);
nand U8302 (N_8302,N_4336,N_1668);
nor U8303 (N_8303,N_2894,N_1547);
xnor U8304 (N_8304,N_3622,N_1061);
and U8305 (N_8305,N_3404,N_3849);
nand U8306 (N_8306,N_4724,N_4498);
or U8307 (N_8307,N_4808,N_468);
xor U8308 (N_8308,N_2538,N_1718);
nand U8309 (N_8309,N_4744,N_11);
and U8310 (N_8310,N_4755,N_3973);
xor U8311 (N_8311,N_4188,N_3108);
or U8312 (N_8312,N_164,N_4647);
nand U8313 (N_8313,N_4993,N_468);
nor U8314 (N_8314,N_2316,N_2318);
xor U8315 (N_8315,N_4422,N_3155);
and U8316 (N_8316,N_1825,N_1749);
xnor U8317 (N_8317,N_1321,N_2504);
nor U8318 (N_8318,N_738,N_2862);
nand U8319 (N_8319,N_3293,N_3679);
xnor U8320 (N_8320,N_3972,N_1176);
nand U8321 (N_8321,N_1401,N_967);
and U8322 (N_8322,N_944,N_1800);
and U8323 (N_8323,N_1682,N_1607);
nand U8324 (N_8324,N_1375,N_4038);
or U8325 (N_8325,N_4885,N_4750);
xor U8326 (N_8326,N_4522,N_1199);
or U8327 (N_8327,N_4527,N_225);
nand U8328 (N_8328,N_94,N_3399);
or U8329 (N_8329,N_4220,N_1563);
and U8330 (N_8330,N_944,N_756);
nor U8331 (N_8331,N_4036,N_1254);
and U8332 (N_8332,N_1396,N_1045);
nand U8333 (N_8333,N_4107,N_793);
or U8334 (N_8334,N_376,N_1575);
or U8335 (N_8335,N_4999,N_747);
nand U8336 (N_8336,N_4348,N_2261);
and U8337 (N_8337,N_2345,N_1921);
and U8338 (N_8338,N_2860,N_630);
and U8339 (N_8339,N_214,N_990);
xor U8340 (N_8340,N_1149,N_77);
xnor U8341 (N_8341,N_2280,N_684);
and U8342 (N_8342,N_1262,N_4410);
or U8343 (N_8343,N_1468,N_1857);
nor U8344 (N_8344,N_2177,N_2380);
xor U8345 (N_8345,N_4620,N_1030);
nand U8346 (N_8346,N_2066,N_4765);
and U8347 (N_8347,N_4970,N_3515);
or U8348 (N_8348,N_4054,N_4796);
or U8349 (N_8349,N_1918,N_241);
nor U8350 (N_8350,N_3477,N_4377);
xnor U8351 (N_8351,N_3163,N_1004);
nand U8352 (N_8352,N_1410,N_4766);
nand U8353 (N_8353,N_3825,N_2988);
and U8354 (N_8354,N_2161,N_1670);
xnor U8355 (N_8355,N_3064,N_4522);
nand U8356 (N_8356,N_2820,N_127);
nand U8357 (N_8357,N_3187,N_3775);
and U8358 (N_8358,N_3088,N_3158);
nor U8359 (N_8359,N_313,N_2883);
xor U8360 (N_8360,N_1725,N_1382);
and U8361 (N_8361,N_4034,N_3310);
or U8362 (N_8362,N_2227,N_629);
nor U8363 (N_8363,N_4508,N_3794);
or U8364 (N_8364,N_4932,N_753);
xor U8365 (N_8365,N_636,N_4819);
nand U8366 (N_8366,N_1258,N_4011);
and U8367 (N_8367,N_2131,N_540);
or U8368 (N_8368,N_4305,N_4209);
or U8369 (N_8369,N_4780,N_1168);
and U8370 (N_8370,N_3917,N_4390);
or U8371 (N_8371,N_2004,N_2567);
and U8372 (N_8372,N_4735,N_2942);
or U8373 (N_8373,N_4993,N_4764);
and U8374 (N_8374,N_1633,N_4439);
or U8375 (N_8375,N_1274,N_3796);
nor U8376 (N_8376,N_3454,N_2233);
and U8377 (N_8377,N_3894,N_3215);
and U8378 (N_8378,N_4944,N_1757);
nor U8379 (N_8379,N_4521,N_1154);
nand U8380 (N_8380,N_1184,N_161);
xnor U8381 (N_8381,N_482,N_491);
nor U8382 (N_8382,N_2542,N_3148);
nand U8383 (N_8383,N_3213,N_3050);
nand U8384 (N_8384,N_1852,N_3637);
or U8385 (N_8385,N_3144,N_1800);
nand U8386 (N_8386,N_3579,N_1839);
nand U8387 (N_8387,N_3227,N_172);
xnor U8388 (N_8388,N_2870,N_1781);
and U8389 (N_8389,N_4528,N_942);
nor U8390 (N_8390,N_3158,N_1391);
nor U8391 (N_8391,N_3614,N_1339);
nor U8392 (N_8392,N_665,N_2410);
xor U8393 (N_8393,N_2323,N_2654);
nand U8394 (N_8394,N_2698,N_3293);
nand U8395 (N_8395,N_4194,N_213);
or U8396 (N_8396,N_1720,N_1651);
nand U8397 (N_8397,N_2629,N_2619);
and U8398 (N_8398,N_726,N_520);
and U8399 (N_8399,N_4013,N_3870);
nor U8400 (N_8400,N_1681,N_957);
or U8401 (N_8401,N_2881,N_278);
or U8402 (N_8402,N_3176,N_3677);
and U8403 (N_8403,N_750,N_1055);
or U8404 (N_8404,N_356,N_3131);
xor U8405 (N_8405,N_1287,N_941);
nor U8406 (N_8406,N_903,N_4762);
nor U8407 (N_8407,N_2344,N_210);
nor U8408 (N_8408,N_3787,N_3336);
and U8409 (N_8409,N_1236,N_1831);
xnor U8410 (N_8410,N_2860,N_667);
nor U8411 (N_8411,N_4186,N_4396);
and U8412 (N_8412,N_1697,N_2628);
xnor U8413 (N_8413,N_2752,N_3873);
nor U8414 (N_8414,N_3767,N_1886);
nor U8415 (N_8415,N_2016,N_87);
xor U8416 (N_8416,N_1346,N_1149);
xnor U8417 (N_8417,N_3883,N_4038);
nor U8418 (N_8418,N_2344,N_4799);
or U8419 (N_8419,N_2422,N_4871);
and U8420 (N_8420,N_1270,N_4357);
nand U8421 (N_8421,N_3078,N_4084);
nor U8422 (N_8422,N_1971,N_2897);
nor U8423 (N_8423,N_3735,N_1555);
nand U8424 (N_8424,N_1902,N_1179);
nand U8425 (N_8425,N_1482,N_4688);
nand U8426 (N_8426,N_2189,N_915);
nor U8427 (N_8427,N_9,N_2704);
and U8428 (N_8428,N_2209,N_367);
and U8429 (N_8429,N_1155,N_1531);
or U8430 (N_8430,N_37,N_3909);
or U8431 (N_8431,N_3064,N_424);
and U8432 (N_8432,N_4793,N_1071);
nor U8433 (N_8433,N_4055,N_167);
or U8434 (N_8434,N_4443,N_3536);
and U8435 (N_8435,N_3639,N_2379);
nand U8436 (N_8436,N_3535,N_105);
nand U8437 (N_8437,N_942,N_4979);
nor U8438 (N_8438,N_479,N_4384);
or U8439 (N_8439,N_4572,N_2530);
xnor U8440 (N_8440,N_3002,N_3464);
nor U8441 (N_8441,N_1890,N_1639);
xor U8442 (N_8442,N_3940,N_3353);
or U8443 (N_8443,N_4477,N_286);
nor U8444 (N_8444,N_2999,N_3957);
xnor U8445 (N_8445,N_51,N_2765);
and U8446 (N_8446,N_4083,N_1877);
or U8447 (N_8447,N_61,N_3459);
nand U8448 (N_8448,N_1632,N_3338);
or U8449 (N_8449,N_30,N_4535);
nand U8450 (N_8450,N_4199,N_2976);
nand U8451 (N_8451,N_1412,N_4272);
nor U8452 (N_8452,N_2536,N_396);
nand U8453 (N_8453,N_3013,N_3201);
and U8454 (N_8454,N_776,N_4860);
and U8455 (N_8455,N_428,N_1267);
nand U8456 (N_8456,N_2154,N_4756);
xnor U8457 (N_8457,N_514,N_2364);
xnor U8458 (N_8458,N_3546,N_2036);
xor U8459 (N_8459,N_4130,N_3575);
nand U8460 (N_8460,N_3766,N_1308);
nor U8461 (N_8461,N_3372,N_1170);
or U8462 (N_8462,N_3519,N_1921);
nand U8463 (N_8463,N_1890,N_4224);
or U8464 (N_8464,N_3161,N_4650);
or U8465 (N_8465,N_4957,N_1835);
xnor U8466 (N_8466,N_2594,N_727);
and U8467 (N_8467,N_4735,N_3166);
xor U8468 (N_8468,N_2044,N_3212);
nor U8469 (N_8469,N_4853,N_1090);
nand U8470 (N_8470,N_1054,N_3838);
nor U8471 (N_8471,N_725,N_4769);
nor U8472 (N_8472,N_2582,N_972);
and U8473 (N_8473,N_1363,N_2798);
xnor U8474 (N_8474,N_732,N_4542);
and U8475 (N_8475,N_4340,N_2744);
and U8476 (N_8476,N_4334,N_1218);
nor U8477 (N_8477,N_3982,N_3344);
and U8478 (N_8478,N_3994,N_2517);
and U8479 (N_8479,N_2512,N_1992);
and U8480 (N_8480,N_179,N_1522);
or U8481 (N_8481,N_4386,N_663);
xnor U8482 (N_8482,N_4606,N_2630);
or U8483 (N_8483,N_214,N_2898);
or U8484 (N_8484,N_3263,N_3777);
or U8485 (N_8485,N_4476,N_113);
or U8486 (N_8486,N_4400,N_1243);
and U8487 (N_8487,N_2985,N_706);
and U8488 (N_8488,N_3079,N_3909);
and U8489 (N_8489,N_513,N_4552);
or U8490 (N_8490,N_2565,N_4498);
nor U8491 (N_8491,N_2117,N_4285);
and U8492 (N_8492,N_2027,N_109);
and U8493 (N_8493,N_4571,N_375);
or U8494 (N_8494,N_259,N_2538);
nand U8495 (N_8495,N_3187,N_1460);
nor U8496 (N_8496,N_2616,N_72);
and U8497 (N_8497,N_3709,N_3235);
and U8498 (N_8498,N_3693,N_1430);
nand U8499 (N_8499,N_506,N_3956);
xnor U8500 (N_8500,N_1967,N_971);
nor U8501 (N_8501,N_3293,N_4447);
nor U8502 (N_8502,N_1001,N_4843);
or U8503 (N_8503,N_715,N_3882);
nor U8504 (N_8504,N_2041,N_764);
and U8505 (N_8505,N_684,N_1003);
or U8506 (N_8506,N_1533,N_3080);
xor U8507 (N_8507,N_531,N_2463);
and U8508 (N_8508,N_81,N_3953);
nand U8509 (N_8509,N_2264,N_3525);
xor U8510 (N_8510,N_3143,N_2878);
nor U8511 (N_8511,N_4323,N_222);
and U8512 (N_8512,N_3654,N_658);
or U8513 (N_8513,N_2823,N_1734);
or U8514 (N_8514,N_2139,N_830);
nand U8515 (N_8515,N_1921,N_3441);
nor U8516 (N_8516,N_3792,N_2936);
nand U8517 (N_8517,N_2659,N_4117);
xor U8518 (N_8518,N_3044,N_1589);
or U8519 (N_8519,N_1524,N_1392);
nor U8520 (N_8520,N_3531,N_1747);
xnor U8521 (N_8521,N_669,N_4233);
or U8522 (N_8522,N_1010,N_2801);
nand U8523 (N_8523,N_1798,N_3097);
xnor U8524 (N_8524,N_4337,N_1737);
and U8525 (N_8525,N_2074,N_2803);
nor U8526 (N_8526,N_1520,N_2239);
nor U8527 (N_8527,N_4271,N_4727);
or U8528 (N_8528,N_3258,N_4515);
or U8529 (N_8529,N_3244,N_2664);
nor U8530 (N_8530,N_1416,N_2104);
and U8531 (N_8531,N_1917,N_735);
nor U8532 (N_8532,N_241,N_1028);
and U8533 (N_8533,N_3984,N_302);
or U8534 (N_8534,N_4754,N_1038);
xor U8535 (N_8535,N_2388,N_2757);
xor U8536 (N_8536,N_312,N_1318);
xnor U8537 (N_8537,N_3358,N_2714);
or U8538 (N_8538,N_991,N_90);
or U8539 (N_8539,N_139,N_2218);
or U8540 (N_8540,N_3424,N_1498);
and U8541 (N_8541,N_3902,N_4090);
xnor U8542 (N_8542,N_197,N_2743);
nor U8543 (N_8543,N_1158,N_1819);
xor U8544 (N_8544,N_697,N_1282);
xor U8545 (N_8545,N_2892,N_456);
xor U8546 (N_8546,N_2534,N_640);
xor U8547 (N_8547,N_4681,N_1611);
xnor U8548 (N_8548,N_747,N_2380);
nand U8549 (N_8549,N_4055,N_3411);
xor U8550 (N_8550,N_817,N_2932);
nor U8551 (N_8551,N_3267,N_1358);
and U8552 (N_8552,N_2220,N_1491);
nor U8553 (N_8553,N_892,N_1435);
nor U8554 (N_8554,N_457,N_3501);
nand U8555 (N_8555,N_705,N_1279);
xor U8556 (N_8556,N_4376,N_874);
nand U8557 (N_8557,N_902,N_4168);
xor U8558 (N_8558,N_1980,N_3481);
nor U8559 (N_8559,N_4153,N_1161);
nand U8560 (N_8560,N_2151,N_1472);
nand U8561 (N_8561,N_1346,N_2687);
and U8562 (N_8562,N_3372,N_2807);
nor U8563 (N_8563,N_3272,N_1882);
xnor U8564 (N_8564,N_2692,N_2351);
xnor U8565 (N_8565,N_303,N_2473);
or U8566 (N_8566,N_543,N_126);
nor U8567 (N_8567,N_758,N_114);
nand U8568 (N_8568,N_672,N_4848);
nor U8569 (N_8569,N_2765,N_3431);
nor U8570 (N_8570,N_3609,N_2422);
or U8571 (N_8571,N_3752,N_1434);
nor U8572 (N_8572,N_1013,N_798);
and U8573 (N_8573,N_2083,N_4970);
or U8574 (N_8574,N_994,N_3483);
nor U8575 (N_8575,N_2143,N_3405);
and U8576 (N_8576,N_3790,N_3976);
nor U8577 (N_8577,N_2023,N_2436);
xnor U8578 (N_8578,N_3696,N_4684);
nand U8579 (N_8579,N_3850,N_1451);
or U8580 (N_8580,N_1940,N_4434);
or U8581 (N_8581,N_4252,N_2936);
nand U8582 (N_8582,N_1509,N_4398);
xor U8583 (N_8583,N_4129,N_2829);
nand U8584 (N_8584,N_4964,N_2046);
nand U8585 (N_8585,N_176,N_4234);
and U8586 (N_8586,N_2191,N_1202);
and U8587 (N_8587,N_1561,N_4129);
or U8588 (N_8588,N_4679,N_2750);
or U8589 (N_8589,N_204,N_3335);
and U8590 (N_8590,N_4550,N_375);
or U8591 (N_8591,N_1406,N_3807);
xor U8592 (N_8592,N_1228,N_3209);
and U8593 (N_8593,N_1161,N_217);
nand U8594 (N_8594,N_942,N_3454);
and U8595 (N_8595,N_4512,N_3488);
or U8596 (N_8596,N_4951,N_4395);
nor U8597 (N_8597,N_4373,N_1831);
or U8598 (N_8598,N_1802,N_856);
and U8599 (N_8599,N_4520,N_1014);
and U8600 (N_8600,N_3836,N_1649);
and U8601 (N_8601,N_4713,N_3044);
nor U8602 (N_8602,N_1341,N_2154);
and U8603 (N_8603,N_2863,N_3846);
xor U8604 (N_8604,N_1714,N_1549);
xnor U8605 (N_8605,N_2849,N_3925);
or U8606 (N_8606,N_3528,N_1745);
nand U8607 (N_8607,N_2907,N_2331);
or U8608 (N_8608,N_193,N_2672);
and U8609 (N_8609,N_4967,N_4245);
nor U8610 (N_8610,N_3118,N_3149);
and U8611 (N_8611,N_3941,N_1889);
and U8612 (N_8612,N_4506,N_2020);
or U8613 (N_8613,N_3700,N_2429);
xnor U8614 (N_8614,N_1170,N_3782);
and U8615 (N_8615,N_4562,N_935);
nor U8616 (N_8616,N_4685,N_3687);
xnor U8617 (N_8617,N_4164,N_597);
and U8618 (N_8618,N_116,N_4928);
xor U8619 (N_8619,N_3492,N_3410);
or U8620 (N_8620,N_531,N_881);
nand U8621 (N_8621,N_594,N_129);
xor U8622 (N_8622,N_235,N_111);
nor U8623 (N_8623,N_4557,N_1191);
or U8624 (N_8624,N_3669,N_2671);
and U8625 (N_8625,N_4421,N_1552);
nand U8626 (N_8626,N_3841,N_3852);
nor U8627 (N_8627,N_3275,N_2161);
or U8628 (N_8628,N_743,N_2847);
xor U8629 (N_8629,N_2230,N_1270);
xnor U8630 (N_8630,N_2634,N_3012);
nor U8631 (N_8631,N_1298,N_1839);
and U8632 (N_8632,N_863,N_580);
or U8633 (N_8633,N_4656,N_2065);
or U8634 (N_8634,N_2256,N_2135);
nor U8635 (N_8635,N_1414,N_3033);
or U8636 (N_8636,N_1064,N_671);
nand U8637 (N_8637,N_683,N_4147);
and U8638 (N_8638,N_536,N_3187);
and U8639 (N_8639,N_2662,N_2234);
xor U8640 (N_8640,N_4202,N_3891);
nand U8641 (N_8641,N_4196,N_3613);
or U8642 (N_8642,N_3698,N_53);
nor U8643 (N_8643,N_358,N_538);
xor U8644 (N_8644,N_3445,N_3114);
or U8645 (N_8645,N_4341,N_2482);
xnor U8646 (N_8646,N_4342,N_4469);
nand U8647 (N_8647,N_2955,N_3930);
nor U8648 (N_8648,N_4220,N_4614);
or U8649 (N_8649,N_2916,N_4544);
xnor U8650 (N_8650,N_1673,N_339);
or U8651 (N_8651,N_3338,N_1093);
xnor U8652 (N_8652,N_4923,N_658);
or U8653 (N_8653,N_3078,N_3734);
or U8654 (N_8654,N_2031,N_2640);
nor U8655 (N_8655,N_1566,N_717);
or U8656 (N_8656,N_256,N_2027);
or U8657 (N_8657,N_1348,N_3429);
nand U8658 (N_8658,N_1542,N_4349);
nor U8659 (N_8659,N_406,N_4445);
nand U8660 (N_8660,N_498,N_850);
and U8661 (N_8661,N_563,N_4014);
xor U8662 (N_8662,N_3204,N_3917);
xor U8663 (N_8663,N_1902,N_524);
nand U8664 (N_8664,N_813,N_3147);
nand U8665 (N_8665,N_4396,N_3623);
and U8666 (N_8666,N_4165,N_2124);
and U8667 (N_8667,N_4851,N_3722);
nand U8668 (N_8668,N_761,N_324);
xnor U8669 (N_8669,N_2597,N_1138);
nand U8670 (N_8670,N_2525,N_2818);
and U8671 (N_8671,N_1795,N_912);
and U8672 (N_8672,N_1356,N_312);
xor U8673 (N_8673,N_2088,N_4591);
nand U8674 (N_8674,N_1634,N_112);
nand U8675 (N_8675,N_4473,N_1563);
nand U8676 (N_8676,N_4303,N_3869);
and U8677 (N_8677,N_1557,N_4335);
nand U8678 (N_8678,N_3256,N_4291);
nor U8679 (N_8679,N_2880,N_1075);
nor U8680 (N_8680,N_4501,N_4601);
nand U8681 (N_8681,N_758,N_2267);
nor U8682 (N_8682,N_2092,N_2786);
nor U8683 (N_8683,N_1768,N_1644);
xnor U8684 (N_8684,N_2560,N_187);
xor U8685 (N_8685,N_2175,N_289);
xnor U8686 (N_8686,N_2870,N_3512);
nor U8687 (N_8687,N_2828,N_2291);
or U8688 (N_8688,N_381,N_2323);
nor U8689 (N_8689,N_698,N_1795);
nor U8690 (N_8690,N_2495,N_2546);
nand U8691 (N_8691,N_4110,N_345);
nand U8692 (N_8692,N_307,N_2484);
nor U8693 (N_8693,N_1920,N_4268);
and U8694 (N_8694,N_1790,N_1800);
nor U8695 (N_8695,N_3643,N_18);
and U8696 (N_8696,N_81,N_2880);
and U8697 (N_8697,N_4853,N_1533);
or U8698 (N_8698,N_1657,N_2438);
nand U8699 (N_8699,N_3654,N_2738);
and U8700 (N_8700,N_1866,N_1894);
nor U8701 (N_8701,N_3391,N_2274);
or U8702 (N_8702,N_4999,N_3180);
nand U8703 (N_8703,N_2199,N_195);
or U8704 (N_8704,N_1442,N_2050);
xnor U8705 (N_8705,N_418,N_3197);
and U8706 (N_8706,N_1127,N_642);
xor U8707 (N_8707,N_451,N_4183);
and U8708 (N_8708,N_2876,N_3880);
and U8709 (N_8709,N_392,N_3191);
xnor U8710 (N_8710,N_2467,N_3773);
or U8711 (N_8711,N_249,N_4632);
nor U8712 (N_8712,N_1080,N_1508);
and U8713 (N_8713,N_4975,N_212);
xor U8714 (N_8714,N_3863,N_216);
nor U8715 (N_8715,N_1685,N_4185);
or U8716 (N_8716,N_2706,N_512);
xnor U8717 (N_8717,N_3146,N_2977);
nor U8718 (N_8718,N_2410,N_1761);
and U8719 (N_8719,N_3118,N_477);
xor U8720 (N_8720,N_1162,N_4349);
or U8721 (N_8721,N_1996,N_4578);
nor U8722 (N_8722,N_1160,N_2425);
xor U8723 (N_8723,N_3318,N_4111);
or U8724 (N_8724,N_1764,N_1637);
nor U8725 (N_8725,N_4498,N_1329);
and U8726 (N_8726,N_4247,N_4161);
xnor U8727 (N_8727,N_4277,N_3202);
and U8728 (N_8728,N_4263,N_1049);
nor U8729 (N_8729,N_1369,N_4325);
xor U8730 (N_8730,N_3771,N_701);
and U8731 (N_8731,N_3062,N_1708);
nand U8732 (N_8732,N_4979,N_3422);
nor U8733 (N_8733,N_4717,N_3928);
nor U8734 (N_8734,N_1573,N_4078);
and U8735 (N_8735,N_4177,N_1874);
or U8736 (N_8736,N_4787,N_4664);
or U8737 (N_8737,N_2266,N_3103);
nand U8738 (N_8738,N_1709,N_2160);
nand U8739 (N_8739,N_3530,N_417);
and U8740 (N_8740,N_1870,N_2654);
nand U8741 (N_8741,N_3362,N_4120);
nor U8742 (N_8742,N_2152,N_4805);
xnor U8743 (N_8743,N_3970,N_1452);
xor U8744 (N_8744,N_3816,N_478);
xor U8745 (N_8745,N_1174,N_785);
nand U8746 (N_8746,N_4095,N_2874);
xnor U8747 (N_8747,N_4180,N_3049);
and U8748 (N_8748,N_4036,N_4178);
nor U8749 (N_8749,N_1940,N_3258);
and U8750 (N_8750,N_3383,N_1045);
xnor U8751 (N_8751,N_94,N_308);
nand U8752 (N_8752,N_1801,N_3185);
xor U8753 (N_8753,N_3371,N_10);
xnor U8754 (N_8754,N_2544,N_315);
or U8755 (N_8755,N_3839,N_306);
xor U8756 (N_8756,N_1572,N_961);
and U8757 (N_8757,N_4386,N_4362);
nand U8758 (N_8758,N_1328,N_2991);
nor U8759 (N_8759,N_910,N_938);
and U8760 (N_8760,N_1583,N_4700);
nor U8761 (N_8761,N_3200,N_2052);
nand U8762 (N_8762,N_2310,N_4237);
or U8763 (N_8763,N_3363,N_1621);
nor U8764 (N_8764,N_4438,N_198);
nand U8765 (N_8765,N_703,N_3903);
and U8766 (N_8766,N_1953,N_1704);
xnor U8767 (N_8767,N_1244,N_1319);
xor U8768 (N_8768,N_2451,N_3390);
nand U8769 (N_8769,N_4422,N_3962);
and U8770 (N_8770,N_4751,N_4367);
or U8771 (N_8771,N_1106,N_3937);
and U8772 (N_8772,N_4987,N_3336);
nand U8773 (N_8773,N_1848,N_4204);
or U8774 (N_8774,N_1328,N_363);
and U8775 (N_8775,N_1724,N_1522);
nor U8776 (N_8776,N_4779,N_3771);
and U8777 (N_8777,N_1124,N_1445);
or U8778 (N_8778,N_3403,N_1936);
or U8779 (N_8779,N_3000,N_269);
nand U8780 (N_8780,N_405,N_3737);
xor U8781 (N_8781,N_378,N_639);
nand U8782 (N_8782,N_1101,N_1157);
nor U8783 (N_8783,N_206,N_1408);
and U8784 (N_8784,N_4840,N_605);
nand U8785 (N_8785,N_3654,N_1549);
or U8786 (N_8786,N_3800,N_3650);
nor U8787 (N_8787,N_4,N_893);
nand U8788 (N_8788,N_2289,N_3755);
or U8789 (N_8789,N_341,N_2773);
nand U8790 (N_8790,N_1023,N_1669);
nand U8791 (N_8791,N_1127,N_864);
xor U8792 (N_8792,N_2056,N_3695);
nor U8793 (N_8793,N_1595,N_1448);
nor U8794 (N_8794,N_1634,N_3903);
nor U8795 (N_8795,N_4163,N_829);
xor U8796 (N_8796,N_206,N_1931);
and U8797 (N_8797,N_2402,N_4483);
nor U8798 (N_8798,N_3032,N_4479);
nor U8799 (N_8799,N_58,N_2159);
nand U8800 (N_8800,N_2311,N_2693);
or U8801 (N_8801,N_3917,N_4201);
nor U8802 (N_8802,N_3309,N_2640);
nor U8803 (N_8803,N_1349,N_3338);
xor U8804 (N_8804,N_372,N_3894);
or U8805 (N_8805,N_3121,N_3440);
xnor U8806 (N_8806,N_272,N_774);
or U8807 (N_8807,N_3593,N_1939);
nand U8808 (N_8808,N_4957,N_4555);
xor U8809 (N_8809,N_379,N_775);
nor U8810 (N_8810,N_2603,N_3559);
xnor U8811 (N_8811,N_3143,N_4652);
or U8812 (N_8812,N_3448,N_3276);
or U8813 (N_8813,N_3246,N_900);
nor U8814 (N_8814,N_1859,N_85);
or U8815 (N_8815,N_4125,N_3045);
xnor U8816 (N_8816,N_247,N_1451);
nand U8817 (N_8817,N_2259,N_3000);
nand U8818 (N_8818,N_405,N_3501);
xnor U8819 (N_8819,N_2345,N_2891);
or U8820 (N_8820,N_1330,N_2391);
or U8821 (N_8821,N_2619,N_2585);
nor U8822 (N_8822,N_2595,N_4599);
nor U8823 (N_8823,N_1782,N_4814);
or U8824 (N_8824,N_1830,N_4728);
nor U8825 (N_8825,N_3881,N_1466);
or U8826 (N_8826,N_957,N_2726);
or U8827 (N_8827,N_4104,N_2920);
and U8828 (N_8828,N_4793,N_2350);
nand U8829 (N_8829,N_459,N_473);
xor U8830 (N_8830,N_4145,N_770);
nand U8831 (N_8831,N_2098,N_3673);
xor U8832 (N_8832,N_1329,N_66);
or U8833 (N_8833,N_2081,N_1580);
nand U8834 (N_8834,N_3181,N_3049);
nand U8835 (N_8835,N_2100,N_1359);
or U8836 (N_8836,N_4786,N_4434);
xor U8837 (N_8837,N_1757,N_2806);
nand U8838 (N_8838,N_3094,N_230);
and U8839 (N_8839,N_1875,N_4689);
nor U8840 (N_8840,N_4695,N_1316);
nor U8841 (N_8841,N_4592,N_3086);
or U8842 (N_8842,N_2899,N_637);
or U8843 (N_8843,N_3074,N_3430);
nand U8844 (N_8844,N_1366,N_4481);
nor U8845 (N_8845,N_4493,N_794);
nor U8846 (N_8846,N_3480,N_1623);
xor U8847 (N_8847,N_2981,N_4248);
nand U8848 (N_8848,N_4262,N_985);
nand U8849 (N_8849,N_1307,N_4501);
xnor U8850 (N_8850,N_3525,N_3573);
and U8851 (N_8851,N_3390,N_1320);
nor U8852 (N_8852,N_42,N_2041);
or U8853 (N_8853,N_2293,N_4250);
nor U8854 (N_8854,N_3565,N_4111);
nand U8855 (N_8855,N_3229,N_2245);
nor U8856 (N_8856,N_545,N_1519);
nand U8857 (N_8857,N_1920,N_2179);
or U8858 (N_8858,N_1648,N_1895);
or U8859 (N_8859,N_1043,N_4724);
and U8860 (N_8860,N_2826,N_4722);
xor U8861 (N_8861,N_735,N_469);
xnor U8862 (N_8862,N_4547,N_2169);
nor U8863 (N_8863,N_3519,N_3788);
xnor U8864 (N_8864,N_4124,N_1759);
xnor U8865 (N_8865,N_3924,N_3011);
or U8866 (N_8866,N_2748,N_3212);
xor U8867 (N_8867,N_4522,N_3743);
or U8868 (N_8868,N_793,N_3605);
nand U8869 (N_8869,N_3896,N_432);
xor U8870 (N_8870,N_4562,N_2006);
xor U8871 (N_8871,N_1109,N_732);
or U8872 (N_8872,N_2242,N_4191);
nand U8873 (N_8873,N_4230,N_335);
nand U8874 (N_8874,N_1222,N_632);
nand U8875 (N_8875,N_828,N_423);
or U8876 (N_8876,N_2609,N_2302);
nor U8877 (N_8877,N_773,N_2290);
xor U8878 (N_8878,N_4216,N_1925);
xnor U8879 (N_8879,N_524,N_3664);
xor U8880 (N_8880,N_3594,N_4136);
nor U8881 (N_8881,N_3514,N_1183);
nand U8882 (N_8882,N_2695,N_3973);
nor U8883 (N_8883,N_795,N_2451);
nor U8884 (N_8884,N_4381,N_1084);
and U8885 (N_8885,N_4171,N_1303);
or U8886 (N_8886,N_3335,N_3666);
or U8887 (N_8887,N_2375,N_984);
nor U8888 (N_8888,N_2846,N_4526);
or U8889 (N_8889,N_1606,N_3327);
xnor U8890 (N_8890,N_3164,N_1629);
nand U8891 (N_8891,N_2459,N_4138);
nor U8892 (N_8892,N_4903,N_22);
nor U8893 (N_8893,N_1797,N_2305);
xnor U8894 (N_8894,N_3930,N_3931);
and U8895 (N_8895,N_250,N_3469);
and U8896 (N_8896,N_149,N_4392);
and U8897 (N_8897,N_4256,N_3481);
and U8898 (N_8898,N_387,N_1595);
nor U8899 (N_8899,N_246,N_4524);
nand U8900 (N_8900,N_2030,N_1166);
and U8901 (N_8901,N_4564,N_4690);
nand U8902 (N_8902,N_4907,N_4139);
or U8903 (N_8903,N_3324,N_842);
xnor U8904 (N_8904,N_2229,N_3363);
nor U8905 (N_8905,N_4808,N_4719);
nand U8906 (N_8906,N_833,N_2424);
xnor U8907 (N_8907,N_3978,N_291);
or U8908 (N_8908,N_1995,N_1775);
xnor U8909 (N_8909,N_440,N_2791);
nand U8910 (N_8910,N_825,N_1144);
and U8911 (N_8911,N_2979,N_2175);
nand U8912 (N_8912,N_2111,N_2205);
nand U8913 (N_8913,N_3728,N_4152);
nand U8914 (N_8914,N_2202,N_2920);
and U8915 (N_8915,N_1670,N_755);
or U8916 (N_8916,N_3969,N_1094);
xnor U8917 (N_8917,N_3029,N_4306);
and U8918 (N_8918,N_3242,N_3093);
nor U8919 (N_8919,N_4653,N_4710);
nor U8920 (N_8920,N_1963,N_516);
or U8921 (N_8921,N_2412,N_1101);
and U8922 (N_8922,N_933,N_3705);
and U8923 (N_8923,N_2075,N_280);
xnor U8924 (N_8924,N_112,N_2174);
xnor U8925 (N_8925,N_3421,N_645);
and U8926 (N_8926,N_4396,N_2512);
xor U8927 (N_8927,N_2320,N_4706);
or U8928 (N_8928,N_109,N_1588);
and U8929 (N_8929,N_1341,N_1692);
and U8930 (N_8930,N_2943,N_3895);
xnor U8931 (N_8931,N_1870,N_4254);
xnor U8932 (N_8932,N_2514,N_3462);
or U8933 (N_8933,N_1530,N_2692);
or U8934 (N_8934,N_4916,N_3057);
and U8935 (N_8935,N_4648,N_74);
or U8936 (N_8936,N_3975,N_902);
xor U8937 (N_8937,N_2454,N_855);
xor U8938 (N_8938,N_2798,N_238);
xnor U8939 (N_8939,N_2633,N_2139);
nand U8940 (N_8940,N_4695,N_770);
and U8941 (N_8941,N_1987,N_742);
nand U8942 (N_8942,N_541,N_2254);
or U8943 (N_8943,N_2449,N_1215);
or U8944 (N_8944,N_3519,N_1532);
or U8945 (N_8945,N_3315,N_3719);
xnor U8946 (N_8946,N_1671,N_644);
xnor U8947 (N_8947,N_1047,N_1687);
or U8948 (N_8948,N_3484,N_2009);
or U8949 (N_8949,N_2793,N_1871);
nand U8950 (N_8950,N_2963,N_4932);
xor U8951 (N_8951,N_2575,N_4264);
xor U8952 (N_8952,N_3795,N_1350);
and U8953 (N_8953,N_3889,N_2641);
or U8954 (N_8954,N_4853,N_4111);
nor U8955 (N_8955,N_796,N_1949);
nand U8956 (N_8956,N_4675,N_3982);
nand U8957 (N_8957,N_3993,N_2206);
or U8958 (N_8958,N_187,N_305);
nor U8959 (N_8959,N_3539,N_4101);
or U8960 (N_8960,N_233,N_4758);
or U8961 (N_8961,N_4049,N_1788);
nor U8962 (N_8962,N_2461,N_2213);
nor U8963 (N_8963,N_3356,N_3590);
nor U8964 (N_8964,N_4766,N_4114);
xnor U8965 (N_8965,N_3964,N_1652);
xnor U8966 (N_8966,N_3514,N_4169);
and U8967 (N_8967,N_4412,N_3946);
xnor U8968 (N_8968,N_1625,N_247);
xor U8969 (N_8969,N_2091,N_974);
nor U8970 (N_8970,N_2547,N_4870);
nand U8971 (N_8971,N_391,N_4982);
nand U8972 (N_8972,N_370,N_2842);
xnor U8973 (N_8973,N_3816,N_2905);
nand U8974 (N_8974,N_4399,N_333);
nand U8975 (N_8975,N_1853,N_3098);
xor U8976 (N_8976,N_1751,N_124);
nand U8977 (N_8977,N_1706,N_890);
or U8978 (N_8978,N_370,N_2063);
nor U8979 (N_8979,N_3247,N_971);
nor U8980 (N_8980,N_1446,N_2984);
nor U8981 (N_8981,N_3777,N_4656);
xor U8982 (N_8982,N_4102,N_2730);
nand U8983 (N_8983,N_3,N_445);
and U8984 (N_8984,N_879,N_4254);
or U8985 (N_8985,N_2340,N_1868);
nand U8986 (N_8986,N_4233,N_3081);
xor U8987 (N_8987,N_2061,N_3592);
nand U8988 (N_8988,N_892,N_4491);
or U8989 (N_8989,N_4257,N_3954);
or U8990 (N_8990,N_3288,N_4971);
and U8991 (N_8991,N_4221,N_1880);
or U8992 (N_8992,N_59,N_2160);
xnor U8993 (N_8993,N_4487,N_3083);
nor U8994 (N_8994,N_3125,N_355);
nand U8995 (N_8995,N_357,N_3202);
nor U8996 (N_8996,N_4524,N_4714);
and U8997 (N_8997,N_1785,N_3141);
and U8998 (N_8998,N_3609,N_1406);
or U8999 (N_8999,N_1859,N_2196);
nand U9000 (N_9000,N_219,N_3354);
nand U9001 (N_9001,N_1572,N_3889);
nor U9002 (N_9002,N_4579,N_3869);
nand U9003 (N_9003,N_4613,N_1107);
nand U9004 (N_9004,N_2136,N_1338);
and U9005 (N_9005,N_730,N_3677);
and U9006 (N_9006,N_386,N_3833);
and U9007 (N_9007,N_2246,N_2165);
or U9008 (N_9008,N_1873,N_945);
or U9009 (N_9009,N_2360,N_735);
xor U9010 (N_9010,N_1533,N_2371);
nor U9011 (N_9011,N_3843,N_1305);
and U9012 (N_9012,N_2678,N_2626);
and U9013 (N_9013,N_2858,N_4212);
nand U9014 (N_9014,N_479,N_4846);
and U9015 (N_9015,N_1861,N_3889);
nand U9016 (N_9016,N_4254,N_1720);
nor U9017 (N_9017,N_2123,N_2540);
and U9018 (N_9018,N_1952,N_4145);
nor U9019 (N_9019,N_850,N_825);
nand U9020 (N_9020,N_1070,N_1252);
nand U9021 (N_9021,N_1129,N_1724);
nand U9022 (N_9022,N_3736,N_991);
and U9023 (N_9023,N_560,N_859);
and U9024 (N_9024,N_1502,N_962);
or U9025 (N_9025,N_1770,N_4541);
or U9026 (N_9026,N_4643,N_4956);
or U9027 (N_9027,N_2686,N_260);
nor U9028 (N_9028,N_2748,N_292);
nand U9029 (N_9029,N_4507,N_741);
nand U9030 (N_9030,N_433,N_1312);
nand U9031 (N_9031,N_3532,N_1606);
nand U9032 (N_9032,N_4032,N_151);
or U9033 (N_9033,N_2967,N_3273);
or U9034 (N_9034,N_2172,N_4731);
nor U9035 (N_9035,N_2719,N_1496);
xnor U9036 (N_9036,N_4700,N_732);
or U9037 (N_9037,N_3045,N_4695);
nor U9038 (N_9038,N_937,N_3301);
nor U9039 (N_9039,N_2710,N_866);
and U9040 (N_9040,N_3905,N_4064);
xor U9041 (N_9041,N_4685,N_1286);
xor U9042 (N_9042,N_386,N_1209);
nand U9043 (N_9043,N_2358,N_3603);
nand U9044 (N_9044,N_1982,N_2922);
and U9045 (N_9045,N_3725,N_210);
nor U9046 (N_9046,N_3695,N_2086);
or U9047 (N_9047,N_1994,N_1233);
or U9048 (N_9048,N_3741,N_620);
nor U9049 (N_9049,N_63,N_1499);
xor U9050 (N_9050,N_2263,N_2893);
or U9051 (N_9051,N_2192,N_2971);
xor U9052 (N_9052,N_403,N_4786);
and U9053 (N_9053,N_1853,N_3267);
and U9054 (N_9054,N_4138,N_2775);
or U9055 (N_9055,N_2777,N_521);
or U9056 (N_9056,N_3674,N_4918);
or U9057 (N_9057,N_1238,N_2833);
or U9058 (N_9058,N_2384,N_198);
and U9059 (N_9059,N_848,N_1433);
nand U9060 (N_9060,N_320,N_3456);
or U9061 (N_9061,N_1993,N_4115);
nor U9062 (N_9062,N_4275,N_4041);
or U9063 (N_9063,N_1525,N_3115);
nor U9064 (N_9064,N_1385,N_1609);
or U9065 (N_9065,N_2324,N_1738);
nand U9066 (N_9066,N_5,N_1285);
xnor U9067 (N_9067,N_3425,N_3196);
and U9068 (N_9068,N_837,N_2447);
or U9069 (N_9069,N_924,N_3566);
nor U9070 (N_9070,N_4634,N_2773);
xnor U9071 (N_9071,N_4719,N_4817);
and U9072 (N_9072,N_1122,N_1813);
or U9073 (N_9073,N_4786,N_3768);
xnor U9074 (N_9074,N_4706,N_1703);
and U9075 (N_9075,N_3353,N_3230);
and U9076 (N_9076,N_3335,N_4067);
nand U9077 (N_9077,N_4978,N_1921);
or U9078 (N_9078,N_1546,N_2982);
and U9079 (N_9079,N_3224,N_4817);
and U9080 (N_9080,N_2453,N_341);
and U9081 (N_9081,N_3737,N_248);
nor U9082 (N_9082,N_3625,N_4164);
nor U9083 (N_9083,N_3704,N_2019);
xnor U9084 (N_9084,N_2411,N_4715);
nand U9085 (N_9085,N_1306,N_218);
nor U9086 (N_9086,N_2586,N_1369);
and U9087 (N_9087,N_3039,N_4287);
or U9088 (N_9088,N_2764,N_2590);
or U9089 (N_9089,N_1445,N_3659);
nand U9090 (N_9090,N_3254,N_4062);
nor U9091 (N_9091,N_3634,N_124);
xor U9092 (N_9092,N_897,N_2852);
nand U9093 (N_9093,N_555,N_432);
nand U9094 (N_9094,N_1923,N_2009);
or U9095 (N_9095,N_4098,N_2824);
xor U9096 (N_9096,N_4627,N_3671);
or U9097 (N_9097,N_1077,N_1182);
xnor U9098 (N_9098,N_4718,N_1359);
nand U9099 (N_9099,N_3932,N_2734);
and U9100 (N_9100,N_1923,N_4396);
xor U9101 (N_9101,N_4058,N_896);
nor U9102 (N_9102,N_2378,N_3052);
or U9103 (N_9103,N_2454,N_1401);
or U9104 (N_9104,N_1919,N_3414);
xnor U9105 (N_9105,N_693,N_3090);
or U9106 (N_9106,N_4783,N_2233);
nor U9107 (N_9107,N_3301,N_962);
nor U9108 (N_9108,N_4514,N_1066);
or U9109 (N_9109,N_2433,N_2290);
and U9110 (N_9110,N_439,N_4636);
nand U9111 (N_9111,N_2202,N_4904);
and U9112 (N_9112,N_4014,N_2339);
nor U9113 (N_9113,N_2495,N_2455);
nand U9114 (N_9114,N_4832,N_3610);
nor U9115 (N_9115,N_4854,N_100);
or U9116 (N_9116,N_2030,N_4729);
nand U9117 (N_9117,N_3525,N_136);
nor U9118 (N_9118,N_3913,N_2725);
nor U9119 (N_9119,N_2743,N_3308);
xor U9120 (N_9120,N_3590,N_4206);
and U9121 (N_9121,N_1788,N_3640);
or U9122 (N_9122,N_3023,N_2969);
xnor U9123 (N_9123,N_1724,N_2191);
nor U9124 (N_9124,N_3595,N_2260);
and U9125 (N_9125,N_3634,N_4307);
or U9126 (N_9126,N_879,N_3308);
nand U9127 (N_9127,N_705,N_1613);
xor U9128 (N_9128,N_3284,N_4201);
nand U9129 (N_9129,N_2216,N_4773);
nor U9130 (N_9130,N_1810,N_3897);
xor U9131 (N_9131,N_2938,N_3614);
nand U9132 (N_9132,N_1875,N_4477);
nand U9133 (N_9133,N_433,N_3379);
xnor U9134 (N_9134,N_3031,N_170);
xor U9135 (N_9135,N_1025,N_549);
and U9136 (N_9136,N_4409,N_3898);
nor U9137 (N_9137,N_338,N_295);
or U9138 (N_9138,N_1666,N_4551);
xnor U9139 (N_9139,N_1233,N_4379);
nor U9140 (N_9140,N_4320,N_2931);
or U9141 (N_9141,N_4340,N_3890);
nand U9142 (N_9142,N_3774,N_4575);
nor U9143 (N_9143,N_4643,N_4229);
and U9144 (N_9144,N_4333,N_2609);
xnor U9145 (N_9145,N_4423,N_2584);
xnor U9146 (N_9146,N_1607,N_4409);
nor U9147 (N_9147,N_4145,N_4160);
nand U9148 (N_9148,N_222,N_1734);
nor U9149 (N_9149,N_89,N_2348);
and U9150 (N_9150,N_1940,N_4588);
nand U9151 (N_9151,N_723,N_3);
or U9152 (N_9152,N_4078,N_1374);
nand U9153 (N_9153,N_377,N_634);
xor U9154 (N_9154,N_3301,N_2509);
nor U9155 (N_9155,N_3218,N_2711);
and U9156 (N_9156,N_194,N_2279);
nand U9157 (N_9157,N_4530,N_1124);
and U9158 (N_9158,N_2278,N_2934);
xnor U9159 (N_9159,N_2247,N_2104);
xnor U9160 (N_9160,N_4408,N_2315);
xor U9161 (N_9161,N_738,N_2552);
nor U9162 (N_9162,N_452,N_562);
and U9163 (N_9163,N_2969,N_181);
or U9164 (N_9164,N_4105,N_4368);
xor U9165 (N_9165,N_1551,N_468);
nor U9166 (N_9166,N_541,N_2236);
nor U9167 (N_9167,N_3487,N_4930);
nand U9168 (N_9168,N_1585,N_1350);
and U9169 (N_9169,N_4515,N_2859);
or U9170 (N_9170,N_2674,N_2285);
nand U9171 (N_9171,N_2058,N_2649);
nand U9172 (N_9172,N_480,N_813);
and U9173 (N_9173,N_4432,N_988);
or U9174 (N_9174,N_1390,N_2079);
nand U9175 (N_9175,N_4212,N_1201);
xnor U9176 (N_9176,N_654,N_4795);
xnor U9177 (N_9177,N_1916,N_3351);
nand U9178 (N_9178,N_2598,N_4098);
xnor U9179 (N_9179,N_4487,N_4665);
nand U9180 (N_9180,N_1945,N_4993);
nor U9181 (N_9181,N_2559,N_3006);
or U9182 (N_9182,N_4538,N_1923);
xnor U9183 (N_9183,N_4145,N_1355);
and U9184 (N_9184,N_300,N_2761);
nor U9185 (N_9185,N_351,N_4944);
nor U9186 (N_9186,N_903,N_4152);
and U9187 (N_9187,N_2011,N_4570);
nor U9188 (N_9188,N_942,N_1941);
or U9189 (N_9189,N_1039,N_4689);
and U9190 (N_9190,N_1912,N_4648);
xor U9191 (N_9191,N_4084,N_3446);
nand U9192 (N_9192,N_3178,N_2305);
xor U9193 (N_9193,N_4425,N_4771);
nor U9194 (N_9194,N_770,N_3958);
nor U9195 (N_9195,N_3330,N_1806);
nor U9196 (N_9196,N_1105,N_3051);
nor U9197 (N_9197,N_4482,N_2667);
or U9198 (N_9198,N_1607,N_2189);
xor U9199 (N_9199,N_4362,N_2340);
or U9200 (N_9200,N_1750,N_4145);
or U9201 (N_9201,N_2630,N_1129);
or U9202 (N_9202,N_3746,N_2302);
nand U9203 (N_9203,N_335,N_1377);
and U9204 (N_9204,N_2637,N_2762);
nor U9205 (N_9205,N_2186,N_4257);
or U9206 (N_9206,N_844,N_4318);
and U9207 (N_9207,N_4314,N_4195);
and U9208 (N_9208,N_1662,N_3111);
or U9209 (N_9209,N_3530,N_1598);
nand U9210 (N_9210,N_4276,N_4175);
or U9211 (N_9211,N_2883,N_1507);
nor U9212 (N_9212,N_1217,N_3323);
or U9213 (N_9213,N_2341,N_129);
and U9214 (N_9214,N_1115,N_3087);
and U9215 (N_9215,N_396,N_2162);
nor U9216 (N_9216,N_2500,N_3704);
xor U9217 (N_9217,N_4485,N_4728);
nor U9218 (N_9218,N_900,N_4817);
nor U9219 (N_9219,N_4133,N_793);
nand U9220 (N_9220,N_1668,N_4533);
or U9221 (N_9221,N_470,N_1366);
or U9222 (N_9222,N_2307,N_1250);
xnor U9223 (N_9223,N_3875,N_4971);
nor U9224 (N_9224,N_1840,N_2046);
or U9225 (N_9225,N_4449,N_3231);
nor U9226 (N_9226,N_4519,N_2036);
nor U9227 (N_9227,N_3465,N_1522);
and U9228 (N_9228,N_3101,N_252);
nand U9229 (N_9229,N_2624,N_3685);
nand U9230 (N_9230,N_3184,N_2945);
nor U9231 (N_9231,N_3380,N_2207);
or U9232 (N_9232,N_848,N_3141);
nor U9233 (N_9233,N_1965,N_3001);
or U9234 (N_9234,N_4590,N_1778);
or U9235 (N_9235,N_1143,N_4891);
or U9236 (N_9236,N_2571,N_728);
and U9237 (N_9237,N_4794,N_4765);
and U9238 (N_9238,N_1696,N_3418);
nor U9239 (N_9239,N_2379,N_1196);
xor U9240 (N_9240,N_4501,N_1985);
and U9241 (N_9241,N_2616,N_3623);
nand U9242 (N_9242,N_2601,N_952);
xnor U9243 (N_9243,N_2044,N_2965);
nand U9244 (N_9244,N_4595,N_3003);
xnor U9245 (N_9245,N_1463,N_1642);
or U9246 (N_9246,N_1662,N_3821);
or U9247 (N_9247,N_2679,N_4681);
nand U9248 (N_9248,N_3716,N_4238);
or U9249 (N_9249,N_4957,N_1596);
nand U9250 (N_9250,N_2379,N_679);
or U9251 (N_9251,N_4928,N_4643);
nand U9252 (N_9252,N_1959,N_2127);
and U9253 (N_9253,N_4073,N_3407);
xnor U9254 (N_9254,N_1892,N_1738);
xnor U9255 (N_9255,N_1153,N_2164);
and U9256 (N_9256,N_3926,N_3766);
and U9257 (N_9257,N_490,N_33);
or U9258 (N_9258,N_4309,N_4637);
xnor U9259 (N_9259,N_2383,N_3883);
or U9260 (N_9260,N_1784,N_326);
nor U9261 (N_9261,N_1330,N_4430);
or U9262 (N_9262,N_4281,N_1143);
nand U9263 (N_9263,N_709,N_382);
nand U9264 (N_9264,N_4573,N_28);
nor U9265 (N_9265,N_2995,N_1690);
nand U9266 (N_9266,N_1527,N_3109);
nor U9267 (N_9267,N_1945,N_4522);
xnor U9268 (N_9268,N_4836,N_880);
nor U9269 (N_9269,N_1940,N_4487);
or U9270 (N_9270,N_2951,N_2035);
and U9271 (N_9271,N_4408,N_2470);
nor U9272 (N_9272,N_4440,N_1688);
xnor U9273 (N_9273,N_4097,N_2631);
nand U9274 (N_9274,N_1913,N_1771);
and U9275 (N_9275,N_2750,N_1736);
and U9276 (N_9276,N_1905,N_3455);
and U9277 (N_9277,N_2103,N_4478);
nor U9278 (N_9278,N_3884,N_3257);
nand U9279 (N_9279,N_4876,N_4062);
nor U9280 (N_9280,N_183,N_3658);
and U9281 (N_9281,N_1817,N_1318);
nor U9282 (N_9282,N_1447,N_65);
xor U9283 (N_9283,N_1724,N_1056);
or U9284 (N_9284,N_1280,N_1982);
or U9285 (N_9285,N_723,N_1579);
nand U9286 (N_9286,N_79,N_2919);
and U9287 (N_9287,N_141,N_3262);
nor U9288 (N_9288,N_2227,N_591);
or U9289 (N_9289,N_3009,N_3270);
and U9290 (N_9290,N_1848,N_4478);
nand U9291 (N_9291,N_4833,N_629);
and U9292 (N_9292,N_3413,N_4422);
nand U9293 (N_9293,N_174,N_2914);
and U9294 (N_9294,N_174,N_4553);
and U9295 (N_9295,N_2272,N_1191);
and U9296 (N_9296,N_4672,N_4470);
nor U9297 (N_9297,N_492,N_823);
and U9298 (N_9298,N_4311,N_1414);
xnor U9299 (N_9299,N_2673,N_2663);
and U9300 (N_9300,N_1018,N_2223);
and U9301 (N_9301,N_577,N_782);
nor U9302 (N_9302,N_1695,N_3049);
and U9303 (N_9303,N_1887,N_3240);
nor U9304 (N_9304,N_4274,N_3229);
and U9305 (N_9305,N_2821,N_3363);
and U9306 (N_9306,N_2148,N_2547);
xnor U9307 (N_9307,N_1119,N_4502);
nand U9308 (N_9308,N_3080,N_4389);
nor U9309 (N_9309,N_4444,N_988);
and U9310 (N_9310,N_3303,N_979);
and U9311 (N_9311,N_4175,N_2242);
nand U9312 (N_9312,N_2210,N_967);
and U9313 (N_9313,N_3368,N_4141);
nand U9314 (N_9314,N_3501,N_3858);
xor U9315 (N_9315,N_3362,N_4981);
nand U9316 (N_9316,N_4499,N_3229);
nor U9317 (N_9317,N_4895,N_3290);
or U9318 (N_9318,N_834,N_704);
nand U9319 (N_9319,N_2027,N_44);
nand U9320 (N_9320,N_4678,N_2937);
nand U9321 (N_9321,N_2290,N_1981);
xor U9322 (N_9322,N_1168,N_1985);
nand U9323 (N_9323,N_4341,N_183);
nand U9324 (N_9324,N_366,N_3882);
and U9325 (N_9325,N_4648,N_4436);
and U9326 (N_9326,N_807,N_2127);
nor U9327 (N_9327,N_1587,N_468);
nand U9328 (N_9328,N_628,N_4326);
xor U9329 (N_9329,N_2302,N_1691);
xnor U9330 (N_9330,N_179,N_1721);
and U9331 (N_9331,N_2597,N_4946);
nand U9332 (N_9332,N_1407,N_2296);
xnor U9333 (N_9333,N_2491,N_882);
nor U9334 (N_9334,N_4827,N_1444);
xnor U9335 (N_9335,N_3790,N_3012);
nand U9336 (N_9336,N_4983,N_2030);
or U9337 (N_9337,N_1475,N_634);
or U9338 (N_9338,N_3638,N_4527);
nor U9339 (N_9339,N_3821,N_927);
and U9340 (N_9340,N_3313,N_4676);
nand U9341 (N_9341,N_2194,N_3389);
xnor U9342 (N_9342,N_2897,N_1198);
or U9343 (N_9343,N_4156,N_439);
and U9344 (N_9344,N_1563,N_3721);
nor U9345 (N_9345,N_1487,N_829);
xor U9346 (N_9346,N_715,N_1277);
nor U9347 (N_9347,N_437,N_1670);
and U9348 (N_9348,N_2307,N_1766);
xor U9349 (N_9349,N_2111,N_3982);
and U9350 (N_9350,N_956,N_2597);
nand U9351 (N_9351,N_725,N_4036);
nor U9352 (N_9352,N_1363,N_1068);
xor U9353 (N_9353,N_2395,N_1607);
nor U9354 (N_9354,N_2441,N_1265);
or U9355 (N_9355,N_2802,N_3337);
or U9356 (N_9356,N_4397,N_4437);
xor U9357 (N_9357,N_1423,N_3221);
and U9358 (N_9358,N_2568,N_1649);
or U9359 (N_9359,N_826,N_2554);
xor U9360 (N_9360,N_4561,N_1981);
or U9361 (N_9361,N_991,N_2662);
xor U9362 (N_9362,N_3170,N_4235);
or U9363 (N_9363,N_488,N_4467);
nand U9364 (N_9364,N_3219,N_3333);
xnor U9365 (N_9365,N_1030,N_689);
or U9366 (N_9366,N_1697,N_1503);
or U9367 (N_9367,N_720,N_196);
xor U9368 (N_9368,N_4611,N_1883);
nor U9369 (N_9369,N_3554,N_1045);
nand U9370 (N_9370,N_4908,N_1263);
and U9371 (N_9371,N_3308,N_1436);
and U9372 (N_9372,N_3590,N_2384);
xnor U9373 (N_9373,N_1992,N_1322);
or U9374 (N_9374,N_4484,N_2780);
and U9375 (N_9375,N_596,N_1592);
nand U9376 (N_9376,N_2501,N_1020);
and U9377 (N_9377,N_2189,N_21);
xnor U9378 (N_9378,N_433,N_1236);
nand U9379 (N_9379,N_2488,N_2175);
and U9380 (N_9380,N_2608,N_1236);
nand U9381 (N_9381,N_2934,N_2832);
or U9382 (N_9382,N_4145,N_3685);
and U9383 (N_9383,N_3488,N_1484);
xor U9384 (N_9384,N_582,N_4279);
xnor U9385 (N_9385,N_2960,N_4881);
xor U9386 (N_9386,N_4304,N_2255);
and U9387 (N_9387,N_262,N_1939);
nand U9388 (N_9388,N_539,N_1104);
and U9389 (N_9389,N_3038,N_4739);
xor U9390 (N_9390,N_2326,N_2015);
xnor U9391 (N_9391,N_3091,N_4584);
or U9392 (N_9392,N_3337,N_4052);
xor U9393 (N_9393,N_2706,N_3108);
nor U9394 (N_9394,N_2136,N_2815);
nand U9395 (N_9395,N_2249,N_4053);
nor U9396 (N_9396,N_3380,N_644);
and U9397 (N_9397,N_188,N_3762);
nor U9398 (N_9398,N_3678,N_3390);
and U9399 (N_9399,N_987,N_1817);
nor U9400 (N_9400,N_2635,N_3869);
nor U9401 (N_9401,N_210,N_4338);
xor U9402 (N_9402,N_2401,N_2010);
and U9403 (N_9403,N_2129,N_589);
nor U9404 (N_9404,N_622,N_4366);
xor U9405 (N_9405,N_38,N_1912);
nor U9406 (N_9406,N_1027,N_827);
nor U9407 (N_9407,N_3488,N_2484);
xnor U9408 (N_9408,N_4130,N_3782);
xnor U9409 (N_9409,N_2918,N_3625);
xnor U9410 (N_9410,N_4758,N_2916);
nand U9411 (N_9411,N_3696,N_2237);
nor U9412 (N_9412,N_558,N_74);
xnor U9413 (N_9413,N_2240,N_1307);
nand U9414 (N_9414,N_1208,N_753);
xnor U9415 (N_9415,N_11,N_1924);
or U9416 (N_9416,N_3412,N_656);
nand U9417 (N_9417,N_625,N_1416);
or U9418 (N_9418,N_4025,N_1740);
nand U9419 (N_9419,N_4449,N_3590);
nand U9420 (N_9420,N_4677,N_3410);
nor U9421 (N_9421,N_1228,N_2070);
or U9422 (N_9422,N_790,N_2462);
or U9423 (N_9423,N_3252,N_3428);
nand U9424 (N_9424,N_1991,N_1012);
xor U9425 (N_9425,N_1753,N_2392);
xor U9426 (N_9426,N_525,N_2818);
or U9427 (N_9427,N_851,N_3694);
nor U9428 (N_9428,N_836,N_4638);
xor U9429 (N_9429,N_264,N_4519);
and U9430 (N_9430,N_561,N_3926);
xor U9431 (N_9431,N_4014,N_1744);
xnor U9432 (N_9432,N_4989,N_1987);
and U9433 (N_9433,N_3694,N_636);
nand U9434 (N_9434,N_882,N_3910);
and U9435 (N_9435,N_2401,N_2712);
and U9436 (N_9436,N_1967,N_747);
or U9437 (N_9437,N_14,N_1197);
xor U9438 (N_9438,N_527,N_3636);
xnor U9439 (N_9439,N_4390,N_4061);
and U9440 (N_9440,N_1519,N_2934);
and U9441 (N_9441,N_2165,N_1076);
nand U9442 (N_9442,N_340,N_1151);
and U9443 (N_9443,N_4170,N_1593);
or U9444 (N_9444,N_1695,N_3462);
and U9445 (N_9445,N_420,N_4933);
and U9446 (N_9446,N_3863,N_2787);
nand U9447 (N_9447,N_1388,N_2899);
nor U9448 (N_9448,N_3184,N_3600);
or U9449 (N_9449,N_2608,N_1479);
or U9450 (N_9450,N_1269,N_3628);
and U9451 (N_9451,N_2268,N_4089);
nand U9452 (N_9452,N_2724,N_4989);
and U9453 (N_9453,N_145,N_4147);
nand U9454 (N_9454,N_4447,N_1924);
or U9455 (N_9455,N_4183,N_11);
or U9456 (N_9456,N_4171,N_3098);
xor U9457 (N_9457,N_4688,N_4020);
nor U9458 (N_9458,N_2277,N_4680);
nor U9459 (N_9459,N_1057,N_1675);
or U9460 (N_9460,N_1847,N_4061);
xor U9461 (N_9461,N_4775,N_946);
and U9462 (N_9462,N_662,N_4974);
or U9463 (N_9463,N_4654,N_4985);
and U9464 (N_9464,N_2933,N_3041);
or U9465 (N_9465,N_170,N_1045);
xnor U9466 (N_9466,N_640,N_940);
nor U9467 (N_9467,N_2858,N_3057);
xor U9468 (N_9468,N_2088,N_2353);
nor U9469 (N_9469,N_4617,N_4515);
xor U9470 (N_9470,N_2800,N_2054);
and U9471 (N_9471,N_2380,N_4356);
or U9472 (N_9472,N_4066,N_3326);
and U9473 (N_9473,N_2234,N_706);
or U9474 (N_9474,N_3291,N_2140);
or U9475 (N_9475,N_1297,N_3601);
nor U9476 (N_9476,N_2968,N_2686);
xor U9477 (N_9477,N_1523,N_2873);
and U9478 (N_9478,N_390,N_1886);
or U9479 (N_9479,N_4568,N_749);
and U9480 (N_9480,N_1299,N_2011);
xor U9481 (N_9481,N_3638,N_1941);
nor U9482 (N_9482,N_2025,N_3550);
and U9483 (N_9483,N_4030,N_1545);
nor U9484 (N_9484,N_3632,N_1380);
xnor U9485 (N_9485,N_1755,N_467);
nand U9486 (N_9486,N_1271,N_799);
nand U9487 (N_9487,N_4945,N_3887);
nor U9488 (N_9488,N_1487,N_2137);
or U9489 (N_9489,N_4336,N_3251);
and U9490 (N_9490,N_3965,N_1567);
xor U9491 (N_9491,N_2282,N_774);
nor U9492 (N_9492,N_2695,N_43);
nand U9493 (N_9493,N_626,N_4659);
nand U9494 (N_9494,N_1634,N_2122);
nand U9495 (N_9495,N_3248,N_4070);
nand U9496 (N_9496,N_744,N_1418);
and U9497 (N_9497,N_956,N_1689);
nor U9498 (N_9498,N_725,N_3239);
nand U9499 (N_9499,N_2969,N_2464);
nand U9500 (N_9500,N_700,N_4020);
and U9501 (N_9501,N_1688,N_1511);
or U9502 (N_9502,N_4113,N_70);
or U9503 (N_9503,N_2725,N_4638);
and U9504 (N_9504,N_2556,N_767);
and U9505 (N_9505,N_2895,N_1558);
nor U9506 (N_9506,N_3068,N_3665);
and U9507 (N_9507,N_2110,N_1869);
or U9508 (N_9508,N_43,N_3727);
nand U9509 (N_9509,N_3929,N_2536);
or U9510 (N_9510,N_2607,N_1984);
nor U9511 (N_9511,N_1410,N_3936);
and U9512 (N_9512,N_3380,N_4921);
xor U9513 (N_9513,N_3753,N_3113);
or U9514 (N_9514,N_1032,N_4173);
and U9515 (N_9515,N_2958,N_580);
xnor U9516 (N_9516,N_1319,N_2478);
and U9517 (N_9517,N_172,N_4660);
nand U9518 (N_9518,N_1144,N_2933);
xnor U9519 (N_9519,N_1072,N_3543);
nor U9520 (N_9520,N_1987,N_1162);
nor U9521 (N_9521,N_2556,N_1913);
or U9522 (N_9522,N_4515,N_4759);
nor U9523 (N_9523,N_4727,N_3752);
nand U9524 (N_9524,N_1688,N_2013);
or U9525 (N_9525,N_3515,N_2680);
nor U9526 (N_9526,N_2147,N_4995);
xnor U9527 (N_9527,N_1896,N_4407);
nor U9528 (N_9528,N_844,N_3505);
nand U9529 (N_9529,N_2171,N_4128);
and U9530 (N_9530,N_4654,N_4409);
and U9531 (N_9531,N_2452,N_2939);
nand U9532 (N_9532,N_159,N_101);
and U9533 (N_9533,N_1692,N_2912);
nand U9534 (N_9534,N_946,N_3137);
nand U9535 (N_9535,N_1118,N_3202);
xnor U9536 (N_9536,N_1147,N_3683);
nor U9537 (N_9537,N_3029,N_511);
xor U9538 (N_9538,N_3613,N_532);
and U9539 (N_9539,N_949,N_2947);
and U9540 (N_9540,N_538,N_1167);
nand U9541 (N_9541,N_4516,N_3147);
nand U9542 (N_9542,N_2368,N_4589);
and U9543 (N_9543,N_3631,N_1640);
and U9544 (N_9544,N_3035,N_4254);
or U9545 (N_9545,N_3775,N_3036);
or U9546 (N_9546,N_3469,N_4836);
xor U9547 (N_9547,N_1245,N_788);
nand U9548 (N_9548,N_4143,N_3298);
nand U9549 (N_9549,N_2219,N_1059);
nand U9550 (N_9550,N_2428,N_218);
and U9551 (N_9551,N_4933,N_1801);
xor U9552 (N_9552,N_1229,N_2877);
xor U9553 (N_9553,N_1166,N_820);
xnor U9554 (N_9554,N_2272,N_2637);
or U9555 (N_9555,N_1059,N_599);
nor U9556 (N_9556,N_1202,N_2292);
nand U9557 (N_9557,N_457,N_1873);
nand U9558 (N_9558,N_1843,N_771);
nand U9559 (N_9559,N_3331,N_4827);
and U9560 (N_9560,N_1962,N_2633);
or U9561 (N_9561,N_4043,N_650);
xor U9562 (N_9562,N_2949,N_3020);
or U9563 (N_9563,N_2103,N_3482);
nand U9564 (N_9564,N_2697,N_3539);
or U9565 (N_9565,N_4704,N_4530);
nand U9566 (N_9566,N_600,N_74);
nand U9567 (N_9567,N_447,N_2340);
nor U9568 (N_9568,N_2525,N_3091);
and U9569 (N_9569,N_952,N_4981);
nor U9570 (N_9570,N_1507,N_4442);
and U9571 (N_9571,N_39,N_4269);
nor U9572 (N_9572,N_954,N_1636);
nand U9573 (N_9573,N_2166,N_2425);
or U9574 (N_9574,N_1908,N_540);
and U9575 (N_9575,N_3086,N_749);
and U9576 (N_9576,N_448,N_4295);
xnor U9577 (N_9577,N_1733,N_4836);
and U9578 (N_9578,N_4723,N_1511);
xor U9579 (N_9579,N_675,N_3203);
xnor U9580 (N_9580,N_4328,N_3699);
nand U9581 (N_9581,N_3835,N_587);
and U9582 (N_9582,N_3405,N_3831);
xor U9583 (N_9583,N_4923,N_4117);
and U9584 (N_9584,N_2766,N_368);
nand U9585 (N_9585,N_2717,N_4385);
nand U9586 (N_9586,N_4557,N_2664);
xor U9587 (N_9587,N_761,N_478);
or U9588 (N_9588,N_4448,N_1543);
nor U9589 (N_9589,N_3176,N_1157);
nand U9590 (N_9590,N_722,N_2076);
nor U9591 (N_9591,N_3991,N_7);
nand U9592 (N_9592,N_4795,N_4674);
xnor U9593 (N_9593,N_4471,N_4279);
and U9594 (N_9594,N_1228,N_4161);
xor U9595 (N_9595,N_4686,N_1625);
nor U9596 (N_9596,N_2976,N_737);
or U9597 (N_9597,N_1181,N_2987);
nor U9598 (N_9598,N_3979,N_3840);
or U9599 (N_9599,N_893,N_3349);
or U9600 (N_9600,N_3938,N_1429);
and U9601 (N_9601,N_1307,N_2167);
xor U9602 (N_9602,N_103,N_2830);
and U9603 (N_9603,N_3898,N_4232);
nor U9604 (N_9604,N_1161,N_4437);
nand U9605 (N_9605,N_2510,N_1766);
nand U9606 (N_9606,N_3190,N_273);
nor U9607 (N_9607,N_1206,N_4150);
nor U9608 (N_9608,N_4447,N_2765);
and U9609 (N_9609,N_3601,N_2363);
nand U9610 (N_9610,N_145,N_4624);
or U9611 (N_9611,N_3952,N_4566);
nor U9612 (N_9612,N_4856,N_2128);
or U9613 (N_9613,N_4725,N_107);
xnor U9614 (N_9614,N_58,N_55);
or U9615 (N_9615,N_639,N_1508);
and U9616 (N_9616,N_227,N_1883);
xnor U9617 (N_9617,N_452,N_290);
xnor U9618 (N_9618,N_2314,N_1693);
and U9619 (N_9619,N_76,N_2399);
or U9620 (N_9620,N_1223,N_4527);
nor U9621 (N_9621,N_2870,N_4644);
or U9622 (N_9622,N_380,N_3077);
or U9623 (N_9623,N_2839,N_563);
or U9624 (N_9624,N_816,N_1218);
nand U9625 (N_9625,N_4447,N_37);
and U9626 (N_9626,N_4226,N_4779);
xor U9627 (N_9627,N_651,N_3257);
or U9628 (N_9628,N_4005,N_3814);
nand U9629 (N_9629,N_3270,N_3999);
nand U9630 (N_9630,N_2424,N_3882);
xor U9631 (N_9631,N_3255,N_4282);
xnor U9632 (N_9632,N_257,N_717);
xnor U9633 (N_9633,N_1022,N_1163);
or U9634 (N_9634,N_1243,N_1900);
or U9635 (N_9635,N_4666,N_564);
nand U9636 (N_9636,N_3911,N_3334);
and U9637 (N_9637,N_3742,N_4041);
and U9638 (N_9638,N_2600,N_3110);
nand U9639 (N_9639,N_2340,N_2529);
nand U9640 (N_9640,N_3906,N_2415);
nor U9641 (N_9641,N_667,N_971);
or U9642 (N_9642,N_4887,N_4744);
xnor U9643 (N_9643,N_4663,N_387);
xor U9644 (N_9644,N_1061,N_2270);
or U9645 (N_9645,N_3187,N_571);
or U9646 (N_9646,N_2294,N_319);
nor U9647 (N_9647,N_4018,N_2933);
nor U9648 (N_9648,N_2133,N_517);
nand U9649 (N_9649,N_1429,N_2842);
nor U9650 (N_9650,N_1370,N_4226);
xnor U9651 (N_9651,N_806,N_256);
nand U9652 (N_9652,N_933,N_3568);
or U9653 (N_9653,N_2865,N_831);
and U9654 (N_9654,N_3803,N_1527);
or U9655 (N_9655,N_3466,N_1906);
xor U9656 (N_9656,N_474,N_481);
or U9657 (N_9657,N_2256,N_1258);
nor U9658 (N_9658,N_4338,N_3693);
nor U9659 (N_9659,N_594,N_767);
and U9660 (N_9660,N_1054,N_4542);
nor U9661 (N_9661,N_3628,N_3311);
and U9662 (N_9662,N_4900,N_4122);
or U9663 (N_9663,N_1003,N_4590);
xnor U9664 (N_9664,N_826,N_3118);
or U9665 (N_9665,N_1885,N_2033);
or U9666 (N_9666,N_3543,N_2547);
nand U9667 (N_9667,N_691,N_939);
and U9668 (N_9668,N_828,N_3264);
nor U9669 (N_9669,N_2573,N_3621);
and U9670 (N_9670,N_912,N_4836);
or U9671 (N_9671,N_1521,N_1995);
xor U9672 (N_9672,N_2891,N_4929);
xnor U9673 (N_9673,N_2799,N_2907);
or U9674 (N_9674,N_1515,N_3722);
or U9675 (N_9675,N_2801,N_3162);
xnor U9676 (N_9676,N_1788,N_1918);
nand U9677 (N_9677,N_1333,N_4151);
nor U9678 (N_9678,N_3630,N_4001);
and U9679 (N_9679,N_3949,N_2703);
nor U9680 (N_9680,N_4220,N_4942);
nor U9681 (N_9681,N_3490,N_1895);
nor U9682 (N_9682,N_3778,N_179);
nand U9683 (N_9683,N_1074,N_4004);
and U9684 (N_9684,N_562,N_2329);
nor U9685 (N_9685,N_1658,N_3623);
and U9686 (N_9686,N_859,N_2444);
nor U9687 (N_9687,N_1361,N_695);
xor U9688 (N_9688,N_3893,N_4383);
or U9689 (N_9689,N_499,N_2689);
nor U9690 (N_9690,N_989,N_1737);
or U9691 (N_9691,N_2755,N_1019);
nor U9692 (N_9692,N_2214,N_4361);
or U9693 (N_9693,N_2614,N_3408);
nor U9694 (N_9694,N_271,N_2668);
and U9695 (N_9695,N_474,N_2649);
nand U9696 (N_9696,N_2233,N_4272);
and U9697 (N_9697,N_4922,N_1186);
nor U9698 (N_9698,N_1969,N_911);
xnor U9699 (N_9699,N_294,N_1966);
nor U9700 (N_9700,N_1058,N_580);
or U9701 (N_9701,N_383,N_318);
and U9702 (N_9702,N_4402,N_2962);
nand U9703 (N_9703,N_2550,N_1349);
nor U9704 (N_9704,N_2476,N_2771);
or U9705 (N_9705,N_50,N_4585);
and U9706 (N_9706,N_3727,N_2740);
xnor U9707 (N_9707,N_3120,N_4891);
xnor U9708 (N_9708,N_143,N_1410);
nand U9709 (N_9709,N_2862,N_3924);
nor U9710 (N_9710,N_1612,N_1517);
nor U9711 (N_9711,N_2425,N_4355);
or U9712 (N_9712,N_1333,N_4421);
or U9713 (N_9713,N_4946,N_2900);
or U9714 (N_9714,N_205,N_2250);
xor U9715 (N_9715,N_3337,N_3431);
nand U9716 (N_9716,N_45,N_718);
nor U9717 (N_9717,N_2640,N_3757);
nor U9718 (N_9718,N_228,N_4185);
xnor U9719 (N_9719,N_3368,N_1012);
nor U9720 (N_9720,N_2244,N_2211);
and U9721 (N_9721,N_4185,N_795);
nand U9722 (N_9722,N_3593,N_2397);
or U9723 (N_9723,N_2685,N_4145);
nor U9724 (N_9724,N_2965,N_2680);
or U9725 (N_9725,N_4979,N_1421);
or U9726 (N_9726,N_1748,N_2696);
nor U9727 (N_9727,N_373,N_2295);
and U9728 (N_9728,N_2168,N_2282);
xor U9729 (N_9729,N_1884,N_3368);
or U9730 (N_9730,N_3230,N_1312);
nor U9731 (N_9731,N_1976,N_104);
nor U9732 (N_9732,N_3608,N_77);
and U9733 (N_9733,N_4100,N_834);
xor U9734 (N_9734,N_2388,N_3988);
or U9735 (N_9735,N_1648,N_1702);
xor U9736 (N_9736,N_211,N_1830);
xnor U9737 (N_9737,N_1764,N_101);
nand U9738 (N_9738,N_1459,N_3678);
nand U9739 (N_9739,N_1389,N_28);
or U9740 (N_9740,N_686,N_3462);
nor U9741 (N_9741,N_689,N_2208);
and U9742 (N_9742,N_3496,N_3285);
nand U9743 (N_9743,N_3959,N_1219);
nand U9744 (N_9744,N_3757,N_1227);
nand U9745 (N_9745,N_4723,N_2634);
nand U9746 (N_9746,N_1979,N_2114);
nor U9747 (N_9747,N_2018,N_4626);
and U9748 (N_9748,N_2646,N_179);
nand U9749 (N_9749,N_1193,N_2719);
nor U9750 (N_9750,N_2686,N_4501);
nor U9751 (N_9751,N_375,N_2743);
nor U9752 (N_9752,N_3748,N_3214);
or U9753 (N_9753,N_4428,N_3149);
and U9754 (N_9754,N_3421,N_3070);
or U9755 (N_9755,N_3937,N_2292);
and U9756 (N_9756,N_1264,N_3175);
xnor U9757 (N_9757,N_2526,N_158);
xnor U9758 (N_9758,N_4953,N_3378);
nand U9759 (N_9759,N_4681,N_3074);
or U9760 (N_9760,N_472,N_4223);
nand U9761 (N_9761,N_1417,N_3652);
nor U9762 (N_9762,N_2576,N_3779);
and U9763 (N_9763,N_1121,N_719);
nor U9764 (N_9764,N_1753,N_4549);
nor U9765 (N_9765,N_334,N_522);
xnor U9766 (N_9766,N_4947,N_1309);
or U9767 (N_9767,N_4296,N_2042);
and U9768 (N_9768,N_2101,N_2820);
xnor U9769 (N_9769,N_4754,N_3664);
nor U9770 (N_9770,N_2383,N_3981);
or U9771 (N_9771,N_4772,N_3854);
xor U9772 (N_9772,N_775,N_3980);
nand U9773 (N_9773,N_22,N_2819);
or U9774 (N_9774,N_535,N_2983);
nand U9775 (N_9775,N_1465,N_4538);
nor U9776 (N_9776,N_902,N_3219);
xor U9777 (N_9777,N_1252,N_160);
and U9778 (N_9778,N_2821,N_4561);
nor U9779 (N_9779,N_3638,N_4433);
nand U9780 (N_9780,N_4106,N_2431);
or U9781 (N_9781,N_1060,N_4025);
nand U9782 (N_9782,N_2300,N_4197);
or U9783 (N_9783,N_2851,N_343);
xor U9784 (N_9784,N_4099,N_2889);
and U9785 (N_9785,N_1993,N_4345);
nor U9786 (N_9786,N_2384,N_3210);
nand U9787 (N_9787,N_3349,N_2932);
or U9788 (N_9788,N_2116,N_405);
or U9789 (N_9789,N_2866,N_156);
xnor U9790 (N_9790,N_644,N_4197);
and U9791 (N_9791,N_3409,N_3285);
nor U9792 (N_9792,N_4075,N_4575);
and U9793 (N_9793,N_462,N_2847);
nand U9794 (N_9794,N_1691,N_1737);
nand U9795 (N_9795,N_1242,N_2794);
nand U9796 (N_9796,N_2180,N_739);
nor U9797 (N_9797,N_2556,N_4020);
xor U9798 (N_9798,N_1970,N_3646);
nand U9799 (N_9799,N_2088,N_662);
and U9800 (N_9800,N_3828,N_2060);
nand U9801 (N_9801,N_1137,N_3732);
nand U9802 (N_9802,N_1714,N_3980);
nand U9803 (N_9803,N_4287,N_2061);
or U9804 (N_9804,N_1943,N_268);
nand U9805 (N_9805,N_2035,N_1243);
nand U9806 (N_9806,N_390,N_3617);
nand U9807 (N_9807,N_2840,N_2625);
xnor U9808 (N_9808,N_4100,N_2972);
or U9809 (N_9809,N_3076,N_4098);
and U9810 (N_9810,N_2176,N_4576);
xnor U9811 (N_9811,N_4309,N_3813);
nand U9812 (N_9812,N_3063,N_2210);
and U9813 (N_9813,N_4446,N_818);
xor U9814 (N_9814,N_174,N_1619);
nand U9815 (N_9815,N_439,N_1823);
nand U9816 (N_9816,N_4910,N_138);
or U9817 (N_9817,N_1265,N_2477);
nor U9818 (N_9818,N_4634,N_1695);
nand U9819 (N_9819,N_4499,N_1562);
xnor U9820 (N_9820,N_465,N_810);
xor U9821 (N_9821,N_2238,N_3773);
and U9822 (N_9822,N_1571,N_3580);
nor U9823 (N_9823,N_4315,N_1642);
nor U9824 (N_9824,N_4149,N_509);
xnor U9825 (N_9825,N_3210,N_1680);
nand U9826 (N_9826,N_4512,N_2686);
and U9827 (N_9827,N_3958,N_2710);
xor U9828 (N_9828,N_3851,N_4089);
xor U9829 (N_9829,N_1846,N_4167);
or U9830 (N_9830,N_514,N_1006);
nand U9831 (N_9831,N_4564,N_3898);
or U9832 (N_9832,N_3896,N_4405);
xor U9833 (N_9833,N_4579,N_2652);
xor U9834 (N_9834,N_764,N_3638);
nand U9835 (N_9835,N_192,N_1093);
and U9836 (N_9836,N_1749,N_1811);
xnor U9837 (N_9837,N_2721,N_1486);
and U9838 (N_9838,N_3248,N_2228);
xor U9839 (N_9839,N_3189,N_3526);
and U9840 (N_9840,N_325,N_2144);
or U9841 (N_9841,N_2372,N_3952);
nor U9842 (N_9842,N_2384,N_4911);
nand U9843 (N_9843,N_2660,N_2840);
nand U9844 (N_9844,N_2330,N_4208);
xor U9845 (N_9845,N_3101,N_2275);
and U9846 (N_9846,N_1390,N_4514);
nor U9847 (N_9847,N_3456,N_234);
and U9848 (N_9848,N_1989,N_3533);
nor U9849 (N_9849,N_1081,N_1787);
xnor U9850 (N_9850,N_1200,N_4263);
xnor U9851 (N_9851,N_3369,N_1653);
nor U9852 (N_9852,N_2722,N_1767);
xnor U9853 (N_9853,N_4516,N_3921);
nor U9854 (N_9854,N_4585,N_1388);
nor U9855 (N_9855,N_4567,N_4653);
xor U9856 (N_9856,N_213,N_420);
and U9857 (N_9857,N_2726,N_4209);
and U9858 (N_9858,N_308,N_4776);
nor U9859 (N_9859,N_3199,N_1657);
and U9860 (N_9860,N_1507,N_1605);
nor U9861 (N_9861,N_4402,N_4392);
xor U9862 (N_9862,N_18,N_1391);
nand U9863 (N_9863,N_2776,N_1256);
nand U9864 (N_9864,N_1726,N_1244);
nand U9865 (N_9865,N_1511,N_4350);
nand U9866 (N_9866,N_1543,N_3652);
nor U9867 (N_9867,N_4103,N_3511);
and U9868 (N_9868,N_532,N_1452);
nand U9869 (N_9869,N_4259,N_4694);
and U9870 (N_9870,N_4565,N_3090);
nand U9871 (N_9871,N_735,N_2732);
and U9872 (N_9872,N_4444,N_3107);
and U9873 (N_9873,N_3912,N_3774);
xor U9874 (N_9874,N_4344,N_581);
nand U9875 (N_9875,N_855,N_2102);
nor U9876 (N_9876,N_411,N_2443);
or U9877 (N_9877,N_524,N_4559);
or U9878 (N_9878,N_328,N_2708);
and U9879 (N_9879,N_4639,N_3873);
and U9880 (N_9880,N_3648,N_3891);
and U9881 (N_9881,N_479,N_301);
xor U9882 (N_9882,N_220,N_3540);
nand U9883 (N_9883,N_2755,N_3355);
nor U9884 (N_9884,N_304,N_1909);
nand U9885 (N_9885,N_4376,N_2615);
nand U9886 (N_9886,N_2540,N_4029);
and U9887 (N_9887,N_2391,N_143);
nor U9888 (N_9888,N_1696,N_3936);
nand U9889 (N_9889,N_4798,N_4326);
or U9890 (N_9890,N_2461,N_2274);
nand U9891 (N_9891,N_3444,N_2164);
nor U9892 (N_9892,N_367,N_1121);
xnor U9893 (N_9893,N_1930,N_2732);
nand U9894 (N_9894,N_2607,N_1388);
or U9895 (N_9895,N_2164,N_1420);
nand U9896 (N_9896,N_4131,N_2993);
or U9897 (N_9897,N_1709,N_2141);
or U9898 (N_9898,N_1408,N_3567);
or U9899 (N_9899,N_4194,N_4353);
xnor U9900 (N_9900,N_139,N_3221);
nand U9901 (N_9901,N_2383,N_4995);
and U9902 (N_9902,N_4300,N_1616);
and U9903 (N_9903,N_4351,N_4232);
or U9904 (N_9904,N_2528,N_1100);
nand U9905 (N_9905,N_4853,N_1797);
and U9906 (N_9906,N_3086,N_4142);
xnor U9907 (N_9907,N_4117,N_3895);
and U9908 (N_9908,N_3497,N_1833);
or U9909 (N_9909,N_2181,N_3021);
or U9910 (N_9910,N_2175,N_3793);
xnor U9911 (N_9911,N_654,N_3484);
xnor U9912 (N_9912,N_4429,N_1483);
nand U9913 (N_9913,N_2395,N_1842);
nand U9914 (N_9914,N_215,N_2104);
nor U9915 (N_9915,N_251,N_3258);
nor U9916 (N_9916,N_4459,N_1069);
xnor U9917 (N_9917,N_1446,N_3744);
nand U9918 (N_9918,N_2775,N_2434);
and U9919 (N_9919,N_2461,N_2502);
or U9920 (N_9920,N_2918,N_1766);
or U9921 (N_9921,N_3391,N_4504);
xor U9922 (N_9922,N_3814,N_1655);
nor U9923 (N_9923,N_3505,N_3045);
xnor U9924 (N_9924,N_776,N_1418);
nor U9925 (N_9925,N_825,N_259);
xnor U9926 (N_9926,N_532,N_2070);
and U9927 (N_9927,N_4992,N_1868);
and U9928 (N_9928,N_2358,N_673);
nor U9929 (N_9929,N_3705,N_1326);
nor U9930 (N_9930,N_1131,N_1757);
and U9931 (N_9931,N_2358,N_3440);
xnor U9932 (N_9932,N_1482,N_1892);
and U9933 (N_9933,N_3533,N_1237);
or U9934 (N_9934,N_2874,N_1275);
nand U9935 (N_9935,N_4809,N_1220);
or U9936 (N_9936,N_3948,N_4166);
nand U9937 (N_9937,N_3761,N_331);
or U9938 (N_9938,N_4471,N_237);
nor U9939 (N_9939,N_1924,N_1353);
xnor U9940 (N_9940,N_2602,N_94);
nand U9941 (N_9941,N_2373,N_4399);
xor U9942 (N_9942,N_1815,N_2702);
nor U9943 (N_9943,N_3467,N_440);
or U9944 (N_9944,N_3980,N_222);
or U9945 (N_9945,N_2227,N_3574);
and U9946 (N_9946,N_680,N_2771);
xor U9947 (N_9947,N_564,N_3107);
xnor U9948 (N_9948,N_1253,N_156);
and U9949 (N_9949,N_1948,N_296);
xnor U9950 (N_9950,N_433,N_2003);
and U9951 (N_9951,N_3503,N_4449);
nand U9952 (N_9952,N_570,N_1051);
or U9953 (N_9953,N_4854,N_537);
nor U9954 (N_9954,N_1826,N_523);
nand U9955 (N_9955,N_4500,N_1135);
and U9956 (N_9956,N_2043,N_4228);
xnor U9957 (N_9957,N_3221,N_2522);
nand U9958 (N_9958,N_2936,N_3648);
xor U9959 (N_9959,N_4787,N_33);
xor U9960 (N_9960,N_2451,N_4301);
nand U9961 (N_9961,N_1286,N_773);
xnor U9962 (N_9962,N_4702,N_442);
or U9963 (N_9963,N_4447,N_2078);
nor U9964 (N_9964,N_3542,N_4893);
nand U9965 (N_9965,N_1157,N_1638);
xor U9966 (N_9966,N_1661,N_3313);
xor U9967 (N_9967,N_2946,N_3113);
nor U9968 (N_9968,N_4536,N_855);
and U9969 (N_9969,N_3752,N_400);
nor U9970 (N_9970,N_1479,N_1169);
and U9971 (N_9971,N_4852,N_2052);
nor U9972 (N_9972,N_11,N_3039);
xnor U9973 (N_9973,N_1751,N_2057);
and U9974 (N_9974,N_4982,N_1116);
nand U9975 (N_9975,N_1707,N_2866);
nand U9976 (N_9976,N_1218,N_3402);
and U9977 (N_9977,N_1769,N_4540);
nor U9978 (N_9978,N_2912,N_1653);
xnor U9979 (N_9979,N_2317,N_180);
nand U9980 (N_9980,N_2186,N_1469);
nand U9981 (N_9981,N_862,N_1282);
or U9982 (N_9982,N_4713,N_3649);
nor U9983 (N_9983,N_4357,N_4110);
xor U9984 (N_9984,N_4035,N_4326);
xor U9985 (N_9985,N_360,N_1887);
or U9986 (N_9986,N_4260,N_747);
or U9987 (N_9987,N_2999,N_3949);
or U9988 (N_9988,N_1816,N_1418);
and U9989 (N_9989,N_909,N_2925);
nand U9990 (N_9990,N_4247,N_738);
nand U9991 (N_9991,N_867,N_2852);
and U9992 (N_9992,N_1342,N_3722);
or U9993 (N_9993,N_3117,N_1729);
xor U9994 (N_9994,N_3950,N_2697);
xor U9995 (N_9995,N_8,N_2346);
nand U9996 (N_9996,N_2275,N_2025);
xnor U9997 (N_9997,N_654,N_3631);
xor U9998 (N_9998,N_4343,N_3758);
nor U9999 (N_9999,N_4199,N_2117);
xor U10000 (N_10000,N_8431,N_5729);
or U10001 (N_10001,N_7270,N_8364);
xnor U10002 (N_10002,N_8980,N_6560);
or U10003 (N_10003,N_5131,N_7751);
xnor U10004 (N_10004,N_9505,N_9070);
nand U10005 (N_10005,N_7106,N_5981);
and U10006 (N_10006,N_6417,N_9180);
xnor U10007 (N_10007,N_8586,N_6369);
xnor U10008 (N_10008,N_6587,N_9645);
nor U10009 (N_10009,N_6672,N_5835);
nor U10010 (N_10010,N_8571,N_7323);
xnor U10011 (N_10011,N_6289,N_9034);
or U10012 (N_10012,N_8896,N_7836);
and U10013 (N_10013,N_6564,N_7001);
xor U10014 (N_10014,N_8573,N_6820);
xnor U10015 (N_10015,N_9851,N_9488);
xnor U10016 (N_10016,N_8520,N_9668);
nor U10017 (N_10017,N_8578,N_6738);
or U10018 (N_10018,N_9606,N_9967);
or U10019 (N_10019,N_7380,N_9802);
nor U10020 (N_10020,N_7673,N_8822);
or U10021 (N_10021,N_8927,N_7044);
nor U10022 (N_10022,N_6461,N_6965);
or U10023 (N_10023,N_9050,N_8397);
or U10024 (N_10024,N_8873,N_7926);
nor U10025 (N_10025,N_7703,N_9401);
and U10026 (N_10026,N_7211,N_7951);
nor U10027 (N_10027,N_7724,N_7586);
nor U10028 (N_10028,N_6394,N_8061);
and U10029 (N_10029,N_8239,N_5434);
or U10030 (N_10030,N_8048,N_7506);
or U10031 (N_10031,N_9843,N_7755);
nand U10032 (N_10032,N_9278,N_7818);
nor U10033 (N_10033,N_7614,N_7918);
and U10034 (N_10034,N_6575,N_5908);
and U10035 (N_10035,N_5818,N_7432);
nand U10036 (N_10036,N_6987,N_9350);
and U10037 (N_10037,N_7788,N_5970);
xnor U10038 (N_10038,N_7035,N_6411);
or U10039 (N_10039,N_6204,N_5998);
xnor U10040 (N_10040,N_8248,N_6261);
or U10041 (N_10041,N_7539,N_8490);
nor U10042 (N_10042,N_9248,N_5789);
or U10043 (N_10043,N_8416,N_5150);
xnor U10044 (N_10044,N_7004,N_7983);
xor U10045 (N_10045,N_7789,N_7347);
nand U10046 (N_10046,N_9281,N_9461);
nor U10047 (N_10047,N_9101,N_8512);
and U10048 (N_10048,N_9184,N_9059);
nand U10049 (N_10049,N_5192,N_5666);
nand U10050 (N_10050,N_6771,N_9354);
nor U10051 (N_10051,N_7538,N_8700);
and U10052 (N_10052,N_5643,N_7273);
nor U10053 (N_10053,N_7125,N_8173);
and U10054 (N_10054,N_9166,N_9508);
or U10055 (N_10055,N_8461,N_5313);
xnor U10056 (N_10056,N_5253,N_6128);
and U10057 (N_10057,N_9377,N_5285);
xor U10058 (N_10058,N_8645,N_9476);
nand U10059 (N_10059,N_7906,N_5028);
and U10060 (N_10060,N_7337,N_8916);
nor U10061 (N_10061,N_7490,N_5623);
nand U10062 (N_10062,N_8511,N_6397);
xnor U10063 (N_10063,N_6806,N_7435);
or U10064 (N_10064,N_7866,N_9307);
nand U10065 (N_10065,N_9181,N_8079);
nor U10066 (N_10066,N_5006,N_8045);
or U10067 (N_10067,N_7180,N_7953);
nand U10068 (N_10068,N_9300,N_7403);
and U10069 (N_10069,N_5871,N_6915);
and U10070 (N_10070,N_8480,N_5370);
xnor U10071 (N_10071,N_6252,N_5939);
nand U10072 (N_10072,N_9466,N_8517);
or U10073 (N_10073,N_5201,N_7842);
nor U10074 (N_10074,N_9097,N_5771);
nor U10075 (N_10075,N_5026,N_7075);
xor U10076 (N_10076,N_9019,N_6963);
nor U10077 (N_10077,N_8941,N_7037);
and U10078 (N_10078,N_9257,N_8828);
and U10079 (N_10079,N_8699,N_6632);
or U10080 (N_10080,N_7734,N_5436);
or U10081 (N_10081,N_5164,N_9573);
and U10082 (N_10082,N_6920,N_9064);
or U10083 (N_10083,N_7716,N_8414);
nor U10084 (N_10084,N_6666,N_9363);
nor U10085 (N_10085,N_5921,N_5162);
nand U10086 (N_10086,N_9785,N_6079);
and U10087 (N_10087,N_9614,N_5013);
and U10088 (N_10088,N_9976,N_9302);
and U10089 (N_10089,N_8965,N_8006);
xnor U10090 (N_10090,N_8555,N_5504);
or U10091 (N_10091,N_9385,N_6420);
and U10092 (N_10092,N_9663,N_7174);
xor U10093 (N_10093,N_6177,N_7553);
and U10094 (N_10094,N_5378,N_8116);
nand U10095 (N_10095,N_7782,N_5545);
xnor U10096 (N_10096,N_5958,N_8832);
xnor U10097 (N_10097,N_6059,N_6961);
nand U10098 (N_10098,N_9225,N_9456);
nand U10099 (N_10099,N_5293,N_5803);
or U10100 (N_10100,N_5445,N_8479);
or U10101 (N_10101,N_7613,N_8703);
nor U10102 (N_10102,N_7177,N_9211);
nand U10103 (N_10103,N_8805,N_6409);
or U10104 (N_10104,N_9028,N_5922);
nand U10105 (N_10105,N_8887,N_8535);
nor U10106 (N_10106,N_8212,N_5777);
xnor U10107 (N_10107,N_5810,N_6708);
nor U10108 (N_10108,N_8936,N_6041);
nor U10109 (N_10109,N_9590,N_7007);
or U10110 (N_10110,N_8684,N_8647);
xor U10111 (N_10111,N_8168,N_6939);
nor U10112 (N_10112,N_5284,N_8170);
nor U10113 (N_10113,N_5189,N_8504);
nor U10114 (N_10114,N_7253,N_9289);
xor U10115 (N_10115,N_5309,N_8085);
or U10116 (N_10116,N_7960,N_8752);
nand U10117 (N_10117,N_9351,N_5538);
nand U10118 (N_10118,N_7028,N_8346);
nand U10119 (N_10119,N_9039,N_7409);
or U10120 (N_10120,N_7984,N_6233);
and U10121 (N_10121,N_6670,N_7431);
nor U10122 (N_10122,N_9051,N_5694);
nor U10123 (N_10123,N_8676,N_7678);
and U10124 (N_10124,N_9173,N_6626);
and U10125 (N_10125,N_9741,N_8419);
nand U10126 (N_10126,N_5595,N_9693);
or U10127 (N_10127,N_5719,N_9942);
and U10128 (N_10128,N_7038,N_7537);
nand U10129 (N_10129,N_7971,N_7512);
nor U10130 (N_10130,N_7945,N_7376);
xnor U10131 (N_10131,N_6971,N_9006);
or U10132 (N_10132,N_9196,N_6194);
nand U10133 (N_10133,N_9395,N_5271);
nor U10134 (N_10134,N_8682,N_5300);
xnor U10135 (N_10135,N_8797,N_5829);
and U10136 (N_10136,N_7145,N_9356);
nor U10137 (N_10137,N_6362,N_6573);
nand U10138 (N_10138,N_9932,N_7890);
or U10139 (N_10139,N_8333,N_5988);
xnor U10140 (N_10140,N_7563,N_9501);
xor U10141 (N_10141,N_5834,N_8204);
or U10142 (N_10142,N_8279,N_6317);
nor U10143 (N_10143,N_6665,N_6761);
xnor U10144 (N_10144,N_5890,N_9472);
or U10145 (N_10145,N_9332,N_7956);
nor U10146 (N_10146,N_7187,N_6726);
and U10147 (N_10147,N_9644,N_7288);
or U10148 (N_10148,N_5498,N_6984);
or U10149 (N_10149,N_6162,N_7349);
or U10150 (N_10150,N_5550,N_8983);
and U10151 (N_10151,N_5033,N_7662);
and U10152 (N_10152,N_6482,N_5991);
xnor U10153 (N_10153,N_8338,N_7274);
nand U10154 (N_10154,N_6827,N_9067);
nand U10155 (N_10155,N_8677,N_5391);
nand U10156 (N_10156,N_7158,N_6232);
and U10157 (N_10157,N_9022,N_5360);
and U10158 (N_10158,N_7454,N_7902);
and U10159 (N_10159,N_8009,N_5959);
and U10160 (N_10160,N_8412,N_5438);
nor U10161 (N_10161,N_7555,N_9891);
nor U10162 (N_10162,N_6800,N_7025);
or U10163 (N_10163,N_6209,N_8500);
nand U10164 (N_10164,N_5885,N_8293);
nand U10165 (N_10165,N_6346,N_9569);
and U10166 (N_10166,N_6373,N_6911);
or U10167 (N_10167,N_9980,N_5521);
or U10168 (N_10168,N_8518,N_8001);
xnor U10169 (N_10169,N_5449,N_8029);
xor U10170 (N_10170,N_9269,N_9899);
xor U10171 (N_10171,N_9268,N_7880);
or U10172 (N_10172,N_5268,N_6060);
or U10173 (N_10173,N_5488,N_5773);
xor U10174 (N_10174,N_5733,N_6154);
nor U10175 (N_10175,N_6500,N_8104);
nor U10176 (N_10176,N_9429,N_9434);
nor U10177 (N_10177,N_8209,N_8465);
nor U10178 (N_10178,N_8196,N_9483);
or U10179 (N_10179,N_5358,N_8991);
and U10180 (N_10180,N_9430,N_7064);
nand U10181 (N_10181,N_8388,N_8050);
nor U10182 (N_10182,N_8049,N_6088);
nor U10183 (N_10183,N_8025,N_7519);
or U10184 (N_10184,N_6716,N_8532);
xor U10185 (N_10185,N_8275,N_8127);
nor U10186 (N_10186,N_7746,N_7640);
nor U10187 (N_10187,N_7031,N_9123);
and U10188 (N_10188,N_7910,N_5899);
xnor U10189 (N_10189,N_9526,N_5965);
nor U10190 (N_10190,N_7164,N_5081);
nor U10191 (N_10191,N_7333,N_7343);
nand U10192 (N_10192,N_9507,N_6486);
nor U10193 (N_10193,N_6251,N_5527);
or U10194 (N_10194,N_7359,N_9112);
xor U10195 (N_10195,N_6360,N_5173);
or U10196 (N_10196,N_6764,N_7546);
nor U10197 (N_10197,N_7666,N_7205);
or U10198 (N_10198,N_5597,N_7943);
nand U10199 (N_10199,N_8640,N_6923);
nand U10200 (N_10200,N_9951,N_8164);
nand U10201 (N_10201,N_6344,N_9383);
nor U10202 (N_10202,N_9177,N_5073);
nor U10203 (N_10203,N_8451,N_9240);
nand U10204 (N_10204,N_7532,N_8046);
nand U10205 (N_10205,N_8734,N_9771);
nor U10206 (N_10206,N_7072,N_9855);
nor U10207 (N_10207,N_8497,N_9035);
xor U10208 (N_10208,N_5185,N_5451);
xor U10209 (N_10209,N_9599,N_9420);
xnor U10210 (N_10210,N_9737,N_8619);
nor U10211 (N_10211,N_7127,N_9730);
and U10212 (N_10212,N_8224,N_6743);
xnor U10213 (N_10213,N_6563,N_7459);
nor U10214 (N_10214,N_9053,N_7478);
or U10215 (N_10215,N_8719,N_7624);
nor U10216 (N_10216,N_6936,N_7964);
nor U10217 (N_10217,N_8120,N_5049);
nor U10218 (N_10218,N_8235,N_6223);
nand U10219 (N_10219,N_8063,N_8909);
or U10220 (N_10220,N_5134,N_5946);
and U10221 (N_10221,N_8038,N_9953);
and U10222 (N_10222,N_8784,N_7171);
or U10223 (N_10223,N_5487,N_6202);
nor U10224 (N_10224,N_5262,N_9286);
nor U10225 (N_10225,N_8407,N_5663);
nand U10226 (N_10226,N_8770,N_6061);
xor U10227 (N_10227,N_9119,N_8713);
nand U10228 (N_10228,N_8362,N_5016);
nor U10229 (N_10229,N_6945,N_5519);
xnor U10230 (N_10230,N_9054,N_7056);
and U10231 (N_10231,N_8399,N_6065);
nor U10232 (N_10232,N_7086,N_5928);
xnor U10233 (N_10233,N_9000,N_6071);
xor U10234 (N_10234,N_5992,N_6833);
nand U10235 (N_10235,N_6906,N_8839);
or U10236 (N_10236,N_6032,N_8148);
nor U10237 (N_10237,N_6774,N_8004);
xnor U10238 (N_10238,N_7641,N_7388);
xnor U10239 (N_10239,N_7003,N_5259);
xnor U10240 (N_10240,N_5238,N_6912);
or U10241 (N_10241,N_5731,N_8718);
or U10242 (N_10242,N_6504,N_8263);
xor U10243 (N_10243,N_8691,N_9988);
nand U10244 (N_10244,N_7603,N_7781);
and U10245 (N_10245,N_5520,N_9640);
nand U10246 (N_10246,N_6406,N_9099);
and U10247 (N_10247,N_7740,N_5154);
and U10248 (N_10248,N_5227,N_5698);
nor U10249 (N_10249,N_5695,N_9413);
nand U10250 (N_10250,N_8642,N_7429);
or U10251 (N_10251,N_7699,N_9312);
nand U10252 (N_10252,N_7776,N_8501);
xnor U10253 (N_10253,N_5739,N_6122);
or U10254 (N_10254,N_8446,N_5406);
xor U10255 (N_10255,N_6677,N_9744);
or U10256 (N_10256,N_5876,N_7103);
nand U10257 (N_10257,N_9468,N_6271);
or U10258 (N_10258,N_7265,N_5897);
and U10259 (N_10259,N_5514,N_7005);
or U10260 (N_10260,N_6085,N_7188);
or U10261 (N_10261,N_7747,N_7043);
or U10262 (N_10262,N_6803,N_9567);
nand U10263 (N_10263,N_7813,N_8098);
nor U10264 (N_10264,N_6644,N_7973);
nor U10265 (N_10265,N_6157,N_6744);
nand U10266 (N_10266,N_6033,N_6365);
nand U10267 (N_10267,N_5424,N_5891);
xor U10268 (N_10268,N_9441,N_8370);
xnor U10269 (N_10269,N_8486,N_9052);
or U10270 (N_10270,N_7462,N_9755);
nand U10271 (N_10271,N_5592,N_6109);
xnor U10272 (N_10272,N_9778,N_5820);
nor U10273 (N_10273,N_9361,N_7576);
xor U10274 (N_10274,N_7050,N_5264);
and U10275 (N_10275,N_9135,N_5786);
or U10276 (N_10276,N_8312,N_8946);
or U10277 (N_10277,N_5392,N_5674);
nand U10278 (N_10278,N_6453,N_8846);
nor U10279 (N_10279,N_7199,N_5178);
xnor U10280 (N_10280,N_6336,N_9936);
or U10281 (N_10281,N_6405,N_8463);
nor U10282 (N_10282,N_7661,N_9303);
nand U10283 (N_10283,N_8287,N_9360);
and U10284 (N_10284,N_5328,N_7358);
and U10285 (N_10285,N_7936,N_5155);
xor U10286 (N_10286,N_5367,N_6582);
nor U10287 (N_10287,N_8187,N_9410);
or U10288 (N_10288,N_9777,N_9973);
and U10289 (N_10289,N_8914,N_9937);
or U10290 (N_10290,N_7352,N_5767);
nor U10291 (N_10291,N_7848,N_6322);
xor U10292 (N_10292,N_8753,N_5652);
and U10293 (N_10293,N_6341,N_5515);
nor U10294 (N_10294,N_8353,N_8122);
and U10295 (N_10295,N_6952,N_5699);
or U10296 (N_10296,N_6762,N_6144);
and U10297 (N_10297,N_7497,N_8184);
or U10298 (N_10298,N_5644,N_6350);
xor U10299 (N_10299,N_5471,N_7606);
xor U10300 (N_10300,N_5825,N_6320);
and U10301 (N_10301,N_7209,N_6054);
nand U10302 (N_10302,N_8929,N_6922);
xor U10303 (N_10303,N_9224,N_8442);
nand U10304 (N_10304,N_6492,N_8251);
nand U10305 (N_10305,N_7655,N_8039);
or U10306 (N_10306,N_9545,N_5823);
and U10307 (N_10307,N_6509,N_9068);
or U10308 (N_10308,N_9450,N_9477);
and U10309 (N_10309,N_8389,N_9105);
or U10310 (N_10310,N_6046,N_7957);
or U10311 (N_10311,N_5894,N_6520);
or U10312 (N_10312,N_7142,N_8881);
nor U10313 (N_10313,N_6025,N_5127);
nand U10314 (N_10314,N_8956,N_5693);
or U10315 (N_10315,N_6353,N_6794);
or U10316 (N_10316,N_5151,N_6068);
xor U10317 (N_10317,N_6725,N_5034);
or U10318 (N_10318,N_8635,N_8810);
nor U10319 (N_10319,N_5403,N_9427);
nor U10320 (N_10320,N_9345,N_7688);
xnor U10321 (N_10321,N_7420,N_5282);
nor U10322 (N_10322,N_6246,N_8195);
xor U10323 (N_10323,N_7305,N_7146);
nand U10324 (N_10324,N_9909,N_9294);
xor U10325 (N_10325,N_6867,N_8710);
or U10326 (N_10326,N_5179,N_5325);
and U10327 (N_10327,N_7297,N_9672);
xor U10328 (N_10328,N_8175,N_8952);
and U10329 (N_10329,N_6446,N_6524);
or U10330 (N_10330,N_8582,N_6311);
or U10331 (N_10331,N_8308,N_7309);
nor U10332 (N_10332,N_9882,N_5724);
xor U10333 (N_10333,N_7224,N_9699);
nand U10334 (N_10334,N_8189,N_6200);
and U10335 (N_10335,N_8202,N_9977);
or U10336 (N_10336,N_7777,N_9653);
nor U10337 (N_10337,N_5098,N_9848);
nand U10338 (N_10338,N_7503,N_5747);
and U10339 (N_10339,N_7727,N_8339);
nand U10340 (N_10340,N_6823,N_8917);
xor U10341 (N_10341,N_6508,N_8767);
and U10342 (N_10342,N_6408,N_7284);
or U10343 (N_10343,N_8086,N_9830);
nor U10344 (N_10344,N_5923,N_9137);
and U10345 (N_10345,N_5732,N_9382);
nor U10346 (N_10346,N_9283,N_8253);
nand U10347 (N_10347,N_8215,N_7771);
or U10348 (N_10348,N_7484,N_9586);
or U10349 (N_10349,N_8866,N_8089);
and U10350 (N_10350,N_9748,N_8083);
xnor U10351 (N_10351,N_5553,N_6147);
nor U10352 (N_10352,N_6722,N_7258);
nor U10353 (N_10353,N_9875,N_8884);
and U10354 (N_10354,N_8357,N_7660);
or U10355 (N_10355,N_6257,N_8967);
or U10356 (N_10356,N_6592,N_6881);
nand U10357 (N_10357,N_8969,N_5030);
xor U10358 (N_10358,N_7154,N_6866);
nor U10359 (N_10359,N_7394,N_7062);
or U10360 (N_10360,N_8614,N_9502);
or U10361 (N_10361,N_9819,N_5619);
xor U10362 (N_10362,N_7815,N_5811);
nor U10363 (N_10363,N_6048,N_6347);
nor U10364 (N_10364,N_6402,N_6141);
xor U10365 (N_10365,N_7865,N_5346);
nand U10366 (N_10366,N_5919,N_5535);
nor U10367 (N_10367,N_7463,N_8986);
xnor U10368 (N_10368,N_9242,N_6496);
nand U10369 (N_10369,N_8628,N_5654);
xor U10370 (N_10370,N_7442,N_8316);
nor U10371 (N_10371,N_8992,N_5461);
and U10372 (N_10372,N_8985,N_9934);
xnor U10373 (N_10373,N_8728,N_7097);
nand U10374 (N_10374,N_7129,N_7499);
or U10375 (N_10375,N_7451,N_6799);
nand U10376 (N_10376,N_8843,N_7391);
nand U10377 (N_10377,N_6942,N_8247);
xor U10378 (N_10378,N_6951,N_6297);
or U10379 (N_10379,N_7197,N_7545);
xor U10380 (N_10380,N_6283,N_8526);
nand U10381 (N_10381,N_9642,N_5483);
nand U10382 (N_10382,N_5437,N_6301);
and U10383 (N_10383,N_9148,N_9008);
nor U10384 (N_10384,N_6329,N_5165);
xor U10385 (N_10385,N_7115,N_5893);
nor U10386 (N_10386,N_7929,N_5303);
nor U10387 (N_10387,N_5941,N_9418);
and U10388 (N_10388,N_8245,N_8404);
nor U10389 (N_10389,N_9633,N_5421);
nand U10390 (N_10390,N_7679,N_6512);
and U10391 (N_10391,N_6188,N_6156);
or U10392 (N_10392,N_6272,N_8211);
nor U10393 (N_10393,N_9417,N_6681);
xnor U10394 (N_10394,N_6370,N_9658);
and U10395 (N_10395,N_6530,N_7149);
nor U10396 (N_10396,N_8455,N_6171);
or U10397 (N_10397,N_5039,N_8132);
nand U10398 (N_10398,N_5019,N_5990);
or U10399 (N_10399,N_5186,N_9126);
and U10400 (N_10400,N_9821,N_8456);
nor U10401 (N_10401,N_7766,N_9167);
nand U10402 (N_10402,N_6620,N_9238);
and U10403 (N_10403,N_6699,N_7294);
xor U10404 (N_10404,N_8885,N_9800);
nor U10405 (N_10405,N_7602,N_5149);
or U10406 (N_10406,N_9007,N_9816);
nand U10407 (N_10407,N_8424,N_6229);
or U10408 (N_10408,N_5896,N_9540);
nor U10409 (N_10409,N_5426,N_5917);
nor U10410 (N_10410,N_9260,N_5387);
and U10411 (N_10411,N_7893,N_5209);
or U10412 (N_10412,N_9727,N_5327);
and U10413 (N_10413,N_9073,N_9813);
and U10414 (N_10414,N_8380,N_8420);
and U10415 (N_10415,N_9404,N_6163);
nand U10416 (N_10416,N_5280,N_9636);
and U10417 (N_10417,N_8154,N_6221);
and U10418 (N_10418,N_6192,N_9623);
and U10419 (N_10419,N_7235,N_7920);
nand U10420 (N_10420,N_9093,N_9603);
and U10421 (N_10421,N_5856,N_6473);
or U10422 (N_10422,N_5146,N_7159);
xor U10423 (N_10423,N_8694,N_8084);
and U10424 (N_10424,N_6814,N_7374);
nand U10425 (N_10425,N_5587,N_7289);
nor U10426 (N_10426,N_9098,N_7065);
nand U10427 (N_10427,N_8371,N_7859);
nor U10428 (N_10428,N_7382,N_9285);
nand U10429 (N_10429,N_8894,N_6602);
xor U10430 (N_10430,N_6357,N_6478);
or U10431 (N_10431,N_9610,N_6132);
nand U10432 (N_10432,N_6621,N_7286);
nand U10433 (N_10433,N_6487,N_5772);
nor U10434 (N_10434,N_8198,N_5659);
or U10435 (N_10435,N_5689,N_7858);
or U10436 (N_10436,N_7615,N_6225);
nor U10437 (N_10437,N_6310,N_5270);
nand U10438 (N_10438,N_7978,N_6892);
nor U10439 (N_10439,N_9174,N_8320);
and U10440 (N_10440,N_9588,N_6316);
nand U10441 (N_10441,N_8935,N_5516);
nor U10442 (N_10442,N_9994,N_9685);
and U10443 (N_10443,N_8358,N_7634);
nor U10444 (N_10444,N_7172,N_7012);
nand U10445 (N_10445,N_6217,N_9723);
xnor U10446 (N_10446,N_9657,N_6974);
xor U10447 (N_10447,N_5540,N_8716);
and U10448 (N_10448,N_5925,N_7714);
or U10449 (N_10449,N_6377,N_6870);
and U10450 (N_10450,N_9069,N_6006);
and U10451 (N_10451,N_5043,N_9643);
xnor U10452 (N_10452,N_6255,N_7184);
nor U10453 (N_10453,N_5372,N_8179);
or U10454 (N_10454,N_9836,N_9929);
and U10455 (N_10455,N_9110,N_9163);
and U10456 (N_10456,N_6686,N_7098);
or U10457 (N_10457,N_5182,N_7995);
or U10458 (N_10458,N_8849,N_6541);
xnor U10459 (N_10459,N_8997,N_8218);
xor U10460 (N_10460,N_7468,N_7415);
xnor U10461 (N_10461,N_8359,N_5510);
or U10462 (N_10462,N_6327,N_9829);
nor U10463 (N_10463,N_6660,N_5170);
and U10464 (N_10464,N_6026,N_6410);
or U10465 (N_10465,N_7591,N_9339);
and U10466 (N_10466,N_5971,N_9793);
nor U10467 (N_10467,N_8727,N_6052);
and U10468 (N_10468,N_6044,N_9589);
and U10469 (N_10469,N_7534,N_5664);
nand U10470 (N_10470,N_7009,N_7645);
or U10471 (N_10471,N_7874,N_9935);
nor U10472 (N_10472,N_9720,N_9330);
nand U10473 (N_10473,N_7847,N_6523);
and U10474 (N_10474,N_5364,N_6748);
nand U10475 (N_10475,N_8503,N_5730);
or U10476 (N_10476,N_5212,N_5452);
nand U10477 (N_10477,N_5000,N_8448);
xnor U10478 (N_10478,N_6148,N_9570);
or U10479 (N_10479,N_5879,N_9631);
or U10480 (N_10480,N_6028,N_6903);
and U10481 (N_10481,N_7952,N_5561);
or U10482 (N_10482,N_6927,N_6593);
xor U10483 (N_10483,N_8544,N_6544);
nand U10484 (N_10484,N_9889,N_6929);
xor U10485 (N_10485,N_9327,N_9475);
or U10486 (N_10486,N_9766,N_9244);
xor U10487 (N_10487,N_5101,N_7227);
nor U10488 (N_10488,N_9509,N_9872);
or U10489 (N_10489,N_5809,N_7183);
nand U10490 (N_10490,N_7840,N_5277);
or U10491 (N_10491,N_6358,N_9547);
nand U10492 (N_10492,N_5371,N_7113);
or U10493 (N_10493,N_5439,N_8221);
and U10494 (N_10494,N_5566,N_7427);
xor U10495 (N_10495,N_6424,N_5650);
or U10496 (N_10496,N_6597,N_7583);
and U10497 (N_10497,N_9409,N_8989);
or U10498 (N_10498,N_5686,N_9274);
xor U10499 (N_10499,N_7764,N_7095);
nor U10500 (N_10500,N_9313,N_8222);
nor U10501 (N_10501,N_9402,N_9638);
and U10502 (N_10502,N_6418,N_7477);
or U10503 (N_10503,N_6349,N_9139);
and U10504 (N_10504,N_7959,N_9788);
nand U10505 (N_10505,N_8942,N_8435);
or U10506 (N_10506,N_5604,N_5047);
xor U10507 (N_10507,N_9040,N_9597);
xnor U10508 (N_10508,N_9950,N_8595);
xnor U10509 (N_10509,N_7669,N_5211);
and U10510 (N_10510,N_6249,N_7074);
nand U10511 (N_10511,N_8955,N_6635);
and U10512 (N_10512,N_8620,N_9161);
nor U10513 (N_10513,N_6070,N_5631);
or U10514 (N_10514,N_9237,N_5611);
nor U10515 (N_10515,N_7407,N_9120);
nand U10516 (N_10516,N_9258,N_8336);
or U10517 (N_10517,N_9279,N_7271);
nand U10518 (N_10518,N_8260,N_7259);
nand U10519 (N_10519,N_9659,N_8605);
and U10520 (N_10520,N_5092,N_9023);
nor U10521 (N_10521,N_7036,N_8060);
nand U10522 (N_10522,N_6871,N_7016);
and U10523 (N_10523,N_7522,N_5172);
or U10524 (N_10524,N_6642,N_7939);
or U10525 (N_10525,N_9665,N_6467);
and U10526 (N_10526,N_8999,N_9615);
or U10527 (N_10527,N_9349,N_7228);
xnor U10528 (N_10528,N_6943,N_6067);
nor U10529 (N_10529,N_7122,N_8393);
nand U10530 (N_10530,N_9898,N_5472);
xor U10531 (N_10531,N_7802,N_5722);
nor U10532 (N_10532,N_8186,N_9546);
nor U10533 (N_10533,N_7002,N_5077);
or U10534 (N_10534,N_9049,N_9704);
or U10535 (N_10535,N_8951,N_9515);
or U10536 (N_10536,N_6745,N_5827);
nand U10537 (N_10537,N_5607,N_6172);
and U10538 (N_10538,N_7825,N_8641);
nand U10539 (N_10539,N_6925,N_8905);
and U10540 (N_10540,N_6749,N_8105);
or U10541 (N_10541,N_8704,N_6485);
xor U10542 (N_10542,N_5839,N_9992);
or U10543 (N_10543,N_7667,N_8837);
nand U10544 (N_10544,N_9201,N_5502);
or U10545 (N_10545,N_9538,N_7510);
nor U10546 (N_10546,N_6777,N_5748);
xnor U10547 (N_10547,N_8181,N_6047);
nand U10548 (N_10548,N_9550,N_6542);
nand U10549 (N_10549,N_6518,N_7439);
nor U10550 (N_10550,N_9182,N_8696);
and U10551 (N_10551,N_7275,N_9087);
and U10552 (N_10552,N_7711,N_5038);
and U10553 (N_10553,N_6431,N_9527);
xnor U10554 (N_10554,N_9399,N_9883);
or U10555 (N_10555,N_7726,N_7895);
or U10556 (N_10556,N_8433,N_8264);
nand U10557 (N_10557,N_9618,N_5287);
nand U10558 (N_10558,N_5681,N_5859);
or U10559 (N_10559,N_6437,N_6844);
nand U10560 (N_10560,N_5435,N_7153);
nand U10561 (N_10561,N_9751,N_7657);
nor U10562 (N_10562,N_5190,N_9188);
or U10563 (N_10563,N_7649,N_6277);
nand U10564 (N_10564,N_6190,N_6645);
or U10565 (N_10565,N_7402,N_8900);
nand U10566 (N_10566,N_8824,N_7021);
nand U10567 (N_10567,N_9810,N_5275);
nand U10568 (N_10568,N_6051,N_5606);
xor U10569 (N_10569,N_6096,N_6435);
nor U10570 (N_10570,N_8493,N_6150);
nand U10571 (N_10571,N_6835,N_7599);
nor U10572 (N_10572,N_8481,N_6114);
or U10573 (N_10573,N_5982,N_7392);
xnor U10574 (N_10574,N_6538,N_9140);
xor U10575 (N_10575,N_7872,N_5802);
nor U10576 (N_10576,N_5603,N_8067);
nor U10577 (N_10577,N_8096,N_6766);
xor U10578 (N_10578,N_5761,N_8408);
nor U10579 (N_10579,N_8069,N_9113);
nand U10580 (N_10580,N_8325,N_5002);
and U10581 (N_10581,N_8143,N_7479);
nand U10582 (N_10582,N_5608,N_5518);
nand U10583 (N_10583,N_9470,N_7829);
xor U10584 (N_10584,N_6103,N_5063);
nand U10585 (N_10585,N_8008,N_7863);
nand U10586 (N_10586,N_5008,N_6338);
and U10587 (N_10587,N_8530,N_8139);
xor U10588 (N_10588,N_9314,N_7215);
nor U10589 (N_10589,N_5972,N_6514);
nand U10590 (N_10590,N_6414,N_7204);
or U10591 (N_10591,N_5261,N_8982);
xor U10592 (N_10592,N_7552,N_7047);
nor U10593 (N_10593,N_8495,N_8003);
and U10594 (N_10594,N_7718,N_8057);
xnor U10595 (N_10595,N_9043,N_5677);
and U10596 (N_10596,N_8561,N_8484);
nand U10597 (N_10597,N_6412,N_5814);
nand U10598 (N_10598,N_7739,N_8324);
xor U10599 (N_10599,N_9301,N_7136);
nor U10600 (N_10600,N_7067,N_6199);
and U10601 (N_10601,N_8232,N_5852);
nor U10602 (N_10602,N_9598,N_8984);
xnor U10603 (N_10603,N_6661,N_7306);
nand U10604 (N_10604,N_6165,N_6804);
or U10605 (N_10605,N_8545,N_7921);
and U10606 (N_10606,N_6847,N_6480);
or U10607 (N_10607,N_9014,N_9850);
and U10608 (N_10608,N_9045,N_9378);
or U10609 (N_10609,N_5904,N_5843);
or U10610 (N_10610,N_9860,N_6719);
and U10611 (N_10611,N_8160,N_7769);
and U10612 (N_10612,N_7099,N_7256);
nor U10613 (N_10613,N_9516,N_9655);
nor U10614 (N_10614,N_8277,N_9369);
xor U10615 (N_10615,N_9719,N_6086);
nand U10616 (N_10616,N_6187,N_5339);
or U10617 (N_10617,N_5409,N_9996);
nand U10618 (N_10618,N_5203,N_7650);
and U10619 (N_10619,N_8693,N_8883);
and U10620 (N_10620,N_7092,N_5333);
or U10621 (N_10621,N_5083,N_8070);
nand U10622 (N_10622,N_9691,N_9428);
nand U10623 (N_10623,N_5289,N_7148);
or U10624 (N_10624,N_9969,N_8342);
nor U10625 (N_10625,N_9219,N_6622);
nand U10626 (N_10626,N_6970,N_6817);
nand U10627 (N_10627,N_7547,N_7348);
and U10628 (N_10628,N_5968,N_6898);
nand U10629 (N_10629,N_8622,N_8650);
and U10630 (N_10630,N_8609,N_5525);
and U10631 (N_10631,N_5599,N_7445);
or U10632 (N_10632,N_5018,N_8047);
or U10633 (N_10633,N_9577,N_5110);
nand U10634 (N_10634,N_9228,N_8496);
nor U10635 (N_10635,N_5986,N_8249);
or U10636 (N_10636,N_6331,N_6491);
xnor U10637 (N_10637,N_6755,N_5714);
and U10638 (N_10638,N_9835,N_7811);
or U10639 (N_10639,N_9460,N_9071);
nand U10640 (N_10640,N_6940,N_6899);
nand U10641 (N_10641,N_6526,N_9440);
xnor U10642 (N_10642,N_5430,N_9518);
or U10643 (N_10643,N_9874,N_7112);
nor U10644 (N_10644,N_5393,N_5594);
and U10645 (N_10645,N_7412,N_6983);
or U10646 (N_10646,N_9982,N_9080);
or U10647 (N_10647,N_7656,N_6488);
or U10648 (N_10648,N_6641,N_5756);
and U10649 (N_10649,N_8801,N_5590);
or U10650 (N_10650,N_5102,N_5787);
or U10651 (N_10651,N_5312,N_8250);
nor U10652 (N_10652,N_5307,N_9297);
xnor U10653 (N_10653,N_9840,N_6454);
nand U10654 (N_10654,N_6775,N_9805);
xor U10655 (N_10655,N_6972,N_8919);
nand U10656 (N_10656,N_9629,N_8228);
nand U10657 (N_10657,N_5045,N_6825);
xor U10658 (N_10658,N_7166,N_9304);
nor U10659 (N_10659,N_8625,N_8524);
nor U10660 (N_10660,N_6376,N_8771);
xnor U10661 (N_10661,N_8381,N_9713);
xor U10662 (N_10662,N_8812,N_9222);
xnor U10663 (N_10663,N_7827,N_5104);
and U10664 (N_10664,N_5703,N_8521);
xnor U10665 (N_10665,N_8591,N_5184);
and U10666 (N_10666,N_5870,N_9880);
xnor U10667 (N_10667,N_8214,N_5774);
and U10668 (N_10668,N_7700,N_7915);
nor U10669 (N_10669,N_9806,N_6574);
nor U10670 (N_10670,N_7885,N_8192);
and U10671 (N_10671,N_7426,N_6957);
nor U10672 (N_10672,N_8808,N_6037);
nand U10673 (N_10673,N_5225,N_8487);
xor U10674 (N_10674,N_6371,N_8429);
or U10675 (N_10675,N_5536,N_8278);
xnor U10676 (N_10676,N_6789,N_9571);
xnor U10677 (N_10677,N_7147,N_9457);
nand U10678 (N_10678,N_9822,N_9090);
and U10679 (N_10679,N_7659,N_9159);
nand U10680 (N_10680,N_7436,N_8030);
xor U10681 (N_10681,N_6758,N_8665);
nor U10682 (N_10682,N_5555,N_5956);
and U10683 (N_10683,N_9379,N_5230);
and U10684 (N_10684,N_6326,N_5467);
and U10685 (N_10685,N_8550,N_6393);
and U10686 (N_10686,N_5413,N_8705);
nand U10687 (N_10687,N_7878,N_8842);
xnor U10688 (N_10688,N_8947,N_7988);
and U10689 (N_10689,N_5942,N_5861);
xnor U10690 (N_10690,N_5479,N_7834);
nand U10691 (N_10691,N_8823,N_9966);
nor U10692 (N_10692,N_5194,N_7804);
nand U10693 (N_10693,N_8819,N_5004);
nand U10694 (N_10694,N_5757,N_7741);
nand U10695 (N_10695,N_7715,N_8949);
xnor U10696 (N_10696,N_5963,N_6280);
or U10697 (N_10697,N_7464,N_6273);
and U10698 (N_10698,N_7944,N_6861);
and U10699 (N_10699,N_8923,N_5174);
nand U10700 (N_10700,N_8108,N_8476);
nand U10701 (N_10701,N_5877,N_7633);
nor U10702 (N_10702,N_7695,N_6715);
xnor U10703 (N_10703,N_8355,N_7390);
nor U10704 (N_10704,N_7006,N_6101);
xnor U10705 (N_10705,N_5936,N_5199);
nor U10706 (N_10706,N_5754,N_9856);
or U10707 (N_10707,N_8560,N_7922);
nor U10708 (N_10708,N_5764,N_6603);
xnor U10709 (N_10709,N_8216,N_9267);
and U10710 (N_10710,N_8306,N_8243);
nor U10711 (N_10711,N_6605,N_6615);
xnor U10712 (N_10712,N_9187,N_9958);
xor U10713 (N_10713,N_5653,N_5296);
or U10714 (N_10714,N_5021,N_5499);
nor U10715 (N_10715,N_6717,N_5103);
xnor U10716 (N_10716,N_8556,N_8230);
xnor U10717 (N_10717,N_6152,N_7123);
xor U10718 (N_10718,N_5228,N_7063);
nand U10719 (N_10719,N_9863,N_6110);
nand U10720 (N_10720,N_6604,N_6548);
and U10721 (N_10721,N_7856,N_9791);
and U10722 (N_10722,N_8525,N_8594);
or U10723 (N_10723,N_9186,N_6493);
or U10724 (N_10724,N_5912,N_8379);
xor U10725 (N_10725,N_9949,N_8834);
or U10726 (N_10726,N_6017,N_7052);
or U10727 (N_10727,N_5678,N_9370);
nor U10728 (N_10728,N_7251,N_9903);
xor U10729 (N_10729,N_5929,N_5881);
and U10730 (N_10730,N_5642,N_8136);
nand U10731 (N_10731,N_5123,N_7616);
xor U10732 (N_10732,N_6483,N_5222);
xnor U10733 (N_10733,N_6462,N_9913);
and U10734 (N_10734,N_8400,N_7573);
nor U10735 (N_10735,N_6285,N_9500);
xnor U10736 (N_10736,N_6894,N_7728);
or U10737 (N_10737,N_8056,N_6678);
or U10738 (N_10738,N_8621,N_8793);
xor U10739 (N_10739,N_8411,N_6811);
xnor U10740 (N_10740,N_5849,N_5412);
xnor U10741 (N_10741,N_6633,N_5808);
nand U10742 (N_10742,N_8559,N_6584);
and U10743 (N_10743,N_5323,N_5720);
xor U10744 (N_10744,N_5775,N_9375);
nand U10745 (N_10745,N_8011,N_7000);
or U10746 (N_10746,N_8895,N_5530);
nor U10747 (N_10747,N_5613,N_9683);
or U10748 (N_10748,N_9012,N_7828);
nand U10749 (N_10749,N_6243,N_6908);
nor U10750 (N_10750,N_7195,N_5625);
nor U10751 (N_10751,N_9367,N_8163);
or U10752 (N_10752,N_9492,N_6572);
nand U10753 (N_10753,N_5181,N_5696);
and U10754 (N_10754,N_9425,N_7710);
xor U10755 (N_10755,N_8554,N_6469);
and U10756 (N_10756,N_6098,N_6683);
nand U10757 (N_10757,N_9125,N_7341);
xnor U10758 (N_10758,N_9352,N_5402);
and U10759 (N_10759,N_5511,N_5281);
nor U10760 (N_10760,N_6577,N_7750);
nand U10761 (N_10761,N_6422,N_8274);
nor U10762 (N_10762,N_5672,N_5688);
nand U10763 (N_10763,N_9673,N_8678);
nand U10764 (N_10764,N_6980,N_6282);
and U10765 (N_10765,N_9116,N_5838);
nor U10766 (N_10766,N_8791,N_9943);
and U10767 (N_10767,N_5830,N_6918);
nor U10768 (N_10768,N_8798,N_6585);
nand U10769 (N_10769,N_8721,N_7805);
nand U10770 (N_10770,N_7946,N_8311);
nor U10771 (N_10771,N_9439,N_7375);
and U10772 (N_10772,N_5446,N_8611);
nor U10773 (N_10773,N_8707,N_5141);
or U10774 (N_10774,N_6505,N_5326);
xor U10775 (N_10775,N_6034,N_5057);
or U10776 (N_10776,N_9814,N_5302);
and U10777 (N_10777,N_6631,N_5420);
nand U10778 (N_10778,N_8901,N_7932);
xnor U10779 (N_10779,N_9654,N_9894);
xnor U10780 (N_10780,N_7800,N_9394);
xnor U10781 (N_10781,N_9337,N_6813);
and U10782 (N_10782,N_9947,N_9847);
nand U10783 (N_10783,N_5069,N_8933);
or U10784 (N_10784,N_8981,N_8147);
or U10785 (N_10785,N_6007,N_9216);
or U10786 (N_10786,N_6268,N_9828);
nor U10787 (N_10787,N_9001,N_6937);
or U10788 (N_10788,N_8078,N_5064);
nand U10789 (N_10789,N_5089,N_7822);
or U10790 (N_10790,N_7179,N_8199);
nor U10791 (N_10791,N_6464,N_9747);
nor U10792 (N_10792,N_7844,N_6009);
nand U10793 (N_10793,N_9089,N_8551);
nand U10794 (N_10794,N_8155,N_7471);
nor U10795 (N_10795,N_5778,N_9421);
or U10796 (N_10796,N_9081,N_7749);
nand U10797 (N_10797,N_9979,N_5655);
and U10798 (N_10798,N_8256,N_7954);
or U10799 (N_10799,N_9121,N_8102);
or U10800 (N_10800,N_7991,N_9247);
xnor U10801 (N_10801,N_7287,N_7569);
xnor U10802 (N_10802,N_7851,N_9333);
or U10803 (N_10803,N_8395,N_5749);
or U10804 (N_10804,N_5142,N_6019);
xor U10805 (N_10805,N_6941,N_5396);
and U10806 (N_10806,N_8281,N_5648);
or U10807 (N_10807,N_6860,N_6565);
or U10808 (N_10808,N_7504,N_6969);
xor U10809 (N_10809,N_8975,N_9679);
and U10810 (N_10810,N_6288,N_9145);
or U10811 (N_10811,N_9674,N_7200);
nor U10812 (N_10812,N_5679,N_8236);
or U10813 (N_10813,N_8035,N_6590);
or U10814 (N_10814,N_8439,N_6805);
nand U10815 (N_10815,N_5837,N_7027);
xnor U10816 (N_10816,N_9767,N_7330);
nor U10817 (N_10817,N_7557,N_7048);
nor U10818 (N_10818,N_7131,N_7612);
nand U10819 (N_10819,N_8597,N_9652);
nor U10820 (N_10820,N_6606,N_7140);
or U10821 (N_10821,N_6591,N_5969);
nor U10822 (N_10822,N_8723,N_7416);
or U10823 (N_10823,N_8298,N_5470);
xor U10824 (N_10824,N_7059,N_6416);
nor U10825 (N_10825,N_6245,N_8911);
xor U10826 (N_10826,N_7304,N_7793);
and U10827 (N_10827,N_6529,N_7485);
nor U10828 (N_10828,N_9150,N_9076);
and U10829 (N_10829,N_7010,N_9365);
nor U10830 (N_10830,N_5345,N_6930);
or U10831 (N_10831,N_8733,N_6516);
nand U10832 (N_10832,N_7364,N_5628);
nor U10833 (N_10833,N_7948,N_6938);
or U10834 (N_10834,N_8310,N_9449);
or U10835 (N_10835,N_6554,N_5669);
or U10836 (N_10836,N_6262,N_9151);
xor U10837 (N_10837,N_7100,N_9690);
and U10838 (N_10838,N_9986,N_7189);
or U10839 (N_10839,N_7379,N_8300);
nor U10840 (N_10840,N_8234,N_8262);
or U10841 (N_10841,N_6883,N_6382);
and U10842 (N_10842,N_7810,N_8294);
and U10843 (N_10843,N_7116,N_8335);
or U10844 (N_10844,N_8897,N_5493);
nor U10845 (N_10845,N_9252,N_7806);
nand U10846 (N_10846,N_8587,N_8172);
xor U10847 (N_10847,N_8888,N_9353);
and U10848 (N_10848,N_8976,N_5712);
and U10849 (N_10849,N_9901,N_6074);
and U10850 (N_10850,N_9532,N_7933);
nand U10851 (N_10851,N_9092,N_6773);
nand U10852 (N_10852,N_9020,N_7058);
or U10853 (N_10853,N_9046,N_6296);
or U10854 (N_10854,N_9346,N_9861);
and U10855 (N_10855,N_5138,N_9465);
nor U10856 (N_10856,N_5746,N_8724);
or U10857 (N_10857,N_6687,N_6474);
nand U10858 (N_10858,N_5143,N_6684);
nor U10859 (N_10859,N_5091,N_5575);
xnor U10860 (N_10860,N_6788,N_7467);
and U10861 (N_10861,N_8898,N_9374);
and U10862 (N_10862,N_9495,N_5410);
and U10863 (N_10863,N_6993,N_5490);
nand U10864 (N_10864,N_9055,N_7773);
and U10865 (N_10865,N_6846,N_5158);
or U10866 (N_10866,N_5324,N_9650);
or U10867 (N_10867,N_6302,N_7625);
xnor U10868 (N_10868,N_9249,N_5868);
or U10869 (N_10869,N_7237,N_7269);
or U10870 (N_10870,N_5443,N_9553);
xor U10871 (N_10871,N_5853,N_7384);
xnor U10872 (N_10872,N_5256,N_9548);
and U10873 (N_10873,N_5533,N_6275);
xnor U10874 (N_10874,N_9082,N_9776);
and U10875 (N_10875,N_8326,N_5509);
and U10876 (N_10876,N_7527,N_7732);
nor U10877 (N_10877,N_9520,N_5072);
and U10878 (N_10878,N_5926,N_5398);
and U10879 (N_10879,N_5620,N_9442);
nor U10880 (N_10880,N_8788,N_5586);
nor U10881 (N_10881,N_7295,N_7965);
nor U10882 (N_10882,N_5898,N_7054);
xor U10883 (N_10883,N_9462,N_8968);
or U10884 (N_10884,N_5989,N_6977);
and U10885 (N_10885,N_5668,N_8886);
xor U10886 (N_10886,N_8957,N_5682);
nor U10887 (N_10887,N_7623,N_5932);
xnor U10888 (N_10888,N_6064,N_6463);
nor U10889 (N_10889,N_6989,N_7653);
nand U10890 (N_10890,N_7775,N_9694);
or U10891 (N_10891,N_6220,N_8831);
or U10892 (N_10892,N_5901,N_6340);
and U10893 (N_10893,N_6754,N_6368);
and U10894 (N_10894,N_5188,N_8692);
nand U10895 (N_10895,N_7472,N_7162);
nor U10896 (N_10896,N_5875,N_9736);
or U10897 (N_10897,N_8246,N_9316);
xnor U10898 (N_10898,N_5457,N_9368);
nand U10899 (N_10899,N_7417,N_6956);
nand U10900 (N_10900,N_7061,N_7234);
nand U10901 (N_10901,N_6637,N_5052);
and U10902 (N_10902,N_9197,N_7476);
nand U10903 (N_10903,N_5292,N_7670);
and U10904 (N_10904,N_8385,N_5948);
and U10905 (N_10905,N_6345,N_7339);
nand U10906 (N_10906,N_7817,N_5207);
nand U10907 (N_10907,N_9666,N_5740);
and U10908 (N_10908,N_7853,N_5977);
nor U10909 (N_10909,N_6334,N_5465);
or U10910 (N_10910,N_6662,N_8226);
xor U10911 (N_10911,N_9905,N_8536);
and U10912 (N_10912,N_8757,N_5460);
nor U10913 (N_10913,N_5352,N_7785);
xnor U10914 (N_10914,N_8492,N_9775);
or U10915 (N_10915,N_7165,N_8091);
or U10916 (N_10916,N_7437,N_8731);
and U10917 (N_10917,N_8657,N_9340);
nor U10918 (N_10918,N_8178,N_7884);
and U10919 (N_10919,N_6151,N_6962);
xor U10920 (N_10920,N_9318,N_8183);
and U10921 (N_10921,N_6451,N_9759);
nand U10922 (N_10922,N_5136,N_6960);
xor U10923 (N_10923,N_8847,N_9605);
nand U10924 (N_10924,N_6543,N_6978);
or U10925 (N_10925,N_7085,N_7542);
nand U10926 (N_10926,N_9941,N_8286);
or U10927 (N_10927,N_9773,N_9656);
or U10928 (N_10928,N_9998,N_9355);
xnor U10929 (N_10929,N_8144,N_5032);
and U10930 (N_10930,N_5883,N_5541);
xor U10931 (N_10931,N_7401,N_9761);
and U10932 (N_10932,N_5503,N_6456);
or U10933 (N_10933,N_6361,N_7531);
nor U10934 (N_10934,N_9914,N_6569);
nor U10935 (N_10935,N_7461,N_5800);
and U10936 (N_10936,N_6281,N_6428);
nor U10937 (N_10937,N_8537,N_6490);
xor U10938 (N_10938,N_8037,N_7632);
and U10939 (N_10939,N_9795,N_9939);
xnor U10940 (N_10940,N_6778,N_5340);
and U10941 (N_10941,N_5382,N_8637);
or U10942 (N_10942,N_5108,N_8643);
nor U10943 (N_10943,N_9048,N_8756);
or U10944 (N_10944,N_6260,N_7529);
xor U10945 (N_10945,N_7344,N_5612);
xnor U10946 (N_10946,N_5637,N_8783);
xor U10947 (N_10947,N_5676,N_6312);
nor U10948 (N_10948,N_6015,N_7232);
xor U10949 (N_10949,N_9858,N_5684);
or U10950 (N_10950,N_8273,N_5109);
nand U10951 (N_10951,N_5766,N_6216);
nand U10952 (N_10952,N_7925,N_7393);
or U10953 (N_10953,N_5090,N_5135);
or U10954 (N_10954,N_5552,N_5252);
or U10955 (N_10955,N_6089,N_7060);
nor U10956 (N_10956,N_8811,N_7664);
and U10957 (N_10957,N_7736,N_7593);
nand U10958 (N_10958,N_8059,N_6531);
xnor U10959 (N_10959,N_6812,N_5913);
or U10960 (N_10960,N_5662,N_9013);
and U10961 (N_10961,N_9176,N_7443);
nor U10962 (N_10962,N_5310,N_9646);
nor U10963 (N_10963,N_6167,N_5887);
nand U10964 (N_10964,N_7770,N_7220);
nand U10965 (N_10965,N_8972,N_9574);
xnor U10966 (N_10966,N_6430,N_5159);
nor U10967 (N_10967,N_6224,N_9084);
nand U10968 (N_10968,N_7264,N_6786);
nand U10969 (N_10969,N_6471,N_5233);
nor U10970 (N_10970,N_6760,N_9494);
xor U10971 (N_10971,N_9818,N_8661);
and U10972 (N_10972,N_5054,N_8167);
nand U10973 (N_10973,N_5450,N_7150);
xor U10974 (N_10974,N_9519,N_7721);
xnor U10975 (N_10975,N_8410,N_5355);
or U10976 (N_10976,N_5953,N_7759);
or U10977 (N_10977,N_7208,N_6685);
nand U10978 (N_10978,N_8821,N_8563);
and U10979 (N_10979,N_8785,N_8158);
or U10980 (N_10980,N_9796,N_8816);
and U10981 (N_10981,N_5979,N_6834);
nor U10982 (N_10982,N_7424,N_8169);
or U10983 (N_10983,N_5760,N_8080);
xor U10984 (N_10984,N_7592,N_6934);
nor U10985 (N_10985,N_6391,N_7045);
nor U10986 (N_10986,N_9175,N_5624);
xor U10987 (N_10987,N_9983,N_8874);
xnor U10988 (N_10988,N_6091,N_6886);
nor U10989 (N_10989,N_7023,N_8763);
xor U10990 (N_10990,N_7820,N_7170);
or U10991 (N_10991,N_8165,N_7196);
nand U10992 (N_10992,N_6266,N_9717);
xnor U10993 (N_10993,N_9364,N_5321);
and U10994 (N_10994,N_5168,N_7869);
or U10995 (N_10995,N_8922,N_7498);
or U10996 (N_10996,N_8284,N_6429);
or U10997 (N_10997,N_6623,N_8659);
or U10998 (N_10998,N_7222,N_6657);
nand U10999 (N_10999,N_5713,N_6629);
xnor U11000 (N_11000,N_9130,N_7020);
and U11001 (N_11001,N_6372,N_5394);
and U11002 (N_11002,N_5074,N_7693);
nor U11003 (N_11003,N_7176,N_8129);
or U11004 (N_11004,N_7107,N_7262);
xnor U11005 (N_11005,N_5562,N_6038);
and U11006 (N_11006,N_5539,N_7892);
xor U11007 (N_11007,N_8764,N_9405);
nand U11008 (N_11008,N_9415,N_9109);
and U11009 (N_11009,N_9724,N_8658);
or U11010 (N_11010,N_7329,N_8988);
xor U11011 (N_11011,N_8113,N_5070);
and U11012 (N_11012,N_9817,N_6185);
nand U11013 (N_11013,N_7422,N_6191);
and U11014 (N_11014,N_9948,N_7114);
nand U11015 (N_11015,N_7690,N_8577);
or U11016 (N_11016,N_8913,N_8261);
or U11017 (N_11017,N_9393,N_6895);
or U11018 (N_11018,N_6309,N_8624);
nor U11019 (N_11019,N_7513,N_8193);
xor U11020 (N_11020,N_5244,N_6831);
or U11021 (N_11021,N_9584,N_9954);
or U11022 (N_11022,N_6390,N_6443);
and U11023 (N_11023,N_6876,N_7913);
and U11024 (N_11024,N_7126,N_5315);
xor U11025 (N_11025,N_9525,N_5846);
nor U11026 (N_11026,N_8833,N_5951);
nand U11027 (N_11027,N_5573,N_8858);
and U11028 (N_11028,N_9290,N_8112);
nor U11029 (N_11029,N_5369,N_6121);
nand U11030 (N_11030,N_8474,N_8632);
xor U11031 (N_11031,N_6438,N_9443);
and U11032 (N_11032,N_9677,N_7157);
or U11033 (N_11033,N_5206,N_7017);
nand U11034 (N_11034,N_7057,N_7226);
or U11035 (N_11035,N_6521,N_9178);
nor U11036 (N_11036,N_8845,N_6123);
or U11037 (N_11037,N_5667,N_9282);
xor U11038 (N_11038,N_6013,N_6419);
and U11039 (N_11039,N_5831,N_9892);
or U11040 (N_11040,N_6757,N_7846);
or U11041 (N_11041,N_6578,N_7704);
xor U11042 (N_11042,N_9801,N_6100);
nand U11043 (N_11043,N_8427,N_6498);
and U11044 (N_11044,N_8878,N_6988);
nor U11045 (N_11045,N_6112,N_5649);
xor U11046 (N_11046,N_8979,N_6724);
or U11047 (N_11047,N_5082,N_5217);
or U11048 (N_11048,N_7194,N_5076);
xor U11049 (N_11049,N_9412,N_6440);
or U11050 (N_11050,N_9233,N_7175);
or U11051 (N_11051,N_9881,N_7525);
nand U11052 (N_11052,N_5900,N_8674);
nor U11053 (N_11053,N_7096,N_7651);
nor U11054 (N_11054,N_7032,N_9912);
and U11055 (N_11055,N_5762,N_5916);
and U11056 (N_11056,N_9251,N_6547);
or U11057 (N_11057,N_8864,N_5743);
nand U11058 (N_11058,N_7404,N_7683);
and U11059 (N_11059,N_6596,N_6264);
xnor U11060 (N_11060,N_5298,N_6293);
xor U11061 (N_11061,N_8094,N_5226);
xor U11062 (N_11062,N_7608,N_5692);
or U11063 (N_11063,N_5105,N_5191);
xor U11064 (N_11064,N_8867,N_7654);
and U11065 (N_11065,N_7938,N_9815);
xor U11066 (N_11066,N_9620,N_8350);
nor U11067 (N_11067,N_7068,N_6772);
nand U11068 (N_11068,N_8546,N_8714);
and U11069 (N_11069,N_5305,N_6999);
or U11070 (N_11070,N_9625,N_8423);
and U11071 (N_11071,N_7318,N_8737);
nor U11072 (N_11072,N_5609,N_9552);
or U11073 (N_11073,N_6537,N_5376);
and U11074 (N_11074,N_7686,N_7967);
xor U11075 (N_11075,N_6324,N_5961);
xor U11076 (N_11076,N_5469,N_8954);
nor U11077 (N_11077,N_7371,N_5683);
or U11078 (N_11078,N_7774,N_5790);
or U11079 (N_11079,N_6600,N_8519);
xnor U11080 (N_11080,N_9331,N_6115);
nor U11081 (N_11081,N_7691,N_5279);
and U11082 (N_11082,N_7325,N_8702);
and U11083 (N_11083,N_9575,N_9945);
or U11084 (N_11084,N_6540,N_5375);
nor U11085 (N_11085,N_5867,N_5097);
nor U11086 (N_11086,N_7143,N_6479);
nor U11087 (N_11087,N_7998,N_8510);
xor U11088 (N_11088,N_5807,N_6196);
xnor U11089 (N_11089,N_9229,N_8054);
nand U11090 (N_11090,N_9989,N_8437);
and U11091 (N_11091,N_6998,N_9928);
xor U11092 (N_11092,N_6862,N_6837);
or U11093 (N_11093,N_7385,N_7536);
xnor U11094 (N_11094,N_8398,N_9757);
xnor U11095 (N_11095,N_9134,N_6155);
nor U11096 (N_11096,N_9232,N_8945);
xnor U11097 (N_11097,N_9256,N_8863);
xor U11098 (N_11098,N_7119,N_8533);
nor U11099 (N_11099,N_7128,N_5670);
or U11100 (N_11100,N_7701,N_8795);
nor U11101 (N_11101,N_9678,N_8680);
xor U11102 (N_11102,N_6872,N_9193);
and U11103 (N_11103,N_6383,N_6618);
xnor U11104 (N_11104,N_6153,N_5909);
or U11105 (N_11105,N_9728,N_5354);
nand U11106 (N_11106,N_6727,N_6108);
nand U11107 (N_11107,N_5579,N_9292);
and U11108 (N_11108,N_6822,N_6954);
or U11109 (N_11109,N_5949,N_8053);
nand U11110 (N_11110,N_5495,N_5895);
and U11111 (N_11111,N_8356,N_7279);
and U11112 (N_11112,N_9565,N_5094);
nand U11113 (N_11113,N_8760,N_8097);
nor U11114 (N_11114,N_9867,N_6012);
nor U11115 (N_11115,N_8924,N_5432);
and U11116 (N_11116,N_9893,N_7301);
xor U11117 (N_11117,N_8656,N_9005);
xnor U11118 (N_11118,N_5405,N_8241);
xor U11119 (N_11119,N_9528,N_6214);
nor U11120 (N_11120,N_9106,N_7879);
or U11121 (N_11121,N_9853,N_7008);
nand U11122 (N_11122,N_9541,N_7707);
nand U11123 (N_11123,N_9416,N_5974);
nor U11124 (N_11124,N_5836,N_7843);
and U11125 (N_11125,N_5485,N_5884);
nor U11126 (N_11126,N_5401,N_5500);
xnor U11127 (N_11127,N_6619,N_9359);
and U11128 (N_11128,N_5475,N_8780);
or U11129 (N_11129,N_8482,N_6063);
and U11130 (N_11130,N_9647,N_8926);
and U11131 (N_11131,N_9873,N_8283);
and U11132 (N_11132,N_9255,N_7706);
nand U11133 (N_11133,N_9635,N_7937);
and U11134 (N_11134,N_8779,N_7723);
nor U11135 (N_11135,N_5012,N_8159);
nand U11136 (N_11136,N_5041,N_7218);
xor U11137 (N_11137,N_6219,N_8392);
xor U11138 (N_11138,N_6982,N_7414);
xnor U11139 (N_11139,N_5581,N_5646);
and U11140 (N_11140,N_7808,N_8450);
or U11141 (N_11141,N_7470,N_6639);
or U11142 (N_11142,N_8019,N_5610);
nor U11143 (N_11143,N_7618,N_8267);
nor U11144 (N_11144,N_7523,N_8021);
and U11145 (N_11145,N_5554,N_8664);
and U11146 (N_11146,N_6880,N_5258);
xnor U11147 (N_11147,N_5319,N_8566);
nor U11148 (N_11148,N_6840,N_8840);
xnor U11149 (N_11149,N_8806,N_5717);
nor U11150 (N_11150,N_6355,N_5600);
or U11151 (N_11151,N_6830,N_9595);
and U11152 (N_11152,N_9746,N_8133);
nor U11153 (N_11153,N_9498,N_8729);
nand U11154 (N_11154,N_7857,N_6475);
or U11155 (N_11155,N_9042,N_9235);
or U11156 (N_11156,N_8996,N_8036);
nor U11157 (N_11157,N_6752,N_6566);
xor U11158 (N_11158,N_7540,N_7338);
xnor U11159 (N_11159,N_6265,N_6295);
xnor U11160 (N_11160,N_8210,N_6935);
xor U11161 (N_11161,N_8340,N_7387);
nand U11162 (N_11162,N_6853,N_9062);
nand U11163 (N_11163,N_5466,N_8088);
xnor U11164 (N_11164,N_8523,N_9491);
or U11165 (N_11165,N_8265,N_8686);
xnor U11166 (N_11166,N_7446,N_9972);
and U11167 (N_11167,N_7242,N_8099);
or U11168 (N_11168,N_9511,N_9499);
xnor U11169 (N_11169,N_9743,N_5569);
nand U11170 (N_11170,N_6869,N_8616);
nor U11171 (N_11171,N_6583,N_6267);
xnor U11172 (N_11172,N_9681,N_8348);
nand U11173 (N_11173,N_6964,N_5079);
or U11174 (N_11174,N_9397,N_8937);
xnor U11175 (N_11175,N_9513,N_7894);
xor U11176 (N_11176,N_6195,N_6730);
or U11177 (N_11177,N_8301,N_9955);
xor U11178 (N_11178,N_6634,N_9722);
xor U11179 (N_11179,N_9438,N_5350);
xor U11180 (N_11180,N_5121,N_5529);
nor U11181 (N_11181,N_8740,N_6335);
nor U11182 (N_11182,N_6958,N_5017);
nor U11183 (N_11183,N_5368,N_5880);
and U11184 (N_11184,N_8775,N_6279);
and U11185 (N_11185,N_8363,N_6561);
nand U11186 (N_11186,N_8026,N_7481);
xor U11187 (N_11187,N_9687,N_7042);
nand U11188 (N_11188,N_5685,N_9230);
and U11189 (N_11189,N_6090,N_8725);
and U11190 (N_11190,N_6084,N_6986);
xor U11191 (N_11191,N_8592,N_5813);
xor U11192 (N_11192,N_5551,N_8679);
nand U11193 (N_11193,N_8856,N_5994);
nor U11194 (N_11194,N_5118,N_9464);
nor U11195 (N_11195,N_6387,N_5389);
nand U11196 (N_11196,N_5318,N_9888);
xnor U11197 (N_11197,N_7395,N_6484);
nand U11198 (N_11198,N_7308,N_9940);
xnor U11199 (N_11199,N_8092,N_7551);
and U11200 (N_11200,N_7408,N_9675);
nand U11201 (N_11201,N_5059,N_6947);
and U11202 (N_11202,N_6863,N_5208);
and U11203 (N_11203,N_8289,N_5088);
or U11204 (N_11204,N_8436,N_6611);
nor U11205 (N_11205,N_7596,N_9846);
xnor U11206 (N_11206,N_9859,N_9700);
nor U11207 (N_11207,N_6933,N_6690);
xnor U11208 (N_11208,N_9243,N_5160);
and U11209 (N_11209,N_5512,N_9613);
and U11210 (N_11210,N_9834,N_6076);
or U11211 (N_11211,N_5050,N_6477);
xnor U11212 (N_11212,N_5824,N_6392);
and U11213 (N_11213,N_9697,N_5750);
or U11214 (N_11214,N_7033,N_6668);
nand U11215 (N_11215,N_7312,N_8630);
nand U11216 (N_11216,N_6793,N_6319);
nand U11217 (N_11217,N_9044,N_8906);
or U11218 (N_11218,N_7575,N_8134);
nand U11219 (N_11219,N_5497,N_6843);
and U11220 (N_11220,N_6905,N_6222);
nor U11221 (N_11221,N_8065,N_8598);
nor U11222 (N_11222,N_6401,N_6494);
xor U11223 (N_11223,N_6651,N_8440);
or U11224 (N_11224,N_5770,N_7638);
and U11225 (N_11225,N_9231,N_5576);
xnor U11226 (N_11226,N_9319,N_5205);
nor U11227 (N_11227,N_8016,N_6081);
nand U11228 (N_11228,N_7500,N_7400);
and U11229 (N_11229,N_9770,N_5582);
nor U11230 (N_11230,N_6979,N_7908);
or U11231 (N_11231,N_9651,N_5379);
or U11232 (N_11232,N_8796,N_6700);
nand U11233 (N_11233,N_9454,N_7240);
or U11234 (N_11234,N_7905,N_7310);
and U11235 (N_11235,N_5726,N_7977);
and U11236 (N_11236,N_8829,N_5765);
and U11237 (N_11237,N_9729,N_5322);
nand U11238 (N_11238,N_9338,N_6740);
or U11239 (N_11239,N_8893,N_8854);
nand U11240 (N_11240,N_9804,N_8688);
nand U11241 (N_11241,N_6601,N_5776);
and U11242 (N_11242,N_6218,N_8745);
nor U11243 (N_11243,N_7249,N_7642);
nor U11244 (N_11244,N_6653,N_7772);
or U11245 (N_11245,N_6011,N_6023);
nor U11246 (N_11246,N_8564,N_7609);
nor U11247 (N_11247,N_7797,N_9811);
and U11248 (N_11248,N_7080,N_8899);
xnor U11249 (N_11249,N_7819,N_6244);
nand U11250 (N_11250,N_5878,N_8117);
nor U11251 (N_11251,N_8499,N_5806);
or U11252 (N_11252,N_5314,N_5316);
and U11253 (N_11253,N_6291,N_9789);
and U11254 (N_11254,N_9104,N_7942);
and U11255 (N_11255,N_5177,N_7541);
and U11256 (N_11256,N_7871,N_7438);
nand U11257 (N_11257,N_7121,N_6608);
or U11258 (N_11258,N_5680,N_7584);
and U11259 (N_11259,N_6515,N_6364);
and U11260 (N_11260,N_5468,N_5390);
xnor U11261 (N_11261,N_6113,N_5593);
and U11262 (N_11262,N_7246,N_6235);
nand U11263 (N_11263,N_7450,N_8751);
xor U11264 (N_11264,N_6169,N_7719);
xnor U11265 (N_11265,N_6164,N_8354);
or U11266 (N_11266,N_6695,N_7124);
nand U11267 (N_11267,N_9431,N_8639);
or U11268 (N_11268,N_8720,N_5645);
or U11269 (N_11269,N_9566,N_5621);
xnor U11270 (N_11270,N_8469,N_6845);
nor U11271 (N_11271,N_5797,N_6189);
and U11272 (N_11272,N_6627,N_8238);
nand U11273 (N_11273,N_8150,N_6701);
nand U11274 (N_11274,N_9474,N_7521);
nand U11275 (N_11275,N_8066,N_8349);
nand U11276 (N_11276,N_9698,N_9018);
and U11277 (N_11277,N_8601,N_6226);
and U11278 (N_11278,N_7713,N_7784);
and U11279 (N_11279,N_9391,N_6294);
and U11280 (N_11280,N_6299,N_9803);
nand U11281 (N_11281,N_5474,N_8090);
and U11282 (N_11282,N_6043,N_8498);
xnor U11283 (N_11283,N_9129,N_5433);
and U11284 (N_11284,N_8344,N_9871);
or U11285 (N_11285,N_9272,N_5351);
and U11286 (N_11286,N_8266,N_5414);
and U11287 (N_11287,N_6274,N_5933);
nor U11288 (N_11288,N_9419,N_7105);
and U11289 (N_11289,N_6676,N_9765);
nand U11290 (N_11290,N_9131,N_5673);
or U11291 (N_11291,N_7334,N_6513);
and U11292 (N_11292,N_8194,N_5930);
xor U11293 (N_11293,N_5858,N_9234);
nor U11294 (N_11294,N_9564,N_8114);
xnor U11295 (N_11295,N_6556,N_6258);
nor U11296 (N_11296,N_6016,N_9088);
nand U11297 (N_11297,N_8759,N_9445);
xnor U11298 (N_11298,N_6714,N_6705);
and U11299 (N_11299,N_7355,N_6248);
nor U11300 (N_11300,N_7206,N_5418);
or U11301 (N_11301,N_6990,N_9876);
nor U11302 (N_11302,N_7896,N_6093);
nor U11303 (N_11303,N_8128,N_5734);
or U11304 (N_11304,N_9213,N_5914);
nor U11305 (N_11305,N_8012,N_9763);
and U11306 (N_11306,N_6698,N_5758);
or U11307 (N_11307,N_9384,N_5440);
nor U11308 (N_11308,N_9170,N_8000);
and U11309 (N_11309,N_9768,N_8950);
and U11310 (N_11310,N_6476,N_6142);
nor U11311 (N_11311,N_8807,N_9141);
xor U11312 (N_11312,N_9734,N_8903);
or U11313 (N_11313,N_9927,N_7731);
nand U11314 (N_11314,N_9277,N_8618);
xor U11315 (N_11315,N_8460,N_7039);
and U11316 (N_11316,N_6460,N_8043);
or U11317 (N_11317,N_6636,N_8145);
and U11318 (N_11318,N_9960,N_6206);
nand U11319 (N_11319,N_7976,N_6036);
nand U11320 (N_11320,N_9794,N_6495);
nand U11321 (N_11321,N_6875,N_5419);
and U11322 (N_11322,N_8944,N_6363);
and U11323 (N_11323,N_6433,N_8489);
or U11324 (N_11324,N_6640,N_7935);
or U11325 (N_11325,N_6731,N_9463);
nand U11326 (N_11326,N_7207,N_7672);
nand U11327 (N_11327,N_6885,N_5320);
or U11328 (N_11328,N_9725,N_7985);
nand U11329 (N_11329,N_9879,N_6107);
nor U11330 (N_11330,N_9918,N_7923);
nor U11331 (N_11331,N_6447,N_7389);
nand U11332 (N_11332,N_7486,N_9209);
or U11333 (N_11333,N_6896,N_5011);
xnor U11334 (N_11334,N_8548,N_6555);
nor U11335 (N_11335,N_9628,N_5239);
and U11336 (N_11336,N_7082,N_6315);
nor U11337 (N_11337,N_5486,N_6131);
or U11338 (N_11338,N_6237,N_8477);
or U11339 (N_11339,N_9481,N_5374);
xnor U11340 (N_11340,N_7598,N_8191);
and U11341 (N_11341,N_8447,N_8859);
nand U11342 (N_11342,N_6136,N_8654);
nand U11343 (N_11343,N_7508,N_8777);
xor U11344 (N_11344,N_6396,N_7198);
and U11345 (N_11345,N_9661,N_8666);
nand U11346 (N_11346,N_6891,N_7428);
xor U11347 (N_11347,N_5060,N_5348);
or U11348 (N_11348,N_5984,N_6652);
nor U11349 (N_11349,N_8709,N_5976);
and U11350 (N_11350,N_6688,N_9102);
or U11351 (N_11351,N_8396,N_6553);
nand U11352 (N_11352,N_5950,N_8131);
nor U11353 (N_11353,N_7245,N_7798);
nor U11354 (N_11354,N_9143,N_5243);
nand U11355 (N_11355,N_5229,N_9807);
xor U11356 (N_11356,N_6770,N_7572);
nand U11357 (N_11357,N_9664,N_7622);
or U11358 (N_11358,N_7698,N_9455);
nor U11359 (N_11359,N_7900,N_5257);
and U11360 (N_11360,N_8633,N_7399);
nand U11361 (N_11361,N_8369,N_5267);
nor U11362 (N_11362,N_5156,N_5290);
xnor U11363 (N_11363,N_6022,N_8855);
nand U11364 (N_11364,N_6525,N_9078);
nand U11365 (N_11365,N_7340,N_7898);
or U11366 (N_11366,N_7410,N_7496);
and U11367 (N_11367,N_7079,N_7757);
or U11368 (N_11368,N_8153,N_8360);
nand U11369 (N_11369,N_5602,N_7801);
xnor U11370 (N_11370,N_5501,N_8761);
xnor U11371 (N_11371,N_9622,N_9611);
and U11372 (N_11372,N_7473,N_9204);
nor U11373 (N_11373,N_5236,N_6953);
xor U11374 (N_11374,N_8742,N_6848);
xnor U11375 (N_11375,N_7870,N_5638);
xor U11376 (N_11376,N_9733,N_5055);
and U11377 (N_11377,N_7912,N_8103);
xnor U11378 (N_11378,N_8077,N_5570);
and U11379 (N_11379,N_7223,N_5795);
and U11380 (N_11380,N_5708,N_8748);
and U11381 (N_11381,N_6552,N_7849);
xnor U11382 (N_11382,N_8302,N_7619);
nor U11383 (N_11383,N_7229,N_9925);
or U11384 (N_11384,N_5317,N_6723);
xnor U11385 (N_11385,N_9963,N_9660);
nand U11386 (N_11386,N_7263,N_5014);
and U11387 (N_11387,N_7094,N_7134);
nor U11388 (N_11388,N_9696,N_6313);
xnor U11389 (N_11389,N_9649,N_7190);
and U11390 (N_11390,N_7316,N_7909);
or U11391 (N_11391,N_9862,N_8509);
nor U11392 (N_11392,N_7466,N_6995);
or U11393 (N_11393,N_8817,N_8386);
or U11394 (N_11394,N_8850,N_9467);
nand U11395 (N_11395,N_7290,N_6380);
xor U11396 (N_11396,N_6395,N_8827);
or U11397 (N_11397,N_7561,N_9535);
nand U11398 (N_11398,N_5591,N_6646);
xnor U11399 (N_11399,N_8074,N_8651);
nand U11400 (N_11400,N_6607,N_8758);
and U11401 (N_11401,N_6253,N_8583);
nor U11402 (N_11402,N_8126,N_7955);
and U11403 (N_11403,N_9563,N_5626);
or U11404 (N_11404,N_8754,N_7720);
or U11405 (N_11405,N_6674,N_5381);
nor U11406 (N_11406,N_9250,N_7356);
nand U11407 (N_11407,N_5286,N_8014);
or U11408 (N_11408,N_7233,N_5715);
nor U11409 (N_11409,N_8732,N_5588);
nor U11410 (N_11410,N_9305,N_8744);
and U11411 (N_11411,N_7398,N_6594);
nand U11412 (N_11412,N_7444,N_5071);
nor U11413 (N_11413,N_7135,N_8409);
xnor U11414 (N_11414,N_7778,N_9797);
nor U11415 (N_11415,N_8257,N_8600);
xor U11416 (N_11416,N_7425,N_6897);
xor U11417 (N_11417,N_9865,N_9376);
nor U11418 (N_11418,N_6767,N_5931);
nand U11419 (N_11419,N_9608,N_9990);
nor U11420 (N_11420,N_5304,N_9320);
and U11421 (N_11421,N_6887,N_6528);
xnor U11422 (N_11422,N_6610,N_5395);
nand U11423 (N_11423,N_9782,N_6333);
nor U11424 (N_11424,N_9254,N_5334);
nor U11425 (N_11425,N_5815,N_7493);
nand U11426 (N_11426,N_7630,N_7381);
and U11427 (N_11427,N_5133,N_7144);
xor U11428 (N_11428,N_8390,N_6511);
xnor U11429 (N_11429,N_9962,N_8494);
xor U11430 (N_11430,N_9387,N_7665);
nor U11431 (N_11431,N_9978,N_5903);
and U11432 (N_11432,N_7916,N_6557);
and U11433 (N_11433,N_9581,N_5937);
nand U11434 (N_11434,N_7300,N_8307);
nor U11435 (N_11435,N_8925,N_9877);
and U11436 (N_11436,N_9484,N_7752);
nor U11437 (N_11437,N_8141,N_8506);
nor U11438 (N_11438,N_5273,N_8857);
and U11439 (N_11439,N_7350,N_6808);
xnor U11440 (N_11440,N_5792,N_6242);
or U11441 (N_11441,N_5640,N_6792);
xnor U11442 (N_11442,N_9534,N_6465);
nor U11443 (N_11443,N_7744,N_9890);
nand U11444 (N_11444,N_8613,N_8882);
xor U11445 (N_11445,N_9032,N_6821);
or U11446 (N_11446,N_8280,N_9617);
nand U11447 (N_11447,N_6444,N_7587);
or U11448 (N_11448,N_7980,N_8567);
or U11449 (N_11449,N_5397,N_6507);
or U11450 (N_11450,N_7089,N_9002);
or U11451 (N_11451,N_9128,N_5850);
or U11452 (N_11452,N_5214,N_7511);
nor U11453 (N_11453,N_8730,N_5053);
nand U11454 (N_11454,N_6239,N_6729);
and U11455 (N_11455,N_5513,N_8786);
and U11456 (N_11456,N_8862,N_7974);
nor U11457 (N_11457,N_9348,N_9293);
nand U11458 (N_11458,N_9593,N_8318);
nand U11459 (N_11459,N_9085,N_9702);
or U11460 (N_11460,N_7066,N_6173);
nand U11461 (N_11461,N_8140,N_9997);
nor U11462 (N_11462,N_9756,N_8125);
xor U11463 (N_11463,N_9108,N_5113);
nand U11464 (N_11464,N_6404,N_9583);
or U11465 (N_11465,N_8860,N_8483);
and U11466 (N_11466,N_5332,N_9568);
xnor U11467 (N_11467,N_7999,N_7518);
nand U11468 (N_11468,N_9616,N_7845);
nand U11469 (N_11469,N_5605,N_8792);
xnor U11470 (N_11470,N_5598,N_6003);
xor U11471 (N_11471,N_9745,N_8990);
xor U11472 (N_11472,N_7950,N_6586);
and U11473 (N_11473,N_8522,N_7904);
nor U11474 (N_11474,N_7328,N_8804);
nor U11475 (N_11475,N_8213,N_7886);
and U11476 (N_11476,N_9916,N_5819);
or U11477 (N_11477,N_5278,N_5416);
and U11478 (N_11478,N_9380,N_7883);
nand U11479 (N_11479,N_6659,N_6466);
or U11480 (N_11480,N_8073,N_6072);
nand U11481 (N_11481,N_5003,N_5964);
nand U11482 (N_11482,N_5353,N_9774);
xor U11483 (N_11483,N_8229,N_7594);
nand U11484 (N_11484,N_5005,N_7621);
nand U11485 (N_11485,N_6842,N_9452);
xor U11486 (N_11486,N_5359,N_7202);
nor U11487 (N_11487,N_9911,N_6824);
xor U11488 (N_11488,N_5872,N_8602);
nor U11489 (N_11489,N_8928,N_7268);
xnor U11490 (N_11490,N_8072,N_5489);
nand U11491 (N_11491,N_9341,N_6174);
and U11492 (N_11492,N_8068,N_9208);
nor U11493 (N_11493,N_5847,N_8297);
xor U11494 (N_11494,N_9426,N_6470);
nor U11495 (N_11495,N_5037,N_8331);
or U11496 (N_11496,N_8940,N_9907);
nand U11497 (N_11497,N_6035,N_8977);
nand U11498 (N_11498,N_7449,N_9849);
or U11499 (N_11499,N_8904,N_7635);
xor U11500 (N_11500,N_5051,N_7346);
nand U11501 (N_11501,N_7411,N_5193);
nand U11502 (N_11502,N_5547,N_9961);
or U11503 (N_11503,N_9669,N_7994);
nand U11504 (N_11504,N_5845,N_5132);
xnor U11505 (N_11505,N_8584,N_7365);
nand U11506 (N_11506,N_6082,N_6158);
nand U11507 (N_11507,N_7979,N_9580);
nor U11508 (N_11508,N_8715,N_9448);
xnor U11509 (N_11509,N_8203,N_9772);
nand U11510 (N_11510,N_8031,N_9324);
xnor U11511 (N_11511,N_5794,N_9931);
nor U11512 (N_11512,N_9153,N_9827);
xnor U11513 (N_11513,N_7327,N_9749);
nor U11514 (N_11514,N_9587,N_9542);
and U11515 (N_11515,N_7899,N_5737);
nor U11516 (N_11516,N_7272,N_7864);
nand U11517 (N_11517,N_7254,N_8918);
nand U11518 (N_11518,N_6689,N_9908);
nand U11519 (N_11519,N_5176,N_8018);
and U11520 (N_11520,N_6680,N_5431);
xnor U11521 (N_11521,N_7335,N_8581);
and U11522 (N_11522,N_7646,N_8470);
nor U11523 (N_11523,N_6303,N_7709);
or U11524 (N_11524,N_5973,N_6024);
and U11525 (N_11525,N_9061,N_8458);
or U11526 (N_11526,N_7276,N_5508);
nand U11527 (N_11527,N_8002,N_5596);
or U11528 (N_11528,N_9923,N_8652);
or U11529 (N_11529,N_9715,N_5574);
xnor U11530 (N_11530,N_9900,N_6306);
xnor U11531 (N_11531,N_8557,N_7182);
nor U11532 (N_11532,N_8109,N_7185);
nor U11533 (N_11533,N_7441,N_9025);
or U11534 (N_11534,N_6718,N_8891);
nand U11535 (N_11535,N_6893,N_8372);
nand U11536 (N_11536,N_9965,N_7257);
nand U11537 (N_11537,N_6104,N_5522);
nand U11538 (N_11538,N_9712,N_9118);
nand U11539 (N_11539,N_7578,N_8848);
and U11540 (N_11540,N_6836,N_5145);
and U11541 (N_11541,N_8539,N_9922);
nand U11542 (N_11542,N_9227,N_8488);
nor U11543 (N_11543,N_7216,N_9422);
and U11544 (N_11544,N_6159,N_9107);
xnor U11545 (N_11545,N_8365,N_5342);
xnor U11546 (N_11546,N_7102,N_9682);
or U11547 (N_11547,N_6878,N_6882);
nand U11548 (N_11548,N_5701,N_9716);
and U11549 (N_11549,N_8121,N_7947);
nor U11550 (N_11550,N_8462,N_5505);
xor U11551 (N_11551,N_6241,N_7517);
xnor U11552 (N_11552,N_5115,N_5647);
xnor U11553 (N_11553,N_9781,N_6779);
xnor U11554 (N_11554,N_6259,N_5975);
nor U11555 (N_11555,N_6643,N_9895);
nand U11556 (N_11556,N_7867,N_7456);
nor U11557 (N_11557,N_6027,N_6000);
and U11558 (N_11558,N_7876,N_8394);
and U11559 (N_11559,N_9838,N_6859);
nand U11560 (N_11560,N_9198,N_7324);
xnor U11561 (N_11561,N_7803,N_8683);
or U11562 (N_11562,N_8252,N_9612);
nand U11563 (N_11563,N_6175,N_8835);
or U11564 (N_11564,N_5335,N_8220);
nor U11565 (N_11565,N_9676,N_8853);
nor U11566 (N_11566,N_8974,N_6269);
and U11567 (N_11567,N_6713,N_6667);
nor U11568 (N_11568,N_5246,N_5240);
or U11569 (N_11569,N_8660,N_5349);
or U11570 (N_11570,N_6857,N_5702);
or U11571 (N_11571,N_6077,N_8452);
or U11572 (N_11572,N_8576,N_5283);
or U11573 (N_11573,N_9266,N_9075);
and U11574 (N_11574,N_5796,N_6706);
xor U11575 (N_11575,N_7230,N_9808);
and U11576 (N_11576,N_5080,N_7737);
or U11577 (N_11577,N_9390,N_7627);
or U11578 (N_11578,N_6829,N_9185);
nand U11579 (N_11579,N_6078,N_9047);
nand U11580 (N_11580,N_5025,N_9995);
and U11581 (N_11581,N_5785,N_8044);
nand U11582 (N_11582,N_5960,N_5627);
nor U11583 (N_11583,N_9414,N_5120);
xnor U11584 (N_11584,N_8690,N_7434);
and U11585 (N_11585,N_5873,N_6707);
nand U11586 (N_11586,N_7595,N_6040);
and U11587 (N_11587,N_6919,N_5232);
and U11588 (N_11588,N_7303,N_6628);
xnor U11589 (N_11589,N_9692,N_6489);
and U11590 (N_11590,N_6458,N_6178);
or U11591 (N_11591,N_6160,N_8081);
or U11592 (N_11592,N_5546,N_9155);
xor U11593 (N_11593,N_6448,N_6240);
and U11594 (N_11594,N_9884,N_7712);
nor U11595 (N_11595,N_8755,N_5247);
nand U11596 (N_11596,N_9095,N_5167);
nor U11597 (N_11597,N_6546,N_7550);
and U11598 (N_11598,N_6733,N_8717);
nand U11599 (N_11599,N_8473,N_6186);
nor U11600 (N_11600,N_5997,N_6029);
or U11601 (N_11601,N_8623,N_8024);
or U11602 (N_11602,N_6580,N_6616);
xnor U11603 (N_11603,N_7585,N_7580);
and U11604 (N_11604,N_6094,N_9561);
xnor U11605 (N_11605,N_8627,N_9885);
and U11606 (N_11606,N_6057,N_5560);
and U11607 (N_11607,N_7313,N_5962);
xor U11608 (N_11608,N_5705,N_5221);
and U11609 (N_11609,N_5265,N_9543);
nor U11610 (N_11610,N_6018,N_5478);
xnor U11611 (N_11611,N_9127,N_5532);
nor U11612 (N_11612,N_5062,N_8673);
xor U11613 (N_11613,N_7298,N_6459);
or U11614 (N_11614,N_9362,N_7413);
nand U11615 (N_11615,N_9560,N_7861);
xor U11616 (N_11616,N_6080,N_8800);
and U11617 (N_11617,N_8685,N_9536);
nor U11618 (N_11618,N_7860,N_7675);
and U11619 (N_11619,N_7796,N_9424);
or U11620 (N_11620,N_9764,N_6796);
nand U11621 (N_11621,N_9946,N_8010);
xnor U11622 (N_11622,N_8669,N_9114);
or U11623 (N_11623,N_8953,N_8373);
xor U11624 (N_11624,N_8644,N_7034);
and U11625 (N_11625,N_8514,N_8689);
xor U11626 (N_11626,N_7958,N_6378);
xor U11627 (N_11627,N_8305,N_8100);
nor U11628 (N_11628,N_9857,N_5524);
or U11629 (N_11629,N_6468,N_6455);
nor U11630 (N_11630,N_9630,N_6613);
nand U11631 (N_11631,N_6230,N_8803);
xnor U11632 (N_11632,N_6917,N_7548);
nand U11633 (N_11633,N_8299,N_7760);
or U11634 (N_11634,N_8466,N_8889);
and U11635 (N_11635,N_6445,N_5001);
and U11636 (N_11636,N_7875,N_6931);
and U11637 (N_11637,N_9146,N_7419);
or U11638 (N_11638,N_8110,N_8422);
and U11639 (N_11639,N_8319,N_6630);
and U11640 (N_11640,N_7406,N_6400);
xnor U11641 (N_11641,N_7588,N_5549);
and U11642 (N_11642,N_9386,N_6576);
or U11643 (N_11643,N_5388,N_5048);
nand U11644 (N_11644,N_8361,N_8382);
xnor U11645 (N_11645,N_6692,N_5380);
or U11646 (N_11646,N_8869,N_8223);
xor U11647 (N_11647,N_8638,N_6855);
or U11648 (N_11648,N_8604,N_9975);
nand U11649 (N_11649,N_6997,N_5297);
nand U11650 (N_11650,N_5924,N_5084);
or U11651 (N_11651,N_9964,N_7248);
nand U11652 (N_11652,N_9529,N_5015);
nor U11653 (N_11653,N_9944,N_8334);
xor U11654 (N_11654,N_5915,N_6179);
and U11655 (N_11655,N_8668,N_5024);
xor U11656 (N_11656,N_8662,N_7489);
nor U11657 (N_11657,N_7687,N_9226);
xor U11658 (N_11658,N_8005,N_7543);
and U11659 (N_11659,N_7430,N_7440);
nor U11660 (N_11660,N_8217,N_8603);
nand U11661 (N_11661,N_7717,N_9041);
and U11662 (N_11662,N_8041,N_7931);
or U11663 (N_11663,N_9262,N_9710);
nor U11664 (N_11664,N_7152,N_8505);
nand U11665 (N_11665,N_9276,N_5745);
nor U11666 (N_11666,N_5918,N_5066);
xor U11667 (N_11667,N_7457,N_8042);
or U11668 (N_11668,N_8912,N_5632);
or U11669 (N_11669,N_5255,N_5200);
nand U11670 (N_11670,N_8809,N_6183);
xnor U11671 (N_11671,N_5691,N_6105);
or U11672 (N_11672,N_8272,N_8663);
xnor U11673 (N_11673,N_8375,N_7748);
nand U11674 (N_11674,N_5065,N_7986);
nor U11675 (N_11675,N_5023,N_6522);
and U11676 (N_11676,N_6120,N_6769);
nand U11677 (N_11677,N_9639,N_5308);
and U11678 (N_11678,N_7452,N_6211);
xor U11679 (N_11679,N_5742,N_6058);
or U11680 (N_11680,N_8197,N_8258);
nor U11681 (N_11681,N_9343,N_7351);
xnor U11682 (N_11682,N_7940,N_7225);
nor U11683 (N_11683,N_6290,N_8722);
nor U11684 (N_11684,N_7837,N_9389);
xor U11685 (N_11685,N_8146,N_5373);
xnor U11686 (N_11686,N_9158,N_8607);
nand U11687 (N_11687,N_8502,N_9754);
or U11688 (N_11688,N_6890,N_7041);
xnor U11689 (N_11689,N_6536,N_7247);
nor U11690 (N_11690,N_9576,N_5220);
and U11691 (N_11691,N_9512,N_5601);
and U11692 (N_11692,N_8712,N_9321);
nand U11693 (N_11693,N_8572,N_5166);
and U11694 (N_11694,N_8330,N_9010);
nand U11695 (N_11695,N_9493,N_6314);
nor U11696 (N_11696,N_8468,N_5344);
xnor U11697 (N_11697,N_5125,N_7975);
nor U11698 (N_11698,N_6039,N_8877);
xnor U11699 (N_11699,N_8227,N_5558);
nand U11700 (N_11700,N_7278,N_5902);
or U11701 (N_11701,N_9203,N_8405);
and U11702 (N_11702,N_8836,N_5657);
nand U11703 (N_11703,N_6499,N_9641);
and U11704 (N_11704,N_6231,N_8237);
nand U11705 (N_11705,N_8789,N_7366);
and U11706 (N_11706,N_8778,N_7421);
xor U11707 (N_11707,N_8762,N_9601);
nand U11708 (N_11708,N_5404,N_7780);
or U11709 (N_11709,N_6001,N_8880);
and U11710 (N_11710,N_8776,N_9558);
and U11711 (N_11711,N_8787,N_9823);
nor U11712 (N_11712,N_9432,N_9205);
nor U11713 (N_11713,N_8413,N_5068);
nand U11714 (N_11714,N_7753,N_7277);
xnor U11715 (N_11715,N_5661,N_8269);
xor U11716 (N_11716,N_9133,N_9670);
xnor U11717 (N_11717,N_9156,N_6874);
nor U11718 (N_11718,N_5528,N_8023);
xor U11719 (N_11719,N_9403,N_5707);
or U11720 (N_11720,N_5822,N_7266);
xor U11721 (N_11721,N_9400,N_5266);
nand U11722 (N_11722,N_9572,N_7169);
xnor U11723 (N_11723,N_7581,N_7684);
nand U11724 (N_11724,N_8417,N_5180);
and U11725 (N_11725,N_5531,N_5085);
nand U11726 (N_11726,N_7997,N_5046);
or U11727 (N_11727,N_9479,N_7487);
xor U11728 (N_11728,N_8558,N_6083);
xnor U11729 (N_11729,N_6625,N_6532);
nor U11730 (N_11730,N_6318,N_9206);
and U11731 (N_11731,N_7161,N_5331);
or U11732 (N_11732,N_7629,N_8219);
nor U11733 (N_11733,N_8313,N_9870);
nand U11734 (N_11734,N_9037,N_9471);
nor U11735 (N_11735,N_6545,N_5967);
nand U11736 (N_11736,N_7078,N_5782);
nor U11737 (N_11737,N_9473,N_7363);
nand U11738 (N_11738,N_7155,N_8106);
nand U11739 (N_11739,N_7283,N_9549);
nor U11740 (N_11740,N_5799,N_8681);
or U11741 (N_11741,N_9627,N_6140);
nor U11742 (N_11742,N_5697,N_9686);
nand U11743 (N_11743,N_9288,N_5736);
nand U11744 (N_11744,N_8270,N_8058);
nor U11745 (N_11745,N_9632,N_9897);
and U11746 (N_11746,N_5463,N_9915);
nor U11747 (N_11747,N_5248,N_5709);
xnor U11748 (N_11748,N_8457,N_7671);
nor U11749 (N_11749,N_9841,N_5630);
and U11750 (N_11750,N_5171,N_7832);
nand U11751 (N_11751,N_9721,N_5889);
or U11752 (N_11752,N_6588,N_9556);
xnor U11753 (N_11753,N_7453,N_9326);
or U11754 (N_11754,N_6768,N_9839);
or U11755 (N_11755,N_5251,N_9514);
xnor U11756 (N_11756,N_7241,N_8875);
and U11757 (N_11757,N_6212,N_9058);
and U11758 (N_11758,N_7763,N_7117);
nor U11759 (N_11759,N_6802,N_6691);
and U11760 (N_11760,N_9096,N_8151);
and U11761 (N_11761,N_7963,N_7018);
xor U11762 (N_11762,N_6967,N_7502);
and U11763 (N_11763,N_6286,N_8332);
or U11764 (N_11764,N_5557,N_5010);
nor U11765 (N_11765,N_7809,N_8615);
nor U11766 (N_11766,N_5738,N_8629);
xnor U11767 (N_11767,N_8865,N_5741);
xor U11768 (N_11768,N_7841,N_7132);
or U11769 (N_11769,N_5866,N_6877);
and U11770 (N_11770,N_7423,N_9510);
or U11771 (N_11771,N_9212,N_9031);
nand U11772 (N_11772,N_6783,N_8749);
nand U11773 (N_11773,N_7353,N_6589);
xor U11774 (N_11774,N_7636,N_8626);
or U11775 (N_11775,N_8064,N_8963);
xor U11776 (N_11776,N_6841,N_8565);
nand U11777 (N_11777,N_7137,N_6579);
and U11778 (N_11778,N_5347,N_9845);
and U11779 (N_11779,N_6092,N_7221);
nor U11780 (N_11780,N_8687,N_5195);
and U11781 (N_11781,N_9200,N_7345);
xnor U11782 (N_11782,N_6551,N_7887);
nor U11783 (N_11783,N_5523,N_6352);
and U11784 (N_11784,N_8736,N_7738);
or U11785 (N_11785,N_6134,N_6921);
xnor U11786 (N_11786,N_8118,N_8314);
nor U11787 (N_11787,N_7730,N_9003);
and U11788 (N_11788,N_9265,N_5910);
or U11789 (N_11789,N_7674,N_5980);
xnor U11790 (N_11790,N_5728,N_6904);
and U11791 (N_11791,N_7302,N_5107);
nand U11792 (N_11792,N_9930,N_7888);
and U11793 (N_11793,N_9103,N_9218);
or U11794 (N_11794,N_9974,N_9784);
and U11795 (N_11795,N_7930,N_9357);
xnor U11796 (N_11796,N_6432,N_5042);
xnor U11797 (N_11797,N_5087,N_6198);
nand U11798 (N_11798,N_9328,N_5022);
xor U11799 (N_11799,N_7168,N_9021);
xor U11800 (N_11800,N_9971,N_8781);
and U11801 (N_11801,N_6809,N_7088);
xnor U11802 (N_11802,N_5864,N_7941);
nand U11803 (N_11803,N_9311,N_9270);
and U11804 (N_11804,N_8612,N_6818);
nand U11805 (N_11805,N_6337,N_5721);
nand U11806 (N_11806,N_6073,N_6851);
nand U11807 (N_11807,N_9485,N_6852);
or U11808 (N_11808,N_8799,N_7812);
nor U11809 (N_11809,N_7331,N_6436);
xnor U11810 (N_11810,N_5234,N_6865);
xor U11811 (N_11811,N_6884,N_8345);
xor U11812 (N_11812,N_7418,N_5840);
or U11813 (N_11813,N_5456,N_8403);
and U11814 (N_11814,N_8152,N_5086);
and U11815 (N_11815,N_6654,N_9026);
and U11816 (N_11816,N_5559,N_7677);
and U11817 (N_11817,N_9596,N_6810);
nand U11818 (N_11818,N_7814,N_9981);
nand U11819 (N_11819,N_7326,N_7236);
xor U11820 (N_11820,N_8107,N_8343);
xnor U11821 (N_11821,N_8322,N_7725);
nand U11822 (N_11822,N_5952,N_7030);
or U11823 (N_11823,N_7807,N_8774);
or U11824 (N_11824,N_7321,N_9521);
and U11825 (N_11825,N_6907,N_8292);
xnor U11826 (N_11826,N_6955,N_6598);
xor U11827 (N_11827,N_5009,N_6117);
or U11828 (N_11828,N_5153,N_8428);
and U11829 (N_11829,N_8580,N_6124);
or U11830 (N_11830,N_7791,N_7173);
nor U11831 (N_11831,N_5219,N_9183);
or U11832 (N_11832,N_7680,N_8711);
nand U11833 (N_11833,N_7783,N_6781);
nor U11834 (N_11834,N_6780,N_5249);
nor U11835 (N_11835,N_7568,N_5361);
and U11836 (N_11836,N_7433,N_6992);
nand U11837 (N_11837,N_8766,N_6343);
or U11838 (N_11838,N_6184,N_5943);
or U11839 (N_11839,N_8590,N_9831);
nor U11840 (N_11840,N_9906,N_9634);
and U11841 (N_11841,N_7322,N_6510);
or U11842 (N_11842,N_7342,N_7524);
and U11843 (N_11843,N_7501,N_8765);
xor U11844 (N_11844,N_7911,N_9433);
or U11845 (N_11845,N_7217,N_8772);
xnor U11846 (N_11846,N_7792,N_9444);
nand U11847 (N_11847,N_7491,N_8157);
nand U11848 (N_11848,N_8022,N_6161);
and U11849 (N_11849,N_5458,N_6568);
nor U11850 (N_11850,N_5224,N_9864);
and U11851 (N_11851,N_7639,N_5826);
or U11852 (N_11852,N_5816,N_5477);
nand U11853 (N_11853,N_7373,N_5198);
nand U11854 (N_11854,N_6750,N_5276);
and U11855 (N_11855,N_8087,N_7831);
nor U11856 (N_11856,N_9015,N_6828);
and U11857 (N_11857,N_5441,N_8970);
nand U11858 (N_11858,N_9066,N_6609);
nand U11859 (N_11859,N_7767,N_8055);
nor U11860 (N_11860,N_8531,N_5235);
or U11861 (N_11861,N_8958,N_7742);
and U11862 (N_11862,N_6736,N_8366);
xnor U11863 (N_11863,N_9769,N_9487);
or U11864 (N_11864,N_8115,N_8328);
nand U11865 (N_11865,N_9215,N_9217);
nand U11866 (N_11866,N_8123,N_9309);
xor U11867 (N_11867,N_7574,N_8434);
nor U11868 (N_11868,N_6126,N_8815);
nor U11869 (N_11869,N_9517,N_8337);
or U11870 (N_11870,N_5294,N_9117);
or U11871 (N_11871,N_7987,N_8794);
and U11872 (N_11872,N_5911,N_5215);
or U11873 (N_11873,N_8367,N_6900);
and U11874 (N_11874,N_6732,N_8200);
nand U11875 (N_11875,N_7924,N_6973);
and U11876 (N_11876,N_6254,N_6533);
xor U11877 (N_11877,N_6325,N_9956);
nor U11878 (N_11878,N_6413,N_6864);
or U11879 (N_11879,N_7296,N_8743);
xnor U11880 (N_11880,N_9887,N_5254);
nor U11881 (N_11881,N_7026,N_9024);
nand U11882 (N_11882,N_8207,N_6087);
and U11883 (N_11883,N_8964,N_5484);
xor U11884 (N_11884,N_5260,N_9478);
and U11885 (N_11885,N_6663,N_5245);
or U11886 (N_11886,N_5494,N_7648);
and U11887 (N_11887,N_8790,N_8930);
nand U11888 (N_11888,N_9344,N_5763);
nand U11889 (N_11889,N_8161,N_6234);
xor U11890 (N_11890,N_6457,N_9790);
nand U11891 (N_11891,N_9779,N_8921);
nor U11892 (N_11892,N_8174,N_6946);
nand U11893 (N_11893,N_6030,N_5832);
nand U11894 (N_11894,N_6710,N_6168);
nand U11895 (N_11895,N_6649,N_9852);
nand U11896 (N_11896,N_6991,N_5128);
xnor U11897 (N_11897,N_8589,N_5706);
xor U11898 (N_11898,N_5044,N_9637);
nand U11899 (N_11899,N_7181,N_6746);
nand U11900 (N_11900,N_5690,N_8655);
and U11901 (N_11901,N_8206,N_7231);
and U11902 (N_11902,N_6581,N_6949);
nand U11903 (N_11903,N_9291,N_6599);
nand U11904 (N_11904,N_9191,N_9147);
and U11905 (N_11905,N_7474,N_8124);
and U11906 (N_11906,N_6228,N_7465);
or U11907 (N_11907,N_5116,N_5453);
xor U11908 (N_11908,N_9079,N_8907);
xnor U11909 (N_11909,N_7768,N_9100);
nand U11910 (N_11910,N_5805,N_9437);
xnor U11911 (N_11911,N_5534,N_6215);
nor U11912 (N_11912,N_5429,N_5886);
nand U11913 (N_11913,N_6839,N_8994);
or U11914 (N_11914,N_6452,N_9115);
nor U11915 (N_11915,N_9246,N_8271);
and U11916 (N_11916,N_8176,N_6975);
or U11917 (N_11917,N_8347,N_5427);
and U11918 (N_11918,N_9458,N_8095);
nor U11919 (N_11919,N_9780,N_5242);
and U11920 (N_11920,N_8093,N_8527);
nor U11921 (N_11921,N_7482,N_8402);
xnor U11922 (N_11922,N_8746,N_8802);
or U11923 (N_11923,N_5036,N_5399);
nand U11924 (N_11924,N_5169,N_7081);
and U11925 (N_11925,N_7692,N_9411);
or U11926 (N_11926,N_5096,N_5299);
nand U11927 (N_11927,N_9714,N_6873);
or U11928 (N_11928,N_6562,N_8441);
or U11929 (N_11929,N_9408,N_5798);
nor U11930 (N_11930,N_5938,N_8130);
or U11931 (N_11931,N_5330,N_9179);
xnor U11932 (N_11932,N_5343,N_5464);
and U11933 (N_11933,N_7794,N_7854);
and U11934 (N_11934,N_6133,N_7644);
or U11935 (N_11935,N_7361,N_9435);
xnor U11936 (N_11936,N_5841,N_7120);
nand U11937 (N_11937,N_8649,N_6348);
and U11938 (N_11938,N_8876,N_8242);
nor U11939 (N_11939,N_7566,N_7011);
or U11940 (N_11940,N_5114,N_5274);
and U11941 (N_11941,N_6968,N_8890);
or U11942 (N_11942,N_7255,N_8549);
nand U11943 (N_11943,N_5584,N_9667);
xor U11944 (N_11944,N_7252,N_5007);
nor U11945 (N_11945,N_5987,N_9585);
nand U11946 (N_11946,N_9011,N_9072);
or U11947 (N_11947,N_7681,N_5564);
or U11948 (N_11948,N_9695,N_7214);
nand U11949 (N_11949,N_8599,N_7685);
and U11950 (N_11950,N_5175,N_9938);
xor U11951 (N_11951,N_5957,N_8233);
or U11952 (N_11952,N_9984,N_9486);
nand U11953 (N_11953,N_6539,N_8908);
nor U11954 (N_11954,N_8861,N_8478);
or U11955 (N_11955,N_6170,N_7317);
nand U11956 (N_11956,N_8201,N_7141);
nand U11957 (N_11957,N_8818,N_8825);
xnor U11958 (N_11958,N_9739,N_6238);
and U11959 (N_11959,N_5306,N_8459);
nand U11960 (N_11960,N_9554,N_7101);
xor U11961 (N_11961,N_6756,N_8585);
xnor U11962 (N_11962,N_7835,N_6549);
nand U11963 (N_11963,N_5357,N_7193);
nor U11964 (N_11964,N_8596,N_5336);
nand U11965 (N_11965,N_6129,N_5854);
or U11966 (N_11966,N_9582,N_9406);
nor U11967 (N_11967,N_6138,N_9957);
nand U11968 (N_11968,N_7830,N_5636);
xnor U11969 (N_11969,N_8739,N_6696);
or U11970 (N_11970,N_5568,N_9057);
nand U11971 (N_11971,N_9347,N_6102);
nor U11972 (N_11972,N_7821,N_9239);
nor U11973 (N_11973,N_8454,N_7377);
nor U11974 (N_11974,N_9602,N_7320);
or U11975 (N_11975,N_9869,N_5061);
and U11976 (N_11976,N_5095,N_6721);
nor U11977 (N_11977,N_5078,N_8701);
nor U11978 (N_11978,N_8033,N_9171);
or U11979 (N_11979,N_9190,N_5780);
nand U11980 (N_11980,N_9497,N_8071);
xor U11981 (N_11981,N_6116,N_6069);
nor U11982 (N_11982,N_8814,N_7370);
xor U11983 (N_11983,N_9762,N_9263);
or U11984 (N_11984,N_9214,N_9009);
nor U11985 (N_11985,N_6742,N_6403);
nor U11986 (N_11986,N_9358,N_7250);
xor U11987 (N_11987,N_9524,N_9503);
or U11988 (N_11988,N_8240,N_7567);
and U11989 (N_11989,N_9924,N_7873);
nand U11990 (N_11990,N_8959,N_6765);
xor U11991 (N_11991,N_7758,N_5869);
nor U11992 (N_11992,N_8508,N_9221);
or U11993 (N_11993,N_5665,N_6300);
or U11994 (N_11994,N_7560,N_9407);
nor U11995 (N_11995,N_5565,N_6213);
nand U11996 (N_11996,N_9236,N_9315);
or U11997 (N_11997,N_9469,N_9381);
xor U11998 (N_11998,N_7151,N_9207);
nor U11999 (N_11999,N_6332,N_9750);
or U12000 (N_12000,N_8998,N_9787);
or U12001 (N_12001,N_8255,N_9594);
or U12002 (N_12002,N_8383,N_6125);
xnor U12003 (N_12003,N_7315,N_7055);
nor U12004 (N_12004,N_6784,N_6856);
nand U12005 (N_12005,N_9157,N_8149);
or U12006 (N_12006,N_9783,N_5423);
or U12007 (N_12007,N_5995,N_9295);
xor U12008 (N_12008,N_5996,N_6664);
and U12009 (N_12009,N_5385,N_6053);
and U12010 (N_12010,N_8425,N_5218);
nand U12011 (N_12011,N_8119,N_9854);
nand U12012 (N_12012,N_7019,N_7093);
and U12013 (N_12013,N_7765,N_7118);
and U12014 (N_12014,N_6066,N_5882);
and U12015 (N_12015,N_9809,N_8052);
and U12016 (N_12016,N_6197,N_5415);
nor U12017 (N_12017,N_6785,N_5571);
nand U12018 (N_12018,N_6045,N_9030);
xor U12019 (N_12019,N_6850,N_6099);
and U12020 (N_12020,N_6049,N_9392);
or U12021 (N_12021,N_8915,N_8852);
xor U12022 (N_12022,N_5857,N_8538);
xor U12023 (N_12023,N_8516,N_9866);
nor U12024 (N_12024,N_6728,N_8670);
nor U12025 (N_12025,N_5615,N_8327);
and U12026 (N_12026,N_9886,N_6062);
nand U12027 (N_12027,N_6472,N_8443);
or U12028 (N_12028,N_5874,N_8507);
nor U12029 (N_12029,N_8588,N_7192);
and U12030 (N_12030,N_5301,N_6901);
nor U12031 (N_12031,N_6449,N_9926);
nand U12032 (N_12032,N_5140,N_6916);
xor U12033 (N_12033,N_5635,N_7492);
and U12034 (N_12034,N_5658,N_6858);
nor U12035 (N_12035,N_8485,N_8540);
nand U12036 (N_12036,N_8491,N_8268);
xor U12037 (N_12037,N_8205,N_5526);
or U12038 (N_12038,N_8932,N_5556);
and U12039 (N_12039,N_8962,N_6284);
and U12040 (N_12040,N_8430,N_5641);
and U12041 (N_12041,N_6205,N_8007);
or U12042 (N_12042,N_7357,N_6948);
nor U12043 (N_12043,N_8608,N_5725);
nand U12044 (N_12044,N_6944,N_9539);
nor U12045 (N_12045,N_9396,N_6020);
or U12046 (N_12046,N_9322,N_7816);
nand U12047 (N_12047,N_7509,N_8735);
nor U12048 (N_12048,N_5288,N_9074);
xor U12049 (N_12049,N_8653,N_7160);
xnor U12050 (N_12050,N_6307,N_8444);
or U12051 (N_12051,N_8631,N_7405);
or U12052 (N_12052,N_6119,N_5407);
or U12053 (N_12053,N_8515,N_5400);
xor U12054 (N_12054,N_9559,N_8648);
nor U12055 (N_12055,N_7589,N_7507);
and U12056 (N_12056,N_9029,N_5801);
nand U12057 (N_12057,N_5716,N_8851);
and U12058 (N_12058,N_6166,N_7762);
and U12059 (N_12059,N_7201,N_6427);
xor U12060 (N_12060,N_8978,N_9812);
nand U12061 (N_12061,N_9124,N_7281);
or U12062 (N_12062,N_6075,N_5459);
or U12063 (N_12063,N_5157,N_5356);
nand U12064 (N_12064,N_6270,N_5633);
and U12065 (N_12065,N_7077,N_5137);
or U12066 (N_12066,N_6517,N_5462);
or U12067 (N_12067,N_6439,N_9522);
nor U12068 (N_12068,N_5578,N_8051);
nand U12069 (N_12069,N_5408,N_9310);
and U12070 (N_12070,N_7826,N_6751);
or U12071 (N_12071,N_8303,N_8667);
nand U12072 (N_12072,N_7577,N_6381);
xor U12073 (N_12073,N_5341,N_9273);
or U12074 (N_12074,N_7795,N_9245);
nor U12075 (N_12075,N_5660,N_5448);
or U12076 (N_12076,N_7564,N_6650);
or U12077 (N_12077,N_9132,N_5935);
nor U12078 (N_12078,N_9820,N_7488);
or U12079 (N_12079,N_7178,N_5618);
nor U12080 (N_12080,N_5067,N_7779);
and U12081 (N_12081,N_5704,N_8961);
or U12082 (N_12082,N_7299,N_9735);
xor U12083 (N_12083,N_8432,N_8225);
nor U12084 (N_12084,N_6655,N_7605);
and U12085 (N_12085,N_7696,N_9253);
xnor U12086 (N_12086,N_6735,N_7628);
and U12087 (N_12087,N_7069,N_9154);
nor U12088 (N_12088,N_5020,N_7949);
or U12089 (N_12089,N_9999,N_8135);
or U12090 (N_12090,N_6819,N_7130);
or U12091 (N_12091,N_8285,N_9136);
or U12092 (N_12092,N_6558,N_9122);
xor U12093 (N_12093,N_8208,N_7076);
and U12094 (N_12094,N_5791,N_7084);
and U12095 (N_12095,N_6595,N_7637);
or U12096 (N_12096,N_8938,N_6994);
nor U12097 (N_12097,N_8351,N_7448);
xnor U12098 (N_12098,N_5040,N_8467);
or U12099 (N_12099,N_7354,N_9707);
and U12100 (N_12100,N_6763,N_8162);
and U12101 (N_12101,N_8017,N_5366);
or U12102 (N_12102,N_5384,N_5365);
and U12103 (N_12103,N_6276,N_9220);
xnor U12104 (N_12104,N_6753,N_5100);
nor U12105 (N_12105,N_9149,N_8993);
xnor U12106 (N_12106,N_9287,N_5031);
or U12107 (N_12107,N_9562,N_8750);
nand U12108 (N_12108,N_5755,N_9557);
and U12109 (N_12109,N_9648,N_6782);
and U12110 (N_12110,N_6287,N_9083);
nor U12111 (N_12111,N_5496,N_9004);
nand U12112 (N_12112,N_6559,N_6366);
and U12113 (N_12113,N_8844,N_8634);
nand U12114 (N_12114,N_5035,N_7336);
nand U12115 (N_12115,N_7163,N_8747);
or U12116 (N_12116,N_9832,N_6399);
nand U12117 (N_12117,N_6854,N_8672);
and U12118 (N_12118,N_7243,N_7590);
or U12119 (N_12119,N_6614,N_7961);
and U12120 (N_12120,N_6055,N_6501);
nand U12121 (N_12121,N_7604,N_9904);
or U12122 (N_12122,N_5111,N_6711);
nand U12123 (N_12123,N_5905,N_7109);
xor U12124 (N_12124,N_9551,N_7631);
or U12125 (N_12125,N_7475,N_7972);
or U12126 (N_12126,N_6801,N_7611);
or U12127 (N_12127,N_7046,N_8426);
and U12128 (N_12128,N_9223,N_6648);
and U12129 (N_12129,N_5940,N_6042);
or U12130 (N_12130,N_5075,N_8401);
xor U12131 (N_12131,N_8706,N_8569);
nor U12132 (N_12132,N_8291,N_8276);
and U12133 (N_12133,N_9798,N_9619);
or U12134 (N_12134,N_9933,N_8315);
nand U12135 (N_12135,N_5269,N_7549);
nor U12136 (N_12136,N_8296,N_6985);
nor U12137 (N_12137,N_5144,N_5577);
nand U12138 (N_12138,N_7396,N_7579);
nand U12139 (N_12139,N_5589,N_9164);
and U12140 (N_12140,N_9842,N_9027);
nand U12141 (N_12141,N_8391,N_6816);
or U12142 (N_12142,N_8534,N_5842);
and U12143 (N_12143,N_7643,N_9824);
nand U12144 (N_12144,N_7360,N_6656);
nand U12145 (N_12145,N_6759,N_6815);
nor U12146 (N_12146,N_8142,N_9038);
or U12147 (N_12147,N_8570,N_7996);
xnor U12148 (N_12148,N_7070,N_9919);
xor U12149 (N_12149,N_6703,N_7261);
or U12150 (N_12150,N_7530,N_8304);
xor U12151 (N_12151,N_8697,N_5130);
xnor U12152 (N_12152,N_6021,N_5291);
nor U12153 (N_12153,N_8960,N_5223);
nor U12154 (N_12154,N_8034,N_7280);
and U12155 (N_12155,N_6950,N_9453);
and U12156 (N_12156,N_9531,N_6247);
xnor U12157 (N_12157,N_9703,N_6367);
nand U12158 (N_12158,N_5944,N_8782);
or U12159 (N_12159,N_5779,N_7210);
nor U12160 (N_12160,N_7733,N_5863);
or U12161 (N_12161,N_7186,N_7862);
and U12162 (N_12162,N_5744,N_5442);
or U12163 (N_12163,N_9844,N_6697);
and U12164 (N_12164,N_9878,N_7314);
or U12165 (N_12165,N_6407,N_9036);
nand U12166 (N_12166,N_9065,N_9371);
nand U12167 (N_12167,N_5947,N_5851);
nor U12168 (N_12168,N_5862,N_7823);
or U12169 (N_12169,N_9732,N_8082);
or U12170 (N_12170,N_9033,N_6130);
nor U12171 (N_12171,N_9760,N_7108);
nand U12172 (N_12172,N_6966,N_9165);
nand U12173 (N_12173,N_8177,N_8137);
and U12174 (N_12174,N_7694,N_5473);
xor U12175 (N_12175,N_7368,N_7372);
or U12176 (N_12176,N_5237,N_6704);
nand U12177 (N_12177,N_7743,N_8636);
and U12178 (N_12178,N_7889,N_7839);
and U12179 (N_12179,N_7024,N_9299);
or U12180 (N_12180,N_6868,N_7787);
or U12181 (N_12181,N_8288,N_6442);
and U12182 (N_12182,N_9169,N_5455);
and U12183 (N_12183,N_9138,N_6097);
and U12184 (N_12184,N_5752,N_7582);
and U12185 (N_12185,N_8931,N_6323);
and U12186 (N_12186,N_7799,N_6182);
nor U12187 (N_12187,N_6354,N_8449);
and U12188 (N_12188,N_9701,N_6145);
xor U12189 (N_12189,N_8552,N_5907);
or U12190 (N_12190,N_9684,N_9985);
xnor U12191 (N_12191,N_6005,N_5444);
and U12192 (N_12192,N_5616,N_7702);
nand U12193 (N_12193,N_7110,N_9530);
or U12194 (N_12194,N_7267,N_8948);
nor U12195 (N_12195,N_7966,N_6137);
nand U12196 (N_12196,N_8943,N_7891);
nand U12197 (N_12197,N_6388,N_7520);
or U12198 (N_12198,N_7676,N_6298);
nand U12199 (N_12199,N_6441,N_9111);
xor U12200 (N_12200,N_8892,N_5161);
xnor U12201 (N_12201,N_7071,N_7907);
and U12202 (N_12202,N_5723,N_8738);
nand U12203 (N_12203,N_5769,N_9063);
or U12204 (N_12204,N_7029,N_5954);
xnor U12205 (N_12205,N_9296,N_8384);
xor U12206 (N_12206,N_5537,N_5272);
nand U12207 (N_12207,N_6434,N_6330);
xor U12208 (N_12208,N_9334,N_7993);
xnor U12209 (N_12209,N_6879,N_6924);
and U12210 (N_12210,N_8185,N_6567);
and U12211 (N_12211,N_9192,N_8902);
and U12212 (N_12212,N_6624,N_8387);
nor U12213 (N_12213,N_9753,N_6675);
nor U12214 (N_12214,N_9323,N_8418);
nand U12215 (N_12215,N_7528,N_5751);
and U12216 (N_12216,N_5563,N_5422);
or U12217 (N_12217,N_6776,N_7514);
and U12218 (N_12218,N_6996,N_9959);
and U12219 (N_12219,N_9718,N_7897);
and U12220 (N_12220,N_8020,N_7934);
and U12221 (N_12221,N_9592,N_8323);
nand U12222 (N_12222,N_9482,N_6181);
xnor U12223 (N_12223,N_5781,N_7386);
nand U12224 (N_12224,N_5507,N_7928);
and U12225 (N_12225,N_8076,N_7722);
nor U12226 (N_12226,N_6292,N_8695);
or U12227 (N_12227,N_8040,N_7458);
or U12228 (N_12228,N_8028,N_6002);
or U12229 (N_12229,N_7917,N_8377);
and U12230 (N_12230,N_5139,N_7647);
xor U12231 (N_12231,N_5966,N_6658);
nand U12232 (N_12232,N_7559,N_6031);
nand U12233 (N_12233,N_6913,N_5844);
xor U12234 (N_12234,N_5617,N_6008);
nand U12235 (N_12235,N_9705,N_6682);
and U12236 (N_12236,N_6570,N_5700);
xnor U12237 (N_12237,N_6095,N_5543);
xnor U12238 (N_12238,N_5338,N_9738);
nand U12239 (N_12239,N_7626,N_6208);
and U12240 (N_12240,N_6135,N_5888);
or U12241 (N_12241,N_5129,N_9194);
nor U12242 (N_12242,N_7919,N_8726);
xnor U12243 (N_12243,N_6010,N_7565);
nor U12244 (N_12244,N_6712,N_8543);
nor U12245 (N_12245,N_8675,N_5263);
xor U12246 (N_12246,N_9496,N_6571);
xor U12247 (N_12247,N_7104,N_9094);
xor U12248 (N_12248,N_5711,N_7600);
and U12249 (N_12249,N_6359,N_6795);
xnor U12250 (N_12250,N_5411,N_9261);
or U12251 (N_12251,N_9423,N_5213);
nand U12252 (N_12252,N_7658,N_5124);
nor U12253 (N_12253,N_5482,N_6180);
nand U12254 (N_12254,N_6737,N_7505);
xor U12255 (N_12255,N_8568,N_9711);
nand U12256 (N_12256,N_9506,N_5417);
nor U12257 (N_12257,N_6932,N_7494);
xor U12258 (N_12258,N_6503,N_6527);
nor U12259 (N_12259,N_7901,N_9373);
and U12260 (N_12260,N_9537,N_8231);
and U12261 (N_12261,N_9968,N_8841);
and U12262 (N_12262,N_5817,N_7882);
nor U12263 (N_12263,N_9680,N_6210);
nor U12264 (N_12264,N_6798,N_8966);
and U12265 (N_12265,N_7516,N_8826);
xnor U12266 (N_12266,N_8445,N_6497);
and U12267 (N_12267,N_7307,N_7483);
xnor U12268 (N_12268,N_6902,N_9489);
and U12269 (N_12269,N_9987,N_8166);
xnor U12270 (N_12270,N_8813,N_6981);
xnor U12271 (N_12271,N_5056,N_5860);
xnor U12272 (N_12272,N_9271,N_7571);
nand U12273 (N_12273,N_9086,N_9264);
nor U12274 (N_12274,N_8987,N_6278);
nor U12275 (N_12275,N_6797,N_8138);
nand U12276 (N_12276,N_5476,N_6374);
nor U12277 (N_12277,N_7735,N_5833);
nand U12278 (N_12278,N_6926,N_6421);
xnor U12279 (N_12279,N_5491,N_5567);
nand U12280 (N_12280,N_5927,N_5727);
nor U12281 (N_12281,N_6423,N_8708);
or U12282 (N_12282,N_8406,N_6959);
and U12283 (N_12283,N_8027,N_5544);
or U12284 (N_12284,N_9609,N_8156);
xnor U12285 (N_12285,N_5454,N_6534);
nand U12286 (N_12286,N_9621,N_9837);
xnor U12287 (N_12287,N_8282,N_5383);
nand U12288 (N_12288,N_7515,N_7786);
nor U12289 (N_12289,N_6146,N_8934);
or U12290 (N_12290,N_8553,N_8562);
and U12291 (N_12291,N_6647,N_5993);
and U12292 (N_12292,N_8378,N_7292);
nor U12293 (N_12293,N_8254,N_7689);
nor U12294 (N_12294,N_5634,N_8910);
xnor U12295 (N_12295,N_6791,N_7167);
xnor U12296 (N_12296,N_8971,N_9671);
nor U12297 (N_12297,N_6425,N_8259);
nand U12298 (N_12298,N_6201,N_6236);
nor U12299 (N_12299,N_8188,N_7607);
and U12300 (N_12300,N_7191,N_5783);
xnor U12301 (N_12301,N_6612,N_6207);
nor U12302 (N_12302,N_9144,N_9298);
nand U12303 (N_12303,N_5250,N_7383);
and U12304 (N_12304,N_6050,N_9709);
nand U12305 (N_12305,N_6617,N_8472);
nor U12306 (N_12306,N_7022,N_5196);
nand U12307 (N_12307,N_9077,N_5147);
nor U12308 (N_12308,N_9662,N_7238);
nand U12309 (N_12309,N_9308,N_5945);
nor U12310 (N_12310,N_5651,N_5865);
nor U12311 (N_12311,N_9731,N_7087);
or U12312 (N_12312,N_7367,N_7992);
or U12313 (N_12313,N_8329,N_8698);
nor U12314 (N_12314,N_9336,N_6111);
or U12315 (N_12315,N_5428,N_8475);
nor U12316 (N_12316,N_7040,N_5295);
or U12317 (N_12317,N_6550,N_8529);
nand U12318 (N_12318,N_5210,N_6386);
xnor U12319 (N_12319,N_7620,N_6263);
nor U12320 (N_12320,N_9689,N_5906);
and U12321 (N_12321,N_9726,N_8542);
or U12322 (N_12322,N_9195,N_5126);
nor U12323 (N_12323,N_5753,N_5821);
xnor U12324 (N_12324,N_9162,N_6143);
nor U12325 (N_12325,N_8171,N_6375);
nand U12326 (N_12326,N_5362,N_5585);
nor U12327 (N_12327,N_6790,N_7981);
xnor U12328 (N_12328,N_8374,N_9306);
xor U12329 (N_12329,N_8646,N_8244);
and U12330 (N_12330,N_6342,N_9523);
nor U12331 (N_12331,N_6389,N_6702);
xor U12332 (N_12332,N_9199,N_7213);
nor U12333 (N_12333,N_6787,N_9917);
nor U12334 (N_12334,N_7790,N_9317);
and U12335 (N_12335,N_5812,N_5656);
nand U12336 (N_12336,N_7927,N_9504);
xor U12337 (N_12337,N_8838,N_6176);
nor U12338 (N_12338,N_9275,N_6450);
and U12339 (N_12339,N_5329,N_6398);
nand U12340 (N_12340,N_7397,N_6709);
nand U12341 (N_12341,N_7708,N_9902);
nand U12342 (N_12342,N_7989,N_6203);
nor U12343 (N_12343,N_6673,N_9799);
and U12344 (N_12344,N_6227,N_9436);
xnor U12345 (N_12345,N_5122,N_8438);
or U12346 (N_12346,N_9533,N_6679);
nor U12347 (N_12347,N_7533,N_6056);
xnor U12348 (N_12348,N_8471,N_8528);
and U12349 (N_12349,N_5492,N_7962);
nand U12350 (N_12350,N_6149,N_5183);
and U12351 (N_12351,N_9210,N_9786);
and U12352 (N_12352,N_6807,N_7156);
nand U12353 (N_12353,N_7824,N_7610);
or U12354 (N_12354,N_9091,N_5848);
nor U12355 (N_12355,N_8062,N_9607);
or U12356 (N_12356,N_8190,N_7319);
and U12357 (N_12357,N_7990,N_6928);
nor U12358 (N_12358,N_7111,N_8075);
xor U12359 (N_12359,N_7495,N_6426);
nand U12360 (N_12360,N_7969,N_7970);
and U12361 (N_12361,N_8547,N_7051);
nor U12362 (N_12362,N_5099,N_5892);
nand U12363 (N_12363,N_8820,N_6826);
nor U12364 (N_12364,N_9325,N_7282);
and U12365 (N_12365,N_9056,N_5386);
xor U12366 (N_12366,N_8868,N_7260);
nand U12367 (N_12367,N_9398,N_5204);
and U12368 (N_12368,N_7982,N_5447);
nand U12369 (N_12369,N_6720,N_9555);
nand U12370 (N_12370,N_7756,N_8453);
and U12371 (N_12371,N_6379,N_8593);
nand U12372 (N_12372,N_9329,N_7754);
nand U12373 (N_12373,N_9688,N_7447);
and U12374 (N_12374,N_8421,N_8341);
or U12375 (N_12375,N_5117,N_7244);
xnor U12376 (N_12376,N_8513,N_6671);
and U12377 (N_12377,N_9202,N_7558);
nor U12378 (N_12378,N_7617,N_6415);
nand U12379 (N_12379,N_6118,N_5828);
xor U12380 (N_12380,N_9544,N_7014);
nor U12381 (N_12381,N_7212,N_8295);
nand U12382 (N_12382,N_6351,N_7881);
or U12383 (N_12383,N_7601,N_5112);
nand U12384 (N_12384,N_5202,N_7015);
xnor U12385 (N_12385,N_7133,N_7652);
nor U12386 (N_12386,N_5093,N_6506);
nand U12387 (N_12387,N_6014,N_9740);
xor U12388 (N_12388,N_8180,N_5671);
nand U12389 (N_12389,N_9284,N_5481);
or U12390 (N_12390,N_9591,N_9825);
or U12391 (N_12391,N_9335,N_8872);
and U12392 (N_12392,N_7570,N_9017);
or U12393 (N_12393,N_9970,N_9480);
nor U12394 (N_12394,N_9626,N_9372);
or U12395 (N_12395,N_8879,N_9896);
xnor U12396 (N_12396,N_6838,N_6734);
nor U12397 (N_12397,N_6741,N_8376);
or U12398 (N_12398,N_8575,N_7682);
nor U12399 (N_12399,N_7597,N_7852);
nor U12400 (N_12400,N_9708,N_9833);
xor U12401 (N_12401,N_5793,N_8101);
or U12402 (N_12402,N_7877,N_5029);
and U12403 (N_12403,N_5999,N_9600);
and U12404 (N_12404,N_6502,N_8032);
nand U12405 (N_12405,N_5768,N_7139);
nor U12406 (N_12406,N_5197,N_6356);
nor U12407 (N_12407,N_9921,N_5583);
and U12408 (N_12408,N_6693,N_9168);
nor U12409 (N_12409,N_5058,N_6193);
xor U12410 (N_12410,N_9752,N_9706);
or U12411 (N_12411,N_8352,N_5718);
xor U12412 (N_12412,N_9241,N_8741);
or U12413 (N_12413,N_6321,N_6256);
xnor U12414 (N_12414,N_9388,N_7091);
xnor U12415 (N_12415,N_5983,N_9952);
nand U12416 (N_12416,N_5311,N_6308);
nor U12417 (N_12417,N_9172,N_5152);
or U12418 (N_12418,N_7833,N_9016);
or U12419 (N_12419,N_5784,N_6385);
and U12420 (N_12420,N_7838,N_9142);
xnor U12421 (N_12421,N_5978,N_6328);
and U12422 (N_12422,N_9758,N_5614);
xnor U12423 (N_12423,N_6127,N_8321);
xor U12424 (N_12424,N_9868,N_5675);
nor U12425 (N_12425,N_6888,N_8368);
or U12426 (N_12426,N_8610,N_5187);
and U12427 (N_12427,N_8920,N_7369);
nand U12428 (N_12428,N_7729,N_9910);
xnor U12429 (N_12429,N_8111,N_8574);
or U12430 (N_12430,N_6004,N_5542);
and U12431 (N_12431,N_6638,N_7556);
xor U12432 (N_12432,N_5934,N_5216);
nor U12433 (N_12433,N_9920,N_7239);
or U12434 (N_12434,N_7203,N_5572);
xnor U12435 (N_12435,N_7332,N_8317);
and U12436 (N_12436,N_6339,N_6481);
xor U12437 (N_12437,N_5920,N_9280);
nand U12438 (N_12438,N_5106,N_5955);
or U12439 (N_12439,N_7855,N_7073);
xnor U12440 (N_12440,N_9060,N_5027);
or U12441 (N_12441,N_9993,N_7293);
nor U12442 (N_12442,N_8013,N_8309);
and U12443 (N_12443,N_7362,N_9604);
nor U12444 (N_12444,N_9826,N_9578);
nand U12445 (N_12445,N_7526,N_7705);
nor U12446 (N_12446,N_9189,N_6914);
xor U12447 (N_12447,N_6384,N_5548);
nand U12448 (N_12448,N_7668,N_9446);
xor U12449 (N_12449,N_8541,N_9991);
nand U12450 (N_12450,N_7138,N_8015);
and U12451 (N_12451,N_7311,N_6910);
nand U12452 (N_12452,N_7460,N_7285);
nand U12453 (N_12453,N_5687,N_7903);
nor U12454 (N_12454,N_7544,N_5622);
or U12455 (N_12455,N_6250,N_5163);
or U12456 (N_12456,N_8995,N_7053);
nand U12457 (N_12457,N_6519,N_7291);
nand U12458 (N_12458,N_9447,N_6832);
nor U12459 (N_12459,N_6849,N_9624);
nand U12460 (N_12460,N_9152,N_8617);
nor U12461 (N_12461,N_6889,N_6304);
nand U12462 (N_12462,N_7968,N_5710);
nand U12463 (N_12463,N_5629,N_8870);
nand U12464 (N_12464,N_6305,N_5855);
nor U12465 (N_12465,N_8415,N_5804);
nor U12466 (N_12466,N_7554,N_9259);
and U12467 (N_12467,N_8773,N_8830);
and U12468 (N_12468,N_7697,N_8871);
nor U12469 (N_12469,N_6909,N_8671);
nor U12470 (N_12470,N_7480,N_8290);
nor U12471 (N_12471,N_8769,N_5337);
or U12472 (N_12472,N_9342,N_6535);
or U12473 (N_12473,N_9459,N_5759);
and U12474 (N_12474,N_5735,N_8606);
and U12475 (N_12475,N_6739,N_5148);
and U12476 (N_12476,N_7469,N_7013);
and U12477 (N_12477,N_5377,N_5241);
xor U12478 (N_12478,N_9742,N_7049);
or U12479 (N_12479,N_7745,N_7378);
or U12480 (N_12480,N_5363,N_9579);
and U12481 (N_12481,N_8939,N_9366);
or U12482 (N_12482,N_7090,N_6694);
or U12483 (N_12483,N_8768,N_5425);
and U12484 (N_12484,N_9490,N_8182);
or U12485 (N_12485,N_9792,N_5639);
nor U12486 (N_12486,N_5231,N_5480);
nor U12487 (N_12487,N_7663,N_5985);
or U12488 (N_12488,N_5119,N_5788);
and U12489 (N_12489,N_6669,N_7562);
nand U12490 (N_12490,N_6106,N_7535);
nor U12491 (N_12491,N_7219,N_6139);
nor U12492 (N_12492,N_6976,N_7914);
nor U12493 (N_12493,N_7761,N_7850);
nor U12494 (N_12494,N_8579,N_8973);
nor U12495 (N_12495,N_7868,N_9160);
and U12496 (N_12496,N_9451,N_7455);
nand U12497 (N_12497,N_5580,N_7083);
nand U12498 (N_12498,N_5517,N_5506);
xnor U12499 (N_12499,N_8464,N_6747);
or U12500 (N_12500,N_6756,N_9112);
nor U12501 (N_12501,N_7451,N_6309);
and U12502 (N_12502,N_7752,N_5882);
nor U12503 (N_12503,N_6383,N_6583);
or U12504 (N_12504,N_7579,N_7295);
or U12505 (N_12505,N_6264,N_8828);
nor U12506 (N_12506,N_7531,N_6292);
or U12507 (N_12507,N_5236,N_8769);
nor U12508 (N_12508,N_6165,N_9817);
nor U12509 (N_12509,N_9204,N_9056);
xor U12510 (N_12510,N_7593,N_7549);
nor U12511 (N_12511,N_7619,N_9137);
and U12512 (N_12512,N_9524,N_5586);
nor U12513 (N_12513,N_9089,N_7983);
and U12514 (N_12514,N_5243,N_5504);
nand U12515 (N_12515,N_8303,N_8963);
or U12516 (N_12516,N_5711,N_8694);
or U12517 (N_12517,N_8216,N_8124);
nor U12518 (N_12518,N_8156,N_6792);
or U12519 (N_12519,N_7071,N_9306);
xnor U12520 (N_12520,N_8194,N_8138);
nor U12521 (N_12521,N_9937,N_8295);
nor U12522 (N_12522,N_5820,N_8150);
or U12523 (N_12523,N_8205,N_9287);
xor U12524 (N_12524,N_7286,N_5493);
nor U12525 (N_12525,N_8712,N_5018);
xor U12526 (N_12526,N_9893,N_8879);
and U12527 (N_12527,N_6716,N_6337);
nand U12528 (N_12528,N_5308,N_9548);
or U12529 (N_12529,N_6611,N_5124);
and U12530 (N_12530,N_9745,N_8356);
xnor U12531 (N_12531,N_7318,N_9220);
nor U12532 (N_12532,N_5944,N_8452);
nor U12533 (N_12533,N_7990,N_5554);
nand U12534 (N_12534,N_9337,N_8724);
or U12535 (N_12535,N_7303,N_7513);
nand U12536 (N_12536,N_8076,N_7161);
and U12537 (N_12537,N_5291,N_6190);
and U12538 (N_12538,N_9908,N_7504);
nor U12539 (N_12539,N_9966,N_9030);
or U12540 (N_12540,N_9258,N_9574);
or U12541 (N_12541,N_6720,N_9543);
xor U12542 (N_12542,N_8201,N_8662);
or U12543 (N_12543,N_7892,N_8866);
and U12544 (N_12544,N_5663,N_8431);
nand U12545 (N_12545,N_7915,N_9170);
nor U12546 (N_12546,N_9403,N_6073);
or U12547 (N_12547,N_7565,N_9336);
xor U12548 (N_12548,N_5985,N_6984);
nand U12549 (N_12549,N_9770,N_7694);
xor U12550 (N_12550,N_8157,N_8284);
nand U12551 (N_12551,N_5047,N_7899);
or U12552 (N_12552,N_6577,N_7061);
nor U12553 (N_12553,N_9372,N_9571);
nand U12554 (N_12554,N_5681,N_5866);
xnor U12555 (N_12555,N_8020,N_8337);
nand U12556 (N_12556,N_5728,N_5443);
nand U12557 (N_12557,N_7342,N_6645);
nor U12558 (N_12558,N_8880,N_8683);
or U12559 (N_12559,N_5436,N_6740);
nor U12560 (N_12560,N_5406,N_6297);
nor U12561 (N_12561,N_9408,N_6117);
nand U12562 (N_12562,N_8136,N_9052);
or U12563 (N_12563,N_7989,N_7285);
and U12564 (N_12564,N_5953,N_9835);
xnor U12565 (N_12565,N_9886,N_6183);
xor U12566 (N_12566,N_7651,N_8485);
xor U12567 (N_12567,N_5624,N_6221);
nand U12568 (N_12568,N_7769,N_8889);
and U12569 (N_12569,N_9501,N_9759);
xnor U12570 (N_12570,N_6777,N_6825);
nand U12571 (N_12571,N_5549,N_8842);
xor U12572 (N_12572,N_8596,N_6338);
or U12573 (N_12573,N_7101,N_6350);
and U12574 (N_12574,N_5416,N_8222);
or U12575 (N_12575,N_6983,N_9359);
or U12576 (N_12576,N_9955,N_6456);
nand U12577 (N_12577,N_5266,N_5262);
and U12578 (N_12578,N_5185,N_9717);
and U12579 (N_12579,N_8315,N_5933);
xor U12580 (N_12580,N_7883,N_9933);
and U12581 (N_12581,N_8240,N_9569);
and U12582 (N_12582,N_6421,N_9757);
or U12583 (N_12583,N_9411,N_9609);
nand U12584 (N_12584,N_6383,N_5098);
and U12585 (N_12585,N_8859,N_9857);
xor U12586 (N_12586,N_9755,N_5287);
xor U12587 (N_12587,N_8236,N_5748);
or U12588 (N_12588,N_5060,N_5253);
and U12589 (N_12589,N_7938,N_6557);
nor U12590 (N_12590,N_7299,N_8163);
nand U12591 (N_12591,N_9202,N_8469);
and U12592 (N_12592,N_8510,N_9381);
nor U12593 (N_12593,N_5192,N_5888);
nand U12594 (N_12594,N_8756,N_8597);
xor U12595 (N_12595,N_6951,N_7342);
nand U12596 (N_12596,N_8039,N_6482);
and U12597 (N_12597,N_5792,N_7631);
and U12598 (N_12598,N_6387,N_8146);
nand U12599 (N_12599,N_8245,N_7055);
xor U12600 (N_12600,N_6127,N_6785);
nor U12601 (N_12601,N_7369,N_7153);
or U12602 (N_12602,N_6056,N_7146);
or U12603 (N_12603,N_8806,N_7731);
and U12604 (N_12604,N_6260,N_9879);
nor U12605 (N_12605,N_5915,N_7855);
nand U12606 (N_12606,N_8102,N_8865);
xnor U12607 (N_12607,N_7564,N_5454);
nand U12608 (N_12608,N_5435,N_7117);
and U12609 (N_12609,N_7847,N_6638);
and U12610 (N_12610,N_9896,N_7283);
nand U12611 (N_12611,N_5788,N_6565);
nor U12612 (N_12612,N_8596,N_5154);
nor U12613 (N_12613,N_8042,N_6331);
and U12614 (N_12614,N_7772,N_5162);
and U12615 (N_12615,N_8086,N_8974);
and U12616 (N_12616,N_9478,N_7728);
nand U12617 (N_12617,N_6796,N_7631);
and U12618 (N_12618,N_7394,N_6539);
and U12619 (N_12619,N_5296,N_6321);
xnor U12620 (N_12620,N_8664,N_9257);
xor U12621 (N_12621,N_5465,N_7772);
nor U12622 (N_12622,N_6099,N_7329);
or U12623 (N_12623,N_5737,N_7291);
nor U12624 (N_12624,N_9993,N_9931);
xnor U12625 (N_12625,N_7186,N_9328);
and U12626 (N_12626,N_5719,N_7191);
xnor U12627 (N_12627,N_6810,N_7980);
or U12628 (N_12628,N_7611,N_9602);
or U12629 (N_12629,N_5847,N_9559);
nor U12630 (N_12630,N_8093,N_9550);
or U12631 (N_12631,N_9803,N_7137);
or U12632 (N_12632,N_9048,N_7236);
nor U12633 (N_12633,N_6669,N_5693);
nor U12634 (N_12634,N_9236,N_6647);
and U12635 (N_12635,N_8073,N_6173);
and U12636 (N_12636,N_5707,N_7455);
and U12637 (N_12637,N_6987,N_5344);
and U12638 (N_12638,N_5708,N_8108);
xor U12639 (N_12639,N_9272,N_9246);
xor U12640 (N_12640,N_5435,N_6170);
nor U12641 (N_12641,N_7455,N_8791);
or U12642 (N_12642,N_8160,N_9573);
xor U12643 (N_12643,N_7173,N_8859);
nor U12644 (N_12644,N_5613,N_5895);
or U12645 (N_12645,N_9767,N_7170);
nor U12646 (N_12646,N_8801,N_7372);
xnor U12647 (N_12647,N_8876,N_9426);
or U12648 (N_12648,N_8309,N_6294);
xor U12649 (N_12649,N_9341,N_8202);
and U12650 (N_12650,N_6713,N_7093);
nand U12651 (N_12651,N_8808,N_5318);
xnor U12652 (N_12652,N_7862,N_8540);
and U12653 (N_12653,N_5441,N_9498);
nor U12654 (N_12654,N_7177,N_9523);
nand U12655 (N_12655,N_8149,N_8924);
nand U12656 (N_12656,N_7405,N_7263);
and U12657 (N_12657,N_5410,N_5741);
nand U12658 (N_12658,N_9489,N_5714);
xor U12659 (N_12659,N_6426,N_7864);
or U12660 (N_12660,N_5574,N_9013);
or U12661 (N_12661,N_7496,N_7390);
nor U12662 (N_12662,N_7029,N_7641);
or U12663 (N_12663,N_6378,N_5157);
xnor U12664 (N_12664,N_5444,N_9144);
xor U12665 (N_12665,N_6848,N_5376);
or U12666 (N_12666,N_6231,N_6472);
nor U12667 (N_12667,N_7906,N_6774);
and U12668 (N_12668,N_9930,N_5055);
nor U12669 (N_12669,N_9808,N_8635);
nor U12670 (N_12670,N_7581,N_5491);
xnor U12671 (N_12671,N_6194,N_5934);
or U12672 (N_12672,N_7455,N_7145);
nand U12673 (N_12673,N_5394,N_6680);
xor U12674 (N_12674,N_7022,N_9092);
or U12675 (N_12675,N_5295,N_8284);
xor U12676 (N_12676,N_6605,N_7163);
or U12677 (N_12677,N_8387,N_6617);
xor U12678 (N_12678,N_5081,N_5440);
and U12679 (N_12679,N_7370,N_8525);
nand U12680 (N_12680,N_7587,N_8522);
nor U12681 (N_12681,N_6368,N_8084);
xor U12682 (N_12682,N_9662,N_9684);
xnor U12683 (N_12683,N_5801,N_8908);
or U12684 (N_12684,N_5022,N_6922);
and U12685 (N_12685,N_9742,N_5730);
nor U12686 (N_12686,N_6510,N_6160);
and U12687 (N_12687,N_5294,N_5443);
nand U12688 (N_12688,N_8634,N_5166);
nor U12689 (N_12689,N_8016,N_9113);
nor U12690 (N_12690,N_9898,N_7889);
nand U12691 (N_12691,N_9094,N_6795);
xnor U12692 (N_12692,N_7639,N_6310);
xor U12693 (N_12693,N_7938,N_7206);
xnor U12694 (N_12694,N_7172,N_6680);
nor U12695 (N_12695,N_6200,N_9270);
or U12696 (N_12696,N_9259,N_5866);
and U12697 (N_12697,N_8485,N_9140);
xnor U12698 (N_12698,N_9705,N_8409);
or U12699 (N_12699,N_6175,N_9688);
and U12700 (N_12700,N_6888,N_5575);
nand U12701 (N_12701,N_9089,N_8519);
nor U12702 (N_12702,N_7435,N_7530);
xnor U12703 (N_12703,N_7720,N_5949);
or U12704 (N_12704,N_9006,N_5321);
nand U12705 (N_12705,N_8304,N_5603);
xor U12706 (N_12706,N_5444,N_7861);
nor U12707 (N_12707,N_8734,N_7142);
nor U12708 (N_12708,N_7393,N_5243);
and U12709 (N_12709,N_8969,N_5165);
xnor U12710 (N_12710,N_9553,N_5968);
and U12711 (N_12711,N_8368,N_6723);
nor U12712 (N_12712,N_5625,N_5304);
xnor U12713 (N_12713,N_7012,N_5446);
xor U12714 (N_12714,N_8855,N_9123);
and U12715 (N_12715,N_6705,N_9045);
xnor U12716 (N_12716,N_8623,N_6812);
and U12717 (N_12717,N_6409,N_6132);
xor U12718 (N_12718,N_5087,N_5179);
and U12719 (N_12719,N_8026,N_6954);
and U12720 (N_12720,N_5447,N_8748);
or U12721 (N_12721,N_8298,N_6746);
nand U12722 (N_12722,N_6321,N_9907);
and U12723 (N_12723,N_6624,N_5427);
nand U12724 (N_12724,N_7938,N_9495);
and U12725 (N_12725,N_5681,N_9130);
nand U12726 (N_12726,N_8600,N_6702);
or U12727 (N_12727,N_6088,N_9002);
nand U12728 (N_12728,N_5847,N_5966);
nand U12729 (N_12729,N_6869,N_9275);
or U12730 (N_12730,N_8679,N_6335);
nand U12731 (N_12731,N_5634,N_6721);
and U12732 (N_12732,N_9025,N_9291);
nand U12733 (N_12733,N_8864,N_6886);
xor U12734 (N_12734,N_6718,N_9181);
or U12735 (N_12735,N_6944,N_7489);
or U12736 (N_12736,N_6793,N_7617);
xnor U12737 (N_12737,N_8797,N_8479);
nor U12738 (N_12738,N_5023,N_9822);
or U12739 (N_12739,N_6061,N_9697);
nor U12740 (N_12740,N_5129,N_5444);
and U12741 (N_12741,N_5672,N_5608);
xnor U12742 (N_12742,N_8337,N_5074);
xor U12743 (N_12743,N_7791,N_7310);
xnor U12744 (N_12744,N_8819,N_8240);
or U12745 (N_12745,N_9227,N_6549);
nand U12746 (N_12746,N_8274,N_8349);
nor U12747 (N_12747,N_6721,N_9997);
nand U12748 (N_12748,N_7137,N_5279);
and U12749 (N_12749,N_9019,N_8587);
nand U12750 (N_12750,N_8065,N_7834);
and U12751 (N_12751,N_9937,N_9284);
nand U12752 (N_12752,N_5426,N_9271);
nand U12753 (N_12753,N_8304,N_5100);
xnor U12754 (N_12754,N_6583,N_9922);
or U12755 (N_12755,N_5849,N_7430);
and U12756 (N_12756,N_9886,N_6474);
nand U12757 (N_12757,N_7573,N_6182);
or U12758 (N_12758,N_8897,N_5283);
xnor U12759 (N_12759,N_9211,N_5590);
xor U12760 (N_12760,N_6247,N_9902);
and U12761 (N_12761,N_6863,N_7756);
and U12762 (N_12762,N_8114,N_8928);
and U12763 (N_12763,N_9023,N_7684);
nand U12764 (N_12764,N_7137,N_9364);
nand U12765 (N_12765,N_5807,N_6453);
or U12766 (N_12766,N_8112,N_6197);
xor U12767 (N_12767,N_8347,N_7847);
nor U12768 (N_12768,N_6316,N_7557);
and U12769 (N_12769,N_6123,N_9192);
nor U12770 (N_12770,N_6115,N_5666);
or U12771 (N_12771,N_6430,N_8792);
nand U12772 (N_12772,N_9152,N_7632);
nand U12773 (N_12773,N_5215,N_7735);
nor U12774 (N_12774,N_7460,N_6294);
xnor U12775 (N_12775,N_9419,N_8390);
and U12776 (N_12776,N_9733,N_6210);
nor U12777 (N_12777,N_5123,N_6709);
nand U12778 (N_12778,N_7512,N_9415);
or U12779 (N_12779,N_6690,N_9066);
nand U12780 (N_12780,N_9469,N_8901);
or U12781 (N_12781,N_8823,N_6539);
and U12782 (N_12782,N_8201,N_5862);
nor U12783 (N_12783,N_6279,N_5968);
or U12784 (N_12784,N_8386,N_5334);
xnor U12785 (N_12785,N_8463,N_6869);
and U12786 (N_12786,N_6444,N_9878);
and U12787 (N_12787,N_5781,N_8990);
xnor U12788 (N_12788,N_5573,N_7199);
or U12789 (N_12789,N_8465,N_9263);
nand U12790 (N_12790,N_9777,N_7423);
xor U12791 (N_12791,N_6259,N_7030);
or U12792 (N_12792,N_5330,N_7763);
xnor U12793 (N_12793,N_5353,N_5237);
xnor U12794 (N_12794,N_8580,N_8255);
or U12795 (N_12795,N_7631,N_5916);
or U12796 (N_12796,N_6369,N_8137);
nor U12797 (N_12797,N_5027,N_6703);
nand U12798 (N_12798,N_8622,N_9206);
xnor U12799 (N_12799,N_5976,N_9748);
nor U12800 (N_12800,N_5201,N_8345);
xor U12801 (N_12801,N_5488,N_5713);
xor U12802 (N_12802,N_7518,N_7526);
nor U12803 (N_12803,N_8710,N_8081);
nor U12804 (N_12804,N_7078,N_6715);
xnor U12805 (N_12805,N_8178,N_6039);
xnor U12806 (N_12806,N_6972,N_8936);
or U12807 (N_12807,N_7977,N_9964);
or U12808 (N_12808,N_7010,N_7209);
nor U12809 (N_12809,N_9359,N_9810);
or U12810 (N_12810,N_5022,N_7242);
nor U12811 (N_12811,N_8274,N_7130);
and U12812 (N_12812,N_7983,N_6557);
xor U12813 (N_12813,N_7206,N_9770);
nand U12814 (N_12814,N_5808,N_7174);
nor U12815 (N_12815,N_7244,N_9491);
nor U12816 (N_12816,N_9398,N_6198);
or U12817 (N_12817,N_7519,N_8095);
nand U12818 (N_12818,N_9450,N_7841);
and U12819 (N_12819,N_8384,N_6861);
nor U12820 (N_12820,N_7408,N_6758);
xor U12821 (N_12821,N_7530,N_9874);
or U12822 (N_12822,N_5446,N_9712);
xor U12823 (N_12823,N_7838,N_9495);
nand U12824 (N_12824,N_9113,N_6353);
nor U12825 (N_12825,N_7138,N_7599);
nor U12826 (N_12826,N_8571,N_9506);
nand U12827 (N_12827,N_7571,N_7726);
or U12828 (N_12828,N_8733,N_7785);
and U12829 (N_12829,N_7682,N_6459);
nand U12830 (N_12830,N_8570,N_7314);
and U12831 (N_12831,N_6857,N_8165);
nor U12832 (N_12832,N_9567,N_5634);
xnor U12833 (N_12833,N_8421,N_7158);
nor U12834 (N_12834,N_7390,N_5051);
xor U12835 (N_12835,N_9102,N_5398);
nand U12836 (N_12836,N_7730,N_5652);
or U12837 (N_12837,N_7808,N_7809);
nor U12838 (N_12838,N_5758,N_5850);
nand U12839 (N_12839,N_5331,N_8385);
nor U12840 (N_12840,N_8163,N_9498);
nand U12841 (N_12841,N_7591,N_8006);
xor U12842 (N_12842,N_8981,N_6165);
and U12843 (N_12843,N_8686,N_6287);
xnor U12844 (N_12844,N_5582,N_9044);
nor U12845 (N_12845,N_7929,N_5004);
or U12846 (N_12846,N_7784,N_8619);
nand U12847 (N_12847,N_9213,N_8183);
xnor U12848 (N_12848,N_6277,N_8579);
and U12849 (N_12849,N_8395,N_9498);
xor U12850 (N_12850,N_5920,N_7034);
or U12851 (N_12851,N_6488,N_9069);
and U12852 (N_12852,N_6822,N_7934);
nor U12853 (N_12853,N_6007,N_7823);
or U12854 (N_12854,N_9704,N_6184);
nand U12855 (N_12855,N_7197,N_9908);
and U12856 (N_12856,N_6746,N_9213);
or U12857 (N_12857,N_7785,N_7189);
xor U12858 (N_12858,N_5916,N_9374);
nand U12859 (N_12859,N_9158,N_5095);
nor U12860 (N_12860,N_6187,N_9885);
nor U12861 (N_12861,N_9586,N_9347);
nor U12862 (N_12862,N_8664,N_8149);
xor U12863 (N_12863,N_7421,N_5932);
and U12864 (N_12864,N_7890,N_6067);
nand U12865 (N_12865,N_8488,N_5592);
or U12866 (N_12866,N_9983,N_6888);
xor U12867 (N_12867,N_9621,N_9964);
xor U12868 (N_12868,N_6971,N_8028);
and U12869 (N_12869,N_7170,N_7432);
nor U12870 (N_12870,N_6514,N_9940);
and U12871 (N_12871,N_8569,N_7223);
nor U12872 (N_12872,N_5736,N_7545);
or U12873 (N_12873,N_5358,N_8509);
nand U12874 (N_12874,N_7464,N_7765);
nor U12875 (N_12875,N_5910,N_8669);
nor U12876 (N_12876,N_6455,N_6893);
or U12877 (N_12877,N_7593,N_9056);
and U12878 (N_12878,N_7291,N_7601);
nand U12879 (N_12879,N_9097,N_8649);
xnor U12880 (N_12880,N_9713,N_6792);
and U12881 (N_12881,N_8250,N_7208);
and U12882 (N_12882,N_9612,N_5421);
or U12883 (N_12883,N_8470,N_6006);
nor U12884 (N_12884,N_9846,N_6336);
or U12885 (N_12885,N_5317,N_7156);
nor U12886 (N_12886,N_7864,N_7612);
nor U12887 (N_12887,N_9930,N_5811);
or U12888 (N_12888,N_6684,N_8388);
nor U12889 (N_12889,N_6083,N_7324);
and U12890 (N_12890,N_6113,N_8025);
nand U12891 (N_12891,N_5974,N_6209);
and U12892 (N_12892,N_6839,N_7139);
or U12893 (N_12893,N_9050,N_5733);
and U12894 (N_12894,N_6866,N_8839);
and U12895 (N_12895,N_7081,N_5602);
nand U12896 (N_12896,N_9889,N_8071);
nor U12897 (N_12897,N_9995,N_8092);
nand U12898 (N_12898,N_9171,N_6933);
nor U12899 (N_12899,N_6565,N_7901);
xnor U12900 (N_12900,N_7297,N_5213);
nor U12901 (N_12901,N_8591,N_5909);
and U12902 (N_12902,N_6172,N_7492);
nand U12903 (N_12903,N_6990,N_9815);
xnor U12904 (N_12904,N_9273,N_7421);
nand U12905 (N_12905,N_9916,N_9769);
or U12906 (N_12906,N_9542,N_6036);
nand U12907 (N_12907,N_6650,N_9304);
nor U12908 (N_12908,N_6291,N_7526);
nor U12909 (N_12909,N_8577,N_9833);
or U12910 (N_12910,N_8077,N_7668);
nor U12911 (N_12911,N_6025,N_6818);
xnor U12912 (N_12912,N_8292,N_9695);
nand U12913 (N_12913,N_5236,N_5094);
nor U12914 (N_12914,N_6310,N_7761);
or U12915 (N_12915,N_5729,N_9122);
xor U12916 (N_12916,N_9809,N_5022);
or U12917 (N_12917,N_9718,N_9710);
xnor U12918 (N_12918,N_5352,N_8753);
nand U12919 (N_12919,N_7147,N_8938);
xor U12920 (N_12920,N_7108,N_6030);
nor U12921 (N_12921,N_7561,N_8999);
nor U12922 (N_12922,N_8568,N_5497);
xor U12923 (N_12923,N_6960,N_6107);
nand U12924 (N_12924,N_7505,N_6530);
nand U12925 (N_12925,N_5271,N_6793);
or U12926 (N_12926,N_7806,N_8433);
nor U12927 (N_12927,N_5487,N_9161);
or U12928 (N_12928,N_8271,N_6324);
nand U12929 (N_12929,N_7301,N_5351);
nor U12930 (N_12930,N_6962,N_9880);
nor U12931 (N_12931,N_9119,N_7433);
or U12932 (N_12932,N_9784,N_6937);
and U12933 (N_12933,N_7949,N_6797);
xnor U12934 (N_12934,N_9610,N_6182);
nand U12935 (N_12935,N_9565,N_5788);
nor U12936 (N_12936,N_9866,N_7909);
nand U12937 (N_12937,N_5958,N_5257);
and U12938 (N_12938,N_7088,N_8581);
xnor U12939 (N_12939,N_8620,N_8749);
xor U12940 (N_12940,N_5675,N_5084);
nor U12941 (N_12941,N_7309,N_8396);
or U12942 (N_12942,N_5532,N_7246);
xor U12943 (N_12943,N_5378,N_8872);
nand U12944 (N_12944,N_7819,N_7089);
nor U12945 (N_12945,N_5604,N_5687);
and U12946 (N_12946,N_5506,N_6680);
nor U12947 (N_12947,N_8439,N_5708);
or U12948 (N_12948,N_7755,N_7428);
xor U12949 (N_12949,N_5239,N_7871);
or U12950 (N_12950,N_8423,N_5512);
and U12951 (N_12951,N_7674,N_8602);
nor U12952 (N_12952,N_5848,N_9047);
xnor U12953 (N_12953,N_6235,N_5777);
nor U12954 (N_12954,N_6037,N_9310);
nor U12955 (N_12955,N_8551,N_7212);
nor U12956 (N_12956,N_8160,N_9615);
nand U12957 (N_12957,N_6090,N_6668);
nor U12958 (N_12958,N_5643,N_8906);
nand U12959 (N_12959,N_8477,N_8885);
xor U12960 (N_12960,N_5940,N_8571);
and U12961 (N_12961,N_6684,N_5937);
and U12962 (N_12962,N_5409,N_5628);
nor U12963 (N_12963,N_5399,N_9444);
nand U12964 (N_12964,N_6420,N_6915);
nand U12965 (N_12965,N_8888,N_8108);
nand U12966 (N_12966,N_6993,N_5601);
xor U12967 (N_12967,N_6867,N_5088);
and U12968 (N_12968,N_7239,N_6346);
xor U12969 (N_12969,N_5433,N_9583);
xor U12970 (N_12970,N_7127,N_5291);
xor U12971 (N_12971,N_5548,N_9094);
nor U12972 (N_12972,N_7298,N_9373);
nor U12973 (N_12973,N_8792,N_5695);
nand U12974 (N_12974,N_8945,N_8479);
xnor U12975 (N_12975,N_7844,N_5393);
xnor U12976 (N_12976,N_5309,N_7171);
or U12977 (N_12977,N_7133,N_8348);
nand U12978 (N_12978,N_6616,N_7676);
nor U12979 (N_12979,N_6123,N_8994);
or U12980 (N_12980,N_6463,N_6364);
or U12981 (N_12981,N_7482,N_9182);
nand U12982 (N_12982,N_6352,N_6241);
and U12983 (N_12983,N_9204,N_5691);
or U12984 (N_12984,N_9135,N_6715);
and U12985 (N_12985,N_8961,N_9013);
and U12986 (N_12986,N_8385,N_7770);
xor U12987 (N_12987,N_5333,N_9669);
nand U12988 (N_12988,N_7753,N_6335);
nand U12989 (N_12989,N_6633,N_9953);
and U12990 (N_12990,N_9515,N_9310);
xnor U12991 (N_12991,N_8220,N_7312);
and U12992 (N_12992,N_5135,N_6176);
or U12993 (N_12993,N_5934,N_6658);
and U12994 (N_12994,N_5698,N_5859);
and U12995 (N_12995,N_5931,N_6506);
or U12996 (N_12996,N_9657,N_7226);
nor U12997 (N_12997,N_5753,N_9768);
or U12998 (N_12998,N_7878,N_5404);
nand U12999 (N_12999,N_5103,N_9924);
nand U13000 (N_13000,N_7704,N_9708);
and U13001 (N_13001,N_7810,N_5375);
xnor U13002 (N_13002,N_8729,N_9321);
nand U13003 (N_13003,N_9612,N_6182);
nand U13004 (N_13004,N_5838,N_5072);
xor U13005 (N_13005,N_7934,N_7569);
or U13006 (N_13006,N_5322,N_8397);
xnor U13007 (N_13007,N_9318,N_6771);
or U13008 (N_13008,N_8703,N_5985);
nor U13009 (N_13009,N_9922,N_8708);
or U13010 (N_13010,N_9178,N_8619);
or U13011 (N_13011,N_6940,N_8144);
nor U13012 (N_13012,N_6113,N_7622);
nor U13013 (N_13013,N_6959,N_8292);
nand U13014 (N_13014,N_6351,N_5052);
xor U13015 (N_13015,N_8182,N_8091);
and U13016 (N_13016,N_8458,N_7439);
and U13017 (N_13017,N_6446,N_5032);
nor U13018 (N_13018,N_7458,N_6249);
nand U13019 (N_13019,N_5666,N_8008);
nor U13020 (N_13020,N_7697,N_6702);
nand U13021 (N_13021,N_5784,N_5036);
nor U13022 (N_13022,N_5123,N_5673);
nor U13023 (N_13023,N_8327,N_8968);
xor U13024 (N_13024,N_9787,N_8373);
nand U13025 (N_13025,N_7737,N_7241);
and U13026 (N_13026,N_6771,N_9015);
nor U13027 (N_13027,N_9235,N_8030);
nand U13028 (N_13028,N_6605,N_9501);
and U13029 (N_13029,N_7631,N_6903);
and U13030 (N_13030,N_7713,N_9916);
or U13031 (N_13031,N_8985,N_7499);
or U13032 (N_13032,N_5310,N_6594);
nand U13033 (N_13033,N_8405,N_6520);
nand U13034 (N_13034,N_9185,N_6423);
or U13035 (N_13035,N_6123,N_9648);
nor U13036 (N_13036,N_8011,N_5942);
or U13037 (N_13037,N_5655,N_5234);
nand U13038 (N_13038,N_5805,N_8642);
xor U13039 (N_13039,N_7980,N_5808);
and U13040 (N_13040,N_6191,N_9189);
nand U13041 (N_13041,N_6064,N_5395);
nor U13042 (N_13042,N_8483,N_8104);
and U13043 (N_13043,N_5486,N_9078);
nand U13044 (N_13044,N_6506,N_9616);
nand U13045 (N_13045,N_8485,N_9975);
and U13046 (N_13046,N_6162,N_5927);
or U13047 (N_13047,N_6218,N_5633);
or U13048 (N_13048,N_5473,N_9420);
xor U13049 (N_13049,N_8009,N_9336);
xnor U13050 (N_13050,N_6010,N_9132);
nor U13051 (N_13051,N_5284,N_8871);
xnor U13052 (N_13052,N_6997,N_7106);
or U13053 (N_13053,N_7963,N_6871);
nand U13054 (N_13054,N_8709,N_8376);
or U13055 (N_13055,N_8581,N_5577);
nor U13056 (N_13056,N_5906,N_5741);
and U13057 (N_13057,N_9912,N_8660);
or U13058 (N_13058,N_7987,N_7283);
nand U13059 (N_13059,N_9791,N_5489);
nor U13060 (N_13060,N_7458,N_8470);
xnor U13061 (N_13061,N_5328,N_7970);
nand U13062 (N_13062,N_7554,N_7870);
nor U13063 (N_13063,N_5280,N_8185);
xor U13064 (N_13064,N_7701,N_5080);
nand U13065 (N_13065,N_9464,N_7609);
nand U13066 (N_13066,N_8691,N_8894);
nand U13067 (N_13067,N_7854,N_8868);
nand U13068 (N_13068,N_7037,N_6063);
nand U13069 (N_13069,N_8765,N_7427);
and U13070 (N_13070,N_7541,N_6996);
nand U13071 (N_13071,N_6946,N_6249);
nand U13072 (N_13072,N_6690,N_6779);
nand U13073 (N_13073,N_8004,N_5512);
nor U13074 (N_13074,N_9151,N_7862);
and U13075 (N_13075,N_7520,N_7316);
nand U13076 (N_13076,N_6341,N_7701);
or U13077 (N_13077,N_6619,N_9354);
and U13078 (N_13078,N_6659,N_9560);
or U13079 (N_13079,N_8571,N_7418);
nand U13080 (N_13080,N_8203,N_6125);
xor U13081 (N_13081,N_8974,N_5356);
and U13082 (N_13082,N_6555,N_9414);
nor U13083 (N_13083,N_8743,N_5497);
or U13084 (N_13084,N_7204,N_8531);
xor U13085 (N_13085,N_8190,N_5300);
and U13086 (N_13086,N_8342,N_7726);
nor U13087 (N_13087,N_8150,N_6056);
and U13088 (N_13088,N_8052,N_9587);
or U13089 (N_13089,N_9749,N_6345);
and U13090 (N_13090,N_7445,N_8331);
and U13091 (N_13091,N_8600,N_9794);
or U13092 (N_13092,N_9906,N_5099);
xor U13093 (N_13093,N_7128,N_6275);
or U13094 (N_13094,N_8401,N_5247);
nand U13095 (N_13095,N_7719,N_8724);
xor U13096 (N_13096,N_5437,N_7344);
nand U13097 (N_13097,N_7137,N_5712);
nor U13098 (N_13098,N_8499,N_9513);
or U13099 (N_13099,N_9053,N_5046);
or U13100 (N_13100,N_9570,N_7356);
nor U13101 (N_13101,N_8113,N_9903);
and U13102 (N_13102,N_9079,N_5808);
nand U13103 (N_13103,N_7976,N_9669);
nand U13104 (N_13104,N_8590,N_5415);
or U13105 (N_13105,N_8117,N_9808);
or U13106 (N_13106,N_7521,N_5551);
nor U13107 (N_13107,N_7403,N_6688);
nor U13108 (N_13108,N_6332,N_9720);
and U13109 (N_13109,N_6457,N_6701);
and U13110 (N_13110,N_9239,N_5883);
xor U13111 (N_13111,N_6721,N_7906);
nand U13112 (N_13112,N_9651,N_6572);
nand U13113 (N_13113,N_6966,N_8340);
and U13114 (N_13114,N_6427,N_6498);
and U13115 (N_13115,N_8376,N_5402);
nor U13116 (N_13116,N_6833,N_8740);
nand U13117 (N_13117,N_6892,N_8376);
and U13118 (N_13118,N_9061,N_6245);
nor U13119 (N_13119,N_7467,N_6286);
and U13120 (N_13120,N_9814,N_5872);
xor U13121 (N_13121,N_5842,N_7011);
nand U13122 (N_13122,N_8456,N_5502);
and U13123 (N_13123,N_7204,N_5694);
or U13124 (N_13124,N_6250,N_6597);
nand U13125 (N_13125,N_6130,N_6023);
or U13126 (N_13126,N_7793,N_5365);
nand U13127 (N_13127,N_8906,N_6402);
or U13128 (N_13128,N_5835,N_7141);
nor U13129 (N_13129,N_6767,N_5701);
or U13130 (N_13130,N_7974,N_6420);
xnor U13131 (N_13131,N_9514,N_7902);
or U13132 (N_13132,N_9522,N_7434);
or U13133 (N_13133,N_6230,N_9550);
nor U13134 (N_13134,N_6956,N_5542);
xnor U13135 (N_13135,N_6648,N_8184);
xnor U13136 (N_13136,N_8810,N_7662);
nand U13137 (N_13137,N_8119,N_8351);
xor U13138 (N_13138,N_8822,N_6755);
nor U13139 (N_13139,N_7917,N_9720);
and U13140 (N_13140,N_7091,N_8326);
nand U13141 (N_13141,N_9604,N_5192);
xor U13142 (N_13142,N_7212,N_9215);
xnor U13143 (N_13143,N_6854,N_6875);
and U13144 (N_13144,N_5808,N_8837);
nand U13145 (N_13145,N_5406,N_5472);
nor U13146 (N_13146,N_8748,N_7836);
or U13147 (N_13147,N_6158,N_9904);
nand U13148 (N_13148,N_6208,N_5065);
and U13149 (N_13149,N_9717,N_5313);
or U13150 (N_13150,N_8900,N_9047);
nor U13151 (N_13151,N_9106,N_6585);
nor U13152 (N_13152,N_8875,N_9989);
nand U13153 (N_13153,N_5242,N_8427);
and U13154 (N_13154,N_7435,N_5433);
nand U13155 (N_13155,N_6007,N_5972);
xor U13156 (N_13156,N_6121,N_6194);
nand U13157 (N_13157,N_6827,N_7432);
and U13158 (N_13158,N_5697,N_7364);
and U13159 (N_13159,N_7387,N_5438);
and U13160 (N_13160,N_9689,N_8903);
xnor U13161 (N_13161,N_7736,N_9026);
nor U13162 (N_13162,N_7019,N_7542);
and U13163 (N_13163,N_5946,N_6819);
nor U13164 (N_13164,N_7385,N_9278);
xnor U13165 (N_13165,N_9904,N_7032);
and U13166 (N_13166,N_6409,N_8560);
or U13167 (N_13167,N_7846,N_7362);
nor U13168 (N_13168,N_7466,N_9678);
nand U13169 (N_13169,N_7122,N_5480);
and U13170 (N_13170,N_9171,N_6809);
xnor U13171 (N_13171,N_8661,N_9882);
and U13172 (N_13172,N_5965,N_5653);
and U13173 (N_13173,N_7884,N_5155);
and U13174 (N_13174,N_7028,N_6893);
nor U13175 (N_13175,N_8909,N_5277);
and U13176 (N_13176,N_9385,N_7240);
xor U13177 (N_13177,N_9025,N_8232);
nand U13178 (N_13178,N_5528,N_8576);
xor U13179 (N_13179,N_7043,N_8387);
nor U13180 (N_13180,N_6016,N_8250);
xor U13181 (N_13181,N_5499,N_5598);
nor U13182 (N_13182,N_7767,N_8231);
xnor U13183 (N_13183,N_7718,N_8977);
or U13184 (N_13184,N_5419,N_9202);
nand U13185 (N_13185,N_8716,N_7418);
xor U13186 (N_13186,N_6444,N_7907);
or U13187 (N_13187,N_7486,N_5353);
nand U13188 (N_13188,N_8544,N_8078);
nand U13189 (N_13189,N_8896,N_9342);
and U13190 (N_13190,N_9260,N_6373);
and U13191 (N_13191,N_8735,N_5472);
xnor U13192 (N_13192,N_6360,N_8971);
nor U13193 (N_13193,N_9833,N_5641);
and U13194 (N_13194,N_5764,N_6125);
xor U13195 (N_13195,N_7466,N_8173);
xnor U13196 (N_13196,N_9357,N_6336);
xnor U13197 (N_13197,N_8547,N_7781);
or U13198 (N_13198,N_8648,N_9935);
nor U13199 (N_13199,N_7200,N_9895);
and U13200 (N_13200,N_8761,N_9061);
nand U13201 (N_13201,N_5810,N_6554);
and U13202 (N_13202,N_9355,N_9929);
nor U13203 (N_13203,N_8824,N_7247);
xnor U13204 (N_13204,N_8123,N_9925);
nor U13205 (N_13205,N_5151,N_5268);
or U13206 (N_13206,N_7877,N_7535);
or U13207 (N_13207,N_9094,N_8799);
nor U13208 (N_13208,N_5074,N_5290);
nand U13209 (N_13209,N_8544,N_5866);
nand U13210 (N_13210,N_9322,N_7120);
or U13211 (N_13211,N_6131,N_5903);
nand U13212 (N_13212,N_5914,N_6784);
nor U13213 (N_13213,N_6547,N_5720);
xnor U13214 (N_13214,N_5449,N_7942);
xor U13215 (N_13215,N_9718,N_6952);
and U13216 (N_13216,N_6084,N_6737);
nand U13217 (N_13217,N_9346,N_9073);
nand U13218 (N_13218,N_8170,N_7749);
and U13219 (N_13219,N_9993,N_5935);
xor U13220 (N_13220,N_7160,N_7588);
nor U13221 (N_13221,N_6660,N_5540);
or U13222 (N_13222,N_5933,N_6219);
or U13223 (N_13223,N_9313,N_9483);
xor U13224 (N_13224,N_7901,N_8911);
xnor U13225 (N_13225,N_5323,N_5161);
nand U13226 (N_13226,N_8211,N_6675);
nand U13227 (N_13227,N_7794,N_7277);
or U13228 (N_13228,N_9102,N_9932);
nand U13229 (N_13229,N_8705,N_6206);
nor U13230 (N_13230,N_8431,N_6063);
xor U13231 (N_13231,N_5957,N_7127);
or U13232 (N_13232,N_7962,N_6801);
nor U13233 (N_13233,N_8445,N_7125);
or U13234 (N_13234,N_9534,N_5688);
nor U13235 (N_13235,N_5648,N_6116);
and U13236 (N_13236,N_6079,N_6006);
and U13237 (N_13237,N_8709,N_6149);
nor U13238 (N_13238,N_8064,N_8286);
nand U13239 (N_13239,N_6810,N_7198);
nor U13240 (N_13240,N_9479,N_8744);
nand U13241 (N_13241,N_9930,N_5489);
and U13242 (N_13242,N_7830,N_7963);
nor U13243 (N_13243,N_6715,N_6449);
xnor U13244 (N_13244,N_8493,N_8536);
or U13245 (N_13245,N_5233,N_9931);
or U13246 (N_13246,N_9315,N_6667);
nand U13247 (N_13247,N_8955,N_9233);
xnor U13248 (N_13248,N_6766,N_7053);
nor U13249 (N_13249,N_7711,N_9868);
and U13250 (N_13250,N_5201,N_7289);
nor U13251 (N_13251,N_7783,N_8900);
nand U13252 (N_13252,N_8050,N_9852);
or U13253 (N_13253,N_8255,N_9532);
and U13254 (N_13254,N_9116,N_6979);
and U13255 (N_13255,N_7922,N_7930);
and U13256 (N_13256,N_5851,N_6985);
and U13257 (N_13257,N_7405,N_7688);
xnor U13258 (N_13258,N_6342,N_9464);
nor U13259 (N_13259,N_5697,N_7154);
xnor U13260 (N_13260,N_9732,N_5720);
xnor U13261 (N_13261,N_7040,N_8473);
xnor U13262 (N_13262,N_9203,N_7397);
nor U13263 (N_13263,N_7507,N_6276);
or U13264 (N_13264,N_6077,N_6876);
xnor U13265 (N_13265,N_6026,N_9878);
nor U13266 (N_13266,N_8666,N_5091);
and U13267 (N_13267,N_8295,N_7591);
xor U13268 (N_13268,N_9372,N_9729);
xor U13269 (N_13269,N_9816,N_8608);
xnor U13270 (N_13270,N_9076,N_9449);
nand U13271 (N_13271,N_6971,N_6239);
or U13272 (N_13272,N_5917,N_8274);
and U13273 (N_13273,N_8465,N_7509);
and U13274 (N_13274,N_8830,N_5502);
and U13275 (N_13275,N_9394,N_8026);
and U13276 (N_13276,N_5601,N_6959);
nor U13277 (N_13277,N_5601,N_8082);
and U13278 (N_13278,N_8909,N_5387);
and U13279 (N_13279,N_7146,N_9272);
nor U13280 (N_13280,N_8526,N_7562);
and U13281 (N_13281,N_8260,N_8867);
and U13282 (N_13282,N_5782,N_5471);
or U13283 (N_13283,N_5240,N_6714);
xor U13284 (N_13284,N_9871,N_5086);
or U13285 (N_13285,N_8290,N_6370);
xor U13286 (N_13286,N_7010,N_6144);
and U13287 (N_13287,N_9931,N_6812);
nand U13288 (N_13288,N_7236,N_9542);
nor U13289 (N_13289,N_7203,N_7324);
nor U13290 (N_13290,N_5484,N_9056);
and U13291 (N_13291,N_5971,N_5645);
nand U13292 (N_13292,N_7082,N_7875);
and U13293 (N_13293,N_6591,N_8365);
nand U13294 (N_13294,N_6653,N_9508);
xor U13295 (N_13295,N_8970,N_5329);
xnor U13296 (N_13296,N_7555,N_7913);
nor U13297 (N_13297,N_7833,N_6141);
nand U13298 (N_13298,N_5466,N_7473);
xor U13299 (N_13299,N_7684,N_9719);
nor U13300 (N_13300,N_9942,N_7341);
nor U13301 (N_13301,N_5236,N_7212);
and U13302 (N_13302,N_9691,N_5992);
nor U13303 (N_13303,N_9503,N_7850);
and U13304 (N_13304,N_6452,N_9616);
or U13305 (N_13305,N_5585,N_5410);
nor U13306 (N_13306,N_8715,N_7964);
nand U13307 (N_13307,N_7441,N_7853);
and U13308 (N_13308,N_7908,N_9928);
nand U13309 (N_13309,N_7915,N_8528);
xor U13310 (N_13310,N_5067,N_8934);
or U13311 (N_13311,N_5585,N_9384);
or U13312 (N_13312,N_8214,N_6845);
nand U13313 (N_13313,N_5481,N_6818);
and U13314 (N_13314,N_6847,N_5101);
nand U13315 (N_13315,N_7616,N_5869);
nor U13316 (N_13316,N_8403,N_5766);
nand U13317 (N_13317,N_8499,N_8893);
and U13318 (N_13318,N_6772,N_5192);
nand U13319 (N_13319,N_5674,N_7176);
or U13320 (N_13320,N_9013,N_9251);
and U13321 (N_13321,N_8580,N_9958);
or U13322 (N_13322,N_5472,N_6717);
or U13323 (N_13323,N_7580,N_8182);
and U13324 (N_13324,N_9825,N_8363);
xor U13325 (N_13325,N_8839,N_7761);
nand U13326 (N_13326,N_7972,N_9293);
xnor U13327 (N_13327,N_7999,N_7768);
or U13328 (N_13328,N_9696,N_9941);
or U13329 (N_13329,N_5063,N_9110);
nor U13330 (N_13330,N_7673,N_5681);
xnor U13331 (N_13331,N_5815,N_8095);
or U13332 (N_13332,N_8059,N_7619);
nor U13333 (N_13333,N_8185,N_6341);
nand U13334 (N_13334,N_9350,N_8635);
or U13335 (N_13335,N_6834,N_7883);
nand U13336 (N_13336,N_9422,N_8584);
or U13337 (N_13337,N_5314,N_5571);
nor U13338 (N_13338,N_7557,N_5363);
nor U13339 (N_13339,N_5004,N_5137);
nand U13340 (N_13340,N_7449,N_8049);
nor U13341 (N_13341,N_6033,N_7099);
and U13342 (N_13342,N_5487,N_6207);
nand U13343 (N_13343,N_8824,N_6196);
xnor U13344 (N_13344,N_9418,N_7640);
xor U13345 (N_13345,N_6777,N_9643);
or U13346 (N_13346,N_9887,N_5656);
and U13347 (N_13347,N_9925,N_6270);
nand U13348 (N_13348,N_7301,N_7778);
nand U13349 (N_13349,N_9784,N_8271);
and U13350 (N_13350,N_9418,N_8603);
and U13351 (N_13351,N_7560,N_5250);
and U13352 (N_13352,N_5407,N_5833);
nor U13353 (N_13353,N_8380,N_5527);
or U13354 (N_13354,N_9357,N_8014);
nor U13355 (N_13355,N_7125,N_5777);
nor U13356 (N_13356,N_7047,N_9082);
xor U13357 (N_13357,N_8160,N_9327);
nand U13358 (N_13358,N_9384,N_9731);
nor U13359 (N_13359,N_8224,N_8142);
or U13360 (N_13360,N_9650,N_6601);
and U13361 (N_13361,N_6532,N_8976);
nor U13362 (N_13362,N_8982,N_5238);
and U13363 (N_13363,N_8100,N_9478);
and U13364 (N_13364,N_8890,N_7693);
and U13365 (N_13365,N_8431,N_6862);
nand U13366 (N_13366,N_7420,N_7039);
nor U13367 (N_13367,N_7172,N_7351);
xor U13368 (N_13368,N_5677,N_8425);
xnor U13369 (N_13369,N_8742,N_6387);
nand U13370 (N_13370,N_9777,N_8475);
xor U13371 (N_13371,N_9118,N_5405);
nand U13372 (N_13372,N_9147,N_8728);
and U13373 (N_13373,N_5287,N_7818);
or U13374 (N_13374,N_8356,N_9037);
xor U13375 (N_13375,N_6179,N_6713);
nor U13376 (N_13376,N_7881,N_6078);
xor U13377 (N_13377,N_7107,N_6460);
xnor U13378 (N_13378,N_5232,N_6828);
nand U13379 (N_13379,N_6755,N_7291);
xnor U13380 (N_13380,N_9420,N_9318);
or U13381 (N_13381,N_8995,N_8599);
nor U13382 (N_13382,N_7146,N_6023);
or U13383 (N_13383,N_5082,N_8608);
nand U13384 (N_13384,N_7835,N_9305);
nand U13385 (N_13385,N_6142,N_8818);
and U13386 (N_13386,N_9055,N_8206);
xnor U13387 (N_13387,N_8853,N_8135);
nor U13388 (N_13388,N_7782,N_9862);
or U13389 (N_13389,N_7999,N_8269);
or U13390 (N_13390,N_5587,N_6950);
nand U13391 (N_13391,N_6733,N_7040);
xnor U13392 (N_13392,N_7665,N_6243);
nor U13393 (N_13393,N_7682,N_6805);
and U13394 (N_13394,N_6674,N_8787);
or U13395 (N_13395,N_9943,N_5671);
xnor U13396 (N_13396,N_9637,N_6572);
nor U13397 (N_13397,N_9662,N_7236);
nor U13398 (N_13398,N_9596,N_5237);
and U13399 (N_13399,N_5551,N_5534);
and U13400 (N_13400,N_5360,N_8843);
nor U13401 (N_13401,N_7633,N_7048);
nor U13402 (N_13402,N_9249,N_9194);
nor U13403 (N_13403,N_7931,N_7324);
xnor U13404 (N_13404,N_6887,N_5240);
nand U13405 (N_13405,N_7726,N_9093);
and U13406 (N_13406,N_8766,N_8858);
or U13407 (N_13407,N_5031,N_7957);
nor U13408 (N_13408,N_8305,N_6715);
xor U13409 (N_13409,N_8013,N_9781);
nor U13410 (N_13410,N_6198,N_9851);
nor U13411 (N_13411,N_5848,N_8088);
xnor U13412 (N_13412,N_8976,N_7488);
nand U13413 (N_13413,N_7046,N_9265);
or U13414 (N_13414,N_9043,N_9045);
xnor U13415 (N_13415,N_6713,N_9814);
xnor U13416 (N_13416,N_7777,N_9442);
and U13417 (N_13417,N_8523,N_6711);
or U13418 (N_13418,N_8063,N_5801);
xnor U13419 (N_13419,N_8234,N_5528);
and U13420 (N_13420,N_6700,N_6904);
nor U13421 (N_13421,N_7333,N_7384);
or U13422 (N_13422,N_6223,N_7214);
nand U13423 (N_13423,N_6580,N_7035);
nand U13424 (N_13424,N_6230,N_6292);
nand U13425 (N_13425,N_7687,N_8023);
and U13426 (N_13426,N_5280,N_5512);
and U13427 (N_13427,N_8712,N_7593);
xnor U13428 (N_13428,N_6864,N_7067);
or U13429 (N_13429,N_8125,N_9733);
xor U13430 (N_13430,N_8006,N_9782);
nand U13431 (N_13431,N_6951,N_6810);
nand U13432 (N_13432,N_7676,N_7690);
and U13433 (N_13433,N_5431,N_7336);
xnor U13434 (N_13434,N_9384,N_5454);
or U13435 (N_13435,N_8368,N_5959);
nand U13436 (N_13436,N_7905,N_9485);
xnor U13437 (N_13437,N_6877,N_7035);
or U13438 (N_13438,N_5069,N_9526);
and U13439 (N_13439,N_9371,N_5671);
nor U13440 (N_13440,N_5571,N_5684);
nand U13441 (N_13441,N_7273,N_7218);
xor U13442 (N_13442,N_7463,N_6983);
nor U13443 (N_13443,N_9799,N_6109);
nor U13444 (N_13444,N_9651,N_8778);
nand U13445 (N_13445,N_5694,N_5322);
nor U13446 (N_13446,N_6016,N_9318);
nor U13447 (N_13447,N_5729,N_8249);
xor U13448 (N_13448,N_6133,N_5068);
nand U13449 (N_13449,N_8247,N_6535);
or U13450 (N_13450,N_7507,N_9164);
nor U13451 (N_13451,N_6613,N_8690);
or U13452 (N_13452,N_9321,N_5764);
or U13453 (N_13453,N_6927,N_9244);
nor U13454 (N_13454,N_5723,N_5140);
and U13455 (N_13455,N_9683,N_8487);
or U13456 (N_13456,N_8913,N_6011);
nand U13457 (N_13457,N_7536,N_6159);
xnor U13458 (N_13458,N_5746,N_7303);
and U13459 (N_13459,N_9866,N_6787);
and U13460 (N_13460,N_6002,N_6606);
nor U13461 (N_13461,N_5215,N_9572);
xnor U13462 (N_13462,N_8184,N_9250);
xor U13463 (N_13463,N_7936,N_5245);
nand U13464 (N_13464,N_6796,N_7852);
nand U13465 (N_13465,N_5402,N_8068);
nand U13466 (N_13466,N_5874,N_5800);
and U13467 (N_13467,N_6788,N_5341);
or U13468 (N_13468,N_5959,N_8353);
and U13469 (N_13469,N_6804,N_8975);
or U13470 (N_13470,N_8936,N_5834);
and U13471 (N_13471,N_6988,N_8620);
nand U13472 (N_13472,N_6637,N_6312);
and U13473 (N_13473,N_8095,N_5164);
and U13474 (N_13474,N_7626,N_5923);
and U13475 (N_13475,N_8474,N_9763);
or U13476 (N_13476,N_7348,N_8740);
and U13477 (N_13477,N_7774,N_9286);
or U13478 (N_13478,N_8624,N_6476);
xnor U13479 (N_13479,N_9668,N_7971);
xor U13480 (N_13480,N_8211,N_9401);
and U13481 (N_13481,N_7256,N_6730);
xor U13482 (N_13482,N_7439,N_6480);
or U13483 (N_13483,N_7981,N_6630);
and U13484 (N_13484,N_6713,N_8456);
xor U13485 (N_13485,N_5080,N_7290);
xnor U13486 (N_13486,N_9046,N_8519);
or U13487 (N_13487,N_9333,N_7882);
or U13488 (N_13488,N_8198,N_8789);
xnor U13489 (N_13489,N_5275,N_5081);
xor U13490 (N_13490,N_6082,N_8279);
or U13491 (N_13491,N_7038,N_6668);
or U13492 (N_13492,N_8663,N_7370);
nand U13493 (N_13493,N_5954,N_5697);
nor U13494 (N_13494,N_7475,N_6151);
nor U13495 (N_13495,N_6323,N_5766);
and U13496 (N_13496,N_9763,N_8940);
xor U13497 (N_13497,N_7269,N_9506);
and U13498 (N_13498,N_5009,N_6523);
and U13499 (N_13499,N_7475,N_9546);
xor U13500 (N_13500,N_5602,N_6100);
nand U13501 (N_13501,N_8441,N_5529);
xnor U13502 (N_13502,N_7721,N_7695);
nand U13503 (N_13503,N_8752,N_7379);
or U13504 (N_13504,N_9708,N_8031);
nand U13505 (N_13505,N_6236,N_8556);
xnor U13506 (N_13506,N_8740,N_5461);
nand U13507 (N_13507,N_9509,N_5067);
nor U13508 (N_13508,N_9468,N_7221);
and U13509 (N_13509,N_7179,N_5926);
nand U13510 (N_13510,N_9877,N_8541);
xnor U13511 (N_13511,N_8977,N_9067);
nor U13512 (N_13512,N_9578,N_9038);
or U13513 (N_13513,N_9979,N_5346);
nand U13514 (N_13514,N_8933,N_6020);
nand U13515 (N_13515,N_7768,N_6896);
xor U13516 (N_13516,N_9988,N_6564);
nor U13517 (N_13517,N_5940,N_5957);
or U13518 (N_13518,N_7158,N_5617);
nor U13519 (N_13519,N_7037,N_6406);
xnor U13520 (N_13520,N_5808,N_7978);
and U13521 (N_13521,N_8335,N_6382);
nor U13522 (N_13522,N_7538,N_6644);
or U13523 (N_13523,N_6865,N_7010);
or U13524 (N_13524,N_9372,N_9644);
nand U13525 (N_13525,N_6001,N_7381);
nor U13526 (N_13526,N_7015,N_9328);
xnor U13527 (N_13527,N_6402,N_5245);
nor U13528 (N_13528,N_8092,N_6187);
or U13529 (N_13529,N_5465,N_5640);
xnor U13530 (N_13530,N_7604,N_8568);
xor U13531 (N_13531,N_7992,N_6525);
nand U13532 (N_13532,N_6615,N_5430);
and U13533 (N_13533,N_6480,N_7000);
nor U13534 (N_13534,N_7932,N_8020);
nor U13535 (N_13535,N_7516,N_7132);
or U13536 (N_13536,N_6978,N_8302);
nor U13537 (N_13537,N_8612,N_5590);
and U13538 (N_13538,N_5513,N_5942);
nand U13539 (N_13539,N_5570,N_6636);
nand U13540 (N_13540,N_7393,N_5840);
xor U13541 (N_13541,N_5380,N_7926);
or U13542 (N_13542,N_5163,N_5808);
xnor U13543 (N_13543,N_6992,N_7591);
and U13544 (N_13544,N_9699,N_7571);
and U13545 (N_13545,N_6184,N_9499);
xnor U13546 (N_13546,N_9601,N_9443);
nand U13547 (N_13547,N_8538,N_6800);
xor U13548 (N_13548,N_6777,N_6435);
xor U13549 (N_13549,N_8771,N_8471);
xnor U13550 (N_13550,N_9629,N_6508);
and U13551 (N_13551,N_9038,N_6088);
xnor U13552 (N_13552,N_8824,N_9364);
and U13553 (N_13553,N_8277,N_5838);
nand U13554 (N_13554,N_9097,N_6255);
or U13555 (N_13555,N_6647,N_6220);
xnor U13556 (N_13556,N_9701,N_5813);
nor U13557 (N_13557,N_6354,N_9821);
and U13558 (N_13558,N_8519,N_5544);
nor U13559 (N_13559,N_9003,N_6917);
or U13560 (N_13560,N_6512,N_5641);
or U13561 (N_13561,N_6461,N_8146);
nand U13562 (N_13562,N_7468,N_5159);
nor U13563 (N_13563,N_8550,N_7000);
nand U13564 (N_13564,N_6900,N_8246);
nor U13565 (N_13565,N_6962,N_8317);
xor U13566 (N_13566,N_9976,N_9128);
or U13567 (N_13567,N_6015,N_9274);
nand U13568 (N_13568,N_6930,N_9884);
xnor U13569 (N_13569,N_6131,N_7796);
nand U13570 (N_13570,N_9341,N_5771);
nor U13571 (N_13571,N_5302,N_9972);
xnor U13572 (N_13572,N_7429,N_6158);
and U13573 (N_13573,N_9909,N_8972);
and U13574 (N_13574,N_6000,N_9089);
xnor U13575 (N_13575,N_5370,N_7935);
and U13576 (N_13576,N_7700,N_5452);
xnor U13577 (N_13577,N_9550,N_8229);
xnor U13578 (N_13578,N_8072,N_8127);
nor U13579 (N_13579,N_6626,N_9201);
or U13580 (N_13580,N_8486,N_5192);
and U13581 (N_13581,N_5290,N_6315);
xor U13582 (N_13582,N_6361,N_6992);
nand U13583 (N_13583,N_7790,N_8470);
xnor U13584 (N_13584,N_9218,N_7968);
xnor U13585 (N_13585,N_6235,N_9039);
xnor U13586 (N_13586,N_6477,N_9538);
xor U13587 (N_13587,N_6375,N_8864);
xor U13588 (N_13588,N_6670,N_5329);
xor U13589 (N_13589,N_9865,N_7713);
nor U13590 (N_13590,N_9991,N_6867);
nor U13591 (N_13591,N_9902,N_5409);
xnor U13592 (N_13592,N_5575,N_9911);
nor U13593 (N_13593,N_6401,N_8215);
and U13594 (N_13594,N_9210,N_8811);
nor U13595 (N_13595,N_9739,N_6454);
xnor U13596 (N_13596,N_7065,N_6214);
nand U13597 (N_13597,N_6003,N_9138);
and U13598 (N_13598,N_5747,N_9637);
nor U13599 (N_13599,N_8341,N_5722);
nor U13600 (N_13600,N_5513,N_8529);
xnor U13601 (N_13601,N_7928,N_7545);
xor U13602 (N_13602,N_9999,N_7422);
nor U13603 (N_13603,N_9196,N_8253);
and U13604 (N_13604,N_6975,N_9655);
nor U13605 (N_13605,N_6305,N_5627);
xor U13606 (N_13606,N_8847,N_9307);
nor U13607 (N_13607,N_6007,N_9420);
or U13608 (N_13608,N_5005,N_9448);
nor U13609 (N_13609,N_7923,N_6752);
or U13610 (N_13610,N_8473,N_9393);
and U13611 (N_13611,N_7036,N_7149);
nand U13612 (N_13612,N_7188,N_9397);
or U13613 (N_13613,N_6057,N_7025);
and U13614 (N_13614,N_8812,N_9986);
nor U13615 (N_13615,N_8676,N_6201);
nor U13616 (N_13616,N_5578,N_6944);
and U13617 (N_13617,N_6425,N_6598);
or U13618 (N_13618,N_8607,N_9911);
xnor U13619 (N_13619,N_6952,N_6021);
nand U13620 (N_13620,N_9776,N_9981);
or U13621 (N_13621,N_7023,N_9707);
or U13622 (N_13622,N_9798,N_8186);
nor U13623 (N_13623,N_8526,N_5084);
xnor U13624 (N_13624,N_7092,N_6564);
or U13625 (N_13625,N_7241,N_6258);
xor U13626 (N_13626,N_9393,N_8528);
nand U13627 (N_13627,N_6003,N_5637);
nand U13628 (N_13628,N_5299,N_5997);
nand U13629 (N_13629,N_7085,N_8018);
nand U13630 (N_13630,N_5273,N_9415);
and U13631 (N_13631,N_7574,N_7425);
or U13632 (N_13632,N_9908,N_6008);
nor U13633 (N_13633,N_7033,N_9544);
nand U13634 (N_13634,N_9470,N_8064);
or U13635 (N_13635,N_9711,N_6110);
nor U13636 (N_13636,N_5697,N_5259);
and U13637 (N_13637,N_6064,N_7005);
nand U13638 (N_13638,N_8168,N_7725);
nor U13639 (N_13639,N_5039,N_5251);
and U13640 (N_13640,N_9954,N_8815);
and U13641 (N_13641,N_8712,N_6818);
and U13642 (N_13642,N_6700,N_9180);
xor U13643 (N_13643,N_5966,N_7628);
or U13644 (N_13644,N_6263,N_9484);
nor U13645 (N_13645,N_5225,N_6021);
and U13646 (N_13646,N_9010,N_7445);
nor U13647 (N_13647,N_7797,N_7931);
and U13648 (N_13648,N_8813,N_9329);
or U13649 (N_13649,N_9925,N_7564);
nand U13650 (N_13650,N_7918,N_8000);
nor U13651 (N_13651,N_6296,N_7386);
nand U13652 (N_13652,N_9598,N_7033);
nand U13653 (N_13653,N_9319,N_5009);
nand U13654 (N_13654,N_5625,N_9868);
xor U13655 (N_13655,N_8239,N_9808);
and U13656 (N_13656,N_8168,N_5943);
nand U13657 (N_13657,N_8046,N_9005);
and U13658 (N_13658,N_7337,N_6169);
xnor U13659 (N_13659,N_8860,N_9752);
xnor U13660 (N_13660,N_9822,N_7153);
nor U13661 (N_13661,N_7614,N_8400);
nor U13662 (N_13662,N_8760,N_7662);
and U13663 (N_13663,N_8097,N_9423);
nor U13664 (N_13664,N_7883,N_7096);
nor U13665 (N_13665,N_7373,N_6645);
nor U13666 (N_13666,N_9831,N_9318);
or U13667 (N_13667,N_6882,N_7420);
nor U13668 (N_13668,N_6563,N_7743);
xor U13669 (N_13669,N_9521,N_7706);
xor U13670 (N_13670,N_8764,N_6661);
xor U13671 (N_13671,N_6934,N_7997);
nand U13672 (N_13672,N_9858,N_8364);
nand U13673 (N_13673,N_8782,N_5216);
nand U13674 (N_13674,N_6603,N_5794);
xor U13675 (N_13675,N_6125,N_6248);
xnor U13676 (N_13676,N_8825,N_9957);
xnor U13677 (N_13677,N_9390,N_5985);
xor U13678 (N_13678,N_7275,N_7939);
nand U13679 (N_13679,N_7977,N_9354);
and U13680 (N_13680,N_7708,N_6221);
or U13681 (N_13681,N_7079,N_8267);
and U13682 (N_13682,N_6428,N_9438);
xnor U13683 (N_13683,N_5297,N_7417);
nand U13684 (N_13684,N_6536,N_7921);
and U13685 (N_13685,N_8385,N_8007);
nor U13686 (N_13686,N_6372,N_9851);
and U13687 (N_13687,N_5227,N_8869);
xor U13688 (N_13688,N_5487,N_6869);
xor U13689 (N_13689,N_7103,N_6153);
nand U13690 (N_13690,N_5534,N_8804);
and U13691 (N_13691,N_7970,N_9400);
xor U13692 (N_13692,N_9202,N_7517);
nor U13693 (N_13693,N_7539,N_7476);
or U13694 (N_13694,N_9614,N_6362);
nor U13695 (N_13695,N_9848,N_8880);
nor U13696 (N_13696,N_7519,N_9639);
xnor U13697 (N_13697,N_6627,N_7488);
nand U13698 (N_13698,N_6446,N_9061);
or U13699 (N_13699,N_8958,N_8911);
nand U13700 (N_13700,N_9118,N_7170);
and U13701 (N_13701,N_8557,N_6175);
nand U13702 (N_13702,N_6666,N_9876);
nor U13703 (N_13703,N_6911,N_6190);
or U13704 (N_13704,N_6034,N_7473);
xor U13705 (N_13705,N_7311,N_6480);
xnor U13706 (N_13706,N_9859,N_9361);
nand U13707 (N_13707,N_9131,N_7252);
nor U13708 (N_13708,N_6456,N_9389);
or U13709 (N_13709,N_6194,N_6617);
nand U13710 (N_13710,N_5367,N_8109);
nand U13711 (N_13711,N_9729,N_8944);
xor U13712 (N_13712,N_5737,N_6299);
or U13713 (N_13713,N_7241,N_8660);
and U13714 (N_13714,N_7841,N_8767);
xnor U13715 (N_13715,N_5229,N_6116);
xnor U13716 (N_13716,N_8069,N_9224);
and U13717 (N_13717,N_6887,N_5698);
xnor U13718 (N_13718,N_6744,N_5876);
nand U13719 (N_13719,N_7505,N_9634);
nand U13720 (N_13720,N_6617,N_8108);
nand U13721 (N_13721,N_9312,N_9976);
xor U13722 (N_13722,N_6410,N_6289);
or U13723 (N_13723,N_6867,N_5842);
or U13724 (N_13724,N_9922,N_6929);
xor U13725 (N_13725,N_8050,N_9850);
xnor U13726 (N_13726,N_9225,N_5090);
and U13727 (N_13727,N_8122,N_7491);
or U13728 (N_13728,N_6897,N_6501);
and U13729 (N_13729,N_7546,N_8744);
nand U13730 (N_13730,N_5999,N_6642);
or U13731 (N_13731,N_6726,N_6335);
nand U13732 (N_13732,N_9607,N_8597);
nand U13733 (N_13733,N_9267,N_6959);
xor U13734 (N_13734,N_8542,N_8279);
nor U13735 (N_13735,N_9504,N_8649);
or U13736 (N_13736,N_5337,N_7396);
nand U13737 (N_13737,N_8246,N_5698);
nor U13738 (N_13738,N_6148,N_9046);
or U13739 (N_13739,N_7280,N_9200);
nand U13740 (N_13740,N_9336,N_7095);
or U13741 (N_13741,N_9368,N_8867);
xor U13742 (N_13742,N_5037,N_6530);
and U13743 (N_13743,N_6572,N_9171);
nor U13744 (N_13744,N_7006,N_9828);
xnor U13745 (N_13745,N_5487,N_5690);
nand U13746 (N_13746,N_5565,N_6572);
and U13747 (N_13747,N_7499,N_9567);
nand U13748 (N_13748,N_9286,N_6417);
nand U13749 (N_13749,N_6362,N_7587);
xnor U13750 (N_13750,N_8145,N_9427);
xor U13751 (N_13751,N_6614,N_9547);
nor U13752 (N_13752,N_9825,N_9941);
or U13753 (N_13753,N_6925,N_7804);
xnor U13754 (N_13754,N_7218,N_5530);
xor U13755 (N_13755,N_5850,N_9432);
and U13756 (N_13756,N_9010,N_9400);
nor U13757 (N_13757,N_5513,N_6115);
nand U13758 (N_13758,N_5157,N_6904);
nand U13759 (N_13759,N_6031,N_8291);
nor U13760 (N_13760,N_5261,N_5109);
or U13761 (N_13761,N_5099,N_8931);
nor U13762 (N_13762,N_5144,N_7531);
xnor U13763 (N_13763,N_7129,N_9217);
or U13764 (N_13764,N_8881,N_8113);
nor U13765 (N_13765,N_6231,N_6211);
nor U13766 (N_13766,N_5038,N_6102);
and U13767 (N_13767,N_9914,N_6556);
xnor U13768 (N_13768,N_8307,N_5152);
xnor U13769 (N_13769,N_8747,N_5962);
xor U13770 (N_13770,N_9908,N_9915);
nand U13771 (N_13771,N_6850,N_9040);
or U13772 (N_13772,N_9323,N_8447);
xnor U13773 (N_13773,N_5019,N_9583);
and U13774 (N_13774,N_7805,N_8037);
and U13775 (N_13775,N_8592,N_9593);
or U13776 (N_13776,N_9590,N_8678);
xnor U13777 (N_13777,N_5627,N_5877);
and U13778 (N_13778,N_8323,N_9394);
and U13779 (N_13779,N_8286,N_8453);
xnor U13780 (N_13780,N_7749,N_9026);
or U13781 (N_13781,N_8151,N_6575);
xor U13782 (N_13782,N_7855,N_9716);
nand U13783 (N_13783,N_6953,N_8700);
nor U13784 (N_13784,N_6190,N_6446);
xor U13785 (N_13785,N_9345,N_7212);
and U13786 (N_13786,N_7747,N_7971);
xor U13787 (N_13787,N_7616,N_6978);
xor U13788 (N_13788,N_8519,N_5838);
xnor U13789 (N_13789,N_9896,N_9492);
or U13790 (N_13790,N_8856,N_9789);
nor U13791 (N_13791,N_9620,N_9823);
nand U13792 (N_13792,N_8209,N_6243);
nor U13793 (N_13793,N_5890,N_6183);
nand U13794 (N_13794,N_5114,N_5364);
or U13795 (N_13795,N_6075,N_6567);
nand U13796 (N_13796,N_6333,N_8894);
nor U13797 (N_13797,N_7094,N_8975);
nor U13798 (N_13798,N_8262,N_5881);
xnor U13799 (N_13799,N_8722,N_6356);
nand U13800 (N_13800,N_6851,N_7690);
nor U13801 (N_13801,N_8743,N_7262);
nand U13802 (N_13802,N_6878,N_7401);
xnor U13803 (N_13803,N_6082,N_5823);
nand U13804 (N_13804,N_7400,N_9647);
and U13805 (N_13805,N_7328,N_6844);
xnor U13806 (N_13806,N_7117,N_9783);
nand U13807 (N_13807,N_5853,N_6439);
xor U13808 (N_13808,N_6052,N_7036);
or U13809 (N_13809,N_8952,N_9012);
xor U13810 (N_13810,N_6673,N_9224);
xor U13811 (N_13811,N_9830,N_5910);
nand U13812 (N_13812,N_9144,N_7030);
nand U13813 (N_13813,N_7875,N_5341);
nor U13814 (N_13814,N_5643,N_5999);
nand U13815 (N_13815,N_8635,N_9311);
and U13816 (N_13816,N_8184,N_7263);
xnor U13817 (N_13817,N_6214,N_7320);
xnor U13818 (N_13818,N_8174,N_9912);
nor U13819 (N_13819,N_5320,N_7011);
nor U13820 (N_13820,N_6154,N_8037);
and U13821 (N_13821,N_5886,N_7053);
nand U13822 (N_13822,N_7610,N_6298);
nor U13823 (N_13823,N_6441,N_6802);
nor U13824 (N_13824,N_7571,N_9430);
nand U13825 (N_13825,N_8402,N_7243);
nand U13826 (N_13826,N_6172,N_5654);
or U13827 (N_13827,N_8557,N_9626);
nor U13828 (N_13828,N_5025,N_6966);
xor U13829 (N_13829,N_9339,N_9785);
and U13830 (N_13830,N_7267,N_9202);
and U13831 (N_13831,N_8167,N_8977);
or U13832 (N_13832,N_7058,N_9250);
xor U13833 (N_13833,N_5953,N_7543);
xor U13834 (N_13834,N_7432,N_8848);
xnor U13835 (N_13835,N_6347,N_9205);
and U13836 (N_13836,N_5204,N_8333);
nor U13837 (N_13837,N_6702,N_5490);
or U13838 (N_13838,N_5093,N_7734);
xnor U13839 (N_13839,N_5766,N_6677);
nand U13840 (N_13840,N_5469,N_9094);
and U13841 (N_13841,N_9180,N_5786);
xor U13842 (N_13842,N_9921,N_7767);
and U13843 (N_13843,N_8669,N_8401);
or U13844 (N_13844,N_6104,N_8583);
or U13845 (N_13845,N_6930,N_7972);
nor U13846 (N_13846,N_9221,N_7659);
xnor U13847 (N_13847,N_7696,N_8504);
nor U13848 (N_13848,N_6109,N_9734);
and U13849 (N_13849,N_5027,N_7249);
and U13850 (N_13850,N_7267,N_5274);
or U13851 (N_13851,N_6424,N_8998);
nor U13852 (N_13852,N_9834,N_9205);
xor U13853 (N_13853,N_8011,N_8106);
xor U13854 (N_13854,N_6980,N_6207);
nor U13855 (N_13855,N_6488,N_7056);
or U13856 (N_13856,N_8612,N_8346);
xnor U13857 (N_13857,N_7813,N_9282);
xnor U13858 (N_13858,N_8899,N_9371);
xor U13859 (N_13859,N_5111,N_6496);
nand U13860 (N_13860,N_5581,N_7268);
xor U13861 (N_13861,N_7097,N_9068);
and U13862 (N_13862,N_6394,N_8658);
and U13863 (N_13863,N_8840,N_8646);
nor U13864 (N_13864,N_6904,N_7960);
nand U13865 (N_13865,N_9353,N_7749);
or U13866 (N_13866,N_5569,N_9566);
nor U13867 (N_13867,N_9786,N_8314);
or U13868 (N_13868,N_8299,N_9755);
xnor U13869 (N_13869,N_7620,N_6240);
nor U13870 (N_13870,N_5368,N_8512);
and U13871 (N_13871,N_6843,N_6472);
nand U13872 (N_13872,N_7661,N_6282);
or U13873 (N_13873,N_6794,N_6110);
or U13874 (N_13874,N_8861,N_9266);
or U13875 (N_13875,N_6073,N_8388);
xor U13876 (N_13876,N_8422,N_9738);
xnor U13877 (N_13877,N_5431,N_9667);
nand U13878 (N_13878,N_7831,N_7144);
or U13879 (N_13879,N_9305,N_5756);
xnor U13880 (N_13880,N_5448,N_9871);
and U13881 (N_13881,N_5624,N_9448);
nor U13882 (N_13882,N_9336,N_5847);
xnor U13883 (N_13883,N_6473,N_7527);
nor U13884 (N_13884,N_6016,N_8590);
nand U13885 (N_13885,N_9778,N_8903);
and U13886 (N_13886,N_5691,N_9628);
and U13887 (N_13887,N_6613,N_6959);
and U13888 (N_13888,N_5598,N_5397);
and U13889 (N_13889,N_7005,N_7185);
or U13890 (N_13890,N_8461,N_8405);
nor U13891 (N_13891,N_8709,N_7733);
xnor U13892 (N_13892,N_8234,N_6061);
nor U13893 (N_13893,N_9055,N_8610);
or U13894 (N_13894,N_9897,N_6855);
xnor U13895 (N_13895,N_9435,N_8836);
and U13896 (N_13896,N_7917,N_6862);
xor U13897 (N_13897,N_5881,N_9261);
xnor U13898 (N_13898,N_8609,N_5526);
nand U13899 (N_13899,N_9677,N_8586);
xnor U13900 (N_13900,N_7698,N_9720);
nor U13901 (N_13901,N_8760,N_9577);
xor U13902 (N_13902,N_7766,N_7931);
xnor U13903 (N_13903,N_5877,N_5057);
nor U13904 (N_13904,N_8359,N_6145);
or U13905 (N_13905,N_8102,N_5340);
and U13906 (N_13906,N_7857,N_7186);
xor U13907 (N_13907,N_7203,N_6830);
or U13908 (N_13908,N_5997,N_9774);
or U13909 (N_13909,N_6143,N_9302);
and U13910 (N_13910,N_8160,N_6470);
and U13911 (N_13911,N_6948,N_5722);
nand U13912 (N_13912,N_9430,N_8695);
xor U13913 (N_13913,N_8503,N_5157);
xnor U13914 (N_13914,N_6304,N_5436);
and U13915 (N_13915,N_5752,N_7433);
nand U13916 (N_13916,N_8742,N_5219);
xor U13917 (N_13917,N_9310,N_8439);
nor U13918 (N_13918,N_9990,N_5005);
and U13919 (N_13919,N_7954,N_9241);
and U13920 (N_13920,N_8413,N_9212);
nor U13921 (N_13921,N_9576,N_6627);
nor U13922 (N_13922,N_6818,N_7683);
nor U13923 (N_13923,N_7076,N_8283);
and U13924 (N_13924,N_8724,N_6834);
and U13925 (N_13925,N_7950,N_5813);
xnor U13926 (N_13926,N_6350,N_5054);
and U13927 (N_13927,N_7373,N_7563);
xor U13928 (N_13928,N_9752,N_5471);
or U13929 (N_13929,N_6641,N_6150);
and U13930 (N_13930,N_7523,N_5307);
nor U13931 (N_13931,N_8674,N_9240);
nand U13932 (N_13932,N_5351,N_5645);
or U13933 (N_13933,N_8166,N_8792);
and U13934 (N_13934,N_8949,N_7101);
nand U13935 (N_13935,N_9041,N_5738);
nand U13936 (N_13936,N_5867,N_5172);
or U13937 (N_13937,N_6901,N_8347);
nor U13938 (N_13938,N_5536,N_9995);
xor U13939 (N_13939,N_5809,N_8280);
nor U13940 (N_13940,N_9525,N_9676);
nor U13941 (N_13941,N_5446,N_7915);
and U13942 (N_13942,N_5904,N_5267);
nand U13943 (N_13943,N_9218,N_7794);
xnor U13944 (N_13944,N_5075,N_7710);
xnor U13945 (N_13945,N_5073,N_6995);
and U13946 (N_13946,N_6261,N_5167);
nor U13947 (N_13947,N_8019,N_8533);
and U13948 (N_13948,N_8360,N_6576);
or U13949 (N_13949,N_8752,N_7223);
or U13950 (N_13950,N_8902,N_6442);
or U13951 (N_13951,N_9906,N_7051);
or U13952 (N_13952,N_8460,N_8781);
nand U13953 (N_13953,N_7549,N_9696);
nor U13954 (N_13954,N_6415,N_8756);
or U13955 (N_13955,N_9822,N_5805);
xor U13956 (N_13956,N_5460,N_5514);
nor U13957 (N_13957,N_9810,N_6305);
xor U13958 (N_13958,N_5614,N_9198);
xnor U13959 (N_13959,N_8323,N_9072);
xnor U13960 (N_13960,N_7221,N_5372);
and U13961 (N_13961,N_5537,N_5704);
nor U13962 (N_13962,N_5785,N_8297);
or U13963 (N_13963,N_6460,N_8187);
xor U13964 (N_13964,N_9859,N_9948);
and U13965 (N_13965,N_5588,N_9776);
xor U13966 (N_13966,N_5661,N_8575);
nor U13967 (N_13967,N_5395,N_8259);
or U13968 (N_13968,N_5523,N_5725);
nor U13969 (N_13969,N_9912,N_7328);
and U13970 (N_13970,N_6569,N_6562);
xor U13971 (N_13971,N_9939,N_5075);
or U13972 (N_13972,N_5051,N_8781);
xnor U13973 (N_13973,N_9946,N_6142);
and U13974 (N_13974,N_8631,N_5358);
nand U13975 (N_13975,N_6922,N_5827);
nor U13976 (N_13976,N_8899,N_7621);
nor U13977 (N_13977,N_8373,N_7353);
nand U13978 (N_13978,N_7233,N_6687);
xnor U13979 (N_13979,N_9094,N_6983);
xnor U13980 (N_13980,N_7233,N_7517);
and U13981 (N_13981,N_7982,N_5912);
xor U13982 (N_13982,N_9083,N_6828);
nor U13983 (N_13983,N_7739,N_8443);
or U13984 (N_13984,N_7590,N_7891);
nor U13985 (N_13985,N_6489,N_9607);
or U13986 (N_13986,N_8355,N_9988);
nor U13987 (N_13987,N_5842,N_8721);
and U13988 (N_13988,N_9442,N_8116);
nor U13989 (N_13989,N_6777,N_7017);
or U13990 (N_13990,N_6966,N_6450);
nand U13991 (N_13991,N_7886,N_6319);
and U13992 (N_13992,N_6675,N_9832);
and U13993 (N_13993,N_7369,N_7623);
nand U13994 (N_13994,N_6914,N_5265);
xor U13995 (N_13995,N_5047,N_9276);
or U13996 (N_13996,N_6545,N_6604);
or U13997 (N_13997,N_8559,N_5185);
xnor U13998 (N_13998,N_5307,N_8043);
nor U13999 (N_13999,N_8999,N_9264);
xnor U14000 (N_14000,N_7022,N_6827);
and U14001 (N_14001,N_7680,N_6463);
nand U14002 (N_14002,N_7303,N_7436);
and U14003 (N_14003,N_6059,N_7335);
nand U14004 (N_14004,N_8025,N_9582);
and U14005 (N_14005,N_7689,N_9342);
and U14006 (N_14006,N_8202,N_5617);
nand U14007 (N_14007,N_9913,N_7569);
and U14008 (N_14008,N_5454,N_8404);
xnor U14009 (N_14009,N_6716,N_8669);
nor U14010 (N_14010,N_8715,N_7812);
or U14011 (N_14011,N_9529,N_5308);
xor U14012 (N_14012,N_9849,N_9506);
or U14013 (N_14013,N_9235,N_9243);
or U14014 (N_14014,N_8439,N_5981);
xor U14015 (N_14015,N_7643,N_9486);
or U14016 (N_14016,N_6594,N_9759);
or U14017 (N_14017,N_7991,N_8404);
nand U14018 (N_14018,N_8708,N_8533);
or U14019 (N_14019,N_5194,N_9096);
or U14020 (N_14020,N_6733,N_6116);
nor U14021 (N_14021,N_9082,N_6780);
nand U14022 (N_14022,N_6655,N_9672);
or U14023 (N_14023,N_6276,N_7801);
xor U14024 (N_14024,N_9757,N_8696);
or U14025 (N_14025,N_9546,N_7945);
and U14026 (N_14026,N_7628,N_8231);
and U14027 (N_14027,N_5942,N_7787);
or U14028 (N_14028,N_6974,N_7533);
xor U14029 (N_14029,N_5958,N_5271);
xnor U14030 (N_14030,N_5960,N_8464);
xor U14031 (N_14031,N_6091,N_9641);
nor U14032 (N_14032,N_5042,N_9112);
nand U14033 (N_14033,N_7503,N_7456);
and U14034 (N_14034,N_6246,N_9817);
or U14035 (N_14035,N_5694,N_9101);
or U14036 (N_14036,N_5616,N_8965);
and U14037 (N_14037,N_6762,N_6026);
and U14038 (N_14038,N_8210,N_9309);
and U14039 (N_14039,N_8550,N_9510);
nand U14040 (N_14040,N_6867,N_7321);
nor U14041 (N_14041,N_7711,N_6137);
nand U14042 (N_14042,N_5648,N_6963);
and U14043 (N_14043,N_9833,N_6505);
or U14044 (N_14044,N_8464,N_9550);
or U14045 (N_14045,N_9850,N_6825);
or U14046 (N_14046,N_6295,N_6497);
nand U14047 (N_14047,N_7745,N_7551);
or U14048 (N_14048,N_8921,N_7934);
nor U14049 (N_14049,N_6960,N_8135);
and U14050 (N_14050,N_7236,N_5570);
xor U14051 (N_14051,N_6054,N_5000);
and U14052 (N_14052,N_6574,N_6629);
and U14053 (N_14053,N_5508,N_9789);
and U14054 (N_14054,N_6281,N_8259);
xnor U14055 (N_14055,N_8230,N_6204);
xor U14056 (N_14056,N_8773,N_6724);
xnor U14057 (N_14057,N_7998,N_7996);
nand U14058 (N_14058,N_6678,N_6233);
nand U14059 (N_14059,N_6207,N_9740);
xnor U14060 (N_14060,N_5812,N_9335);
and U14061 (N_14061,N_7132,N_9628);
or U14062 (N_14062,N_9141,N_7156);
and U14063 (N_14063,N_8912,N_5994);
and U14064 (N_14064,N_8977,N_8759);
and U14065 (N_14065,N_9614,N_5171);
and U14066 (N_14066,N_8050,N_5755);
and U14067 (N_14067,N_8259,N_5889);
and U14068 (N_14068,N_9736,N_5861);
xnor U14069 (N_14069,N_7887,N_8716);
or U14070 (N_14070,N_5426,N_5259);
xor U14071 (N_14071,N_5701,N_7568);
nand U14072 (N_14072,N_8891,N_7331);
xnor U14073 (N_14073,N_6236,N_8299);
and U14074 (N_14074,N_6748,N_9313);
nand U14075 (N_14075,N_8494,N_8082);
or U14076 (N_14076,N_5619,N_7108);
or U14077 (N_14077,N_5293,N_5861);
nand U14078 (N_14078,N_5325,N_9135);
and U14079 (N_14079,N_6223,N_8500);
nand U14080 (N_14080,N_9538,N_9387);
or U14081 (N_14081,N_9356,N_8285);
nor U14082 (N_14082,N_6342,N_6738);
xnor U14083 (N_14083,N_6005,N_7304);
nand U14084 (N_14084,N_9140,N_5341);
xnor U14085 (N_14085,N_9958,N_9754);
or U14086 (N_14086,N_6393,N_6412);
and U14087 (N_14087,N_7775,N_8057);
nor U14088 (N_14088,N_8642,N_9201);
xor U14089 (N_14089,N_9243,N_8273);
nand U14090 (N_14090,N_9982,N_8365);
nor U14091 (N_14091,N_5531,N_7548);
or U14092 (N_14092,N_6607,N_7193);
nand U14093 (N_14093,N_7287,N_9927);
or U14094 (N_14094,N_7880,N_7572);
nand U14095 (N_14095,N_7676,N_5167);
nor U14096 (N_14096,N_7328,N_6634);
xor U14097 (N_14097,N_7423,N_8075);
or U14098 (N_14098,N_8233,N_7968);
nand U14099 (N_14099,N_8732,N_9020);
xor U14100 (N_14100,N_5558,N_8587);
nand U14101 (N_14101,N_5774,N_6917);
nor U14102 (N_14102,N_7807,N_7164);
nand U14103 (N_14103,N_8179,N_6073);
and U14104 (N_14104,N_6779,N_6407);
nand U14105 (N_14105,N_5745,N_9165);
nor U14106 (N_14106,N_9497,N_6882);
and U14107 (N_14107,N_9683,N_5805);
xnor U14108 (N_14108,N_7500,N_7686);
xor U14109 (N_14109,N_5530,N_8198);
and U14110 (N_14110,N_8970,N_5155);
nand U14111 (N_14111,N_7460,N_6602);
or U14112 (N_14112,N_9799,N_8465);
nor U14113 (N_14113,N_6069,N_9515);
nor U14114 (N_14114,N_8347,N_5395);
xnor U14115 (N_14115,N_6289,N_5721);
and U14116 (N_14116,N_5473,N_5166);
or U14117 (N_14117,N_5130,N_9266);
or U14118 (N_14118,N_8261,N_7920);
or U14119 (N_14119,N_5408,N_7055);
and U14120 (N_14120,N_8918,N_5489);
nand U14121 (N_14121,N_6493,N_5849);
and U14122 (N_14122,N_9806,N_7633);
or U14123 (N_14123,N_8727,N_6822);
nand U14124 (N_14124,N_7398,N_8557);
xor U14125 (N_14125,N_7638,N_6990);
nand U14126 (N_14126,N_9163,N_7121);
nand U14127 (N_14127,N_9344,N_7002);
nor U14128 (N_14128,N_8934,N_5202);
or U14129 (N_14129,N_6277,N_5717);
nor U14130 (N_14130,N_5957,N_6533);
xnor U14131 (N_14131,N_7463,N_7010);
xor U14132 (N_14132,N_6907,N_9066);
nand U14133 (N_14133,N_7957,N_9490);
nor U14134 (N_14134,N_7151,N_5265);
nor U14135 (N_14135,N_8805,N_5800);
or U14136 (N_14136,N_9706,N_7494);
and U14137 (N_14137,N_9873,N_9857);
nand U14138 (N_14138,N_6284,N_7109);
and U14139 (N_14139,N_7360,N_5934);
nor U14140 (N_14140,N_9933,N_9622);
nand U14141 (N_14141,N_6689,N_9390);
nand U14142 (N_14142,N_8995,N_8371);
xnor U14143 (N_14143,N_7991,N_9788);
nand U14144 (N_14144,N_5640,N_7880);
or U14145 (N_14145,N_7737,N_7946);
and U14146 (N_14146,N_7077,N_5846);
and U14147 (N_14147,N_5306,N_9472);
and U14148 (N_14148,N_5478,N_8555);
and U14149 (N_14149,N_5921,N_9082);
xor U14150 (N_14150,N_6230,N_5206);
nand U14151 (N_14151,N_7690,N_7580);
xor U14152 (N_14152,N_9949,N_8969);
nand U14153 (N_14153,N_6682,N_5469);
or U14154 (N_14154,N_6514,N_5324);
nor U14155 (N_14155,N_6930,N_5922);
or U14156 (N_14156,N_5911,N_9294);
xor U14157 (N_14157,N_7586,N_9184);
nand U14158 (N_14158,N_9278,N_8267);
xor U14159 (N_14159,N_9058,N_7909);
and U14160 (N_14160,N_7150,N_8975);
nor U14161 (N_14161,N_5865,N_6757);
xnor U14162 (N_14162,N_9874,N_9365);
nor U14163 (N_14163,N_8210,N_5791);
nor U14164 (N_14164,N_8422,N_7498);
and U14165 (N_14165,N_5713,N_8146);
nand U14166 (N_14166,N_9844,N_8242);
nand U14167 (N_14167,N_5355,N_6183);
or U14168 (N_14168,N_7795,N_6427);
xor U14169 (N_14169,N_8323,N_7226);
or U14170 (N_14170,N_7934,N_7708);
nand U14171 (N_14171,N_9453,N_7072);
nand U14172 (N_14172,N_5499,N_8857);
nor U14173 (N_14173,N_8343,N_6210);
xnor U14174 (N_14174,N_9117,N_5633);
nor U14175 (N_14175,N_5270,N_6815);
or U14176 (N_14176,N_9849,N_6023);
and U14177 (N_14177,N_9477,N_8526);
nand U14178 (N_14178,N_9177,N_7180);
and U14179 (N_14179,N_7145,N_9924);
nor U14180 (N_14180,N_6496,N_7126);
nand U14181 (N_14181,N_9078,N_8414);
or U14182 (N_14182,N_7134,N_6007);
xnor U14183 (N_14183,N_8483,N_6593);
nor U14184 (N_14184,N_9159,N_9160);
nand U14185 (N_14185,N_6029,N_7272);
xnor U14186 (N_14186,N_6826,N_9181);
and U14187 (N_14187,N_6397,N_7877);
xor U14188 (N_14188,N_5884,N_7344);
or U14189 (N_14189,N_5131,N_9296);
xor U14190 (N_14190,N_7616,N_6939);
xor U14191 (N_14191,N_5842,N_7367);
and U14192 (N_14192,N_6709,N_8807);
nor U14193 (N_14193,N_5992,N_7721);
and U14194 (N_14194,N_7721,N_7990);
or U14195 (N_14195,N_8399,N_5730);
nor U14196 (N_14196,N_5728,N_7258);
or U14197 (N_14197,N_8726,N_6530);
nor U14198 (N_14198,N_6580,N_9705);
xor U14199 (N_14199,N_7395,N_9721);
and U14200 (N_14200,N_8494,N_5680);
or U14201 (N_14201,N_5318,N_8783);
and U14202 (N_14202,N_8649,N_7424);
or U14203 (N_14203,N_6191,N_5683);
nand U14204 (N_14204,N_9025,N_5718);
xor U14205 (N_14205,N_6404,N_8121);
nor U14206 (N_14206,N_6138,N_9832);
nand U14207 (N_14207,N_6147,N_5901);
nand U14208 (N_14208,N_5869,N_8528);
nor U14209 (N_14209,N_7341,N_5330);
nand U14210 (N_14210,N_7493,N_9553);
and U14211 (N_14211,N_7356,N_9501);
or U14212 (N_14212,N_7505,N_8368);
and U14213 (N_14213,N_9886,N_7682);
nor U14214 (N_14214,N_7649,N_7026);
or U14215 (N_14215,N_5125,N_6257);
xnor U14216 (N_14216,N_9777,N_9897);
xnor U14217 (N_14217,N_5351,N_9795);
nor U14218 (N_14218,N_8068,N_7700);
nor U14219 (N_14219,N_9473,N_5014);
nor U14220 (N_14220,N_8532,N_9320);
xor U14221 (N_14221,N_9136,N_6780);
and U14222 (N_14222,N_9291,N_8472);
and U14223 (N_14223,N_9333,N_6830);
and U14224 (N_14224,N_6587,N_6150);
nor U14225 (N_14225,N_5900,N_9527);
and U14226 (N_14226,N_9542,N_7657);
or U14227 (N_14227,N_8114,N_7047);
nor U14228 (N_14228,N_7232,N_5602);
nand U14229 (N_14229,N_5014,N_5755);
nand U14230 (N_14230,N_9638,N_7151);
xnor U14231 (N_14231,N_9719,N_9333);
or U14232 (N_14232,N_7852,N_8002);
and U14233 (N_14233,N_9342,N_9088);
xor U14234 (N_14234,N_7032,N_5956);
nor U14235 (N_14235,N_8984,N_8319);
xnor U14236 (N_14236,N_6750,N_6627);
xnor U14237 (N_14237,N_9186,N_8398);
or U14238 (N_14238,N_9494,N_7888);
or U14239 (N_14239,N_8203,N_7572);
nor U14240 (N_14240,N_7066,N_9004);
nor U14241 (N_14241,N_6642,N_7280);
and U14242 (N_14242,N_5945,N_8521);
xnor U14243 (N_14243,N_6541,N_5170);
xnor U14244 (N_14244,N_7844,N_8781);
nand U14245 (N_14245,N_6232,N_9493);
xor U14246 (N_14246,N_5882,N_7690);
xnor U14247 (N_14247,N_8613,N_8896);
nand U14248 (N_14248,N_7775,N_6963);
nand U14249 (N_14249,N_8089,N_9979);
xor U14250 (N_14250,N_6917,N_9623);
or U14251 (N_14251,N_8911,N_6246);
xnor U14252 (N_14252,N_7626,N_9478);
or U14253 (N_14253,N_5728,N_6586);
or U14254 (N_14254,N_9779,N_8345);
xnor U14255 (N_14255,N_8198,N_8716);
and U14256 (N_14256,N_8729,N_5101);
nor U14257 (N_14257,N_7136,N_9357);
and U14258 (N_14258,N_5173,N_7149);
nor U14259 (N_14259,N_8319,N_8911);
xnor U14260 (N_14260,N_6263,N_6715);
and U14261 (N_14261,N_5310,N_6221);
xor U14262 (N_14262,N_6174,N_9000);
nor U14263 (N_14263,N_8413,N_6612);
nand U14264 (N_14264,N_9451,N_7265);
nand U14265 (N_14265,N_7839,N_6744);
nor U14266 (N_14266,N_8718,N_6952);
xnor U14267 (N_14267,N_9507,N_8030);
nor U14268 (N_14268,N_8590,N_6644);
and U14269 (N_14269,N_6990,N_6681);
or U14270 (N_14270,N_8048,N_8409);
and U14271 (N_14271,N_9768,N_8416);
or U14272 (N_14272,N_7747,N_7373);
xnor U14273 (N_14273,N_5253,N_5777);
and U14274 (N_14274,N_6881,N_8888);
nand U14275 (N_14275,N_8389,N_5918);
and U14276 (N_14276,N_6884,N_6600);
or U14277 (N_14277,N_6498,N_8635);
xor U14278 (N_14278,N_7110,N_7270);
or U14279 (N_14279,N_7448,N_9135);
or U14280 (N_14280,N_9766,N_8957);
or U14281 (N_14281,N_7486,N_6792);
xnor U14282 (N_14282,N_5822,N_9510);
and U14283 (N_14283,N_6484,N_5499);
and U14284 (N_14284,N_7168,N_6164);
or U14285 (N_14285,N_5976,N_6962);
and U14286 (N_14286,N_6692,N_7997);
nor U14287 (N_14287,N_5884,N_6411);
nand U14288 (N_14288,N_6188,N_6253);
xnor U14289 (N_14289,N_6420,N_5885);
nand U14290 (N_14290,N_5809,N_6181);
nor U14291 (N_14291,N_5514,N_6873);
and U14292 (N_14292,N_8382,N_6084);
or U14293 (N_14293,N_5382,N_5340);
or U14294 (N_14294,N_5106,N_6998);
nor U14295 (N_14295,N_9614,N_6406);
nor U14296 (N_14296,N_5562,N_8238);
or U14297 (N_14297,N_6415,N_6599);
nand U14298 (N_14298,N_5124,N_7980);
or U14299 (N_14299,N_9901,N_8433);
and U14300 (N_14300,N_5906,N_6137);
xor U14301 (N_14301,N_9678,N_6624);
nand U14302 (N_14302,N_8059,N_7346);
nor U14303 (N_14303,N_7418,N_6971);
nand U14304 (N_14304,N_7496,N_6562);
xnor U14305 (N_14305,N_6308,N_9501);
and U14306 (N_14306,N_9551,N_5958);
or U14307 (N_14307,N_6685,N_8877);
or U14308 (N_14308,N_8833,N_5491);
nor U14309 (N_14309,N_8848,N_9204);
nor U14310 (N_14310,N_8564,N_7633);
nand U14311 (N_14311,N_5396,N_5404);
nand U14312 (N_14312,N_6180,N_8935);
or U14313 (N_14313,N_9055,N_8335);
xnor U14314 (N_14314,N_7217,N_7645);
or U14315 (N_14315,N_5711,N_6417);
xnor U14316 (N_14316,N_8766,N_5694);
or U14317 (N_14317,N_8875,N_8897);
or U14318 (N_14318,N_5955,N_7676);
nor U14319 (N_14319,N_8718,N_7018);
xnor U14320 (N_14320,N_5211,N_8827);
or U14321 (N_14321,N_8029,N_8474);
xnor U14322 (N_14322,N_9347,N_8374);
or U14323 (N_14323,N_6384,N_9303);
and U14324 (N_14324,N_9758,N_7662);
nor U14325 (N_14325,N_9331,N_9551);
and U14326 (N_14326,N_9908,N_9159);
xnor U14327 (N_14327,N_9878,N_9625);
and U14328 (N_14328,N_7312,N_7185);
xor U14329 (N_14329,N_8200,N_5964);
nand U14330 (N_14330,N_7148,N_5821);
and U14331 (N_14331,N_6163,N_9390);
nor U14332 (N_14332,N_7883,N_5812);
xor U14333 (N_14333,N_8298,N_7263);
nand U14334 (N_14334,N_7895,N_6294);
or U14335 (N_14335,N_8096,N_7823);
or U14336 (N_14336,N_5594,N_8004);
nor U14337 (N_14337,N_8861,N_8063);
nand U14338 (N_14338,N_7847,N_7386);
and U14339 (N_14339,N_6542,N_7817);
nand U14340 (N_14340,N_8874,N_8667);
nor U14341 (N_14341,N_9308,N_5989);
xor U14342 (N_14342,N_6616,N_8038);
xor U14343 (N_14343,N_5287,N_8372);
nor U14344 (N_14344,N_7277,N_6449);
xnor U14345 (N_14345,N_7449,N_7604);
and U14346 (N_14346,N_7979,N_8517);
nand U14347 (N_14347,N_9939,N_5426);
nand U14348 (N_14348,N_6866,N_9219);
nor U14349 (N_14349,N_5460,N_7387);
or U14350 (N_14350,N_7371,N_5795);
xnor U14351 (N_14351,N_6338,N_6781);
nand U14352 (N_14352,N_8797,N_8203);
nor U14353 (N_14353,N_5295,N_9388);
and U14354 (N_14354,N_9556,N_5022);
and U14355 (N_14355,N_5647,N_8527);
nor U14356 (N_14356,N_9633,N_8164);
xnor U14357 (N_14357,N_5673,N_8041);
xnor U14358 (N_14358,N_9993,N_7484);
or U14359 (N_14359,N_7298,N_8009);
nand U14360 (N_14360,N_8331,N_7758);
nor U14361 (N_14361,N_8072,N_7708);
xor U14362 (N_14362,N_8443,N_6615);
or U14363 (N_14363,N_7209,N_6443);
xnor U14364 (N_14364,N_7278,N_5045);
and U14365 (N_14365,N_7039,N_5195);
nor U14366 (N_14366,N_5484,N_9023);
xnor U14367 (N_14367,N_6835,N_7338);
or U14368 (N_14368,N_9301,N_9155);
and U14369 (N_14369,N_9030,N_8250);
or U14370 (N_14370,N_9262,N_9786);
and U14371 (N_14371,N_9370,N_6126);
nor U14372 (N_14372,N_8194,N_7424);
xnor U14373 (N_14373,N_6997,N_5868);
nand U14374 (N_14374,N_5085,N_7471);
nand U14375 (N_14375,N_5982,N_8147);
nor U14376 (N_14376,N_8657,N_5949);
and U14377 (N_14377,N_9470,N_9349);
and U14378 (N_14378,N_7533,N_6708);
or U14379 (N_14379,N_5541,N_6524);
xnor U14380 (N_14380,N_9078,N_5550);
nor U14381 (N_14381,N_7198,N_9423);
and U14382 (N_14382,N_5966,N_7013);
or U14383 (N_14383,N_5928,N_9687);
nand U14384 (N_14384,N_6675,N_6921);
or U14385 (N_14385,N_9588,N_8763);
nand U14386 (N_14386,N_7741,N_5222);
nand U14387 (N_14387,N_8163,N_7829);
xnor U14388 (N_14388,N_9722,N_8062);
and U14389 (N_14389,N_5624,N_9152);
nand U14390 (N_14390,N_5175,N_5477);
nand U14391 (N_14391,N_7416,N_8641);
xor U14392 (N_14392,N_6071,N_8438);
xnor U14393 (N_14393,N_5853,N_6058);
nand U14394 (N_14394,N_5956,N_8693);
xor U14395 (N_14395,N_5909,N_6117);
or U14396 (N_14396,N_8309,N_8794);
nand U14397 (N_14397,N_8324,N_6099);
and U14398 (N_14398,N_6733,N_8498);
nor U14399 (N_14399,N_6263,N_9041);
nor U14400 (N_14400,N_7752,N_9538);
xor U14401 (N_14401,N_6997,N_5316);
nor U14402 (N_14402,N_7578,N_8114);
xnor U14403 (N_14403,N_5440,N_9015);
and U14404 (N_14404,N_5271,N_9885);
nor U14405 (N_14405,N_9044,N_8189);
or U14406 (N_14406,N_7052,N_5363);
and U14407 (N_14407,N_5245,N_6465);
or U14408 (N_14408,N_7715,N_7433);
xnor U14409 (N_14409,N_5911,N_9429);
nand U14410 (N_14410,N_5181,N_8163);
nor U14411 (N_14411,N_7496,N_8928);
nand U14412 (N_14412,N_6070,N_7776);
xnor U14413 (N_14413,N_9039,N_9002);
or U14414 (N_14414,N_6388,N_5440);
nand U14415 (N_14415,N_9909,N_5048);
or U14416 (N_14416,N_9210,N_8623);
and U14417 (N_14417,N_7838,N_6970);
nand U14418 (N_14418,N_5739,N_5030);
or U14419 (N_14419,N_7453,N_6719);
and U14420 (N_14420,N_6685,N_5969);
or U14421 (N_14421,N_8095,N_8516);
xnor U14422 (N_14422,N_6844,N_8888);
nor U14423 (N_14423,N_5676,N_6318);
nor U14424 (N_14424,N_6079,N_9051);
xnor U14425 (N_14425,N_8969,N_7036);
or U14426 (N_14426,N_6475,N_7693);
or U14427 (N_14427,N_7876,N_8737);
xor U14428 (N_14428,N_8955,N_9320);
xnor U14429 (N_14429,N_5810,N_7651);
or U14430 (N_14430,N_7055,N_5843);
or U14431 (N_14431,N_8587,N_8602);
nor U14432 (N_14432,N_9526,N_9160);
and U14433 (N_14433,N_5447,N_7563);
xor U14434 (N_14434,N_9804,N_6300);
nand U14435 (N_14435,N_7792,N_8901);
xnor U14436 (N_14436,N_5554,N_7888);
nor U14437 (N_14437,N_5441,N_5495);
nand U14438 (N_14438,N_7133,N_8441);
xnor U14439 (N_14439,N_8736,N_9270);
nor U14440 (N_14440,N_7286,N_9670);
or U14441 (N_14441,N_7461,N_6960);
and U14442 (N_14442,N_8874,N_8508);
and U14443 (N_14443,N_8805,N_8993);
and U14444 (N_14444,N_9902,N_6265);
nor U14445 (N_14445,N_5719,N_8916);
or U14446 (N_14446,N_8715,N_6754);
xnor U14447 (N_14447,N_7489,N_5752);
nand U14448 (N_14448,N_8199,N_5015);
or U14449 (N_14449,N_8058,N_8052);
nand U14450 (N_14450,N_6257,N_6086);
and U14451 (N_14451,N_5407,N_8576);
xor U14452 (N_14452,N_7846,N_6835);
or U14453 (N_14453,N_5640,N_9892);
nand U14454 (N_14454,N_9613,N_5922);
or U14455 (N_14455,N_8933,N_7581);
or U14456 (N_14456,N_5725,N_5962);
and U14457 (N_14457,N_6364,N_8681);
and U14458 (N_14458,N_8657,N_9060);
nor U14459 (N_14459,N_7845,N_9490);
nand U14460 (N_14460,N_9532,N_9460);
xor U14461 (N_14461,N_5813,N_7505);
nand U14462 (N_14462,N_6669,N_6536);
and U14463 (N_14463,N_5246,N_7636);
nor U14464 (N_14464,N_5277,N_7125);
or U14465 (N_14465,N_9050,N_8197);
or U14466 (N_14466,N_5752,N_8786);
xnor U14467 (N_14467,N_9762,N_9771);
or U14468 (N_14468,N_7935,N_6080);
or U14469 (N_14469,N_6411,N_5172);
or U14470 (N_14470,N_7346,N_8612);
nor U14471 (N_14471,N_8543,N_7472);
nor U14472 (N_14472,N_5843,N_5084);
nor U14473 (N_14473,N_8607,N_9656);
nand U14474 (N_14474,N_9605,N_6203);
nand U14475 (N_14475,N_6489,N_8086);
or U14476 (N_14476,N_5609,N_9092);
xor U14477 (N_14477,N_7942,N_7376);
or U14478 (N_14478,N_7224,N_6038);
nand U14479 (N_14479,N_5154,N_7624);
xnor U14480 (N_14480,N_8611,N_9534);
nor U14481 (N_14481,N_8981,N_8182);
xor U14482 (N_14482,N_7138,N_9027);
and U14483 (N_14483,N_5493,N_5203);
nor U14484 (N_14484,N_9586,N_7121);
nor U14485 (N_14485,N_6548,N_8084);
and U14486 (N_14486,N_8692,N_9561);
xor U14487 (N_14487,N_5949,N_6492);
xor U14488 (N_14488,N_6757,N_7608);
and U14489 (N_14489,N_6081,N_5278);
or U14490 (N_14490,N_5382,N_7776);
nand U14491 (N_14491,N_6950,N_8502);
or U14492 (N_14492,N_8774,N_7319);
nor U14493 (N_14493,N_5861,N_9661);
or U14494 (N_14494,N_8371,N_8743);
nand U14495 (N_14495,N_8171,N_5546);
nand U14496 (N_14496,N_6690,N_5478);
nor U14497 (N_14497,N_8559,N_6864);
and U14498 (N_14498,N_7181,N_9723);
nand U14499 (N_14499,N_8173,N_8907);
and U14500 (N_14500,N_7745,N_6322);
and U14501 (N_14501,N_8320,N_7885);
xnor U14502 (N_14502,N_9759,N_9410);
nor U14503 (N_14503,N_8104,N_5490);
xor U14504 (N_14504,N_9651,N_7919);
xor U14505 (N_14505,N_5148,N_8432);
nor U14506 (N_14506,N_8102,N_8925);
nor U14507 (N_14507,N_7032,N_9062);
nor U14508 (N_14508,N_8023,N_8967);
xnor U14509 (N_14509,N_8777,N_8974);
and U14510 (N_14510,N_5200,N_9404);
or U14511 (N_14511,N_9509,N_8173);
or U14512 (N_14512,N_9172,N_9494);
and U14513 (N_14513,N_6618,N_5148);
or U14514 (N_14514,N_7256,N_8141);
nand U14515 (N_14515,N_9618,N_7856);
nor U14516 (N_14516,N_9435,N_8455);
nand U14517 (N_14517,N_9070,N_5289);
and U14518 (N_14518,N_5096,N_7378);
nor U14519 (N_14519,N_7666,N_7664);
and U14520 (N_14520,N_5590,N_7483);
nand U14521 (N_14521,N_9619,N_6505);
xor U14522 (N_14522,N_7349,N_9550);
and U14523 (N_14523,N_9620,N_7492);
nor U14524 (N_14524,N_5159,N_5399);
or U14525 (N_14525,N_9353,N_8502);
xor U14526 (N_14526,N_8422,N_5166);
and U14527 (N_14527,N_8832,N_8309);
nand U14528 (N_14528,N_5487,N_8790);
or U14529 (N_14529,N_8272,N_9292);
nand U14530 (N_14530,N_6340,N_9645);
nor U14531 (N_14531,N_7643,N_9222);
nand U14532 (N_14532,N_9457,N_5630);
and U14533 (N_14533,N_9983,N_5999);
or U14534 (N_14534,N_8006,N_8266);
nand U14535 (N_14535,N_9180,N_6500);
nor U14536 (N_14536,N_7123,N_6888);
xnor U14537 (N_14537,N_5477,N_9888);
or U14538 (N_14538,N_7786,N_9028);
nor U14539 (N_14539,N_9758,N_5340);
xor U14540 (N_14540,N_8665,N_9126);
nand U14541 (N_14541,N_6630,N_5243);
xnor U14542 (N_14542,N_6965,N_8419);
and U14543 (N_14543,N_6494,N_6630);
nor U14544 (N_14544,N_7388,N_9798);
and U14545 (N_14545,N_9174,N_9155);
or U14546 (N_14546,N_5059,N_6892);
or U14547 (N_14547,N_6915,N_7211);
nand U14548 (N_14548,N_7969,N_7632);
nor U14549 (N_14549,N_5029,N_5986);
and U14550 (N_14550,N_8133,N_9974);
nor U14551 (N_14551,N_7492,N_6233);
and U14552 (N_14552,N_8754,N_6904);
and U14553 (N_14553,N_7842,N_8648);
xnor U14554 (N_14554,N_7525,N_9093);
nor U14555 (N_14555,N_9912,N_5375);
or U14556 (N_14556,N_9027,N_8107);
xor U14557 (N_14557,N_8534,N_9005);
and U14558 (N_14558,N_6557,N_8462);
and U14559 (N_14559,N_8466,N_8077);
or U14560 (N_14560,N_6580,N_6944);
or U14561 (N_14561,N_9108,N_5095);
nor U14562 (N_14562,N_6458,N_7083);
xor U14563 (N_14563,N_8941,N_8413);
or U14564 (N_14564,N_9532,N_6464);
or U14565 (N_14565,N_9462,N_7705);
nand U14566 (N_14566,N_6088,N_6733);
and U14567 (N_14567,N_7723,N_5993);
xnor U14568 (N_14568,N_6685,N_8169);
xor U14569 (N_14569,N_8622,N_6966);
nand U14570 (N_14570,N_6856,N_5865);
and U14571 (N_14571,N_6634,N_7115);
or U14572 (N_14572,N_9164,N_5759);
and U14573 (N_14573,N_8931,N_6721);
xor U14574 (N_14574,N_5462,N_7918);
or U14575 (N_14575,N_7431,N_5299);
xnor U14576 (N_14576,N_9011,N_7219);
and U14577 (N_14577,N_5365,N_7343);
xor U14578 (N_14578,N_7594,N_7395);
nand U14579 (N_14579,N_8381,N_7795);
xor U14580 (N_14580,N_8086,N_9109);
and U14581 (N_14581,N_7004,N_7169);
nand U14582 (N_14582,N_5382,N_7884);
and U14583 (N_14583,N_6855,N_8796);
xor U14584 (N_14584,N_8640,N_8540);
nand U14585 (N_14585,N_6271,N_7034);
nand U14586 (N_14586,N_5031,N_6984);
and U14587 (N_14587,N_9557,N_5285);
nor U14588 (N_14588,N_9616,N_6479);
and U14589 (N_14589,N_5977,N_5465);
nor U14590 (N_14590,N_8758,N_7136);
and U14591 (N_14591,N_8665,N_5227);
nor U14592 (N_14592,N_7595,N_7611);
or U14593 (N_14593,N_8901,N_7416);
nor U14594 (N_14594,N_6646,N_5976);
and U14595 (N_14595,N_8448,N_7625);
nand U14596 (N_14596,N_7481,N_9383);
and U14597 (N_14597,N_9218,N_5769);
xor U14598 (N_14598,N_6210,N_8981);
xor U14599 (N_14599,N_8507,N_7994);
or U14600 (N_14600,N_7886,N_8356);
and U14601 (N_14601,N_8802,N_6317);
nor U14602 (N_14602,N_7231,N_8446);
and U14603 (N_14603,N_6301,N_7951);
and U14604 (N_14604,N_7229,N_9341);
and U14605 (N_14605,N_8841,N_9145);
nand U14606 (N_14606,N_7102,N_6438);
xor U14607 (N_14607,N_6798,N_6280);
nand U14608 (N_14608,N_5602,N_6356);
nand U14609 (N_14609,N_5804,N_7030);
and U14610 (N_14610,N_8732,N_9524);
nand U14611 (N_14611,N_8531,N_7029);
nand U14612 (N_14612,N_9892,N_5004);
nand U14613 (N_14613,N_6072,N_6677);
and U14614 (N_14614,N_6048,N_9788);
or U14615 (N_14615,N_5995,N_8281);
nand U14616 (N_14616,N_9565,N_5361);
nand U14617 (N_14617,N_5588,N_5472);
xnor U14618 (N_14618,N_5403,N_8578);
or U14619 (N_14619,N_8551,N_5807);
or U14620 (N_14620,N_5159,N_9307);
nor U14621 (N_14621,N_6740,N_7132);
or U14622 (N_14622,N_8616,N_7477);
xnor U14623 (N_14623,N_6386,N_6335);
xor U14624 (N_14624,N_7764,N_8404);
nand U14625 (N_14625,N_6358,N_5030);
nand U14626 (N_14626,N_7579,N_5622);
and U14627 (N_14627,N_6307,N_6646);
xnor U14628 (N_14628,N_5076,N_5815);
xor U14629 (N_14629,N_9478,N_8659);
nand U14630 (N_14630,N_6033,N_9381);
nor U14631 (N_14631,N_6184,N_7265);
nor U14632 (N_14632,N_7927,N_9415);
nor U14633 (N_14633,N_7992,N_7246);
nor U14634 (N_14634,N_9550,N_9161);
or U14635 (N_14635,N_7128,N_5679);
or U14636 (N_14636,N_6557,N_9321);
nor U14637 (N_14637,N_9233,N_7417);
nand U14638 (N_14638,N_9246,N_5434);
nor U14639 (N_14639,N_8924,N_9113);
nor U14640 (N_14640,N_9906,N_9249);
and U14641 (N_14641,N_7538,N_6820);
nand U14642 (N_14642,N_5917,N_9083);
or U14643 (N_14643,N_5582,N_5387);
nor U14644 (N_14644,N_9280,N_6735);
nor U14645 (N_14645,N_7451,N_9459);
nor U14646 (N_14646,N_8625,N_9696);
and U14647 (N_14647,N_5473,N_7725);
xor U14648 (N_14648,N_9897,N_9814);
and U14649 (N_14649,N_8701,N_8427);
xnor U14650 (N_14650,N_9035,N_5619);
nand U14651 (N_14651,N_6533,N_5130);
nand U14652 (N_14652,N_8497,N_7369);
xor U14653 (N_14653,N_5302,N_6172);
and U14654 (N_14654,N_9869,N_9705);
xnor U14655 (N_14655,N_8050,N_6527);
and U14656 (N_14656,N_7487,N_8690);
nor U14657 (N_14657,N_9954,N_6576);
nor U14658 (N_14658,N_7616,N_7938);
nand U14659 (N_14659,N_7600,N_5240);
nor U14660 (N_14660,N_9091,N_6302);
and U14661 (N_14661,N_7135,N_6880);
xnor U14662 (N_14662,N_7196,N_8624);
nor U14663 (N_14663,N_7686,N_5785);
xnor U14664 (N_14664,N_5230,N_7152);
and U14665 (N_14665,N_5506,N_8336);
or U14666 (N_14666,N_5606,N_9791);
nand U14667 (N_14667,N_5326,N_9953);
or U14668 (N_14668,N_7492,N_5406);
xnor U14669 (N_14669,N_8345,N_5106);
and U14670 (N_14670,N_6560,N_5910);
xnor U14671 (N_14671,N_9792,N_9050);
xnor U14672 (N_14672,N_8535,N_7917);
nor U14673 (N_14673,N_9717,N_6858);
nand U14674 (N_14674,N_7664,N_9153);
nand U14675 (N_14675,N_9254,N_5855);
xnor U14676 (N_14676,N_8324,N_8382);
or U14677 (N_14677,N_8590,N_5422);
and U14678 (N_14678,N_6594,N_9863);
xnor U14679 (N_14679,N_8167,N_7853);
xnor U14680 (N_14680,N_8846,N_5882);
xnor U14681 (N_14681,N_5728,N_8071);
nand U14682 (N_14682,N_5603,N_5369);
nor U14683 (N_14683,N_9058,N_7450);
xor U14684 (N_14684,N_8891,N_5591);
xor U14685 (N_14685,N_8506,N_7580);
nand U14686 (N_14686,N_9941,N_7785);
nand U14687 (N_14687,N_7082,N_6283);
nor U14688 (N_14688,N_6428,N_9159);
and U14689 (N_14689,N_5172,N_5656);
xor U14690 (N_14690,N_9490,N_8364);
xor U14691 (N_14691,N_9742,N_9826);
nor U14692 (N_14692,N_5059,N_6456);
nor U14693 (N_14693,N_8680,N_9812);
nor U14694 (N_14694,N_7148,N_7271);
nor U14695 (N_14695,N_9256,N_5213);
xnor U14696 (N_14696,N_8810,N_9912);
or U14697 (N_14697,N_6841,N_8246);
or U14698 (N_14698,N_6173,N_9524);
xor U14699 (N_14699,N_8253,N_7447);
nor U14700 (N_14700,N_8413,N_5489);
and U14701 (N_14701,N_6726,N_8262);
xnor U14702 (N_14702,N_8460,N_5133);
or U14703 (N_14703,N_9143,N_7012);
nand U14704 (N_14704,N_8499,N_8319);
xnor U14705 (N_14705,N_9516,N_9234);
and U14706 (N_14706,N_9748,N_8949);
nor U14707 (N_14707,N_9304,N_9946);
nand U14708 (N_14708,N_9301,N_5125);
or U14709 (N_14709,N_7404,N_6010);
and U14710 (N_14710,N_8384,N_7361);
nor U14711 (N_14711,N_9131,N_6052);
xnor U14712 (N_14712,N_9071,N_8082);
xnor U14713 (N_14713,N_6378,N_5635);
or U14714 (N_14714,N_7002,N_7116);
nand U14715 (N_14715,N_5293,N_8007);
nand U14716 (N_14716,N_9091,N_8639);
and U14717 (N_14717,N_8655,N_7646);
nor U14718 (N_14718,N_9093,N_7220);
and U14719 (N_14719,N_5625,N_9200);
nor U14720 (N_14720,N_8939,N_9177);
nand U14721 (N_14721,N_5575,N_9206);
nor U14722 (N_14722,N_5871,N_9798);
nor U14723 (N_14723,N_6209,N_9123);
xor U14724 (N_14724,N_5119,N_5057);
or U14725 (N_14725,N_5202,N_7719);
nor U14726 (N_14726,N_7427,N_8233);
or U14727 (N_14727,N_6624,N_6425);
nand U14728 (N_14728,N_6068,N_5108);
nand U14729 (N_14729,N_9106,N_9063);
and U14730 (N_14730,N_6277,N_5015);
or U14731 (N_14731,N_8693,N_5859);
nor U14732 (N_14732,N_7556,N_8861);
nor U14733 (N_14733,N_7410,N_7919);
nand U14734 (N_14734,N_8376,N_8115);
xnor U14735 (N_14735,N_7651,N_9223);
nand U14736 (N_14736,N_9977,N_7411);
or U14737 (N_14737,N_5380,N_9024);
nand U14738 (N_14738,N_8676,N_6817);
xor U14739 (N_14739,N_9511,N_7188);
xor U14740 (N_14740,N_7174,N_6153);
nor U14741 (N_14741,N_5137,N_9250);
or U14742 (N_14742,N_6390,N_8842);
or U14743 (N_14743,N_9589,N_7366);
nand U14744 (N_14744,N_8001,N_9543);
xor U14745 (N_14745,N_6505,N_8860);
nor U14746 (N_14746,N_5291,N_8087);
nor U14747 (N_14747,N_7815,N_9810);
xnor U14748 (N_14748,N_6629,N_9535);
or U14749 (N_14749,N_8841,N_9823);
nand U14750 (N_14750,N_5689,N_7087);
xor U14751 (N_14751,N_6790,N_7278);
or U14752 (N_14752,N_8601,N_5082);
nor U14753 (N_14753,N_7970,N_7630);
and U14754 (N_14754,N_5135,N_8359);
nand U14755 (N_14755,N_7641,N_8185);
nor U14756 (N_14756,N_7051,N_9696);
xnor U14757 (N_14757,N_6886,N_7115);
xor U14758 (N_14758,N_5277,N_8937);
or U14759 (N_14759,N_5309,N_6268);
xnor U14760 (N_14760,N_9401,N_7423);
nand U14761 (N_14761,N_7618,N_9936);
xor U14762 (N_14762,N_8084,N_6044);
xnor U14763 (N_14763,N_9445,N_8930);
nand U14764 (N_14764,N_6075,N_8056);
nand U14765 (N_14765,N_5523,N_8213);
nand U14766 (N_14766,N_6489,N_8674);
nand U14767 (N_14767,N_9459,N_5844);
nand U14768 (N_14768,N_7951,N_5719);
or U14769 (N_14769,N_6739,N_7475);
nor U14770 (N_14770,N_5955,N_9019);
nor U14771 (N_14771,N_6227,N_8693);
and U14772 (N_14772,N_5849,N_5949);
nand U14773 (N_14773,N_9436,N_8153);
xor U14774 (N_14774,N_5266,N_8494);
or U14775 (N_14775,N_6171,N_6211);
nand U14776 (N_14776,N_6634,N_7180);
xnor U14777 (N_14777,N_9597,N_6139);
xnor U14778 (N_14778,N_9424,N_7144);
nor U14779 (N_14779,N_7436,N_5713);
xor U14780 (N_14780,N_9528,N_9058);
nand U14781 (N_14781,N_5249,N_5338);
nand U14782 (N_14782,N_8795,N_9296);
and U14783 (N_14783,N_6362,N_9111);
nor U14784 (N_14784,N_6269,N_7395);
or U14785 (N_14785,N_6439,N_9883);
and U14786 (N_14786,N_5299,N_8567);
xnor U14787 (N_14787,N_9851,N_7699);
or U14788 (N_14788,N_9912,N_9012);
nand U14789 (N_14789,N_8716,N_5188);
and U14790 (N_14790,N_8718,N_9528);
and U14791 (N_14791,N_5152,N_7834);
xor U14792 (N_14792,N_9781,N_5856);
and U14793 (N_14793,N_9095,N_5993);
or U14794 (N_14794,N_5793,N_8259);
xor U14795 (N_14795,N_7544,N_5495);
and U14796 (N_14796,N_9629,N_5306);
nand U14797 (N_14797,N_5487,N_5570);
and U14798 (N_14798,N_5965,N_7321);
and U14799 (N_14799,N_9459,N_9101);
nand U14800 (N_14800,N_7232,N_5075);
xor U14801 (N_14801,N_5838,N_9833);
xor U14802 (N_14802,N_6988,N_6746);
nor U14803 (N_14803,N_6243,N_7035);
nand U14804 (N_14804,N_6471,N_7790);
or U14805 (N_14805,N_5149,N_7443);
or U14806 (N_14806,N_7603,N_9100);
xor U14807 (N_14807,N_8041,N_8515);
and U14808 (N_14808,N_5507,N_6052);
xnor U14809 (N_14809,N_7365,N_9185);
nand U14810 (N_14810,N_8738,N_5856);
and U14811 (N_14811,N_9915,N_6899);
xnor U14812 (N_14812,N_5118,N_6663);
nor U14813 (N_14813,N_5119,N_9783);
xnor U14814 (N_14814,N_5446,N_8599);
xor U14815 (N_14815,N_6196,N_6168);
nand U14816 (N_14816,N_9941,N_6517);
xnor U14817 (N_14817,N_7248,N_9318);
nor U14818 (N_14818,N_5704,N_7519);
or U14819 (N_14819,N_8067,N_8414);
nor U14820 (N_14820,N_6333,N_7582);
or U14821 (N_14821,N_7979,N_7283);
nor U14822 (N_14822,N_9329,N_7105);
and U14823 (N_14823,N_5115,N_7966);
or U14824 (N_14824,N_9112,N_8639);
and U14825 (N_14825,N_6946,N_9827);
nor U14826 (N_14826,N_6683,N_9963);
nor U14827 (N_14827,N_7353,N_5456);
or U14828 (N_14828,N_6051,N_5036);
nand U14829 (N_14829,N_6849,N_7940);
xor U14830 (N_14830,N_6184,N_5765);
xor U14831 (N_14831,N_5988,N_5471);
and U14832 (N_14832,N_9254,N_8928);
and U14833 (N_14833,N_7663,N_7575);
xnor U14834 (N_14834,N_6391,N_5104);
nor U14835 (N_14835,N_8371,N_5267);
xnor U14836 (N_14836,N_8736,N_9610);
xor U14837 (N_14837,N_5379,N_6913);
nor U14838 (N_14838,N_8025,N_9795);
nand U14839 (N_14839,N_9718,N_5062);
xor U14840 (N_14840,N_5879,N_5773);
nand U14841 (N_14841,N_5651,N_9233);
xnor U14842 (N_14842,N_5635,N_6296);
nor U14843 (N_14843,N_7215,N_9742);
and U14844 (N_14844,N_9215,N_9354);
nor U14845 (N_14845,N_7506,N_7496);
nor U14846 (N_14846,N_6132,N_9221);
and U14847 (N_14847,N_7548,N_5945);
or U14848 (N_14848,N_8307,N_9763);
nand U14849 (N_14849,N_8928,N_9827);
xor U14850 (N_14850,N_6963,N_8959);
or U14851 (N_14851,N_5230,N_8778);
nand U14852 (N_14852,N_5388,N_9044);
nor U14853 (N_14853,N_5174,N_9317);
xor U14854 (N_14854,N_9164,N_9222);
nor U14855 (N_14855,N_7023,N_8560);
xor U14856 (N_14856,N_9405,N_7149);
and U14857 (N_14857,N_9299,N_6157);
nor U14858 (N_14858,N_5836,N_8544);
or U14859 (N_14859,N_8266,N_5811);
or U14860 (N_14860,N_7527,N_6091);
or U14861 (N_14861,N_9671,N_6404);
or U14862 (N_14862,N_7880,N_8054);
xnor U14863 (N_14863,N_5410,N_7871);
or U14864 (N_14864,N_6493,N_5173);
xnor U14865 (N_14865,N_7041,N_9706);
and U14866 (N_14866,N_5384,N_5389);
xnor U14867 (N_14867,N_6712,N_7191);
xor U14868 (N_14868,N_8783,N_6131);
or U14869 (N_14869,N_7821,N_7395);
and U14870 (N_14870,N_7869,N_5860);
or U14871 (N_14871,N_6109,N_6069);
xnor U14872 (N_14872,N_9661,N_5461);
nor U14873 (N_14873,N_8431,N_7490);
and U14874 (N_14874,N_8283,N_7793);
xor U14875 (N_14875,N_5408,N_8600);
nand U14876 (N_14876,N_7508,N_9809);
nor U14877 (N_14877,N_8138,N_6443);
nor U14878 (N_14878,N_9170,N_6207);
nand U14879 (N_14879,N_5348,N_6076);
nand U14880 (N_14880,N_6001,N_7670);
nor U14881 (N_14881,N_5795,N_6670);
xnor U14882 (N_14882,N_9172,N_8476);
or U14883 (N_14883,N_8154,N_7168);
or U14884 (N_14884,N_8933,N_7235);
xor U14885 (N_14885,N_5639,N_8397);
nor U14886 (N_14886,N_9154,N_9699);
nand U14887 (N_14887,N_6762,N_7206);
xor U14888 (N_14888,N_8197,N_8617);
or U14889 (N_14889,N_6743,N_9181);
nand U14890 (N_14890,N_5807,N_5359);
or U14891 (N_14891,N_6363,N_9291);
or U14892 (N_14892,N_7021,N_5389);
nand U14893 (N_14893,N_7969,N_8768);
and U14894 (N_14894,N_7712,N_6428);
xnor U14895 (N_14895,N_8728,N_7947);
nand U14896 (N_14896,N_5791,N_8630);
xnor U14897 (N_14897,N_8602,N_7583);
xor U14898 (N_14898,N_8378,N_6819);
xor U14899 (N_14899,N_6667,N_7744);
nand U14900 (N_14900,N_9526,N_7450);
or U14901 (N_14901,N_7050,N_7091);
nand U14902 (N_14902,N_9571,N_5890);
xor U14903 (N_14903,N_6256,N_5590);
xor U14904 (N_14904,N_5042,N_5776);
nor U14905 (N_14905,N_7748,N_9994);
nand U14906 (N_14906,N_5973,N_9248);
or U14907 (N_14907,N_8491,N_6402);
and U14908 (N_14908,N_6949,N_5115);
xor U14909 (N_14909,N_8275,N_8841);
xnor U14910 (N_14910,N_5872,N_7589);
or U14911 (N_14911,N_6037,N_7496);
nor U14912 (N_14912,N_9073,N_5394);
xnor U14913 (N_14913,N_8687,N_8880);
and U14914 (N_14914,N_5561,N_7126);
nand U14915 (N_14915,N_8280,N_5218);
nor U14916 (N_14916,N_5133,N_9336);
nand U14917 (N_14917,N_8470,N_9624);
xor U14918 (N_14918,N_5738,N_7844);
xor U14919 (N_14919,N_9775,N_5446);
xor U14920 (N_14920,N_9386,N_9060);
nand U14921 (N_14921,N_9468,N_9740);
or U14922 (N_14922,N_9641,N_5233);
and U14923 (N_14923,N_8144,N_5317);
xnor U14924 (N_14924,N_5597,N_5219);
xnor U14925 (N_14925,N_7920,N_7301);
xor U14926 (N_14926,N_8916,N_8167);
nand U14927 (N_14927,N_6160,N_5977);
xor U14928 (N_14928,N_7865,N_5081);
xor U14929 (N_14929,N_7324,N_7265);
xnor U14930 (N_14930,N_5840,N_6894);
and U14931 (N_14931,N_8221,N_8591);
or U14932 (N_14932,N_7242,N_9546);
xor U14933 (N_14933,N_8241,N_6037);
nand U14934 (N_14934,N_7702,N_8488);
or U14935 (N_14935,N_5865,N_8539);
and U14936 (N_14936,N_7510,N_7363);
and U14937 (N_14937,N_5758,N_6382);
nor U14938 (N_14938,N_7900,N_7792);
or U14939 (N_14939,N_9295,N_9285);
xor U14940 (N_14940,N_6027,N_8055);
or U14941 (N_14941,N_5769,N_8572);
nand U14942 (N_14942,N_5363,N_9779);
xor U14943 (N_14943,N_9442,N_5229);
and U14944 (N_14944,N_6103,N_6905);
nand U14945 (N_14945,N_5152,N_5213);
nor U14946 (N_14946,N_9069,N_8111);
nand U14947 (N_14947,N_5313,N_6065);
nor U14948 (N_14948,N_6155,N_8010);
nand U14949 (N_14949,N_7180,N_7442);
nor U14950 (N_14950,N_7911,N_6633);
and U14951 (N_14951,N_5680,N_6089);
nand U14952 (N_14952,N_7569,N_8149);
or U14953 (N_14953,N_7852,N_6001);
nand U14954 (N_14954,N_6955,N_9644);
nand U14955 (N_14955,N_9455,N_7685);
nor U14956 (N_14956,N_9118,N_9878);
nand U14957 (N_14957,N_7956,N_9519);
or U14958 (N_14958,N_7890,N_9858);
nand U14959 (N_14959,N_5692,N_7897);
xor U14960 (N_14960,N_7563,N_6275);
nand U14961 (N_14961,N_6381,N_7625);
nor U14962 (N_14962,N_7975,N_5591);
xnor U14963 (N_14963,N_6321,N_7144);
nor U14964 (N_14964,N_9848,N_7888);
xor U14965 (N_14965,N_9676,N_8202);
or U14966 (N_14966,N_7401,N_9910);
nand U14967 (N_14967,N_9828,N_7854);
nand U14968 (N_14968,N_6879,N_7851);
nand U14969 (N_14969,N_5944,N_5867);
and U14970 (N_14970,N_6009,N_5680);
nand U14971 (N_14971,N_8110,N_6203);
and U14972 (N_14972,N_9832,N_8072);
xnor U14973 (N_14973,N_7977,N_5561);
or U14974 (N_14974,N_9089,N_7928);
or U14975 (N_14975,N_9704,N_8885);
and U14976 (N_14976,N_6151,N_5270);
or U14977 (N_14977,N_5626,N_9682);
and U14978 (N_14978,N_8557,N_8158);
nor U14979 (N_14979,N_7610,N_7217);
xnor U14980 (N_14980,N_6935,N_6644);
and U14981 (N_14981,N_8874,N_7685);
and U14982 (N_14982,N_5674,N_9655);
or U14983 (N_14983,N_6290,N_9039);
or U14984 (N_14984,N_5162,N_6339);
and U14985 (N_14985,N_5659,N_7495);
nor U14986 (N_14986,N_5514,N_8571);
and U14987 (N_14987,N_8654,N_8070);
xor U14988 (N_14988,N_5442,N_7252);
and U14989 (N_14989,N_9062,N_8384);
or U14990 (N_14990,N_8237,N_7253);
nor U14991 (N_14991,N_8939,N_5726);
and U14992 (N_14992,N_9578,N_8668);
xor U14993 (N_14993,N_8438,N_8829);
nand U14994 (N_14994,N_8016,N_9906);
and U14995 (N_14995,N_8449,N_7878);
and U14996 (N_14996,N_8751,N_8722);
and U14997 (N_14997,N_7025,N_7473);
xor U14998 (N_14998,N_7220,N_5591);
nor U14999 (N_14999,N_6035,N_8973);
or U15000 (N_15000,N_10340,N_12362);
nor U15001 (N_15001,N_10110,N_10753);
nor U15002 (N_15002,N_10204,N_13660);
nand U15003 (N_15003,N_10149,N_12853);
and U15004 (N_15004,N_10623,N_11078);
and U15005 (N_15005,N_10937,N_12579);
xnor U15006 (N_15006,N_11372,N_12428);
xor U15007 (N_15007,N_10010,N_11749);
and U15008 (N_15008,N_14810,N_13340);
nand U15009 (N_15009,N_13692,N_14232);
nand U15010 (N_15010,N_10516,N_10769);
nand U15011 (N_15011,N_11659,N_13084);
nand U15012 (N_15012,N_14778,N_11275);
and U15013 (N_15013,N_10543,N_11323);
and U15014 (N_15014,N_11314,N_12928);
nand U15015 (N_15015,N_13865,N_10674);
or U15016 (N_15016,N_14420,N_13133);
nand U15017 (N_15017,N_10739,N_13507);
or U15018 (N_15018,N_14352,N_10459);
or U15019 (N_15019,N_11752,N_10185);
nand U15020 (N_15020,N_10033,N_12472);
or U15021 (N_15021,N_10875,N_10154);
or U15022 (N_15022,N_11972,N_12888);
xnor U15023 (N_15023,N_11953,N_13763);
and U15024 (N_15024,N_11181,N_11765);
xnor U15025 (N_15025,N_13860,N_13758);
or U15026 (N_15026,N_12628,N_13969);
nor U15027 (N_15027,N_12064,N_12829);
xor U15028 (N_15028,N_13360,N_12606);
xnor U15029 (N_15029,N_10494,N_12059);
nand U15030 (N_15030,N_10917,N_12661);
nand U15031 (N_15031,N_11412,N_13687);
or U15032 (N_15032,N_13427,N_12484);
or U15033 (N_15033,N_10272,N_10467);
nor U15034 (N_15034,N_10828,N_11886);
nor U15035 (N_15035,N_11766,N_10750);
xnor U15036 (N_15036,N_13423,N_11384);
xor U15037 (N_15037,N_14645,N_10034);
nand U15038 (N_15038,N_14834,N_11205);
or U15039 (N_15039,N_13734,N_13998);
or U15040 (N_15040,N_11464,N_11396);
or U15041 (N_15041,N_12728,N_11948);
nor U15042 (N_15042,N_11890,N_10121);
and U15043 (N_15043,N_12274,N_13509);
xor U15044 (N_15044,N_13454,N_14535);
or U15045 (N_15045,N_10525,N_14924);
or U15046 (N_15046,N_11695,N_11495);
nor U15047 (N_15047,N_13887,N_13718);
and U15048 (N_15048,N_11176,N_11018);
or U15049 (N_15049,N_14942,N_14564);
or U15050 (N_15050,N_11658,N_13450);
or U15051 (N_15051,N_14307,N_11798);
and U15052 (N_15052,N_14584,N_10539);
nor U15053 (N_15053,N_10305,N_12151);
nand U15054 (N_15054,N_12838,N_14050);
or U15055 (N_15055,N_11194,N_11135);
nor U15056 (N_15056,N_12264,N_13873);
nor U15057 (N_15057,N_13749,N_10571);
xor U15058 (N_15058,N_12974,N_11029);
nand U15059 (N_15059,N_10732,N_11125);
xor U15060 (N_15060,N_13521,N_12494);
nor U15061 (N_15061,N_10704,N_14479);
xor U15062 (N_15062,N_12907,N_14573);
xnor U15063 (N_15063,N_13961,N_11344);
nand U15064 (N_15064,N_11224,N_13292);
and U15065 (N_15065,N_11967,N_10225);
nand U15066 (N_15066,N_14657,N_14663);
nor U15067 (N_15067,N_11044,N_13201);
nand U15068 (N_15068,N_14684,N_12052);
nand U15069 (N_15069,N_14046,N_11005);
and U15070 (N_15070,N_14056,N_14636);
nand U15071 (N_15071,N_13033,N_14255);
xor U15072 (N_15072,N_10883,N_12298);
nor U15073 (N_15073,N_11607,N_14516);
nor U15074 (N_15074,N_10406,N_10288);
and U15075 (N_15075,N_12900,N_13676);
xnor U15076 (N_15076,N_14514,N_13220);
xnor U15077 (N_15077,N_11951,N_14257);
nor U15078 (N_15078,N_11883,N_10952);
nor U15079 (N_15079,N_14559,N_10684);
and U15080 (N_15080,N_10632,N_10138);
nor U15081 (N_15081,N_14758,N_11368);
nor U15082 (N_15082,N_14945,N_10797);
nor U15083 (N_15083,N_13547,N_14768);
or U15084 (N_15084,N_14033,N_13845);
xnor U15085 (N_15085,N_10766,N_14868);
nand U15086 (N_15086,N_11192,N_11800);
xnor U15087 (N_15087,N_13834,N_12410);
nand U15088 (N_15088,N_14268,N_11515);
xnor U15089 (N_15089,N_13601,N_12164);
or U15090 (N_15090,N_14315,N_10823);
and U15091 (N_15091,N_10546,N_12327);
and U15092 (N_15092,N_12778,N_12012);
nand U15093 (N_15093,N_14245,N_13376);
or U15094 (N_15094,N_10462,N_11359);
xor U15095 (N_15095,N_14204,N_13200);
xor U15096 (N_15096,N_13207,N_10230);
xor U15097 (N_15097,N_13142,N_13334);
nor U15098 (N_15098,N_12535,N_12003);
nor U15099 (N_15099,N_10142,N_10680);
nor U15100 (N_15100,N_14226,N_11263);
and U15101 (N_15101,N_12857,N_11006);
nand U15102 (N_15102,N_13569,N_13003);
nand U15103 (N_15103,N_10866,N_13812);
and U15104 (N_15104,N_14958,N_14067);
nor U15105 (N_15105,N_13818,N_11310);
and U15106 (N_15106,N_11492,N_14458);
or U15107 (N_15107,N_11682,N_14493);
nor U15108 (N_15108,N_14335,N_11411);
nor U15109 (N_15109,N_12748,N_14836);
nor U15110 (N_15110,N_11012,N_13743);
and U15111 (N_15111,N_13032,N_10556);
and U15112 (N_15112,N_12948,N_14682);
nor U15113 (N_15113,N_10175,N_10846);
nor U15114 (N_15114,N_14926,N_10384);
nand U15115 (N_15115,N_14716,N_14691);
nor U15116 (N_15116,N_14963,N_12211);
and U15117 (N_15117,N_11404,N_10805);
xnor U15118 (N_15118,N_12166,N_12419);
and U15119 (N_15119,N_13786,N_10511);
and U15120 (N_15120,N_14146,N_13439);
xnor U15121 (N_15121,N_13821,N_11385);
xnor U15122 (N_15122,N_14787,N_10727);
and U15123 (N_15123,N_13036,N_11417);
xor U15124 (N_15124,N_12726,N_10057);
nand U15125 (N_15125,N_11295,N_13807);
or U15126 (N_15126,N_11994,N_13977);
xnor U15127 (N_15127,N_10194,N_14852);
and U15128 (N_15128,N_12294,N_13584);
xor U15129 (N_15129,N_14041,N_12574);
nand U15130 (N_15130,N_12011,N_14861);
xnor U15131 (N_15131,N_14111,N_11260);
nor U15132 (N_15132,N_11197,N_12476);
and U15133 (N_15133,N_14314,N_14741);
nor U15134 (N_15134,N_14103,N_12334);
or U15135 (N_15135,N_10620,N_11097);
or U15136 (N_15136,N_13504,N_13937);
and U15137 (N_15137,N_11387,N_11598);
nand U15138 (N_15138,N_13952,N_10346);
nor U15139 (N_15139,N_14739,N_14609);
and U15140 (N_15140,N_13492,N_10755);
nand U15141 (N_15141,N_12608,N_11362);
nor U15142 (N_15142,N_14605,N_10545);
and U15143 (N_15143,N_12507,N_10878);
and U15144 (N_15144,N_11661,N_11882);
nand U15145 (N_15145,N_13076,N_11638);
nand U15146 (N_15146,N_13122,N_14260);
nand U15147 (N_15147,N_12429,N_14976);
or U15148 (N_15148,N_11085,N_14017);
xor U15149 (N_15149,N_11028,N_13377);
nand U15150 (N_15150,N_10255,N_13510);
xor U15151 (N_15151,N_11380,N_13208);
or U15152 (N_15152,N_11735,N_14927);
xor U15153 (N_15153,N_11833,N_14038);
xor U15154 (N_15154,N_13674,N_14598);
nor U15155 (N_15155,N_13609,N_14404);
xor U15156 (N_15156,N_10134,N_11774);
nor U15157 (N_15157,N_12030,N_10446);
and U15158 (N_15158,N_10763,N_11755);
xor U15159 (N_15159,N_13737,N_11978);
nor U15160 (N_15160,N_11154,N_13101);
or U15161 (N_15161,N_14365,N_11191);
nand U15162 (N_15162,N_14272,N_12146);
nand U15163 (N_15163,N_10061,N_14813);
or U15164 (N_15164,N_11347,N_13481);
nand U15165 (N_15165,N_14387,N_11927);
nand U15166 (N_15166,N_13310,N_10504);
nand U15167 (N_15167,N_12941,N_14993);
nor U15168 (N_15168,N_10757,N_11829);
or U15169 (N_15169,N_10964,N_10053);
and U15170 (N_15170,N_11113,N_13617);
xnor U15171 (N_15171,N_11393,N_14597);
xor U15172 (N_15172,N_14150,N_14986);
and U15173 (N_15173,N_11803,N_10224);
or U15174 (N_15174,N_10103,N_11738);
xor U15175 (N_15175,N_13940,N_11955);
xor U15176 (N_15176,N_12277,N_14552);
or U15177 (N_15177,N_14974,N_12315);
xor U15178 (N_15178,N_14793,N_11488);
and U15179 (N_15179,N_11742,N_14385);
nor U15180 (N_15180,N_12717,N_12385);
xnor U15181 (N_15181,N_14862,N_10635);
xor U15182 (N_15182,N_13506,N_10938);
or U15183 (N_15183,N_13877,N_13105);
nand U15184 (N_15184,N_13627,N_12955);
or U15185 (N_15185,N_10710,N_13452);
and U15186 (N_15186,N_12831,N_10021);
nand U15187 (N_15187,N_10013,N_13703);
or U15188 (N_15188,N_11108,N_14959);
nand U15189 (N_15189,N_12510,N_10017);
xnor U15190 (N_15190,N_12015,N_14014);
xnor U15191 (N_15191,N_12964,N_13104);
or U15192 (N_15192,N_11068,N_10362);
nor U15193 (N_15193,N_11778,N_11276);
or U15194 (N_15194,N_11054,N_11535);
nor U15195 (N_15195,N_10093,N_14646);
or U15196 (N_15196,N_11203,N_13026);
or U15197 (N_15197,N_13429,N_13422);
and U15198 (N_15198,N_12947,N_12988);
and U15199 (N_15199,N_14745,N_12055);
xor U15200 (N_15200,N_10508,N_14074);
or U15201 (N_15201,N_13438,N_11485);
nor U15202 (N_15202,N_11437,N_12361);
xor U15203 (N_15203,N_14702,N_14360);
and U15204 (N_15204,N_13193,N_12039);
and U15205 (N_15205,N_11024,N_12806);
nor U15206 (N_15206,N_13619,N_11484);
or U15207 (N_15207,N_14081,N_11573);
xnor U15208 (N_15208,N_14421,N_11242);
nor U15209 (N_15209,N_13960,N_10169);
xnor U15210 (N_15210,N_13802,N_13318);
nand U15211 (N_15211,N_10321,N_12825);
xor U15212 (N_15212,N_12196,N_10082);
and U15213 (N_15213,N_13012,N_12391);
nand U15214 (N_15214,N_12513,N_10649);
nor U15215 (N_15215,N_10997,N_12587);
xor U15216 (N_15216,N_14275,N_14614);
nand U15217 (N_15217,N_10312,N_10977);
xor U15218 (N_15218,N_10583,N_11353);
nand U15219 (N_15219,N_13551,N_10709);
nor U15220 (N_15220,N_14794,N_11812);
xnor U15221 (N_15221,N_12404,N_11988);
and U15222 (N_15222,N_11046,N_13369);
or U15223 (N_15223,N_12783,N_14631);
and U15224 (N_15224,N_13275,N_14051);
or U15225 (N_15225,N_13565,N_10834);
and U15226 (N_15226,N_13349,N_14890);
or U15227 (N_15227,N_14715,N_10063);
nor U15228 (N_15228,N_11164,N_10817);
xnor U15229 (N_15229,N_10113,N_13090);
and U15230 (N_15230,N_10024,N_12545);
and U15231 (N_15231,N_14685,N_13889);
xor U15232 (N_15232,N_11151,N_12412);
nor U15233 (N_15233,N_13278,N_10311);
xor U15234 (N_15234,N_11261,N_11872);
and U15235 (N_15235,N_14444,N_13790);
xnor U15236 (N_15236,N_10374,N_13162);
or U15237 (N_15237,N_13339,N_14846);
nor U15238 (N_15238,N_11400,N_11581);
or U15239 (N_15239,N_14374,N_11633);
and U15240 (N_15240,N_12503,N_11590);
xnor U15241 (N_15241,N_10588,N_13679);
and U15242 (N_15242,N_12205,N_12051);
nor U15243 (N_15243,N_10337,N_11834);
nor U15244 (N_15244,N_14087,N_11976);
or U15245 (N_15245,N_14606,N_11835);
xor U15246 (N_15246,N_11616,N_14991);
nand U15247 (N_15247,N_10810,N_11900);
xor U15248 (N_15248,N_11991,N_14877);
nor U15249 (N_15249,N_13820,N_12359);
nor U15250 (N_15250,N_14107,N_12733);
and U15251 (N_15251,N_10835,N_10733);
xnor U15252 (N_15252,N_10333,N_10485);
nor U15253 (N_15253,N_12635,N_12650);
and U15254 (N_15254,N_12025,N_12667);
nor U15255 (N_15255,N_11286,N_13698);
xor U15256 (N_15256,N_14367,N_10574);
nor U15257 (N_15257,N_14343,N_11142);
xnor U15258 (N_15258,N_12720,N_12906);
or U15259 (N_15259,N_12155,N_12331);
xor U15260 (N_15260,N_11600,N_13091);
nor U15261 (N_15261,N_14531,N_12275);
nor U15262 (N_15262,N_10076,N_13638);
or U15263 (N_15263,N_13533,N_14950);
xnor U15264 (N_15264,N_12345,N_14357);
and U15265 (N_15265,N_14030,N_13585);
or U15266 (N_15266,N_12553,N_13519);
nand U15267 (N_15267,N_14833,N_10612);
xor U15268 (N_15268,N_13596,N_12204);
xnor U15269 (N_15269,N_13707,N_14160);
or U15270 (N_15270,N_12668,N_11462);
and U15271 (N_15271,N_11451,N_12420);
nor U15272 (N_15272,N_10136,N_10568);
or U15273 (N_15273,N_12208,N_14929);
nand U15274 (N_15274,N_13525,N_14553);
and U15275 (N_15275,N_11719,N_12341);
xor U15276 (N_15276,N_10438,N_13684);
xnor U15277 (N_15277,N_12256,N_12103);
xnor U15278 (N_15278,N_14034,N_13906);
xnor U15279 (N_15279,N_14453,N_14086);
nand U15280 (N_15280,N_12687,N_14220);
xnor U15281 (N_15281,N_12532,N_13579);
and U15282 (N_15282,N_10278,N_11264);
nor U15283 (N_15283,N_10716,N_12394);
nor U15284 (N_15284,N_14289,N_14110);
or U15285 (N_15285,N_14490,N_13295);
or U15286 (N_15286,N_13885,N_12525);
nand U15287 (N_15287,N_14743,N_14995);
xnor U15288 (N_15288,N_11888,N_11623);
and U15289 (N_15289,N_13226,N_13994);
or U15290 (N_15290,N_13963,N_13414);
or U15291 (N_15291,N_10644,N_12489);
xor U15292 (N_15292,N_13361,N_13260);
xnor U15293 (N_15293,N_13232,N_14057);
xnor U15294 (N_15294,N_10125,N_14388);
nand U15295 (N_15295,N_12550,N_13120);
and U15296 (N_15296,N_12214,N_14960);
nor U15297 (N_15297,N_14258,N_12267);
or U15298 (N_15298,N_13756,N_12581);
nand U15299 (N_15299,N_11156,N_10735);
xnor U15300 (N_15300,N_13591,N_12908);
or U15301 (N_15301,N_13555,N_14376);
or U15302 (N_15302,N_13726,N_13110);
and U15303 (N_15303,N_11069,N_14709);
nand U15304 (N_15304,N_10648,N_13497);
nand U15305 (N_15305,N_14148,N_13253);
nor U15306 (N_15306,N_13313,N_14353);
and U15307 (N_15307,N_12916,N_11392);
nand U15308 (N_15308,N_12980,N_12056);
nand U15309 (N_15309,N_12010,N_13534);
or U15310 (N_15310,N_14049,N_14707);
and U15311 (N_15311,N_10873,N_11440);
xor U15312 (N_15312,N_12261,N_13308);
and U15313 (N_15313,N_13686,N_11289);
nand U15314 (N_15314,N_14529,N_11618);
or U15315 (N_15315,N_11258,N_13801);
or U15316 (N_15316,N_13092,N_14733);
or U15317 (N_15317,N_10297,N_12811);
or U15318 (N_15318,N_11060,N_11330);
nand U15319 (N_15319,N_12803,N_10655);
nand U15320 (N_15320,N_12221,N_14708);
and U15321 (N_15321,N_11525,N_12035);
nand U15322 (N_15322,N_12626,N_14219);
or U15323 (N_15323,N_14690,N_11799);
and U15324 (N_15324,N_12839,N_13789);
nor U15325 (N_15325,N_14263,N_14306);
xor U15326 (N_15326,N_10394,N_14457);
xor U15327 (N_15327,N_12502,N_13018);
and U15328 (N_15328,N_14015,N_12772);
nand U15329 (N_15329,N_13071,N_14678);
and U15330 (N_15330,N_12442,N_12674);
and U15331 (N_15331,N_12411,N_10816);
xnor U15332 (N_15332,N_12771,N_13849);
nand U15333 (N_15333,N_11360,N_12586);
nor U15334 (N_15334,N_14802,N_13975);
and U15335 (N_15335,N_11397,N_14456);
nor U15336 (N_15336,N_13128,N_14888);
nor U15337 (N_15337,N_12648,N_10106);
nor U15338 (N_15338,N_13389,N_13293);
and U15339 (N_15339,N_10885,N_10178);
or U15340 (N_15340,N_10074,N_12738);
nand U15341 (N_15341,N_13513,N_11849);
or U15342 (N_15342,N_10144,N_12913);
nor U15343 (N_15343,N_14892,N_12631);
nand U15344 (N_15344,N_11469,N_11183);
and U15345 (N_15345,N_12346,N_11291);
nand U15346 (N_15346,N_12367,N_12505);
nor U15347 (N_15347,N_13413,N_13327);
nor U15348 (N_15348,N_12449,N_12705);
xor U15349 (N_15349,N_14189,N_11839);
nand U15350 (N_15350,N_12396,N_13938);
nor U15351 (N_15351,N_13421,N_13113);
and U15352 (N_15352,N_13274,N_13847);
nor U15353 (N_15353,N_14936,N_12110);
or U15354 (N_15354,N_12477,N_10856);
nor U15355 (N_15355,N_12165,N_12885);
nor U15356 (N_15356,N_14692,N_11855);
nor U15357 (N_15357,N_14988,N_14572);
and U15358 (N_15358,N_12006,N_12301);
and U15359 (N_15359,N_13165,N_14170);
nand U15360 (N_15360,N_14031,N_10804);
xor U15361 (N_15361,N_10398,N_12401);
nor U15362 (N_15362,N_12271,N_11157);
nor U15363 (N_15363,N_13793,N_14472);
nor U15364 (N_15364,N_13851,N_10818);
nand U15365 (N_15365,N_14473,N_12000);
xnor U15366 (N_15366,N_14125,N_14932);
or U15367 (N_15367,N_10018,N_14323);
or U15368 (N_15368,N_10527,N_12827);
or U15369 (N_15369,N_14012,N_13240);
or U15370 (N_15370,N_10075,N_14063);
or U15371 (N_15371,N_10558,N_14876);
nand U15372 (N_15372,N_14720,N_13483);
and U15373 (N_15373,N_11216,N_10347);
xnor U15374 (N_15374,N_12533,N_12021);
and U15375 (N_15375,N_12843,N_10884);
and U15376 (N_15376,N_11521,N_12414);
nand U15377 (N_15377,N_14369,N_12363);
or U15378 (N_15378,N_12500,N_10016);
and U15379 (N_15379,N_10500,N_12570);
xor U15380 (N_15380,N_11269,N_14548);
nor U15381 (N_15381,N_11042,N_14541);
nand U15382 (N_15382,N_10170,N_13826);
and U15383 (N_15383,N_11034,N_14344);
nand U15384 (N_15384,N_11713,N_11748);
nand U15385 (N_15385,N_11065,N_10461);
and U15386 (N_15386,N_12927,N_10089);
and U15387 (N_15387,N_14774,N_14455);
nand U15388 (N_15388,N_11305,N_11631);
and U15389 (N_15389,N_12437,N_13283);
or U15390 (N_15390,N_10068,N_14659);
and U15391 (N_15391,N_11655,N_12817);
nand U15392 (N_15392,N_10864,N_11675);
and U15393 (N_15393,N_14235,N_14380);
or U15394 (N_15394,N_13949,N_11115);
and U15395 (N_15395,N_11916,N_10538);
and U15396 (N_15396,N_12680,N_14539);
and U15397 (N_15397,N_14904,N_11499);
or U15398 (N_15398,N_12337,N_12695);
nor U15399 (N_15399,N_10152,N_14126);
and U15400 (N_15400,N_13904,N_12092);
xnor U15401 (N_15401,N_13632,N_14326);
nand U15402 (N_15402,N_11743,N_11739);
xor U15403 (N_15403,N_11428,N_10771);
nand U15404 (N_15404,N_12559,N_11716);
and U15405 (N_15405,N_13404,N_13114);
xnor U15406 (N_15406,N_11536,N_10667);
nor U15407 (N_15407,N_11697,N_10778);
and U15408 (N_15408,N_14815,N_12440);
and U15409 (N_15409,N_11938,N_13967);
nor U15410 (N_15410,N_11202,N_13155);
or U15411 (N_15411,N_13470,N_10930);
nor U15412 (N_15412,N_12675,N_12037);
xor U15413 (N_15413,N_14338,N_10777);
nor U15414 (N_15414,N_13270,N_11138);
xnor U15415 (N_15415,N_10940,N_13444);
and U15416 (N_15416,N_10231,N_14085);
nor U15417 (N_15417,N_10815,N_13051);
nand U15418 (N_15418,N_12338,N_12923);
and U15419 (N_15419,N_12050,N_11996);
xor U15420 (N_15420,N_14485,N_14223);
and U15421 (N_15421,N_10662,N_12349);
nor U15422 (N_15422,N_10259,N_12152);
and U15423 (N_15423,N_10879,N_10825);
or U15424 (N_15424,N_10209,N_10829);
nand U15425 (N_15425,N_12381,N_13798);
or U15426 (N_15426,N_12787,N_13522);
or U15427 (N_15427,N_10791,N_14714);
nor U15428 (N_15428,N_12543,N_10368);
and U15429 (N_15429,N_10429,N_13899);
xor U15430 (N_15430,N_11639,N_10665);
or U15431 (N_15431,N_12218,N_10317);
or U15432 (N_15432,N_11231,N_10325);
nand U15433 (N_15433,N_12178,N_13989);
nor U15434 (N_15434,N_11403,N_14035);
nand U15435 (N_15435,N_11228,N_12023);
nand U15436 (N_15436,N_13267,N_11929);
or U15437 (N_15437,N_11811,N_12802);
nor U15438 (N_15438,N_11997,N_12048);
or U15439 (N_15439,N_10318,N_13137);
or U15440 (N_15440,N_11879,N_12393);
or U15441 (N_15441,N_13095,N_10307);
nand U15442 (N_15442,N_11595,N_12922);
xor U15443 (N_15443,N_14414,N_10150);
xnor U15444 (N_15444,N_11911,N_12090);
xor U15445 (N_15445,N_11287,N_11906);
nor U15446 (N_15446,N_11349,N_10505);
nand U15447 (N_15447,N_14825,N_13457);
or U15448 (N_15448,N_13002,N_12800);
nor U15449 (N_15449,N_10245,N_12751);
xor U15450 (N_15450,N_11940,N_12044);
and U15451 (N_15451,N_13944,N_14746);
nor U15452 (N_15452,N_11580,N_10987);
nand U15453 (N_15453,N_12816,N_11706);
nor U15454 (N_15454,N_14303,N_13939);
xor U15455 (N_15455,N_12254,N_14688);
nor U15456 (N_15456,N_12529,N_13603);
or U15457 (N_15457,N_11377,N_12511);
or U15458 (N_15458,N_10237,N_13867);
nor U15459 (N_15459,N_13093,N_10301);
nor U15460 (N_15460,N_13800,N_14026);
xor U15461 (N_15461,N_10931,N_14144);
nor U15462 (N_15462,N_11180,N_12666);
nand U15463 (N_15463,N_13412,N_11009);
nor U15464 (N_15464,N_10487,N_13243);
xnor U15465 (N_15465,N_13666,N_14786);
and U15466 (N_15466,N_14349,N_11629);
or U15467 (N_15467,N_13107,N_11100);
nand U15468 (N_15468,N_14673,N_11208);
xnor U15469 (N_15469,N_14560,N_11053);
and U15470 (N_15470,N_14019,N_10313);
nor U15471 (N_15471,N_14438,N_13765);
xor U15472 (N_15472,N_14354,N_10303);
nor U15473 (N_15473,N_11381,N_11917);
nand U15474 (N_15474,N_14434,N_11601);
nand U15475 (N_15475,N_14024,N_14703);
nor U15476 (N_15476,N_12548,N_10880);
nor U15477 (N_15477,N_13843,N_11134);
or U15478 (N_15478,N_11136,N_12847);
or U15479 (N_15479,N_10677,N_12149);
xor U15480 (N_15480,N_12764,N_10315);
or U15481 (N_15481,N_12259,N_12891);
and U15482 (N_15482,N_14491,N_11328);
nand U15483 (N_15483,N_10962,N_12965);
xnor U15484 (N_15484,N_13735,N_14363);
and U15485 (N_15485,N_11599,N_13082);
nand U15486 (N_15486,N_13266,N_12558);
or U15487 (N_15487,N_10266,N_12307);
nor U15488 (N_15488,N_11498,N_14808);
or U15489 (N_15489,N_10071,N_14515);
nor U15490 (N_15490,N_10471,N_10642);
nor U15491 (N_15491,N_11319,N_10172);
xor U15492 (N_15492,N_12135,N_12365);
nand U15493 (N_15493,N_12607,N_14154);
nand U15494 (N_15494,N_10950,N_10035);
or U15495 (N_15495,N_11321,N_11075);
and U15496 (N_15496,N_11491,N_10122);
or U15497 (N_15497,N_13391,N_14629);
nand U15498 (N_15498,N_12008,N_12711);
nand U15499 (N_15499,N_11039,N_12697);
and U15500 (N_15500,N_11267,N_12335);
xnor U15501 (N_15501,N_13416,N_10983);
and U15502 (N_15502,N_14652,N_11664);
nand U15503 (N_15503,N_12276,N_12740);
xnor U15504 (N_15504,N_14395,N_11653);
nor U15505 (N_15505,N_13976,N_12493);
nand U15506 (N_15506,N_12539,N_11722);
xnor U15507 (N_15507,N_10694,N_13258);
and U15508 (N_15508,N_13624,N_13066);
or U15509 (N_15509,N_12192,N_10552);
or U15510 (N_15510,N_14831,N_11144);
xnor U15511 (N_15511,N_12002,N_10409);
nor U15512 (N_15512,N_11597,N_13311);
nand U15513 (N_15513,N_11455,N_10196);
xnor U15514 (N_15514,N_14439,N_11147);
nand U15515 (N_15515,N_13286,N_10578);
nand U15516 (N_15516,N_11646,N_10198);
nand U15517 (N_15517,N_10396,N_11889);
xor U15518 (N_15518,N_12114,N_11961);
nor U15519 (N_15519,N_12408,N_14225);
or U15520 (N_15520,N_14466,N_13247);
or U15521 (N_15521,N_12722,N_13235);
and U15522 (N_15522,N_11503,N_12209);
xnor U15523 (N_15523,N_11243,N_14803);
nand U15524 (N_15524,N_14578,N_11170);
and U15525 (N_15525,N_14429,N_12433);
nand U15526 (N_15526,N_14477,N_11233);
nor U15527 (N_15527,N_14467,N_13182);
or U15528 (N_15528,N_10715,N_12920);
nand U15529 (N_15529,N_14627,N_14644);
nand U15530 (N_15530,N_13564,N_14092);
or U15531 (N_15531,N_12911,N_10328);
nand U15532 (N_15532,N_14249,N_14003);
nand U15533 (N_15533,N_14129,N_10375);
xor U15534 (N_15534,N_10476,N_11059);
and U15535 (N_15535,N_14964,N_10836);
or U15536 (N_15536,N_13690,N_13731);
nand U15537 (N_15537,N_11761,N_14858);
nor U15538 (N_15538,N_14309,N_14253);
and U15539 (N_15539,N_11934,N_12566);
and U15540 (N_15540,N_11201,N_13739);
or U15541 (N_15541,N_13922,N_11280);
or U15542 (N_15542,N_14433,N_13590);
and U15543 (N_15543,N_11807,N_12481);
and U15544 (N_15544,N_13841,N_10939);
xor U15545 (N_15545,N_12483,N_10415);
nor U15546 (N_15546,N_14208,N_10986);
nor U15547 (N_15547,N_13556,N_10207);
nor U15548 (N_15548,N_12552,N_11175);
or U15549 (N_15549,N_10509,N_10894);
nand U15550 (N_15550,N_13322,N_10808);
and U15551 (N_15551,N_11797,N_14378);
or U15552 (N_15552,N_10128,N_11582);
nand U15553 (N_15553,N_11546,N_10413);
xnor U15554 (N_15554,N_10860,N_11845);
nor U15555 (N_15555,N_10819,N_11533);
or U15556 (N_15556,N_10267,N_13576);
and U15557 (N_15557,N_12774,N_12320);
nand U15558 (N_15558,N_14853,N_12485);
or U15559 (N_15559,N_11087,N_14310);
nor U15560 (N_15560,N_12475,N_14076);
nor U15561 (N_15561,N_12905,N_12084);
nand U15562 (N_15562,N_12518,N_12157);
or U15563 (N_15563,N_10062,N_12079);
nand U15564 (N_15564,N_12424,N_11975);
xnor U15565 (N_15565,N_12822,N_13685);
xnor U15566 (N_15566,N_13229,N_12611);
and U15567 (N_15567,N_14566,N_14601);
and U15568 (N_15568,N_13471,N_14348);
and U15569 (N_15569,N_10354,N_14120);
nor U15570 (N_15570,N_14186,N_12430);
or U15571 (N_15571,N_14413,N_12257);
and U15572 (N_15572,N_14581,N_10155);
nor U15573 (N_15573,N_12386,N_14277);
and U15574 (N_15574,N_11248,N_12131);
or U15575 (N_15575,N_10629,N_12102);
and U15576 (N_15576,N_10759,N_13503);
or U15577 (N_15577,N_12388,N_14694);
nor U15578 (N_15578,N_12121,N_13148);
and U15579 (N_15579,N_10425,N_14969);
and U15580 (N_15580,N_11504,N_10664);
or U15581 (N_15581,N_10027,N_12837);
xnor U15582 (N_15582,N_10699,N_13077);
or U15583 (N_15583,N_12633,N_10332);
nand U15584 (N_15584,N_10430,N_10165);
or U15585 (N_15585,N_11624,N_12583);
nand U15586 (N_15586,N_13501,N_13846);
xnor U15587 (N_15587,N_12951,N_11840);
nand U15588 (N_15588,N_14885,N_12470);
nand U15589 (N_15589,N_11999,N_14416);
nor U15590 (N_15590,N_11720,N_11676);
and U15591 (N_15591,N_12246,N_12782);
nand U15592 (N_15592,N_12499,N_11984);
xor U15593 (N_15593,N_13118,N_13909);
and U15594 (N_15594,N_13187,N_14313);
nor U15595 (N_15595,N_12959,N_11885);
xor U15596 (N_15596,N_10622,N_13752);
nor U15597 (N_15597,N_10386,N_10615);
nor U15598 (N_15598,N_14603,N_13086);
and U15599 (N_15599,N_11255,N_14897);
nor U15600 (N_15600,N_11805,N_10465);
or U15601 (N_15601,N_13869,N_14710);
nor U15602 (N_15602,N_12241,N_14006);
or U15603 (N_15603,N_12815,N_10114);
or U15604 (N_15604,N_10306,N_10350);
and U15605 (N_15605,N_14791,N_11707);
and U15606 (N_15606,N_13810,N_13417);
nor U15607 (N_15607,N_14782,N_10898);
nand U15608 (N_15608,N_12262,N_14650);
xnor U15609 (N_15609,N_13970,N_12330);
and U15610 (N_15610,N_12791,N_14625);
xnor U15611 (N_15611,N_11063,N_13030);
xor U15612 (N_15612,N_14970,N_11223);
nand U15613 (N_15613,N_14585,N_12202);
nor U15614 (N_15614,N_11406,N_12496);
and U15615 (N_15615,N_14143,N_13437);
and U15616 (N_15616,N_14955,N_12669);
and U15617 (N_15617,N_10351,N_13265);
xnor U15618 (N_15618,N_10951,N_12066);
or U15619 (N_15619,N_12898,N_13931);
nand U15620 (N_15620,N_14662,N_14863);
and U15621 (N_15621,N_13067,N_13183);
or U15622 (N_15622,N_13934,N_11303);
nand U15623 (N_15623,N_13803,N_13455);
or U15624 (N_15624,N_13566,N_11846);
or U15625 (N_15625,N_13781,N_13612);
nor U15626 (N_15626,N_11270,N_11390);
and U15627 (N_15627,N_14322,N_12845);
and U15628 (N_15628,N_13681,N_13581);
nor U15629 (N_15629,N_10673,N_14913);
nor U15630 (N_15630,N_10619,N_13245);
nor U15631 (N_15631,N_11901,N_10176);
or U15632 (N_15632,N_11083,N_14934);
and U15633 (N_15633,N_14840,N_13694);
nand U15634 (N_15634,N_11410,N_10717);
and U15635 (N_15635,N_10336,N_11438);
and U15636 (N_15636,N_13982,N_11635);
xnor U15637 (N_15637,N_14028,N_11672);
or U15638 (N_15638,N_10822,N_14228);
or U15639 (N_15639,N_12143,N_10985);
nor U15640 (N_15640,N_10256,N_10238);
and U15641 (N_15641,N_10756,N_12379);
nor U15642 (N_15642,N_14576,N_14753);
or U15643 (N_15643,N_13830,N_14972);
xor U15644 (N_15644,N_13857,N_10135);
nor U15645 (N_15645,N_10290,N_10847);
nand U15646 (N_15646,N_11557,N_10081);
or U15647 (N_15647,N_12045,N_11952);
and U15648 (N_15648,N_13657,N_12350);
nand U15649 (N_15649,N_14522,N_13838);
or U15650 (N_15650,N_14250,N_10848);
nor U15651 (N_15651,N_14191,N_12319);
xor U15652 (N_15652,N_10844,N_12305);
or U15653 (N_15653,N_14407,N_13954);
and U15654 (N_15654,N_13297,N_10323);
and U15655 (N_15655,N_12521,N_11348);
xnor U15656 (N_15656,N_10946,N_12921);
nand U15657 (N_15657,N_14593,N_12285);
and U15658 (N_15658,N_13933,N_13575);
or U15659 (N_15659,N_10314,N_10404);
nor U15660 (N_15660,N_10582,N_12723);
nand U15661 (N_15661,N_12491,N_13835);
nor U15662 (N_15662,N_11663,N_11058);
or U15663 (N_15663,N_11189,N_13463);
nand U15664 (N_15664,N_11251,N_12887);
nor U15665 (N_15665,N_13085,N_11332);
nor U15666 (N_15666,N_11737,N_12200);
nand U15667 (N_15667,N_14023,N_12028);
nand U15668 (N_15668,N_12290,N_12933);
nand U15669 (N_15669,N_14214,N_11678);
nand U15670 (N_15670,N_12644,N_11933);
xor U15671 (N_15671,N_13211,N_12101);
nor U15672 (N_15672,N_13345,N_13268);
nand U15673 (N_15673,N_13608,N_11775);
or U15674 (N_15674,N_11562,N_13096);
and U15675 (N_15675,N_10108,N_14138);
nor U15676 (N_15676,N_14701,N_14630);
nand U15677 (N_15677,N_14450,N_12132);
and U15678 (N_15678,N_10945,N_12994);
or U15679 (N_15679,N_10605,N_13374);
nor U15680 (N_15680,N_11493,N_12854);
xnor U15681 (N_15681,N_12944,N_13042);
nand U15682 (N_15682,N_14405,N_13664);
nor U15683 (N_15683,N_10868,N_10423);
nand U15684 (N_15684,N_12657,N_11081);
nand U15685 (N_15685,N_13210,N_13806);
nand U15686 (N_15686,N_11061,N_10133);
or U15687 (N_15687,N_13396,N_14854);
nor U15688 (N_15688,N_13323,N_12739);
nor U15689 (N_15689,N_14484,N_10261);
and U15690 (N_15690,N_11516,N_13589);
nor U15691 (N_15691,N_10174,N_13358);
or U15692 (N_15692,N_11780,N_14612);
nor U15693 (N_15693,N_12654,N_12977);
or U15694 (N_15694,N_14580,N_13188);
nand U15695 (N_15695,N_14112,N_13252);
nand U15696 (N_15696,N_10131,N_10472);
or U15697 (N_15697,N_12970,N_12183);
xnor U15698 (N_15698,N_11817,N_13779);
nor U15699 (N_15699,N_10807,N_13075);
nor U15700 (N_15700,N_14943,N_11041);
nand U15701 (N_15701,N_13356,N_11632);
xor U15702 (N_15702,N_10402,N_12754);
or U15703 (N_15703,N_11808,N_13400);
and U15704 (N_15704,N_11430,N_10304);
nand U15705 (N_15705,N_12034,N_13173);
xnor U15706 (N_15706,N_13535,N_12929);
xor U15707 (N_15707,N_13953,N_13023);
xor U15708 (N_15708,N_10040,N_13695);
nand U15709 (N_15709,N_10281,N_10249);
and U15710 (N_15710,N_12810,N_13972);
and U15711 (N_15711,N_11587,N_12874);
nand U15712 (N_15712,N_12120,N_14565);
and U15713 (N_15713,N_12169,N_10153);
xor U15714 (N_15714,N_12652,N_12547);
or U15715 (N_15715,N_11881,N_10004);
and U15716 (N_15716,N_14447,N_10783);
and U15717 (N_15717,N_14010,N_12284);
or U15718 (N_15718,N_13580,N_11563);
or U15719 (N_15719,N_11423,N_11825);
xor U15720 (N_15720,N_11490,N_12761);
xor U15721 (N_15721,N_10517,N_12956);
and U15722 (N_15722,N_13927,N_10335);
or U15723 (N_15723,N_12744,N_10364);
nand U15724 (N_15724,N_11072,N_10562);
xnor U15725 (N_15725,N_10210,N_13577);
nand U15726 (N_15726,N_10344,N_11777);
and U15727 (N_15727,N_12159,N_12292);
and U15728 (N_15728,N_11754,N_11329);
or U15729 (N_15729,N_13858,N_14654);
nor U15730 (N_15730,N_11970,N_12153);
nor U15731 (N_15731,N_11691,N_10992);
or U15732 (N_15732,N_12145,N_11526);
xnor U15733 (N_15733,N_10646,N_12297);
or U15734 (N_15734,N_13864,N_10349);
or U15735 (N_15735,N_14118,N_12142);
nand U15736 (N_15736,N_13407,N_13771);
xor U15737 (N_15737,N_12371,N_10980);
nand U15738 (N_15738,N_13705,N_10842);
xor U15739 (N_15739,N_11220,N_10867);
xnor U15740 (N_15740,N_14296,N_10270);
or U15741 (N_15741,N_14661,N_14282);
or U15742 (N_15742,N_10299,N_12111);
nor U15743 (N_15743,N_13343,N_13099);
or U15744 (N_15744,N_13342,N_14996);
or U15745 (N_15745,N_14933,N_11182);
xnor U15746 (N_15746,N_13418,N_10779);
xor U15747 (N_15747,N_12228,N_11173);
or U15748 (N_15748,N_14124,N_14771);
and U15749 (N_15749,N_13246,N_11448);
and U15750 (N_15750,N_11904,N_10859);
xnor U15751 (N_15751,N_13587,N_11271);
nor U15752 (N_15752,N_12745,N_10246);
or U15753 (N_15753,N_14468,N_12555);
nor U15754 (N_15754,N_11919,N_14422);
or U15755 (N_15755,N_13811,N_10881);
xnor U15756 (N_15756,N_14497,N_12795);
xnor U15757 (N_15757,N_10240,N_13500);
nor U15758 (N_15758,N_12303,N_14621);
xnor U15759 (N_15759,N_12935,N_10206);
and U15760 (N_15760,N_14660,N_14446);
nor U15761 (N_15761,N_13626,N_10714);
nand U15762 (N_15762,N_11094,N_14665);
nor U15763 (N_15763,N_11225,N_13041);
and U15764 (N_15764,N_14875,N_11401);
nand U15765 (N_15765,N_13924,N_11355);
nand U15766 (N_15766,N_11398,N_14878);
or U15767 (N_15767,N_10037,N_12762);
nand U15768 (N_15768,N_13202,N_10631);
nor U15769 (N_15769,N_13309,N_13132);
nor U15770 (N_15770,N_12604,N_13502);
or U15771 (N_15771,N_11000,N_10533);
nand U15772 (N_15772,N_10658,N_14234);
xor U15773 (N_15773,N_13651,N_14489);
or U15774 (N_15774,N_14577,N_13347);
nor U15775 (N_15775,N_11079,N_14169);
nand U15776 (N_15776,N_13956,N_10060);
nor U15777 (N_15777,N_11217,N_12598);
xor U15778 (N_15778,N_10050,N_13748);
and U15779 (N_15779,N_12252,N_10728);
nor U15780 (N_15780,N_13016,N_11586);
xnor U15781 (N_15781,N_12194,N_13383);
xor U15782 (N_15782,N_13675,N_11426);
xnor U15783 (N_15783,N_14717,N_12427);
and U15784 (N_15784,N_10236,N_12753);
nand U15785 (N_15785,N_10749,N_11454);
xnor U15786 (N_15786,N_12368,N_10262);
and U15787 (N_15787,N_10279,N_12060);
or U15788 (N_15788,N_14183,N_14174);
nor U15789 (N_15789,N_10501,N_14618);
and U15790 (N_15790,N_10479,N_14623);
nand U15791 (N_15791,N_10098,N_10008);
nor U15792 (N_15792,N_10712,N_10918);
or U15793 (N_15793,N_11979,N_13729);
nor U15794 (N_15794,N_11290,N_12639);
or U15795 (N_15795,N_12474,N_11593);
and U15796 (N_15796,N_13971,N_10077);
xnor U15797 (N_15797,N_13287,N_12040);
xnor U15798 (N_15798,N_14998,N_12075);
and U15799 (N_15799,N_14480,N_13098);
xor U15800 (N_15800,N_11331,N_14905);
nand U15801 (N_15801,N_11734,N_11571);
xnor U15802 (N_15802,N_14128,N_12690);
nand U15803 (N_15803,N_12043,N_11823);
xor U15804 (N_15804,N_13230,N_10234);
nand U15805 (N_15805,N_10327,N_11222);
or U15806 (N_15806,N_14864,N_11884);
nand U15807 (N_15807,N_13131,N_12119);
xor U15808 (N_15808,N_12168,N_12380);
xor U15809 (N_15809,N_11654,N_14524);
and U15810 (N_15810,N_12653,N_10643);
or U15811 (N_15811,N_13134,N_12046);
and U15812 (N_15812,N_12969,N_12080);
or U15813 (N_15813,N_11647,N_14212);
xor U15814 (N_15814,N_10760,N_11944);
xnor U15815 (N_15815,N_11285,N_12871);
xnor U15816 (N_15816,N_14163,N_14042);
nand U15817 (N_15817,N_14305,N_10721);
nand U15818 (N_15818,N_13866,N_12582);
nor U15819 (N_15819,N_13419,N_14428);
and U15820 (N_15820,N_13561,N_10653);
and U15821 (N_15821,N_13330,N_14132);
and U15822 (N_15822,N_12556,N_10410);
and U15823 (N_15823,N_11369,N_13415);
nor U15824 (N_15824,N_11973,N_14002);
or U15825 (N_15825,N_12136,N_12323);
nor U15826 (N_15826,N_10718,N_12390);
and U15827 (N_15827,N_10971,N_13387);
nor U15828 (N_15828,N_14361,N_14874);
nor U15829 (N_15829,N_10132,N_10949);
and U15830 (N_15830,N_10638,N_12038);
nor U15831 (N_15831,N_14819,N_12403);
or U15832 (N_15832,N_10379,N_14562);
nor U15833 (N_15833,N_11687,N_11420);
xnor U15834 (N_15834,N_13915,N_10187);
or U15835 (N_15835,N_12640,N_13061);
nand U15836 (N_15836,N_11963,N_12501);
xnor U15837 (N_15837,N_13039,N_11977);
and U15838 (N_15838,N_13993,N_14294);
nor U15839 (N_15839,N_11862,N_11447);
and U15840 (N_15840,N_14448,N_12005);
and U15841 (N_15841,N_12982,N_13472);
or U15842 (N_15842,N_10148,N_10397);
xnor U15843 (N_15843,N_13025,N_10942);
xnor U15844 (N_15844,N_13009,N_10591);
nor U15845 (N_15845,N_12863,N_14287);
and U15846 (N_15846,N_11252,N_14083);
or U15847 (N_15847,N_14776,N_12673);
or U15848 (N_15848,N_10775,N_14022);
nand U15849 (N_15849,N_11794,N_14082);
nand U15850 (N_15850,N_13656,N_13079);
or U15851 (N_15851,N_12531,N_10776);
nor U15852 (N_15852,N_11762,N_14096);
nor U15853 (N_15853,N_10999,N_12962);
and U15854 (N_15854,N_14339,N_12492);
and U15855 (N_15855,N_12322,N_14329);
nand U15856 (N_15856,N_12182,N_10208);
nor U15857 (N_15857,N_10630,N_12482);
xor U15858 (N_15858,N_12296,N_11160);
nor U15859 (N_15859,N_13637,N_12161);
nor U15860 (N_15860,N_10518,N_12926);
nand U15861 (N_15861,N_13926,N_10405);
nor U15862 (N_15862,N_10263,N_11705);
nor U15863 (N_15863,N_14465,N_14526);
and U15864 (N_15864,N_13144,N_10495);
nor U15865 (N_15865,N_13750,N_10843);
or U15866 (N_15866,N_11893,N_14563);
nand U15867 (N_15867,N_14080,N_13315);
and U15868 (N_15868,N_14247,N_14318);
nor U15869 (N_15869,N_14504,N_13379);
xor U15870 (N_15870,N_13661,N_14377);
nor U15871 (N_15871,N_10803,N_12383);
xor U15872 (N_15872,N_13020,N_10535);
and U15873 (N_15873,N_11853,N_12398);
and U15874 (N_15874,N_12519,N_10854);
nand U15875 (N_15875,N_10066,N_14521);
nor U15876 (N_15876,N_10265,N_10726);
and U15877 (N_15877,N_10747,N_11341);
xor U15878 (N_15878,N_14203,N_14511);
and U15879 (N_15879,N_10737,N_13335);
xnor U15880 (N_15880,N_14045,N_14867);
or U15881 (N_15881,N_14719,N_12938);
nand U15882 (N_15882,N_13831,N_14801);
or U15883 (N_15883,N_13233,N_10572);
xnor U15884 (N_15884,N_13121,N_12175);
nor U15885 (N_15885,N_10345,N_10781);
or U15886 (N_15886,N_12917,N_14764);
and U15887 (N_15887,N_14193,N_14523);
xor U15888 (N_15888,N_10469,N_10293);
nor U15889 (N_15889,N_10358,N_12425);
or U15890 (N_15890,N_13212,N_10746);
nand U15891 (N_15891,N_10378,N_12373);
nand U15892 (N_15892,N_10502,N_13256);
nor U15893 (N_15893,N_11728,N_12377);
or U15894 (N_15894,N_12729,N_13672);
and U15895 (N_15895,N_10813,N_10899);
xor U15896 (N_15896,N_12895,N_11528);
xor U15897 (N_15897,N_14938,N_10767);
and U15898 (N_15898,N_10443,N_11806);
xor U15899 (N_15899,N_14342,N_13968);
nor U15900 (N_15900,N_10058,N_14977);
nand U15901 (N_15901,N_12478,N_13263);
and U15902 (N_15902,N_12721,N_14332);
xnor U15903 (N_15903,N_14944,N_11689);
nor U15904 (N_15904,N_11989,N_14317);
or U15905 (N_15905,N_10698,N_13301);
nand U15906 (N_15906,N_10466,N_10690);
nand U15907 (N_15907,N_10352,N_13218);
and U15908 (N_15908,N_14647,N_11686);
or U15909 (N_15909,N_12207,N_13613);
xor U15910 (N_15910,N_12107,N_10672);
and U15911 (N_15911,N_10851,N_13257);
nor U15912 (N_15912,N_12616,N_11148);
or U15913 (N_15913,N_13294,N_10490);
and U15914 (N_15914,N_12154,N_14181);
nor U15915 (N_15915,N_13331,N_11502);
nor U15916 (N_15916,N_12300,N_10120);
and U15917 (N_15917,N_11300,N_13725);
xor U15918 (N_15918,N_14392,N_10603);
or U15919 (N_15919,N_14617,N_12625);
xor U15920 (N_15920,N_10725,N_14594);
or U15921 (N_15921,N_14039,N_14168);
nand U15922 (N_15922,N_10936,N_11357);
nor U15923 (N_15923,N_12173,N_13498);
or U15924 (N_15924,N_11930,N_10701);
nand U15925 (N_15925,N_14104,N_14721);
and U15926 (N_15926,N_12880,N_12954);
xnor U15927 (N_15927,N_11981,N_11399);
nand U15928 (N_15928,N_11594,N_13056);
or U15929 (N_15929,N_10554,N_13250);
and U15930 (N_15930,N_12643,N_13563);
or U15931 (N_15931,N_12989,N_12255);
or U15932 (N_15932,N_14788,N_11923);
xor U15933 (N_15933,N_14760,N_12508);
nand U15934 (N_15934,N_11859,N_12758);
and U15935 (N_15935,N_12019,N_13683);
and U15936 (N_15936,N_11693,N_11373);
nand U15937 (N_15937,N_12097,N_13197);
xor U15938 (N_15938,N_11486,N_11688);
and U15939 (N_15939,N_11854,N_10289);
xor U15940 (N_15940,N_12415,N_12749);
nor U15941 (N_15941,N_14817,N_11324);
nor U15942 (N_15942,N_10581,N_11764);
or U15943 (N_15943,N_12081,N_14769);
and U15944 (N_15944,N_14384,N_14048);
nand U15945 (N_15945,N_14844,N_13043);
xor U15946 (N_15946,N_13038,N_11939);
xnor U15947 (N_15947,N_11864,N_12049);
and U15948 (N_15948,N_13199,N_11320);
xnor U15949 (N_15949,N_10343,N_14589);
xnor U15950 (N_15950,N_10028,N_13991);
nand U15951 (N_15951,N_11790,N_11524);
nand U15952 (N_15952,N_13527,N_14425);
or U15953 (N_15953,N_12418,N_10929);
nand U15954 (N_15954,N_14194,N_12963);
xnor U15955 (N_15955,N_10298,N_10676);
nand U15956 (N_15956,N_12569,N_14582);
or U15957 (N_15957,N_13428,N_10534);
nor U15958 (N_15958,N_11603,N_12174);
nor U15959 (N_15959,N_12129,N_11605);
or U15960 (N_15960,N_10657,N_11476);
nand U15961 (N_15961,N_12985,N_12699);
xnor U15962 (N_15962,N_11782,N_10953);
and U15963 (N_15963,N_14009,N_11425);
nor U15964 (N_15964,N_14966,N_11732);
nor U15965 (N_15965,N_12316,N_11389);
nand U15966 (N_15966,N_12859,N_12902);
nand U15967 (N_15967,N_14567,N_10671);
nor U15968 (N_15968,N_12376,N_10445);
nand U15969 (N_15969,N_13962,N_14330);
or U15970 (N_15970,N_14843,N_14449);
nor U15971 (N_15971,N_10498,N_14824);
or U15972 (N_15972,N_10308,N_14173);
xnor U15973 (N_15973,N_11708,N_14408);
nor U15974 (N_15974,N_11340,N_12987);
xor U15975 (N_15975,N_14216,N_14909);
nand U15976 (N_15976,N_13530,N_10801);
xnor U15977 (N_15977,N_14931,N_12223);
nand U15978 (N_15978,N_13986,N_14857);
and U15979 (N_15979,N_14611,N_14820);
nand U15980 (N_15980,N_10488,N_11592);
nor U15981 (N_15981,N_14797,N_11445);
and U15982 (N_15982,N_12647,N_11346);
xor U15983 (N_15983,N_13842,N_13181);
and U15984 (N_15984,N_14382,N_11429);
xnor U15985 (N_15985,N_10526,N_12992);
nor U15986 (N_15986,N_11206,N_12432);
or U15987 (N_15987,N_14227,N_13194);
and U15988 (N_15988,N_12088,N_13289);
and U15989 (N_15989,N_13951,N_11363);
or U15990 (N_15990,N_12250,N_13013);
or U15991 (N_15991,N_10532,N_10703);
or U15992 (N_15992,N_10216,N_14908);
or U15993 (N_15993,N_14188,N_13307);
xnor U15994 (N_15994,N_11841,N_13368);
and U15995 (N_15995,N_10140,N_12930);
and U15996 (N_15996,N_14902,N_10529);
nand U15997 (N_15997,N_11986,N_10158);
and U15998 (N_15998,N_10146,N_12212);
nor U15999 (N_15999,N_14494,N_10650);
xnor U16000 (N_16000,N_12850,N_12455);
or U16001 (N_16001,N_12313,N_12190);
nor U16002 (N_16002,N_14686,N_13524);
nor U16003 (N_16003,N_13635,N_14172);
xnor U16004 (N_16004,N_14971,N_13582);
nand U16005 (N_16005,N_13942,N_10392);
and U16006 (N_16006,N_13691,N_11121);
or U16007 (N_16007,N_14040,N_13185);
or U16008 (N_16008,N_12240,N_13932);
and U16009 (N_16009,N_12270,N_11482);
nand U16010 (N_16010,N_13050,N_13269);
xnor U16011 (N_16011,N_10464,N_10036);
nand U16012 (N_16012,N_11998,N_13754);
nand U16013 (N_16013,N_14855,N_14987);
nor U16014 (N_16014,N_10764,N_11792);
xnor U16015 (N_16015,N_14544,N_13117);
xnor U16016 (N_16016,N_13541,N_10145);
or U16017 (N_16017,N_13902,N_11772);
nor U16018 (N_16018,N_10407,N_11273);
or U16019 (N_16019,N_13822,N_10784);
xnor U16020 (N_16020,N_11681,N_12855);
nor U16021 (N_16021,N_11796,N_11139);
and U16022 (N_16022,N_14321,N_11895);
or U16023 (N_16023,N_11662,N_11109);
or U16024 (N_16024,N_10503,N_14137);
nand U16025 (N_16025,N_10449,N_13119);
or U16026 (N_16026,N_12742,N_11033);
nand U16027 (N_16027,N_13442,N_10609);
or U16028 (N_16028,N_14291,N_11161);
and U16029 (N_16029,N_14704,N_10296);
nor U16030 (N_16030,N_10014,N_12813);
or U16031 (N_16031,N_10322,N_14655);
nand U16032 (N_16032,N_14624,N_13172);
xnor U16033 (N_16033,N_12266,N_12562);
nand U16034 (N_16034,N_10512,N_11957);
or U16035 (N_16035,N_14418,N_10593);
xor U16036 (N_16036,N_12984,N_13836);
or U16037 (N_16037,N_11221,N_13984);
nand U16038 (N_16038,N_13616,N_10450);
or U16039 (N_16039,N_10979,N_11992);
nand U16040 (N_16040,N_10190,N_13143);
xor U16041 (N_16041,N_14533,N_14241);
nand U16042 (N_16042,N_14341,N_11074);
xor U16043 (N_16043,N_10618,N_10943);
or U16044 (N_16044,N_13028,N_12814);
nor U16045 (N_16045,N_10724,N_10886);
xnor U16046 (N_16046,N_14981,N_11787);
or U16047 (N_16047,N_13740,N_10247);
nand U16048 (N_16048,N_11758,N_12537);
or U16049 (N_16049,N_13078,N_10613);
xor U16050 (N_16050,N_14324,N_12251);
nor U16051 (N_16051,N_10269,N_14806);
nor U16052 (N_16052,N_12950,N_13653);
or U16053 (N_16053,N_11928,N_14262);
or U16054 (N_16054,N_13948,N_14962);
nand U16055 (N_16055,N_14873,N_13462);
nand U16056 (N_16056,N_14359,N_14956);
xor U16057 (N_16057,N_13390,N_11416);
and U16058 (N_16058,N_12517,N_10668);
or U16059 (N_16059,N_13108,N_11579);
xor U16060 (N_16060,N_13196,N_14903);
nor U16061 (N_16061,N_12567,N_13985);
or U16062 (N_16062,N_10639,N_11922);
nand U16063 (N_16063,N_10356,N_14543);
or U16064 (N_16064,N_11257,N_11842);
and U16065 (N_16065,N_11779,N_13065);
or U16066 (N_16066,N_10156,N_14488);
nand U16067 (N_16067,N_10627,N_14155);
xnor U16068 (N_16068,N_11140,N_14265);
nor U16069 (N_16069,N_10934,N_10624);
xnor U16070 (N_16070,N_11104,N_13723);
xnor U16071 (N_16071,N_13116,N_10697);
and U16072 (N_16072,N_13663,N_10047);
nor U16073 (N_16073,N_14222,N_13321);
xnor U16074 (N_16074,N_11621,N_12958);
nor U16075 (N_16075,N_12186,N_10537);
xnor U16076 (N_16076,N_13059,N_11723);
nor U16077 (N_16077,N_13550,N_14004);
nand U16078 (N_16078,N_12473,N_14767);
or U16079 (N_16079,N_11110,N_11352);
or U16080 (N_16080,N_10044,N_10845);
xnor U16081 (N_16081,N_10510,N_10720);
or U16082 (N_16082,N_14116,N_13326);
nor U16083 (N_16083,N_11960,N_13929);
nand U16084 (N_16084,N_12515,N_14044);
nand U16085 (N_16085,N_11549,N_11936);
xnor U16086 (N_16086,N_10659,N_13027);
and U16087 (N_16087,N_10369,N_13170);
nand U16088 (N_16088,N_11473,N_14880);
nand U16089 (N_16089,N_11902,N_12058);
xor U16090 (N_16090,N_13721,N_10484);
or U16091 (N_16091,N_11729,N_11788);
nor U16092 (N_16092,N_10838,N_12737);
xnor U16093 (N_16093,N_10693,N_12568);
and U16094 (N_16094,N_10440,N_11912);
and U16095 (N_16095,N_14723,N_13460);
and U16096 (N_16096,N_13863,N_11768);
nand U16097 (N_16097,N_11302,N_14304);
and U16098 (N_16098,N_13870,N_11001);
nor U16099 (N_16099,N_10957,N_12488);
or U16100 (N_16100,N_12877,N_10096);
nor U16101 (N_16101,N_13159,N_13403);
nor U16102 (N_16102,N_12407,N_11518);
or U16103 (N_16103,N_14557,N_11128);
xor U16104 (N_16104,N_10385,N_13325);
xor U16105 (N_16105,N_11378,N_13491);
or U16106 (N_16106,N_14001,N_13536);
nor U16107 (N_16107,N_11622,N_11118);
nand U16108 (N_16108,N_10331,N_14761);
xor U16109 (N_16109,N_12083,N_13775);
and U16110 (N_16110,N_13224,N_10920);
or U16111 (N_16111,N_14829,N_12702);
xor U16112 (N_16112,N_11008,N_11512);
or U16113 (N_16113,N_11037,N_13213);
nand U16114 (N_16114,N_12623,N_13621);
and U16115 (N_16115,N_12247,N_10260);
nand U16116 (N_16116,N_13958,N_13823);
nand U16117 (N_16117,N_10547,N_11941);
and U16118 (N_16118,N_14165,N_12775);
or U16119 (N_16119,N_14537,N_14653);
nand U16120 (N_16120,N_12601,N_10435);
or U16121 (N_16121,N_13100,N_10227);
nand U16122 (N_16122,N_12961,N_14765);
or U16123 (N_16123,N_10978,N_11480);
xor U16124 (N_16124,N_14242,N_14417);
nor U16125 (N_16125,N_10264,N_11475);
xor U16126 (N_16126,N_13871,N_13604);
or U16127 (N_16127,N_12236,N_13878);
and U16128 (N_16128,N_13348,N_14135);
nand U16129 (N_16129,N_12670,N_13879);
nor U16130 (N_16130,N_12351,N_14814);
and U16131 (N_16131,N_13981,N_13261);
or U16132 (N_16132,N_11847,N_13055);
nor U16133 (N_16133,N_11439,N_11591);
nand U16134 (N_16134,N_12967,N_13875);
nand U16135 (N_16135,N_14509,N_13517);
xnor U16136 (N_16136,N_13112,N_13163);
and U16137 (N_16137,N_11155,N_10101);
and U16138 (N_16138,N_10168,N_12078);
nand U16139 (N_16139,N_10239,N_10849);
or U16140 (N_16140,N_10177,N_13223);
nor U16141 (N_16141,N_12820,N_14658);
nand U16142 (N_16142,N_12715,N_13001);
or U16143 (N_16143,N_13518,N_14748);
nand U16144 (N_16144,N_10486,N_14134);
and U16145 (N_16145,N_14072,N_12118);
xnor U16146 (N_16146,N_12830,N_12588);
nor U16147 (N_16147,N_10048,N_10042);
xnor U16148 (N_16148,N_10559,N_10112);
nand U16149 (N_16149,N_10889,N_11828);
nor U16150 (N_16150,N_13531,N_13276);
and U16151 (N_16151,N_14556,N_10073);
and U16152 (N_16152,N_14267,N_14891);
or U16153 (N_16153,N_13402,N_11288);
and U16154 (N_16154,N_11740,N_11370);
nand U16155 (N_16155,N_10651,N_14859);
and U16156 (N_16156,N_10941,N_10026);
nor U16157 (N_16157,N_14512,N_14054);
nand U16158 (N_16158,N_13248,N_13005);
nand U16159 (N_16159,N_14648,N_12352);
nand U16160 (N_16160,N_11238,N_13650);
nor U16161 (N_16161,N_13943,N_12400);
xnor U16162 (N_16162,N_14008,N_14441);
or U16163 (N_16163,N_13365,N_10408);
nand U16164 (N_16164,N_14153,N_11896);
xnor U16165 (N_16165,N_14887,N_10993);
nor U16166 (N_16166,N_12128,N_14513);
and U16167 (N_16167,N_12747,N_14921);
xnor U16168 (N_16168,N_14099,N_10359);
and U16169 (N_16169,N_11861,N_11982);
xnor U16170 (N_16170,N_14728,N_12329);
or U16171 (N_16171,N_13015,N_12602);
nand U16172 (N_16172,N_11218,N_11198);
or U16173 (N_16173,N_11382,N_13430);
nand U16174 (N_16174,N_12637,N_11602);
or U16175 (N_16175,N_14337,N_10252);
nand U16176 (N_16176,N_14406,N_13532);
and U16177 (N_16177,N_10181,N_11943);
nor U16178 (N_16178,N_11830,N_12869);
and U16179 (N_16179,N_10706,N_14930);
nand U16180 (N_16180,N_13316,N_10656);
nor U16181 (N_16181,N_13914,N_14570);
nand U16182 (N_16182,N_11642,N_14941);
xor U16183 (N_16183,N_11628,N_14410);
xnor U16184 (N_16184,N_14053,N_13828);
nand U16185 (N_16185,N_12861,N_12716);
or U16186 (N_16186,N_11918,N_14069);
and U16187 (N_16187,N_11442,N_12960);
nor U16188 (N_16188,N_10800,N_14239);
and U16189 (N_16189,N_10052,N_12224);
nand U16190 (N_16190,N_10291,N_13011);
nor U16191 (N_16191,N_13151,N_13175);
nand U16192 (N_16192,N_12203,N_10319);
or U16193 (N_16193,N_11529,N_13512);
and U16194 (N_16194,N_11174,N_12459);
nand U16195 (N_16195,N_14389,N_12734);
nand U16196 (N_16196,N_12571,N_14261);
or U16197 (N_16197,N_14071,N_10890);
nor U16198 (N_16198,N_13595,N_14568);
and U16199 (N_16199,N_12191,N_13973);
nor U16200 (N_16200,N_11338,N_14292);
or U16201 (N_16201,N_12219,N_12243);
nand U16202 (N_16202,N_14114,N_12879);
nor U16203 (N_16203,N_11560,N_14426);
or U16204 (N_16204,N_13426,N_14670);
xnor U16205 (N_16205,N_12343,N_10399);
xor U16206 (N_16206,N_11227,N_13649);
nor U16207 (N_16207,N_12998,N_14182);
xor U16208 (N_16208,N_14411,N_13644);
xor U16209 (N_16209,N_13054,N_11246);
or U16210 (N_16210,N_12610,N_10316);
xnor U16211 (N_16211,N_10295,N_11651);
nand U16212 (N_16212,N_12304,N_12936);
or U16213 (N_16213,N_14828,N_11964);
xor U16214 (N_16214,N_13668,N_10541);
nand U16215 (N_16215,N_13814,N_12812);
or U16216 (N_16216,N_14518,N_13572);
and U16217 (N_16217,N_11070,N_14795);
xor U16218 (N_16218,N_13908,N_10348);
and U16219 (N_16219,N_12809,N_11212);
and U16220 (N_16220,N_14984,N_10506);
xor U16221 (N_16221,N_12557,N_11795);
and U16222 (N_16222,N_13045,N_10215);
nand U16223 (N_16223,N_14105,N_11643);
xor U16224 (N_16224,N_12975,N_14218);
nor U16225 (N_16225,N_11172,N_10515);
nor U16226 (N_16226,N_13520,N_13611);
or U16227 (N_16227,N_14192,N_12799);
nand U16228 (N_16228,N_13241,N_12234);
and U16229 (N_16229,N_11213,N_12216);
nand U16230 (N_16230,N_12591,N_10991);
xnor U16231 (N_16231,N_10589,N_12014);
and U16232 (N_16232,N_13179,N_12698);
nor U16233 (N_16233,N_12314,N_14184);
nor U16234 (N_16234,N_14311,N_11937);
xor U16235 (N_16235,N_10540,N_13060);
nand U16236 (N_16236,N_12952,N_10663);
or U16237 (N_16237,N_13554,N_11517);
or U16238 (N_16238,N_10682,N_13730);
and U16239 (N_16239,N_12942,N_11925);
xnor U16240 (N_16240,N_12909,N_13458);
nand U16241 (N_16241,N_14386,N_12193);
or U16242 (N_16242,N_10069,N_14910);
xor U16243 (N_16243,N_10211,N_14269);
or U16244 (N_16244,N_10360,N_10483);
and U16245 (N_16245,N_13180,N_14860);
nand U16246 (N_16246,N_13192,N_14632);
nor U16247 (N_16247,N_13514,N_11345);
nand U16248 (N_16248,N_12897,N_14499);
or U16249 (N_16249,N_14626,N_12480);
and U16250 (N_16250,N_12177,N_10411);
and U16251 (N_16251,N_14620,N_12551);
or U16252 (N_16252,N_12724,N_12289);
and U16253 (N_16253,N_12701,N_10092);
xnor U16254 (N_16254,N_14293,N_10383);
nand U16255 (N_16255,N_13296,N_11558);
xnor U16256 (N_16256,N_13074,N_12139);
xnor U16257 (N_16257,N_13832,N_11067);
or U16258 (N_16258,N_12185,N_14032);
nor U16259 (N_16259,N_10389,N_13623);
and U16260 (N_16260,N_11102,N_11096);
nor U16261 (N_16261,N_12333,N_11283);
nor U16262 (N_16262,N_12179,N_12033);
or U16263 (N_16263,N_14752,N_12779);
xnor U16264 (N_16264,N_14676,N_10654);
nor U16265 (N_16265,N_10045,N_14616);
or U16266 (N_16266,N_14483,N_13231);
xnor U16267 (N_16267,N_12122,N_13063);
xnor U16268 (N_16268,N_10191,N_11040);
xnor U16269 (N_16269,N_13140,N_11184);
nor U16270 (N_16270,N_14121,N_13894);
or U16271 (N_16271,N_12924,N_11235);
nand U16272 (N_16272,N_14368,N_11610);
or U16273 (N_16273,N_11365,N_14059);
or U16274 (N_16274,N_12018,N_13854);
or U16275 (N_16275,N_12009,N_10064);
nor U16276 (N_16276,N_14336,N_10173);
or U16277 (N_16277,N_14350,N_14712);
or U16278 (N_16278,N_11724,N_12423);
nor U16279 (N_16279,N_10975,N_11545);
xnor U16280 (N_16280,N_12328,N_10412);
nand U16281 (N_16281,N_14495,N_11709);
nand U16282 (N_16282,N_11776,N_11987);
and U16283 (N_16283,N_11844,N_10961);
or U16284 (N_16284,N_13156,N_11910);
nand U16285 (N_16285,N_12868,N_11865);
nand U16286 (N_16286,N_14792,N_10606);
nand U16287 (N_16287,N_14850,N_11826);
and U16288 (N_16288,N_11554,N_10200);
xor U16289 (N_16289,N_13424,N_10280);
and U16290 (N_16290,N_14895,N_12785);
nor U16291 (N_16291,N_12712,N_11080);
or U16292 (N_16292,N_13000,N_14569);
or U16293 (N_16293,N_13446,N_10431);
xnor U16294 (N_16294,N_12158,N_12096);
and U16295 (N_16295,N_14784,N_13352);
xnor U16296 (N_16296,N_14394,N_11496);
nor U16297 (N_16297,N_11507,N_12007);
or U16298 (N_16298,N_12225,N_10579);
nand U16299 (N_16299,N_14596,N_10183);
xor U16300 (N_16300,N_11692,N_11483);
and U16301 (N_16301,N_12618,N_12968);
nand U16302 (N_16302,N_13558,N_10708);
nand U16303 (N_16303,N_14729,N_10865);
and U16304 (N_16304,N_13184,N_13759);
or U16305 (N_16305,N_14327,N_12725);
nor U16306 (N_16306,N_11167,N_11897);
and U16307 (N_16307,N_13646,N_10217);
and U16308 (N_16308,N_13480,N_12509);
nand U16309 (N_16309,N_13633,N_14940);
nand U16310 (N_16310,N_13542,N_10587);
or U16311 (N_16311,N_13021,N_10514);
nor U16312 (N_16312,N_12308,N_10116);
and U16313 (N_16313,N_12364,N_11700);
nor U16314 (N_16314,N_12612,N_10250);
nand U16315 (N_16315,N_13303,N_13872);
nor U16316 (N_16316,N_13277,N_12017);
and U16317 (N_16317,N_10094,N_13868);
xnor U16318 (N_16318,N_11187,N_11374);
nor U16319 (N_16319,N_10000,N_13408);
nor U16320 (N_16320,N_10115,N_14454);
and U16321 (N_16321,N_14595,N_12076);
or U16322 (N_16322,N_14000,N_13205);
nor U16323 (N_16323,N_11014,N_10548);
nand U16324 (N_16324,N_11119,N_13047);
nand U16325 (N_16325,N_12245,N_12760);
nor U16326 (N_16326,N_10223,N_12526);
or U16327 (N_16327,N_13363,N_13198);
nand U16328 (N_16328,N_10426,N_11665);
or U16329 (N_16329,N_12781,N_12873);
xor U16330 (N_16330,N_11763,N_11434);
and U16331 (N_16331,N_14830,N_14749);
or U16332 (N_16332,N_13583,N_10723);
or U16333 (N_16333,N_13792,N_11259);
nor U16334 (N_16334,N_10277,N_14949);
or U16335 (N_16335,N_11819,N_14037);
nand U16336 (N_16336,N_12067,N_14281);
nor U16337 (N_16337,N_11891,N_14101);
nor U16338 (N_16338,N_11745,N_13995);
nand U16339 (N_16339,N_13614,N_13804);
xor U16340 (N_16340,N_10895,N_10403);
nor U16341 (N_16341,N_13540,N_10998);
or U16342 (N_16342,N_11894,N_12957);
or U16343 (N_16343,N_12934,N_11117);
xor U16344 (N_16344,N_11284,N_10597);
and U16345 (N_16345,N_12991,N_10164);
or U16346 (N_16346,N_10422,N_13559);
xor U16347 (N_16347,N_10908,N_14142);
or U16348 (N_16348,N_14079,N_12689);
and U16349 (N_16349,N_12226,N_14106);
xor U16350 (N_16350,N_13432,N_10143);
nor U16351 (N_16351,N_13755,N_12389);
and U16352 (N_16352,N_11773,N_12679);
nor U16353 (N_16353,N_13850,N_13861);
xnor U16354 (N_16354,N_12807,N_12856);
nor U16355 (N_16355,N_10195,N_13693);
nand U16356 (N_16356,N_10959,N_13152);
and U16357 (N_16357,N_11821,N_11750);
xnor U16358 (N_16358,N_13753,N_14400);
or U16359 (N_16359,N_11753,N_14221);
xor U16360 (N_16360,N_10157,N_11644);
xor U16361 (N_16361,N_11666,N_12085);
nor U16362 (N_16362,N_12686,N_12996);
or U16363 (N_16363,N_12524,N_12864);
xnor U16364 (N_16364,N_13367,N_12915);
and U16365 (N_16365,N_12849,N_12918);
nand U16366 (N_16366,N_13809,N_11585);
and U16367 (N_16367,N_13618,N_12105);
nand U16368 (N_16368,N_14841,N_10730);
and U16369 (N_16369,N_10390,N_10493);
or U16370 (N_16370,N_10922,N_13560);
and U16371 (N_16371,N_14935,N_12268);
or U16372 (N_16372,N_13736,N_12858);
and U16373 (N_16373,N_12780,N_12925);
nand U16374 (N_16374,N_14109,N_10901);
or U16375 (N_16375,N_10419,N_11047);
or U16376 (N_16376,N_12439,N_11415);
xnor U16377 (N_16377,N_12731,N_12180);
or U16378 (N_16378,N_12089,N_13434);
nand U16379 (N_16379,N_10338,N_12031);
nand U16380 (N_16380,N_13488,N_11099);
nor U16381 (N_16381,N_13111,N_10006);
and U16382 (N_16382,N_12013,N_11466);
nor U16383 (N_16383,N_14807,N_11791);
or U16384 (N_16384,N_10468,N_12293);
or U16385 (N_16385,N_10119,N_13598);
nand U16386 (N_16386,N_12310,N_11030);
and U16387 (N_16387,N_13493,N_13272);
xor U16388 (N_16388,N_11127,N_14818);
nor U16389 (N_16389,N_10565,N_11863);
nand U16390 (N_16390,N_13925,N_14982);
nand U16391 (N_16391,N_10400,N_12282);
or U16392 (N_16392,N_14285,N_13346);
or U16393 (N_16393,N_12372,N_14238);
nor U16394 (N_16394,N_13496,N_10577);
and U16395 (N_16395,N_11265,N_10752);
and U16396 (N_16396,N_12072,N_10976);
nor U16397 (N_16397,N_11089,N_13219);
xnor U16398 (N_16398,N_14431,N_11615);
or U16399 (N_16399,N_13049,N_11566);
xor U16400 (N_16400,N_12141,N_11920);
nand U16401 (N_16401,N_10377,N_12466);
nand U16402 (N_16402,N_11017,N_12889);
nor U16403 (N_16403,N_12339,N_12777);
nor U16404 (N_16404,N_13420,N_12797);
and U16405 (N_16405,N_10926,N_14671);
nand U16406 (N_16406,N_11673,N_10324);
nor U16407 (N_16407,N_11942,N_14346);
nor U16408 (N_16408,N_11129,N_11905);
or U16409 (N_16409,N_13435,N_12678);
xnor U16410 (N_16410,N_11036,N_10221);
nor U16411 (N_16411,N_12708,N_10420);
nor U16412 (N_16412,N_12993,N_10984);
nand U16413 (N_16413,N_14301,N_12746);
nor U16414 (N_16414,N_13094,N_12901);
or U16415 (N_16415,N_11003,N_12890);
and U16416 (N_16416,N_11367,N_13203);
xnor U16417 (N_16417,N_14047,N_10055);
nor U16418 (N_16418,N_12981,N_11519);
nor U16419 (N_16419,N_14979,N_11282);
nand U16420 (N_16420,N_10162,N_10696);
nor U16421 (N_16421,N_11376,N_13154);
or U16422 (N_16422,N_11822,N_12651);
nor U16423 (N_16423,N_13568,N_10913);
and U16424 (N_16424,N_12575,N_10628);
xnor U16425 (N_16425,N_12789,N_11583);
xnor U16426 (N_16426,N_14233,N_13667);
and U16427 (N_16427,N_13242,N_14763);
xor U16428 (N_16428,N_14622,N_13127);
or U16429 (N_16429,N_12659,N_13332);
nand U16430 (N_16430,N_14790,N_13677);
nand U16431 (N_16431,N_12683,N_14476);
nand U16432 (N_16432,N_10086,N_14978);
and U16433 (N_16433,N_10056,N_12201);
or U16434 (N_16434,N_10382,N_10166);
or U16435 (N_16435,N_13946,N_12068);
and U16436 (N_16436,N_11395,N_11538);
xnor U16437 (N_16437,N_11253,N_13671);
nand U16438 (N_16438,N_12069,N_14052);
nor U16439 (N_16439,N_14381,N_12239);
xnor U16440 (N_16440,N_12971,N_13699);
xor U16441 (N_16441,N_11141,N_14619);
and U16442 (N_16442,N_14487,N_12870);
xor U16443 (N_16443,N_10041,N_12603);
or U16444 (N_16444,N_11277,N_11510);
nor U16445 (N_16445,N_13920,N_12645);
xor U16446 (N_16446,N_11460,N_11307);
nor U16447 (N_16447,N_13171,N_14957);
nor U16448 (N_16448,N_10015,N_14147);
and U16449 (N_16449,N_14992,N_10300);
nand U16450 (N_16450,N_12113,N_10100);
nand U16451 (N_16451,N_12233,N_12042);
nand U16452 (N_16452,N_14178,N_11312);
nor U16453 (N_16453,N_10683,N_12750);
or U16454 (N_16454,N_11715,N_11813);
nor U16455 (N_16455,N_11508,N_13006);
nor U16456 (N_16456,N_12790,N_10054);
nor U16457 (N_16457,N_14587,N_14681);
or U16458 (N_16458,N_10965,N_13713);
xnor U16459 (N_16459,N_10111,N_10126);
or U16460 (N_16460,N_14613,N_10388);
nor U16461 (N_16461,N_14157,N_14679);
xor U16462 (N_16462,N_11611,N_12004);
or U16463 (N_16463,N_13549,N_13761);
and U16464 (N_16464,N_10871,N_13588);
xnor U16465 (N_16465,N_12685,N_13945);
and U16466 (N_16466,N_13459,N_11913);
xnor U16467 (N_16467,N_12572,N_14196);
and U16468 (N_16468,N_11871,N_10686);
xor U16469 (N_16469,N_14762,N_10192);
or U16470 (N_16470,N_12642,N_10273);
and U16471 (N_16471,N_13537,N_12546);
nor U16472 (N_16472,N_11506,N_12808);
nand U16473 (N_16473,N_12053,N_11149);
or U16474 (N_16474,N_12457,N_10220);
and U16475 (N_16475,N_14783,N_10956);
and U16476 (N_16476,N_12220,N_13905);
nand U16477 (N_16477,N_12801,N_11449);
and U16478 (N_16478,N_13445,N_14427);
nand U16479 (N_16479,N_12117,N_12070);
nor U16480 (N_16480,N_10367,N_10049);
xor U16481 (N_16481,N_13724,N_14845);
nand U16482 (N_16482,N_11670,N_10788);
nor U16483 (N_16483,N_13153,N_13328);
nand U16484 (N_16484,N_13912,N_13992);
nand U16485 (N_16485,N_14098,N_13957);
or U16486 (N_16486,N_12392,N_10011);
or U16487 (N_16487,N_13936,N_11757);
nand U16488 (N_16488,N_14879,N_10905);
nand U16489 (N_16489,N_13124,N_14906);
or U16490 (N_16490,N_14508,N_10366);
and U16491 (N_16491,N_12116,N_10441);
and U16492 (N_16492,N_13876,N_10966);
or U16493 (N_16493,N_12378,N_12528);
and U16494 (N_16494,N_11318,N_13306);
xor U16495 (N_16495,N_14070,N_12456);
nand U16496 (N_16496,N_14759,N_11409);
nor U16497 (N_16497,N_10107,N_10105);
xor U16498 (N_16498,N_10550,N_14530);
xnor U16499 (N_16499,N_14687,N_10219);
nor U16500 (N_16500,N_11038,N_10897);
or U16501 (N_16501,N_14849,N_12375);
and U16502 (N_16502,N_10711,N_14215);
nand U16503 (N_16503,N_11232,N_10184);
and U16504 (N_16504,N_13037,N_11683);
nand U16505 (N_16505,N_10569,N_10870);
or U16506 (N_16506,N_12767,N_14699);
nor U16507 (N_16507,N_10147,N_13745);
or U16508 (N_16508,N_11898,N_11056);
or U16509 (N_16509,N_10907,N_14571);
or U16510 (N_16510,N_10070,N_10007);
and U16511 (N_16511,N_10302,N_11055);
xor U16512 (N_16512,N_13636,N_10795);
and U16513 (N_16513,N_11195,N_10768);
nor U16514 (N_16514,N_10608,N_14816);
or U16515 (N_16515,N_13489,N_13166);
and U16516 (N_16516,N_10713,N_11892);
xnor U16517 (N_16517,N_13024,N_10852);
nand U16518 (N_16518,N_12605,N_14060);
and U16519 (N_16519,N_11588,N_14827);
or U16520 (N_16520,N_13764,N_11668);
nand U16521 (N_16521,N_13150,N_14599);
xnor U16522 (N_16522,N_12878,N_11470);
or U16523 (N_16523,N_11584,N_14822);
and U16524 (N_16524,N_13714,N_11166);
or U16525 (N_16525,N_12672,N_14835);
and U16526 (N_16526,N_12655,N_10874);
xor U16527 (N_16527,N_12062,N_12450);
or U16528 (N_16528,N_11694,N_12972);
or U16529 (N_16529,N_13805,N_13799);
and U16530 (N_16530,N_12589,N_11366);
and U16531 (N_16531,N_14136,N_10614);
xor U16532 (N_16532,N_12600,N_14207);
and U16533 (N_16533,N_14090,N_10276);
and U16534 (N_16534,N_13597,N_11511);
or U16535 (N_16535,N_10271,N_11721);
or U16536 (N_16536,N_11256,N_10833);
xnor U16537 (N_16537,N_10575,N_12819);
nand U16538 (N_16538,N_14122,N_13712);
nand U16539 (N_16539,N_12095,N_10104);
or U16540 (N_16540,N_12629,N_10212);
nor U16541 (N_16541,N_13570,N_11296);
or U16542 (N_16542,N_14811,N_14100);
or U16543 (N_16543,N_11802,N_13639);
xor U16544 (N_16544,N_12106,N_14027);
nand U16545 (N_16545,N_14899,N_11468);
nand U16546 (N_16546,N_11576,N_13344);
nand U16547 (N_16547,N_11336,N_11095);
and U16548 (N_16548,N_10734,N_13678);
xor U16549 (N_16549,N_11559,N_14379);
nor U16550 (N_16550,N_13353,N_10994);
and U16551 (N_16551,N_13441,N_12544);
nor U16552 (N_16552,N_10320,N_11116);
nor U16553 (N_16553,N_11914,N_14973);
nand U16554 (N_16554,N_14113,N_13447);
or U16555 (N_16555,N_12140,N_11784);
and U16556 (N_16556,N_13468,N_14470);
nor U16557 (N_16557,N_12649,N_12943);
xnor U16558 (N_16558,N_13433,N_12299);
nand U16559 (N_16559,N_13708,N_14399);
or U16560 (N_16560,N_14127,N_14775);
nand U16561 (N_16561,N_12677,N_10738);
nand U16562 (N_16562,N_12054,N_13125);
or U16563 (N_16563,N_13411,N_14308);
and U16564 (N_16564,N_10826,N_12741);
nor U16565 (N_16565,N_13186,N_10091);
xor U16566 (N_16566,N_12832,N_13281);
nor U16567 (N_16567,N_12886,N_10661);
or U16568 (N_16568,N_10329,N_10009);
nor U16569 (N_16569,N_11552,N_12903);
nand U16570 (N_16570,N_14968,N_14254);
nand U16571 (N_16571,N_10002,N_11868);
xnor U16572 (N_16572,N_14800,N_10522);
nor U16573 (N_16573,N_12086,N_14498);
nand U16574 (N_16574,N_13538,N_11570);
nand U16575 (N_16575,N_10566,N_11474);
xor U16576 (N_16576,N_10902,N_10432);
and U16577 (N_16577,N_14271,N_12272);
and U16578 (N_16578,N_10284,N_11733);
nor U16579 (N_16579,N_13495,N_13482);
or U16580 (N_16580,N_12765,N_14278);
xor U16581 (N_16581,N_14744,N_13485);
and U16582 (N_16582,N_11617,N_13950);
nand U16583 (N_16583,N_13251,N_13955);
nor U16584 (N_16584,N_11965,N_14462);
xor U16585 (N_16585,N_10812,N_10059);
nand U16586 (N_16586,N_10641,N_13890);
and U16587 (N_16587,N_12522,N_12634);
and U16588 (N_16588,N_11903,N_11703);
or U16589 (N_16589,N_12026,N_10678);
nor U16590 (N_16590,N_10551,N_10877);
nor U16591 (N_16591,N_14638,N_14297);
and U16592 (N_16592,N_12283,N_13262);
xnor U16593 (N_16593,N_10634,N_12130);
nor U16594 (N_16594,N_10457,N_14961);
nor U16595 (N_16595,N_14994,N_10679);
or U16596 (N_16596,N_12001,N_13478);
or U16597 (N_16597,N_13141,N_12336);
nand U16598 (N_16598,N_10199,N_11857);
xnor U16599 (N_16599,N_13069,N_10660);
xor U16600 (N_16600,N_10201,N_10850);
xor U16601 (N_16601,N_12232,N_10602);
xor U16602 (N_16602,N_14872,N_13602);
nor U16603 (N_16603,N_12495,N_10167);
nand U16604 (N_16604,N_11171,N_11107);
xor U16605 (N_16605,N_10519,N_11162);
nor U16606 (N_16606,N_11177,N_14316);
or U16607 (N_16607,N_12098,N_13769);
or U16608 (N_16608,N_10896,N_14325);
nand U16609 (N_16609,N_11674,N_12279);
or U16610 (N_16610,N_13742,N_11974);
nand U16611 (N_16611,N_12860,N_13088);
nand U16612 (N_16612,N_14280,N_12147);
xnor U16613 (N_16613,N_11086,N_12818);
nor U16614 (N_16614,N_11837,N_14077);
nor U16615 (N_16615,N_11301,N_13782);
xnor U16616 (N_16616,N_13168,N_13606);
or U16617 (N_16617,N_11178,N_10839);
and U16618 (N_16618,N_12727,N_14507);
and U16619 (N_16619,N_13528,N_10882);
nand U16620 (N_16620,N_13670,N_11744);
xor U16621 (N_16621,N_10189,N_14351);
xnor U16622 (N_16622,N_10473,N_13217);
nand U16623 (N_16623,N_14471,N_10729);
xnor U16624 (N_16624,N_11690,N_10275);
or U16625 (N_16625,N_13634,N_12467);
xnor U16626 (N_16626,N_11022,N_10373);
or U16627 (N_16627,N_11614,N_10283);
nor U16628 (N_16628,N_11274,N_11424);
and U16629 (N_16629,N_13160,N_10731);
or U16630 (N_16630,N_14756,N_11569);
and U16631 (N_16631,N_11718,N_12700);
xnor U16632 (N_16632,N_10370,N_12318);
or U16633 (N_16633,N_11781,N_13285);
nand U16634 (N_16634,N_12332,N_12431);
or U16635 (N_16635,N_11467,N_11852);
nor U16636 (N_16636,N_10480,N_13333);
or U16637 (N_16637,N_11297,N_13607);
and U16638 (N_16638,N_10376,N_13543);
nand U16639 (N_16639,N_14201,N_13359);
nand U16640 (N_16640,N_14698,N_13410);
nand U16641 (N_16641,N_11379,N_14725);
or U16642 (N_16642,N_14669,N_12743);
or U16643 (N_16643,N_11343,N_12614);
nor U16644 (N_16644,N_14020,N_14545);
or U16645 (N_16645,N_14689,N_10688);
nand U16646 (N_16646,N_11441,N_12949);
nand U16647 (N_16647,N_14643,N_10762);
nor U16648 (N_16648,N_12882,N_13921);
nand U16649 (N_16649,N_12244,N_10421);
xnor U16650 (N_16650,N_12321,N_13523);
and U16651 (N_16651,N_10840,N_14592);
xnor U16652 (N_16652,N_10689,N_10640);
and U16653 (N_16653,N_11606,N_12353);
nor U16654 (N_16654,N_11980,N_10163);
nor U16655 (N_16655,N_14312,N_12162);
nor U16656 (N_16656,N_14722,N_10787);
nand U16657 (N_16657,N_10600,N_14333);
and U16658 (N_16658,N_10292,N_11836);
nor U16659 (N_16659,N_11315,N_10287);
nand U16660 (N_16660,N_14551,N_13913);
nor U16661 (N_16661,N_12732,N_13918);
or U16662 (N_16662,N_12823,N_13655);
or U16663 (N_16663,N_12104,N_14274);
nor U16664 (N_16664,N_13784,N_11860);
or U16665 (N_16665,N_13370,N_13362);
nand U16666 (N_16666,N_13605,N_10564);
or U16667 (N_16667,N_14989,N_11230);
nand U16668 (N_16668,N_14547,N_12156);
nand U16669 (N_16669,N_12199,N_13479);
nand U16670 (N_16670,N_11574,N_11035);
or U16671 (N_16671,N_10078,N_10705);
and U16672 (N_16672,N_14319,N_12016);
nand U16673 (N_16673,N_11858,N_12260);
or U16674 (N_16674,N_14946,N_13630);
nand U16675 (N_16675,N_12317,N_14675);
nand U16676 (N_16676,N_11921,N_11152);
xnor U16677 (N_16677,N_11626,N_12565);
xnor U16678 (N_16678,N_10652,N_12273);
nor U16679 (N_16679,N_11555,N_11408);
nor U16680 (N_16680,N_13586,N_14901);
nor U16681 (N_16681,N_10099,N_10988);
xnor U16682 (N_16682,N_11513,N_12265);
nand U16683 (N_16683,N_14837,N_11541);
or U16684 (N_16684,N_13896,N_10130);
nor U16685 (N_16685,N_14156,N_11145);
nor U16686 (N_16686,N_11751,N_12593);
xnor U16687 (N_16687,N_13599,N_13625);
nand U16688 (N_16688,N_13035,N_13139);
and U16689 (N_16689,N_10824,N_14804);
xor U16690 (N_16690,N_14402,N_13409);
and U16691 (N_16691,N_11237,N_10171);
and U16692 (N_16692,N_10751,N_12828);
xor U16693 (N_16693,N_10039,N_12249);
or U16694 (N_16694,N_14005,N_11049);
nand U16695 (N_16695,N_11785,N_11266);
nor U16696 (N_16696,N_10669,N_11604);
nor U16697 (N_16697,N_13711,N_10633);
or U16698 (N_16698,N_12940,N_13702);
nand U16699 (N_16699,N_12821,N_11375);
xor U16700 (N_16700,N_11019,N_14066);
nor U16701 (N_16701,N_12595,N_10647);
and U16702 (N_16702,N_10924,N_11358);
or U16703 (N_16703,N_11402,N_11122);
xor U16704 (N_16704,N_10357,N_13965);
and U16705 (N_16705,N_12973,N_10586);
and U16706 (N_16706,N_11021,N_14390);
or U16707 (N_16707,N_14674,N_11575);
nor U16708 (N_16708,N_13884,N_11043);
and U16709 (N_16709,N_13405,N_11418);
nand U16710 (N_16710,N_13083,N_10912);
nand U16711 (N_16711,N_13336,N_13797);
or U16712 (N_16712,N_14478,N_12506);
nor U16713 (N_16713,N_12134,N_14094);
nor U16714 (N_16714,N_13895,N_10911);
nor U16715 (N_16715,N_10626,N_13573);
nor U16716 (N_16716,N_11143,N_10387);
nor U16717 (N_16717,N_10330,N_13302);
or U16718 (N_16718,N_13709,N_12585);
nor U16719 (N_16719,N_13855,N_10782);
xor U16720 (N_16720,N_12148,N_12227);
and U16721 (N_16721,N_13436,N_11887);
and U16722 (N_16722,N_10232,N_10401);
or U16723 (N_16723,N_12624,N_12486);
and U16724 (N_16724,N_11254,N_10030);
and U16725 (N_16725,N_12768,N_12434);
and U16726 (N_16726,N_11497,N_10611);
xnor U16727 (N_16727,N_12664,N_10933);
nor U16728 (N_16728,N_12248,N_14288);
xor U16729 (N_16729,N_12881,N_13717);
nor U16730 (N_16730,N_13357,N_12796);
xor U16731 (N_16731,N_13829,N_13539);
nor U16732 (N_16732,N_11188,N_14460);
or U16733 (N_16733,N_11947,N_12834);
nand U16734 (N_16734,N_13704,N_11186);
nor U16735 (N_16735,N_14740,N_12833);
nand U16736 (N_16736,N_13629,N_11875);
and U16737 (N_16737,N_10197,N_11596);
or U16738 (N_16738,N_13174,N_11641);
and U16739 (N_16739,N_14252,N_13856);
nand U16740 (N_16740,N_12836,N_10592);
nor U16741 (N_16741,N_10182,N_11204);
or U16742 (N_16742,N_14334,N_11814);
nor U16743 (N_16743,N_14600,N_14534);
nand U16744 (N_16744,N_10257,N_11435);
or U16745 (N_16745,N_13526,N_13214);
or U16746 (N_16746,N_13373,N_13072);
and U16747 (N_16747,N_14754,N_10032);
nand U16748 (N_16748,N_11949,N_11543);
or U16749 (N_16749,N_11874,N_12027);
and U16750 (N_16750,N_12893,N_13227);
and U16751 (N_16751,N_14482,N_12752);
xnor U16752 (N_16752,N_11436,N_12170);
nand U16753 (N_16753,N_14246,N_14634);
and U16754 (N_16754,N_14391,N_13126);
or U16755 (N_16755,N_12824,N_10139);
or U16756 (N_16756,N_11431,N_14965);
xnor U16757 (N_16757,N_13578,N_13980);
nand U16758 (N_16758,N_12342,N_14496);
and U16759 (N_16759,N_11867,N_14371);
nand U16760 (N_16760,N_10914,N_14766);
nor U16761 (N_16761,N_11544,N_13046);
nand U16762 (N_16762,N_14437,N_10496);
xnor U16763 (N_16763,N_13355,N_14883);
and U16764 (N_16764,N_10012,N_14140);
nor U16765 (N_16765,N_14206,N_11680);
nor U16766 (N_16766,N_12904,N_12206);
xnor U16767 (N_16767,N_11548,N_10065);
or U16768 (N_16768,N_11481,N_13785);
and U16769 (N_16769,N_11278,N_12237);
nor U16770 (N_16770,N_14209,N_14706);
nand U16771 (N_16771,N_12707,N_11091);
or U16772 (N_16772,N_11809,N_14871);
nand U16773 (N_16773,N_11878,N_10741);
xor U16774 (N_16774,N_10097,N_12580);
and U16775 (N_16775,N_13622,N_10470);
xnor U16776 (N_16776,N_11193,N_13974);
nor U16777 (N_16777,N_13988,N_11660);
or U16778 (N_16778,N_11190,N_14889);
nor U16779 (N_16779,N_14925,N_11207);
xnor U16780 (N_16780,N_10363,N_12464);
xnor U16781 (N_16781,N_13553,N_14167);
and U16782 (N_16782,N_11612,N_11534);
xnor U16783 (N_16783,N_10202,N_14016);
xor U16784 (N_16784,N_14078,N_11371);
xor U16785 (N_16785,N_13206,N_12691);
xnor U16786 (N_16786,N_10372,N_14286);
nor U16787 (N_16787,N_13384,N_11215);
or U16788 (N_16788,N_11578,N_10492);
or U16789 (N_16789,N_14583,N_11356);
nand U16790 (N_16790,N_12399,N_11827);
nand U16791 (N_16791,N_12356,N_13029);
nor U16792 (N_16792,N_11472,N_12646);
nor U16793 (N_16793,N_14967,N_10948);
and U16794 (N_16794,N_14370,N_14061);
or U16795 (N_16795,N_13916,N_10625);
xor U16796 (N_16796,N_14366,N_14018);
nand U16797 (N_16797,N_12238,N_10242);
and U16798 (N_16798,N_11294,N_12123);
xor U16799 (N_16799,N_13305,N_12438);
nor U16800 (N_16800,N_10758,N_14198);
nand U16801 (N_16801,N_13897,N_11684);
nand U16802 (N_16802,N_12326,N_10205);
nand U16803 (N_16803,N_14064,N_10159);
and U16804 (N_16804,N_14502,N_13643);
nor U16805 (N_16805,N_14300,N_11640);
nor U16806 (N_16806,N_13654,N_12138);
xor U16807 (N_16807,N_12846,N_14951);
or U16808 (N_16808,N_11619,N_12413);
nor U16809 (N_16809,N_13064,N_12253);
and U16810 (N_16810,N_14290,N_14299);
and U16811 (N_16811,N_10474,N_14403);
or U16812 (N_16812,N_12311,N_11456);
nand U16813 (N_16813,N_12704,N_11405);
xnor U16814 (N_16814,N_14179,N_14697);
xor U16815 (N_16815,N_12288,N_14916);
nor U16816 (N_16816,N_11711,N_14954);
xor U16817 (N_16817,N_12709,N_10707);
xnor U16818 (N_16818,N_12230,N_10919);
nor U16819 (N_16819,N_12710,N_11657);
nor U16820 (N_16820,N_11011,N_10090);
xnor U16821 (N_16821,N_10831,N_13776);
nand U16822 (N_16822,N_12047,N_10967);
xor U16823 (N_16823,N_10745,N_11211);
and U16824 (N_16824,N_13780,N_10561);
nand U16825 (N_16825,N_12784,N_11539);
nor U16826 (N_16826,N_14812,N_11667);
nor U16827 (N_16827,N_12573,N_12435);
or U16828 (N_16828,N_14073,N_10798);
or U16829 (N_16829,N_12794,N_12057);
and U16830 (N_16830,N_13652,N_12215);
xnor U16831 (N_16831,N_13880,N_11146);
xnor U16832 (N_16832,N_13228,N_12590);
nand U16833 (N_16833,N_14549,N_14240);
xnor U16834 (N_16834,N_10681,N_11677);
xor U16835 (N_16835,N_14542,N_11350);
or U16836 (N_16836,N_11489,N_14266);
and U16837 (N_16837,N_14145,N_10765);
and U16838 (N_16838,N_11281,N_10869);
nand U16839 (N_16839,N_10229,N_12137);
nor U16840 (N_16840,N_12883,N_13115);
nor U16841 (N_16841,N_13930,N_12912);
nor U16842 (N_16842,N_11698,N_10427);
xor U16843 (N_16843,N_12074,N_11789);
nor U16844 (N_16844,N_10282,N_10326);
xor U16845 (N_16845,N_13157,N_12460);
or U16846 (N_16846,N_12446,N_14693);
nor U16847 (N_16847,N_13448,N_14340);
nand U16848 (N_16848,N_12497,N_12184);
or U16849 (N_16849,N_13146,N_13658);
xor U16850 (N_16850,N_14486,N_14607);
xnor U16851 (N_16851,N_14527,N_10748);
and U16852 (N_16852,N_14742,N_12195);
xor U16853 (N_16853,N_11051,N_14525);
nor U16854 (N_16854,N_13979,N_11103);
and U16855 (N_16855,N_13874,N_13062);
and U16856 (N_16856,N_14865,N_11627);
xnor U16857 (N_16857,N_10416,N_13161);
xnor U16858 (N_16858,N_14058,N_12109);
or U16859 (N_16859,N_13386,N_11093);
nand U16860 (N_16860,N_12632,N_11421);
and U16861 (N_16861,N_14870,N_11550);
or U16862 (N_16862,N_10968,N_11824);
nor U16863 (N_16863,N_12884,N_13034);
nor U16864 (N_16864,N_11945,N_14713);
and U16865 (N_16865,N_11985,N_12842);
xnor U16866 (N_16866,N_11446,N_12445);
nand U16867 (N_16867,N_11831,N_10087);
and U16868 (N_16868,N_11309,N_14180);
or U16869 (N_16869,N_10029,N_13881);
nor U16870 (N_16870,N_14373,N_14554);
or U16871 (N_16871,N_11105,N_13022);
or U16872 (N_16872,N_13058,N_14975);
nand U16873 (N_16873,N_11725,N_14065);
and U16874 (N_16874,N_10452,N_10754);
xnor U16875 (N_16875,N_11272,N_13592);
nand U16876 (N_16876,N_11669,N_11214);
nor U16877 (N_16877,N_11015,N_12065);
xnor U16878 (N_16878,N_13574,N_12024);
nor U16879 (N_16879,N_10513,N_10621);
nor U16880 (N_16880,N_12899,N_12100);
nand U16881 (N_16881,N_12554,N_10046);
nor U16882 (N_16882,N_13017,N_12187);
nand U16883 (N_16883,N_12536,N_11701);
and U16884 (N_16884,N_10499,N_14131);
or U16885 (N_16885,N_10127,N_13486);
xnor U16886 (N_16886,N_14195,N_13888);
nand U16887 (N_16887,N_13080,N_14396);
nor U16888 (N_16888,N_10491,N_11567);
nor U16889 (N_16889,N_13515,N_11244);
and U16890 (N_16890,N_10218,N_10861);
or U16891 (N_16891,N_10862,N_14922);
nand U16892 (N_16892,N_10974,N_11351);
and U16893 (N_16893,N_10887,N_12713);
xnor U16894 (N_16894,N_14328,N_13848);
nor U16895 (N_16895,N_13964,N_12999);
or U16896 (N_16896,N_14424,N_11531);
nor U16897 (N_16897,N_14894,N_13648);
or U16898 (N_16898,N_11500,N_10796);
or U16899 (N_16899,N_13273,N_14770);
or U16900 (N_16900,N_14151,N_11450);
or U16901 (N_16901,N_10958,N_13004);
or U16902 (N_16902,N_12402,N_12995);
xor U16903 (N_16903,N_11126,N_13249);
nor U16904 (N_16904,N_11856,N_11873);
nor U16905 (N_16905,N_14177,N_14500);
xnor U16906 (N_16906,N_14777,N_10080);
or U16907 (N_16907,N_13097,N_10137);
and U16908 (N_16908,N_13282,N_12384);
nand U16909 (N_16909,N_10253,N_13176);
and U16910 (N_16910,N_11747,N_12592);
and U16911 (N_16911,N_12295,N_14375);
nor U16912 (N_16912,N_11101,N_13642);
and U16913 (N_16913,N_11032,N_13244);
xor U16914 (N_16914,N_14914,N_14190);
and U16915 (N_16915,N_14217,N_10341);
and U16916 (N_16916,N_13073,N_13783);
xnor U16917 (N_16917,N_11671,N_11050);
nand U16918 (N_16918,N_13701,N_11572);
nand U16919 (N_16919,N_11066,N_12217);
or U16920 (N_16920,N_12939,N_13354);
nor U16921 (N_16921,N_14823,N_14347);
or U16922 (N_16922,N_14695,N_12387);
or U16923 (N_16923,N_11322,N_11926);
or U16924 (N_16924,N_10636,N_14772);
or U16925 (N_16925,N_14115,N_13385);
nand U16926 (N_16926,N_12835,N_10203);
xor U16927 (N_16927,N_14730,N_14896);
or U16928 (N_16928,N_13312,N_13862);
xnor U16929 (N_16929,N_14503,N_13136);
nand U16930 (N_16930,N_12302,N_14579);
xor U16931 (N_16931,N_14750,N_11736);
or U16932 (N_16932,N_10161,N_12022);
nand U16933 (N_16933,N_13089,N_13813);
nor U16934 (N_16934,N_10837,N_13978);
xnor U16935 (N_16935,N_10123,N_12235);
nor U16936 (N_16936,N_10458,N_13631);
and U16937 (N_16937,N_11150,N_11710);
xor U16938 (N_16938,N_14656,N_10477);
nand U16939 (N_16939,N_11459,N_11111);
or U16940 (N_16940,N_12374,N_11971);
nor U16941 (N_16941,N_12719,N_13794);
and U16942 (N_16942,N_13893,N_13891);
nor U16943 (N_16943,N_14546,N_14243);
or U16944 (N_16944,N_10455,N_13700);
nor U16945 (N_16945,N_13044,N_11804);
xnor U16946 (N_16946,N_11306,N_12841);
or U16947 (N_16947,N_14166,N_14062);
and U16948 (N_16948,N_13778,N_10736);
or U16949 (N_16949,N_10598,N_12448);
nand U16950 (N_16950,N_14724,N_11530);
nor U16951 (N_16951,N_11354,N_14091);
nand U16952 (N_16952,N_13222,N_12534);
and U16953 (N_16953,N_12405,N_11909);
or U16954 (N_16954,N_13766,N_13593);
or U16955 (N_16955,N_10395,N_10743);
or U16956 (N_16956,N_12325,N_12281);
xnor U16957 (N_16957,N_11325,N_12073);
xnor U16958 (N_16958,N_14898,N_13529);
nand U16959 (N_16959,N_13544,N_14161);
nand U16960 (N_16960,N_14036,N_14213);
and U16961 (N_16961,N_11339,N_12755);
nand U16962 (N_16962,N_10691,N_13236);
nand U16963 (N_16963,N_11247,N_10604);
or U16964 (N_16964,N_11337,N_12171);
nor U16965 (N_16965,N_11007,N_14517);
nor U16966 (N_16966,N_10932,N_11609);
and U16967 (N_16967,N_12181,N_13941);
xor U16968 (N_16968,N_11956,N_14798);
and U16969 (N_16969,N_10553,N_10580);
or U16970 (N_16970,N_10243,N_10792);
nor U16971 (N_16971,N_10809,N_14799);
xnor U16972 (N_16972,N_14412,N_12504);
and U16973 (N_16973,N_13796,N_10186);
xor U16974 (N_16974,N_13259,N_11556);
and U16975 (N_16975,N_11727,N_12694);
nor U16976 (N_16976,N_10342,N_12229);
and U16977 (N_16977,N_10972,N_14947);
or U16978 (N_16978,N_13279,N_10222);
nor U16979 (N_16979,N_10447,N_13381);
or U16980 (N_16980,N_13014,N_10248);
and U16981 (N_16981,N_12718,N_14097);
nand U16982 (N_16982,N_11783,N_10853);
and U16983 (N_16983,N_14187,N_12465);
xnor U16984 (N_16984,N_11958,N_13907);
and U16985 (N_16985,N_14785,N_12706);
nand U16986 (N_16986,N_10955,N_10785);
nand U16987 (N_16987,N_10687,N_11746);
xor U16988 (N_16988,N_10863,N_11386);
nand U16989 (N_16989,N_11769,N_14919);
and U16990 (N_16990,N_10005,N_13477);
nand U16991 (N_16991,N_13008,N_11756);
xor U16992 (N_16992,N_10489,N_10700);
or U16993 (N_16993,N_11962,N_10001);
nand U16994 (N_16994,N_12805,N_10670);
nor U16995 (N_16995,N_12578,N_13341);
and U16996 (N_16996,N_10365,N_14538);
xnor U16997 (N_16997,N_13040,N_12306);
or U16998 (N_16998,N_10960,N_12656);
xnor U16999 (N_16999,N_11114,N_13689);
nor U17000 (N_17000,N_11551,N_10802);
nand U17001 (N_17001,N_13788,N_12036);
or U17002 (N_17002,N_13319,N_11540);
nand U17003 (N_17003,N_10244,N_13010);
xnor U17004 (N_17004,N_13147,N_13911);
xor U17005 (N_17005,N_11137,N_14451);
nand U17006 (N_17006,N_12020,N_12286);
nor U17007 (N_17007,N_12682,N_12417);
and U17008 (N_17008,N_10740,N_13600);
nor U17009 (N_17009,N_13760,N_10793);
nand U17010 (N_17010,N_12347,N_14608);
nand U17011 (N_17011,N_11313,N_11648);
and U17012 (N_17012,N_14842,N_13990);
nor U17013 (N_17013,N_10381,N_13757);
xnor U17014 (N_17014,N_10996,N_13337);
xor U17015 (N_17015,N_10904,N_14236);
xor U17016 (N_17016,N_11443,N_10595);
nand U17017 (N_17017,N_11326,N_13719);
nand U17018 (N_17018,N_10355,N_14917);
xnor U17019 (N_17019,N_10906,N_13081);
xor U17020 (N_17020,N_10530,N_10109);
and U17021 (N_17021,N_14302,N_14826);
nor U17022 (N_17022,N_10214,N_11995);
xor U17023 (N_17023,N_14700,N_11589);
nor U17024 (N_17024,N_10921,N_12099);
xor U17025 (N_17025,N_13372,N_14923);
xor U17026 (N_17026,N_14805,N_14364);
nand U17027 (N_17027,N_14779,N_11866);
nor U17028 (N_17028,N_10857,N_10947);
or U17029 (N_17029,N_12756,N_11810);
nor U17030 (N_17030,N_11577,N_14983);
and U17031 (N_17031,N_12564,N_14757);
or U17032 (N_17032,N_11565,N_12188);
nor U17033 (N_17033,N_14884,N_10414);
xor U17034 (N_17034,N_11714,N_14443);
or U17035 (N_17035,N_11444,N_12197);
xor U17036 (N_17036,N_11656,N_11699);
nor U17037 (N_17037,N_10916,N_14084);
xor U17038 (N_17038,N_10594,N_13238);
and U17039 (N_17039,N_11071,N_12627);
nand U17040 (N_17040,N_13910,N_12676);
or U17041 (N_17041,N_10213,N_14999);
or U17042 (N_17042,N_12563,N_14475);
nor U17043 (N_17043,N_13255,N_13883);
and U17044 (N_17044,N_14393,N_13068);
nor U17045 (N_17045,N_12462,N_11317);
xor U17046 (N_17046,N_14270,N_12763);
nand U17047 (N_17047,N_10601,N_10928);
or U17048 (N_17048,N_11832,N_13620);
and U17049 (N_17049,N_10129,N_12615);
nor U17050 (N_17050,N_10497,N_14224);
and U17051 (N_17051,N_10523,N_13819);
nand U17052 (N_17052,N_13791,N_10584);
and U17053 (N_17053,N_11057,N_14089);
nand U17054 (N_17054,N_11759,N_13300);
and U17055 (N_17055,N_14997,N_12714);
xor U17056 (N_17056,N_12597,N_12867);
nor U17057 (N_17057,N_12983,N_12979);
nor U17058 (N_17058,N_10079,N_10567);
xor U17059 (N_17059,N_13900,N_10025);
nor U17060 (N_17060,N_11422,N_11304);
and U17061 (N_17061,N_13392,N_13291);
nor U17062 (N_17062,N_11388,N_13149);
nor U17063 (N_17063,N_14141,N_14773);
nor U17064 (N_17064,N_14985,N_12421);
nand U17065 (N_17065,N_13254,N_10521);
xor U17066 (N_17066,N_13280,N_11364);
and U17067 (N_17067,N_11801,N_11465);
or U17068 (N_17068,N_14726,N_11250);
nand U17069 (N_17069,N_12071,N_11494);
or U17070 (N_17070,N_12242,N_11818);
nand U17071 (N_17071,N_11786,N_14751);
nand U17072 (N_17072,N_13189,N_11487);
xor U17073 (N_17073,N_11625,N_12798);
and U17074 (N_17074,N_11553,N_14436);
nand U17075 (N_17075,N_10888,N_12087);
and U17076 (N_17076,N_12093,N_13647);
nand U17077 (N_17077,N_11876,N_14900);
nor U17078 (N_17078,N_13665,N_10371);
xnor U17079 (N_17079,N_11850,N_14591);
and U17080 (N_17080,N_12684,N_11702);
nand U17081 (N_17081,N_14435,N_14013);
or U17082 (N_17082,N_12914,N_12189);
xnor U17083 (N_17083,N_14866,N_14397);
xor U17084 (N_17084,N_10841,N_13225);
and U17085 (N_17085,N_10235,N_10434);
or U17086 (N_17086,N_13552,N_13840);
or U17087 (N_17087,N_12458,N_11649);
nor U17088 (N_17088,N_11196,N_14068);
or U17089 (N_17089,N_12125,N_14851);
and U17090 (N_17090,N_10557,N_14532);
or U17091 (N_17091,N_11394,N_12041);
nand U17092 (N_17092,N_10003,N_10773);
nand U17093 (N_17093,N_12360,N_12409);
nand U17094 (N_17094,N_11880,N_11501);
and U17095 (N_17095,N_10524,N_11461);
and U17096 (N_17096,N_14510,N_10820);
xor U17097 (N_17097,N_11946,N_10915);
nand U17098 (N_17098,N_11453,N_14952);
nor U17099 (N_17099,N_13466,N_11704);
xnor U17100 (N_17100,N_12576,N_10188);
or U17101 (N_17101,N_14152,N_14423);
xor U17102 (N_17102,N_12454,N_12231);
or U17103 (N_17103,N_14095,N_11452);
and U17104 (N_17104,N_13545,N_14229);
nor U17105 (N_17105,N_12866,N_11179);
nor U17106 (N_17106,N_12527,N_13744);
nand U17107 (N_17107,N_11163,N_11279);
or U17108 (N_17108,N_11568,N_14264);
or U17109 (N_17109,N_12516,N_12770);
or U17110 (N_17110,N_12773,N_13696);
and U17111 (N_17111,N_10361,N_13469);
nand U17112 (N_17112,N_14200,N_10891);
and U17113 (N_17113,N_11004,N_12124);
nor U17114 (N_17114,N_12620,N_11316);
and U17115 (N_17115,N_12560,N_13999);
nor U17116 (N_17116,N_13741,N_11077);
nand U17117 (N_17117,N_10439,N_14231);
nand U17118 (N_17118,N_13499,N_14540);
xor U17119 (N_17119,N_13816,N_14615);
xnor U17120 (N_17120,N_12966,N_11696);
and U17121 (N_17121,N_11234,N_10585);
xnor U17122 (N_17122,N_11159,N_12263);
nand U17123 (N_17123,N_14953,N_13728);
or U17124 (N_17124,N_10923,N_14937);
xnor U17125 (N_17125,N_13919,N_11013);
and U17126 (N_17126,N_14832,N_12471);
nor U17127 (N_17127,N_13824,N_11712);
nand U17128 (N_17128,N_12599,N_10180);
nor U17129 (N_17129,N_13264,N_12172);
and U17130 (N_17130,N_10463,N_11236);
nor U17131 (N_17131,N_14911,N_11645);
xnor U17132 (N_17132,N_14117,N_10228);
and U17133 (N_17133,N_11620,N_14869);
nand U17134 (N_17134,N_14123,N_10596);
xor U17135 (N_17135,N_14519,N_12324);
and U17136 (N_17136,N_10482,N_12693);
nand U17137 (N_17137,N_12160,N_13177);
and U17138 (N_17138,N_12498,N_14907);
nor U17139 (N_17139,N_10020,N_14298);
xor U17140 (N_17140,N_11523,N_11130);
xor U17141 (N_17141,N_14738,N_11479);
nor U17142 (N_17142,N_11335,N_10858);
nor U17143 (N_17143,N_14501,N_13615);
xnor U17144 (N_17144,N_10590,N_14711);
nor U17145 (N_17145,N_10241,N_12703);
nor U17146 (N_17146,N_11168,N_14736);
nand U17147 (N_17147,N_12662,N_12163);
or U17148 (N_17148,N_12468,N_14505);
nor U17149 (N_17149,N_14651,N_10023);
or U17150 (N_17150,N_14459,N_13456);
nor U17151 (N_17151,N_10806,N_14809);
and U17152 (N_17152,N_11741,N_11298);
nor U17153 (N_17153,N_11966,N_14588);
nand U17154 (N_17154,N_14734,N_10268);
or U17155 (N_17155,N_10832,N_14886);
nor U17156 (N_17156,N_14211,N_12061);
or U17157 (N_17157,N_12530,N_11407);
or U17158 (N_17158,N_12452,N_11851);
nand U17159 (N_17159,N_11073,N_14356);
and U17160 (N_17160,N_13762,N_11899);
or U17161 (N_17161,N_12788,N_14602);
or U17162 (N_17162,N_11870,N_11413);
xor U17163 (N_17163,N_14130,N_10067);
or U17164 (N_17164,N_13562,N_13825);
or U17165 (N_17165,N_14383,N_12108);
and U17166 (N_17166,N_11076,N_14881);
nor U17167 (N_17167,N_10799,N_12735);
and U17168 (N_17168,N_12127,N_14276);
or U17169 (N_17169,N_12692,N_14642);
nor U17170 (N_17170,N_14320,N_10855);
nand U17171 (N_17171,N_14838,N_10702);
nand U17172 (N_17172,N_11026,N_14372);
or U17173 (N_17173,N_13774,N_12344);
xnor U17174 (N_17174,N_10454,N_10542);
and U17175 (N_17175,N_13351,N_14677);
nand U17176 (N_17176,N_13048,N_14590);
nand U17177 (N_17177,N_14442,N_13380);
nor U17178 (N_17178,N_11968,N_12665);
xor U17179 (N_17179,N_11935,N_11062);
xnor U17180 (N_17180,N_13221,N_11342);
nor U17181 (N_17181,N_14796,N_10811);
nand U17182 (N_17182,N_12730,N_12520);
nand U17183 (N_17183,N_13271,N_12091);
xnor U17184 (N_17184,N_11471,N_14640);
nand U17185 (N_17185,N_13304,N_13487);
and U17186 (N_17186,N_14641,N_14780);
and U17187 (N_17187,N_14283,N_13640);
nor U17188 (N_17188,N_10117,N_10780);
and U17189 (N_17189,N_13923,N_11542);
or U17190 (N_17190,N_14561,N_13138);
nand U17191 (N_17191,N_11025,N_12150);
or U17192 (N_17192,N_11457,N_13808);
nand U17193 (N_17193,N_10982,N_12382);
and U17194 (N_17194,N_11292,N_12986);
and U17195 (N_17195,N_12422,N_14732);
and U17196 (N_17196,N_11419,N_14520);
nor U17197 (N_17197,N_14162,N_11120);
xnor U17198 (N_17198,N_11843,N_11414);
xnor U17199 (N_17199,N_14649,N_13109);
xor U17200 (N_17200,N_11685,N_10310);
nor U17201 (N_17201,N_11158,N_11838);
nor U17202 (N_17202,N_14839,N_12671);
nand U17203 (N_17203,N_13787,N_10944);
nor U17204 (N_17204,N_13777,N_13375);
and U17205 (N_17205,N_14847,N_12596);
or U17206 (N_17206,N_10772,N_12490);
nor U17207 (N_17207,N_13190,N_13928);
nand U17208 (N_17208,N_13720,N_14912);
and U17209 (N_17209,N_13464,N_10549);
and U17210 (N_17210,N_11760,N_13935);
or U17211 (N_17211,N_14244,N_11311);
and U17212 (N_17212,N_11090,N_12077);
nand U17213 (N_17213,N_14696,N_10927);
and U17214 (N_17214,N_13853,N_13167);
nand U17215 (N_17215,N_11770,N_11532);
or U17216 (N_17216,N_14432,N_11262);
xnor U17217 (N_17217,N_13135,N_10821);
xnor U17218 (N_17218,N_11509,N_10990);
or U17219 (N_17219,N_12636,N_10233);
nand U17220 (N_17220,N_13473,N_14355);
nand U17221 (N_17221,N_10830,N_14043);
xor U17222 (N_17222,N_14256,N_11132);
or U17223 (N_17223,N_13474,N_13052);
and U17224 (N_17224,N_11547,N_11505);
xnor U17225 (N_17225,N_14461,N_10442);
and U17226 (N_17226,N_13516,N_14237);
nor U17227 (N_17227,N_12176,N_14856);
or U17228 (N_17228,N_14021,N_10970);
nor U17229 (N_17229,N_14747,N_10531);
xnor U17230 (N_17230,N_10774,N_10570);
nand U17231 (N_17231,N_12126,N_14007);
nand U17232 (N_17232,N_10088,N_11088);
and U17233 (N_17233,N_13688,N_14680);
nor U17234 (N_17234,N_12736,N_11993);
nor U17235 (N_17235,N_13476,N_13130);
nor U17236 (N_17236,N_12340,N_13898);
or U17237 (N_17237,N_11637,N_13178);
nand U17238 (N_17238,N_13697,N_10380);
xnor U17239 (N_17239,N_13641,N_13164);
and U17240 (N_17240,N_11717,N_14574);
and U17241 (N_17241,N_14398,N_10309);
xor U17242 (N_17242,N_11959,N_10827);
nor U17243 (N_17243,N_14980,N_10478);
xnor U17244 (N_17244,N_10417,N_10391);
nor U17245 (N_17245,N_11123,N_11932);
or U17246 (N_17246,N_11169,N_13204);
xnor U17247 (N_17247,N_14158,N_14075);
or U17248 (N_17248,N_10286,N_13371);
or U17249 (N_17249,N_14628,N_14683);
and U17250 (N_17250,N_11293,N_13959);
or U17251 (N_17251,N_13773,N_12696);
nor U17252 (N_17252,N_11848,N_10761);
nand U17253 (N_17253,N_13123,N_13903);
xnor U17254 (N_17254,N_14251,N_14735);
nand U17255 (N_17255,N_11634,N_11131);
and U17256 (N_17256,N_10334,N_11092);
nand U17257 (N_17257,N_11983,N_11020);
nor U17258 (N_17258,N_14821,N_12953);
nand U17259 (N_17259,N_12997,N_13732);
nor U17260 (N_17260,N_13917,N_13449);
and U17261 (N_17261,N_13852,N_13645);
or U17262 (N_17262,N_13031,N_12577);
xor U17263 (N_17263,N_11954,N_14610);
nand U17264 (N_17264,N_13329,N_10528);
nor U17265 (N_17265,N_13837,N_14259);
nor U17266 (N_17266,N_11209,N_10692);
xnor U17267 (N_17267,N_13191,N_13548);
nor U17268 (N_17268,N_12357,N_14119);
or U17269 (N_17269,N_12082,N_14463);
or U17270 (N_17270,N_11226,N_13216);
nand U17271 (N_17271,N_14149,N_12312);
nor U17272 (N_17272,N_12291,N_12348);
or U17273 (N_17273,N_13770,N_14230);
nand U17274 (N_17274,N_10258,N_11333);
nor U17275 (N_17275,N_13746,N_13833);
xnor U17276 (N_17276,N_11877,N_14469);
xor U17277 (N_17277,N_10675,N_12619);
nand U17278 (N_17278,N_10925,N_12766);
xnor U17279 (N_17279,N_14536,N_13388);
and U17280 (N_17280,N_12876,N_12115);
nand U17281 (N_17281,N_11084,N_12932);
nand U17282 (N_17282,N_13901,N_10910);
nand U17283 (N_17283,N_11239,N_13288);
xor U17284 (N_17284,N_14055,N_10607);
xnor U17285 (N_17285,N_13284,N_11432);
and U17286 (N_17286,N_13987,N_13398);
nand U17287 (N_17287,N_14284,N_12549);
nand U17288 (N_17288,N_12931,N_12198);
xor U17289 (N_17289,N_13461,N_10339);
xor U17290 (N_17290,N_10645,N_12063);
nor U17291 (N_17291,N_10555,N_11002);
and U17292 (N_17292,N_13490,N_12759);
nand U17293 (N_17293,N_13290,N_12487);
nand U17294 (N_17294,N_13882,N_13366);
and U17295 (N_17295,N_13019,N_14419);
or U17296 (N_17296,N_12258,N_12688);
xor U17297 (N_17297,N_11613,N_12617);
and U17298 (N_17298,N_13382,N_10294);
and U17299 (N_17299,N_13314,N_13057);
xor U17300 (N_17300,N_10424,N_11650);
xor U17301 (N_17301,N_13839,N_13715);
xor U17302 (N_17302,N_12660,N_14666);
nand U17303 (N_17303,N_14506,N_12406);
or U17304 (N_17304,N_10954,N_13324);
xnor U17305 (N_17305,N_13399,N_12354);
nor U17306 (N_17306,N_10563,N_13299);
or U17307 (N_17307,N_14727,N_12443);
nand U17308 (N_17308,N_12512,N_14185);
or U17309 (N_17309,N_13158,N_14199);
xor U17310 (N_17310,N_13594,N_14202);
nand U17311 (N_17311,N_12776,N_13106);
or U17312 (N_17312,N_11240,N_14345);
xor U17313 (N_17313,N_11268,N_14604);
xor U17314 (N_17314,N_14164,N_10444);
or U17315 (N_17315,N_13571,N_13680);
nand U17316 (N_17316,N_13007,N_13747);
or U17317 (N_17317,N_13070,N_14550);
and U17318 (N_17318,N_14481,N_12144);
nand U17319 (N_17319,N_14362,N_12937);
xnor U17320 (N_17320,N_10022,N_13817);
nor U17321 (N_17321,N_12416,N_12280);
nand U17322 (N_17322,N_10742,N_14664);
or U17323 (N_17323,N_11361,N_12910);
xnor U17324 (N_17324,N_14528,N_14331);
and U17325 (N_17325,N_12852,N_14279);
and U17326 (N_17326,N_12945,N_11731);
nand U17327 (N_17327,N_13397,N_13546);
nor U17328 (N_17328,N_11969,N_11561);
or U17329 (N_17329,N_10544,N_10790);
nor U17330 (N_17330,N_11106,N_14920);
nand U17331 (N_17331,N_14575,N_10576);
xnor U17332 (N_17332,N_10083,N_13682);
xor U17333 (N_17333,N_14918,N_13467);
nor U17334 (N_17334,N_10872,N_12210);
and U17335 (N_17335,N_10909,N_10900);
and U17336 (N_17336,N_11767,N_10226);
nor U17337 (N_17337,N_14440,N_13453);
xnor U17338 (N_17338,N_11924,N_13465);
xor U17339 (N_17339,N_13209,N_12621);
xnor U17340 (N_17340,N_11391,N_12609);
nand U17341 (N_17341,N_12872,N_12436);
xnor U17342 (N_17342,N_10573,N_10193);
and U17343 (N_17343,N_10031,N_11241);
or U17344 (N_17344,N_12461,N_12514);
or U17345 (N_17345,N_14755,N_11327);
xor U17346 (N_17346,N_14639,N_11334);
nor U17347 (N_17347,N_10418,N_10151);
nand U17348 (N_17348,N_10610,N_10084);
or U17349 (N_17349,N_12786,N_14093);
nand U17350 (N_17350,N_11199,N_11112);
xnor U17351 (N_17351,N_13338,N_13431);
nand U17352 (N_17352,N_10520,N_13706);
xnor U17353 (N_17353,N_13738,N_12946);
and U17354 (N_17354,N_13320,N_11820);
nor U17355 (N_17355,N_13215,N_10285);
xor U17356 (N_17356,N_11816,N_14415);
nand U17357 (N_17357,N_11098,N_10451);
and U17358 (N_17358,N_12133,N_10353);
nor U17359 (N_17359,N_12094,N_12865);
nand U17360 (N_17360,N_13567,N_13966);
and U17361 (N_17361,N_10814,N_10695);
xnor U17362 (N_17362,N_12793,N_10051);
and U17363 (N_17363,N_11027,N_12792);
xor U17364 (N_17364,N_14295,N_14133);
xnor U17365 (N_17365,N_11165,N_12441);
or U17366 (N_17366,N_10995,N_14108);
and U17367 (N_17367,N_12469,N_13733);
xnor U17368 (N_17368,N_13239,N_13395);
or U17369 (N_17369,N_14401,N_13727);
nor U17370 (N_17370,N_11915,N_11133);
nor U17371 (N_17371,N_12663,N_10460);
or U17372 (N_17372,N_13669,N_11477);
nor U17373 (N_17373,N_13751,N_10160);
xor U17374 (N_17374,N_13443,N_10179);
or U17375 (N_17375,N_13451,N_13440);
xor U17376 (N_17376,N_12892,N_10453);
xnor U17377 (N_17377,N_13662,N_10560);
nand U17378 (N_17378,N_13767,N_13145);
and U17379 (N_17379,N_10448,N_12369);
or U17380 (N_17380,N_13364,N_10666);
or U17381 (N_17381,N_14205,N_13892);
nand U17382 (N_17382,N_12896,N_14025);
and U17383 (N_17383,N_10981,N_13844);
nor U17384 (N_17384,N_11608,N_10436);
and U17385 (N_17385,N_14492,N_14893);
or U17386 (N_17386,N_14672,N_13087);
or U17387 (N_17387,N_10617,N_12894);
nor U17388 (N_17388,N_14635,N_12919);
nor U17389 (N_17389,N_11383,N_10903);
xor U17390 (N_17390,N_13129,N_10393);
nor U17391 (N_17391,N_11185,N_13610);
or U17392 (N_17392,N_10095,N_12453);
or U17393 (N_17393,N_11869,N_11427);
nand U17394 (N_17394,N_12584,N_12875);
nand U17395 (N_17395,N_10251,N_11082);
and U17396 (N_17396,N_11023,N_14430);
nor U17397 (N_17397,N_11124,N_12658);
and U17398 (N_17398,N_13815,N_10274);
and U17399 (N_17399,N_13996,N_11016);
nand U17400 (N_17400,N_11064,N_13710);
or U17401 (N_17401,N_11537,N_11527);
xnor U17402 (N_17402,N_11522,N_12463);
nand U17403 (N_17403,N_10599,N_11031);
nand U17404 (N_17404,N_12757,N_11793);
nor U17405 (N_17405,N_10141,N_10481);
xor U17406 (N_17406,N_14088,N_10989);
xnor U17407 (N_17407,N_12032,N_12622);
and U17408 (N_17408,N_12426,N_14445);
nor U17409 (N_17409,N_14159,N_10876);
nand U17410 (N_17410,N_10892,N_11514);
nand U17411 (N_17411,N_12844,N_14474);
nand U17412 (N_17412,N_13886,N_10794);
and U17413 (N_17413,N_10019,N_12542);
and U17414 (N_17414,N_13859,N_10428);
and U17415 (N_17415,N_11219,N_11730);
xnor U17416 (N_17416,N_11630,N_12613);
and U17417 (N_17417,N_10043,N_12167);
or U17418 (N_17418,N_13722,N_10102);
or U17419 (N_17419,N_12358,N_12990);
nor U17420 (N_17420,N_14718,N_12287);
xnor U17421 (N_17421,N_10254,N_14737);
xor U17422 (N_17422,N_11463,N_10637);
nor U17423 (N_17423,N_10072,N_12029);
nand U17424 (N_17424,N_14789,N_11299);
nand U17425 (N_17425,N_11679,N_13505);
xnor U17426 (N_17426,N_12540,N_13406);
xor U17427 (N_17427,N_13195,N_12395);
nand U17428 (N_17428,N_13716,N_11010);
and U17429 (N_17429,N_13768,N_14705);
xnor U17430 (N_17430,N_11652,N_14248);
or U17431 (N_17431,N_11200,N_14928);
xor U17432 (N_17432,N_11308,N_14555);
or U17433 (N_17433,N_13425,N_12370);
and U17434 (N_17434,N_11245,N_13494);
and U17435 (N_17435,N_10893,N_11931);
xor U17436 (N_17436,N_11433,N_12769);
and U17437 (N_17437,N_11771,N_14848);
or U17438 (N_17438,N_10118,N_10685);
xor U17439 (N_17439,N_12479,N_13103);
xor U17440 (N_17440,N_10433,N_11990);
nor U17441 (N_17441,N_12594,N_10969);
and U17442 (N_17442,N_12222,N_14558);
nand U17443 (N_17443,N_12366,N_12397);
nand U17444 (N_17444,N_14731,N_14139);
nor U17445 (N_17445,N_14939,N_10536);
nand U17446 (N_17446,N_13484,N_13169);
nor U17447 (N_17447,N_14990,N_14171);
nor U17448 (N_17448,N_14273,N_13947);
and U17449 (N_17449,N_10973,N_12451);
nor U17450 (N_17450,N_13401,N_13508);
xnor U17451 (N_17451,N_12840,N_12851);
or U17452 (N_17452,N_11636,N_13997);
or U17453 (N_17453,N_12978,N_14210);
and U17454 (N_17454,N_12269,N_12309);
or U17455 (N_17455,N_12862,N_10437);
or U17456 (N_17456,N_12804,N_13659);
and U17457 (N_17457,N_13317,N_12561);
xor U17458 (N_17458,N_10963,N_10616);
or U17459 (N_17459,N_14197,N_13298);
xnor U17460 (N_17460,N_11520,N_11052);
xnor U17461 (N_17461,N_14176,N_13350);
and U17462 (N_17462,N_10507,N_12447);
and U17463 (N_17463,N_14668,N_10719);
or U17464 (N_17464,N_11045,N_14358);
nand U17465 (N_17465,N_10744,N_13237);
nor U17466 (N_17466,N_14586,N_10770);
and U17467 (N_17467,N_10786,N_11048);
nand U17468 (N_17468,N_14667,N_12976);
and U17469 (N_17469,N_14882,N_13772);
or U17470 (N_17470,N_12848,N_12541);
nor U17471 (N_17471,N_11908,N_11210);
xor U17472 (N_17472,N_12444,N_14409);
or U17473 (N_17473,N_12630,N_13378);
xor U17474 (N_17474,N_14011,N_13234);
nor U17475 (N_17475,N_13394,N_12538);
and U17476 (N_17476,N_13393,N_13673);
nand U17477 (N_17477,N_12523,N_14464);
nor U17478 (N_17478,N_13102,N_14029);
xor U17479 (N_17479,N_11907,N_11249);
xor U17480 (N_17480,N_13983,N_12641);
and U17481 (N_17481,N_14452,N_12112);
nand U17482 (N_17482,N_10722,N_11229);
or U17483 (N_17483,N_10085,N_14102);
nor U17484 (N_17484,N_10456,N_11950);
or U17485 (N_17485,N_10789,N_14781);
nand U17486 (N_17486,N_13475,N_13557);
xnor U17487 (N_17487,N_11153,N_10475);
nand U17488 (N_17488,N_13511,N_12826);
nor U17489 (N_17489,N_11726,N_14175);
nor U17490 (N_17490,N_12681,N_13827);
nand U17491 (N_17491,N_10935,N_13795);
nand U17492 (N_17492,N_12638,N_14633);
xor U17493 (N_17493,N_10124,N_11478);
or U17494 (N_17494,N_14637,N_12355);
or U17495 (N_17495,N_11458,N_13628);
nand U17496 (N_17496,N_11564,N_10038);
or U17497 (N_17497,N_12278,N_13053);
and U17498 (N_17498,N_12213,N_11815);
and U17499 (N_17499,N_14915,N_14948);
or U17500 (N_17500,N_11958,N_12572);
xnor U17501 (N_17501,N_10976,N_11929);
nand U17502 (N_17502,N_13339,N_10773);
or U17503 (N_17503,N_11566,N_11894);
xnor U17504 (N_17504,N_13884,N_11766);
and U17505 (N_17505,N_12277,N_12035);
xnor U17506 (N_17506,N_11193,N_12724);
xor U17507 (N_17507,N_14726,N_13253);
nand U17508 (N_17508,N_11657,N_12754);
xor U17509 (N_17509,N_14762,N_11572);
and U17510 (N_17510,N_13396,N_14227);
or U17511 (N_17511,N_11284,N_14045);
nor U17512 (N_17512,N_14069,N_13910);
or U17513 (N_17513,N_10997,N_12832);
nand U17514 (N_17514,N_11521,N_12323);
and U17515 (N_17515,N_11395,N_12895);
xor U17516 (N_17516,N_12773,N_12843);
xnor U17517 (N_17517,N_13813,N_11614);
nand U17518 (N_17518,N_10989,N_13405);
nand U17519 (N_17519,N_14120,N_12770);
xor U17520 (N_17520,N_11157,N_10107);
nand U17521 (N_17521,N_12503,N_12054);
and U17522 (N_17522,N_13598,N_14954);
nor U17523 (N_17523,N_14956,N_10727);
and U17524 (N_17524,N_14062,N_13159);
nand U17525 (N_17525,N_10406,N_10675);
xor U17526 (N_17526,N_10625,N_14590);
or U17527 (N_17527,N_11704,N_10158);
nor U17528 (N_17528,N_10348,N_10856);
nor U17529 (N_17529,N_10699,N_12507);
nor U17530 (N_17530,N_13692,N_12384);
or U17531 (N_17531,N_13785,N_10623);
nand U17532 (N_17532,N_14863,N_13554);
xor U17533 (N_17533,N_13710,N_13944);
nor U17534 (N_17534,N_11023,N_11848);
nand U17535 (N_17535,N_13939,N_10138);
or U17536 (N_17536,N_13609,N_10182);
and U17537 (N_17537,N_10623,N_11287);
nor U17538 (N_17538,N_10935,N_10174);
nand U17539 (N_17539,N_13934,N_14121);
nand U17540 (N_17540,N_14805,N_12538);
or U17541 (N_17541,N_13838,N_11339);
or U17542 (N_17542,N_10032,N_13117);
and U17543 (N_17543,N_14237,N_10725);
or U17544 (N_17544,N_13108,N_11478);
xnor U17545 (N_17545,N_11590,N_10773);
and U17546 (N_17546,N_10592,N_14275);
nor U17547 (N_17547,N_14823,N_10053);
nor U17548 (N_17548,N_13025,N_12318);
and U17549 (N_17549,N_14196,N_14153);
or U17550 (N_17550,N_11999,N_12389);
or U17551 (N_17551,N_12060,N_11718);
nor U17552 (N_17552,N_10302,N_12742);
xnor U17553 (N_17553,N_10465,N_12465);
nor U17554 (N_17554,N_10536,N_11960);
xor U17555 (N_17555,N_10114,N_14994);
and U17556 (N_17556,N_14078,N_11029);
or U17557 (N_17557,N_14089,N_10921);
and U17558 (N_17558,N_13069,N_13115);
xor U17559 (N_17559,N_12120,N_13840);
or U17560 (N_17560,N_12339,N_14294);
xnor U17561 (N_17561,N_13696,N_14550);
and U17562 (N_17562,N_10699,N_14844);
nor U17563 (N_17563,N_11448,N_12494);
nor U17564 (N_17564,N_13619,N_13642);
nor U17565 (N_17565,N_13500,N_10192);
nand U17566 (N_17566,N_13315,N_10255);
nand U17567 (N_17567,N_11139,N_12413);
nand U17568 (N_17568,N_11855,N_12476);
xnor U17569 (N_17569,N_12574,N_10519);
and U17570 (N_17570,N_12843,N_14117);
nor U17571 (N_17571,N_14131,N_10515);
and U17572 (N_17572,N_10047,N_11579);
and U17573 (N_17573,N_14271,N_11527);
xor U17574 (N_17574,N_13562,N_13377);
and U17575 (N_17575,N_10489,N_11242);
or U17576 (N_17576,N_12764,N_10800);
and U17577 (N_17577,N_13667,N_13480);
xnor U17578 (N_17578,N_11505,N_13998);
or U17579 (N_17579,N_11302,N_13942);
or U17580 (N_17580,N_11745,N_11050);
and U17581 (N_17581,N_11273,N_12515);
nand U17582 (N_17582,N_11397,N_12793);
or U17583 (N_17583,N_12019,N_13445);
nand U17584 (N_17584,N_10329,N_10099);
xor U17585 (N_17585,N_10274,N_13742);
or U17586 (N_17586,N_12683,N_11186);
xnor U17587 (N_17587,N_10553,N_14778);
xnor U17588 (N_17588,N_13842,N_12107);
or U17589 (N_17589,N_10173,N_11657);
and U17590 (N_17590,N_14370,N_13091);
nand U17591 (N_17591,N_12821,N_10998);
nand U17592 (N_17592,N_12388,N_13282);
nor U17593 (N_17593,N_14622,N_13403);
xor U17594 (N_17594,N_11853,N_13417);
nand U17595 (N_17595,N_14928,N_11636);
and U17596 (N_17596,N_13588,N_11591);
xnor U17597 (N_17597,N_14857,N_12602);
and U17598 (N_17598,N_12007,N_13506);
and U17599 (N_17599,N_14867,N_11049);
xor U17600 (N_17600,N_12551,N_10915);
nand U17601 (N_17601,N_13668,N_14359);
or U17602 (N_17602,N_14473,N_11403);
and U17603 (N_17603,N_13258,N_14770);
and U17604 (N_17604,N_10505,N_14899);
nand U17605 (N_17605,N_11039,N_14037);
and U17606 (N_17606,N_12508,N_14246);
xnor U17607 (N_17607,N_12258,N_14884);
nand U17608 (N_17608,N_11970,N_14499);
nand U17609 (N_17609,N_10126,N_14732);
nand U17610 (N_17610,N_14198,N_10761);
xor U17611 (N_17611,N_10517,N_10846);
or U17612 (N_17612,N_11153,N_12463);
nor U17613 (N_17613,N_10060,N_12880);
or U17614 (N_17614,N_12185,N_14904);
nor U17615 (N_17615,N_13917,N_14264);
or U17616 (N_17616,N_10500,N_14083);
or U17617 (N_17617,N_10456,N_11466);
xnor U17618 (N_17618,N_14557,N_11571);
or U17619 (N_17619,N_11113,N_11297);
and U17620 (N_17620,N_14992,N_13057);
nand U17621 (N_17621,N_13389,N_14002);
xor U17622 (N_17622,N_13047,N_12201);
and U17623 (N_17623,N_14103,N_14264);
and U17624 (N_17624,N_14168,N_12903);
nand U17625 (N_17625,N_10094,N_13776);
nand U17626 (N_17626,N_10938,N_12642);
or U17627 (N_17627,N_14467,N_14513);
or U17628 (N_17628,N_14963,N_12098);
nor U17629 (N_17629,N_13746,N_11529);
xor U17630 (N_17630,N_10844,N_13326);
or U17631 (N_17631,N_10741,N_14538);
xor U17632 (N_17632,N_11990,N_11446);
and U17633 (N_17633,N_14801,N_14515);
xor U17634 (N_17634,N_10907,N_10803);
or U17635 (N_17635,N_13803,N_14209);
and U17636 (N_17636,N_13932,N_13491);
nand U17637 (N_17637,N_14777,N_11775);
nand U17638 (N_17638,N_11723,N_13079);
nand U17639 (N_17639,N_13314,N_13906);
nand U17640 (N_17640,N_11754,N_14861);
nand U17641 (N_17641,N_10158,N_14548);
or U17642 (N_17642,N_11965,N_13939);
and U17643 (N_17643,N_14452,N_10417);
and U17644 (N_17644,N_14725,N_12453);
nor U17645 (N_17645,N_13071,N_12744);
nand U17646 (N_17646,N_11824,N_13188);
xor U17647 (N_17647,N_12275,N_11936);
xnor U17648 (N_17648,N_14002,N_13884);
nor U17649 (N_17649,N_14158,N_13765);
or U17650 (N_17650,N_11834,N_14758);
or U17651 (N_17651,N_13368,N_12309);
or U17652 (N_17652,N_13487,N_13787);
or U17653 (N_17653,N_12733,N_13856);
xor U17654 (N_17654,N_13788,N_14091);
nor U17655 (N_17655,N_14028,N_10241);
nand U17656 (N_17656,N_14108,N_14274);
or U17657 (N_17657,N_10673,N_14859);
or U17658 (N_17658,N_14777,N_11804);
nor U17659 (N_17659,N_14879,N_11871);
xnor U17660 (N_17660,N_11288,N_11596);
and U17661 (N_17661,N_12711,N_12565);
nor U17662 (N_17662,N_12336,N_11718);
and U17663 (N_17663,N_10933,N_10789);
nor U17664 (N_17664,N_11827,N_14498);
nand U17665 (N_17665,N_13687,N_11540);
and U17666 (N_17666,N_11229,N_11158);
or U17667 (N_17667,N_10339,N_11563);
nand U17668 (N_17668,N_14497,N_13733);
xor U17669 (N_17669,N_11385,N_11313);
nor U17670 (N_17670,N_14200,N_14569);
and U17671 (N_17671,N_10603,N_10254);
or U17672 (N_17672,N_14353,N_13596);
nor U17673 (N_17673,N_14888,N_11478);
and U17674 (N_17674,N_13005,N_10411);
nand U17675 (N_17675,N_10765,N_13477);
and U17676 (N_17676,N_11391,N_13655);
or U17677 (N_17677,N_13256,N_10252);
nor U17678 (N_17678,N_12091,N_12973);
and U17679 (N_17679,N_11132,N_14222);
nor U17680 (N_17680,N_10973,N_10727);
and U17681 (N_17681,N_12397,N_13274);
and U17682 (N_17682,N_11184,N_12758);
xnor U17683 (N_17683,N_11751,N_11422);
nor U17684 (N_17684,N_10045,N_10840);
and U17685 (N_17685,N_13569,N_12145);
xnor U17686 (N_17686,N_10924,N_14232);
nand U17687 (N_17687,N_12014,N_13749);
and U17688 (N_17688,N_12301,N_12685);
and U17689 (N_17689,N_14745,N_13980);
nor U17690 (N_17690,N_13130,N_13587);
or U17691 (N_17691,N_11649,N_10926);
xor U17692 (N_17692,N_10135,N_11494);
and U17693 (N_17693,N_13310,N_12745);
and U17694 (N_17694,N_13642,N_12845);
xor U17695 (N_17695,N_11362,N_13866);
nor U17696 (N_17696,N_13005,N_11793);
nor U17697 (N_17697,N_11369,N_12056);
and U17698 (N_17698,N_14920,N_11222);
nor U17699 (N_17699,N_14317,N_10429);
xnor U17700 (N_17700,N_10101,N_12406);
nand U17701 (N_17701,N_14110,N_11512);
nor U17702 (N_17702,N_14396,N_14903);
or U17703 (N_17703,N_12350,N_11276);
nor U17704 (N_17704,N_13332,N_12201);
or U17705 (N_17705,N_12848,N_13144);
or U17706 (N_17706,N_10026,N_12319);
nor U17707 (N_17707,N_13612,N_13334);
nor U17708 (N_17708,N_10267,N_11879);
nor U17709 (N_17709,N_14010,N_10409);
and U17710 (N_17710,N_12262,N_14596);
nor U17711 (N_17711,N_12943,N_10444);
and U17712 (N_17712,N_10864,N_12723);
and U17713 (N_17713,N_12153,N_11602);
xnor U17714 (N_17714,N_11770,N_12935);
nand U17715 (N_17715,N_11927,N_14839);
or U17716 (N_17716,N_12953,N_11092);
xor U17717 (N_17717,N_10092,N_10720);
xnor U17718 (N_17718,N_12114,N_10516);
xor U17719 (N_17719,N_12605,N_11458);
xor U17720 (N_17720,N_10001,N_14976);
or U17721 (N_17721,N_13414,N_13170);
nor U17722 (N_17722,N_10553,N_14653);
xnor U17723 (N_17723,N_10134,N_10913);
nor U17724 (N_17724,N_12934,N_12020);
xnor U17725 (N_17725,N_11316,N_12906);
or U17726 (N_17726,N_13178,N_13756);
nor U17727 (N_17727,N_10318,N_10389);
nand U17728 (N_17728,N_10776,N_11736);
nand U17729 (N_17729,N_11298,N_13866);
and U17730 (N_17730,N_14871,N_13682);
xor U17731 (N_17731,N_10588,N_11313);
or U17732 (N_17732,N_13971,N_11711);
and U17733 (N_17733,N_11371,N_11584);
nor U17734 (N_17734,N_12597,N_12467);
nor U17735 (N_17735,N_10765,N_12553);
or U17736 (N_17736,N_12887,N_12330);
xor U17737 (N_17737,N_14509,N_11690);
xor U17738 (N_17738,N_14872,N_11952);
xor U17739 (N_17739,N_14731,N_12586);
xnor U17740 (N_17740,N_12823,N_10255);
nand U17741 (N_17741,N_11629,N_11468);
xnor U17742 (N_17742,N_14358,N_10256);
nand U17743 (N_17743,N_11842,N_14307);
nor U17744 (N_17744,N_13176,N_11254);
xnor U17745 (N_17745,N_10514,N_11001);
xnor U17746 (N_17746,N_11401,N_12493);
nand U17747 (N_17747,N_14258,N_10227);
nand U17748 (N_17748,N_12141,N_11271);
or U17749 (N_17749,N_14815,N_12403);
or U17750 (N_17750,N_13951,N_13323);
and U17751 (N_17751,N_14772,N_10944);
xnor U17752 (N_17752,N_10798,N_13615);
nor U17753 (N_17753,N_12865,N_14491);
xor U17754 (N_17754,N_11168,N_11991);
and U17755 (N_17755,N_13927,N_10362);
nor U17756 (N_17756,N_13220,N_10052);
or U17757 (N_17757,N_11648,N_11347);
and U17758 (N_17758,N_10209,N_10726);
nor U17759 (N_17759,N_14556,N_10244);
nor U17760 (N_17760,N_11406,N_13762);
nor U17761 (N_17761,N_12718,N_13769);
xor U17762 (N_17762,N_14726,N_14672);
nand U17763 (N_17763,N_10351,N_13685);
or U17764 (N_17764,N_13147,N_13404);
and U17765 (N_17765,N_13745,N_13866);
nor U17766 (N_17766,N_13912,N_11288);
xor U17767 (N_17767,N_11628,N_10704);
xor U17768 (N_17768,N_11965,N_12446);
and U17769 (N_17769,N_10995,N_14199);
nand U17770 (N_17770,N_10975,N_11689);
and U17771 (N_17771,N_13668,N_10145);
nor U17772 (N_17772,N_14023,N_11782);
nand U17773 (N_17773,N_11259,N_14981);
xor U17774 (N_17774,N_12908,N_13189);
and U17775 (N_17775,N_12176,N_12981);
nor U17776 (N_17776,N_10538,N_13916);
nand U17777 (N_17777,N_11692,N_12737);
nand U17778 (N_17778,N_14579,N_13390);
and U17779 (N_17779,N_10850,N_10053);
or U17780 (N_17780,N_14656,N_10365);
nor U17781 (N_17781,N_12744,N_14659);
nand U17782 (N_17782,N_11537,N_13276);
and U17783 (N_17783,N_14611,N_11299);
and U17784 (N_17784,N_11419,N_14617);
nor U17785 (N_17785,N_11440,N_14492);
nand U17786 (N_17786,N_14983,N_11944);
or U17787 (N_17787,N_12150,N_11549);
nand U17788 (N_17788,N_11585,N_12127);
nor U17789 (N_17789,N_11355,N_10880);
nor U17790 (N_17790,N_12544,N_10030);
nand U17791 (N_17791,N_13975,N_10443);
or U17792 (N_17792,N_14253,N_10680);
or U17793 (N_17793,N_14879,N_14216);
or U17794 (N_17794,N_13174,N_12431);
xor U17795 (N_17795,N_12805,N_13820);
and U17796 (N_17796,N_13251,N_10804);
xor U17797 (N_17797,N_13755,N_13482);
xor U17798 (N_17798,N_13948,N_12394);
nor U17799 (N_17799,N_12617,N_12268);
xnor U17800 (N_17800,N_14922,N_12711);
and U17801 (N_17801,N_11127,N_10133);
nand U17802 (N_17802,N_12545,N_14165);
nand U17803 (N_17803,N_11623,N_14564);
xnor U17804 (N_17804,N_14417,N_12976);
or U17805 (N_17805,N_10584,N_14090);
xnor U17806 (N_17806,N_10808,N_11990);
xnor U17807 (N_17807,N_14538,N_14760);
nor U17808 (N_17808,N_12100,N_13399);
and U17809 (N_17809,N_10547,N_11697);
and U17810 (N_17810,N_14364,N_12175);
xnor U17811 (N_17811,N_12036,N_11399);
xnor U17812 (N_17812,N_13666,N_10294);
nor U17813 (N_17813,N_13797,N_14329);
xor U17814 (N_17814,N_13668,N_10013);
nand U17815 (N_17815,N_11119,N_11344);
nor U17816 (N_17816,N_13907,N_12562);
xnor U17817 (N_17817,N_10098,N_11071);
nor U17818 (N_17818,N_14896,N_13501);
and U17819 (N_17819,N_12322,N_11489);
and U17820 (N_17820,N_14718,N_12054);
nand U17821 (N_17821,N_11404,N_13975);
xnor U17822 (N_17822,N_11654,N_11279);
nor U17823 (N_17823,N_13498,N_13362);
nor U17824 (N_17824,N_12649,N_10236);
and U17825 (N_17825,N_12750,N_13957);
xnor U17826 (N_17826,N_14198,N_13950);
nand U17827 (N_17827,N_10383,N_11992);
nand U17828 (N_17828,N_13730,N_12609);
xor U17829 (N_17829,N_14747,N_12433);
nor U17830 (N_17830,N_12546,N_14556);
nor U17831 (N_17831,N_12624,N_11365);
or U17832 (N_17832,N_14374,N_12801);
and U17833 (N_17833,N_12149,N_14008);
nor U17834 (N_17834,N_13385,N_14914);
nor U17835 (N_17835,N_13574,N_14766);
or U17836 (N_17836,N_12884,N_13542);
nand U17837 (N_17837,N_10585,N_10726);
and U17838 (N_17838,N_14649,N_14276);
xor U17839 (N_17839,N_11753,N_11274);
nand U17840 (N_17840,N_10057,N_10578);
or U17841 (N_17841,N_12004,N_14658);
or U17842 (N_17842,N_10517,N_10409);
xor U17843 (N_17843,N_14410,N_14102);
xor U17844 (N_17844,N_10817,N_13650);
and U17845 (N_17845,N_14291,N_13180);
xor U17846 (N_17846,N_12376,N_10242);
nand U17847 (N_17847,N_13374,N_14220);
nor U17848 (N_17848,N_10435,N_11151);
nand U17849 (N_17849,N_13963,N_13351);
nor U17850 (N_17850,N_10387,N_11707);
xnor U17851 (N_17851,N_10956,N_11677);
nand U17852 (N_17852,N_13677,N_14739);
and U17853 (N_17853,N_12605,N_11749);
xnor U17854 (N_17854,N_11021,N_13703);
nor U17855 (N_17855,N_14890,N_12250);
nand U17856 (N_17856,N_14932,N_10843);
xnor U17857 (N_17857,N_14679,N_14580);
or U17858 (N_17858,N_10385,N_11949);
or U17859 (N_17859,N_13956,N_10629);
nor U17860 (N_17860,N_10514,N_10876);
or U17861 (N_17861,N_10161,N_13879);
or U17862 (N_17862,N_12164,N_11797);
xnor U17863 (N_17863,N_14229,N_12930);
nor U17864 (N_17864,N_13308,N_14823);
nor U17865 (N_17865,N_11687,N_13941);
and U17866 (N_17866,N_13350,N_13461);
nand U17867 (N_17867,N_11712,N_13449);
nand U17868 (N_17868,N_12536,N_14798);
nand U17869 (N_17869,N_12365,N_11567);
nor U17870 (N_17870,N_10387,N_10035);
or U17871 (N_17871,N_10696,N_14378);
or U17872 (N_17872,N_12689,N_12337);
or U17873 (N_17873,N_10938,N_11410);
or U17874 (N_17874,N_14816,N_13768);
or U17875 (N_17875,N_12765,N_13974);
nand U17876 (N_17876,N_14166,N_13107);
nor U17877 (N_17877,N_11510,N_11153);
xnor U17878 (N_17878,N_12558,N_11675);
and U17879 (N_17879,N_13524,N_11048);
xor U17880 (N_17880,N_14653,N_14465);
or U17881 (N_17881,N_10525,N_12825);
xnor U17882 (N_17882,N_13698,N_12860);
or U17883 (N_17883,N_10418,N_10736);
xnor U17884 (N_17884,N_14986,N_12874);
nor U17885 (N_17885,N_12062,N_11473);
or U17886 (N_17886,N_10199,N_11625);
xor U17887 (N_17887,N_10536,N_14121);
or U17888 (N_17888,N_12574,N_10603);
nand U17889 (N_17889,N_13385,N_10210);
or U17890 (N_17890,N_11855,N_10177);
nor U17891 (N_17891,N_12444,N_14901);
nor U17892 (N_17892,N_13059,N_12881);
nor U17893 (N_17893,N_12633,N_13379);
nand U17894 (N_17894,N_13241,N_14827);
or U17895 (N_17895,N_13738,N_12172);
xor U17896 (N_17896,N_13533,N_11851);
nand U17897 (N_17897,N_12203,N_10649);
nor U17898 (N_17898,N_13561,N_14518);
nand U17899 (N_17899,N_13025,N_14627);
nand U17900 (N_17900,N_13474,N_12000);
or U17901 (N_17901,N_10785,N_11222);
or U17902 (N_17902,N_11167,N_14237);
and U17903 (N_17903,N_13728,N_11094);
xor U17904 (N_17904,N_13917,N_12937);
or U17905 (N_17905,N_10827,N_14835);
or U17906 (N_17906,N_12190,N_12525);
and U17907 (N_17907,N_10137,N_14816);
and U17908 (N_17908,N_13862,N_13807);
and U17909 (N_17909,N_11972,N_11313);
nand U17910 (N_17910,N_11506,N_10749);
or U17911 (N_17911,N_13590,N_11797);
and U17912 (N_17912,N_10638,N_13576);
or U17913 (N_17913,N_14856,N_13853);
xnor U17914 (N_17914,N_12757,N_13428);
or U17915 (N_17915,N_10838,N_13623);
nor U17916 (N_17916,N_12034,N_12866);
and U17917 (N_17917,N_11688,N_10900);
and U17918 (N_17918,N_14644,N_13427);
or U17919 (N_17919,N_14346,N_10165);
xor U17920 (N_17920,N_13166,N_14591);
nand U17921 (N_17921,N_13439,N_11251);
nor U17922 (N_17922,N_10848,N_14663);
or U17923 (N_17923,N_13178,N_12206);
nor U17924 (N_17924,N_12070,N_10633);
nand U17925 (N_17925,N_12554,N_12661);
and U17926 (N_17926,N_12961,N_14807);
nand U17927 (N_17927,N_12085,N_10023);
nand U17928 (N_17928,N_11463,N_13166);
or U17929 (N_17929,N_13043,N_12389);
nand U17930 (N_17930,N_11538,N_13658);
and U17931 (N_17931,N_14621,N_11069);
xnor U17932 (N_17932,N_10383,N_11558);
and U17933 (N_17933,N_11733,N_12698);
nand U17934 (N_17934,N_10029,N_14792);
or U17935 (N_17935,N_14250,N_14470);
and U17936 (N_17936,N_10235,N_13123);
or U17937 (N_17937,N_12542,N_13561);
xnor U17938 (N_17938,N_14677,N_11240);
and U17939 (N_17939,N_12726,N_13550);
nor U17940 (N_17940,N_14874,N_12685);
or U17941 (N_17941,N_11438,N_13414);
xnor U17942 (N_17942,N_14977,N_10300);
and U17943 (N_17943,N_11906,N_13623);
nor U17944 (N_17944,N_14952,N_11106);
and U17945 (N_17945,N_14105,N_10019);
or U17946 (N_17946,N_12528,N_11573);
nand U17947 (N_17947,N_10202,N_14187);
nor U17948 (N_17948,N_12282,N_11700);
nor U17949 (N_17949,N_12157,N_14436);
nand U17950 (N_17950,N_13689,N_14689);
nor U17951 (N_17951,N_14631,N_12747);
xor U17952 (N_17952,N_13513,N_11199);
nor U17953 (N_17953,N_13690,N_13129);
and U17954 (N_17954,N_13655,N_10560);
xor U17955 (N_17955,N_11514,N_14226);
xnor U17956 (N_17956,N_12484,N_13212);
nand U17957 (N_17957,N_14022,N_12040);
and U17958 (N_17958,N_10014,N_12488);
nand U17959 (N_17959,N_13249,N_10453);
nor U17960 (N_17960,N_11506,N_14678);
or U17961 (N_17961,N_10670,N_12188);
nor U17962 (N_17962,N_11708,N_12239);
and U17963 (N_17963,N_10663,N_14562);
nand U17964 (N_17964,N_14240,N_13214);
nand U17965 (N_17965,N_13655,N_11967);
or U17966 (N_17966,N_11674,N_11645);
nor U17967 (N_17967,N_10785,N_11542);
and U17968 (N_17968,N_12967,N_10267);
xor U17969 (N_17969,N_10420,N_13724);
nor U17970 (N_17970,N_12266,N_10489);
or U17971 (N_17971,N_14448,N_13965);
nand U17972 (N_17972,N_14496,N_12370);
and U17973 (N_17973,N_14719,N_14587);
nand U17974 (N_17974,N_10498,N_14245);
nand U17975 (N_17975,N_12619,N_13820);
xnor U17976 (N_17976,N_11975,N_12040);
or U17977 (N_17977,N_11978,N_13741);
nor U17978 (N_17978,N_14261,N_10287);
nand U17979 (N_17979,N_14724,N_13960);
or U17980 (N_17980,N_11955,N_14097);
nor U17981 (N_17981,N_12056,N_14662);
or U17982 (N_17982,N_11371,N_13784);
nand U17983 (N_17983,N_13989,N_14244);
xor U17984 (N_17984,N_10602,N_12292);
and U17985 (N_17985,N_12286,N_13125);
and U17986 (N_17986,N_14209,N_10247);
nor U17987 (N_17987,N_10101,N_10377);
nand U17988 (N_17988,N_14841,N_10817);
xor U17989 (N_17989,N_13212,N_12927);
xor U17990 (N_17990,N_12292,N_13645);
nor U17991 (N_17991,N_11271,N_14865);
and U17992 (N_17992,N_12053,N_11347);
nand U17993 (N_17993,N_12874,N_13999);
xnor U17994 (N_17994,N_13159,N_13916);
xnor U17995 (N_17995,N_10635,N_14825);
xor U17996 (N_17996,N_13177,N_12133);
nand U17997 (N_17997,N_13698,N_12581);
and U17998 (N_17998,N_11774,N_12643);
and U17999 (N_17999,N_12464,N_11073);
nand U18000 (N_18000,N_14993,N_12032);
nand U18001 (N_18001,N_12000,N_10563);
nand U18002 (N_18002,N_13058,N_12035);
xor U18003 (N_18003,N_14367,N_14760);
and U18004 (N_18004,N_13196,N_10408);
and U18005 (N_18005,N_13387,N_13843);
or U18006 (N_18006,N_11840,N_13520);
nand U18007 (N_18007,N_11728,N_12567);
nor U18008 (N_18008,N_12345,N_11543);
and U18009 (N_18009,N_10702,N_12592);
and U18010 (N_18010,N_11540,N_10750);
and U18011 (N_18011,N_13128,N_13497);
or U18012 (N_18012,N_11781,N_14345);
xnor U18013 (N_18013,N_12010,N_13914);
xnor U18014 (N_18014,N_12972,N_11211);
nand U18015 (N_18015,N_10462,N_10420);
nand U18016 (N_18016,N_12105,N_11889);
or U18017 (N_18017,N_10912,N_14029);
or U18018 (N_18018,N_10641,N_12183);
and U18019 (N_18019,N_11831,N_14812);
nand U18020 (N_18020,N_12370,N_11823);
nor U18021 (N_18021,N_10360,N_12800);
nand U18022 (N_18022,N_13153,N_11675);
nand U18023 (N_18023,N_11404,N_11484);
xnor U18024 (N_18024,N_13263,N_13860);
nand U18025 (N_18025,N_10724,N_12759);
or U18026 (N_18026,N_13488,N_12547);
xnor U18027 (N_18027,N_13308,N_13821);
and U18028 (N_18028,N_10915,N_10330);
or U18029 (N_18029,N_12742,N_13889);
or U18030 (N_18030,N_11016,N_12699);
xor U18031 (N_18031,N_10423,N_13704);
and U18032 (N_18032,N_14064,N_11227);
xnor U18033 (N_18033,N_11185,N_10458);
and U18034 (N_18034,N_13239,N_12478);
and U18035 (N_18035,N_10620,N_14173);
nor U18036 (N_18036,N_10296,N_12950);
or U18037 (N_18037,N_13401,N_10428);
xor U18038 (N_18038,N_10752,N_13407);
nand U18039 (N_18039,N_13709,N_10785);
xnor U18040 (N_18040,N_11440,N_12247);
nand U18041 (N_18041,N_10876,N_11671);
nor U18042 (N_18042,N_11447,N_14234);
nor U18043 (N_18043,N_12805,N_13025);
nand U18044 (N_18044,N_12535,N_14531);
or U18045 (N_18045,N_11253,N_11837);
or U18046 (N_18046,N_10519,N_11489);
xor U18047 (N_18047,N_10208,N_12989);
and U18048 (N_18048,N_11384,N_10505);
and U18049 (N_18049,N_13623,N_14858);
xor U18050 (N_18050,N_11297,N_13107);
xnor U18051 (N_18051,N_10682,N_11215);
or U18052 (N_18052,N_10225,N_13732);
and U18053 (N_18053,N_13242,N_14402);
and U18054 (N_18054,N_14150,N_11094);
nand U18055 (N_18055,N_11521,N_10384);
and U18056 (N_18056,N_13163,N_10990);
nor U18057 (N_18057,N_14005,N_11298);
xnor U18058 (N_18058,N_12482,N_11243);
xnor U18059 (N_18059,N_12124,N_10665);
nand U18060 (N_18060,N_13888,N_10257);
nor U18061 (N_18061,N_11368,N_12286);
nor U18062 (N_18062,N_14269,N_11339);
and U18063 (N_18063,N_14639,N_12007);
nor U18064 (N_18064,N_14369,N_10946);
nand U18065 (N_18065,N_12059,N_10701);
and U18066 (N_18066,N_10172,N_10260);
nand U18067 (N_18067,N_11986,N_12232);
or U18068 (N_18068,N_10201,N_13618);
or U18069 (N_18069,N_11373,N_13196);
and U18070 (N_18070,N_10073,N_10928);
or U18071 (N_18071,N_12862,N_10691);
nor U18072 (N_18072,N_13510,N_12015);
nand U18073 (N_18073,N_11962,N_11634);
or U18074 (N_18074,N_14825,N_10845);
nand U18075 (N_18075,N_11295,N_14433);
or U18076 (N_18076,N_10460,N_14454);
or U18077 (N_18077,N_11429,N_10674);
nand U18078 (N_18078,N_11233,N_12822);
xnor U18079 (N_18079,N_12724,N_13271);
nor U18080 (N_18080,N_11961,N_11641);
or U18081 (N_18081,N_10873,N_13592);
xor U18082 (N_18082,N_12964,N_11361);
xor U18083 (N_18083,N_11319,N_10679);
or U18084 (N_18084,N_14012,N_11615);
nor U18085 (N_18085,N_11144,N_14212);
nand U18086 (N_18086,N_12439,N_13829);
xnor U18087 (N_18087,N_13928,N_12328);
or U18088 (N_18088,N_12925,N_12063);
xor U18089 (N_18089,N_10667,N_11180);
nand U18090 (N_18090,N_12973,N_13593);
nand U18091 (N_18091,N_11328,N_12678);
nor U18092 (N_18092,N_11559,N_11900);
nand U18093 (N_18093,N_13467,N_14240);
nand U18094 (N_18094,N_13819,N_11363);
nor U18095 (N_18095,N_13319,N_12574);
nor U18096 (N_18096,N_12180,N_10422);
nand U18097 (N_18097,N_10146,N_13148);
and U18098 (N_18098,N_12565,N_12057);
nor U18099 (N_18099,N_12990,N_14852);
nor U18100 (N_18100,N_14710,N_14590);
or U18101 (N_18101,N_12377,N_14202);
xnor U18102 (N_18102,N_13530,N_14605);
nor U18103 (N_18103,N_14801,N_14798);
nand U18104 (N_18104,N_11414,N_14729);
or U18105 (N_18105,N_13435,N_14126);
nand U18106 (N_18106,N_13265,N_13588);
nand U18107 (N_18107,N_14360,N_14656);
nand U18108 (N_18108,N_13125,N_12296);
nand U18109 (N_18109,N_11279,N_10093);
or U18110 (N_18110,N_10930,N_13376);
nor U18111 (N_18111,N_13343,N_12279);
xnor U18112 (N_18112,N_13052,N_13568);
xnor U18113 (N_18113,N_13481,N_14841);
nor U18114 (N_18114,N_13849,N_13857);
nand U18115 (N_18115,N_12233,N_12909);
xor U18116 (N_18116,N_14832,N_11321);
nand U18117 (N_18117,N_13604,N_10038);
and U18118 (N_18118,N_14060,N_11516);
nand U18119 (N_18119,N_10538,N_10908);
and U18120 (N_18120,N_12644,N_11708);
nor U18121 (N_18121,N_14748,N_12559);
or U18122 (N_18122,N_13973,N_10318);
xnor U18123 (N_18123,N_10050,N_11720);
or U18124 (N_18124,N_11307,N_14813);
and U18125 (N_18125,N_11726,N_14226);
nor U18126 (N_18126,N_10396,N_10630);
and U18127 (N_18127,N_14035,N_12202);
and U18128 (N_18128,N_11596,N_13501);
nor U18129 (N_18129,N_11768,N_12234);
and U18130 (N_18130,N_11900,N_11647);
nand U18131 (N_18131,N_11721,N_12355);
nor U18132 (N_18132,N_13381,N_13833);
or U18133 (N_18133,N_10057,N_10720);
and U18134 (N_18134,N_10640,N_11146);
or U18135 (N_18135,N_14714,N_11952);
nand U18136 (N_18136,N_14051,N_13316);
nand U18137 (N_18137,N_12053,N_14809);
nor U18138 (N_18138,N_11490,N_14897);
nor U18139 (N_18139,N_14567,N_12273);
nor U18140 (N_18140,N_12817,N_10208);
and U18141 (N_18141,N_10338,N_13912);
or U18142 (N_18142,N_11131,N_12171);
or U18143 (N_18143,N_11985,N_14409);
nand U18144 (N_18144,N_14216,N_10484);
nor U18145 (N_18145,N_12956,N_14190);
and U18146 (N_18146,N_10281,N_11784);
nor U18147 (N_18147,N_12258,N_11066);
nor U18148 (N_18148,N_14274,N_11788);
nand U18149 (N_18149,N_14656,N_12436);
nand U18150 (N_18150,N_14156,N_13163);
xnor U18151 (N_18151,N_10461,N_10810);
and U18152 (N_18152,N_12647,N_10447);
nor U18153 (N_18153,N_11945,N_14333);
or U18154 (N_18154,N_13062,N_13191);
nor U18155 (N_18155,N_11931,N_14041);
nand U18156 (N_18156,N_12574,N_10475);
or U18157 (N_18157,N_14471,N_14836);
xor U18158 (N_18158,N_14238,N_13197);
nor U18159 (N_18159,N_11420,N_10779);
or U18160 (N_18160,N_12132,N_11877);
and U18161 (N_18161,N_10018,N_13561);
or U18162 (N_18162,N_14191,N_12760);
or U18163 (N_18163,N_10678,N_11657);
nand U18164 (N_18164,N_10632,N_13074);
nor U18165 (N_18165,N_12592,N_10614);
xnor U18166 (N_18166,N_14294,N_14565);
xor U18167 (N_18167,N_10643,N_10745);
or U18168 (N_18168,N_14790,N_11082);
xnor U18169 (N_18169,N_12780,N_14951);
nand U18170 (N_18170,N_12515,N_14610);
or U18171 (N_18171,N_11178,N_14697);
nand U18172 (N_18172,N_14827,N_13919);
nand U18173 (N_18173,N_10976,N_13454);
nand U18174 (N_18174,N_11125,N_13123);
and U18175 (N_18175,N_11189,N_13959);
xnor U18176 (N_18176,N_10958,N_14913);
nand U18177 (N_18177,N_12649,N_10336);
xnor U18178 (N_18178,N_12322,N_12394);
nor U18179 (N_18179,N_13970,N_10396);
or U18180 (N_18180,N_11204,N_10207);
xor U18181 (N_18181,N_13537,N_10292);
and U18182 (N_18182,N_12060,N_12164);
or U18183 (N_18183,N_13010,N_14981);
or U18184 (N_18184,N_12893,N_10707);
and U18185 (N_18185,N_13176,N_10649);
nand U18186 (N_18186,N_13102,N_12754);
and U18187 (N_18187,N_13498,N_10058);
and U18188 (N_18188,N_10125,N_13466);
nor U18189 (N_18189,N_13375,N_12354);
nor U18190 (N_18190,N_11279,N_12516);
nand U18191 (N_18191,N_14592,N_14310);
nor U18192 (N_18192,N_10595,N_11700);
nand U18193 (N_18193,N_11548,N_10248);
nor U18194 (N_18194,N_11256,N_10217);
and U18195 (N_18195,N_13870,N_10422);
or U18196 (N_18196,N_14806,N_11239);
or U18197 (N_18197,N_14075,N_11215);
and U18198 (N_18198,N_10448,N_10502);
xnor U18199 (N_18199,N_11039,N_12073);
xnor U18200 (N_18200,N_10439,N_10671);
nor U18201 (N_18201,N_11253,N_14894);
nor U18202 (N_18202,N_13284,N_11538);
or U18203 (N_18203,N_12352,N_14060);
xor U18204 (N_18204,N_14204,N_14460);
nor U18205 (N_18205,N_13167,N_11598);
or U18206 (N_18206,N_11332,N_12990);
and U18207 (N_18207,N_10198,N_12341);
and U18208 (N_18208,N_12009,N_10269);
or U18209 (N_18209,N_12007,N_12135);
nand U18210 (N_18210,N_10840,N_12259);
nor U18211 (N_18211,N_10600,N_10166);
xnor U18212 (N_18212,N_14735,N_13769);
nor U18213 (N_18213,N_14212,N_13544);
xnor U18214 (N_18214,N_14123,N_11138);
nor U18215 (N_18215,N_14874,N_14107);
and U18216 (N_18216,N_13499,N_10577);
or U18217 (N_18217,N_14633,N_10481);
nor U18218 (N_18218,N_10526,N_13303);
xnor U18219 (N_18219,N_12374,N_14731);
and U18220 (N_18220,N_13239,N_14830);
or U18221 (N_18221,N_13330,N_13574);
and U18222 (N_18222,N_10988,N_11497);
xnor U18223 (N_18223,N_11894,N_12712);
xnor U18224 (N_18224,N_10407,N_10217);
xor U18225 (N_18225,N_14716,N_14713);
nor U18226 (N_18226,N_11055,N_14264);
nand U18227 (N_18227,N_12062,N_11082);
nand U18228 (N_18228,N_12843,N_13039);
xnor U18229 (N_18229,N_10390,N_13310);
nor U18230 (N_18230,N_13945,N_11235);
xor U18231 (N_18231,N_10778,N_14077);
or U18232 (N_18232,N_10270,N_14777);
nand U18233 (N_18233,N_14760,N_11026);
nand U18234 (N_18234,N_12382,N_14847);
nand U18235 (N_18235,N_11807,N_10038);
nor U18236 (N_18236,N_10298,N_14464);
nand U18237 (N_18237,N_14539,N_13512);
nor U18238 (N_18238,N_13917,N_10044);
nor U18239 (N_18239,N_14741,N_13989);
xor U18240 (N_18240,N_10188,N_10662);
or U18241 (N_18241,N_14321,N_14063);
nand U18242 (N_18242,N_12646,N_10662);
nand U18243 (N_18243,N_10131,N_13777);
xor U18244 (N_18244,N_11230,N_14293);
nor U18245 (N_18245,N_14820,N_13565);
or U18246 (N_18246,N_12550,N_10709);
nor U18247 (N_18247,N_10645,N_13908);
xnor U18248 (N_18248,N_13720,N_14830);
or U18249 (N_18249,N_12726,N_11226);
nand U18250 (N_18250,N_10159,N_14576);
and U18251 (N_18251,N_10691,N_11005);
or U18252 (N_18252,N_12646,N_13589);
nand U18253 (N_18253,N_14808,N_10440);
and U18254 (N_18254,N_13395,N_11880);
or U18255 (N_18255,N_10038,N_12326);
or U18256 (N_18256,N_14078,N_12485);
xnor U18257 (N_18257,N_10209,N_12545);
or U18258 (N_18258,N_10214,N_13618);
nor U18259 (N_18259,N_13449,N_12864);
and U18260 (N_18260,N_14052,N_14836);
nor U18261 (N_18261,N_13443,N_12981);
or U18262 (N_18262,N_12671,N_11491);
xor U18263 (N_18263,N_13458,N_10792);
nand U18264 (N_18264,N_11358,N_11090);
nand U18265 (N_18265,N_10445,N_13439);
and U18266 (N_18266,N_13100,N_12732);
xnor U18267 (N_18267,N_11331,N_14121);
and U18268 (N_18268,N_13531,N_14343);
nand U18269 (N_18269,N_13307,N_10221);
nor U18270 (N_18270,N_14912,N_11245);
and U18271 (N_18271,N_11382,N_13764);
and U18272 (N_18272,N_11325,N_13166);
nor U18273 (N_18273,N_11009,N_14405);
xnor U18274 (N_18274,N_10212,N_13231);
and U18275 (N_18275,N_10587,N_11180);
nor U18276 (N_18276,N_13483,N_12724);
xnor U18277 (N_18277,N_13129,N_11796);
xnor U18278 (N_18278,N_14612,N_14450);
xor U18279 (N_18279,N_12888,N_12872);
and U18280 (N_18280,N_10844,N_11406);
nand U18281 (N_18281,N_12400,N_10097);
nand U18282 (N_18282,N_11142,N_13759);
nand U18283 (N_18283,N_12912,N_14253);
xor U18284 (N_18284,N_11630,N_11797);
or U18285 (N_18285,N_11418,N_12222);
or U18286 (N_18286,N_11644,N_10912);
xor U18287 (N_18287,N_11473,N_13889);
or U18288 (N_18288,N_10386,N_12177);
and U18289 (N_18289,N_14571,N_14679);
or U18290 (N_18290,N_13818,N_11930);
or U18291 (N_18291,N_11846,N_11229);
or U18292 (N_18292,N_13819,N_12832);
nor U18293 (N_18293,N_10178,N_11219);
nor U18294 (N_18294,N_12305,N_12947);
or U18295 (N_18295,N_12928,N_14873);
nand U18296 (N_18296,N_11550,N_10152);
nor U18297 (N_18297,N_13613,N_13602);
nor U18298 (N_18298,N_11147,N_13325);
or U18299 (N_18299,N_13041,N_12393);
nor U18300 (N_18300,N_12970,N_10128);
and U18301 (N_18301,N_10572,N_13754);
xor U18302 (N_18302,N_14221,N_13778);
nor U18303 (N_18303,N_12949,N_11125);
or U18304 (N_18304,N_11187,N_10257);
and U18305 (N_18305,N_14650,N_11838);
nor U18306 (N_18306,N_10912,N_12954);
or U18307 (N_18307,N_10384,N_12412);
or U18308 (N_18308,N_13514,N_11693);
or U18309 (N_18309,N_14953,N_11216);
or U18310 (N_18310,N_14061,N_12973);
xnor U18311 (N_18311,N_12789,N_10427);
xnor U18312 (N_18312,N_12917,N_14420);
xor U18313 (N_18313,N_14418,N_11513);
nand U18314 (N_18314,N_11194,N_10634);
xnor U18315 (N_18315,N_10603,N_10320);
nand U18316 (N_18316,N_13357,N_11713);
xnor U18317 (N_18317,N_14486,N_13970);
and U18318 (N_18318,N_10722,N_13390);
nand U18319 (N_18319,N_12279,N_12835);
or U18320 (N_18320,N_11965,N_11370);
and U18321 (N_18321,N_10054,N_10800);
nor U18322 (N_18322,N_14343,N_11822);
xnor U18323 (N_18323,N_10939,N_12648);
xnor U18324 (N_18324,N_11550,N_12501);
nor U18325 (N_18325,N_11233,N_12716);
and U18326 (N_18326,N_14807,N_11455);
or U18327 (N_18327,N_10052,N_11340);
and U18328 (N_18328,N_14930,N_13552);
nand U18329 (N_18329,N_11314,N_10308);
nand U18330 (N_18330,N_12947,N_11464);
nand U18331 (N_18331,N_11813,N_14608);
xor U18332 (N_18332,N_14543,N_13384);
and U18333 (N_18333,N_12529,N_10189);
and U18334 (N_18334,N_10154,N_10092);
nand U18335 (N_18335,N_14810,N_14232);
nand U18336 (N_18336,N_13854,N_12906);
xor U18337 (N_18337,N_13681,N_13436);
or U18338 (N_18338,N_11197,N_12014);
nand U18339 (N_18339,N_13953,N_14134);
xor U18340 (N_18340,N_12966,N_12758);
and U18341 (N_18341,N_10785,N_12774);
or U18342 (N_18342,N_12092,N_11031);
xor U18343 (N_18343,N_10971,N_11521);
and U18344 (N_18344,N_11424,N_14749);
nor U18345 (N_18345,N_13528,N_10960);
nor U18346 (N_18346,N_11437,N_10208);
and U18347 (N_18347,N_11516,N_11621);
or U18348 (N_18348,N_11690,N_12985);
nor U18349 (N_18349,N_13310,N_14446);
and U18350 (N_18350,N_13269,N_13360);
or U18351 (N_18351,N_13035,N_11702);
nor U18352 (N_18352,N_12669,N_10480);
xor U18353 (N_18353,N_10441,N_11319);
nor U18354 (N_18354,N_10993,N_11867);
or U18355 (N_18355,N_13364,N_13956);
or U18356 (N_18356,N_12126,N_12555);
nand U18357 (N_18357,N_12602,N_10227);
nand U18358 (N_18358,N_12537,N_12155);
or U18359 (N_18359,N_12598,N_11271);
and U18360 (N_18360,N_14989,N_12855);
or U18361 (N_18361,N_12466,N_10160);
and U18362 (N_18362,N_11040,N_11933);
or U18363 (N_18363,N_10898,N_12838);
or U18364 (N_18364,N_10436,N_10758);
nand U18365 (N_18365,N_11384,N_11992);
nand U18366 (N_18366,N_14563,N_12850);
nand U18367 (N_18367,N_10803,N_13320);
nor U18368 (N_18368,N_12010,N_13389);
nor U18369 (N_18369,N_12248,N_12658);
nand U18370 (N_18370,N_10532,N_12958);
and U18371 (N_18371,N_10791,N_14147);
nor U18372 (N_18372,N_14221,N_11355);
xnor U18373 (N_18373,N_14646,N_12278);
nand U18374 (N_18374,N_12684,N_13010);
nor U18375 (N_18375,N_11031,N_14639);
or U18376 (N_18376,N_12048,N_12457);
nor U18377 (N_18377,N_13613,N_12352);
xor U18378 (N_18378,N_13854,N_13349);
nor U18379 (N_18379,N_13942,N_11813);
and U18380 (N_18380,N_11028,N_10253);
and U18381 (N_18381,N_12206,N_10714);
or U18382 (N_18382,N_11464,N_12454);
nand U18383 (N_18383,N_13539,N_14330);
xor U18384 (N_18384,N_14271,N_12671);
and U18385 (N_18385,N_10345,N_12742);
and U18386 (N_18386,N_14313,N_13185);
nand U18387 (N_18387,N_12663,N_14660);
or U18388 (N_18388,N_14231,N_13422);
or U18389 (N_18389,N_12311,N_11110);
nand U18390 (N_18390,N_11309,N_11016);
nor U18391 (N_18391,N_12099,N_13295);
and U18392 (N_18392,N_11654,N_10658);
nand U18393 (N_18393,N_12795,N_14649);
nand U18394 (N_18394,N_10133,N_10215);
or U18395 (N_18395,N_12785,N_13475);
nand U18396 (N_18396,N_10944,N_11082);
and U18397 (N_18397,N_14833,N_10238);
nand U18398 (N_18398,N_13297,N_10843);
xor U18399 (N_18399,N_13830,N_14663);
nand U18400 (N_18400,N_10188,N_14055);
nor U18401 (N_18401,N_11662,N_14948);
xnor U18402 (N_18402,N_14915,N_10846);
nor U18403 (N_18403,N_13476,N_12010);
and U18404 (N_18404,N_12309,N_11316);
xor U18405 (N_18405,N_12466,N_12052);
nand U18406 (N_18406,N_11626,N_13277);
xor U18407 (N_18407,N_11182,N_10363);
nand U18408 (N_18408,N_13070,N_13494);
nor U18409 (N_18409,N_13198,N_14147);
or U18410 (N_18410,N_14721,N_12511);
or U18411 (N_18411,N_10338,N_11641);
and U18412 (N_18412,N_12301,N_14890);
nand U18413 (N_18413,N_11213,N_11076);
xnor U18414 (N_18414,N_14216,N_14981);
nor U18415 (N_18415,N_11806,N_10015);
xor U18416 (N_18416,N_14400,N_12538);
nor U18417 (N_18417,N_14006,N_10272);
or U18418 (N_18418,N_13518,N_14695);
or U18419 (N_18419,N_10495,N_11167);
or U18420 (N_18420,N_10678,N_12392);
and U18421 (N_18421,N_14318,N_13642);
and U18422 (N_18422,N_12362,N_13307);
nand U18423 (N_18423,N_12379,N_12992);
xnor U18424 (N_18424,N_13705,N_12980);
or U18425 (N_18425,N_10299,N_12626);
nand U18426 (N_18426,N_13235,N_10725);
nand U18427 (N_18427,N_13938,N_14143);
nor U18428 (N_18428,N_14001,N_13575);
xnor U18429 (N_18429,N_11125,N_10925);
or U18430 (N_18430,N_14716,N_12821);
xnor U18431 (N_18431,N_13963,N_14908);
or U18432 (N_18432,N_11257,N_14562);
or U18433 (N_18433,N_13090,N_10444);
xnor U18434 (N_18434,N_12718,N_12987);
and U18435 (N_18435,N_14316,N_14836);
nand U18436 (N_18436,N_14136,N_10193);
nor U18437 (N_18437,N_11474,N_12975);
nor U18438 (N_18438,N_11682,N_14258);
or U18439 (N_18439,N_10854,N_13671);
and U18440 (N_18440,N_14072,N_11637);
nand U18441 (N_18441,N_10878,N_12833);
and U18442 (N_18442,N_11149,N_14486);
or U18443 (N_18443,N_11290,N_12688);
nor U18444 (N_18444,N_10744,N_10376);
and U18445 (N_18445,N_10558,N_11710);
xnor U18446 (N_18446,N_13589,N_10278);
nor U18447 (N_18447,N_14498,N_10806);
and U18448 (N_18448,N_12937,N_10842);
and U18449 (N_18449,N_10788,N_10833);
and U18450 (N_18450,N_10812,N_10202);
nor U18451 (N_18451,N_12901,N_11128);
nor U18452 (N_18452,N_14778,N_13330);
nor U18453 (N_18453,N_12994,N_12657);
nor U18454 (N_18454,N_10987,N_13813);
or U18455 (N_18455,N_12196,N_12347);
or U18456 (N_18456,N_10299,N_14438);
nand U18457 (N_18457,N_14253,N_11673);
nor U18458 (N_18458,N_14311,N_12599);
or U18459 (N_18459,N_10083,N_14711);
xor U18460 (N_18460,N_13383,N_13194);
nor U18461 (N_18461,N_13718,N_10822);
xnor U18462 (N_18462,N_13608,N_12422);
and U18463 (N_18463,N_11349,N_14982);
and U18464 (N_18464,N_12606,N_10915);
xnor U18465 (N_18465,N_10098,N_10973);
xnor U18466 (N_18466,N_13601,N_13823);
nor U18467 (N_18467,N_14067,N_11394);
or U18468 (N_18468,N_10346,N_13134);
nor U18469 (N_18469,N_14725,N_12703);
nor U18470 (N_18470,N_14155,N_14896);
and U18471 (N_18471,N_12574,N_10811);
nor U18472 (N_18472,N_12147,N_13612);
and U18473 (N_18473,N_13119,N_10846);
nand U18474 (N_18474,N_10228,N_11816);
and U18475 (N_18475,N_14005,N_13911);
or U18476 (N_18476,N_10649,N_13661);
nor U18477 (N_18477,N_10305,N_11266);
or U18478 (N_18478,N_13221,N_10513);
xnor U18479 (N_18479,N_14720,N_12822);
or U18480 (N_18480,N_14717,N_11952);
xor U18481 (N_18481,N_13759,N_14413);
nand U18482 (N_18482,N_14306,N_11290);
and U18483 (N_18483,N_10842,N_10924);
and U18484 (N_18484,N_11398,N_14054);
nand U18485 (N_18485,N_13073,N_13542);
nand U18486 (N_18486,N_12809,N_14611);
and U18487 (N_18487,N_14679,N_11894);
xor U18488 (N_18488,N_11024,N_11402);
nand U18489 (N_18489,N_11529,N_14853);
and U18490 (N_18490,N_14423,N_11140);
xor U18491 (N_18491,N_11552,N_10275);
and U18492 (N_18492,N_11561,N_13611);
or U18493 (N_18493,N_12583,N_10391);
xnor U18494 (N_18494,N_12127,N_14575);
xor U18495 (N_18495,N_13270,N_11357);
or U18496 (N_18496,N_11462,N_14913);
nand U18497 (N_18497,N_10525,N_10625);
nand U18498 (N_18498,N_14968,N_11075);
or U18499 (N_18499,N_12015,N_11794);
xnor U18500 (N_18500,N_11852,N_12856);
nor U18501 (N_18501,N_14952,N_11970);
nand U18502 (N_18502,N_14677,N_11122);
or U18503 (N_18503,N_13225,N_10974);
or U18504 (N_18504,N_13445,N_14318);
nand U18505 (N_18505,N_11702,N_14146);
xor U18506 (N_18506,N_12703,N_10274);
nand U18507 (N_18507,N_13925,N_13433);
nor U18508 (N_18508,N_10977,N_10713);
and U18509 (N_18509,N_11478,N_10660);
xnor U18510 (N_18510,N_13371,N_10844);
and U18511 (N_18511,N_11191,N_14381);
nor U18512 (N_18512,N_10199,N_13861);
nand U18513 (N_18513,N_10000,N_10262);
nand U18514 (N_18514,N_13686,N_11190);
xnor U18515 (N_18515,N_10621,N_14501);
xnor U18516 (N_18516,N_12950,N_12856);
nor U18517 (N_18517,N_13451,N_12334);
nor U18518 (N_18518,N_14839,N_13236);
nand U18519 (N_18519,N_14454,N_10164);
nand U18520 (N_18520,N_13460,N_12992);
or U18521 (N_18521,N_11463,N_13814);
nand U18522 (N_18522,N_13459,N_14276);
xnor U18523 (N_18523,N_12070,N_14579);
xnor U18524 (N_18524,N_12166,N_11494);
and U18525 (N_18525,N_10406,N_13379);
xnor U18526 (N_18526,N_13262,N_12186);
xnor U18527 (N_18527,N_10946,N_10813);
nand U18528 (N_18528,N_13861,N_14356);
nand U18529 (N_18529,N_14444,N_11008);
nand U18530 (N_18530,N_13572,N_11696);
and U18531 (N_18531,N_10196,N_12259);
xor U18532 (N_18532,N_11546,N_12899);
and U18533 (N_18533,N_10893,N_13729);
nand U18534 (N_18534,N_11611,N_13673);
xor U18535 (N_18535,N_12908,N_13279);
and U18536 (N_18536,N_11697,N_13919);
nor U18537 (N_18537,N_14610,N_13505);
nand U18538 (N_18538,N_10107,N_14431);
nand U18539 (N_18539,N_10432,N_14323);
or U18540 (N_18540,N_11808,N_10213);
and U18541 (N_18541,N_10412,N_11553);
nand U18542 (N_18542,N_10867,N_11858);
or U18543 (N_18543,N_13063,N_10395);
nor U18544 (N_18544,N_10088,N_14478);
or U18545 (N_18545,N_14271,N_11851);
or U18546 (N_18546,N_13585,N_11616);
or U18547 (N_18547,N_11992,N_11479);
and U18548 (N_18548,N_11930,N_13585);
and U18549 (N_18549,N_14556,N_10606);
xor U18550 (N_18550,N_11052,N_10873);
or U18551 (N_18551,N_11255,N_11259);
xnor U18552 (N_18552,N_11634,N_10999);
nor U18553 (N_18553,N_11362,N_14291);
and U18554 (N_18554,N_11105,N_14689);
nand U18555 (N_18555,N_10448,N_10198);
or U18556 (N_18556,N_10367,N_14521);
or U18557 (N_18557,N_12571,N_14157);
or U18558 (N_18558,N_10355,N_14489);
and U18559 (N_18559,N_12984,N_11085);
nor U18560 (N_18560,N_11850,N_11545);
xnor U18561 (N_18561,N_14348,N_11100);
xor U18562 (N_18562,N_12259,N_13915);
xor U18563 (N_18563,N_10839,N_11439);
and U18564 (N_18564,N_13951,N_13971);
nor U18565 (N_18565,N_14360,N_14353);
nor U18566 (N_18566,N_10922,N_11750);
and U18567 (N_18567,N_12674,N_14168);
nor U18568 (N_18568,N_10027,N_14188);
nor U18569 (N_18569,N_10871,N_14876);
or U18570 (N_18570,N_13561,N_10086);
and U18571 (N_18571,N_12632,N_10428);
nand U18572 (N_18572,N_13484,N_14296);
nand U18573 (N_18573,N_14006,N_11014);
nand U18574 (N_18574,N_10560,N_13814);
xor U18575 (N_18575,N_12368,N_14794);
or U18576 (N_18576,N_13469,N_12863);
xnor U18577 (N_18577,N_11197,N_12136);
xnor U18578 (N_18578,N_11182,N_10917);
nor U18579 (N_18579,N_14541,N_12384);
nor U18580 (N_18580,N_11807,N_14404);
xnor U18581 (N_18581,N_11688,N_10924);
xor U18582 (N_18582,N_11947,N_11205);
nand U18583 (N_18583,N_13313,N_10541);
nor U18584 (N_18584,N_13265,N_13563);
or U18585 (N_18585,N_14259,N_13795);
and U18586 (N_18586,N_12580,N_14003);
and U18587 (N_18587,N_11866,N_11898);
nor U18588 (N_18588,N_13586,N_11499);
or U18589 (N_18589,N_10520,N_14272);
nand U18590 (N_18590,N_14196,N_14853);
or U18591 (N_18591,N_10571,N_13399);
and U18592 (N_18592,N_10284,N_14858);
nand U18593 (N_18593,N_14209,N_12170);
and U18594 (N_18594,N_14149,N_12334);
or U18595 (N_18595,N_10455,N_14744);
xor U18596 (N_18596,N_11015,N_13255);
xnor U18597 (N_18597,N_11291,N_12030);
or U18598 (N_18598,N_13040,N_10602);
nand U18599 (N_18599,N_14613,N_13055);
and U18600 (N_18600,N_11085,N_10446);
xnor U18601 (N_18601,N_10818,N_13971);
xor U18602 (N_18602,N_13685,N_14069);
or U18603 (N_18603,N_11728,N_13386);
xor U18604 (N_18604,N_10050,N_11197);
and U18605 (N_18605,N_13594,N_10951);
or U18606 (N_18606,N_12749,N_11250);
or U18607 (N_18607,N_11874,N_13050);
and U18608 (N_18608,N_11620,N_14752);
nand U18609 (N_18609,N_13158,N_14940);
nor U18610 (N_18610,N_12899,N_12767);
nor U18611 (N_18611,N_13698,N_11701);
nand U18612 (N_18612,N_10098,N_12156);
or U18613 (N_18613,N_14131,N_14058);
nand U18614 (N_18614,N_14075,N_10603);
and U18615 (N_18615,N_12684,N_10898);
and U18616 (N_18616,N_11456,N_11327);
or U18617 (N_18617,N_10776,N_10804);
or U18618 (N_18618,N_12108,N_13432);
xor U18619 (N_18619,N_12856,N_11370);
nand U18620 (N_18620,N_13800,N_12103);
or U18621 (N_18621,N_11000,N_13361);
and U18622 (N_18622,N_13545,N_11758);
nand U18623 (N_18623,N_14224,N_14038);
nor U18624 (N_18624,N_14413,N_13828);
or U18625 (N_18625,N_12376,N_10145);
nor U18626 (N_18626,N_11434,N_13083);
nor U18627 (N_18627,N_11879,N_11097);
or U18628 (N_18628,N_11712,N_14351);
nor U18629 (N_18629,N_12281,N_10098);
nand U18630 (N_18630,N_14797,N_10088);
xnor U18631 (N_18631,N_11197,N_11893);
or U18632 (N_18632,N_14470,N_12178);
or U18633 (N_18633,N_12040,N_10337);
xor U18634 (N_18634,N_13720,N_13551);
or U18635 (N_18635,N_13984,N_10508);
nand U18636 (N_18636,N_12055,N_13983);
and U18637 (N_18637,N_11648,N_10807);
nand U18638 (N_18638,N_11140,N_13992);
nand U18639 (N_18639,N_13453,N_11371);
nand U18640 (N_18640,N_12848,N_12673);
or U18641 (N_18641,N_11544,N_13517);
or U18642 (N_18642,N_14900,N_11510);
xnor U18643 (N_18643,N_10025,N_11238);
or U18644 (N_18644,N_12419,N_10631);
or U18645 (N_18645,N_11497,N_12922);
and U18646 (N_18646,N_10993,N_11548);
and U18647 (N_18647,N_10056,N_13310);
nand U18648 (N_18648,N_12107,N_13973);
and U18649 (N_18649,N_11898,N_14310);
xor U18650 (N_18650,N_12419,N_12591);
nor U18651 (N_18651,N_13068,N_11319);
and U18652 (N_18652,N_11899,N_14043);
and U18653 (N_18653,N_13132,N_12524);
xor U18654 (N_18654,N_13192,N_10519);
nand U18655 (N_18655,N_10276,N_12502);
or U18656 (N_18656,N_11422,N_10804);
or U18657 (N_18657,N_14230,N_14640);
and U18658 (N_18658,N_14074,N_12310);
xor U18659 (N_18659,N_14516,N_13340);
nor U18660 (N_18660,N_10760,N_12460);
or U18661 (N_18661,N_12855,N_13043);
or U18662 (N_18662,N_14143,N_12186);
nand U18663 (N_18663,N_12044,N_13900);
or U18664 (N_18664,N_11422,N_13476);
or U18665 (N_18665,N_13036,N_11731);
or U18666 (N_18666,N_11193,N_11715);
nor U18667 (N_18667,N_11776,N_11580);
or U18668 (N_18668,N_14217,N_10850);
or U18669 (N_18669,N_14944,N_12032);
and U18670 (N_18670,N_11436,N_10272);
nand U18671 (N_18671,N_12661,N_10024);
nor U18672 (N_18672,N_10773,N_10566);
and U18673 (N_18673,N_14585,N_13090);
and U18674 (N_18674,N_13717,N_14559);
xor U18675 (N_18675,N_10777,N_11717);
nand U18676 (N_18676,N_10313,N_13622);
nand U18677 (N_18677,N_10714,N_13859);
and U18678 (N_18678,N_14160,N_12108);
xor U18679 (N_18679,N_11885,N_13643);
nand U18680 (N_18680,N_13696,N_11288);
or U18681 (N_18681,N_11555,N_10541);
and U18682 (N_18682,N_13536,N_10800);
and U18683 (N_18683,N_14752,N_13994);
nand U18684 (N_18684,N_13912,N_12113);
and U18685 (N_18685,N_14350,N_12527);
or U18686 (N_18686,N_11400,N_12209);
nand U18687 (N_18687,N_12393,N_10702);
and U18688 (N_18688,N_11802,N_10120);
nor U18689 (N_18689,N_14887,N_10594);
xor U18690 (N_18690,N_14054,N_10736);
nand U18691 (N_18691,N_14334,N_11697);
xor U18692 (N_18692,N_10514,N_13963);
nand U18693 (N_18693,N_14221,N_13555);
xnor U18694 (N_18694,N_14091,N_12673);
nand U18695 (N_18695,N_14238,N_10147);
nand U18696 (N_18696,N_13610,N_12354);
nand U18697 (N_18697,N_12918,N_10305);
or U18698 (N_18698,N_11013,N_11466);
nor U18699 (N_18699,N_14853,N_11383);
xor U18700 (N_18700,N_14958,N_11475);
nor U18701 (N_18701,N_12453,N_11272);
or U18702 (N_18702,N_14850,N_12110);
xor U18703 (N_18703,N_12011,N_13983);
and U18704 (N_18704,N_14426,N_14373);
or U18705 (N_18705,N_10769,N_12390);
xnor U18706 (N_18706,N_11555,N_12918);
xnor U18707 (N_18707,N_10063,N_14397);
and U18708 (N_18708,N_11989,N_14881);
or U18709 (N_18709,N_11959,N_14278);
or U18710 (N_18710,N_14955,N_11811);
or U18711 (N_18711,N_14409,N_12868);
nand U18712 (N_18712,N_12510,N_14360);
xor U18713 (N_18713,N_12678,N_10147);
nor U18714 (N_18714,N_14564,N_14804);
nand U18715 (N_18715,N_13933,N_13584);
nor U18716 (N_18716,N_12453,N_12563);
nor U18717 (N_18717,N_13111,N_14275);
nand U18718 (N_18718,N_12124,N_14062);
nor U18719 (N_18719,N_14895,N_13957);
nor U18720 (N_18720,N_12154,N_10946);
nor U18721 (N_18721,N_14251,N_13886);
xnor U18722 (N_18722,N_11955,N_12998);
nor U18723 (N_18723,N_13191,N_11838);
and U18724 (N_18724,N_13609,N_12915);
nor U18725 (N_18725,N_13540,N_14187);
xnor U18726 (N_18726,N_13685,N_14116);
xor U18727 (N_18727,N_10942,N_13596);
nor U18728 (N_18728,N_11583,N_13937);
or U18729 (N_18729,N_13251,N_14122);
xor U18730 (N_18730,N_10492,N_10081);
xor U18731 (N_18731,N_10202,N_13069);
xnor U18732 (N_18732,N_10596,N_13901);
or U18733 (N_18733,N_10662,N_11745);
and U18734 (N_18734,N_11805,N_14056);
and U18735 (N_18735,N_10092,N_12291);
or U18736 (N_18736,N_11576,N_13433);
or U18737 (N_18737,N_14879,N_14810);
and U18738 (N_18738,N_10837,N_14873);
or U18739 (N_18739,N_13219,N_13437);
xnor U18740 (N_18740,N_11472,N_11579);
or U18741 (N_18741,N_11623,N_13924);
and U18742 (N_18742,N_11895,N_10486);
nor U18743 (N_18743,N_14394,N_12912);
or U18744 (N_18744,N_14495,N_12542);
nor U18745 (N_18745,N_10668,N_11667);
nor U18746 (N_18746,N_12979,N_12694);
nand U18747 (N_18747,N_10293,N_12437);
nor U18748 (N_18748,N_12562,N_11458);
xor U18749 (N_18749,N_14484,N_11427);
and U18750 (N_18750,N_12421,N_13601);
nand U18751 (N_18751,N_11264,N_14730);
or U18752 (N_18752,N_13410,N_12486);
and U18753 (N_18753,N_12949,N_10123);
xor U18754 (N_18754,N_14315,N_11113);
and U18755 (N_18755,N_12151,N_10831);
or U18756 (N_18756,N_11617,N_14137);
nor U18757 (N_18757,N_10254,N_10207);
nor U18758 (N_18758,N_11327,N_14906);
xnor U18759 (N_18759,N_12714,N_10948);
xnor U18760 (N_18760,N_11633,N_12943);
nor U18761 (N_18761,N_11232,N_12012);
nor U18762 (N_18762,N_12693,N_13619);
or U18763 (N_18763,N_12954,N_14469);
nor U18764 (N_18764,N_10439,N_12028);
or U18765 (N_18765,N_13509,N_11954);
and U18766 (N_18766,N_11766,N_10611);
nand U18767 (N_18767,N_12895,N_12415);
nor U18768 (N_18768,N_10997,N_12948);
and U18769 (N_18769,N_10751,N_14677);
xnor U18770 (N_18770,N_10267,N_14409);
nand U18771 (N_18771,N_10764,N_10499);
nand U18772 (N_18772,N_11983,N_14857);
or U18773 (N_18773,N_12649,N_12405);
or U18774 (N_18774,N_13514,N_13180);
nor U18775 (N_18775,N_10074,N_14644);
nand U18776 (N_18776,N_10860,N_12317);
xnor U18777 (N_18777,N_10362,N_10963);
nand U18778 (N_18778,N_13208,N_12802);
nand U18779 (N_18779,N_12867,N_12014);
and U18780 (N_18780,N_13942,N_10753);
and U18781 (N_18781,N_10345,N_11654);
nand U18782 (N_18782,N_12054,N_13335);
nand U18783 (N_18783,N_10647,N_10061);
and U18784 (N_18784,N_14035,N_10569);
xor U18785 (N_18785,N_10417,N_10441);
nand U18786 (N_18786,N_12053,N_10162);
nor U18787 (N_18787,N_12855,N_12415);
nor U18788 (N_18788,N_13214,N_13262);
or U18789 (N_18789,N_12205,N_11634);
xor U18790 (N_18790,N_11934,N_12578);
xor U18791 (N_18791,N_11690,N_12005);
xnor U18792 (N_18792,N_14944,N_13690);
xor U18793 (N_18793,N_14347,N_14940);
xnor U18794 (N_18794,N_11797,N_10696);
nor U18795 (N_18795,N_13561,N_14956);
nor U18796 (N_18796,N_13218,N_13408);
or U18797 (N_18797,N_10126,N_13887);
or U18798 (N_18798,N_10499,N_14786);
and U18799 (N_18799,N_13345,N_10017);
and U18800 (N_18800,N_12334,N_11735);
nor U18801 (N_18801,N_10555,N_11095);
xnor U18802 (N_18802,N_12080,N_14775);
xor U18803 (N_18803,N_10644,N_13135);
and U18804 (N_18804,N_12477,N_13638);
nor U18805 (N_18805,N_10222,N_10617);
nand U18806 (N_18806,N_14728,N_11176);
xnor U18807 (N_18807,N_13853,N_14671);
or U18808 (N_18808,N_11502,N_11772);
nand U18809 (N_18809,N_11600,N_14857);
nor U18810 (N_18810,N_13032,N_12383);
or U18811 (N_18811,N_14898,N_13033);
nor U18812 (N_18812,N_13279,N_14405);
xor U18813 (N_18813,N_13574,N_10766);
and U18814 (N_18814,N_10325,N_11526);
nor U18815 (N_18815,N_14396,N_13633);
nand U18816 (N_18816,N_11592,N_13863);
nor U18817 (N_18817,N_11922,N_14446);
nand U18818 (N_18818,N_10810,N_14679);
and U18819 (N_18819,N_11866,N_11989);
nand U18820 (N_18820,N_14900,N_14800);
xnor U18821 (N_18821,N_14964,N_13002);
nor U18822 (N_18822,N_14363,N_13313);
nand U18823 (N_18823,N_13418,N_10427);
or U18824 (N_18824,N_12185,N_14512);
nor U18825 (N_18825,N_11738,N_12201);
or U18826 (N_18826,N_14588,N_12771);
nor U18827 (N_18827,N_10008,N_13937);
nor U18828 (N_18828,N_12290,N_13894);
xor U18829 (N_18829,N_11273,N_14788);
xor U18830 (N_18830,N_13788,N_13184);
xnor U18831 (N_18831,N_11710,N_10229);
xor U18832 (N_18832,N_10689,N_10820);
xor U18833 (N_18833,N_11436,N_14645);
nor U18834 (N_18834,N_12998,N_11156);
and U18835 (N_18835,N_13342,N_10560);
nor U18836 (N_18836,N_12093,N_10117);
or U18837 (N_18837,N_12707,N_10763);
nand U18838 (N_18838,N_14917,N_12745);
nand U18839 (N_18839,N_12238,N_12635);
and U18840 (N_18840,N_13857,N_14818);
nand U18841 (N_18841,N_14899,N_11835);
nand U18842 (N_18842,N_11852,N_12784);
and U18843 (N_18843,N_12425,N_12489);
and U18844 (N_18844,N_12973,N_14680);
or U18845 (N_18845,N_11619,N_13446);
and U18846 (N_18846,N_14246,N_14784);
and U18847 (N_18847,N_12261,N_13492);
nor U18848 (N_18848,N_13513,N_10036);
nor U18849 (N_18849,N_11338,N_11292);
xor U18850 (N_18850,N_11530,N_14545);
and U18851 (N_18851,N_14097,N_14326);
and U18852 (N_18852,N_10906,N_14726);
or U18853 (N_18853,N_12864,N_12492);
xnor U18854 (N_18854,N_13756,N_12343);
xnor U18855 (N_18855,N_13803,N_13389);
nor U18856 (N_18856,N_11316,N_10739);
nor U18857 (N_18857,N_13271,N_14631);
and U18858 (N_18858,N_14529,N_13353);
or U18859 (N_18859,N_13517,N_13991);
xnor U18860 (N_18860,N_10208,N_12335);
nand U18861 (N_18861,N_11086,N_11183);
or U18862 (N_18862,N_14151,N_13047);
xnor U18863 (N_18863,N_12452,N_14893);
or U18864 (N_18864,N_14686,N_12727);
nor U18865 (N_18865,N_14477,N_14421);
xor U18866 (N_18866,N_11539,N_12390);
nor U18867 (N_18867,N_12067,N_12913);
and U18868 (N_18868,N_13299,N_13388);
or U18869 (N_18869,N_12940,N_12290);
xnor U18870 (N_18870,N_13602,N_13371);
nor U18871 (N_18871,N_12412,N_14215);
xnor U18872 (N_18872,N_11455,N_14334);
nand U18873 (N_18873,N_10526,N_11221);
or U18874 (N_18874,N_14592,N_14101);
or U18875 (N_18875,N_11016,N_13389);
nor U18876 (N_18876,N_12440,N_13140);
xor U18877 (N_18877,N_12224,N_13565);
nor U18878 (N_18878,N_11418,N_14846);
nor U18879 (N_18879,N_13461,N_12245);
nand U18880 (N_18880,N_12939,N_11708);
xor U18881 (N_18881,N_12548,N_12607);
nor U18882 (N_18882,N_12602,N_10801);
or U18883 (N_18883,N_10328,N_10953);
xnor U18884 (N_18884,N_11098,N_10901);
and U18885 (N_18885,N_10473,N_10542);
xor U18886 (N_18886,N_14345,N_12633);
xor U18887 (N_18887,N_12303,N_11791);
xnor U18888 (N_18888,N_14780,N_11481);
xor U18889 (N_18889,N_14069,N_14828);
and U18890 (N_18890,N_13507,N_14469);
or U18891 (N_18891,N_11527,N_14114);
xor U18892 (N_18892,N_13529,N_11322);
nor U18893 (N_18893,N_12490,N_13260);
or U18894 (N_18894,N_12507,N_10797);
or U18895 (N_18895,N_11150,N_10877);
and U18896 (N_18896,N_10061,N_10454);
xor U18897 (N_18897,N_10368,N_10232);
and U18898 (N_18898,N_10923,N_11533);
xor U18899 (N_18899,N_12032,N_11826);
or U18900 (N_18900,N_12294,N_12386);
and U18901 (N_18901,N_11088,N_13185);
nor U18902 (N_18902,N_14856,N_14497);
nor U18903 (N_18903,N_10542,N_12416);
nor U18904 (N_18904,N_12344,N_14657);
xor U18905 (N_18905,N_10139,N_13797);
xnor U18906 (N_18906,N_10925,N_10158);
xor U18907 (N_18907,N_13769,N_11634);
nand U18908 (N_18908,N_14098,N_13740);
nor U18909 (N_18909,N_10849,N_11212);
xnor U18910 (N_18910,N_12837,N_13997);
or U18911 (N_18911,N_10876,N_12498);
nor U18912 (N_18912,N_14822,N_12697);
nor U18913 (N_18913,N_14920,N_11078);
or U18914 (N_18914,N_10177,N_12200);
nor U18915 (N_18915,N_12260,N_12504);
nand U18916 (N_18916,N_13590,N_11005);
nor U18917 (N_18917,N_10799,N_13087);
nor U18918 (N_18918,N_12558,N_13368);
or U18919 (N_18919,N_13463,N_13640);
xnor U18920 (N_18920,N_13212,N_10036);
nand U18921 (N_18921,N_10358,N_14934);
nor U18922 (N_18922,N_12328,N_14946);
nand U18923 (N_18923,N_12284,N_11897);
and U18924 (N_18924,N_12050,N_10539);
nand U18925 (N_18925,N_14834,N_14343);
nor U18926 (N_18926,N_11138,N_11855);
nand U18927 (N_18927,N_12216,N_11937);
or U18928 (N_18928,N_12880,N_11343);
and U18929 (N_18929,N_13286,N_13256);
and U18930 (N_18930,N_11602,N_13468);
and U18931 (N_18931,N_12849,N_14051);
or U18932 (N_18932,N_10928,N_12616);
xor U18933 (N_18933,N_12927,N_12610);
or U18934 (N_18934,N_12337,N_14257);
nand U18935 (N_18935,N_13107,N_10524);
or U18936 (N_18936,N_12568,N_11466);
or U18937 (N_18937,N_13080,N_10778);
nand U18938 (N_18938,N_12234,N_13319);
nand U18939 (N_18939,N_14481,N_14784);
xor U18940 (N_18940,N_12651,N_14124);
and U18941 (N_18941,N_14323,N_13909);
nand U18942 (N_18942,N_12955,N_11650);
nand U18943 (N_18943,N_12154,N_14987);
or U18944 (N_18944,N_10744,N_14851);
xnor U18945 (N_18945,N_14193,N_13377);
and U18946 (N_18946,N_10928,N_11383);
xor U18947 (N_18947,N_11457,N_12697);
nor U18948 (N_18948,N_13586,N_13691);
nor U18949 (N_18949,N_14637,N_11714);
nor U18950 (N_18950,N_14864,N_13437);
xnor U18951 (N_18951,N_12196,N_14539);
xor U18952 (N_18952,N_11603,N_14226);
and U18953 (N_18953,N_11899,N_14919);
nor U18954 (N_18954,N_13221,N_13121);
xnor U18955 (N_18955,N_14393,N_13606);
and U18956 (N_18956,N_14904,N_12182);
xor U18957 (N_18957,N_14427,N_14335);
xor U18958 (N_18958,N_12049,N_12172);
and U18959 (N_18959,N_12588,N_13963);
nor U18960 (N_18960,N_13451,N_13035);
nor U18961 (N_18961,N_10513,N_11458);
nor U18962 (N_18962,N_11745,N_13266);
or U18963 (N_18963,N_11658,N_13992);
and U18964 (N_18964,N_10640,N_12629);
xor U18965 (N_18965,N_12895,N_13775);
xnor U18966 (N_18966,N_10975,N_10378);
and U18967 (N_18967,N_11611,N_12617);
or U18968 (N_18968,N_11312,N_13224);
nor U18969 (N_18969,N_11942,N_13624);
nand U18970 (N_18970,N_10165,N_11010);
nand U18971 (N_18971,N_14486,N_13167);
nand U18972 (N_18972,N_13200,N_12836);
and U18973 (N_18973,N_12898,N_12473);
and U18974 (N_18974,N_11336,N_12717);
and U18975 (N_18975,N_10943,N_10415);
or U18976 (N_18976,N_13310,N_10480);
and U18977 (N_18977,N_11695,N_11329);
nor U18978 (N_18978,N_11816,N_12311);
xor U18979 (N_18979,N_14109,N_12257);
nand U18980 (N_18980,N_10590,N_13825);
and U18981 (N_18981,N_14808,N_10912);
nor U18982 (N_18982,N_13914,N_10304);
nand U18983 (N_18983,N_14220,N_10257);
xnor U18984 (N_18984,N_13896,N_10982);
or U18985 (N_18985,N_10474,N_12718);
nand U18986 (N_18986,N_12068,N_12284);
nor U18987 (N_18987,N_13347,N_10239);
nor U18988 (N_18988,N_11820,N_13590);
or U18989 (N_18989,N_11106,N_10978);
and U18990 (N_18990,N_13273,N_13447);
nor U18991 (N_18991,N_12152,N_13213);
nor U18992 (N_18992,N_14678,N_14256);
or U18993 (N_18993,N_14450,N_14514);
nand U18994 (N_18994,N_12392,N_10152);
xor U18995 (N_18995,N_13431,N_11881);
or U18996 (N_18996,N_13806,N_13002);
or U18997 (N_18997,N_11130,N_10654);
or U18998 (N_18998,N_11549,N_12142);
xnor U18999 (N_18999,N_11924,N_10868);
and U19000 (N_19000,N_14026,N_14774);
nand U19001 (N_19001,N_13907,N_13667);
nand U19002 (N_19002,N_10069,N_11967);
nand U19003 (N_19003,N_13066,N_12011);
xor U19004 (N_19004,N_10188,N_10037);
or U19005 (N_19005,N_14711,N_13261);
xnor U19006 (N_19006,N_10450,N_11063);
nor U19007 (N_19007,N_14890,N_12783);
nor U19008 (N_19008,N_12199,N_10918);
nor U19009 (N_19009,N_12727,N_13864);
nor U19010 (N_19010,N_13014,N_12890);
nor U19011 (N_19011,N_13874,N_12889);
xor U19012 (N_19012,N_10842,N_10357);
nand U19013 (N_19013,N_13819,N_10897);
nor U19014 (N_19014,N_13671,N_10924);
nor U19015 (N_19015,N_11016,N_11404);
nand U19016 (N_19016,N_14274,N_13704);
nor U19017 (N_19017,N_12439,N_12732);
xnor U19018 (N_19018,N_11024,N_14830);
nor U19019 (N_19019,N_11011,N_11754);
nand U19020 (N_19020,N_11472,N_14891);
and U19021 (N_19021,N_13735,N_14448);
xor U19022 (N_19022,N_12728,N_13394);
nor U19023 (N_19023,N_12299,N_10897);
and U19024 (N_19024,N_13752,N_11507);
and U19025 (N_19025,N_10419,N_13948);
xor U19026 (N_19026,N_12863,N_11043);
nor U19027 (N_19027,N_12861,N_14353);
and U19028 (N_19028,N_12797,N_10173);
nand U19029 (N_19029,N_11202,N_13399);
and U19030 (N_19030,N_11744,N_10945);
xnor U19031 (N_19031,N_14675,N_11630);
nand U19032 (N_19032,N_13996,N_14518);
and U19033 (N_19033,N_13728,N_10721);
nand U19034 (N_19034,N_12252,N_13856);
nand U19035 (N_19035,N_10307,N_11456);
xor U19036 (N_19036,N_13723,N_10875);
nand U19037 (N_19037,N_10086,N_12885);
or U19038 (N_19038,N_14907,N_11068);
or U19039 (N_19039,N_12470,N_11219);
xnor U19040 (N_19040,N_11520,N_12135);
or U19041 (N_19041,N_11034,N_12441);
and U19042 (N_19042,N_10069,N_10538);
nand U19043 (N_19043,N_10169,N_14121);
nor U19044 (N_19044,N_12855,N_14186);
nor U19045 (N_19045,N_11126,N_14388);
nor U19046 (N_19046,N_10004,N_11489);
and U19047 (N_19047,N_11150,N_10318);
nand U19048 (N_19048,N_10147,N_12701);
nor U19049 (N_19049,N_14139,N_12945);
nor U19050 (N_19050,N_12788,N_13824);
nand U19051 (N_19051,N_13586,N_11529);
or U19052 (N_19052,N_14321,N_14928);
and U19053 (N_19053,N_12530,N_14470);
nand U19054 (N_19054,N_11862,N_10683);
nor U19055 (N_19055,N_12573,N_14204);
and U19056 (N_19056,N_12586,N_12701);
or U19057 (N_19057,N_12527,N_12815);
nand U19058 (N_19058,N_12007,N_12726);
xnor U19059 (N_19059,N_11282,N_13119);
nor U19060 (N_19060,N_11087,N_11186);
or U19061 (N_19061,N_11367,N_13458);
nor U19062 (N_19062,N_11733,N_11853);
nor U19063 (N_19063,N_12393,N_10116);
xor U19064 (N_19064,N_14978,N_13603);
xnor U19065 (N_19065,N_10643,N_11965);
or U19066 (N_19066,N_12709,N_10696);
nand U19067 (N_19067,N_13749,N_12844);
nand U19068 (N_19068,N_10684,N_13876);
nor U19069 (N_19069,N_10189,N_13579);
xor U19070 (N_19070,N_12412,N_14519);
nor U19071 (N_19071,N_10068,N_13320);
xor U19072 (N_19072,N_10401,N_11397);
and U19073 (N_19073,N_14847,N_10976);
nand U19074 (N_19074,N_12907,N_12390);
nand U19075 (N_19075,N_14700,N_10995);
nor U19076 (N_19076,N_12998,N_11144);
nand U19077 (N_19077,N_13228,N_10434);
nor U19078 (N_19078,N_13938,N_10874);
nand U19079 (N_19079,N_11005,N_11810);
nand U19080 (N_19080,N_13875,N_10109);
and U19081 (N_19081,N_13016,N_13084);
nor U19082 (N_19082,N_14449,N_11169);
xnor U19083 (N_19083,N_11205,N_11322);
nand U19084 (N_19084,N_10686,N_13138);
and U19085 (N_19085,N_14852,N_11016);
or U19086 (N_19086,N_11077,N_10122);
or U19087 (N_19087,N_12685,N_13410);
xor U19088 (N_19088,N_12547,N_14012);
and U19089 (N_19089,N_14821,N_12178);
nor U19090 (N_19090,N_10313,N_11985);
and U19091 (N_19091,N_12197,N_11288);
xor U19092 (N_19092,N_10691,N_13920);
nand U19093 (N_19093,N_10508,N_14479);
and U19094 (N_19094,N_10354,N_10934);
nand U19095 (N_19095,N_14921,N_13176);
or U19096 (N_19096,N_10893,N_12536);
xor U19097 (N_19097,N_14105,N_13358);
or U19098 (N_19098,N_14250,N_13599);
nand U19099 (N_19099,N_11415,N_12038);
and U19100 (N_19100,N_10523,N_12817);
nand U19101 (N_19101,N_12313,N_11551);
or U19102 (N_19102,N_14379,N_14766);
nor U19103 (N_19103,N_14123,N_12243);
nand U19104 (N_19104,N_12585,N_13380);
xor U19105 (N_19105,N_12133,N_10156);
nor U19106 (N_19106,N_14682,N_14989);
xor U19107 (N_19107,N_13057,N_10467);
nor U19108 (N_19108,N_13756,N_14431);
and U19109 (N_19109,N_12468,N_11239);
or U19110 (N_19110,N_10427,N_14396);
nand U19111 (N_19111,N_10849,N_14735);
or U19112 (N_19112,N_14276,N_12539);
nor U19113 (N_19113,N_13773,N_13272);
xnor U19114 (N_19114,N_13692,N_12065);
and U19115 (N_19115,N_12042,N_10984);
and U19116 (N_19116,N_14415,N_13433);
nand U19117 (N_19117,N_10726,N_13749);
and U19118 (N_19118,N_10598,N_11314);
xor U19119 (N_19119,N_14077,N_13099);
nor U19120 (N_19120,N_10392,N_12490);
nor U19121 (N_19121,N_13462,N_12486);
and U19122 (N_19122,N_12096,N_11737);
nand U19123 (N_19123,N_11154,N_11853);
or U19124 (N_19124,N_12271,N_11180);
xor U19125 (N_19125,N_11012,N_10814);
xor U19126 (N_19126,N_10379,N_11954);
or U19127 (N_19127,N_11821,N_12000);
nand U19128 (N_19128,N_10391,N_10863);
xor U19129 (N_19129,N_13112,N_11258);
xnor U19130 (N_19130,N_12868,N_11762);
nor U19131 (N_19131,N_11387,N_12564);
nand U19132 (N_19132,N_12862,N_12431);
xor U19133 (N_19133,N_10475,N_14956);
or U19134 (N_19134,N_10288,N_12203);
or U19135 (N_19135,N_12699,N_11394);
or U19136 (N_19136,N_13460,N_11939);
xor U19137 (N_19137,N_14619,N_14688);
nor U19138 (N_19138,N_13587,N_13008);
and U19139 (N_19139,N_10193,N_13322);
xnor U19140 (N_19140,N_10772,N_14758);
xor U19141 (N_19141,N_11745,N_10127);
and U19142 (N_19142,N_14185,N_13256);
nand U19143 (N_19143,N_12160,N_14700);
and U19144 (N_19144,N_13262,N_10949);
xor U19145 (N_19145,N_10515,N_13751);
nor U19146 (N_19146,N_10173,N_14426);
or U19147 (N_19147,N_13337,N_10706);
xor U19148 (N_19148,N_11266,N_10844);
nor U19149 (N_19149,N_12436,N_12138);
nand U19150 (N_19150,N_13300,N_14428);
or U19151 (N_19151,N_12799,N_10121);
xnor U19152 (N_19152,N_12064,N_10617);
nand U19153 (N_19153,N_11976,N_13872);
nand U19154 (N_19154,N_12692,N_11655);
and U19155 (N_19155,N_10982,N_12712);
and U19156 (N_19156,N_11465,N_13625);
and U19157 (N_19157,N_10775,N_13113);
xnor U19158 (N_19158,N_11856,N_14842);
or U19159 (N_19159,N_10577,N_10849);
or U19160 (N_19160,N_13003,N_14091);
nand U19161 (N_19161,N_12707,N_10384);
nor U19162 (N_19162,N_11341,N_10970);
nor U19163 (N_19163,N_12694,N_13352);
xnor U19164 (N_19164,N_12286,N_13190);
nor U19165 (N_19165,N_12712,N_11259);
nor U19166 (N_19166,N_11571,N_11787);
or U19167 (N_19167,N_13657,N_10519);
nor U19168 (N_19168,N_11781,N_10619);
nand U19169 (N_19169,N_11185,N_11440);
and U19170 (N_19170,N_14737,N_13753);
nand U19171 (N_19171,N_10282,N_11549);
nor U19172 (N_19172,N_10791,N_13738);
nand U19173 (N_19173,N_14553,N_13468);
nand U19174 (N_19174,N_13740,N_14639);
xor U19175 (N_19175,N_10612,N_11429);
or U19176 (N_19176,N_13408,N_12261);
xnor U19177 (N_19177,N_14174,N_10672);
nor U19178 (N_19178,N_14315,N_14977);
and U19179 (N_19179,N_11566,N_13726);
and U19180 (N_19180,N_12265,N_11447);
nand U19181 (N_19181,N_12809,N_14009);
or U19182 (N_19182,N_10740,N_14463);
or U19183 (N_19183,N_12379,N_11649);
nand U19184 (N_19184,N_10352,N_11956);
nand U19185 (N_19185,N_12842,N_13684);
nand U19186 (N_19186,N_14411,N_12017);
nor U19187 (N_19187,N_12537,N_14127);
and U19188 (N_19188,N_12074,N_12270);
nand U19189 (N_19189,N_10076,N_12911);
or U19190 (N_19190,N_14806,N_10611);
nor U19191 (N_19191,N_10854,N_11052);
or U19192 (N_19192,N_11442,N_14069);
nand U19193 (N_19193,N_14865,N_11231);
xnor U19194 (N_19194,N_14829,N_10219);
xor U19195 (N_19195,N_14548,N_12330);
xnor U19196 (N_19196,N_12443,N_10338);
xor U19197 (N_19197,N_13787,N_10855);
nand U19198 (N_19198,N_10247,N_10628);
nand U19199 (N_19199,N_11040,N_11453);
nand U19200 (N_19200,N_13445,N_13201);
nor U19201 (N_19201,N_13253,N_11259);
xnor U19202 (N_19202,N_13571,N_10517);
nand U19203 (N_19203,N_13955,N_14349);
nor U19204 (N_19204,N_12794,N_11778);
nand U19205 (N_19205,N_11512,N_13720);
nand U19206 (N_19206,N_14428,N_10950);
and U19207 (N_19207,N_13279,N_14039);
nand U19208 (N_19208,N_13373,N_10932);
xnor U19209 (N_19209,N_10788,N_11361);
nor U19210 (N_19210,N_13547,N_14991);
and U19211 (N_19211,N_11847,N_12371);
nor U19212 (N_19212,N_10200,N_10219);
xnor U19213 (N_19213,N_11748,N_13752);
and U19214 (N_19214,N_12250,N_10755);
nand U19215 (N_19215,N_14609,N_13051);
and U19216 (N_19216,N_14778,N_13111);
and U19217 (N_19217,N_12748,N_10960);
nand U19218 (N_19218,N_11264,N_10697);
or U19219 (N_19219,N_10365,N_14662);
nand U19220 (N_19220,N_14885,N_11146);
xor U19221 (N_19221,N_10219,N_13263);
or U19222 (N_19222,N_11060,N_13591);
nand U19223 (N_19223,N_11756,N_11331);
nand U19224 (N_19224,N_11030,N_10973);
nor U19225 (N_19225,N_13226,N_11225);
or U19226 (N_19226,N_10143,N_11065);
xnor U19227 (N_19227,N_12546,N_13015);
xnor U19228 (N_19228,N_10014,N_14843);
or U19229 (N_19229,N_13244,N_12186);
nand U19230 (N_19230,N_10364,N_10049);
nor U19231 (N_19231,N_13740,N_10587);
nand U19232 (N_19232,N_14723,N_13867);
or U19233 (N_19233,N_10061,N_12171);
nand U19234 (N_19234,N_11936,N_10646);
xor U19235 (N_19235,N_10378,N_14917);
nand U19236 (N_19236,N_14986,N_11732);
nand U19237 (N_19237,N_14818,N_12816);
nor U19238 (N_19238,N_12537,N_12501);
or U19239 (N_19239,N_12453,N_12783);
xnor U19240 (N_19240,N_10727,N_12315);
xnor U19241 (N_19241,N_11216,N_11427);
and U19242 (N_19242,N_10702,N_12373);
nor U19243 (N_19243,N_12172,N_14926);
xnor U19244 (N_19244,N_11136,N_11968);
or U19245 (N_19245,N_14309,N_10899);
xor U19246 (N_19246,N_13028,N_13429);
and U19247 (N_19247,N_14391,N_13524);
and U19248 (N_19248,N_11589,N_11559);
and U19249 (N_19249,N_14368,N_12185);
nand U19250 (N_19250,N_10436,N_14279);
nor U19251 (N_19251,N_14086,N_10475);
nor U19252 (N_19252,N_14518,N_12387);
nor U19253 (N_19253,N_13271,N_11260);
nor U19254 (N_19254,N_11609,N_13637);
nand U19255 (N_19255,N_13265,N_11044);
or U19256 (N_19256,N_14872,N_10495);
xnor U19257 (N_19257,N_13013,N_12377);
nor U19258 (N_19258,N_14264,N_12952);
or U19259 (N_19259,N_13193,N_13113);
or U19260 (N_19260,N_10281,N_13514);
nor U19261 (N_19261,N_14625,N_13267);
nor U19262 (N_19262,N_11996,N_14402);
nor U19263 (N_19263,N_12611,N_12722);
and U19264 (N_19264,N_13677,N_11377);
xor U19265 (N_19265,N_10929,N_13906);
or U19266 (N_19266,N_14444,N_10948);
nand U19267 (N_19267,N_11088,N_13428);
or U19268 (N_19268,N_14363,N_14400);
and U19269 (N_19269,N_12597,N_13191);
and U19270 (N_19270,N_14449,N_11314);
nand U19271 (N_19271,N_10498,N_13340);
nor U19272 (N_19272,N_14831,N_14552);
and U19273 (N_19273,N_14269,N_14840);
nand U19274 (N_19274,N_14378,N_12336);
nand U19275 (N_19275,N_11385,N_10935);
and U19276 (N_19276,N_12232,N_11649);
nor U19277 (N_19277,N_12038,N_13618);
and U19278 (N_19278,N_11740,N_13199);
and U19279 (N_19279,N_10255,N_13580);
nand U19280 (N_19280,N_10025,N_12377);
nand U19281 (N_19281,N_13875,N_12379);
nor U19282 (N_19282,N_10528,N_14806);
and U19283 (N_19283,N_11607,N_10032);
nand U19284 (N_19284,N_12926,N_11370);
nand U19285 (N_19285,N_12504,N_12889);
nand U19286 (N_19286,N_13190,N_11830);
nor U19287 (N_19287,N_11915,N_10660);
nor U19288 (N_19288,N_14212,N_10126);
nor U19289 (N_19289,N_13736,N_11363);
nand U19290 (N_19290,N_14818,N_12787);
nand U19291 (N_19291,N_13077,N_14291);
nor U19292 (N_19292,N_14523,N_13133);
xor U19293 (N_19293,N_12055,N_11957);
and U19294 (N_19294,N_13954,N_14271);
nand U19295 (N_19295,N_14120,N_13501);
and U19296 (N_19296,N_11516,N_10320);
and U19297 (N_19297,N_11046,N_11589);
xor U19298 (N_19298,N_12321,N_14617);
xnor U19299 (N_19299,N_11566,N_10581);
xnor U19300 (N_19300,N_14719,N_14004);
or U19301 (N_19301,N_13915,N_11158);
or U19302 (N_19302,N_11286,N_12897);
xor U19303 (N_19303,N_10425,N_12227);
nand U19304 (N_19304,N_13401,N_10002);
nor U19305 (N_19305,N_12788,N_11469);
or U19306 (N_19306,N_11172,N_11472);
nor U19307 (N_19307,N_11548,N_12367);
xor U19308 (N_19308,N_14049,N_14082);
xnor U19309 (N_19309,N_13125,N_11057);
nor U19310 (N_19310,N_13890,N_11811);
or U19311 (N_19311,N_12036,N_10896);
xnor U19312 (N_19312,N_10137,N_10594);
xnor U19313 (N_19313,N_10740,N_12903);
nor U19314 (N_19314,N_11548,N_10973);
xor U19315 (N_19315,N_13341,N_13781);
or U19316 (N_19316,N_11986,N_13744);
and U19317 (N_19317,N_11861,N_10049);
nor U19318 (N_19318,N_14104,N_14747);
or U19319 (N_19319,N_14018,N_14645);
nand U19320 (N_19320,N_10186,N_14862);
nand U19321 (N_19321,N_11285,N_11415);
nor U19322 (N_19322,N_10290,N_10521);
nand U19323 (N_19323,N_10660,N_12754);
nor U19324 (N_19324,N_14817,N_11776);
and U19325 (N_19325,N_14719,N_10074);
or U19326 (N_19326,N_10630,N_13410);
nor U19327 (N_19327,N_12119,N_14728);
nand U19328 (N_19328,N_10718,N_14893);
nor U19329 (N_19329,N_12329,N_12178);
nor U19330 (N_19330,N_11373,N_14033);
or U19331 (N_19331,N_11983,N_14596);
nand U19332 (N_19332,N_10442,N_10233);
nor U19333 (N_19333,N_11801,N_13602);
or U19334 (N_19334,N_14089,N_11334);
and U19335 (N_19335,N_12925,N_14650);
nor U19336 (N_19336,N_13402,N_12358);
nor U19337 (N_19337,N_13907,N_13487);
or U19338 (N_19338,N_11156,N_12568);
xnor U19339 (N_19339,N_14114,N_11619);
nor U19340 (N_19340,N_10440,N_11829);
and U19341 (N_19341,N_11611,N_10312);
or U19342 (N_19342,N_14419,N_10129);
or U19343 (N_19343,N_13005,N_13701);
or U19344 (N_19344,N_12483,N_13707);
or U19345 (N_19345,N_10389,N_14862);
and U19346 (N_19346,N_12457,N_13232);
or U19347 (N_19347,N_14067,N_14759);
nor U19348 (N_19348,N_13346,N_12898);
or U19349 (N_19349,N_12161,N_11979);
or U19350 (N_19350,N_13756,N_13600);
xnor U19351 (N_19351,N_10039,N_13368);
or U19352 (N_19352,N_14910,N_13524);
and U19353 (N_19353,N_10401,N_13631);
nor U19354 (N_19354,N_10228,N_13526);
and U19355 (N_19355,N_10805,N_11211);
nand U19356 (N_19356,N_13349,N_14589);
or U19357 (N_19357,N_14809,N_13871);
or U19358 (N_19358,N_12312,N_13143);
or U19359 (N_19359,N_13099,N_14182);
xnor U19360 (N_19360,N_10597,N_13598);
and U19361 (N_19361,N_10237,N_11569);
nor U19362 (N_19362,N_13853,N_10309);
nand U19363 (N_19363,N_10053,N_13126);
nand U19364 (N_19364,N_11996,N_13687);
xor U19365 (N_19365,N_13768,N_13172);
nor U19366 (N_19366,N_10262,N_10312);
nand U19367 (N_19367,N_10836,N_11975);
nand U19368 (N_19368,N_14895,N_11007);
xor U19369 (N_19369,N_12671,N_10291);
nor U19370 (N_19370,N_10317,N_13000);
or U19371 (N_19371,N_14303,N_12662);
and U19372 (N_19372,N_11454,N_12948);
nand U19373 (N_19373,N_13801,N_12965);
and U19374 (N_19374,N_13982,N_13275);
nand U19375 (N_19375,N_14044,N_12794);
or U19376 (N_19376,N_12413,N_14380);
and U19377 (N_19377,N_12328,N_12771);
xnor U19378 (N_19378,N_11359,N_10513);
and U19379 (N_19379,N_13869,N_13337);
nor U19380 (N_19380,N_12438,N_12720);
nand U19381 (N_19381,N_13910,N_12064);
or U19382 (N_19382,N_13750,N_13124);
xor U19383 (N_19383,N_14907,N_13604);
or U19384 (N_19384,N_11882,N_12856);
and U19385 (N_19385,N_13149,N_11895);
nor U19386 (N_19386,N_13999,N_11209);
xor U19387 (N_19387,N_14003,N_13269);
nand U19388 (N_19388,N_10038,N_10350);
xnor U19389 (N_19389,N_11465,N_13309);
xnor U19390 (N_19390,N_12652,N_14174);
and U19391 (N_19391,N_11191,N_14001);
nor U19392 (N_19392,N_12819,N_10638);
nand U19393 (N_19393,N_10853,N_12715);
nor U19394 (N_19394,N_11468,N_11311);
or U19395 (N_19395,N_10202,N_13545);
and U19396 (N_19396,N_11535,N_14755);
nor U19397 (N_19397,N_10555,N_14521);
nor U19398 (N_19398,N_13686,N_11460);
xnor U19399 (N_19399,N_12634,N_10142);
and U19400 (N_19400,N_12625,N_10890);
and U19401 (N_19401,N_13854,N_14806);
nand U19402 (N_19402,N_11007,N_10178);
nor U19403 (N_19403,N_11957,N_11036);
and U19404 (N_19404,N_12624,N_13730);
or U19405 (N_19405,N_13255,N_11479);
and U19406 (N_19406,N_12353,N_14568);
nand U19407 (N_19407,N_14082,N_12020);
nand U19408 (N_19408,N_14052,N_11933);
and U19409 (N_19409,N_14271,N_11342);
or U19410 (N_19410,N_11165,N_10666);
nor U19411 (N_19411,N_10536,N_13728);
and U19412 (N_19412,N_10920,N_14795);
and U19413 (N_19413,N_10961,N_13715);
xnor U19414 (N_19414,N_10221,N_10607);
nand U19415 (N_19415,N_10018,N_12802);
xnor U19416 (N_19416,N_11287,N_13896);
or U19417 (N_19417,N_13817,N_10261);
nor U19418 (N_19418,N_14648,N_14986);
and U19419 (N_19419,N_11929,N_13822);
or U19420 (N_19420,N_11747,N_10656);
xnor U19421 (N_19421,N_13581,N_12947);
xnor U19422 (N_19422,N_13411,N_11789);
or U19423 (N_19423,N_12346,N_14757);
nor U19424 (N_19424,N_11462,N_12702);
nor U19425 (N_19425,N_11778,N_13733);
xnor U19426 (N_19426,N_10968,N_10343);
and U19427 (N_19427,N_11383,N_11045);
or U19428 (N_19428,N_10054,N_12988);
xor U19429 (N_19429,N_11951,N_12757);
nand U19430 (N_19430,N_11657,N_11072);
and U19431 (N_19431,N_13521,N_13484);
or U19432 (N_19432,N_14714,N_13837);
xnor U19433 (N_19433,N_14956,N_13681);
nor U19434 (N_19434,N_13009,N_10259);
and U19435 (N_19435,N_14584,N_11295);
or U19436 (N_19436,N_11559,N_12237);
xnor U19437 (N_19437,N_12944,N_10285);
and U19438 (N_19438,N_12441,N_13627);
nand U19439 (N_19439,N_11357,N_11171);
and U19440 (N_19440,N_11932,N_12037);
or U19441 (N_19441,N_11982,N_14227);
nor U19442 (N_19442,N_13202,N_12321);
nand U19443 (N_19443,N_13084,N_10618);
and U19444 (N_19444,N_11823,N_14232);
nor U19445 (N_19445,N_12612,N_12888);
and U19446 (N_19446,N_12292,N_10096);
nor U19447 (N_19447,N_11696,N_11020);
nand U19448 (N_19448,N_11425,N_10185);
nor U19449 (N_19449,N_13065,N_11411);
and U19450 (N_19450,N_14013,N_13213);
nor U19451 (N_19451,N_10540,N_11499);
nand U19452 (N_19452,N_10201,N_11725);
or U19453 (N_19453,N_13924,N_11265);
nand U19454 (N_19454,N_14608,N_12129);
nand U19455 (N_19455,N_10921,N_14617);
or U19456 (N_19456,N_10783,N_11028);
xor U19457 (N_19457,N_11057,N_11403);
xnor U19458 (N_19458,N_14870,N_14537);
and U19459 (N_19459,N_14351,N_10226);
and U19460 (N_19460,N_10712,N_11802);
nand U19461 (N_19461,N_13320,N_12766);
nand U19462 (N_19462,N_10852,N_10057);
nor U19463 (N_19463,N_13323,N_13200);
or U19464 (N_19464,N_14080,N_13393);
and U19465 (N_19465,N_10887,N_12066);
or U19466 (N_19466,N_14912,N_13480);
nor U19467 (N_19467,N_11193,N_10131);
or U19468 (N_19468,N_13608,N_10930);
and U19469 (N_19469,N_12182,N_11477);
and U19470 (N_19470,N_11054,N_12662);
xor U19471 (N_19471,N_12753,N_13213);
xnor U19472 (N_19472,N_12391,N_13610);
and U19473 (N_19473,N_13192,N_11328);
nand U19474 (N_19474,N_12010,N_14843);
and U19475 (N_19475,N_12545,N_11865);
nor U19476 (N_19476,N_11081,N_11881);
nor U19477 (N_19477,N_12346,N_11419);
and U19478 (N_19478,N_14045,N_10366);
xnor U19479 (N_19479,N_14493,N_13346);
nor U19480 (N_19480,N_11057,N_14278);
xnor U19481 (N_19481,N_12120,N_12913);
nor U19482 (N_19482,N_14256,N_13178);
nand U19483 (N_19483,N_11708,N_10411);
xor U19484 (N_19484,N_12385,N_12616);
nand U19485 (N_19485,N_10260,N_13788);
or U19486 (N_19486,N_11562,N_12455);
and U19487 (N_19487,N_11543,N_12209);
nand U19488 (N_19488,N_11872,N_10007);
or U19489 (N_19489,N_14491,N_11879);
and U19490 (N_19490,N_13948,N_13613);
nand U19491 (N_19491,N_14914,N_10909);
or U19492 (N_19492,N_10501,N_14570);
xor U19493 (N_19493,N_12904,N_12695);
nand U19494 (N_19494,N_12596,N_14833);
nor U19495 (N_19495,N_13814,N_11510);
and U19496 (N_19496,N_11969,N_13335);
nand U19497 (N_19497,N_10552,N_13815);
or U19498 (N_19498,N_12739,N_12394);
or U19499 (N_19499,N_14921,N_11446);
nor U19500 (N_19500,N_11767,N_11759);
nand U19501 (N_19501,N_13056,N_13880);
xnor U19502 (N_19502,N_14457,N_13171);
xnor U19503 (N_19503,N_11754,N_11381);
and U19504 (N_19504,N_13282,N_12790);
nand U19505 (N_19505,N_13049,N_10168);
nor U19506 (N_19506,N_11249,N_10885);
xor U19507 (N_19507,N_14960,N_11328);
and U19508 (N_19508,N_13882,N_12448);
and U19509 (N_19509,N_11620,N_10762);
and U19510 (N_19510,N_10905,N_11554);
nor U19511 (N_19511,N_13932,N_11602);
nor U19512 (N_19512,N_10120,N_12950);
xor U19513 (N_19513,N_12203,N_12814);
or U19514 (N_19514,N_12413,N_10656);
xnor U19515 (N_19515,N_13647,N_13093);
or U19516 (N_19516,N_13792,N_13736);
xor U19517 (N_19517,N_11571,N_10345);
xor U19518 (N_19518,N_14329,N_10779);
and U19519 (N_19519,N_13339,N_10749);
nand U19520 (N_19520,N_12423,N_12134);
and U19521 (N_19521,N_12814,N_12986);
nor U19522 (N_19522,N_14894,N_13509);
nor U19523 (N_19523,N_10907,N_13389);
xor U19524 (N_19524,N_14145,N_12398);
nand U19525 (N_19525,N_11684,N_10456);
and U19526 (N_19526,N_10842,N_12935);
xnor U19527 (N_19527,N_11447,N_14450);
and U19528 (N_19528,N_14598,N_11649);
nand U19529 (N_19529,N_13928,N_12098);
and U19530 (N_19530,N_14471,N_13292);
or U19531 (N_19531,N_12112,N_13835);
xnor U19532 (N_19532,N_12650,N_11408);
nand U19533 (N_19533,N_14352,N_11371);
nand U19534 (N_19534,N_13270,N_14586);
or U19535 (N_19535,N_12022,N_14106);
nand U19536 (N_19536,N_10516,N_14102);
nor U19537 (N_19537,N_13981,N_12922);
nor U19538 (N_19538,N_13777,N_10989);
and U19539 (N_19539,N_13660,N_11150);
nand U19540 (N_19540,N_12076,N_12970);
nand U19541 (N_19541,N_12906,N_13679);
xor U19542 (N_19542,N_10181,N_13825);
nor U19543 (N_19543,N_13797,N_12219);
or U19544 (N_19544,N_12809,N_11444);
xor U19545 (N_19545,N_14365,N_14890);
nor U19546 (N_19546,N_10256,N_10784);
xnor U19547 (N_19547,N_13699,N_12662);
nor U19548 (N_19548,N_12735,N_13052);
nand U19549 (N_19549,N_12437,N_12939);
nand U19550 (N_19550,N_13414,N_13943);
or U19551 (N_19551,N_13513,N_14089);
or U19552 (N_19552,N_13061,N_11126);
nor U19553 (N_19553,N_14872,N_13915);
and U19554 (N_19554,N_12718,N_10682);
nor U19555 (N_19555,N_13131,N_13486);
or U19556 (N_19556,N_14297,N_14238);
and U19557 (N_19557,N_11687,N_11906);
xor U19558 (N_19558,N_14701,N_11847);
or U19559 (N_19559,N_13367,N_14609);
xnor U19560 (N_19560,N_11296,N_13978);
nand U19561 (N_19561,N_12048,N_13845);
nand U19562 (N_19562,N_12713,N_12636);
nor U19563 (N_19563,N_12863,N_13260);
xor U19564 (N_19564,N_14533,N_10095);
nand U19565 (N_19565,N_10308,N_14501);
nand U19566 (N_19566,N_10578,N_12143);
xnor U19567 (N_19567,N_11339,N_12700);
xnor U19568 (N_19568,N_10753,N_13018);
nor U19569 (N_19569,N_11852,N_10762);
nor U19570 (N_19570,N_13018,N_14871);
nand U19571 (N_19571,N_13059,N_10692);
and U19572 (N_19572,N_12378,N_12767);
nand U19573 (N_19573,N_14241,N_11114);
nor U19574 (N_19574,N_13464,N_11197);
or U19575 (N_19575,N_11020,N_13804);
or U19576 (N_19576,N_13592,N_10122);
and U19577 (N_19577,N_10160,N_12488);
xnor U19578 (N_19578,N_12002,N_13635);
xnor U19579 (N_19579,N_12869,N_11135);
or U19580 (N_19580,N_13467,N_10414);
xnor U19581 (N_19581,N_12734,N_10404);
and U19582 (N_19582,N_13018,N_12773);
xnor U19583 (N_19583,N_11788,N_14113);
nand U19584 (N_19584,N_12886,N_11365);
and U19585 (N_19585,N_14201,N_11943);
xor U19586 (N_19586,N_13211,N_14183);
xor U19587 (N_19587,N_11763,N_14840);
or U19588 (N_19588,N_10722,N_10505);
nand U19589 (N_19589,N_12342,N_10821);
nor U19590 (N_19590,N_12578,N_14526);
or U19591 (N_19591,N_14894,N_14224);
nand U19592 (N_19592,N_12996,N_10733);
nand U19593 (N_19593,N_13266,N_10570);
nand U19594 (N_19594,N_13353,N_10142);
and U19595 (N_19595,N_14412,N_13318);
nor U19596 (N_19596,N_13692,N_12347);
nor U19597 (N_19597,N_10072,N_11034);
nand U19598 (N_19598,N_13568,N_12939);
and U19599 (N_19599,N_14642,N_12995);
xnor U19600 (N_19600,N_13089,N_14356);
nor U19601 (N_19601,N_10922,N_10200);
nor U19602 (N_19602,N_10991,N_11135);
nor U19603 (N_19603,N_13735,N_11820);
xnor U19604 (N_19604,N_13226,N_11601);
nand U19605 (N_19605,N_10923,N_11079);
nor U19606 (N_19606,N_13217,N_14026);
and U19607 (N_19607,N_11687,N_14712);
xor U19608 (N_19608,N_13766,N_12211);
nor U19609 (N_19609,N_13009,N_11830);
xor U19610 (N_19610,N_14225,N_14471);
or U19611 (N_19611,N_14387,N_14657);
nor U19612 (N_19612,N_13164,N_13707);
and U19613 (N_19613,N_14231,N_10766);
nor U19614 (N_19614,N_12772,N_12670);
and U19615 (N_19615,N_11051,N_13470);
and U19616 (N_19616,N_13592,N_12084);
or U19617 (N_19617,N_13979,N_10355);
xor U19618 (N_19618,N_10141,N_13569);
nor U19619 (N_19619,N_12626,N_11675);
nand U19620 (N_19620,N_12467,N_12240);
nand U19621 (N_19621,N_11860,N_14249);
xnor U19622 (N_19622,N_10076,N_10614);
nor U19623 (N_19623,N_12722,N_13341);
or U19624 (N_19624,N_13188,N_12235);
nand U19625 (N_19625,N_13282,N_12852);
nor U19626 (N_19626,N_12857,N_10883);
or U19627 (N_19627,N_13256,N_14384);
or U19628 (N_19628,N_12623,N_14585);
nor U19629 (N_19629,N_10859,N_10308);
nand U19630 (N_19630,N_13825,N_12117);
xor U19631 (N_19631,N_10068,N_10077);
xnor U19632 (N_19632,N_14358,N_11047);
nand U19633 (N_19633,N_11776,N_14800);
and U19634 (N_19634,N_12023,N_13464);
nor U19635 (N_19635,N_11703,N_11473);
or U19636 (N_19636,N_11971,N_14829);
or U19637 (N_19637,N_13033,N_10846);
or U19638 (N_19638,N_14098,N_10062);
nor U19639 (N_19639,N_13468,N_12477);
or U19640 (N_19640,N_13781,N_10859);
or U19641 (N_19641,N_14529,N_10568);
and U19642 (N_19642,N_11122,N_13465);
xor U19643 (N_19643,N_12221,N_13835);
nor U19644 (N_19644,N_11832,N_11384);
nor U19645 (N_19645,N_12402,N_14900);
nor U19646 (N_19646,N_13892,N_10962);
nand U19647 (N_19647,N_14204,N_12322);
or U19648 (N_19648,N_13324,N_11501);
nand U19649 (N_19649,N_12181,N_10781);
nor U19650 (N_19650,N_11217,N_12199);
nor U19651 (N_19651,N_11127,N_14681);
xnor U19652 (N_19652,N_14977,N_12695);
nor U19653 (N_19653,N_10208,N_13003);
nor U19654 (N_19654,N_10743,N_12652);
and U19655 (N_19655,N_14011,N_10146);
and U19656 (N_19656,N_12160,N_12702);
or U19657 (N_19657,N_12782,N_13030);
and U19658 (N_19658,N_13243,N_12501);
xor U19659 (N_19659,N_11528,N_10336);
nand U19660 (N_19660,N_10060,N_14312);
nor U19661 (N_19661,N_14356,N_14311);
and U19662 (N_19662,N_13979,N_11765);
xor U19663 (N_19663,N_13492,N_13223);
and U19664 (N_19664,N_11224,N_13563);
xor U19665 (N_19665,N_13563,N_13382);
nor U19666 (N_19666,N_10119,N_14759);
and U19667 (N_19667,N_10363,N_10665);
or U19668 (N_19668,N_12639,N_12157);
xor U19669 (N_19669,N_13901,N_12864);
nand U19670 (N_19670,N_13521,N_14952);
nand U19671 (N_19671,N_12481,N_12739);
or U19672 (N_19672,N_13982,N_11877);
or U19673 (N_19673,N_10921,N_11998);
nand U19674 (N_19674,N_13699,N_10218);
nand U19675 (N_19675,N_11438,N_10816);
or U19676 (N_19676,N_11643,N_14771);
and U19677 (N_19677,N_12250,N_10908);
xnor U19678 (N_19678,N_11677,N_12389);
xor U19679 (N_19679,N_11369,N_11767);
and U19680 (N_19680,N_12555,N_14515);
nor U19681 (N_19681,N_14772,N_11989);
and U19682 (N_19682,N_13681,N_11810);
and U19683 (N_19683,N_12290,N_14938);
nand U19684 (N_19684,N_10995,N_14752);
and U19685 (N_19685,N_10343,N_11443);
and U19686 (N_19686,N_11344,N_11230);
and U19687 (N_19687,N_13343,N_12609);
or U19688 (N_19688,N_13076,N_10539);
xor U19689 (N_19689,N_10258,N_12892);
or U19690 (N_19690,N_14879,N_12785);
nor U19691 (N_19691,N_10475,N_12877);
or U19692 (N_19692,N_12729,N_13648);
xor U19693 (N_19693,N_12935,N_12404);
nand U19694 (N_19694,N_13543,N_14197);
or U19695 (N_19695,N_12007,N_13595);
and U19696 (N_19696,N_13190,N_10794);
nand U19697 (N_19697,N_13060,N_12885);
or U19698 (N_19698,N_13593,N_11577);
nand U19699 (N_19699,N_12622,N_13733);
nand U19700 (N_19700,N_13726,N_11845);
nand U19701 (N_19701,N_11101,N_14791);
and U19702 (N_19702,N_14675,N_14811);
xnor U19703 (N_19703,N_14605,N_13387);
xor U19704 (N_19704,N_13511,N_12124);
and U19705 (N_19705,N_13459,N_12612);
and U19706 (N_19706,N_13819,N_10314);
or U19707 (N_19707,N_12531,N_11821);
xnor U19708 (N_19708,N_14287,N_13768);
xor U19709 (N_19709,N_13385,N_12089);
and U19710 (N_19710,N_13914,N_13862);
or U19711 (N_19711,N_11402,N_14730);
nor U19712 (N_19712,N_13968,N_13309);
xnor U19713 (N_19713,N_10392,N_11438);
or U19714 (N_19714,N_13058,N_12381);
nand U19715 (N_19715,N_10313,N_12883);
or U19716 (N_19716,N_13487,N_14502);
nand U19717 (N_19717,N_10423,N_13345);
nand U19718 (N_19718,N_10536,N_12501);
nor U19719 (N_19719,N_14150,N_14644);
nand U19720 (N_19720,N_13835,N_14933);
nor U19721 (N_19721,N_10095,N_12829);
or U19722 (N_19722,N_14667,N_13231);
nor U19723 (N_19723,N_12139,N_10331);
nand U19724 (N_19724,N_13267,N_13409);
nor U19725 (N_19725,N_14108,N_14225);
nand U19726 (N_19726,N_10841,N_14861);
nor U19727 (N_19727,N_14242,N_12027);
or U19728 (N_19728,N_14589,N_11705);
nor U19729 (N_19729,N_10659,N_12349);
and U19730 (N_19730,N_10587,N_10787);
or U19731 (N_19731,N_10609,N_10209);
or U19732 (N_19732,N_13961,N_12605);
xnor U19733 (N_19733,N_14260,N_12705);
or U19734 (N_19734,N_13210,N_12334);
nor U19735 (N_19735,N_13180,N_14143);
or U19736 (N_19736,N_12628,N_13892);
xor U19737 (N_19737,N_14425,N_13621);
xor U19738 (N_19738,N_13862,N_10666);
nand U19739 (N_19739,N_10565,N_13519);
or U19740 (N_19740,N_14894,N_12253);
xor U19741 (N_19741,N_14642,N_11914);
nor U19742 (N_19742,N_13678,N_12576);
nand U19743 (N_19743,N_13200,N_12495);
nor U19744 (N_19744,N_13030,N_13059);
xor U19745 (N_19745,N_10649,N_10813);
nand U19746 (N_19746,N_14601,N_13300);
nor U19747 (N_19747,N_11961,N_14673);
or U19748 (N_19748,N_10350,N_12134);
and U19749 (N_19749,N_11470,N_13698);
and U19750 (N_19750,N_12646,N_10968);
or U19751 (N_19751,N_13663,N_11672);
nor U19752 (N_19752,N_12590,N_10054);
and U19753 (N_19753,N_13080,N_10366);
or U19754 (N_19754,N_12846,N_11174);
or U19755 (N_19755,N_11808,N_10793);
xnor U19756 (N_19756,N_13470,N_11020);
or U19757 (N_19757,N_12651,N_13940);
nand U19758 (N_19758,N_13108,N_14915);
xnor U19759 (N_19759,N_12037,N_11587);
or U19760 (N_19760,N_12590,N_12654);
nand U19761 (N_19761,N_11095,N_10325);
nor U19762 (N_19762,N_12514,N_11959);
nand U19763 (N_19763,N_11419,N_12007);
nor U19764 (N_19764,N_14670,N_12532);
nand U19765 (N_19765,N_12440,N_13055);
and U19766 (N_19766,N_14352,N_10332);
and U19767 (N_19767,N_13900,N_11453);
nand U19768 (N_19768,N_13429,N_11609);
or U19769 (N_19769,N_11649,N_10699);
nor U19770 (N_19770,N_13889,N_13658);
and U19771 (N_19771,N_14710,N_14072);
or U19772 (N_19772,N_11037,N_11911);
nand U19773 (N_19773,N_13640,N_10487);
nor U19774 (N_19774,N_11248,N_13059);
xor U19775 (N_19775,N_14512,N_12171);
and U19776 (N_19776,N_10351,N_14483);
nand U19777 (N_19777,N_10415,N_11015);
nand U19778 (N_19778,N_12524,N_11796);
xnor U19779 (N_19779,N_12316,N_11002);
or U19780 (N_19780,N_11099,N_11511);
xor U19781 (N_19781,N_10019,N_11321);
nor U19782 (N_19782,N_12069,N_10216);
xnor U19783 (N_19783,N_13674,N_12226);
xnor U19784 (N_19784,N_13241,N_12008);
nor U19785 (N_19785,N_13723,N_14724);
nand U19786 (N_19786,N_13068,N_14400);
nor U19787 (N_19787,N_14346,N_10617);
nor U19788 (N_19788,N_12182,N_11375);
xor U19789 (N_19789,N_10597,N_14371);
and U19790 (N_19790,N_10269,N_13506);
nor U19791 (N_19791,N_12522,N_12225);
and U19792 (N_19792,N_14677,N_14733);
nand U19793 (N_19793,N_11661,N_10604);
nor U19794 (N_19794,N_11629,N_13485);
or U19795 (N_19795,N_13614,N_12220);
or U19796 (N_19796,N_11830,N_10073);
nand U19797 (N_19797,N_12195,N_12718);
xor U19798 (N_19798,N_10898,N_12392);
or U19799 (N_19799,N_12415,N_12807);
nor U19800 (N_19800,N_12061,N_10990);
xor U19801 (N_19801,N_11525,N_14250);
or U19802 (N_19802,N_13987,N_11561);
nand U19803 (N_19803,N_13928,N_13147);
or U19804 (N_19804,N_14959,N_14702);
xor U19805 (N_19805,N_10271,N_11175);
nor U19806 (N_19806,N_12235,N_12418);
xor U19807 (N_19807,N_10213,N_13353);
nor U19808 (N_19808,N_12640,N_10541);
or U19809 (N_19809,N_14480,N_12090);
or U19810 (N_19810,N_10000,N_14410);
nand U19811 (N_19811,N_12489,N_13318);
or U19812 (N_19812,N_10498,N_13687);
nand U19813 (N_19813,N_12260,N_11626);
xnor U19814 (N_19814,N_14920,N_10934);
and U19815 (N_19815,N_14590,N_11279);
or U19816 (N_19816,N_10484,N_10373);
nand U19817 (N_19817,N_14045,N_10259);
xor U19818 (N_19818,N_14575,N_12649);
nand U19819 (N_19819,N_13745,N_14297);
nor U19820 (N_19820,N_12970,N_10472);
nor U19821 (N_19821,N_10399,N_13230);
xnor U19822 (N_19822,N_11404,N_14963);
or U19823 (N_19823,N_10240,N_11209);
and U19824 (N_19824,N_10414,N_14842);
nor U19825 (N_19825,N_12993,N_13891);
or U19826 (N_19826,N_12208,N_14926);
and U19827 (N_19827,N_11884,N_10219);
and U19828 (N_19828,N_14731,N_12442);
nor U19829 (N_19829,N_13742,N_10266);
or U19830 (N_19830,N_12444,N_10121);
nor U19831 (N_19831,N_12517,N_14857);
xor U19832 (N_19832,N_12741,N_11964);
nor U19833 (N_19833,N_11970,N_11073);
nand U19834 (N_19834,N_11416,N_11533);
nor U19835 (N_19835,N_14530,N_11892);
nor U19836 (N_19836,N_14882,N_12493);
nor U19837 (N_19837,N_13987,N_14295);
and U19838 (N_19838,N_10491,N_10530);
xnor U19839 (N_19839,N_10837,N_11908);
and U19840 (N_19840,N_13687,N_13826);
and U19841 (N_19841,N_13214,N_12723);
nor U19842 (N_19842,N_12225,N_10631);
or U19843 (N_19843,N_14366,N_13721);
nand U19844 (N_19844,N_13206,N_13183);
xor U19845 (N_19845,N_14492,N_11673);
nand U19846 (N_19846,N_12722,N_10716);
or U19847 (N_19847,N_12294,N_12030);
xnor U19848 (N_19848,N_14591,N_10689);
nor U19849 (N_19849,N_11725,N_10855);
nor U19850 (N_19850,N_11132,N_10131);
nand U19851 (N_19851,N_13816,N_10628);
nand U19852 (N_19852,N_10887,N_10171);
or U19853 (N_19853,N_14571,N_13846);
nor U19854 (N_19854,N_13191,N_10566);
or U19855 (N_19855,N_13084,N_13838);
xor U19856 (N_19856,N_12177,N_14983);
and U19857 (N_19857,N_13250,N_12053);
xnor U19858 (N_19858,N_10432,N_10387);
nand U19859 (N_19859,N_10143,N_14359);
or U19860 (N_19860,N_13924,N_10220);
xor U19861 (N_19861,N_13980,N_10873);
nand U19862 (N_19862,N_14826,N_10735);
xnor U19863 (N_19863,N_11689,N_12813);
and U19864 (N_19864,N_10664,N_13097);
xnor U19865 (N_19865,N_12864,N_13493);
nor U19866 (N_19866,N_11335,N_10023);
or U19867 (N_19867,N_14159,N_10696);
nand U19868 (N_19868,N_11507,N_14928);
xnor U19869 (N_19869,N_13967,N_10016);
and U19870 (N_19870,N_10291,N_13953);
xnor U19871 (N_19871,N_10477,N_11564);
and U19872 (N_19872,N_10810,N_11428);
xor U19873 (N_19873,N_14206,N_14877);
and U19874 (N_19874,N_12658,N_11660);
nand U19875 (N_19875,N_14351,N_10439);
nor U19876 (N_19876,N_14240,N_13751);
xor U19877 (N_19877,N_13543,N_12089);
nand U19878 (N_19878,N_14525,N_12517);
xor U19879 (N_19879,N_13585,N_14231);
xor U19880 (N_19880,N_13814,N_10381);
nand U19881 (N_19881,N_10723,N_10735);
or U19882 (N_19882,N_14124,N_14899);
xor U19883 (N_19883,N_11684,N_14009);
xnor U19884 (N_19884,N_12809,N_10756);
or U19885 (N_19885,N_13866,N_11634);
nor U19886 (N_19886,N_13543,N_11127);
xor U19887 (N_19887,N_13705,N_12119);
xor U19888 (N_19888,N_13347,N_12450);
nor U19889 (N_19889,N_12457,N_14193);
and U19890 (N_19890,N_14444,N_11894);
nand U19891 (N_19891,N_14453,N_13818);
nor U19892 (N_19892,N_13969,N_11450);
nor U19893 (N_19893,N_12887,N_14637);
or U19894 (N_19894,N_10664,N_14840);
xnor U19895 (N_19895,N_14192,N_13324);
nor U19896 (N_19896,N_14824,N_14614);
and U19897 (N_19897,N_10747,N_10771);
nor U19898 (N_19898,N_12077,N_13438);
and U19899 (N_19899,N_13738,N_12189);
nand U19900 (N_19900,N_14840,N_11612);
xor U19901 (N_19901,N_11849,N_13259);
nor U19902 (N_19902,N_11639,N_13776);
nor U19903 (N_19903,N_12847,N_12872);
xnor U19904 (N_19904,N_11950,N_12207);
nor U19905 (N_19905,N_12790,N_12347);
nand U19906 (N_19906,N_13246,N_13817);
xor U19907 (N_19907,N_14065,N_12921);
xor U19908 (N_19908,N_12138,N_14267);
or U19909 (N_19909,N_14149,N_13105);
or U19910 (N_19910,N_13303,N_12609);
xnor U19911 (N_19911,N_12700,N_11084);
nand U19912 (N_19912,N_10109,N_14396);
xnor U19913 (N_19913,N_10828,N_13713);
xnor U19914 (N_19914,N_14412,N_13888);
xnor U19915 (N_19915,N_14133,N_11774);
nor U19916 (N_19916,N_10463,N_10744);
or U19917 (N_19917,N_11843,N_10955);
xor U19918 (N_19918,N_14376,N_12669);
nand U19919 (N_19919,N_12027,N_14683);
nand U19920 (N_19920,N_14871,N_10235);
or U19921 (N_19921,N_13104,N_14169);
nand U19922 (N_19922,N_14127,N_14071);
nor U19923 (N_19923,N_14932,N_12269);
xnor U19924 (N_19924,N_12364,N_14223);
nand U19925 (N_19925,N_14605,N_10724);
nor U19926 (N_19926,N_12327,N_10880);
nor U19927 (N_19927,N_14376,N_11649);
xor U19928 (N_19928,N_12168,N_12206);
nand U19929 (N_19929,N_14817,N_10734);
nor U19930 (N_19930,N_10192,N_13899);
and U19931 (N_19931,N_13565,N_13197);
or U19932 (N_19932,N_12615,N_14066);
and U19933 (N_19933,N_12381,N_10819);
xor U19934 (N_19934,N_10448,N_14323);
nand U19935 (N_19935,N_13652,N_14786);
xor U19936 (N_19936,N_12918,N_13224);
or U19937 (N_19937,N_12301,N_10467);
and U19938 (N_19938,N_10421,N_13584);
nor U19939 (N_19939,N_10812,N_13902);
or U19940 (N_19940,N_13684,N_12221);
or U19941 (N_19941,N_13710,N_10442);
and U19942 (N_19942,N_12928,N_14744);
and U19943 (N_19943,N_12320,N_12650);
nand U19944 (N_19944,N_13398,N_11995);
xor U19945 (N_19945,N_12750,N_13832);
xor U19946 (N_19946,N_14120,N_10905);
and U19947 (N_19947,N_13486,N_13242);
xnor U19948 (N_19948,N_11210,N_10021);
xnor U19949 (N_19949,N_13358,N_13482);
nor U19950 (N_19950,N_11448,N_11294);
nor U19951 (N_19951,N_13452,N_10200);
nand U19952 (N_19952,N_10998,N_13932);
or U19953 (N_19953,N_10894,N_13725);
and U19954 (N_19954,N_12723,N_12140);
and U19955 (N_19955,N_10436,N_12770);
nand U19956 (N_19956,N_13534,N_11890);
nand U19957 (N_19957,N_12048,N_10977);
or U19958 (N_19958,N_12819,N_14908);
nand U19959 (N_19959,N_11352,N_13959);
and U19960 (N_19960,N_14856,N_10711);
and U19961 (N_19961,N_13077,N_10618);
nor U19962 (N_19962,N_14204,N_12606);
and U19963 (N_19963,N_13481,N_12270);
nand U19964 (N_19964,N_11931,N_10110);
and U19965 (N_19965,N_10273,N_14792);
nand U19966 (N_19966,N_12899,N_13546);
nor U19967 (N_19967,N_10344,N_13304);
nand U19968 (N_19968,N_10899,N_11836);
and U19969 (N_19969,N_14480,N_14309);
and U19970 (N_19970,N_12435,N_13777);
nand U19971 (N_19971,N_12351,N_11545);
or U19972 (N_19972,N_10145,N_13554);
xnor U19973 (N_19973,N_13984,N_14256);
or U19974 (N_19974,N_10958,N_10363);
and U19975 (N_19975,N_11703,N_12083);
and U19976 (N_19976,N_14083,N_11225);
and U19977 (N_19977,N_10663,N_11260);
and U19978 (N_19978,N_12063,N_14490);
nor U19979 (N_19979,N_11248,N_11775);
xnor U19980 (N_19980,N_11263,N_12158);
and U19981 (N_19981,N_10750,N_13935);
nor U19982 (N_19982,N_14452,N_11697);
nor U19983 (N_19983,N_12160,N_12420);
and U19984 (N_19984,N_12522,N_10155);
nor U19985 (N_19985,N_12500,N_10955);
and U19986 (N_19986,N_12594,N_13989);
or U19987 (N_19987,N_12323,N_11198);
or U19988 (N_19988,N_12078,N_11769);
nor U19989 (N_19989,N_11218,N_13820);
xor U19990 (N_19990,N_13206,N_14231);
xnor U19991 (N_19991,N_12861,N_14324);
or U19992 (N_19992,N_14406,N_10285);
xor U19993 (N_19993,N_11592,N_13035);
xnor U19994 (N_19994,N_11839,N_13143);
and U19995 (N_19995,N_13624,N_10888);
or U19996 (N_19996,N_10527,N_14475);
and U19997 (N_19997,N_12277,N_12504);
nor U19998 (N_19998,N_13147,N_12367);
nor U19999 (N_19999,N_11772,N_14111);
xnor U20000 (N_20000,N_15828,N_17257);
nand U20001 (N_20001,N_16126,N_17462);
and U20002 (N_20002,N_16394,N_15080);
nor U20003 (N_20003,N_17033,N_17305);
and U20004 (N_20004,N_17306,N_17669);
nor U20005 (N_20005,N_15806,N_15062);
nor U20006 (N_20006,N_18131,N_15341);
and U20007 (N_20007,N_18606,N_18956);
nor U20008 (N_20008,N_16578,N_19177);
nand U20009 (N_20009,N_17429,N_15006);
nand U20010 (N_20010,N_19517,N_16015);
and U20011 (N_20011,N_15183,N_17722);
or U20012 (N_20012,N_16145,N_16908);
nor U20013 (N_20013,N_15135,N_18079);
xor U20014 (N_20014,N_17707,N_15695);
xor U20015 (N_20015,N_19127,N_17977);
nand U20016 (N_20016,N_18050,N_16116);
xnor U20017 (N_20017,N_18226,N_18347);
nand U20018 (N_20018,N_17232,N_19534);
and U20019 (N_20019,N_19468,N_18355);
nand U20020 (N_20020,N_19744,N_19384);
xor U20021 (N_20021,N_17592,N_16541);
and U20022 (N_20022,N_19324,N_16942);
nor U20023 (N_20023,N_17616,N_17629);
nand U20024 (N_20024,N_17425,N_19240);
nor U20025 (N_20025,N_16437,N_17087);
or U20026 (N_20026,N_15603,N_17471);
nand U20027 (N_20027,N_18857,N_16156);
or U20028 (N_20028,N_19942,N_17521);
xor U20029 (N_20029,N_15969,N_19603);
or U20030 (N_20030,N_19228,N_16695);
and U20031 (N_20031,N_15994,N_17350);
nor U20032 (N_20032,N_16353,N_15844);
and U20033 (N_20033,N_19952,N_17825);
or U20034 (N_20034,N_18900,N_19274);
or U20035 (N_20035,N_17203,N_19890);
nor U20036 (N_20036,N_17703,N_19577);
or U20037 (N_20037,N_16893,N_16043);
or U20038 (N_20038,N_19141,N_16177);
and U20039 (N_20039,N_18498,N_19895);
or U20040 (N_20040,N_19773,N_16565);
nand U20041 (N_20041,N_19040,N_19082);
xnor U20042 (N_20042,N_16768,N_17795);
and U20043 (N_20043,N_16740,N_19333);
xnor U20044 (N_20044,N_19278,N_18640);
or U20045 (N_20045,N_18584,N_17240);
and U20046 (N_20046,N_19451,N_18962);
or U20047 (N_20047,N_19041,N_18631);
nand U20048 (N_20048,N_19501,N_18400);
or U20049 (N_20049,N_18294,N_18968);
nor U20050 (N_20050,N_16775,N_19339);
xor U20051 (N_20051,N_15978,N_15993);
or U20052 (N_20052,N_19039,N_17134);
and U20053 (N_20053,N_19677,N_18500);
nand U20054 (N_20054,N_19230,N_16932);
and U20055 (N_20055,N_19899,N_16644);
and U20056 (N_20056,N_18946,N_17765);
nand U20057 (N_20057,N_19802,N_16602);
nor U20058 (N_20058,N_15666,N_16431);
or U20059 (N_20059,N_18978,N_15626);
nand U20060 (N_20060,N_19365,N_16767);
nor U20061 (N_20061,N_19212,N_15084);
nand U20062 (N_20062,N_15032,N_15344);
and U20063 (N_20063,N_18685,N_17009);
nand U20064 (N_20064,N_15177,N_18883);
nor U20065 (N_20065,N_19017,N_19107);
or U20066 (N_20066,N_16389,N_16570);
nor U20067 (N_20067,N_16914,N_19815);
nand U20068 (N_20068,N_15000,N_18981);
xor U20069 (N_20069,N_17981,N_17072);
nand U20070 (N_20070,N_16397,N_17205);
nor U20071 (N_20071,N_18613,N_15742);
and U20072 (N_20072,N_18239,N_17299);
and U20073 (N_20073,N_15625,N_17901);
or U20074 (N_20074,N_17896,N_18053);
and U20075 (N_20075,N_15448,N_18545);
and U20076 (N_20076,N_15877,N_16297);
or U20077 (N_20077,N_18320,N_17782);
and U20078 (N_20078,N_16623,N_15759);
nand U20079 (N_20079,N_18394,N_19345);
and U20080 (N_20080,N_17097,N_15332);
and U20081 (N_20081,N_16113,N_17856);
or U20082 (N_20082,N_19977,N_15165);
and U20083 (N_20083,N_15789,N_16037);
or U20084 (N_20084,N_18417,N_15951);
or U20085 (N_20085,N_19659,N_19200);
nor U20086 (N_20086,N_17950,N_16948);
nor U20087 (N_20087,N_16143,N_19223);
or U20088 (N_20088,N_19596,N_17530);
xor U20089 (N_20089,N_15971,N_17958);
nand U20090 (N_20090,N_15280,N_19676);
xor U20091 (N_20091,N_19221,N_19442);
xor U20092 (N_20092,N_19767,N_17286);
nand U20093 (N_20093,N_16757,N_15707);
and U20094 (N_20094,N_17103,N_17060);
and U20095 (N_20095,N_18015,N_19612);
nor U20096 (N_20096,N_19555,N_18650);
nand U20097 (N_20097,N_17415,N_18827);
or U20098 (N_20098,N_19715,N_16918);
or U20099 (N_20099,N_16165,N_16664);
nor U20100 (N_20100,N_15967,N_16419);
and U20101 (N_20101,N_15073,N_17440);
nand U20102 (N_20102,N_19825,N_17720);
xor U20103 (N_20103,N_16737,N_18469);
nor U20104 (N_20104,N_15437,N_19997);
nor U20105 (N_20105,N_17672,N_17442);
nand U20106 (N_20106,N_19858,N_17389);
xnor U20107 (N_20107,N_16211,N_17322);
nand U20108 (N_20108,N_19428,N_18295);
xor U20109 (N_20109,N_19933,N_16373);
xnor U20110 (N_20110,N_16702,N_18281);
xor U20111 (N_20111,N_18728,N_15316);
and U20112 (N_20112,N_19377,N_19828);
xnor U20113 (N_20113,N_15433,N_17964);
or U20114 (N_20114,N_17690,N_18527);
and U20115 (N_20115,N_15069,N_17576);
nand U20116 (N_20116,N_15168,N_16903);
and U20117 (N_20117,N_15431,N_19335);
nand U20118 (N_20118,N_19382,N_19764);
nor U20119 (N_20119,N_19235,N_18261);
nand U20120 (N_20120,N_15892,N_16136);
and U20121 (N_20121,N_18162,N_18308);
nor U20122 (N_20122,N_17968,N_16386);
or U20123 (N_20123,N_19803,N_19196);
and U20124 (N_20124,N_16745,N_19188);
and U20125 (N_20125,N_19669,N_15455);
and U20126 (N_20126,N_18198,N_17413);
or U20127 (N_20127,N_16503,N_18032);
and U20128 (N_20128,N_17477,N_19700);
nand U20129 (N_20129,N_18003,N_19472);
nand U20130 (N_20130,N_16473,N_18448);
and U20131 (N_20131,N_19558,N_16657);
xor U20132 (N_20132,N_16176,N_17225);
and U20133 (N_20133,N_17379,N_16945);
and U20134 (N_20134,N_18271,N_18621);
nand U20135 (N_20135,N_15458,N_16417);
and U20136 (N_20136,N_16264,N_16205);
xor U20137 (N_20137,N_18174,N_15182);
and U20138 (N_20138,N_17279,N_15764);
xor U20139 (N_20139,N_18642,N_16303);
and U20140 (N_20140,N_15560,N_18231);
or U20141 (N_20141,N_17952,N_19594);
and U20142 (N_20142,N_18412,N_15247);
and U20143 (N_20143,N_18307,N_18878);
xnor U20144 (N_20144,N_16208,N_19046);
or U20145 (N_20145,N_18585,N_16554);
or U20146 (N_20146,N_19503,N_17406);
xor U20147 (N_20147,N_19537,N_16278);
nand U20148 (N_20148,N_18887,N_18848);
and U20149 (N_20149,N_19824,N_19128);
or U20150 (N_20150,N_16754,N_16593);
nor U20151 (N_20151,N_19661,N_18430);
or U20152 (N_20152,N_15788,N_19795);
xor U20153 (N_20153,N_18392,N_17126);
or U20154 (N_20154,N_17417,N_16468);
xnor U20155 (N_20155,N_15596,N_19204);
nor U20156 (N_20156,N_16484,N_18866);
nand U20157 (N_20157,N_19598,N_15571);
or U20158 (N_20158,N_17011,N_15819);
and U20159 (N_20159,N_15675,N_18672);
xnor U20160 (N_20160,N_17271,N_16069);
nor U20161 (N_20161,N_15685,N_18507);
nand U20162 (N_20162,N_15623,N_16817);
and U20163 (N_20163,N_19801,N_15134);
xnor U20164 (N_20164,N_17872,N_15852);
or U20165 (N_20165,N_17817,N_19882);
or U20166 (N_20166,N_15882,N_16694);
or U20167 (N_20167,N_17906,N_16319);
nor U20168 (N_20168,N_16540,N_15397);
and U20169 (N_20169,N_19863,N_15331);
nand U20170 (N_20170,N_18305,N_15770);
and U20171 (N_20171,N_16689,N_18403);
xnor U20172 (N_20172,N_19610,N_16543);
or U20173 (N_20173,N_15992,N_19009);
or U20174 (N_20174,N_15412,N_17553);
xnor U20175 (N_20175,N_15519,N_17273);
or U20176 (N_20176,N_18599,N_18197);
nor U20177 (N_20177,N_16349,N_19967);
or U20178 (N_20178,N_19341,N_18370);
nor U20179 (N_20179,N_18321,N_16718);
nand U20180 (N_20180,N_17432,N_19330);
nor U20181 (N_20181,N_17976,N_16998);
and U20182 (N_20182,N_19742,N_19607);
xnor U20183 (N_20183,N_19735,N_17633);
or U20184 (N_20184,N_15867,N_15775);
nor U20185 (N_20185,N_18068,N_15481);
nor U20186 (N_20186,N_19761,N_18770);
nand U20187 (N_20187,N_19402,N_16844);
or U20188 (N_20188,N_15320,N_16339);
xor U20189 (N_20189,N_15120,N_16697);
or U20190 (N_20190,N_17280,N_17871);
and U20191 (N_20191,N_15900,N_16666);
or U20192 (N_20192,N_18628,N_16151);
nor U20193 (N_20193,N_16010,N_18011);
and U20194 (N_20194,N_16816,N_17724);
or U20195 (N_20195,N_18562,N_17176);
and U20196 (N_20196,N_17171,N_15615);
or U20197 (N_20197,N_15715,N_18526);
and U20198 (N_20198,N_15096,N_16904);
or U20199 (N_20199,N_16446,N_18762);
xnor U20200 (N_20200,N_16510,N_17207);
xnor U20201 (N_20201,N_18105,N_15921);
and U20202 (N_20202,N_15386,N_17730);
or U20203 (N_20203,N_19785,N_15029);
nor U20204 (N_20204,N_16239,N_15104);
or U20205 (N_20205,N_17465,N_19937);
nor U20206 (N_20206,N_15855,N_15093);
xnor U20207 (N_20207,N_15935,N_15224);
and U20208 (N_20208,N_18961,N_16036);
nand U20209 (N_20209,N_18021,N_19894);
nand U20210 (N_20210,N_17885,N_19461);
and U20211 (N_20211,N_19794,N_15474);
or U20212 (N_20212,N_19300,N_19826);
nor U20213 (N_20213,N_18004,N_18429);
or U20214 (N_20214,N_17975,N_17942);
xnor U20215 (N_20215,N_19456,N_15003);
or U20216 (N_20216,N_18066,N_17926);
nand U20217 (N_20217,N_15575,N_18408);
or U20218 (N_20218,N_16430,N_17927);
and U20219 (N_20219,N_16444,N_16246);
nor U20220 (N_20220,N_16714,N_19478);
or U20221 (N_20221,N_17581,N_15310);
or U20222 (N_20222,N_17555,N_16636);
xor U20223 (N_20223,N_19689,N_15799);
nand U20224 (N_20224,N_15010,N_18907);
nor U20225 (N_20225,N_19851,N_15576);
and U20226 (N_20226,N_19307,N_19615);
xor U20227 (N_20227,N_17626,N_15534);
xor U20228 (N_20228,N_15972,N_19736);
or U20229 (N_20229,N_17188,N_15905);
and U20230 (N_20230,N_17735,N_16777);
nand U20231 (N_20231,N_17229,N_19780);
nor U20232 (N_20232,N_17421,N_17371);
xnor U20233 (N_20233,N_15249,N_19315);
nand U20234 (N_20234,N_17740,N_18084);
or U20235 (N_20235,N_16392,N_15434);
nand U20236 (N_20236,N_17061,N_18283);
nor U20237 (N_20237,N_16162,N_19508);
xnor U20238 (N_20238,N_16438,N_18476);
and U20239 (N_20239,N_17805,N_16832);
nand U20240 (N_20240,N_15542,N_18553);
xor U20241 (N_20241,N_18675,N_16995);
and U20242 (N_20242,N_18252,N_15917);
nor U20243 (N_20243,N_17456,N_16361);
xnor U20244 (N_20244,N_16171,N_19309);
or U20245 (N_20245,N_18279,N_19163);
xnor U20246 (N_20246,N_17838,N_18451);
xor U20247 (N_20247,N_15698,N_17353);
xnor U20248 (N_20248,N_15863,N_16423);
xor U20249 (N_20249,N_17631,N_19550);
nor U20250 (N_20250,N_19004,N_18348);
xor U20251 (N_20251,N_17044,N_15377);
xnor U20252 (N_20252,N_18738,N_18737);
or U20253 (N_20253,N_18285,N_18077);
nor U20254 (N_20254,N_16288,N_19648);
nand U20255 (N_20255,N_19605,N_18707);
nand U20256 (N_20256,N_15952,N_17598);
nor U20257 (N_20257,N_16333,N_15837);
and U20258 (N_20258,N_18176,N_18472);
or U20259 (N_20259,N_16838,N_19155);
and U20260 (N_20260,N_16121,N_15725);
nand U20261 (N_20261,N_15447,N_15758);
nand U20262 (N_20262,N_17049,N_19123);
or U20263 (N_20263,N_15420,N_18572);
and U20264 (N_20264,N_16490,N_15628);
and U20265 (N_20265,N_18413,N_17219);
nand U20266 (N_20266,N_15955,N_17113);
nand U20267 (N_20267,N_15800,N_17727);
or U20268 (N_20268,N_15903,N_16317);
or U20269 (N_20269,N_18892,N_18835);
or U20270 (N_20270,N_17936,N_18288);
and U20271 (N_20271,N_16003,N_17632);
or U20272 (N_20272,N_15147,N_17258);
nand U20273 (N_20273,N_17201,N_16704);
or U20274 (N_20274,N_18504,N_19674);
xor U20275 (N_20275,N_17121,N_17332);
and U20276 (N_20276,N_18998,N_17818);
xnor U20277 (N_20277,N_17954,N_15573);
nor U20278 (N_20278,N_16684,N_19088);
and U20279 (N_20279,N_19246,N_17062);
or U20280 (N_20280,N_15213,N_18262);
and U20281 (N_20281,N_17947,N_16762);
or U20282 (N_20282,N_17863,N_17491);
nor U20283 (N_20283,N_15973,N_17552);
nand U20284 (N_20284,N_17184,N_19632);
or U20285 (N_20285,N_18116,N_17233);
nor U20286 (N_20286,N_18576,N_19003);
xnor U20287 (N_20287,N_16830,N_15220);
and U20288 (N_20288,N_19255,N_17197);
or U20289 (N_20289,N_15647,N_19509);
nand U20290 (N_20290,N_18859,N_15704);
xor U20291 (N_20291,N_16577,N_17910);
and U20292 (N_20292,N_19265,N_18273);
nand U20293 (N_20293,N_17928,N_18521);
nor U20294 (N_20294,N_16861,N_19385);
nand U20295 (N_20295,N_18722,N_18618);
xnor U20296 (N_20296,N_19258,N_16294);
and U20297 (N_20297,N_19019,N_19301);
and U20298 (N_20298,N_15527,N_16994);
or U20299 (N_20299,N_15879,N_16743);
xor U20300 (N_20300,N_17120,N_19624);
nor U20301 (N_20301,N_18363,N_15208);
or U20302 (N_20302,N_19599,N_18950);
nor U20303 (N_20303,N_19282,N_17995);
nand U20304 (N_20304,N_18712,N_15400);
xor U20305 (N_20305,N_15008,N_15278);
or U20306 (N_20306,N_18677,N_19580);
nand U20307 (N_20307,N_18118,N_19688);
or U20308 (N_20308,N_19470,N_18756);
nand U20309 (N_20309,N_18780,N_17221);
xor U20310 (N_20310,N_19374,N_15621);
nand U20311 (N_20311,N_17094,N_19343);
xor U20312 (N_20312,N_16677,N_17574);
nor U20313 (N_20313,N_19419,N_19471);
or U20314 (N_20314,N_15588,N_15736);
and U20315 (N_20315,N_18838,N_17348);
or U20316 (N_20316,N_17937,N_19914);
xnor U20317 (N_20317,N_16659,N_17766);
nand U20318 (N_20318,N_16669,N_16035);
nor U20319 (N_20319,N_18212,N_19299);
xor U20320 (N_20320,N_18888,N_15276);
and U20321 (N_20321,N_18164,N_18577);
or U20322 (N_20322,N_16911,N_19367);
xnor U20323 (N_20323,N_17250,N_17640);
or U20324 (N_20324,N_19955,N_16026);
nand U20325 (N_20325,N_16011,N_17495);
xor U20326 (N_20326,N_16594,N_16481);
xor U20327 (N_20327,N_15059,N_18735);
and U20328 (N_20328,N_17401,N_17627);
xor U20329 (N_20329,N_16849,N_15470);
or U20330 (N_20330,N_18227,N_18616);
or U20331 (N_20331,N_16933,N_18991);
xnor U20332 (N_20332,N_16382,N_18902);
or U20333 (N_20333,N_19837,N_16040);
xnor U20334 (N_20334,N_16452,N_18366);
and U20335 (N_20335,N_15257,N_17122);
nand U20336 (N_20336,N_18201,N_16814);
and U20337 (N_20337,N_16915,N_18985);
or U20338 (N_20338,N_16358,N_16158);
nor U20339 (N_20339,N_19245,N_15579);
xnor U20340 (N_20340,N_16458,N_15078);
nand U20341 (N_20341,N_18692,N_16321);
and U20342 (N_20342,N_15030,N_17510);
xor U20343 (N_20343,N_19636,N_19835);
xnor U20344 (N_20344,N_18155,N_16440);
xor U20345 (N_20345,N_18027,N_19027);
xor U20346 (N_20346,N_19467,N_17951);
nor U20347 (N_20347,N_15307,N_16189);
nor U20348 (N_20348,N_17677,N_18699);
xnor U20349 (N_20349,N_19585,N_17961);
nand U20350 (N_20350,N_19668,N_19005);
nor U20351 (N_20351,N_16277,N_16831);
or U20352 (N_20352,N_18525,N_19465);
nor U20353 (N_20353,N_17617,N_18942);
xnor U20354 (N_20354,N_17535,N_17761);
and U20355 (N_20355,N_19956,N_15347);
nor U20356 (N_20356,N_16075,N_19368);
nor U20357 (N_20357,N_17738,N_16407);
and U20358 (N_20358,N_15670,N_19125);
nand U20359 (N_20359,N_19076,N_15506);
xor U20360 (N_20360,N_16311,N_17959);
nor U20361 (N_20361,N_17053,N_17443);
nor U20362 (N_20362,N_17355,N_19947);
or U20363 (N_20363,N_16390,N_15658);
xnor U20364 (N_20364,N_15569,N_15211);
or U20365 (N_20365,N_15330,N_15430);
nand U20366 (N_20366,N_19173,N_16885);
or U20367 (N_20367,N_15997,N_15097);
and U20368 (N_20368,N_19342,N_18767);
or U20369 (N_20369,N_15387,N_17948);
nor U20370 (N_20370,N_19812,N_17822);
and U20371 (N_20371,N_19178,N_17015);
nor U20372 (N_20372,N_19813,N_15604);
nor U20373 (N_20373,N_16429,N_15733);
or U20374 (N_20374,N_19552,N_15530);
xor U20375 (N_20375,N_18852,N_19533);
or U20376 (N_20376,N_17316,N_19256);
nand U20377 (N_20377,N_18223,N_19151);
and U20378 (N_20378,N_19182,N_16693);
and U20379 (N_20379,N_17281,N_19216);
or U20380 (N_20380,N_18931,N_15755);
nand U20381 (N_20381,N_16715,N_19346);
or U20382 (N_20382,N_16675,N_19816);
nor U20383 (N_20383,N_16204,N_16272);
nand U20384 (N_20384,N_19433,N_15501);
nand U20385 (N_20385,N_17602,N_17043);
nor U20386 (N_20386,N_18199,N_17372);
or U20387 (N_20387,N_15139,N_19979);
xor U20388 (N_20388,N_18581,N_16557);
nor U20389 (N_20389,N_19980,N_15118);
or U20390 (N_20390,N_18739,N_17891);
xor U20391 (N_20391,N_19353,N_15049);
nor U20392 (N_20392,N_17580,N_15904);
xor U20393 (N_20393,N_19043,N_15500);
xnor U20394 (N_20394,N_16462,N_19165);
nor U20395 (N_20395,N_18668,N_18594);
and U20396 (N_20396,N_15688,N_17151);
and U20397 (N_20397,N_15261,N_17549);
nor U20398 (N_20398,N_18410,N_15061);
or U20399 (N_20399,N_18028,N_15677);
nand U20400 (N_20400,N_18546,N_17594);
xnor U20401 (N_20401,N_19189,N_18567);
nand U20402 (N_20402,N_16730,N_16878);
or U20403 (N_20403,N_19941,N_19793);
nand U20404 (N_20404,N_15174,N_18938);
or U20405 (N_20405,N_19650,N_16793);
xor U20406 (N_20406,N_19035,N_19719);
and U20407 (N_20407,N_16504,N_15730);
and U20408 (N_20408,N_18851,N_19628);
nand U20409 (N_20409,N_17635,N_16905);
nor U20410 (N_20410,N_16365,N_17636);
and U20411 (N_20411,N_15729,N_17068);
nand U20412 (N_20412,N_18399,N_17347);
xnor U20413 (N_20413,N_15805,N_15929);
xnor U20414 (N_20414,N_18751,N_19732);
nor U20415 (N_20415,N_18067,N_19755);
or U20416 (N_20416,N_19587,N_15306);
nor U20417 (N_20417,N_16665,N_15954);
nand U20418 (N_20418,N_18119,N_15846);
nand U20419 (N_20419,N_17064,N_18580);
or U20420 (N_20420,N_15265,N_17212);
or U20421 (N_20421,N_16810,N_19388);
or U20422 (N_20422,N_18871,N_17892);
nor U20423 (N_20423,N_17460,N_16614);
nand U20424 (N_20424,N_19254,N_16424);
nand U20425 (N_20425,N_15121,N_17601);
or U20426 (N_20426,N_18579,N_19194);
nand U20427 (N_20427,N_19772,N_17275);
or U20428 (N_20428,N_17558,N_17014);
and U20429 (N_20429,N_15373,N_15262);
xor U20430 (N_20430,N_15482,N_15998);
xnor U20431 (N_20431,N_15129,N_15300);
nand U20432 (N_20432,N_18454,N_16313);
nor U20433 (N_20433,N_16865,N_17801);
nor U20434 (N_20434,N_19724,N_17793);
and U20435 (N_20435,N_18954,N_17994);
nand U20436 (N_20436,N_15081,N_18841);
xor U20437 (N_20437,N_15406,N_15283);
nor U20438 (N_20438,N_19693,N_17485);
and U20439 (N_20439,N_16428,N_18208);
or U20440 (N_20440,N_16985,N_17702);
or U20441 (N_20441,N_17753,N_17074);
nand U20442 (N_20442,N_16927,N_17705);
xor U20443 (N_20443,N_16142,N_16555);
and U20444 (N_20444,N_16085,N_19014);
nor U20445 (N_20445,N_19403,N_17701);
nand U20446 (N_20446,N_19690,N_17249);
or U20447 (N_20447,N_16184,N_17887);
nor U20448 (N_20448,N_19443,N_15175);
nand U20449 (N_20449,N_15614,N_16667);
nand U20450 (N_20450,N_16094,N_19294);
and U20451 (N_20451,N_15547,N_15378);
nor U20452 (N_20452,N_15925,N_18132);
nand U20453 (N_20453,N_15453,N_17422);
nor U20454 (N_20454,N_17373,N_17605);
nor U20455 (N_20455,N_16977,N_15637);
nand U20456 (N_20456,N_18427,N_17777);
and U20457 (N_20457,N_19413,N_19539);
and U20458 (N_20458,N_17459,N_16608);
or U20459 (N_20459,N_18639,N_17092);
nand U20460 (N_20460,N_18025,N_19175);
xor U20461 (N_20461,N_18730,N_15950);
xnor U20462 (N_20462,N_19934,N_15610);
nand U20463 (N_20463,N_17695,N_15056);
nor U20464 (N_20464,N_17454,N_17699);
nor U20465 (N_20465,N_19758,N_17609);
and U20466 (N_20466,N_18682,N_18783);
or U20467 (N_20467,N_18528,N_19568);
nand U20468 (N_20468,N_15618,N_16248);
nand U20469 (N_20469,N_19821,N_16856);
nor U20470 (N_20470,N_17827,N_17129);
xor U20471 (N_20471,N_18817,N_18860);
xor U20472 (N_20472,N_16898,N_17056);
and U20473 (N_20473,N_18194,N_16955);
nand U20474 (N_20474,N_18893,N_15878);
xnor U20475 (N_20475,N_16042,N_18957);
nor U20476 (N_20476,N_15605,N_16161);
nand U20477 (N_20477,N_15766,N_17828);
nor U20478 (N_20478,N_19257,N_15485);
nor U20479 (N_20479,N_15350,N_18578);
nor U20480 (N_20480,N_19789,N_16169);
or U20481 (N_20481,N_19065,N_18424);
nor U20482 (N_20482,N_17369,N_18123);
nor U20483 (N_20483,N_16725,N_19707);
or U20484 (N_20484,N_17354,N_17969);
xor U20485 (N_20485,N_15566,N_19407);
and U20486 (N_20486,N_18996,N_17577);
nand U20487 (N_20487,N_18072,N_17375);
nor U20488 (N_20488,N_17464,N_18135);
and U20489 (N_20489,N_18235,N_16393);
and U20490 (N_20490,N_16513,N_18372);
xor U20491 (N_20491,N_17813,N_17802);
and U20492 (N_20492,N_15737,N_17269);
nand U20493 (N_20493,N_18040,N_16147);
xor U20494 (N_20494,N_19024,N_16811);
nor U20495 (N_20495,N_16652,N_18651);
xor U20496 (N_20496,N_17161,N_19106);
nand U20497 (N_20497,N_18301,N_17693);
or U20498 (N_20498,N_18115,N_19412);
xor U20499 (N_20499,N_19126,N_16127);
and U20500 (N_20500,N_15502,N_17309);
xor U20501 (N_20501,N_18051,N_16640);
or U20502 (N_20502,N_17527,N_18541);
xnor U20503 (N_20503,N_15577,N_15325);
nand U20504 (N_20504,N_19132,N_19843);
nand U20505 (N_20505,N_16414,N_18010);
or U20506 (N_20506,N_19492,N_18849);
and U20507 (N_20507,N_19092,N_19809);
or U20508 (N_20508,N_19769,N_18736);
nand U20509 (N_20509,N_18204,N_17774);
and U20510 (N_20510,N_16864,N_15740);
and U20511 (N_20511,N_17451,N_17063);
or U20512 (N_20512,N_17096,N_17665);
or U20513 (N_20513,N_19518,N_18390);
xnor U20514 (N_20514,N_15918,N_16187);
nand U20515 (N_20515,N_18339,N_17963);
xor U20516 (N_20516,N_18192,N_19649);
xor U20517 (N_20517,N_15098,N_17715);
nor U20518 (N_20518,N_15239,N_16750);
xnor U20519 (N_20519,N_15808,N_19875);
nor U20520 (N_20520,N_16897,N_19960);
and U20521 (N_20521,N_18901,N_17550);
or U20522 (N_20522,N_18760,N_15411);
and U20523 (N_20523,N_17798,N_19572);
xor U20524 (N_20524,N_15977,N_18104);
or U20525 (N_20525,N_19010,N_17482);
or U20526 (N_20526,N_15233,N_18552);
and U20527 (N_20527,N_17143,N_15889);
and U20528 (N_20528,N_19919,N_16820);
nor U20529 (N_20529,N_15238,N_18912);
or U20530 (N_20530,N_19954,N_15234);
or U20531 (N_20531,N_15439,N_18565);
nor U20532 (N_20532,N_18514,N_16101);
xnor U20533 (N_20533,N_15367,N_19372);
xnor U20534 (N_20534,N_15505,N_16732);
xnor U20535 (N_20535,N_19531,N_16906);
nor U20536 (N_20536,N_17854,N_15333);
nand U20537 (N_20537,N_18471,N_17814);
and U20538 (N_20538,N_19383,N_15624);
nand U20539 (N_20539,N_16509,N_16213);
or U20540 (N_20540,N_18933,N_19766);
xnor U20541 (N_20541,N_18563,N_16781);
or U20542 (N_20542,N_17725,N_18516);
nor U20543 (N_20543,N_15457,N_16344);
or U20544 (N_20544,N_18943,N_18401);
xnor U20545 (N_20545,N_16783,N_15902);
xor U20546 (N_20546,N_18648,N_16526);
and U20547 (N_20547,N_19268,N_19847);
nor U20548 (N_20548,N_18600,N_17328);
or U20549 (N_20549,N_17528,N_18653);
and U20550 (N_20550,N_17775,N_17755);
or U20551 (N_20551,N_16708,N_18515);
or U20552 (N_20552,N_16108,N_15612);
nand U20553 (N_20553,N_19945,N_19381);
and U20554 (N_20554,N_15649,N_15021);
nor U20555 (N_20555,N_17559,N_18955);
and U20556 (N_20556,N_19994,N_19768);
or U20557 (N_20557,N_15317,N_18922);
xor U20558 (N_20558,N_18278,N_19595);
or U20559 (N_20559,N_17537,N_19202);
and U20560 (N_20560,N_18660,N_16801);
nor U20561 (N_20561,N_18512,N_19829);
xor U20562 (N_20562,N_17742,N_19015);
xor U20563 (N_20563,N_19239,N_17663);
nor U20564 (N_20564,N_16114,N_16448);
xnor U20565 (N_20565,N_17895,N_19654);
nand U20566 (N_20566,N_16658,N_15285);
nor U20567 (N_20567,N_16978,N_19340);
nor U20568 (N_20568,N_17533,N_18657);
or U20569 (N_20569,N_17127,N_15113);
xor U20570 (N_20570,N_16013,N_17523);
or U20571 (N_20571,N_18964,N_18326);
and U20572 (N_20572,N_19143,N_16135);
or U20573 (N_20573,N_15901,N_18329);
nand U20574 (N_20574,N_18406,N_19562);
or U20575 (N_20575,N_17189,N_15706);
nand U20576 (N_20576,N_17915,N_17595);
or U20577 (N_20577,N_18771,N_17048);
and U20578 (N_20578,N_17358,N_15150);
and U20579 (N_20579,N_15802,N_15741);
and U20580 (N_20580,N_18869,N_17603);
or U20581 (N_20581,N_18937,N_19020);
or U20582 (N_20582,N_17089,N_16599);
or U20583 (N_20583,N_19697,N_18254);
nor U20584 (N_20584,N_16427,N_17539);
nor U20585 (N_20585,N_18276,N_17943);
nor U20586 (N_20586,N_15845,N_18102);
xor U20587 (N_20587,N_15231,N_18464);
or U20588 (N_20588,N_19214,N_15692);
xor U20589 (N_20589,N_16131,N_18275);
nor U20590 (N_20590,N_15410,N_17772);
and U20591 (N_20591,N_16155,N_19331);
nand U20592 (N_20592,N_18814,N_15363);
or U20593 (N_20593,N_17771,N_18139);
nor U20594 (N_20594,N_15840,N_18853);
nor U20595 (N_20595,N_16221,N_19034);
xor U20596 (N_20596,N_17668,N_19298);
nor U20597 (N_20597,N_15319,N_18016);
nand U20598 (N_20598,N_16218,N_16776);
xor U20599 (N_20599,N_17119,N_15125);
nand U20600 (N_20600,N_18882,N_16241);
or U20601 (N_20601,N_15087,N_19756);
nor U20602 (N_20602,N_15751,N_18485);
and U20603 (N_20603,N_17327,N_16454);
nand U20604 (N_20604,N_18543,N_18744);
xor U20605 (N_20605,N_19946,N_18868);
and U20606 (N_20606,N_16456,N_17680);
xnor U20607 (N_20607,N_15348,N_17239);
nor U20608 (N_20608,N_15732,N_18941);
nand U20609 (N_20609,N_15620,N_16366);
or U20610 (N_20610,N_16167,N_16045);
nor U20611 (N_20611,N_19720,N_16639);
nor U20612 (N_20612,N_18409,N_15214);
nor U20613 (N_20613,N_17704,N_15197);
and U20614 (N_20614,N_18716,N_16283);
nand U20615 (N_20615,N_15767,N_18179);
nand U20616 (N_20616,N_16739,N_18256);
nor U20617 (N_20617,N_18490,N_17055);
nand U20618 (N_20618,N_16712,N_19989);
nor U20619 (N_20619,N_16613,N_15063);
and U20620 (N_20620,N_19459,N_16930);
xnor U20621 (N_20621,N_16687,N_15601);
and U20622 (N_20622,N_17167,N_18062);
and U20623 (N_20623,N_16546,N_15743);
nand U20624 (N_20624,N_17093,N_19117);
xnor U20625 (N_20625,N_16012,N_18260);
xnor U20626 (N_20626,N_19287,N_19376);
nor U20627 (N_20627,N_17153,N_16848);
or U20628 (N_20628,N_16356,N_16223);
nor U20629 (N_20629,N_18870,N_15219);
and U20630 (N_20630,N_19502,N_15240);
and U20631 (N_20631,N_17021,N_16600);
xnor U20632 (N_20632,N_19709,N_19757);
and U20633 (N_20633,N_16274,N_16713);
xnor U20634 (N_20634,N_17979,N_19704);
nand U20635 (N_20635,N_17248,N_16764);
xnor U20636 (N_20636,N_17728,N_18920);
or U20637 (N_20637,N_16959,N_19430);
and U20638 (N_20638,N_16092,N_19119);
nand U20639 (N_20639,N_15535,N_16335);
and U20640 (N_20640,N_19681,N_18436);
nor U20641 (N_20641,N_15380,N_15731);
or U20642 (N_20642,N_16269,N_16080);
nand U20643 (N_20643,N_15498,N_17430);
or U20644 (N_20644,N_15536,N_17960);
nand U20645 (N_20645,N_16785,N_17035);
nor U20646 (N_20646,N_16141,N_17295);
or U20647 (N_20647,N_19663,N_17208);
xnor U20648 (N_20648,N_18975,N_19679);
and U20649 (N_20649,N_17002,N_16471);
xnor U20650 (N_20650,N_17941,N_17847);
or U20651 (N_20651,N_16589,N_17411);
or U20652 (N_20652,N_17211,N_18665);
nor U20653 (N_20653,N_16926,N_17100);
and U20654 (N_20654,N_18786,N_17760);
nor U20655 (N_20655,N_18328,N_18414);
xor U20656 (N_20656,N_19739,N_15866);
nand U20657 (N_20657,N_18395,N_16398);
and U20658 (N_20658,N_19056,N_18804);
nand U20659 (N_20659,N_17517,N_16402);
and U20660 (N_20660,N_18322,N_15074);
nor U20661 (N_20661,N_19718,N_18894);
nor U20662 (N_20662,N_16572,N_18936);
and U20663 (N_20663,N_17058,N_15776);
nand U20664 (N_20664,N_15115,N_15026);
and U20665 (N_20665,N_15442,N_16952);
or U20666 (N_20666,N_16862,N_19510);
or U20667 (N_20667,N_18615,N_18564);
and U20668 (N_20668,N_17557,N_19423);
or U20669 (N_20669,N_19495,N_19932);
nor U20670 (N_20670,N_16773,N_18219);
and U20671 (N_20671,N_19526,N_17758);
xnor U20672 (N_20672,N_16808,N_19747);
and U20673 (N_20673,N_19929,N_15324);
xor U20674 (N_20674,N_17514,N_18874);
nand U20675 (N_20675,N_17418,N_16792);
or U20676 (N_20676,N_19665,N_17247);
or U20677 (N_20677,N_19187,N_19359);
or U20678 (N_20678,N_16784,N_15399);
and U20679 (N_20679,N_16710,N_18586);
nand U20680 (N_20680,N_17091,N_18847);
and U20681 (N_20681,N_19206,N_15040);
nand U20682 (N_20682,N_17090,N_18391);
xnor U20683 (N_20683,N_15826,N_17152);
xnor U20684 (N_20684,N_15641,N_18818);
nand U20685 (N_20685,N_15968,N_18625);
nand U20686 (N_20686,N_18713,N_19708);
xnor U20687 (N_20687,N_19957,N_17261);
nor U20688 (N_20688,N_15046,N_17792);
nor U20689 (N_20689,N_15757,N_15503);
and U20690 (N_20690,N_16609,N_16921);
xnor U20691 (N_20691,N_15369,N_16825);
nand U20692 (N_20692,N_16464,N_15172);
nand U20693 (N_20693,N_19917,N_17681);
and U20694 (N_20694,N_19564,N_19251);
and U20695 (N_20695,N_16005,N_16357);
and U20696 (N_20696,N_17660,N_15450);
nor U20697 (N_20697,N_16370,N_18732);
nor U20698 (N_20698,N_15223,N_19753);
nor U20699 (N_20699,N_19519,N_16564);
nor U20700 (N_20700,N_16273,N_17955);
nand U20701 (N_20701,N_17809,N_15110);
xor U20702 (N_20702,N_15148,N_17084);
nand U20703 (N_20703,N_17643,N_17455);
xor U20704 (N_20704,N_15714,N_18045);
nand U20705 (N_20705,N_15252,N_19168);
xor U20706 (N_20706,N_15717,N_17541);
nand U20707 (N_20707,N_17604,N_17732);
and U20708 (N_20708,N_19366,N_18556);
or U20709 (N_20709,N_17832,N_18063);
or U20710 (N_20710,N_17787,N_16795);
nor U20711 (N_20711,N_19623,N_18559);
xor U20712 (N_20712,N_15607,N_16050);
nor U20713 (N_20713,N_19507,N_18719);
nand U20714 (N_20714,N_19542,N_19996);
and U20715 (N_20715,N_18474,N_18979);
nand U20716 (N_20716,N_18125,N_18314);
and U20717 (N_20717,N_19896,N_16359);
xnor U20718 (N_20718,N_18168,N_15456);
nand U20719 (N_20719,N_15644,N_17815);
nand U20720 (N_20720,N_17177,N_17370);
or U20721 (N_20721,N_16262,N_17785);
xor U20722 (N_20722,N_18232,N_19449);
or U20723 (N_20723,N_19590,N_16046);
nand U20724 (N_20724,N_16822,N_16592);
nor U20725 (N_20725,N_19490,N_17343);
and U20726 (N_20726,N_19926,N_17839);
or U20727 (N_20727,N_17642,N_18537);
or U20728 (N_20728,N_15507,N_19738);
xnor U20729 (N_20729,N_15287,N_16829);
nand U20730 (N_20730,N_15792,N_19325);
xor U20731 (N_20731,N_19703,N_15192);
and U20732 (N_20732,N_15760,N_16826);
and U20733 (N_20733,N_15028,N_16122);
or U20734 (N_20734,N_15005,N_16511);
or U20735 (N_20735,N_19285,N_16835);
and U20736 (N_20736,N_17412,N_18608);
nand U20737 (N_20737,N_18317,N_19701);
xor U20738 (N_20738,N_18779,N_19390);
or U20739 (N_20739,N_17277,N_16220);
or U20740 (N_20740,N_16797,N_15484);
or U20741 (N_20741,N_16641,N_18548);
nand U20742 (N_20742,N_15354,N_16534);
or U20743 (N_20743,N_17365,N_15199);
nor U20744 (N_20744,N_19726,N_18896);
nor U20745 (N_20745,N_16362,N_19845);
nand U20746 (N_20746,N_19405,N_19897);
nand U20747 (N_20747,N_17536,N_15206);
or U20748 (N_20748,N_19401,N_17433);
and U20749 (N_20749,N_17700,N_15297);
and U20750 (N_20750,N_18180,N_19392);
nor U20751 (N_20751,N_17041,N_15613);
nand U20752 (N_20752,N_19488,N_16287);
xor U20753 (N_20753,N_19289,N_15164);
nor U20754 (N_20754,N_16200,N_16616);
and U20755 (N_20755,N_16160,N_18890);
or U20756 (N_20756,N_19975,N_18807);
xnor U20757 (N_20757,N_18747,N_15215);
or U20758 (N_20758,N_15678,N_16722);
nand U20759 (N_20759,N_15031,N_18133);
and U20760 (N_20760,N_16350,N_17905);
xor U20761 (N_20761,N_17990,N_19292);
nand U20762 (N_20762,N_16827,N_17911);
and U20763 (N_20763,N_15163,N_15424);
and U20764 (N_20764,N_19839,N_16336);
xnor U20765 (N_20765,N_15857,N_16173);
or U20766 (N_20766,N_15162,N_18984);
nand U20767 (N_20767,N_15681,N_15886);
or U20768 (N_20768,N_16916,N_17116);
xnor U20769 (N_20769,N_18324,N_18473);
or U20770 (N_20770,N_15833,N_18558);
nand U20771 (N_20771,N_15986,N_16191);
or U20772 (N_20772,N_15356,N_16420);
or U20773 (N_20773,N_16196,N_17245);
nor U20774 (N_20774,N_16671,N_17956);
nor U20775 (N_20775,N_15777,N_17980);
or U20776 (N_20776,N_19078,N_17242);
or U20777 (N_20777,N_15496,N_18466);
nand U20778 (N_20778,N_19397,N_15508);
and U20779 (N_20779,N_16175,N_15275);
or U20780 (N_20780,N_16633,N_15258);
nand U20781 (N_20781,N_17419,N_19486);
nor U20782 (N_20782,N_18723,N_15242);
nor U20783 (N_20783,N_15176,N_17263);
xor U20784 (N_20784,N_15691,N_19441);
nand U20785 (N_20785,N_15668,N_17107);
nor U20786 (N_20786,N_19971,N_16892);
nor U20787 (N_20787,N_16138,N_16065);
or U20788 (N_20788,N_17071,N_17163);
nor U20789 (N_20789,N_15512,N_18036);
nand U20790 (N_20790,N_19867,N_18478);
nand U20791 (N_20791,N_17834,N_18662);
nor U20792 (N_20792,N_15048,N_15746);
xor U20793 (N_20793,N_15472,N_16254);
nor U20794 (N_20794,N_18554,N_18935);
or U20795 (N_20795,N_16477,N_16182);
and U20796 (N_20796,N_19311,N_15171);
and U20797 (N_20797,N_16836,N_18623);
and U20798 (N_20798,N_19930,N_15014);
xor U20799 (N_20799,N_16632,N_16281);
or U20800 (N_20800,N_18056,N_17621);
nor U20801 (N_20801,N_18829,N_15723);
nand U20802 (N_20802,N_17858,N_19846);
xor U20803 (N_20803,N_19777,N_19538);
nand U20804 (N_20804,N_16699,N_19093);
and U20805 (N_20805,N_19122,N_16185);
or U20806 (N_20806,N_15368,N_15847);
nor U20807 (N_20807,N_19786,N_18169);
xnor U20808 (N_20808,N_18142,N_17849);
or U20809 (N_20809,N_17080,N_19008);
or U20810 (N_20810,N_18012,N_15862);
xor U20811 (N_20811,N_16771,N_18461);
nor U20812 (N_20812,N_16285,N_17483);
or U20813 (N_20813,N_16000,N_19903);
nor U20814 (N_20814,N_16960,N_18160);
and U20815 (N_20815,N_16755,N_19699);
xnor U20816 (N_20816,N_16323,N_15102);
nor U20817 (N_20817,N_16598,N_15036);
nand U20818 (N_20818,N_19678,N_18741);
nor U20819 (N_20819,N_17186,N_17141);
or U20820 (N_20820,N_18806,N_19481);
nor U20821 (N_20821,N_18972,N_17600);
and U20822 (N_20822,N_15018,N_15689);
and U20823 (N_20823,N_17622,N_16077);
and U20824 (N_20824,N_15816,N_15462);
and U20825 (N_20825,N_15851,N_16247);
or U20826 (N_20826,N_17256,N_18715);
xor U20827 (N_20827,N_17391,N_15157);
xor U20828 (N_20828,N_15159,N_18035);
nor U20829 (N_20829,N_17525,N_16987);
xor U20830 (N_20830,N_19347,N_19838);
and U20831 (N_20831,N_18568,N_16233);
nand U20832 (N_20832,N_16855,N_16535);
or U20833 (N_20833,N_16234,N_15103);
or U20834 (N_20834,N_18173,N_16243);
or U20835 (N_20835,N_17150,N_19030);
xor U20836 (N_20836,N_18557,N_18385);
and U20837 (N_20837,N_19608,N_19183);
or U20838 (N_20838,N_19589,N_18114);
and U20839 (N_20839,N_18691,N_16990);
nand U20840 (N_20840,N_15937,N_15835);
nor U20841 (N_20841,N_18149,N_15964);
nand U20842 (N_20842,N_16459,N_19276);
or U20843 (N_20843,N_18134,N_19184);
nor U20844 (N_20844,N_19528,N_15254);
nor U20845 (N_20845,N_19460,N_18593);
xor U20846 (N_20846,N_17984,N_18349);
xnor U20847 (N_20847,N_15629,N_15744);
and U20848 (N_20848,N_19631,N_17351);
nand U20849 (N_20849,N_17841,N_16581);
xnor U20850 (N_20850,N_16071,N_15394);
nor U20851 (N_20851,N_15091,N_18495);
and U20852 (N_20852,N_19439,N_16799);
or U20853 (N_20853,N_16660,N_18842);
nor U20854 (N_20854,N_19164,N_15067);
nand U20855 (N_20855,N_17685,N_15101);
nor U20856 (N_20856,N_18670,N_19243);
and U20857 (N_20857,N_18483,N_16940);
xnor U20858 (N_20858,N_18582,N_17781);
and U20859 (N_20859,N_15887,N_19609);
nor U20860 (N_20860,N_18666,N_18336);
nand U20861 (N_20861,N_15292,N_19080);
or U20862 (N_20862,N_17110,N_16934);
and U20863 (N_20863,N_19848,N_18315);
nand U20864 (N_20864,N_16819,N_19702);
or U20865 (N_20865,N_15592,N_16340);
and U20866 (N_20866,N_19427,N_19545);
nor U20867 (N_20867,N_18636,N_18834);
or U20868 (N_20868,N_15109,N_19541);
nand U20869 (N_20869,N_17136,N_19604);
nand U20870 (N_20870,N_18620,N_16859);
nand U20871 (N_20871,N_19166,N_19118);
and U20872 (N_20872,N_19849,N_15340);
and U20873 (N_20873,N_19808,N_18018);
nor U20874 (N_20874,N_15927,N_16874);
nor U20875 (N_20875,N_19549,N_15557);
xnor U20876 (N_20876,N_15346,N_15336);
and U20877 (N_20877,N_18238,N_18470);
nor U20878 (N_20878,N_16374,N_15822);
and U20879 (N_20879,N_15980,N_16225);
or U20880 (N_20880,N_19915,N_16907);
nor U20881 (N_20881,N_17065,N_18916);
nand U20882 (N_20882,N_16946,N_17836);
xnor U20883 (N_20883,N_18508,N_17420);
nand U20884 (N_20884,N_19559,N_17651);
nor U20885 (N_20885,N_19506,N_15229);
nor U20886 (N_20886,N_17696,N_18237);
and U20887 (N_20887,N_15824,N_16588);
xor U20888 (N_20888,N_15436,N_16306);
nand U20889 (N_20889,N_18960,N_19560);
and U20890 (N_20890,N_17428,N_16331);
and U20891 (N_20891,N_19582,N_15246);
or U20892 (N_20892,N_16327,N_18652);
nor U20893 (N_20893,N_19883,N_19634);
nor U20894 (N_20894,N_17426,N_16920);
or U20895 (N_20895,N_19248,N_19063);
nand U20896 (N_20896,N_17861,N_16338);
nand U20897 (N_20897,N_19364,N_19713);
nand U20898 (N_20898,N_15769,N_15632);
nand U20899 (N_20899,N_19120,N_19226);
xnor U20900 (N_20900,N_17749,N_18992);
nand U20901 (N_20901,N_16656,N_16309);
and U20902 (N_20902,N_15271,N_19921);
and U20903 (N_20903,N_15302,N_16388);
nand U20904 (N_20904,N_18122,N_15694);
and U20905 (N_20905,N_19362,N_17708);
or U20906 (N_20906,N_15106,N_15149);
nand U20907 (N_20907,N_16129,N_16654);
nand U20908 (N_20908,N_15445,N_15001);
nand U20909 (N_20909,N_18519,N_15916);
nor U20910 (N_20910,N_17561,N_17396);
xor U20911 (N_20911,N_19031,N_17488);
and U20912 (N_20912,N_16190,N_18209);
and U20913 (N_20913,N_16032,N_17889);
nor U20914 (N_20914,N_17545,N_15345);
and U20915 (N_20915,N_19633,N_18217);
and U20916 (N_20916,N_18081,N_17751);
or U20917 (N_20917,N_16347,N_18418);
nand U20918 (N_20918,N_16787,N_19483);
xnor U20919 (N_20919,N_16134,N_15930);
and U20920 (N_20920,N_16631,N_17123);
nand U20921 (N_20921,N_18945,N_15137);
or U20922 (N_20922,N_19888,N_19613);
and U20923 (N_20923,N_16079,N_16956);
xnor U20924 (N_20924,N_17182,N_16630);
or U20925 (N_20925,N_19201,N_16982);
or U20926 (N_20926,N_17179,N_16840);
nor U20927 (N_20927,N_19210,N_17352);
xor U20928 (N_20928,N_19936,N_15454);
xnor U20929 (N_20929,N_19232,N_19696);
or U20930 (N_20930,N_16928,N_16183);
and U20931 (N_20931,N_19984,N_19234);
nor U20932 (N_20932,N_15942,N_18906);
and U20933 (N_20933,N_17206,N_17925);
and U20934 (N_20934,N_19350,N_18268);
xnor U20935 (N_20935,N_16532,N_15982);
nor U20936 (N_20936,N_16780,N_16224);
and U20937 (N_20937,N_16705,N_17573);
nand U20938 (N_20938,N_17364,N_19840);
nand U20939 (N_20939,N_18496,N_16197);
or U20940 (N_20940,N_19319,N_18850);
xnor U20941 (N_20941,N_17446,N_16873);
xnor U20942 (N_20942,N_15705,N_17246);
xnor U20943 (N_20943,N_19075,N_15780);
and U20944 (N_20944,N_18434,N_17325);
or U20945 (N_20945,N_16691,N_16571);
nor U20946 (N_20946,N_16168,N_17001);
and U20947 (N_20947,N_15181,N_17165);
xor U20948 (N_20948,N_15513,N_16352);
and U20949 (N_20949,N_18740,N_15598);
nand U20950 (N_20950,N_16001,N_19484);
nor U20951 (N_20951,N_16726,N_16276);
or U20952 (N_20952,N_18043,N_19686);
and U20953 (N_20953,N_18637,N_16500);
or U20954 (N_20954,N_18073,N_16794);
xor U20955 (N_20955,N_19658,N_18087);
nand U20956 (N_20956,N_17808,N_19060);
xnor U20957 (N_20957,N_16999,N_16493);
or U20958 (N_20958,N_16604,N_18141);
nand U20959 (N_20959,N_15815,N_18229);
nor U20960 (N_20960,N_16886,N_17788);
xor U20961 (N_20961,N_16929,N_15263);
nor U20962 (N_20962,N_16455,N_15988);
xor U20963 (N_20963,N_15308,N_17666);
xnor U20964 (N_20964,N_19620,N_16499);
or U20965 (N_20965,N_16251,N_18419);
xor U20966 (N_20966,N_19112,N_19313);
and U20967 (N_20967,N_17117,N_17569);
nand U20968 (N_20968,N_17563,N_18976);
nand U20969 (N_20969,N_16265,N_17086);
nor U20970 (N_20970,N_19479,N_19778);
xor U20971 (N_20971,N_17564,N_19110);
xnor U20972 (N_20972,N_18904,N_16261);
or U20973 (N_20973,N_15094,N_17804);
nand U20974 (N_20974,N_16749,N_16422);
or U20975 (N_20975,N_16888,N_17480);
nor U20976 (N_20976,N_15946,N_18833);
nor U20977 (N_20977,N_18086,N_15153);
or U20978 (N_20978,N_15216,N_17731);
nor U20979 (N_20979,N_19734,N_18977);
or U20980 (N_20980,N_19279,N_15076);
nand U20981 (N_20981,N_17473,N_16674);
nor U20982 (N_20982,N_15602,N_15221);
and U20983 (N_20983,N_19079,N_18111);
and U20984 (N_20984,N_15894,N_19473);
xor U20985 (N_20985,N_18583,N_17932);
nor U20986 (N_20986,N_19940,N_17138);
nor U20987 (N_20987,N_19242,N_16091);
xor U20988 (N_20988,N_19418,N_16332);
xnor U20989 (N_20989,N_15979,N_16858);
and U20990 (N_20990,N_18520,N_15256);
xnor U20991 (N_20991,N_16413,N_15105);
xnor U20992 (N_20992,N_17551,N_19907);
nand U20993 (N_20993,N_17402,N_19134);
or U20994 (N_20994,N_19115,N_19086);
xor U20995 (N_20995,N_16488,N_15016);
xnor U20996 (N_20996,N_17985,N_19869);
or U20997 (N_20997,N_15965,N_17414);
xnor U20998 (N_20998,N_18533,N_16385);
xor U20999 (N_20999,N_15749,N_15052);
xnor U21000 (N_21000,N_16478,N_15716);
nand U21001 (N_21001,N_15841,N_17083);
and U21002 (N_21002,N_18100,N_15493);
and U21003 (N_21003,N_19647,N_16881);
and U21004 (N_21004,N_17694,N_19062);
nor U21005 (N_21005,N_17291,N_19356);
and U21006 (N_21006,N_19643,N_16531);
nand U21007 (N_21007,N_18649,N_19900);
nand U21008 (N_21008,N_19574,N_15609);
nand U21009 (N_21009,N_16779,N_16821);
nor U21010 (N_21010,N_16368,N_15630);
nor U21011 (N_21011,N_18452,N_18259);
nand U21012 (N_21012,N_19991,N_18988);
or U21013 (N_21013,N_19892,N_19139);
xnor U21014 (N_21014,N_16133,N_15651);
xnor U21015 (N_21015,N_18791,N_18630);
nand U21016 (N_21016,N_15124,N_18213);
xor U21017 (N_21017,N_15364,N_18867);
nand U21018 (N_21018,N_18855,N_17338);
nand U21019 (N_21019,N_17046,N_17824);
and U21020 (N_21020,N_17181,N_17278);
xor U21021 (N_21021,N_15718,N_15587);
or U21022 (N_21022,N_19579,N_15908);
nand U21023 (N_21023,N_16179,N_18196);
or U21024 (N_21024,N_17416,N_17513);
nand U21025 (N_21025,N_17323,N_18790);
or U21026 (N_21026,N_17363,N_17734);
nor U21027 (N_21027,N_19379,N_17566);
or U21028 (N_21028,N_19097,N_18927);
or U21029 (N_21029,N_15663,N_16935);
or U21030 (N_21030,N_15703,N_16993);
nor U21031 (N_21031,N_19622,N_17913);
nand U21032 (N_21032,N_18724,N_15045);
and U21033 (N_21033,N_15303,N_19312);
xor U21034 (N_21034,N_16576,N_19211);
xnor U21035 (N_21035,N_15112,N_18013);
and U21036 (N_21036,N_18428,N_17337);
nor U21037 (N_21037,N_19530,N_19444);
xnor U21038 (N_21038,N_16207,N_16953);
xnor U21039 (N_21039,N_18207,N_18421);
and U21040 (N_21040,N_19420,N_18447);
xor U21041 (N_21041,N_18351,N_16583);
nor U21042 (N_21042,N_17266,N_18680);
or U21043 (N_21043,N_16252,N_17534);
xnor U21044 (N_21044,N_15392,N_16947);
xnor U21045 (N_21045,N_16270,N_17670);
nor U21046 (N_21046,N_19923,N_18220);
xor U21047 (N_21047,N_17624,N_17532);
and U21048 (N_21048,N_16495,N_15664);
and U21049 (N_21049,N_17671,N_18517);
nor U21050 (N_21050,N_15119,N_17791);
and U21051 (N_21051,N_19554,N_15933);
and U21052 (N_21052,N_16214,N_17568);
nor U21053 (N_21053,N_16648,N_18993);
and U21054 (N_21054,N_17307,N_17864);
nor U21055 (N_21055,N_15189,N_18967);
nand U21056 (N_21056,N_17992,N_19591);
xor U21057 (N_21057,N_16662,N_18311);
and U21058 (N_21058,N_17965,N_19976);
nand U21059 (N_21059,N_19329,N_15898);
xnor U21060 (N_21060,N_15583,N_16539);
nor U21061 (N_21061,N_19855,N_18255);
or U21062 (N_21062,N_17800,N_15441);
and U21063 (N_21063,N_18438,N_16560);
xnor U21064 (N_21064,N_19121,N_18800);
nand U21065 (N_21065,N_19600,N_16547);
xor U21066 (N_21066,N_17881,N_19485);
nor U21067 (N_21067,N_19961,N_17268);
xor U21068 (N_21068,N_18877,N_15170);
nor U21069 (N_21069,N_19138,N_15797);
or U21070 (N_21070,N_17843,N_17466);
nand U21071 (N_21071,N_19712,N_18607);
xor U21072 (N_21072,N_17767,N_16095);
nand U21073 (N_21073,N_16605,N_15404);
nand U21074 (N_21074,N_16202,N_16476);
xnor U21075 (N_21075,N_15282,N_18731);
or U21076 (N_21076,N_19306,N_15268);
and U21077 (N_21077,N_16690,N_16884);
and U21078 (N_21078,N_19181,N_18538);
and U21079 (N_21079,N_17989,N_15584);
nor U21080 (N_21080,N_19597,N_18113);
nand U21081 (N_21081,N_18903,N_16263);
nor U21082 (N_21082,N_18948,N_15202);
nor U21083 (N_21083,N_18109,N_17036);
nand U21084 (N_21084,N_18605,N_18592);
nand U21085 (N_21085,N_15264,N_18234);
xnor U21086 (N_21086,N_17169,N_16522);
nor U21087 (N_21087,N_19190,N_17737);
xnor U21088 (N_21088,N_16970,N_19055);
nor U21089 (N_21089,N_19363,N_15362);
nand U21090 (N_21090,N_18396,N_15418);
nand U21091 (N_21091,N_19489,N_19074);
nand U21092 (N_21092,N_18188,N_16436);
or U21093 (N_21093,N_16087,N_17155);
nor U21094 (N_21094,N_17368,N_16919);
and U21095 (N_21095,N_19090,N_17638);
or U21096 (N_21096,N_16379,N_19499);
xnor U21097 (N_21097,N_16716,N_19970);
nor U21098 (N_21098,N_16320,N_16404);
nor U21099 (N_21099,N_19641,N_19084);
and U21100 (N_21100,N_15243,N_18126);
nor U21101 (N_21101,N_17003,N_15393);
nand U21102 (N_21102,N_15108,N_19057);
or U21103 (N_21103,N_19746,N_18065);
and U21104 (N_21104,N_16216,N_17852);
or U21105 (N_21105,N_18193,N_15339);
or U21106 (N_21106,N_15709,N_17183);
or U21107 (N_21107,N_16412,N_16863);
or U21108 (N_21108,N_16612,N_15561);
or U21109 (N_21109,N_18187,N_16528);
xnor U21110 (N_21110,N_17020,N_16299);
and U21111 (N_21111,N_16813,N_16957);
nand U21112 (N_21112,N_17865,N_19844);
nand U21113 (N_21113,N_19692,N_15304);
xnor U21114 (N_21114,N_15222,N_17226);
or U21115 (N_21115,N_16067,N_15646);
and U21116 (N_21116,N_19614,N_17339);
or U21117 (N_21117,N_19209,N_15142);
or U21118 (N_21118,N_16720,N_17654);
and U21119 (N_21119,N_16595,N_19804);
and U21120 (N_21120,N_18561,N_15966);
and U21121 (N_21121,N_15178,N_15987);
nand U21122 (N_21122,N_17684,N_17712);
or U21123 (N_21123,N_15509,N_17497);
xor U21124 (N_21124,N_17027,N_19290);
and U21125 (N_21125,N_17374,N_18889);
nand U21126 (N_21126,N_18203,N_15559);
nand U21127 (N_21127,N_17682,N_19272);
nor U21128 (N_21128,N_17723,N_19640);
or U21129 (N_21129,N_15827,N_15765);
and U21130 (N_21130,N_18423,N_16620);
and U21131 (N_21131,N_16078,N_17437);
xnor U21132 (N_21132,N_15361,N_16729);
nor U21133 (N_21133,N_15734,N_17930);
or U21134 (N_21134,N_17878,N_18898);
nor U21135 (N_21135,N_18215,N_16290);
nor U21136 (N_21136,N_15581,N_15154);
nor U21137 (N_21137,N_16479,N_18983);
nor U21138 (N_21138,N_16019,N_17320);
nand U21139 (N_21139,N_16292,N_18837);
nor U21140 (N_21140,N_15203,N_17474);
and U21141 (N_21141,N_16939,N_15326);
nand U21142 (N_21142,N_15919,N_18566);
xnor U21143 (N_21143,N_18420,N_16585);
nand U21144 (N_21144,N_15880,N_15395);
xnor U21145 (N_21145,N_19095,N_18107);
or U21146 (N_21146,N_18205,N_16025);
nand U21147 (N_21147,N_19805,N_18671);
or U21148 (N_21148,N_19137,N_18112);
xor U21149 (N_21149,N_15673,N_19264);
xor U21150 (N_21150,N_19191,N_19852);
nand U21151 (N_21151,N_16449,N_15158);
or U21152 (N_21152,N_16818,N_18151);
xor U21153 (N_21153,N_19781,N_15661);
xor U21154 (N_21154,N_17287,N_17366);
xor U21155 (N_21155,N_17194,N_16466);
nand U21156 (N_21156,N_19399,N_15327);
xnor U21157 (N_21157,N_16877,N_18061);
nor U21158 (N_21158,N_15335,N_18750);
or U21159 (N_21159,N_15236,N_15680);
and U21160 (N_21160,N_17006,N_19085);
or U21161 (N_21161,N_19355,N_17478);
xor U21162 (N_21162,N_19147,N_16259);
and U21163 (N_21163,N_17726,N_17917);
xnor U21164 (N_21164,N_16193,N_18644);
nor U21165 (N_21165,N_16051,N_16401);
and U21166 (N_21166,N_18402,N_16537);
nand U21167 (N_21167,N_17175,N_16472);
nor U21168 (N_21168,N_15883,N_17938);
xor U21169 (N_21169,N_15713,N_15565);
and U21170 (N_21170,N_18655,N_18222);
and U21171 (N_21171,N_18539,N_19037);
nor U21172 (N_21172,N_17867,N_15791);
and U21173 (N_21173,N_15328,N_17345);
and U21174 (N_21174,N_19229,N_16707);
or U21175 (N_21175,N_18437,N_15684);
or U21176 (N_21176,N_16525,N_17040);
xor U21177 (N_21177,N_18041,N_15423);
xnor U21178 (N_21178,N_19749,N_19006);
nor U21179 (N_21179,N_18378,N_15248);
nand U21180 (N_21180,N_17190,N_18269);
and U21181 (N_21181,N_19497,N_19627);
nor U21182 (N_21182,N_17431,N_17265);
xor U21183 (N_21183,N_16847,N_19253);
nor U21184 (N_21184,N_17253,N_18819);
and U21185 (N_21185,N_17606,N_16567);
or U21186 (N_21186,N_17860,N_16425);
and U21187 (N_21187,N_17623,N_16210);
and U21188 (N_21188,N_16508,N_18688);
or U21189 (N_21189,N_19308,N_15656);
and U21190 (N_21190,N_19969,N_17698);
and U21191 (N_21191,N_19361,N_15702);
nand U21192 (N_21192,N_15752,N_19231);
nor U21193 (N_21193,N_18290,N_16972);
xnor U21194 (N_21194,N_17900,N_17807);
and U21195 (N_21195,N_17614,N_15562);
xor U21196 (N_21196,N_15483,N_16017);
or U21197 (N_21197,N_16416,N_17691);
nor U21198 (N_21198,N_19394,N_15499);
or U21199 (N_21199,N_15323,N_18795);
xnor U21200 (N_21200,N_18792,N_16021);
nand U21201 (N_21201,N_18356,N_15198);
and U21202 (N_21202,N_18689,N_17986);
xor U21203 (N_21203,N_18006,N_18679);
and U21204 (N_21204,N_17145,N_19513);
nand U21205 (N_21205,N_19963,N_15510);
and U21206 (N_21206,N_16520,N_16098);
and U21207 (N_21207,N_18686,N_17503);
xor U21208 (N_21208,N_19901,N_16328);
nand U21209 (N_21209,N_15999,N_18353);
nand U21210 (N_21210,N_15787,N_18360);
and U21211 (N_21211,N_16342,N_16253);
and U21212 (N_21212,N_19149,N_18383);
xor U21213 (N_21213,N_18755,N_16198);
and U21214 (N_21214,N_17490,N_18617);
xor U21215 (N_21215,N_16703,N_18776);
and U21216 (N_21216,N_16711,N_19540);
nand U21217 (N_21217,N_18532,N_16553);
and U21218 (N_21218,N_18136,N_17757);
and U21219 (N_21219,N_19521,N_17973);
xor U21220 (N_21220,N_19639,N_19044);
nor U21221 (N_21221,N_18076,N_19334);
nand U21222 (N_21222,N_19660,N_16022);
nor U21223 (N_21223,N_15116,N_17676);
and U21224 (N_21224,N_18569,N_17591);
nand U21225 (N_21225,N_17763,N_15924);
or U21226 (N_21226,N_18982,N_16673);
and U21227 (N_21227,N_19617,N_19950);
and U21228 (N_21228,N_15133,N_15720);
nor U21229 (N_21229,N_17264,N_17799);
nor U21230 (N_21230,N_19811,N_17897);
nand U21231 (N_21231,N_15487,N_18788);
or U21232 (N_21232,N_18224,N_19831);
nand U21233 (N_21233,N_19007,N_19856);
or U21234 (N_21234,N_19013,N_18718);
or U21235 (N_21235,N_15638,N_15794);
nor U21236 (N_21236,N_18918,N_17360);
nand U21237 (N_21237,N_19100,N_15057);
and U21238 (N_21238,N_15293,N_17059);
nand U21239 (N_21239,N_15940,N_17216);
nor U21240 (N_21240,N_17597,N_17154);
nor U21241 (N_21241,N_17970,N_15200);
or U21242 (N_21242,N_15763,N_17610);
nor U21243 (N_21243,N_19073,N_17251);
xor U21244 (N_21244,N_17585,N_17890);
xor U21245 (N_21245,N_19721,N_16944);
nand U21246 (N_21246,N_17274,N_15085);
or U21247 (N_21247,N_15459,N_18696);
xnor U21248 (N_21248,N_16958,N_17130);
or U21249 (N_21249,N_16487,N_17840);
or U21250 (N_21250,N_17873,N_17987);
or U21251 (N_21251,N_18243,N_18505);
nand U21252 (N_21252,N_17646,N_15738);
xor U21253 (N_21253,N_16851,N_19524);
nor U21254 (N_21254,N_16409,N_19652);
xnor U21255 (N_21255,N_17538,N_16086);
nand U21256 (N_21256,N_16728,N_15039);
xnor U21257 (N_21257,N_19238,N_16159);
xor U21258 (N_21258,N_18687,N_16506);
or U21259 (N_21259,N_18535,N_18729);
nand U21260 (N_21260,N_15522,N_15277);
or U21261 (N_21261,N_18381,N_15146);
and U21262 (N_21262,N_19601,N_15870);
nand U21263 (N_21263,N_19157,N_15151);
nor U21264 (N_21264,N_17996,N_16489);
or U21265 (N_21265,N_15428,N_18206);
nor U21266 (N_21266,N_15516,N_15425);
or U21267 (N_21267,N_16346,N_19457);
nand U21268 (N_21268,N_18368,N_18758);
xnor U21269 (N_21269,N_15622,N_15699);
or U21270 (N_21270,N_19281,N_16582);
xnor U21271 (N_21271,N_16117,N_15869);
nand U21272 (N_21272,N_19241,N_15288);
or U21273 (N_21273,N_16850,N_16181);
nand U21274 (N_21274,N_17816,N_18247);
nand U21275 (N_21275,N_15756,N_16318);
and U21276 (N_21276,N_17826,N_15537);
nor U21277 (N_21277,N_16367,N_15936);
nor U21278 (N_21278,N_18772,N_15724);
nand U21279 (N_21279,N_16376,N_15891);
nand U21280 (N_21280,N_15920,N_18610);
and U21281 (N_21281,N_19878,N_15546);
and U21282 (N_21282,N_19993,N_17908);
nor U21283 (N_21283,N_15071,N_15931);
xnor U21284 (N_21284,N_15100,N_19931);
and U21285 (N_21285,N_17524,N_16524);
or U21286 (N_21286,N_15034,N_18646);
nand U21287 (N_21287,N_18019,N_17945);
nor U21288 (N_21288,N_17289,N_19186);
and U21289 (N_21289,N_16066,N_16501);
and U21290 (N_21290,N_15152,N_15858);
or U21291 (N_21291,N_19236,N_18994);
nand U21292 (N_21292,N_15795,N_16527);
xnor U21293 (N_21293,N_17296,N_15913);
or U21294 (N_21294,N_17180,N_16649);
or U21295 (N_21295,N_19142,N_19284);
nand U21296 (N_21296,N_18327,N_17050);
nand U21297 (N_21297,N_18928,N_18108);
and U21298 (N_21298,N_18694,N_15072);
nand U21299 (N_21299,N_19146,N_15365);
and U21300 (N_21300,N_19948,N_17988);
xnor U21301 (N_21301,N_18673,N_19797);
nor U21302 (N_21302,N_17148,N_17098);
or U21303 (N_21303,N_18009,N_18879);
nor U21304 (N_21304,N_16018,N_17135);
xor U21305 (N_21305,N_15772,N_18595);
xnor U21306 (N_21306,N_15834,N_19927);
and U21307 (N_21307,N_18282,N_15868);
xor U21308 (N_21308,N_16627,N_15272);
nor U21309 (N_21309,N_19910,N_15796);
nand U21310 (N_21310,N_19207,N_17140);
or U21311 (N_21311,N_15352,N_18280);
or U21312 (N_21312,N_19288,N_19884);
nor U21313 (N_21313,N_18865,N_17144);
nor U21314 (N_21314,N_19874,N_15187);
or U21315 (N_21315,N_18484,N_18165);
or U21316 (N_21316,N_16312,N_17031);
xor U21317 (N_21317,N_15012,N_17283);
or U21318 (N_21318,N_18812,N_15250);
and U21319 (N_21319,N_15654,N_16351);
xnor U21320 (N_21320,N_16883,N_15697);
nor U21321 (N_21321,N_16828,N_18764);
and U21322 (N_21322,N_18573,N_19981);
or U21323 (N_21323,N_18924,N_17998);
nand U21324 (N_21324,N_17656,N_16676);
xor U21325 (N_21325,N_17102,N_15038);
nor U21326 (N_21326,N_19619,N_16747);
and U21327 (N_21327,N_17223,N_17217);
and U21328 (N_21328,N_16496,N_15995);
nand U21329 (N_21329,N_16326,N_17812);
nor U21330 (N_21330,N_19064,N_17469);
xnor U21331 (N_21331,N_19411,N_15473);
and U21332 (N_21332,N_18411,N_17649);
or U21333 (N_21333,N_16383,N_15475);
or U21334 (N_21334,N_16611,N_15047);
nor U21335 (N_21335,N_15555,N_18944);
xor U21336 (N_21336,N_18202,N_19425);
nand U21337 (N_21337,N_19198,N_17904);
nor U21338 (N_21338,N_19469,N_19316);
nand U21339 (N_21339,N_15141,N_16763);
nor U21340 (N_21340,N_15051,N_18439);
or U21341 (N_21341,N_15593,N_16983);
nand U21342 (N_21342,N_16686,N_17215);
nand U21343 (N_21343,N_19072,N_16061);
or U21344 (N_21344,N_19853,N_16742);
and U21345 (N_21345,N_19584,N_15885);
and U21346 (N_21346,N_19375,N_17128);
xnor U21347 (N_21347,N_17022,N_15015);
nand U21348 (N_21348,N_15079,N_15385);
nand U21349 (N_21349,N_16284,N_17214);
and U21350 (N_21350,N_15594,N_15409);
nor U21351 (N_21351,N_19762,N_17922);
nand U21352 (N_21352,N_16212,N_18784);
nor U21353 (N_21353,N_16016,N_16688);
or U21354 (N_21354,N_18293,N_15662);
nor U21355 (N_21355,N_16770,N_15388);
or U21356 (N_21356,N_17026,N_16721);
nand U21357 (N_21357,N_15665,N_17010);
nand U21358 (N_21358,N_16483,N_16195);
or U21359 (N_21359,N_16109,N_16257);
xnor U21360 (N_21360,N_18959,N_15669);
or U21361 (N_21361,N_18049,N_16447);
or U21362 (N_21362,N_16917,N_18459);
and U21363 (N_21363,N_18475,N_15291);
nor U21364 (N_21364,N_16206,N_15060);
nand U21365 (N_21365,N_18120,N_19237);
or U21366 (N_21366,N_18820,N_15861);
and U21367 (N_21367,N_19939,N_16474);
nor U21368 (N_21368,N_16302,N_15334);
xor U21369 (N_21369,N_16044,N_17504);
xor U21370 (N_21370,N_17579,N_15095);
and U21371 (N_21371,N_15314,N_18026);
or U21372 (N_21372,N_19972,N_16002);
nor U21373 (N_21373,N_18331,N_19435);
nand U21374 (N_21374,N_19414,N_16267);
or U21375 (N_21375,N_16823,N_18030);
nor U21376 (N_21376,N_16064,N_16096);
or U21377 (N_21377,N_15023,N_17034);
nand U21378 (N_21378,N_18332,N_19098);
nor U21379 (N_21379,N_19380,N_19464);
nor U21380 (N_21380,N_16530,N_15682);
nor U21381 (N_21381,N_17030,N_17803);
or U21382 (N_21382,N_18373,N_16637);
nor U21383 (N_21383,N_18632,N_19358);
and U21384 (N_21384,N_16569,N_17393);
nand U21385 (N_21385,N_16240,N_17634);
or U21386 (N_21386,N_15990,N_17615);
nand U21387 (N_21387,N_18684,N_15693);
or U21388 (N_21388,N_15659,N_18291);
nand U21389 (N_21389,N_19556,N_18492);
xor U21390 (N_21390,N_16857,N_16790);
and U21391 (N_21391,N_15912,N_18711);
nor U21392 (N_21392,N_18458,N_19304);
nand U21393 (N_21393,N_16997,N_19136);
nand U21394 (N_21394,N_18422,N_15294);
nand U21395 (N_21395,N_19680,N_17170);
nand U21396 (N_21396,N_17185,N_18465);
or U21397 (N_21397,N_15619,N_19130);
nor U21398 (N_21398,N_18690,N_16377);
nor U21399 (N_21399,N_17562,N_19566);
nand U21400 (N_21400,N_18661,N_15099);
nand U21401 (N_21401,N_17526,N_17773);
and U21402 (N_21402,N_16192,N_17918);
nor U21403 (N_21403,N_19621,N_18986);
nor U21404 (N_21404,N_18106,N_18547);
and U21405 (N_21405,N_18766,N_17070);
xor U21406 (N_21406,N_15785,N_15783);
nand U21407 (N_21407,N_16842,N_16551);
nand U21408 (N_21408,N_17272,N_16943);
nand U21409 (N_21409,N_19458,N_16761);
xor U21410 (N_21410,N_17655,N_15747);
or U21411 (N_21411,N_17547,N_19328);
nor U21412 (N_21412,N_19798,N_15226);
or U21413 (N_21413,N_19038,N_18441);
nand U21414 (N_21414,N_18083,N_19790);
xnor U21415 (N_21415,N_17999,N_19924);
nor U21416 (N_21416,N_17476,N_17224);
and U21417 (N_21417,N_15778,N_18809);
nand U21418 (N_21418,N_17997,N_19638);
or U21419 (N_21419,N_15315,N_15180);
nor U21420 (N_21420,N_19148,N_15541);
xnor U21421 (N_21421,N_17095,N_16979);
and U21422 (N_21422,N_17502,N_15128);
xor U21423 (N_21423,N_16381,N_16966);
nor U21424 (N_21424,N_18909,N_17475);
and U21425 (N_21425,N_16461,N_19818);
or U21426 (N_21426,N_15745,N_18542);
or U21427 (N_21427,N_15881,N_18778);
xnor U21428 (N_21428,N_16556,N_18575);
or U21429 (N_21429,N_18300,N_19395);
or U21430 (N_21430,N_19876,N_15349);
xnor U21431 (N_21431,N_16027,N_16186);
xnor U21432 (N_21432,N_17729,N_18503);
nand U21433 (N_21433,N_19269,N_19332);
or U21434 (N_21434,N_18191,N_16364);
xnor U21435 (N_21435,N_17857,N_19410);
or U21436 (N_21436,N_19096,N_19070);
or U21437 (N_21437,N_17453,N_16170);
nor U21438 (N_21438,N_17661,N_17821);
or U21439 (N_21439,N_17571,N_17304);
nor U21440 (N_21440,N_16076,N_17962);
or U21441 (N_21441,N_18480,N_18836);
nor U21442 (N_21442,N_19263,N_15655);
and U21443 (N_21443,N_16242,N_16772);
nand U21444 (N_21444,N_19787,N_19920);
nand U21445 (N_21445,N_15865,N_16132);
nand U21446 (N_21446,N_16174,N_15322);
xnor U21447 (N_21447,N_17487,N_16482);
and U21448 (N_21448,N_16282,N_17037);
or U21449 (N_21449,N_18609,N_19782);
nor U21450 (N_21450,N_19854,N_18734);
and U21451 (N_21451,N_17692,N_15953);
and U21452 (N_21452,N_15390,N_17903);
nand U21453 (N_21453,N_15089,N_19326);
xor U21454 (N_21454,N_18929,N_18530);
and U21455 (N_21455,N_19827,N_15657);
nand U21456 (N_21456,N_19978,N_17829);
and U21457 (N_21457,N_18101,N_16523);
or U21458 (N_21458,N_19474,N_18374);
nand U21459 (N_21459,N_15123,N_16188);
xor U21460 (N_21460,N_16149,N_17884);
or U21461 (N_21461,N_17554,N_15589);
and U21462 (N_21462,N_15580,N_17957);
xnor U21463 (N_21463,N_18634,N_17241);
and U21464 (N_21464,N_18338,N_15068);
nor U21465 (N_21465,N_19891,N_18717);
and U21466 (N_21466,N_17721,N_16286);
xor U21467 (N_21467,N_15711,N_19305);
nand U21468 (N_21468,N_17909,N_18038);
nand U21469 (N_21469,N_18899,N_18797);
xor U21470 (N_21470,N_17540,N_18970);
or U21471 (N_21471,N_15318,N_17498);
nand U21472 (N_21472,N_15201,N_18822);
xor U21473 (N_21473,N_16852,N_19544);
or U21474 (N_21474,N_17866,N_17069);
or U21475 (N_21475,N_16597,N_16271);
nand U21476 (N_21476,N_19741,N_18340);
and U21477 (N_21477,N_17405,N_15372);
xnor U21478 (N_21478,N_16199,N_19918);
or U21479 (N_21479,N_16249,N_19842);
nand U21480 (N_21480,N_16231,N_15290);
nor U21481 (N_21481,N_16144,N_17931);
nand U21482 (N_21482,N_15520,N_18297);
nor U21483 (N_21483,N_18658,N_17324);
nor U21484 (N_21484,N_16266,N_16442);
xor U21485 (N_21485,N_18494,N_15218);
and U21486 (N_21486,N_15922,N_17139);
or U21487 (N_21487,N_19731,N_16492);
nand U21488 (N_21488,N_15083,N_15311);
or U21489 (N_21489,N_15376,N_16514);
and U21490 (N_21490,N_19670,N_15949);
nor U21491 (N_21491,N_18075,N_17118);
and U21492 (N_21492,N_17231,N_16733);
nor U21493 (N_21493,N_16399,N_15554);
xor U21494 (N_21494,N_18042,N_17298);
xnor U21495 (N_21495,N_18181,N_19966);
or U21496 (N_21496,N_16786,N_15161);
nor U21497 (N_21497,N_17978,N_17736);
xor U21498 (N_21498,N_19099,N_18210);
and U21499 (N_21499,N_19776,N_15476);
nand U21500 (N_21500,N_18911,N_15526);
xnor U21501 (N_21501,N_17608,N_16209);
nand U21502 (N_21502,N_17923,N_15371);
xor U21503 (N_21503,N_19512,N_19751);
nor U21504 (N_21504,N_19968,N_19902);
nand U21505 (N_21505,N_17934,N_16039);
nand U21506 (N_21506,N_16083,N_15722);
or U21507 (N_21507,N_18488,N_16965);
nor U21508 (N_21508,N_16869,N_17747);
or U21509 (N_21509,N_19454,N_19429);
nand U21510 (N_21510,N_16237,N_17575);
and U21511 (N_21511,N_15342,N_17444);
or U21512 (N_21512,N_19260,N_17939);
xor U21513 (N_21513,N_19081,N_15884);
and U21514 (N_21514,N_19267,N_16866);
nand U21515 (N_21515,N_15810,N_17159);
or U21516 (N_21516,N_16860,N_19089);
xnor U21517 (N_21517,N_18886,N_16902);
nor U21518 (N_21518,N_15230,N_16041);
and U21519 (N_21519,N_15467,N_17733);
or U21520 (N_21520,N_15963,N_19881);
nand U21521 (N_21521,N_15943,N_17717);
nor U21522 (N_21522,N_18047,N_16316);
and U21523 (N_21523,N_18099,N_18365);
or U21524 (N_21524,N_15811,N_15464);
nand U21525 (N_21525,N_16901,N_18667);
and U21526 (N_21526,N_16153,N_16314);
and U21527 (N_21527,N_17449,N_15179);
xnor U21528 (N_21528,N_18092,N_17797);
nand U21529 (N_21529,N_15444,N_17678);
xor U21530 (N_21530,N_17711,N_15874);
nand U21531 (N_21531,N_18995,N_17844);
or U21532 (N_21532,N_17754,N_16426);
xor U21533 (N_21533,N_19796,N_16343);
nand U21534 (N_21534,N_17333,N_19527);
nor U21535 (N_21535,N_16330,N_19021);
and U21536 (N_21536,N_16748,N_19565);
nor U21537 (N_21537,N_18813,N_18023);
nand U21538 (N_21538,N_15086,N_15875);
or U21539 (N_21539,N_16760,N_18624);
nand U21540 (N_21540,N_19836,N_16692);
or U21541 (N_21541,N_16307,N_15830);
and U21542 (N_21542,N_15191,N_17874);
nand U21543 (N_21543,N_19179,N_17109);
xor U21544 (N_21544,N_19904,N_15244);
nand U21545 (N_21545,N_16550,N_18761);
or U21546 (N_21546,N_15194,N_16651);
nand U21547 (N_21547,N_19494,N_15289);
and U21548 (N_21548,N_16230,N_17794);
nor U21549 (N_21549,N_17845,N_15814);
xor U21550 (N_21550,N_17088,N_16548);
nand U21551 (N_21551,N_18266,N_16900);
or U21552 (N_21552,N_17501,N_19048);
nand U21553 (N_21553,N_19664,N_17584);
xnor U21554 (N_21554,N_17982,N_17613);
xnor U21555 (N_21555,N_15923,N_18681);
or U21556 (N_21556,N_17196,N_15871);
or U21557 (N_21557,N_16099,N_17326);
or U21558 (N_21558,N_16634,N_19893);
xnor U21559 (N_21559,N_16563,N_19922);
nand U21560 (N_21560,N_17641,N_18676);
or U21561 (N_21561,N_18129,N_15025);
and U21562 (N_21562,N_17367,N_16635);
xor U21563 (N_21563,N_16809,N_18854);
xnor U21564 (N_21564,N_15974,N_17929);
or U21565 (N_21565,N_19912,N_16962);
and U21566 (N_21566,N_15533,N_19051);
or U21567 (N_21567,N_15540,N_17543);
nand U21568 (N_21568,N_15370,N_15667);
xor U21569 (N_21569,N_17132,N_15719);
xnor U21570 (N_21570,N_18091,N_18656);
or U21571 (N_21571,N_15209,N_16088);
or U21572 (N_21572,N_19140,N_16354);
nand U21573 (N_21573,N_18145,N_17673);
nor U21574 (N_21574,N_17146,N_15599);
or U21575 (N_21575,N_16872,N_19944);
or U21576 (N_21576,N_18544,N_16991);
nand U21577 (N_21577,N_15255,N_15136);
or U21578 (N_21578,N_15970,N_17318);
xor U21579 (N_21579,N_16973,N_19557);
xnor U21580 (N_21580,N_16154,N_19646);
nand U21581 (N_21581,N_17868,N_18709);
or U21582 (N_21582,N_15551,N_16280);
xnor U21583 (N_21583,N_18808,N_19360);
xnor U21584 (N_21584,N_19462,N_18093);
nor U21585 (N_21585,N_15914,N_16296);
nand U21586 (N_21586,N_18163,N_18128);
and U21587 (N_21587,N_15696,N_15408);
nor U21588 (N_21588,N_15801,N_19520);
nand U21589 (N_21589,N_19233,N_16853);
xor U21590 (N_21590,N_19532,N_16395);
and U21591 (N_21591,N_18550,N_18597);
nor U21592 (N_21592,N_19247,N_19111);
nand U21593 (N_21593,N_18233,N_17252);
nand U21594 (N_21594,N_18635,N_16441);
xor U21595 (N_21595,N_16107,N_17434);
nor U21596 (N_21596,N_15131,N_17381);
nor U21597 (N_21597,N_18277,N_17213);
nand U21598 (N_21598,N_16867,N_17164);
or U21599 (N_21599,N_15007,N_16698);
and U21600 (N_21600,N_17427,N_15281);
nand U21601 (N_21601,N_18140,N_19626);
xnor U21602 (N_21602,N_17017,N_15983);
and U21603 (N_21603,N_19999,N_18748);
xor U21604 (N_21604,N_18828,N_19389);
nor U21605 (N_21605,N_16164,N_19135);
nand U21606 (N_21606,N_17395,N_19170);
nor U21607 (N_21607,N_16606,N_16610);
and U21608 (N_21608,N_18371,N_18551);
xor U21609 (N_21609,N_15650,N_17507);
nand U21610 (N_21610,N_18522,N_18150);
nand U21611 (N_21611,N_15676,N_16643);
nand U21612 (N_21612,N_18380,N_15821);
nor U21613 (N_21613,N_15253,N_15708);
or U21614 (N_21614,N_17893,N_17384);
or U21615 (N_21615,N_18745,N_15895);
xnor U21616 (N_21616,N_15944,N_18501);
nand U21617 (N_21617,N_17410,N_18008);
nor U21618 (N_21618,N_16115,N_17946);
nand U21619 (N_21619,N_18862,N_16052);
nand U21620 (N_21620,N_18352,N_19985);
and U21621 (N_21621,N_19807,N_18345);
nor U21622 (N_21622,N_16646,N_19548);
and U21623 (N_21623,N_17588,N_18117);
nand U21624 (N_21624,N_17300,N_19864);
nand U21625 (N_21625,N_17230,N_17512);
and U21626 (N_21626,N_19515,N_15286);
and U21627 (N_21627,N_16059,N_16980);
and U21628 (N_21628,N_18017,N_18826);
nor U21629 (N_21629,N_16655,N_17862);
or U21630 (N_21630,N_18240,N_19861);
xor U21631 (N_21631,N_16573,N_15558);
xor U21632 (N_21632,N_15517,N_15671);
nand U21633 (N_21633,N_15402,N_18811);
and U21634 (N_21634,N_18622,N_18334);
nor U21635 (N_21635,N_15539,N_18154);
nand U21636 (N_21636,N_16590,N_16048);
or U21637 (N_21637,N_18432,N_16056);
and U21638 (N_21638,N_15531,N_16068);
or U21639 (N_21639,N_16081,N_16552);
or U21640 (N_21640,N_18386,N_15907);
nand U21641 (N_21641,N_19406,N_18482);
and U21642 (N_21642,N_18782,N_18939);
or U21643 (N_21643,N_15893,N_18880);
nand U21644 (N_21644,N_15212,N_16152);
nor U21645 (N_21645,N_17879,N_16110);
and U21646 (N_21646,N_19913,N_16443);
and U21647 (N_21647,N_15391,N_17435);
and U21648 (N_21648,N_16723,N_18054);
xor U21649 (N_21649,N_15701,N_19889);
or U21650 (N_21650,N_19286,N_17359);
nand U21651 (N_21651,N_18872,N_16008);
nand U21652 (N_21652,N_19354,N_19171);
or U21653 (N_21653,N_17645,N_19102);
nor U21654 (N_21654,N_17424,N_17888);
or U21655 (N_21655,N_18350,N_15043);
and U21656 (N_21656,N_16625,N_18647);
nand U21657 (N_21657,N_19727,N_16895);
nor U21658 (N_21658,N_18683,N_16093);
xnor U21659 (N_21659,N_17162,N_17933);
xor U21660 (N_21660,N_15107,N_15495);
and U21661 (N_21661,N_18218,N_15232);
nand U21662 (N_21662,N_16647,N_15690);
or U21663 (N_21663,N_16337,N_17005);
and U21664 (N_21664,N_16305,N_17317);
xor U21665 (N_21665,N_18103,N_19477);
nor U21666 (N_21666,N_15896,N_17467);
nor U21667 (N_21667,N_18693,N_15299);
and U21668 (N_21668,N_18700,N_15296);
or U21669 (N_21669,N_19156,N_19705);
xor U21670 (N_21670,N_18753,N_17301);
and U21671 (N_21671,N_17688,N_18298);
xnor U21672 (N_21672,N_17883,N_18491);
and U21673 (N_21673,N_16744,N_15672);
nand U21674 (N_21674,N_16734,N_19982);
or U21675 (N_21675,N_18839,N_18453);
nor U21676 (N_21676,N_19691,N_19748);
or U21677 (N_21677,N_19028,N_17032);
xnor U21678 (N_21678,N_16882,N_18022);
and U21679 (N_21679,N_15355,N_19763);
and U21680 (N_21680,N_19180,N_15396);
xnor U21681 (N_21681,N_18251,N_15899);
nand U21682 (N_21682,N_18426,N_17137);
xor U21683 (N_21683,N_18257,N_17362);
nor U21684 (N_21684,N_15414,N_17407);
nand U21685 (N_21685,N_15616,N_19317);
xor U21686 (N_21686,N_17789,N_16457);
nand U21687 (N_21687,N_15195,N_16834);
xor U21688 (N_21688,N_17921,N_19422);
nand U21689 (N_21689,N_19154,N_18816);
and U21690 (N_21690,N_19453,N_17714);
xnor U21691 (N_21691,N_19522,N_19438);
nor U21692 (N_21692,N_19016,N_15491);
or U21693 (N_21693,N_18052,N_16890);
nor U21694 (N_21694,N_15033,N_17806);
and U21695 (N_21695,N_18253,N_18952);
nor U21696 (N_21696,N_18225,N_18449);
xor U21697 (N_21697,N_17830,N_18643);
and U21698 (N_21698,N_15578,N_15037);
nand U21699 (N_21699,N_16841,N_17741);
xnor U21700 (N_21700,N_18801,N_19068);
nand U21701 (N_21701,N_16400,N_18183);
or U21702 (N_21702,N_18973,N_18861);
or U21703 (N_21703,N_17556,N_15511);
or U21704 (N_21704,N_19398,N_15939);
xnor U21705 (N_21705,N_15452,N_18166);
xnor U21706 (N_21706,N_16058,N_17679);
and U21707 (N_21707,N_17619,N_18571);
nor U21708 (N_21708,N_15009,N_18949);
or U21709 (N_21709,N_17016,N_19259);
xor U21710 (N_21710,N_17716,N_17764);
xor U21711 (N_21711,N_18148,N_17518);
and U21712 (N_21712,N_15768,N_16215);
nor U21713 (N_21713,N_17486,N_18425);
nand U21714 (N_21714,N_15938,N_18200);
nor U21715 (N_21715,N_16536,N_18258);
or U21716 (N_21716,N_15478,N_18144);
nand U21717 (N_21717,N_16544,N_15762);
nor U21718 (N_21718,N_17357,N_19938);
or U21719 (N_21719,N_15295,N_16880);
nand U21720 (N_21720,N_19053,N_18611);
and U21721 (N_21721,N_18127,N_17618);
xor U21722 (N_21722,N_18309,N_17267);
xnor U21723 (N_21723,N_18773,N_16521);
nand U21724 (N_21724,N_19525,N_15443);
and U21725 (N_21725,N_15013,N_18614);
nor U21726 (N_21726,N_15652,N_17081);
xnor U21727 (N_21727,N_19770,N_17029);
nor U21728 (N_21728,N_19104,N_16679);
xor U21729 (N_21729,N_18296,N_17450);
xor U21730 (N_21730,N_17290,N_19995);
xor U21731 (N_21731,N_18468,N_16020);
or U21732 (N_21732,N_17042,N_16931);
nor U21733 (N_21733,N_17522,N_18463);
xor U21734 (N_21734,N_19487,N_16245);
or U21735 (N_21735,N_19400,N_19336);
xnor U21736 (N_21736,N_19760,N_18249);
xnor U21737 (N_21737,N_18153,N_15130);
or U21738 (N_21738,N_17971,N_18158);
or U21739 (N_21739,N_15590,N_19871);
and U21740 (N_21740,N_16854,N_19822);
nand U21741 (N_21741,N_17191,N_16219);
or U21742 (N_21742,N_17227,N_16236);
and U21743 (N_21743,N_17548,N_19806);
and U21744 (N_21744,N_15753,N_16765);
nand U21745 (N_21745,N_19998,N_15451);
xor U21746 (N_21746,N_18754,N_17898);
nand U21747 (N_21747,N_17330,N_17111);
nand U21748 (N_21748,N_17710,N_16574);
nor U21749 (N_21749,N_17441,N_15525);
or U21750 (N_21750,N_16062,N_17377);
xnor U21751 (N_21751,N_17404,N_17940);
nor U21752 (N_21752,N_19047,N_17234);
nand U21753 (N_21753,N_18914,N_18323);
xor U21754 (N_21754,N_18965,N_18055);
or U21755 (N_21755,N_19193,N_15528);
or U21756 (N_21756,N_17342,N_18926);
nand U21757 (N_21757,N_19225,N_15155);
nor U21758 (N_21758,N_17750,N_19581);
xor U21759 (N_21759,N_17142,N_17284);
nor U21760 (N_21760,N_16727,N_17786);
nand U21761 (N_21761,N_16363,N_16033);
or U21762 (N_21762,N_15267,N_16244);
or U21763 (N_21763,N_18246,N_19167);
and U21764 (N_21764,N_15143,N_18825);
xor U21765 (N_21765,N_16222,N_18265);
xor U21766 (N_21766,N_19108,N_18303);
nor U21767 (N_21767,N_19431,N_19133);
xnor U21768 (N_21768,N_18031,N_16405);
nand U21769 (N_21769,N_17297,N_18211);
nand U21770 (N_21770,N_15490,N_19197);
nand U21771 (N_21771,N_16871,N_18440);
nor U21772 (N_21772,N_16753,N_17875);
xnor U21773 (N_21773,N_18397,N_16255);
nand U21774 (N_21774,N_18769,N_19667);
xor U21775 (N_21775,N_15274,N_15823);
and U21776 (N_21776,N_18509,N_16120);
xor U21777 (N_21777,N_15027,N_18953);
and U21778 (N_21778,N_15958,N_16796);
xor U21779 (N_21779,N_18875,N_19091);
or U21780 (N_21780,N_17293,N_17667);
or U21781 (N_21781,N_15058,N_18934);
nand U21782 (N_21782,N_18619,N_16894);
nand U21783 (N_21783,N_15832,N_16954);
nand U21784 (N_21784,N_16812,N_17744);
and U21785 (N_21785,N_16030,N_19987);
or U21786 (N_21786,N_16355,N_15471);
xor U21787 (N_21787,N_17067,N_19523);
xor U21788 (N_21788,N_17334,N_19302);
or U21789 (N_21789,N_15167,N_16738);
and U21790 (N_21790,N_18589,N_16507);
and U21791 (N_21791,N_15492,N_16112);
and U21792 (N_21792,N_16746,N_16451);
nor U21793 (N_21793,N_15301,N_17386);
or U21794 (N_21794,N_17147,N_16896);
nor U21795 (N_21795,N_17823,N_16293);
or U21796 (N_21796,N_18034,N_18641);
xnor U21797 (N_21797,N_15518,N_16301);
or U21798 (N_21798,N_18214,N_15585);
nor U21799 (N_21799,N_15427,N_17520);
and U21800 (N_21800,N_19415,N_18130);
or U21801 (N_21801,N_19446,N_18167);
and U21802 (N_21802,N_19625,N_19671);
nor U21803 (N_21803,N_19475,N_17292);
xnor U21804 (N_21804,N_16268,N_16125);
nand U21805 (N_21805,N_17709,N_18759);
xor U21806 (N_21806,N_17953,N_17718);
and U21807 (N_21807,N_15803,N_19344);
or U21808 (N_21808,N_15486,N_17400);
xnor U21809 (N_21809,N_19323,N_18863);
nor U21810 (N_21810,N_16558,N_15429);
and U21811 (N_21811,N_19109,N_16791);
xor U21812 (N_21812,N_15956,N_19199);
nor U21813 (N_21813,N_15185,N_18727);
nor U21814 (N_21814,N_16118,N_16345);
and U21815 (N_21815,N_18885,N_16913);
nor U21816 (N_21816,N_15144,N_18726);
xnor U21817 (N_21817,N_15854,N_18455);
xnor U21818 (N_21818,N_18757,N_15064);
and U21819 (N_21819,N_19943,N_16629);
nor U21820 (N_21820,N_18940,N_19161);
nand U21821 (N_21821,N_17131,N_19371);
nand U21822 (N_21822,N_18221,N_18897);
and U21823 (N_21823,N_16387,N_19105);
nand U21824 (N_21824,N_15548,N_16678);
and U21825 (N_21825,N_18990,N_17378);
or U21826 (N_21826,N_18499,N_18404);
xnor U21827 (N_21827,N_17314,N_16505);
and U21828 (N_21828,N_19463,N_19722);
nand U21829 (N_21829,N_18306,N_19925);
or U21830 (N_21830,N_19706,N_19023);
nand U21831 (N_21831,N_17719,N_19349);
xor U21832 (N_21832,N_18654,N_19493);
nand U21833 (N_21833,N_15611,N_19965);
nand U21834 (N_21834,N_16584,N_19338);
nand U21835 (N_21835,N_19321,N_17652);
nand U21836 (N_21836,N_17361,N_15375);
nand U21837 (N_21837,N_18184,N_17706);
and U21838 (N_21838,N_17222,N_18433);
nand U21839 (N_21839,N_17254,N_15909);
xor U21840 (N_21840,N_18913,N_18242);
or U21841 (N_21841,N_18645,N_17340);
or U21842 (N_21842,N_17713,N_19262);
and U21843 (N_21843,N_15235,N_19905);
nand U21844 (N_21844,N_17079,N_16250);
nor U21845 (N_21845,N_18250,N_18037);
and U21846 (N_21846,N_15432,N_18951);
nand U21847 (N_21847,N_15228,N_18316);
xor U21848 (N_21848,N_16909,N_18810);
or U21849 (N_21849,N_17810,N_19737);
xor U21850 (N_21850,N_15831,N_17850);
nor U21851 (N_21851,N_19131,N_19417);
or U21852 (N_21852,N_15065,N_15421);
nor U21853 (N_21853,N_17133,N_19629);
nor U21854 (N_21854,N_19152,N_15856);
nand U21855 (N_21855,N_17156,N_18489);
and U21856 (N_21856,N_17193,N_18098);
or U21857 (N_21857,N_19491,N_18781);
xnor U21858 (N_21858,N_16146,N_15225);
or U21859 (N_21859,N_19730,N_17008);
xor U21860 (N_21860,N_19378,N_19219);
xor U21861 (N_21861,N_19779,N_18362);
or U21862 (N_21862,N_17880,N_19642);
nor U21863 (N_21863,N_18598,N_18333);
or U21864 (N_21864,N_19698,N_19546);
xnor U21865 (N_21865,N_16923,N_17869);
and U21866 (N_21866,N_17675,N_19868);
or U21867 (N_21867,N_17519,N_16766);
nand U21868 (N_21868,N_17349,N_17583);
xor U21869 (N_21869,N_16518,N_15494);
or U21870 (N_21870,N_19745,N_15132);
nor U21871 (N_21871,N_19026,N_18044);
nand U21872 (N_21872,N_19563,N_18536);
nor U21873 (N_21873,N_16070,N_18765);
and U21874 (N_21874,N_15564,N_18481);
or U21875 (N_21875,N_17000,N_19733);
nand U21876 (N_21876,N_18159,N_16006);
nand U21877 (N_21877,N_19203,N_15957);
and U21878 (N_21878,N_16645,N_16621);
and U21879 (N_21879,N_17859,N_19496);
and U21880 (N_21880,N_18341,N_18669);
nand U21881 (N_21881,N_16938,N_16260);
xnor U21882 (N_21882,N_18627,N_16622);
or U21883 (N_21883,N_17907,N_17899);
and U21884 (N_21884,N_16788,N_18513);
nor U21885 (N_21885,N_15850,N_18708);
nor U21886 (N_21886,N_19396,N_15438);
and U21887 (N_21887,N_16148,N_15126);
nor U21888 (N_21888,N_18831,N_19500);
and U21889 (N_21889,N_17484,N_19870);
and U21890 (N_21890,N_17944,N_16706);
and U21891 (N_21891,N_17639,N_16628);
or U21892 (N_21892,N_17542,N_17209);
or U21893 (N_21893,N_19159,N_18337);
or U21894 (N_21894,N_15838,N_19025);
nor U21895 (N_21895,N_18450,N_15782);
xnor U21896 (N_21896,N_17607,N_17505);
and U21897 (N_21897,N_18089,N_18146);
or U21898 (N_21898,N_15337,N_15054);
xnor U21899 (N_21899,N_19452,N_17683);
nand U21900 (N_21900,N_19059,N_17768);
nand U21901 (N_21901,N_15419,N_16969);
xnor U21902 (N_21902,N_17949,N_17294);
or U21903 (N_21903,N_16670,N_16380);
xnor U21904 (N_21904,N_17114,N_15572);
and U21905 (N_21905,N_15082,N_16226);
or U21906 (N_21906,N_15417,N_15497);
xor U21907 (N_21907,N_18518,N_16683);
xnor U21908 (N_21908,N_16238,N_15945);
or U21909 (N_21909,N_16421,N_19859);
or U21910 (N_21910,N_18398,N_19094);
and U21911 (N_21911,N_17160,N_17423);
nor U21912 (N_21912,N_16391,N_15338);
and U21913 (N_21913,N_15050,N_18923);
xor U21914 (N_21914,N_19505,N_19351);
or U21915 (N_21915,N_19213,N_18701);
xor U21916 (N_21916,N_16951,N_15786);
xnor U21917 (N_21917,N_15053,N_18721);
nor U21918 (N_21918,N_16922,N_19820);
xnor U21919 (N_21919,N_15843,N_17115);
nor U21920 (N_21920,N_17457,N_19694);
xor U21921 (N_21921,N_15488,N_17382);
and U21922 (N_21922,N_19618,N_19113);
xor U21923 (N_21923,N_16465,N_15820);
or U21924 (N_21924,N_16178,N_19067);
nor U21925 (N_21925,N_16304,N_17376);
and U21926 (N_21926,N_19448,N_15210);
nand U21927 (N_21927,N_15700,N_17388);
or U21928 (N_21928,N_15890,N_17746);
and U21929 (N_21929,N_15947,N_17912);
xnor U21930 (N_21930,N_19819,N_17479);
or U21931 (N_21931,N_15329,N_17202);
nand U21932 (N_21932,N_17302,N_16372);
and U21933 (N_21933,N_18467,N_16950);
and U21934 (N_21934,N_15728,N_15582);
or U21935 (N_21935,N_15996,N_17894);
xor U21936 (N_21936,N_16180,N_15976);
xor U21937 (N_21937,N_19012,N_15608);
nor U21938 (N_21938,N_17531,N_16229);
and U21939 (N_21939,N_15754,N_18335);
nor U21940 (N_21940,N_15312,N_15959);
nand U21941 (N_21941,N_18864,N_19504);
xor U21942 (N_21942,N_17882,N_18156);
or U21943 (N_21943,N_16889,N_17392);
nor U21944 (N_21944,N_18457,N_17399);
nand U21945 (N_21945,N_19416,N_19602);
or U21946 (N_21946,N_17047,N_16709);
or U21947 (N_21947,N_19032,N_18840);
and U21948 (N_21948,N_19879,N_17674);
xor U21949 (N_21949,N_16741,N_15070);
xnor U21950 (N_21950,N_18742,N_15748);
nand U21951 (N_21951,N_18245,N_16054);
xnor U21952 (N_21952,N_17983,N_18171);
nor U21953 (N_21953,N_19791,N_17776);
xor U21954 (N_21954,N_19293,N_16700);
or U21955 (N_21955,N_16870,N_18523);
and U21956 (N_21956,N_19630,N_18947);
nand U21957 (N_21957,N_18789,N_17833);
or U21958 (N_21958,N_19592,N_17057);
xnor U21959 (N_21959,N_15055,N_18590);
nor U21960 (N_21960,N_17168,N_18059);
or U21961 (N_21961,N_17390,N_16217);
and U21962 (N_21962,N_18549,N_16009);
or U21963 (N_21963,N_16460,N_18286);
xnor U21964 (N_21964,N_15873,N_15207);
xnor U21965 (N_21965,N_16756,N_16467);
xnor U21966 (N_21966,N_16024,N_16663);
or U21967 (N_21967,N_19373,N_16949);
and U21968 (N_21968,N_16937,N_18330);
xnor U21969 (N_21969,N_17496,N_19788);
and U21970 (N_21970,N_15504,N_19445);
or U21971 (N_21971,N_17238,N_17780);
nor U21972 (N_21972,N_15636,N_17259);
and U21973 (N_21973,N_15383,N_16759);
or U21974 (N_21974,N_15524,N_16824);
xor U21975 (N_21975,N_15915,N_18799);
or U21976 (N_21976,N_17625,N_17648);
and U21977 (N_21977,N_19158,N_16802);
or U21978 (N_21978,N_16415,N_16049);
nand U21979 (N_21979,N_16047,N_17319);
nor U21980 (N_21980,N_19862,N_18915);
and U21981 (N_21981,N_15435,N_15793);
xor U21982 (N_21982,N_19370,N_18304);
and U21983 (N_21983,N_17570,N_18270);
or U21984 (N_21984,N_16701,N_16063);
xor U21985 (N_21985,N_16418,N_16082);
nand U21986 (N_21986,N_16839,N_19873);
nand U21987 (N_21987,N_18768,N_18529);
and U21988 (N_21988,N_16104,N_18905);
and U21989 (N_21989,N_19682,N_19810);
and U21990 (N_21990,N_18787,N_16100);
or U21991 (N_21991,N_19129,N_17439);
xnor U21992 (N_21992,N_18048,N_17472);
nor U21993 (N_21993,N_18846,N_18560);
xor U21994 (N_21994,N_17445,N_19337);
nor U21995 (N_21995,N_15567,N_16432);
or U21996 (N_21996,N_15859,N_15381);
and U21997 (N_21997,N_16128,N_18170);
or U21998 (N_21998,N_18344,N_15712);
or U21999 (N_21999,N_17572,N_17492);
nor U22000 (N_22000,N_16976,N_17173);
or U22001 (N_22001,N_18910,N_17515);
nor U22002 (N_22002,N_15991,N_18777);
and U22003 (N_22003,N_19765,N_16529);
nor U22004 (N_22004,N_19959,N_17784);
xor U22005 (N_22005,N_15468,N_16497);
and U22006 (N_22006,N_15446,N_19150);
nor U22007 (N_22007,N_16778,N_15686);
or U22008 (N_22008,N_19409,N_19220);
nand U22009 (N_22009,N_16653,N_18798);
nand U22010 (N_22010,N_15237,N_16227);
nor U22011 (N_22011,N_19958,N_17770);
and U22012 (N_22012,N_17966,N_17172);
nand U22013 (N_22013,N_16157,N_15726);
and U22014 (N_22014,N_19535,N_16360);
or U22015 (N_22015,N_19637,N_15413);
xnor U22016 (N_22016,N_16023,N_18014);
xnor U22017 (N_22017,N_15075,N_18917);
nand U22018 (N_22018,N_17397,N_16910);
nand U22019 (N_22019,N_15204,N_17468);
or U22020 (N_22020,N_19685,N_19511);
or U22021 (N_22021,N_16291,N_18574);
xor U22022 (N_22022,N_16403,N_18264);
and U22023 (N_22023,N_17243,N_19160);
nor U22024 (N_22024,N_16833,N_16256);
nor U22025 (N_22025,N_15773,N_19817);
nor U22026 (N_22026,N_19814,N_18456);
nor U22027 (N_22027,N_17329,N_19215);
nand U22028 (N_22028,N_17819,N_16469);
nor U22029 (N_22029,N_19683,N_15989);
and U22030 (N_22030,N_17108,N_19725);
and U22031 (N_22031,N_16111,N_16106);
nor U22032 (N_22032,N_17052,N_17587);
xor U22033 (N_22033,N_16575,N_19218);
nor U22034 (N_22034,N_16031,N_17438);
nor U22035 (N_22035,N_16275,N_18236);
or U22036 (N_22036,N_16989,N_16731);
nand U22037 (N_22037,N_15839,N_15948);
and U22038 (N_22038,N_19261,N_18074);
and U22039 (N_22039,N_16073,N_15617);
nor U22040 (N_22040,N_16315,N_15633);
nor U22041 (N_22041,N_16566,N_15984);
or U22042 (N_22042,N_18313,N_16804);
nand U22043 (N_22043,N_16807,N_15479);
or U22044 (N_22044,N_18997,N_17013);
or U22045 (N_22045,N_19322,N_17077);
nand U22046 (N_22046,N_17820,N_18510);
or U22047 (N_22047,N_15127,N_19775);
or U22048 (N_22048,N_17023,N_19250);
xnor U22049 (N_22049,N_15193,N_16619);
or U22050 (N_22050,N_18725,N_15544);
and U22051 (N_22051,N_17499,N_18312);
or U22052 (N_22052,N_16545,N_15549);
or U22053 (N_22053,N_18094,N_16029);
xnor U22054 (N_22054,N_19880,N_17837);
nor U22055 (N_22055,N_16102,N_17260);
nand U22056 (N_22056,N_19714,N_18001);
and U22057 (N_22057,N_16591,N_19964);
nor U22058 (N_22058,N_18493,N_19588);
and U22059 (N_22059,N_18186,N_16232);
xor U22060 (N_22060,N_17028,N_17312);
xnor U22061 (N_22061,N_17051,N_19387);
nand U22062 (N_22062,N_19066,N_19830);
or U22063 (N_22063,N_17054,N_18161);
nand U22064 (N_22064,N_18749,N_16789);
or U22065 (N_22065,N_19283,N_15245);
nand U22066 (N_22066,N_15309,N_15710);
or U22067 (N_22067,N_18039,N_18325);
xor U22068 (N_22068,N_16491,N_17687);
or U22069 (N_22069,N_15489,N_18930);
xor U22070 (N_22070,N_17024,N_15679);
and U22071 (N_22071,N_17653,N_15227);
or U22072 (N_22072,N_19962,N_17582);
nand U22073 (N_22073,N_15359,N_19567);
nor U22074 (N_22074,N_16434,N_16325);
xor U22075 (N_22075,N_19436,N_15660);
nor U22076 (N_22076,N_19296,N_16014);
or U22077 (N_22077,N_16322,N_18823);
and U22078 (N_22078,N_16475,N_16607);
and U22079 (N_22079,N_17811,N_17174);
nor U22080 (N_22080,N_18963,N_15298);
or U22081 (N_22081,N_19318,N_19953);
nor U22082 (N_22082,N_15523,N_16055);
xor U22083 (N_22083,N_17331,N_15836);
nor U22084 (N_22084,N_18881,N_16941);
nand U22085 (N_22085,N_19717,N_17762);
nand U22086 (N_22086,N_16235,N_19860);
and U22087 (N_22087,N_17105,N_17007);
nand U22088 (N_22088,N_19551,N_17461);
and U22089 (N_22089,N_18702,N_18591);
nor U22090 (N_22090,N_16806,N_18487);
nor U22091 (N_22091,N_16680,N_19576);
nand U22092 (N_22092,N_18884,N_17796);
or U22093 (N_22093,N_19249,N_15017);
xnor U22094 (N_22094,N_15122,N_17045);
or U22095 (N_22095,N_17974,N_17321);
nand U22096 (N_22096,N_15825,N_16975);
or U22097 (N_22097,N_19750,N_16445);
nand U22098 (N_22098,N_15761,N_17303);
nor U22099 (N_22099,N_15343,N_18763);
nand U22100 (N_22100,N_19586,N_15888);
nor U22101 (N_22101,N_16334,N_19434);
or U22102 (N_22102,N_15809,N_19935);
nor U22103 (N_22103,N_19651,N_19297);
or U22104 (N_22104,N_15173,N_17387);
nor U22105 (N_22105,N_18678,N_18531);
or U22106 (N_22106,N_16879,N_17967);
xor U22107 (N_22107,N_18987,N_17149);
nor U22108 (N_22108,N_18497,N_18704);
nand U22109 (N_22109,N_17493,N_15114);
xnor U22110 (N_22110,N_16034,N_15727);
nand U22111 (N_22111,N_17073,N_19011);
nand U22112 (N_22112,N_19077,N_17112);
xor U22113 (N_22113,N_19547,N_16868);
and U22114 (N_22114,N_19866,N_18876);
nand U22115 (N_22115,N_16308,N_15804);
and U22116 (N_22116,N_15813,N_15415);
nor U22117 (N_22117,N_15631,N_18925);
xor U22118 (N_22118,N_16172,N_18289);
nor U22119 (N_22119,N_18774,N_19217);
nor U22120 (N_22120,N_15645,N_17756);
or U22121 (N_22121,N_18596,N_18376);
xor U22122 (N_22122,N_19393,N_16038);
or U22123 (N_22123,N_16201,N_19992);
and U22124 (N_22124,N_18974,N_15480);
nand U22125 (N_22125,N_19054,N_15357);
xor U22126 (N_22126,N_19114,N_18157);
and U22127 (N_22127,N_18080,N_15842);
xor U22128 (N_22128,N_16124,N_19000);
nor U22129 (N_22129,N_17783,N_18524);
and U22130 (N_22130,N_17658,N_16967);
and U22131 (N_22131,N_16736,N_16450);
nand U22132 (N_22132,N_19898,N_17158);
nor U22133 (N_22133,N_17012,N_15798);
xnor U22134 (N_22134,N_18587,N_17085);
xnor U22135 (N_22135,N_15864,N_19716);
nand U22136 (N_22136,N_19799,N_16279);
nor U22137 (N_22137,N_18460,N_15735);
nor U22138 (N_22138,N_19103,N_18969);
xor U22139 (N_22139,N_18919,N_19144);
nor U22140 (N_22140,N_15932,N_16887);
nand U22141 (N_22141,N_17739,N_19973);
and U22142 (N_22142,N_15269,N_17630);
and U22143 (N_22143,N_18070,N_16624);
xnor U22144 (N_22144,N_18147,N_16650);
and U22145 (N_22145,N_17166,N_17187);
nor U22146 (N_22146,N_16805,N_18096);
nor U22147 (N_22147,N_16638,N_16642);
nand U22148 (N_22148,N_16140,N_15351);
nand U22149 (N_22149,N_15465,N_15910);
or U22150 (N_22150,N_19310,N_15066);
and U22151 (N_22151,N_16341,N_16258);
nand U22152 (N_22152,N_16130,N_17842);
xor U22153 (N_22153,N_18189,N_18177);
xnor U22154 (N_22154,N_18843,N_17509);
xor U22155 (N_22155,N_18502,N_16984);
nor U22156 (N_22156,N_19711,N_15011);
xor U22157 (N_22157,N_17567,N_15077);
and U22158 (N_22158,N_17664,N_15739);
nor U22159 (N_22159,N_15521,N_16406);
nor U22160 (N_22160,N_17356,N_17516);
xor U22161 (N_22161,N_16846,N_16371);
xnor U22162 (N_22162,N_16668,N_19885);
nor U22163 (N_22163,N_18832,N_19872);
nor U22164 (N_22164,N_19723,N_18602);
and U22165 (N_22165,N_19800,N_17846);
nor U22166 (N_22166,N_15374,N_15552);
xnor U22167 (N_22167,N_15586,N_16963);
and U22168 (N_22168,N_15515,N_16876);
nand U22169 (N_22169,N_16453,N_19514);
nor U22170 (N_22170,N_18071,N_19061);
xnor U22171 (N_22171,N_19553,N_19877);
xor U22172 (N_22172,N_19391,N_18272);
or U22173 (N_22173,N_19440,N_15653);
or U22174 (N_22174,N_15853,N_16559);
xor U22175 (N_22175,N_15961,N_17288);
and U22176 (N_22176,N_18152,N_19455);
or U22177 (N_22177,N_19169,N_17038);
and U22178 (N_22178,N_15145,N_19573);
or U22179 (N_22179,N_18830,N_19058);
nor U22180 (N_22180,N_17157,N_16992);
or U22181 (N_22181,N_16498,N_17935);
nand U22182 (N_22182,N_17018,N_19424);
nand U22183 (N_22183,N_15366,N_17916);
and U22184 (N_22184,N_17920,N_17335);
nor U22185 (N_22185,N_18357,N_17914);
and U22186 (N_22186,N_19653,N_18354);
nor U22187 (N_22187,N_18698,N_18369);
or U22188 (N_22188,N_16580,N_15600);
or U22189 (N_22189,N_19482,N_16295);
or U22190 (N_22190,N_18185,N_17500);
xnor U22191 (N_22191,N_19823,N_16719);
or U22192 (N_22192,N_18387,N_18292);
nand U22193 (N_22193,N_18230,N_17759);
nand U22194 (N_22194,N_16470,N_15897);
or U22195 (N_22195,N_19740,N_15532);
or U22196 (N_22196,N_17779,N_18555);
xnor U22197 (N_22197,N_19752,N_19771);
and U22198 (N_22198,N_15674,N_18703);
and U22199 (N_22199,N_16981,N_17511);
and U22200 (N_22200,N_19033,N_17104);
and U22201 (N_22201,N_18007,N_15597);
or U22202 (N_22202,N_17276,N_18190);
or U22203 (N_22203,N_17237,N_17039);
or U22204 (N_22204,N_15449,N_19291);
nor U22205 (N_22205,N_17106,N_15382);
and U22206 (N_22206,N_19583,N_16845);
or U22207 (N_22207,N_19280,N_19569);
nand U22208 (N_22208,N_15514,N_17644);
or U22209 (N_22209,N_19295,N_16579);
nor U22210 (N_22210,N_18024,N_19101);
or U22211 (N_22211,N_17991,N_16735);
or U22212 (N_22212,N_15779,N_19145);
or U22213 (N_22213,N_16369,N_15872);
nor U22214 (N_22214,N_15169,N_17689);
or U22215 (N_22215,N_16028,N_18858);
xor U22216 (N_22216,N_18082,N_15750);
and U22217 (N_22217,N_15849,N_16408);
and U22218 (N_22218,N_18095,N_15911);
xnor U22219 (N_22219,N_18908,N_19124);
xnor U22220 (N_22220,N_18659,N_15266);
and U22221 (N_22221,N_18090,N_16924);
or U22222 (N_22222,N_16925,N_15807);
nand U22223 (N_22223,N_16463,N_16769);
and U22224 (N_22224,N_17637,N_15205);
and U22225 (N_22225,N_19656,N_18845);
nand U22226 (N_22226,N_15550,N_17270);
nand U22227 (N_22227,N_16986,N_16533);
nor U22228 (N_22228,N_15634,N_16433);
nand U22229 (N_22229,N_17620,N_15090);
nor U22230 (N_22230,N_18124,N_17218);
nor U22231 (N_22231,N_19928,N_17311);
nand U22232 (N_22232,N_18310,N_18284);
or U22233 (N_22233,N_17255,N_19208);
xnor U22234 (N_22234,N_19606,N_16119);
or U22235 (N_22235,N_18534,N_15019);
nor U22236 (N_22236,N_18182,N_17076);
xor U22237 (N_22237,N_16384,N_17743);
or U22238 (N_22238,N_19666,N_18078);
and U22239 (N_22239,N_19320,N_19271);
nand U22240 (N_22240,N_18097,N_18020);
nor U22241 (N_22241,N_15928,N_18873);
xor U22242 (N_22242,N_15398,N_19695);
nand U22243 (N_22243,N_17612,N_15771);
nand U22244 (N_22244,N_17919,N_18664);
nand U22245 (N_22245,N_17662,N_18710);
and U22246 (N_22246,N_19616,N_19570);
or U22247 (N_22247,N_19645,N_16053);
xor U22248 (N_22248,N_17436,N_17494);
nand U22249 (N_22249,N_17508,N_19543);
and U22250 (N_22250,N_19270,N_16480);
nor U22251 (N_22251,N_15529,N_18241);
nand U22252 (N_22252,N_17244,N_15416);
nor U22253 (N_22253,N_16494,N_16601);
or U22254 (N_22254,N_19087,N_19222);
nor U22255 (N_22255,N_18058,N_15321);
nand U22256 (N_22256,N_18263,N_17877);
nor U22257 (N_22257,N_17848,N_19224);
nor U22258 (N_22258,N_18511,N_17529);
xnor U22259 (N_22259,N_15403,N_16137);
or U22260 (N_22260,N_18805,N_18604);
and U22261 (N_22261,N_19865,N_17078);
xor U22262 (N_22262,N_19036,N_15259);
nor U22263 (N_22263,N_15591,N_16289);
and U22264 (N_22264,N_17235,N_15284);
and U22265 (N_22265,N_18638,N_15401);
and U22266 (N_22266,N_18570,N_17075);
or U22267 (N_22267,N_17344,N_19277);
nor U22268 (N_22268,N_18445,N_15426);
and U22269 (N_22269,N_18367,N_17313);
and U22270 (N_22270,N_19728,N_16300);
nor U22271 (N_22271,N_15117,N_19635);
nor U22272 (N_22272,N_17341,N_18346);
and U22273 (N_22273,N_18706,N_15543);
xnor U22274 (N_22274,N_16517,N_15574);
nor U22275 (N_22275,N_18603,N_16661);
nor U22276 (N_22276,N_19906,N_18343);
nand U22277 (N_22277,N_18342,N_15460);
nor U22278 (N_22278,N_17394,N_15627);
and U22279 (N_22279,N_15360,N_15024);
xnor U22280 (N_22280,N_19850,N_18228);
or U22281 (N_22281,N_15461,N_16782);
and U22282 (N_22282,N_18802,N_18752);
xor U22283 (N_22283,N_17192,N_17778);
nor U22284 (N_22284,N_17993,N_16502);
nor U22285 (N_22285,N_17565,N_15196);
and U22286 (N_22286,N_18267,N_19684);
and U22287 (N_22287,N_19759,N_19071);
xor U22288 (N_22288,N_19404,N_17315);
nor U22289 (N_22289,N_16538,N_19561);
nor U22290 (N_22290,N_18486,N_18733);
nand U22291 (N_22291,N_19466,N_17025);
or U22292 (N_22292,N_17228,N_17210);
xor U22293 (N_22293,N_16681,N_16996);
or U22294 (N_22294,N_18415,N_16587);
xor U22295 (N_22295,N_17470,N_17124);
xnor U22296 (N_22296,N_15035,N_16971);
xor U22297 (N_22297,N_17448,N_15829);
xor U22298 (N_22298,N_15648,N_17835);
nand U22299 (N_22299,N_15469,N_15568);
xor U22300 (N_22300,N_17409,N_17593);
or U22301 (N_22301,N_17611,N_19437);
nand U22302 (N_22302,N_19833,N_18626);
nand U22303 (N_22303,N_19176,N_19792);
nand U22304 (N_22304,N_17481,N_19834);
and U22305 (N_22305,N_19352,N_16961);
xnor U22306 (N_22306,N_16435,N_17282);
and U22307 (N_22307,N_15818,N_17686);
and U22308 (N_22308,N_18060,N_18462);
and U22309 (N_22309,N_18743,N_18856);
or U22310 (N_22310,N_15279,N_18069);
nor U22311 (N_22311,N_18695,N_18601);
nand U22312 (N_22312,N_19002,N_18248);
nor U22313 (N_22313,N_15270,N_16150);
xnor U22314 (N_22314,N_17506,N_18382);
nor U22315 (N_22315,N_19536,N_16626);
nor U22316 (N_22316,N_16090,N_18195);
xnor U22317 (N_22317,N_18299,N_17578);
nand U22318 (N_22318,N_19069,N_19657);
and U22319 (N_22319,N_18431,N_17628);
xnor U22320 (N_22320,N_16060,N_15906);
nor U22321 (N_22321,N_17972,N_16724);
and U22322 (N_22322,N_19001,N_18803);
xnor U22323 (N_22323,N_18033,N_18318);
nor U22324 (N_22324,N_17308,N_15563);
or U22325 (N_22325,N_19951,N_15440);
and U22326 (N_22326,N_17752,N_16310);
nand U22327 (N_22327,N_19644,N_16089);
or U22328 (N_22328,N_18407,N_17748);
nand U22329 (N_22329,N_16875,N_19578);
nor U22330 (N_22330,N_16007,N_19784);
nand U22331 (N_22331,N_19949,N_19348);
nand U22332 (N_22332,N_19916,N_15044);
xnor U22333 (N_22333,N_18319,N_18932);
nand U22334 (N_22334,N_18405,N_15962);
nand U22335 (N_22335,N_18674,N_17790);
and U22336 (N_22336,N_18775,N_19266);
xor U22337 (N_22337,N_18137,N_17870);
and U22338 (N_22338,N_19911,N_17851);
or U22339 (N_22339,N_17463,N_15570);
nand U22340 (N_22340,N_15156,N_18720);
xor U22341 (N_22341,N_19516,N_19426);
or U22342 (N_22342,N_18216,N_15384);
and U22343 (N_22343,N_17697,N_18785);
nand U22344 (N_22344,N_18364,N_18663);
nand U22345 (N_22345,N_15595,N_15817);
and U22346 (N_22346,N_19710,N_19192);
and U22347 (N_22347,N_16348,N_17262);
xnor U22348 (N_22348,N_16057,N_18443);
nand U22349 (N_22349,N_17489,N_17066);
nand U22350 (N_22350,N_19988,N_15553);
nand U22351 (N_22351,N_15721,N_15184);
and U22352 (N_22352,N_16899,N_16549);
nor U22353 (N_22353,N_18477,N_19162);
or U22354 (N_22354,N_16097,N_17383);
nor U22355 (N_22355,N_15042,N_18172);
and U22356 (N_22356,N_17408,N_16751);
or U22357 (N_22357,N_19447,N_19029);
and U22358 (N_22358,N_17458,N_15545);
or U22359 (N_22359,N_19886,N_17853);
or U22360 (N_22360,N_15422,N_19729);
or U22361 (N_22361,N_17886,N_17586);
and U22362 (N_22362,N_18274,N_19273);
or U22363 (N_22363,N_16774,N_15463);
or U22364 (N_22364,N_19783,N_16798);
nand U22365 (N_22365,N_19841,N_19476);
nor U22366 (N_22366,N_18815,N_17924);
or U22367 (N_22367,N_17590,N_19185);
and U22368 (N_22368,N_16615,N_17195);
and U22369 (N_22369,N_16800,N_16803);
nand U22370 (N_22370,N_15004,N_19655);
nor U22371 (N_22371,N_19049,N_16324);
nor U22372 (N_22372,N_19529,N_17019);
nor U22373 (N_22373,N_19672,N_19575);
nand U22374 (N_22374,N_19990,N_15876);
nand U22375 (N_22375,N_15643,N_18379);
nand U22376 (N_22376,N_15186,N_15812);
nand U22377 (N_22377,N_17831,N_18999);
xor U22378 (N_22378,N_19172,N_16596);
nor U22379 (N_22379,N_18966,N_18005);
xnor U22380 (N_22380,N_16103,N_16568);
nand U22381 (N_22381,N_19022,N_18442);
nor U22382 (N_22382,N_19571,N_17546);
nor U22383 (N_22383,N_16837,N_16123);
xor U22384 (N_22384,N_18506,N_17589);
and U22385 (N_22385,N_16912,N_17004);
and U22386 (N_22386,N_19498,N_18612);
nand U22387 (N_22387,N_19244,N_16074);
or U22388 (N_22388,N_16717,N_17380);
nor U22389 (N_22389,N_16378,N_16439);
xor U22390 (N_22390,N_15790,N_19754);
nor U22391 (N_22391,N_18377,N_15358);
or U22392 (N_22392,N_17178,N_19153);
or U22393 (N_22393,N_15138,N_18361);
nor U22394 (N_22394,N_17403,N_17596);
xor U22395 (N_22395,N_15405,N_16685);
xnor U22396 (N_22396,N_16516,N_17310);
xnor U22397 (N_22397,N_17082,N_15305);
nor U22398 (N_22398,N_16072,N_15188);
nand U22399 (N_22399,N_18175,N_17647);
xor U22400 (N_22400,N_16542,N_18540);
nand U22401 (N_22401,N_15981,N_18444);
nand U22402 (N_22402,N_15477,N_19303);
and U22403 (N_22403,N_19408,N_16396);
or U22404 (N_22404,N_19450,N_18178);
xnor U22405 (N_22405,N_16603,N_18821);
xnor U22406 (N_22406,N_18389,N_19611);
nand U22407 (N_22407,N_16891,N_15926);
nor U22408 (N_22408,N_19205,N_16974);
xor U22409 (N_22409,N_18358,N_15934);
or U22410 (N_22410,N_16375,N_16486);
nand U22411 (N_22411,N_18375,N_19386);
and U22412 (N_22412,N_19018,N_17385);
nand U22413 (N_22413,N_18393,N_17657);
or U22414 (N_22414,N_19083,N_17125);
nor U22415 (N_22415,N_18958,N_16752);
and U22416 (N_22416,N_18000,N_16562);
nand U22417 (N_22417,N_15683,N_18057);
nor U22418 (N_22418,N_17876,N_15190);
nor U22419 (N_22419,N_15353,N_18302);
or U22420 (N_22420,N_15313,N_16166);
nor U22421 (N_22421,N_19421,N_15642);
and U22422 (N_22422,N_15687,N_15140);
or U22423 (N_22423,N_16618,N_19887);
or U22424 (N_22424,N_18629,N_16298);
or U22425 (N_22425,N_19045,N_15160);
xnor U22426 (N_22426,N_18796,N_19909);
or U22427 (N_22427,N_16004,N_17599);
nor U22428 (N_22428,N_18921,N_19687);
or U22429 (N_22429,N_15640,N_18891);
xor U22430 (N_22430,N_16964,N_16228);
and U22431 (N_22431,N_19369,N_19908);
xnor U22432 (N_22432,N_19743,N_18824);
and U22433 (N_22433,N_18046,N_15041);
nor U22434 (N_22434,N_17099,N_17346);
and U22435 (N_22435,N_15217,N_15002);
and U22436 (N_22436,N_17236,N_18446);
xor U22437 (N_22437,N_18416,N_18359);
nor U22438 (N_22438,N_18479,N_17560);
nand U22439 (N_22439,N_15273,N_19116);
nand U22440 (N_22440,N_16194,N_17198);
nor U22441 (N_22441,N_16682,N_19986);
nand U22442 (N_22442,N_18138,N_17659);
xor U22443 (N_22443,N_15635,N_17902);
nand U22444 (N_22444,N_16936,N_15088);
and U22445 (N_22445,N_17220,N_16696);
xor U22446 (N_22446,N_15985,N_19314);
xnor U22447 (N_22447,N_19174,N_19227);
or U22448 (N_22448,N_18746,N_18143);
xor U22449 (N_22449,N_15941,N_18697);
nor U22450 (N_22450,N_17101,N_15975);
nand U22451 (N_22451,N_15389,N_15251);
xnor U22452 (N_22452,N_15111,N_16105);
and U22453 (N_22453,N_15466,N_16758);
nor U22454 (N_22454,N_19275,N_16410);
and U22455 (N_22455,N_17447,N_18895);
xor U22456 (N_22456,N_18989,N_19974);
or U22457 (N_22457,N_15166,N_16617);
nand U22458 (N_22458,N_19052,N_19195);
xnor U22459 (N_22459,N_16485,N_17745);
nor U22460 (N_22460,N_18088,N_16329);
or U22461 (N_22461,N_16515,N_17650);
xor U22462 (N_22462,N_18029,N_17199);
xor U22463 (N_22463,N_15260,N_16843);
and U22464 (N_22464,N_17544,N_17285);
nand U22465 (N_22465,N_19857,N_19357);
nor U22466 (N_22466,N_15784,N_16968);
or U22467 (N_22467,N_17204,N_18435);
or U22468 (N_22468,N_16672,N_15556);
and U22469 (N_22469,N_18064,N_19432);
nand U22470 (N_22470,N_17855,N_18980);
nand U22471 (N_22471,N_17336,N_19050);
or U22472 (N_22472,N_16988,N_18110);
nor U22473 (N_22473,N_15606,N_19593);
nand U22474 (N_22474,N_15241,N_18705);
nand U22475 (N_22475,N_15860,N_18244);
xnor U22476 (N_22476,N_19662,N_16519);
nor U22477 (N_22477,N_15538,N_15092);
nand U22478 (N_22478,N_16084,N_18971);
nor U22479 (N_22479,N_16512,N_15781);
nor U22480 (N_22480,N_18388,N_18384);
xor U22481 (N_22481,N_19673,N_15960);
or U22482 (N_22482,N_15022,N_16815);
xnor U22483 (N_22483,N_18085,N_19675);
nor U22484 (N_22484,N_19983,N_16163);
or U22485 (N_22485,N_18588,N_16139);
or U22486 (N_22486,N_15774,N_17398);
nor U22487 (N_22487,N_18287,N_15020);
xor U22488 (N_22488,N_19042,N_16586);
nand U22489 (N_22489,N_18844,N_18793);
xnor U22490 (N_22490,N_15848,N_16411);
nor U22491 (N_22491,N_17200,N_18633);
nor U22492 (N_22492,N_16561,N_19480);
xor U22493 (N_22493,N_15407,N_15379);
nor U22494 (N_22494,N_18002,N_19327);
and U22495 (N_22495,N_19774,N_17452);
nand U22496 (N_22496,N_16203,N_18714);
nand U22497 (N_22497,N_18794,N_19252);
nand U22498 (N_22498,N_17769,N_19832);
or U22499 (N_22499,N_18121,N_15639);
nand U22500 (N_22500,N_17631,N_15090);
nor U22501 (N_22501,N_18908,N_19641);
and U22502 (N_22502,N_17338,N_18209);
nor U22503 (N_22503,N_15449,N_16671);
nand U22504 (N_22504,N_17713,N_19292);
nand U22505 (N_22505,N_15837,N_18957);
nor U22506 (N_22506,N_16769,N_18408);
nor U22507 (N_22507,N_17886,N_19950);
nand U22508 (N_22508,N_18865,N_16253);
or U22509 (N_22509,N_15240,N_16343);
and U22510 (N_22510,N_17274,N_18706);
and U22511 (N_22511,N_19909,N_18155);
xor U22512 (N_22512,N_19080,N_18792);
xor U22513 (N_22513,N_18625,N_15202);
nand U22514 (N_22514,N_17935,N_18863);
or U22515 (N_22515,N_15381,N_19055);
or U22516 (N_22516,N_15684,N_19639);
and U22517 (N_22517,N_15297,N_15798);
nor U22518 (N_22518,N_16766,N_17570);
xnor U22519 (N_22519,N_16838,N_16266);
nand U22520 (N_22520,N_17044,N_18621);
xor U22521 (N_22521,N_15699,N_16845);
or U22522 (N_22522,N_18020,N_19616);
nand U22523 (N_22523,N_17568,N_18913);
xnor U22524 (N_22524,N_17966,N_15090);
xnor U22525 (N_22525,N_16662,N_19754);
nand U22526 (N_22526,N_15281,N_19733);
or U22527 (N_22527,N_17061,N_19062);
nand U22528 (N_22528,N_17971,N_19662);
or U22529 (N_22529,N_19782,N_18162);
xnor U22530 (N_22530,N_19169,N_16464);
xor U22531 (N_22531,N_15440,N_16735);
or U22532 (N_22532,N_15485,N_19608);
xnor U22533 (N_22533,N_15783,N_15521);
nor U22534 (N_22534,N_19884,N_16743);
or U22535 (N_22535,N_17074,N_16687);
nor U22536 (N_22536,N_17892,N_17008);
xnor U22537 (N_22537,N_16207,N_17669);
or U22538 (N_22538,N_18251,N_19457);
and U22539 (N_22539,N_18410,N_17809);
and U22540 (N_22540,N_17430,N_16468);
and U22541 (N_22541,N_17332,N_19141);
and U22542 (N_22542,N_15528,N_15994);
nand U22543 (N_22543,N_16432,N_19678);
nor U22544 (N_22544,N_15927,N_16869);
and U22545 (N_22545,N_19407,N_19633);
xor U22546 (N_22546,N_17228,N_15731);
nor U22547 (N_22547,N_19702,N_15733);
nand U22548 (N_22548,N_18897,N_15795);
nand U22549 (N_22549,N_16098,N_17692);
or U22550 (N_22550,N_16649,N_19086);
nand U22551 (N_22551,N_15371,N_19404);
xor U22552 (N_22552,N_15616,N_15778);
and U22553 (N_22553,N_18722,N_15241);
nor U22554 (N_22554,N_17563,N_16266);
or U22555 (N_22555,N_17961,N_15806);
xnor U22556 (N_22556,N_16998,N_19210);
nor U22557 (N_22557,N_16123,N_16247);
or U22558 (N_22558,N_18870,N_19652);
nor U22559 (N_22559,N_16560,N_18331);
and U22560 (N_22560,N_18145,N_15165);
nor U22561 (N_22561,N_17423,N_19000);
or U22562 (N_22562,N_18593,N_18704);
and U22563 (N_22563,N_15276,N_15430);
nand U22564 (N_22564,N_18507,N_15567);
and U22565 (N_22565,N_15831,N_19978);
nor U22566 (N_22566,N_19384,N_17037);
or U22567 (N_22567,N_19258,N_15157);
nand U22568 (N_22568,N_15563,N_19457);
or U22569 (N_22569,N_15372,N_17495);
or U22570 (N_22570,N_19512,N_16239);
and U22571 (N_22571,N_16380,N_16471);
xor U22572 (N_22572,N_18599,N_16980);
nor U22573 (N_22573,N_18269,N_17381);
and U22574 (N_22574,N_16469,N_15910);
xnor U22575 (N_22575,N_15595,N_19241);
nor U22576 (N_22576,N_16096,N_18978);
or U22577 (N_22577,N_17014,N_19206);
nor U22578 (N_22578,N_15648,N_18239);
or U22579 (N_22579,N_16434,N_15484);
nand U22580 (N_22580,N_19748,N_19628);
nor U22581 (N_22581,N_18677,N_15413);
nor U22582 (N_22582,N_18729,N_18322);
xor U22583 (N_22583,N_17074,N_17670);
nand U22584 (N_22584,N_19711,N_16030);
and U22585 (N_22585,N_16557,N_18071);
and U22586 (N_22586,N_16153,N_16244);
nor U22587 (N_22587,N_19831,N_17187);
nand U22588 (N_22588,N_18596,N_16282);
or U22589 (N_22589,N_18455,N_15289);
xnor U22590 (N_22590,N_19774,N_19349);
xnor U22591 (N_22591,N_15004,N_15106);
and U22592 (N_22592,N_18189,N_18114);
nor U22593 (N_22593,N_18325,N_16630);
nand U22594 (N_22594,N_15479,N_15117);
nor U22595 (N_22595,N_19405,N_19442);
and U22596 (N_22596,N_17192,N_19658);
nand U22597 (N_22597,N_19608,N_17581);
nor U22598 (N_22598,N_17239,N_15886);
and U22599 (N_22599,N_17606,N_18129);
nand U22600 (N_22600,N_16908,N_18288);
and U22601 (N_22601,N_15613,N_15900);
and U22602 (N_22602,N_15786,N_19227);
and U22603 (N_22603,N_19578,N_17390);
nor U22604 (N_22604,N_18530,N_15273);
or U22605 (N_22605,N_19975,N_17657);
nor U22606 (N_22606,N_18959,N_17036);
nor U22607 (N_22607,N_19885,N_18895);
nand U22608 (N_22608,N_18136,N_17589);
xor U22609 (N_22609,N_18259,N_16656);
nand U22610 (N_22610,N_18675,N_15722);
nor U22611 (N_22611,N_17749,N_19002);
and U22612 (N_22612,N_17264,N_18126);
xor U22613 (N_22613,N_19713,N_16403);
or U22614 (N_22614,N_16128,N_16876);
xnor U22615 (N_22615,N_18403,N_16976);
and U22616 (N_22616,N_16605,N_19438);
nand U22617 (N_22617,N_18549,N_19154);
xnor U22618 (N_22618,N_18407,N_18893);
and U22619 (N_22619,N_16573,N_19922);
nand U22620 (N_22620,N_18598,N_16739);
xnor U22621 (N_22621,N_17456,N_16484);
or U22622 (N_22622,N_19831,N_17470);
nand U22623 (N_22623,N_19623,N_17740);
xnor U22624 (N_22624,N_16324,N_18654);
and U22625 (N_22625,N_17310,N_18900);
nor U22626 (N_22626,N_17374,N_15959);
and U22627 (N_22627,N_19250,N_15000);
and U22628 (N_22628,N_15178,N_17511);
nand U22629 (N_22629,N_18767,N_19353);
xor U22630 (N_22630,N_19903,N_16258);
and U22631 (N_22631,N_19871,N_18490);
nand U22632 (N_22632,N_18686,N_16651);
nand U22633 (N_22633,N_17842,N_15415);
nor U22634 (N_22634,N_16986,N_16831);
and U22635 (N_22635,N_17024,N_16898);
nand U22636 (N_22636,N_18091,N_17654);
xnor U22637 (N_22637,N_19325,N_19725);
nand U22638 (N_22638,N_19301,N_19182);
nand U22639 (N_22639,N_19547,N_15104);
nor U22640 (N_22640,N_16471,N_16056);
xnor U22641 (N_22641,N_17817,N_16305);
nor U22642 (N_22642,N_18823,N_16630);
nor U22643 (N_22643,N_16358,N_19927);
and U22644 (N_22644,N_19911,N_19277);
or U22645 (N_22645,N_18034,N_18311);
and U22646 (N_22646,N_16584,N_19732);
nor U22647 (N_22647,N_15480,N_15501);
nand U22648 (N_22648,N_17834,N_18447);
or U22649 (N_22649,N_17765,N_19541);
and U22650 (N_22650,N_16909,N_19615);
nor U22651 (N_22651,N_17997,N_17338);
or U22652 (N_22652,N_17514,N_15817);
nand U22653 (N_22653,N_15433,N_18725);
and U22654 (N_22654,N_15917,N_18475);
nand U22655 (N_22655,N_16385,N_18979);
nor U22656 (N_22656,N_17490,N_15066);
xor U22657 (N_22657,N_17785,N_17172);
nor U22658 (N_22658,N_16193,N_16367);
xor U22659 (N_22659,N_17048,N_15519);
or U22660 (N_22660,N_19200,N_19886);
nor U22661 (N_22661,N_16845,N_18748);
xor U22662 (N_22662,N_17013,N_15185);
or U22663 (N_22663,N_15536,N_18038);
nand U22664 (N_22664,N_19334,N_16290);
nor U22665 (N_22665,N_17916,N_17563);
or U22666 (N_22666,N_19480,N_19507);
nand U22667 (N_22667,N_18963,N_16067);
or U22668 (N_22668,N_17287,N_15462);
and U22669 (N_22669,N_18214,N_18550);
or U22670 (N_22670,N_15194,N_16085);
or U22671 (N_22671,N_17702,N_19861);
xnor U22672 (N_22672,N_17715,N_17322);
nand U22673 (N_22673,N_16791,N_15118);
nand U22674 (N_22674,N_16347,N_17895);
or U22675 (N_22675,N_18620,N_17912);
and U22676 (N_22676,N_16382,N_17005);
xor U22677 (N_22677,N_18317,N_19308);
and U22678 (N_22678,N_18446,N_16529);
nand U22679 (N_22679,N_18954,N_19603);
and U22680 (N_22680,N_18519,N_16663);
nor U22681 (N_22681,N_16176,N_18008);
nor U22682 (N_22682,N_17855,N_18538);
and U22683 (N_22683,N_18177,N_15740);
nand U22684 (N_22684,N_19810,N_17122);
or U22685 (N_22685,N_16835,N_16576);
nand U22686 (N_22686,N_18689,N_15523);
nor U22687 (N_22687,N_18473,N_16235);
and U22688 (N_22688,N_15465,N_19406);
and U22689 (N_22689,N_18135,N_16811);
or U22690 (N_22690,N_16043,N_18908);
and U22691 (N_22691,N_16093,N_15390);
nor U22692 (N_22692,N_17761,N_18588);
xnor U22693 (N_22693,N_18238,N_16942);
and U22694 (N_22694,N_18856,N_16883);
or U22695 (N_22695,N_17249,N_15023);
xor U22696 (N_22696,N_18310,N_17334);
nand U22697 (N_22697,N_16505,N_16338);
or U22698 (N_22698,N_15287,N_17379);
nand U22699 (N_22699,N_18160,N_18559);
nor U22700 (N_22700,N_16670,N_16336);
nor U22701 (N_22701,N_17224,N_19278);
and U22702 (N_22702,N_17375,N_15119);
and U22703 (N_22703,N_17101,N_18136);
nand U22704 (N_22704,N_15602,N_15677);
and U22705 (N_22705,N_16192,N_16116);
nor U22706 (N_22706,N_15471,N_18728);
or U22707 (N_22707,N_15578,N_15085);
and U22708 (N_22708,N_18865,N_16155);
nand U22709 (N_22709,N_19075,N_18500);
or U22710 (N_22710,N_18730,N_18503);
or U22711 (N_22711,N_17238,N_17375);
and U22712 (N_22712,N_16172,N_16489);
xnor U22713 (N_22713,N_17655,N_19386);
or U22714 (N_22714,N_19053,N_17934);
nor U22715 (N_22715,N_17675,N_18259);
nor U22716 (N_22716,N_18502,N_16072);
and U22717 (N_22717,N_16232,N_17612);
nand U22718 (N_22718,N_18346,N_18374);
xnor U22719 (N_22719,N_17572,N_18198);
nand U22720 (N_22720,N_16478,N_15220);
and U22721 (N_22721,N_17825,N_19243);
or U22722 (N_22722,N_16910,N_16448);
nand U22723 (N_22723,N_17363,N_19376);
nand U22724 (N_22724,N_19709,N_15458);
nor U22725 (N_22725,N_19247,N_19180);
nor U22726 (N_22726,N_16219,N_15234);
and U22727 (N_22727,N_17584,N_17538);
nand U22728 (N_22728,N_19760,N_16478);
and U22729 (N_22729,N_18930,N_18112);
xnor U22730 (N_22730,N_15893,N_15880);
nand U22731 (N_22731,N_16634,N_16835);
nand U22732 (N_22732,N_19952,N_17905);
nor U22733 (N_22733,N_19248,N_16758);
nand U22734 (N_22734,N_18025,N_16322);
xor U22735 (N_22735,N_16024,N_17081);
and U22736 (N_22736,N_15143,N_17704);
and U22737 (N_22737,N_19800,N_15777);
xor U22738 (N_22738,N_16088,N_17309);
nand U22739 (N_22739,N_18751,N_16523);
or U22740 (N_22740,N_15236,N_15286);
or U22741 (N_22741,N_17269,N_18373);
and U22742 (N_22742,N_19379,N_18355);
and U22743 (N_22743,N_15669,N_18777);
nand U22744 (N_22744,N_18212,N_15791);
and U22745 (N_22745,N_16344,N_16163);
or U22746 (N_22746,N_18042,N_19224);
or U22747 (N_22747,N_17715,N_15327);
and U22748 (N_22748,N_18663,N_18019);
nor U22749 (N_22749,N_17632,N_19000);
or U22750 (N_22750,N_19340,N_16180);
nor U22751 (N_22751,N_19688,N_19155);
xnor U22752 (N_22752,N_19166,N_17535);
or U22753 (N_22753,N_15892,N_18290);
or U22754 (N_22754,N_16543,N_19267);
or U22755 (N_22755,N_15723,N_15561);
or U22756 (N_22756,N_17167,N_16750);
xor U22757 (N_22757,N_15950,N_19838);
nand U22758 (N_22758,N_16219,N_19161);
nor U22759 (N_22759,N_15940,N_18360);
or U22760 (N_22760,N_19893,N_19743);
xnor U22761 (N_22761,N_16071,N_16138);
or U22762 (N_22762,N_17115,N_19231);
xor U22763 (N_22763,N_16083,N_15769);
or U22764 (N_22764,N_18083,N_17281);
and U22765 (N_22765,N_16689,N_19589);
xnor U22766 (N_22766,N_17820,N_15621);
nor U22767 (N_22767,N_15141,N_15987);
xnor U22768 (N_22768,N_19230,N_19295);
nand U22769 (N_22769,N_16589,N_16039);
or U22770 (N_22770,N_19768,N_18769);
xnor U22771 (N_22771,N_17657,N_17989);
nand U22772 (N_22772,N_15184,N_18366);
and U22773 (N_22773,N_17887,N_18153);
nor U22774 (N_22774,N_15443,N_18804);
xor U22775 (N_22775,N_16348,N_19978);
nor U22776 (N_22776,N_19768,N_18171);
nand U22777 (N_22777,N_15787,N_17908);
nand U22778 (N_22778,N_18828,N_19718);
xor U22779 (N_22779,N_15606,N_19567);
xor U22780 (N_22780,N_16070,N_15685);
and U22781 (N_22781,N_16734,N_15524);
nand U22782 (N_22782,N_16528,N_16148);
nand U22783 (N_22783,N_16791,N_15440);
xnor U22784 (N_22784,N_18783,N_18952);
xor U22785 (N_22785,N_15958,N_18097);
nor U22786 (N_22786,N_18551,N_17942);
or U22787 (N_22787,N_18807,N_19241);
or U22788 (N_22788,N_15683,N_17114);
and U22789 (N_22789,N_15746,N_18680);
xnor U22790 (N_22790,N_17944,N_16502);
nand U22791 (N_22791,N_16884,N_19411);
and U22792 (N_22792,N_15971,N_19221);
xnor U22793 (N_22793,N_15683,N_18218);
xor U22794 (N_22794,N_17095,N_16717);
nor U22795 (N_22795,N_16686,N_18850);
or U22796 (N_22796,N_18263,N_19423);
and U22797 (N_22797,N_16084,N_16276);
nor U22798 (N_22798,N_19429,N_16624);
nand U22799 (N_22799,N_18909,N_18284);
or U22800 (N_22800,N_19319,N_19734);
or U22801 (N_22801,N_15556,N_19046);
nor U22802 (N_22802,N_19874,N_17950);
nor U22803 (N_22803,N_16178,N_15323);
nand U22804 (N_22804,N_17098,N_18880);
nor U22805 (N_22805,N_17761,N_16136);
xnor U22806 (N_22806,N_15070,N_15607);
or U22807 (N_22807,N_15177,N_18226);
and U22808 (N_22808,N_16154,N_19690);
nor U22809 (N_22809,N_15147,N_16652);
nor U22810 (N_22810,N_15200,N_17250);
and U22811 (N_22811,N_17274,N_18931);
or U22812 (N_22812,N_15290,N_18102);
or U22813 (N_22813,N_15482,N_17228);
xor U22814 (N_22814,N_16745,N_16873);
xnor U22815 (N_22815,N_16430,N_19942);
nand U22816 (N_22816,N_19579,N_15193);
nand U22817 (N_22817,N_16706,N_18424);
nor U22818 (N_22818,N_16202,N_18740);
and U22819 (N_22819,N_19283,N_15363);
or U22820 (N_22820,N_18648,N_17519);
nor U22821 (N_22821,N_19148,N_19466);
xnor U22822 (N_22822,N_19606,N_19624);
nor U22823 (N_22823,N_15534,N_17068);
nand U22824 (N_22824,N_15029,N_15177);
nor U22825 (N_22825,N_17916,N_17697);
nor U22826 (N_22826,N_18421,N_18362);
nand U22827 (N_22827,N_15579,N_19641);
nor U22828 (N_22828,N_15295,N_18668);
nand U22829 (N_22829,N_17040,N_16927);
nand U22830 (N_22830,N_16301,N_18053);
xor U22831 (N_22831,N_19156,N_17688);
nand U22832 (N_22832,N_19882,N_15044);
xor U22833 (N_22833,N_18654,N_15300);
nand U22834 (N_22834,N_15863,N_15740);
xnor U22835 (N_22835,N_17695,N_19741);
xor U22836 (N_22836,N_16809,N_16648);
or U22837 (N_22837,N_15245,N_18861);
and U22838 (N_22838,N_15406,N_16585);
nand U22839 (N_22839,N_16751,N_19364);
and U22840 (N_22840,N_19088,N_18867);
and U22841 (N_22841,N_19455,N_15311);
nand U22842 (N_22842,N_18371,N_19824);
and U22843 (N_22843,N_15252,N_19552);
nor U22844 (N_22844,N_17781,N_18265);
nand U22845 (N_22845,N_15897,N_15314);
or U22846 (N_22846,N_17469,N_17288);
nor U22847 (N_22847,N_18404,N_16865);
nand U22848 (N_22848,N_19679,N_18989);
xor U22849 (N_22849,N_19270,N_18853);
or U22850 (N_22850,N_19956,N_19297);
or U22851 (N_22851,N_18457,N_19640);
and U22852 (N_22852,N_17070,N_18335);
xnor U22853 (N_22853,N_18199,N_16513);
or U22854 (N_22854,N_18225,N_19301);
and U22855 (N_22855,N_19870,N_18957);
and U22856 (N_22856,N_16290,N_17160);
nand U22857 (N_22857,N_18568,N_18056);
nand U22858 (N_22858,N_19395,N_18586);
and U22859 (N_22859,N_15189,N_18504);
and U22860 (N_22860,N_19790,N_18528);
nor U22861 (N_22861,N_18742,N_19884);
nor U22862 (N_22862,N_18366,N_19916);
nand U22863 (N_22863,N_17134,N_18739);
nor U22864 (N_22864,N_19508,N_19551);
and U22865 (N_22865,N_19074,N_15119);
xor U22866 (N_22866,N_16608,N_16958);
and U22867 (N_22867,N_15390,N_18760);
and U22868 (N_22868,N_16780,N_15633);
and U22869 (N_22869,N_19183,N_17251);
and U22870 (N_22870,N_15993,N_18480);
or U22871 (N_22871,N_19136,N_19792);
nand U22872 (N_22872,N_19988,N_19838);
and U22873 (N_22873,N_15131,N_16744);
nand U22874 (N_22874,N_17016,N_17332);
or U22875 (N_22875,N_16908,N_17151);
and U22876 (N_22876,N_17710,N_16380);
or U22877 (N_22877,N_18792,N_17971);
nor U22878 (N_22878,N_15195,N_17960);
xor U22879 (N_22879,N_19237,N_16825);
nor U22880 (N_22880,N_17725,N_16913);
xor U22881 (N_22881,N_15596,N_19598);
xor U22882 (N_22882,N_15444,N_19911);
and U22883 (N_22883,N_19844,N_17262);
and U22884 (N_22884,N_16250,N_18246);
and U22885 (N_22885,N_17661,N_17399);
xnor U22886 (N_22886,N_18492,N_16472);
xnor U22887 (N_22887,N_15014,N_19300);
nand U22888 (N_22888,N_18070,N_19663);
and U22889 (N_22889,N_17671,N_17424);
nand U22890 (N_22890,N_18950,N_17231);
xor U22891 (N_22891,N_19989,N_17396);
and U22892 (N_22892,N_17493,N_19639);
nand U22893 (N_22893,N_18397,N_19059);
or U22894 (N_22894,N_15479,N_17575);
xor U22895 (N_22895,N_18292,N_18562);
xnor U22896 (N_22896,N_15124,N_18383);
xor U22897 (N_22897,N_18269,N_17778);
nand U22898 (N_22898,N_16690,N_15220);
xor U22899 (N_22899,N_18514,N_17349);
xnor U22900 (N_22900,N_19708,N_18407);
xor U22901 (N_22901,N_18149,N_18129);
nor U22902 (N_22902,N_15040,N_19550);
and U22903 (N_22903,N_15802,N_18470);
and U22904 (N_22904,N_19324,N_19294);
and U22905 (N_22905,N_19120,N_17432);
nor U22906 (N_22906,N_19201,N_19417);
nor U22907 (N_22907,N_19083,N_15523);
nor U22908 (N_22908,N_17365,N_15950);
or U22909 (N_22909,N_16480,N_15356);
nor U22910 (N_22910,N_16384,N_16077);
nand U22911 (N_22911,N_15916,N_15884);
and U22912 (N_22912,N_18940,N_15773);
or U22913 (N_22913,N_16608,N_16752);
xor U22914 (N_22914,N_16973,N_19528);
or U22915 (N_22915,N_16382,N_18437);
xnor U22916 (N_22916,N_18145,N_16363);
and U22917 (N_22917,N_19391,N_16038);
or U22918 (N_22918,N_16821,N_19047);
xnor U22919 (N_22919,N_19645,N_18044);
xnor U22920 (N_22920,N_19727,N_16453);
nand U22921 (N_22921,N_19119,N_15480);
or U22922 (N_22922,N_18113,N_18937);
and U22923 (N_22923,N_17955,N_17741);
nand U22924 (N_22924,N_17901,N_18799);
nand U22925 (N_22925,N_18162,N_17587);
xor U22926 (N_22926,N_18394,N_16956);
and U22927 (N_22927,N_16973,N_19588);
nand U22928 (N_22928,N_18995,N_19583);
nor U22929 (N_22929,N_17808,N_16819);
xnor U22930 (N_22930,N_15028,N_15555);
nand U22931 (N_22931,N_17087,N_18141);
or U22932 (N_22932,N_18393,N_17381);
xor U22933 (N_22933,N_16159,N_16459);
xor U22934 (N_22934,N_17969,N_17089);
and U22935 (N_22935,N_18473,N_18206);
nand U22936 (N_22936,N_19724,N_17692);
xor U22937 (N_22937,N_16098,N_16499);
or U22938 (N_22938,N_15823,N_16605);
xor U22939 (N_22939,N_19403,N_17755);
nand U22940 (N_22940,N_16128,N_16731);
or U22941 (N_22941,N_16476,N_17321);
or U22942 (N_22942,N_19378,N_19588);
nor U22943 (N_22943,N_17230,N_19915);
and U22944 (N_22944,N_15349,N_16764);
or U22945 (N_22945,N_19481,N_16827);
and U22946 (N_22946,N_17920,N_19099);
nand U22947 (N_22947,N_15051,N_19445);
nor U22948 (N_22948,N_17717,N_18452);
xnor U22949 (N_22949,N_18868,N_15731);
nand U22950 (N_22950,N_15656,N_16119);
and U22951 (N_22951,N_17749,N_15931);
nand U22952 (N_22952,N_18070,N_19648);
or U22953 (N_22953,N_16019,N_18393);
xor U22954 (N_22954,N_17738,N_16252);
or U22955 (N_22955,N_19527,N_18332);
or U22956 (N_22956,N_15475,N_15764);
or U22957 (N_22957,N_15257,N_19280);
or U22958 (N_22958,N_18342,N_19677);
nand U22959 (N_22959,N_15070,N_15531);
nor U22960 (N_22960,N_18394,N_19159);
nand U22961 (N_22961,N_18770,N_18338);
xnor U22962 (N_22962,N_17963,N_19154);
nor U22963 (N_22963,N_16350,N_16293);
xor U22964 (N_22964,N_19569,N_15718);
nand U22965 (N_22965,N_15314,N_16867);
xor U22966 (N_22966,N_18873,N_17791);
nand U22967 (N_22967,N_16008,N_19339);
nand U22968 (N_22968,N_15979,N_17422);
nand U22969 (N_22969,N_18313,N_15221);
or U22970 (N_22970,N_17297,N_19175);
nand U22971 (N_22971,N_18046,N_17184);
and U22972 (N_22972,N_18681,N_16693);
xnor U22973 (N_22973,N_19335,N_16216);
or U22974 (N_22974,N_18957,N_18726);
nor U22975 (N_22975,N_16263,N_19742);
nor U22976 (N_22976,N_17817,N_18418);
nor U22977 (N_22977,N_16912,N_18019);
or U22978 (N_22978,N_16549,N_17990);
nand U22979 (N_22979,N_19497,N_15536);
and U22980 (N_22980,N_19911,N_15696);
nor U22981 (N_22981,N_19282,N_16010);
or U22982 (N_22982,N_17193,N_17570);
xnor U22983 (N_22983,N_19275,N_15392);
xnor U22984 (N_22984,N_18797,N_18610);
and U22985 (N_22985,N_19720,N_16085);
nor U22986 (N_22986,N_17616,N_16535);
or U22987 (N_22987,N_19153,N_19948);
and U22988 (N_22988,N_19483,N_15705);
nor U22989 (N_22989,N_15821,N_17551);
or U22990 (N_22990,N_18254,N_15811);
or U22991 (N_22991,N_17134,N_15096);
nand U22992 (N_22992,N_18970,N_19565);
nor U22993 (N_22993,N_16712,N_15537);
and U22994 (N_22994,N_17517,N_15640);
xor U22995 (N_22995,N_18272,N_18076);
nor U22996 (N_22996,N_17648,N_16312);
xor U22997 (N_22997,N_19113,N_16585);
and U22998 (N_22998,N_19057,N_19921);
or U22999 (N_22999,N_16465,N_19993);
and U23000 (N_23000,N_19655,N_17089);
or U23001 (N_23001,N_17229,N_19846);
xnor U23002 (N_23002,N_15351,N_18487);
nor U23003 (N_23003,N_17066,N_16886);
nor U23004 (N_23004,N_17051,N_18605);
and U23005 (N_23005,N_16341,N_17072);
and U23006 (N_23006,N_17186,N_19358);
xnor U23007 (N_23007,N_16328,N_18028);
or U23008 (N_23008,N_16198,N_17836);
and U23009 (N_23009,N_18307,N_19538);
xor U23010 (N_23010,N_16754,N_19865);
xor U23011 (N_23011,N_19476,N_19460);
xnor U23012 (N_23012,N_17321,N_16967);
xor U23013 (N_23013,N_15417,N_15476);
xnor U23014 (N_23014,N_16608,N_16704);
or U23015 (N_23015,N_19109,N_19305);
or U23016 (N_23016,N_15098,N_18082);
xnor U23017 (N_23017,N_18540,N_16499);
nand U23018 (N_23018,N_15307,N_15198);
nand U23019 (N_23019,N_17068,N_18239);
or U23020 (N_23020,N_16758,N_17547);
xnor U23021 (N_23021,N_18057,N_17614);
nor U23022 (N_23022,N_19210,N_15467);
and U23023 (N_23023,N_15775,N_17917);
nand U23024 (N_23024,N_18577,N_18586);
nor U23025 (N_23025,N_16166,N_15833);
xnor U23026 (N_23026,N_17662,N_19779);
xor U23027 (N_23027,N_18999,N_19464);
nor U23028 (N_23028,N_18540,N_18735);
xnor U23029 (N_23029,N_15411,N_17533);
and U23030 (N_23030,N_15568,N_18940);
and U23031 (N_23031,N_17386,N_15933);
nor U23032 (N_23032,N_15083,N_15924);
and U23033 (N_23033,N_15212,N_17284);
and U23034 (N_23034,N_16394,N_15096);
nand U23035 (N_23035,N_17625,N_18695);
xor U23036 (N_23036,N_18937,N_16063);
and U23037 (N_23037,N_18788,N_19100);
and U23038 (N_23038,N_15657,N_15174);
xnor U23039 (N_23039,N_19636,N_16547);
nor U23040 (N_23040,N_19827,N_16294);
nand U23041 (N_23041,N_18241,N_15140);
xor U23042 (N_23042,N_16222,N_16292);
nand U23043 (N_23043,N_19787,N_19521);
or U23044 (N_23044,N_17841,N_19656);
or U23045 (N_23045,N_16386,N_15216);
xor U23046 (N_23046,N_16879,N_17185);
or U23047 (N_23047,N_15326,N_15426);
nand U23048 (N_23048,N_16101,N_15688);
nand U23049 (N_23049,N_15409,N_16615);
and U23050 (N_23050,N_19419,N_19534);
nor U23051 (N_23051,N_15857,N_17641);
or U23052 (N_23052,N_15141,N_17890);
and U23053 (N_23053,N_16339,N_19620);
nor U23054 (N_23054,N_16882,N_18796);
or U23055 (N_23055,N_19883,N_15417);
xnor U23056 (N_23056,N_17391,N_19998);
xnor U23057 (N_23057,N_15920,N_19872);
xnor U23058 (N_23058,N_17002,N_15023);
nor U23059 (N_23059,N_17914,N_17850);
nor U23060 (N_23060,N_18574,N_18052);
and U23061 (N_23061,N_19522,N_19669);
nor U23062 (N_23062,N_16013,N_19277);
xnor U23063 (N_23063,N_19858,N_18770);
xor U23064 (N_23064,N_17870,N_16828);
nor U23065 (N_23065,N_18470,N_17017);
xnor U23066 (N_23066,N_18114,N_19124);
or U23067 (N_23067,N_17003,N_16748);
xnor U23068 (N_23068,N_16641,N_16725);
nand U23069 (N_23069,N_15124,N_17951);
xor U23070 (N_23070,N_18298,N_19722);
or U23071 (N_23071,N_18971,N_17508);
nand U23072 (N_23072,N_17168,N_19765);
nor U23073 (N_23073,N_19331,N_16788);
or U23074 (N_23074,N_15985,N_18345);
xor U23075 (N_23075,N_15090,N_17504);
nand U23076 (N_23076,N_18744,N_17557);
nor U23077 (N_23077,N_16619,N_19795);
and U23078 (N_23078,N_18147,N_18510);
and U23079 (N_23079,N_19426,N_16081);
xnor U23080 (N_23080,N_17205,N_19841);
and U23081 (N_23081,N_18626,N_16199);
or U23082 (N_23082,N_16374,N_15693);
xor U23083 (N_23083,N_17334,N_19895);
or U23084 (N_23084,N_18723,N_16267);
and U23085 (N_23085,N_19051,N_16386);
xor U23086 (N_23086,N_15055,N_16328);
or U23087 (N_23087,N_17064,N_16243);
or U23088 (N_23088,N_15906,N_16809);
nor U23089 (N_23089,N_15531,N_17332);
nand U23090 (N_23090,N_18574,N_19400);
nor U23091 (N_23091,N_17376,N_16547);
xor U23092 (N_23092,N_18893,N_15357);
nand U23093 (N_23093,N_17509,N_19684);
or U23094 (N_23094,N_18045,N_15736);
xnor U23095 (N_23095,N_19996,N_15800);
xor U23096 (N_23096,N_16070,N_16948);
nor U23097 (N_23097,N_18013,N_19719);
xor U23098 (N_23098,N_19758,N_18285);
nor U23099 (N_23099,N_16972,N_17549);
or U23100 (N_23100,N_18273,N_17318);
xnor U23101 (N_23101,N_17227,N_15069);
xnor U23102 (N_23102,N_15817,N_15910);
xnor U23103 (N_23103,N_17875,N_19677);
xnor U23104 (N_23104,N_16124,N_16963);
xnor U23105 (N_23105,N_18655,N_18576);
nor U23106 (N_23106,N_17830,N_16752);
xor U23107 (N_23107,N_17058,N_18239);
xnor U23108 (N_23108,N_17715,N_16509);
xor U23109 (N_23109,N_17308,N_18579);
and U23110 (N_23110,N_19525,N_15560);
xnor U23111 (N_23111,N_16868,N_17289);
xnor U23112 (N_23112,N_17684,N_16138);
and U23113 (N_23113,N_16388,N_18829);
and U23114 (N_23114,N_19343,N_16473);
xnor U23115 (N_23115,N_16093,N_18622);
nor U23116 (N_23116,N_17261,N_16783);
or U23117 (N_23117,N_15139,N_17671);
or U23118 (N_23118,N_15428,N_15172);
nand U23119 (N_23119,N_16111,N_15045);
nor U23120 (N_23120,N_15137,N_18600);
or U23121 (N_23121,N_19909,N_18017);
nand U23122 (N_23122,N_16859,N_16310);
or U23123 (N_23123,N_18222,N_16792);
and U23124 (N_23124,N_15741,N_16777);
xnor U23125 (N_23125,N_19612,N_17093);
or U23126 (N_23126,N_15362,N_15196);
nand U23127 (N_23127,N_16374,N_18928);
and U23128 (N_23128,N_15831,N_15311);
nor U23129 (N_23129,N_19445,N_15434);
xor U23130 (N_23130,N_17822,N_15403);
or U23131 (N_23131,N_15434,N_16751);
and U23132 (N_23132,N_18866,N_16014);
or U23133 (N_23133,N_15777,N_18446);
xor U23134 (N_23134,N_16833,N_16501);
nor U23135 (N_23135,N_16823,N_16715);
xnor U23136 (N_23136,N_18452,N_16179);
and U23137 (N_23137,N_16453,N_16248);
xor U23138 (N_23138,N_19653,N_15470);
nand U23139 (N_23139,N_15679,N_18628);
nor U23140 (N_23140,N_18899,N_15556);
nand U23141 (N_23141,N_19082,N_18794);
and U23142 (N_23142,N_18180,N_18176);
nand U23143 (N_23143,N_18318,N_19708);
or U23144 (N_23144,N_19891,N_19832);
or U23145 (N_23145,N_19055,N_17426);
nand U23146 (N_23146,N_15284,N_19182);
nor U23147 (N_23147,N_18971,N_16423);
or U23148 (N_23148,N_18769,N_16741);
nand U23149 (N_23149,N_15614,N_17613);
xor U23150 (N_23150,N_16108,N_19966);
nand U23151 (N_23151,N_17105,N_16735);
nor U23152 (N_23152,N_18356,N_18333);
nand U23153 (N_23153,N_15216,N_19718);
and U23154 (N_23154,N_15035,N_19740);
and U23155 (N_23155,N_17440,N_15364);
and U23156 (N_23156,N_18051,N_16452);
nor U23157 (N_23157,N_18425,N_16668);
nor U23158 (N_23158,N_15841,N_15487);
nor U23159 (N_23159,N_17910,N_18036);
and U23160 (N_23160,N_15748,N_18244);
xnor U23161 (N_23161,N_15568,N_17016);
xnor U23162 (N_23162,N_17382,N_18353);
or U23163 (N_23163,N_16885,N_16703);
nor U23164 (N_23164,N_19250,N_16318);
xnor U23165 (N_23165,N_18559,N_16314);
or U23166 (N_23166,N_16102,N_15402);
nor U23167 (N_23167,N_19875,N_18825);
xor U23168 (N_23168,N_18213,N_17856);
nand U23169 (N_23169,N_17902,N_16526);
nand U23170 (N_23170,N_19587,N_17190);
and U23171 (N_23171,N_15854,N_18812);
or U23172 (N_23172,N_18208,N_16469);
or U23173 (N_23173,N_18892,N_19752);
or U23174 (N_23174,N_19677,N_15901);
xor U23175 (N_23175,N_16819,N_17882);
or U23176 (N_23176,N_17044,N_18740);
xnor U23177 (N_23177,N_17724,N_17468);
xnor U23178 (N_23178,N_17344,N_16148);
or U23179 (N_23179,N_18912,N_16483);
xnor U23180 (N_23180,N_17372,N_15818);
nand U23181 (N_23181,N_15092,N_15882);
nand U23182 (N_23182,N_15579,N_18244);
xnor U23183 (N_23183,N_15980,N_19340);
xor U23184 (N_23184,N_19218,N_19879);
or U23185 (N_23185,N_18539,N_18321);
nor U23186 (N_23186,N_15363,N_16407);
xnor U23187 (N_23187,N_19413,N_16027);
nand U23188 (N_23188,N_15702,N_15626);
or U23189 (N_23189,N_17383,N_19790);
nor U23190 (N_23190,N_18626,N_17300);
nor U23191 (N_23191,N_16726,N_19187);
nor U23192 (N_23192,N_16224,N_17951);
nand U23193 (N_23193,N_17424,N_19070);
nand U23194 (N_23194,N_15749,N_19064);
nand U23195 (N_23195,N_15890,N_17395);
nand U23196 (N_23196,N_17664,N_17296);
and U23197 (N_23197,N_16067,N_19684);
xnor U23198 (N_23198,N_18799,N_15184);
and U23199 (N_23199,N_17643,N_18044);
xnor U23200 (N_23200,N_17197,N_15413);
nand U23201 (N_23201,N_15880,N_19041);
nand U23202 (N_23202,N_16345,N_18835);
or U23203 (N_23203,N_18968,N_16164);
nor U23204 (N_23204,N_15495,N_16845);
and U23205 (N_23205,N_18588,N_18441);
xnor U23206 (N_23206,N_15330,N_18291);
nor U23207 (N_23207,N_15116,N_19680);
xor U23208 (N_23208,N_18237,N_18954);
or U23209 (N_23209,N_18991,N_15325);
nand U23210 (N_23210,N_18936,N_17827);
and U23211 (N_23211,N_15096,N_16280);
and U23212 (N_23212,N_16872,N_18831);
nand U23213 (N_23213,N_18052,N_16949);
or U23214 (N_23214,N_19862,N_15388);
xnor U23215 (N_23215,N_17320,N_16555);
nand U23216 (N_23216,N_16742,N_17328);
and U23217 (N_23217,N_16570,N_15096);
or U23218 (N_23218,N_18552,N_18192);
and U23219 (N_23219,N_16252,N_17982);
nand U23220 (N_23220,N_17953,N_19120);
nand U23221 (N_23221,N_19496,N_16741);
or U23222 (N_23222,N_19606,N_18518);
nor U23223 (N_23223,N_18155,N_15047);
and U23224 (N_23224,N_19502,N_17273);
and U23225 (N_23225,N_16733,N_15771);
nand U23226 (N_23226,N_17522,N_16199);
and U23227 (N_23227,N_19138,N_19820);
and U23228 (N_23228,N_15853,N_17695);
nand U23229 (N_23229,N_19023,N_18349);
nor U23230 (N_23230,N_15793,N_15739);
xnor U23231 (N_23231,N_18143,N_15767);
nand U23232 (N_23232,N_18182,N_16383);
xnor U23233 (N_23233,N_16733,N_15410);
or U23234 (N_23234,N_18562,N_19248);
and U23235 (N_23235,N_15925,N_15014);
xor U23236 (N_23236,N_18470,N_19912);
xnor U23237 (N_23237,N_15879,N_16057);
or U23238 (N_23238,N_16309,N_15337);
nand U23239 (N_23239,N_15253,N_16769);
and U23240 (N_23240,N_19964,N_18572);
and U23241 (N_23241,N_18539,N_19867);
nor U23242 (N_23242,N_16408,N_19528);
or U23243 (N_23243,N_18191,N_19558);
and U23244 (N_23244,N_18773,N_17505);
nand U23245 (N_23245,N_19755,N_18541);
and U23246 (N_23246,N_15769,N_15033);
xor U23247 (N_23247,N_18736,N_16085);
nand U23248 (N_23248,N_17586,N_15983);
or U23249 (N_23249,N_18401,N_15626);
nor U23250 (N_23250,N_15557,N_19307);
and U23251 (N_23251,N_15375,N_18953);
xnor U23252 (N_23252,N_18956,N_17622);
xnor U23253 (N_23253,N_15721,N_15227);
nor U23254 (N_23254,N_19052,N_15755);
or U23255 (N_23255,N_16027,N_17819);
xnor U23256 (N_23256,N_16479,N_18807);
and U23257 (N_23257,N_19602,N_18017);
nand U23258 (N_23258,N_18056,N_17013);
and U23259 (N_23259,N_17332,N_19893);
nor U23260 (N_23260,N_18852,N_18946);
nor U23261 (N_23261,N_16588,N_19669);
xor U23262 (N_23262,N_19337,N_19003);
nor U23263 (N_23263,N_15906,N_17013);
and U23264 (N_23264,N_18727,N_19670);
xor U23265 (N_23265,N_19246,N_19512);
nor U23266 (N_23266,N_16604,N_18459);
or U23267 (N_23267,N_15929,N_19619);
xor U23268 (N_23268,N_19449,N_17786);
xor U23269 (N_23269,N_18550,N_18244);
or U23270 (N_23270,N_16274,N_18464);
or U23271 (N_23271,N_17057,N_15515);
nor U23272 (N_23272,N_16092,N_19704);
and U23273 (N_23273,N_16901,N_19334);
nand U23274 (N_23274,N_15778,N_17764);
and U23275 (N_23275,N_18161,N_18453);
or U23276 (N_23276,N_18537,N_18327);
xnor U23277 (N_23277,N_16342,N_18048);
xnor U23278 (N_23278,N_19636,N_17489);
and U23279 (N_23279,N_17866,N_19166);
nor U23280 (N_23280,N_18782,N_17921);
nor U23281 (N_23281,N_18213,N_17211);
and U23282 (N_23282,N_17448,N_17235);
xnor U23283 (N_23283,N_16119,N_16104);
nor U23284 (N_23284,N_15039,N_17154);
or U23285 (N_23285,N_16813,N_16678);
nand U23286 (N_23286,N_17924,N_15110);
and U23287 (N_23287,N_19974,N_17252);
xor U23288 (N_23288,N_17157,N_16447);
nand U23289 (N_23289,N_17587,N_17922);
nand U23290 (N_23290,N_18015,N_18035);
nand U23291 (N_23291,N_16615,N_17569);
nor U23292 (N_23292,N_19001,N_16512);
and U23293 (N_23293,N_17082,N_19373);
xor U23294 (N_23294,N_17257,N_18204);
xor U23295 (N_23295,N_16092,N_15677);
and U23296 (N_23296,N_18422,N_15891);
nand U23297 (N_23297,N_17681,N_15333);
or U23298 (N_23298,N_16882,N_15293);
nand U23299 (N_23299,N_19666,N_19146);
xor U23300 (N_23300,N_19713,N_16551);
and U23301 (N_23301,N_15429,N_16823);
and U23302 (N_23302,N_18047,N_17745);
nor U23303 (N_23303,N_16677,N_17941);
xnor U23304 (N_23304,N_16691,N_15386);
nand U23305 (N_23305,N_17285,N_17834);
xor U23306 (N_23306,N_17326,N_16418);
or U23307 (N_23307,N_18615,N_19449);
nand U23308 (N_23308,N_17209,N_15726);
and U23309 (N_23309,N_19631,N_18409);
nor U23310 (N_23310,N_15434,N_17778);
nand U23311 (N_23311,N_19304,N_15193);
nor U23312 (N_23312,N_15361,N_15959);
nand U23313 (N_23313,N_16458,N_15825);
and U23314 (N_23314,N_17385,N_18761);
nor U23315 (N_23315,N_19920,N_16868);
nor U23316 (N_23316,N_15320,N_16039);
or U23317 (N_23317,N_18942,N_19397);
and U23318 (N_23318,N_15361,N_18270);
nand U23319 (N_23319,N_17139,N_18507);
or U23320 (N_23320,N_16352,N_15655);
xor U23321 (N_23321,N_16420,N_17829);
xor U23322 (N_23322,N_16078,N_17420);
nor U23323 (N_23323,N_18290,N_17681);
and U23324 (N_23324,N_17963,N_15631);
or U23325 (N_23325,N_15327,N_17459);
nor U23326 (N_23326,N_15492,N_17764);
or U23327 (N_23327,N_17969,N_15199);
xnor U23328 (N_23328,N_18159,N_19052);
or U23329 (N_23329,N_15575,N_16480);
or U23330 (N_23330,N_16571,N_19146);
and U23331 (N_23331,N_16735,N_15567);
or U23332 (N_23332,N_19973,N_17733);
xor U23333 (N_23333,N_16355,N_19198);
nor U23334 (N_23334,N_18096,N_15066);
xor U23335 (N_23335,N_16761,N_15016);
and U23336 (N_23336,N_15660,N_19049);
or U23337 (N_23337,N_17484,N_15422);
nand U23338 (N_23338,N_17521,N_17646);
xor U23339 (N_23339,N_19219,N_17030);
nor U23340 (N_23340,N_18130,N_15160);
nor U23341 (N_23341,N_16214,N_18650);
or U23342 (N_23342,N_18649,N_19562);
xnor U23343 (N_23343,N_18815,N_15593);
or U23344 (N_23344,N_19445,N_19420);
nor U23345 (N_23345,N_17890,N_19936);
nor U23346 (N_23346,N_16450,N_19130);
nand U23347 (N_23347,N_15097,N_16529);
and U23348 (N_23348,N_17305,N_15895);
or U23349 (N_23349,N_15876,N_18237);
nand U23350 (N_23350,N_19093,N_17179);
and U23351 (N_23351,N_17799,N_15697);
nand U23352 (N_23352,N_18956,N_15639);
and U23353 (N_23353,N_16220,N_16816);
xnor U23354 (N_23354,N_18122,N_15315);
xor U23355 (N_23355,N_15118,N_16127);
nor U23356 (N_23356,N_17276,N_18082);
and U23357 (N_23357,N_17609,N_16125);
nor U23358 (N_23358,N_18113,N_17324);
nand U23359 (N_23359,N_16896,N_19620);
and U23360 (N_23360,N_16932,N_16240);
and U23361 (N_23361,N_18061,N_15403);
nor U23362 (N_23362,N_16422,N_15294);
xor U23363 (N_23363,N_15914,N_15307);
xnor U23364 (N_23364,N_17287,N_15914);
or U23365 (N_23365,N_16822,N_17449);
or U23366 (N_23366,N_15996,N_19150);
nand U23367 (N_23367,N_15651,N_16136);
or U23368 (N_23368,N_15832,N_16399);
or U23369 (N_23369,N_17004,N_15200);
and U23370 (N_23370,N_18993,N_15242);
and U23371 (N_23371,N_16022,N_19708);
xnor U23372 (N_23372,N_15341,N_15855);
nand U23373 (N_23373,N_17372,N_19520);
or U23374 (N_23374,N_19020,N_17051);
nor U23375 (N_23375,N_18040,N_16367);
or U23376 (N_23376,N_18424,N_19027);
and U23377 (N_23377,N_18760,N_17714);
and U23378 (N_23378,N_18001,N_17906);
nor U23379 (N_23379,N_15039,N_18125);
or U23380 (N_23380,N_19772,N_19625);
or U23381 (N_23381,N_17252,N_17327);
nand U23382 (N_23382,N_17797,N_18372);
nor U23383 (N_23383,N_17233,N_16387);
nor U23384 (N_23384,N_18835,N_16481);
nand U23385 (N_23385,N_18375,N_17410);
and U23386 (N_23386,N_16184,N_19680);
nand U23387 (N_23387,N_16202,N_19382);
or U23388 (N_23388,N_15486,N_15757);
nand U23389 (N_23389,N_17959,N_18494);
and U23390 (N_23390,N_16634,N_15785);
xor U23391 (N_23391,N_17051,N_19699);
and U23392 (N_23392,N_18955,N_17587);
or U23393 (N_23393,N_17837,N_17871);
or U23394 (N_23394,N_17573,N_16230);
and U23395 (N_23395,N_18719,N_17928);
nor U23396 (N_23396,N_17129,N_16734);
or U23397 (N_23397,N_19447,N_17874);
nor U23398 (N_23398,N_19614,N_16438);
nor U23399 (N_23399,N_16327,N_19829);
and U23400 (N_23400,N_17713,N_15125);
nand U23401 (N_23401,N_19353,N_17153);
nor U23402 (N_23402,N_16300,N_17093);
nor U23403 (N_23403,N_15675,N_16261);
xnor U23404 (N_23404,N_18079,N_15817);
nand U23405 (N_23405,N_19548,N_15109);
or U23406 (N_23406,N_15858,N_19030);
xor U23407 (N_23407,N_17797,N_18223);
nor U23408 (N_23408,N_18731,N_15176);
nor U23409 (N_23409,N_18758,N_17754);
and U23410 (N_23410,N_19317,N_16341);
or U23411 (N_23411,N_18144,N_16700);
and U23412 (N_23412,N_18036,N_16156);
and U23413 (N_23413,N_17791,N_19839);
or U23414 (N_23414,N_16087,N_15805);
nand U23415 (N_23415,N_19006,N_15369);
nand U23416 (N_23416,N_19142,N_17533);
or U23417 (N_23417,N_18770,N_18914);
nor U23418 (N_23418,N_15403,N_15500);
nand U23419 (N_23419,N_19001,N_18191);
or U23420 (N_23420,N_19783,N_19086);
nand U23421 (N_23421,N_19631,N_18769);
xnor U23422 (N_23422,N_17140,N_19133);
or U23423 (N_23423,N_19844,N_15472);
and U23424 (N_23424,N_18679,N_19423);
xor U23425 (N_23425,N_15336,N_16131);
and U23426 (N_23426,N_17682,N_15114);
and U23427 (N_23427,N_16016,N_19684);
xor U23428 (N_23428,N_17255,N_15544);
nand U23429 (N_23429,N_19076,N_16486);
nand U23430 (N_23430,N_19998,N_19069);
or U23431 (N_23431,N_19037,N_18722);
nand U23432 (N_23432,N_15406,N_19571);
nor U23433 (N_23433,N_18990,N_18260);
nand U23434 (N_23434,N_18625,N_15189);
and U23435 (N_23435,N_19697,N_19424);
nand U23436 (N_23436,N_17762,N_18956);
nand U23437 (N_23437,N_18297,N_15417);
nand U23438 (N_23438,N_15426,N_15923);
and U23439 (N_23439,N_15227,N_19897);
nor U23440 (N_23440,N_18926,N_17180);
nand U23441 (N_23441,N_19465,N_15614);
xnor U23442 (N_23442,N_16006,N_17352);
nand U23443 (N_23443,N_17140,N_15632);
nand U23444 (N_23444,N_18093,N_17119);
nand U23445 (N_23445,N_18363,N_19794);
nor U23446 (N_23446,N_15967,N_19106);
and U23447 (N_23447,N_19312,N_18732);
xor U23448 (N_23448,N_19189,N_15387);
or U23449 (N_23449,N_17789,N_16832);
and U23450 (N_23450,N_18501,N_19026);
nor U23451 (N_23451,N_17257,N_16356);
nor U23452 (N_23452,N_18714,N_16248);
and U23453 (N_23453,N_18898,N_18234);
nor U23454 (N_23454,N_18807,N_18034);
nor U23455 (N_23455,N_15795,N_17805);
or U23456 (N_23456,N_19193,N_16443);
and U23457 (N_23457,N_17229,N_15517);
nor U23458 (N_23458,N_18884,N_18401);
xnor U23459 (N_23459,N_19866,N_18834);
xnor U23460 (N_23460,N_19762,N_17143);
nand U23461 (N_23461,N_18459,N_16841);
xor U23462 (N_23462,N_17226,N_18693);
and U23463 (N_23463,N_15347,N_18312);
xnor U23464 (N_23464,N_19405,N_19443);
or U23465 (N_23465,N_15027,N_18664);
or U23466 (N_23466,N_18288,N_17197);
nand U23467 (N_23467,N_19574,N_19223);
and U23468 (N_23468,N_19690,N_17360);
and U23469 (N_23469,N_16333,N_15815);
xnor U23470 (N_23470,N_19117,N_17666);
nand U23471 (N_23471,N_17913,N_17790);
nand U23472 (N_23472,N_15916,N_18731);
xor U23473 (N_23473,N_18516,N_16019);
xnor U23474 (N_23474,N_16909,N_17709);
xor U23475 (N_23475,N_18380,N_15924);
nand U23476 (N_23476,N_15691,N_16886);
and U23477 (N_23477,N_19034,N_17331);
nor U23478 (N_23478,N_17154,N_18469);
nand U23479 (N_23479,N_17306,N_15247);
or U23480 (N_23480,N_18704,N_19864);
or U23481 (N_23481,N_19456,N_16194);
xnor U23482 (N_23482,N_18938,N_16620);
xor U23483 (N_23483,N_17013,N_16671);
nor U23484 (N_23484,N_16125,N_15876);
and U23485 (N_23485,N_15865,N_19008);
xnor U23486 (N_23486,N_18935,N_19495);
nor U23487 (N_23487,N_15037,N_19964);
nor U23488 (N_23488,N_16522,N_16598);
nor U23489 (N_23489,N_18776,N_17178);
nor U23490 (N_23490,N_15389,N_16674);
nor U23491 (N_23491,N_15622,N_16080);
and U23492 (N_23492,N_18886,N_16697);
nor U23493 (N_23493,N_17626,N_16696);
nor U23494 (N_23494,N_16246,N_19175);
and U23495 (N_23495,N_18131,N_15430);
or U23496 (N_23496,N_15222,N_17374);
or U23497 (N_23497,N_19383,N_18856);
or U23498 (N_23498,N_15369,N_18528);
and U23499 (N_23499,N_18150,N_17075);
nand U23500 (N_23500,N_18455,N_19281);
xor U23501 (N_23501,N_16553,N_19492);
xor U23502 (N_23502,N_16957,N_16464);
or U23503 (N_23503,N_17721,N_18450);
or U23504 (N_23504,N_17047,N_16110);
xnor U23505 (N_23505,N_16385,N_15057);
nor U23506 (N_23506,N_19796,N_18047);
nor U23507 (N_23507,N_17636,N_19945);
xor U23508 (N_23508,N_15522,N_19801);
nor U23509 (N_23509,N_15103,N_16231);
xor U23510 (N_23510,N_18528,N_19350);
and U23511 (N_23511,N_17792,N_18833);
nor U23512 (N_23512,N_18294,N_17861);
and U23513 (N_23513,N_18283,N_19407);
or U23514 (N_23514,N_19593,N_18786);
nand U23515 (N_23515,N_19571,N_19154);
nor U23516 (N_23516,N_15061,N_16364);
nor U23517 (N_23517,N_17062,N_15232);
xor U23518 (N_23518,N_16182,N_15488);
nor U23519 (N_23519,N_16073,N_17830);
nand U23520 (N_23520,N_15544,N_17142);
nor U23521 (N_23521,N_19829,N_15368);
or U23522 (N_23522,N_18601,N_16984);
xor U23523 (N_23523,N_16708,N_17730);
xnor U23524 (N_23524,N_18842,N_16361);
and U23525 (N_23525,N_19980,N_15569);
and U23526 (N_23526,N_16016,N_15596);
xor U23527 (N_23527,N_16919,N_17218);
nand U23528 (N_23528,N_16565,N_18350);
nor U23529 (N_23529,N_19453,N_18503);
and U23530 (N_23530,N_15149,N_17278);
nor U23531 (N_23531,N_16910,N_17255);
and U23532 (N_23532,N_15559,N_15037);
nand U23533 (N_23533,N_16005,N_17643);
xnor U23534 (N_23534,N_15759,N_15566);
nand U23535 (N_23535,N_16105,N_17216);
nor U23536 (N_23536,N_18843,N_16452);
nor U23537 (N_23537,N_17150,N_16083);
nor U23538 (N_23538,N_17925,N_15626);
and U23539 (N_23539,N_16319,N_19381);
nor U23540 (N_23540,N_16351,N_17485);
xor U23541 (N_23541,N_17621,N_19153);
nor U23542 (N_23542,N_17511,N_16769);
nor U23543 (N_23543,N_17191,N_18515);
nand U23544 (N_23544,N_15773,N_15262);
nor U23545 (N_23545,N_16803,N_19704);
and U23546 (N_23546,N_15674,N_15983);
or U23547 (N_23547,N_16655,N_16584);
xor U23548 (N_23548,N_15139,N_18231);
nor U23549 (N_23549,N_15416,N_19861);
xnor U23550 (N_23550,N_19676,N_17667);
or U23551 (N_23551,N_19673,N_15524);
nor U23552 (N_23552,N_17305,N_16513);
or U23553 (N_23553,N_16082,N_16994);
nor U23554 (N_23554,N_19064,N_15118);
and U23555 (N_23555,N_19801,N_16286);
or U23556 (N_23556,N_17561,N_16337);
xor U23557 (N_23557,N_16250,N_18076);
nor U23558 (N_23558,N_17073,N_16598);
nand U23559 (N_23559,N_17082,N_15876);
or U23560 (N_23560,N_17554,N_16195);
xor U23561 (N_23561,N_18377,N_19159);
or U23562 (N_23562,N_19161,N_19330);
and U23563 (N_23563,N_16119,N_16163);
nand U23564 (N_23564,N_18379,N_17154);
and U23565 (N_23565,N_19709,N_18657);
nand U23566 (N_23566,N_18872,N_19357);
nor U23567 (N_23567,N_16981,N_15737);
xnor U23568 (N_23568,N_15625,N_19312);
xor U23569 (N_23569,N_15547,N_18748);
nand U23570 (N_23570,N_16154,N_16685);
or U23571 (N_23571,N_15632,N_15548);
xnor U23572 (N_23572,N_17955,N_19711);
or U23573 (N_23573,N_18102,N_18943);
and U23574 (N_23574,N_15765,N_19076);
xnor U23575 (N_23575,N_17188,N_15578);
and U23576 (N_23576,N_16423,N_17407);
or U23577 (N_23577,N_18243,N_18178);
nand U23578 (N_23578,N_18951,N_17458);
nand U23579 (N_23579,N_16216,N_17087);
xor U23580 (N_23580,N_17399,N_18587);
or U23581 (N_23581,N_15481,N_19234);
and U23582 (N_23582,N_17778,N_16228);
nand U23583 (N_23583,N_18408,N_17221);
nand U23584 (N_23584,N_18712,N_19959);
nor U23585 (N_23585,N_15456,N_15231);
xnor U23586 (N_23586,N_19932,N_16526);
or U23587 (N_23587,N_19921,N_18054);
or U23588 (N_23588,N_15285,N_16472);
xnor U23589 (N_23589,N_16602,N_19701);
or U23590 (N_23590,N_15428,N_18027);
nand U23591 (N_23591,N_16683,N_17889);
nor U23592 (N_23592,N_18171,N_15085);
nand U23593 (N_23593,N_15464,N_19094);
or U23594 (N_23594,N_19034,N_15457);
xor U23595 (N_23595,N_17472,N_18194);
or U23596 (N_23596,N_19788,N_19120);
or U23597 (N_23597,N_19728,N_19314);
nor U23598 (N_23598,N_18902,N_16218);
xor U23599 (N_23599,N_15224,N_17414);
nor U23600 (N_23600,N_19000,N_17464);
and U23601 (N_23601,N_19169,N_15798);
or U23602 (N_23602,N_19411,N_19226);
nand U23603 (N_23603,N_18093,N_19915);
and U23604 (N_23604,N_19627,N_17131);
nor U23605 (N_23605,N_16524,N_15528);
or U23606 (N_23606,N_17277,N_16444);
or U23607 (N_23607,N_18858,N_15091);
or U23608 (N_23608,N_19527,N_18122);
nor U23609 (N_23609,N_17852,N_17487);
or U23610 (N_23610,N_16100,N_16075);
and U23611 (N_23611,N_18916,N_19706);
and U23612 (N_23612,N_17731,N_16413);
nor U23613 (N_23613,N_19395,N_15883);
nor U23614 (N_23614,N_16595,N_15728);
nor U23615 (N_23615,N_17933,N_19469);
or U23616 (N_23616,N_17649,N_16959);
nand U23617 (N_23617,N_16212,N_17720);
nand U23618 (N_23618,N_17384,N_17423);
nor U23619 (N_23619,N_16796,N_17867);
nor U23620 (N_23620,N_16899,N_18307);
nor U23621 (N_23621,N_17921,N_18398);
or U23622 (N_23622,N_16197,N_18392);
nand U23623 (N_23623,N_17013,N_15878);
xnor U23624 (N_23624,N_16328,N_17393);
nor U23625 (N_23625,N_19647,N_18737);
nand U23626 (N_23626,N_17399,N_15336);
and U23627 (N_23627,N_16250,N_18161);
nand U23628 (N_23628,N_17908,N_18868);
and U23629 (N_23629,N_18631,N_17942);
and U23630 (N_23630,N_15157,N_15859);
or U23631 (N_23631,N_18211,N_16282);
nor U23632 (N_23632,N_17787,N_18325);
or U23633 (N_23633,N_17515,N_17193);
and U23634 (N_23634,N_19985,N_16531);
xnor U23635 (N_23635,N_15201,N_15104);
nor U23636 (N_23636,N_16925,N_15522);
nand U23637 (N_23637,N_15324,N_15695);
or U23638 (N_23638,N_17258,N_16549);
and U23639 (N_23639,N_16625,N_18623);
and U23640 (N_23640,N_17558,N_19402);
or U23641 (N_23641,N_18539,N_18670);
or U23642 (N_23642,N_16591,N_18913);
and U23643 (N_23643,N_19264,N_18466);
or U23644 (N_23644,N_17629,N_17281);
nor U23645 (N_23645,N_15464,N_16414);
nor U23646 (N_23646,N_19884,N_17176);
and U23647 (N_23647,N_16955,N_16800);
xnor U23648 (N_23648,N_17713,N_19886);
xor U23649 (N_23649,N_15245,N_16018);
nor U23650 (N_23650,N_17821,N_19128);
and U23651 (N_23651,N_19034,N_16270);
nor U23652 (N_23652,N_15396,N_19480);
nand U23653 (N_23653,N_16003,N_15553);
or U23654 (N_23654,N_15574,N_16952);
or U23655 (N_23655,N_19027,N_19015);
nor U23656 (N_23656,N_19536,N_19417);
nand U23657 (N_23657,N_18701,N_15918);
xnor U23658 (N_23658,N_16348,N_18600);
or U23659 (N_23659,N_17144,N_15704);
xnor U23660 (N_23660,N_17570,N_15560);
or U23661 (N_23661,N_18881,N_16230);
and U23662 (N_23662,N_15369,N_17628);
nor U23663 (N_23663,N_19190,N_16581);
nand U23664 (N_23664,N_18672,N_16360);
nor U23665 (N_23665,N_18971,N_19909);
xor U23666 (N_23666,N_16714,N_15892);
nand U23667 (N_23667,N_19375,N_19446);
nor U23668 (N_23668,N_16218,N_18933);
or U23669 (N_23669,N_16812,N_15352);
nand U23670 (N_23670,N_16542,N_15360);
nand U23671 (N_23671,N_15309,N_15253);
nor U23672 (N_23672,N_15076,N_15660);
or U23673 (N_23673,N_15509,N_17219);
xor U23674 (N_23674,N_18794,N_17959);
nor U23675 (N_23675,N_16226,N_19082);
nor U23676 (N_23676,N_19498,N_19857);
and U23677 (N_23677,N_18110,N_18777);
or U23678 (N_23678,N_15683,N_18407);
and U23679 (N_23679,N_16791,N_17307);
nor U23680 (N_23680,N_19969,N_19654);
xnor U23681 (N_23681,N_18926,N_15252);
nor U23682 (N_23682,N_19045,N_18372);
or U23683 (N_23683,N_18462,N_16176);
xor U23684 (N_23684,N_15739,N_16933);
xor U23685 (N_23685,N_17642,N_18234);
or U23686 (N_23686,N_18488,N_19827);
nand U23687 (N_23687,N_15641,N_18545);
xor U23688 (N_23688,N_15084,N_15797);
xor U23689 (N_23689,N_16239,N_19630);
or U23690 (N_23690,N_16554,N_16013);
or U23691 (N_23691,N_18719,N_18615);
nand U23692 (N_23692,N_18555,N_16917);
and U23693 (N_23693,N_18688,N_18059);
and U23694 (N_23694,N_17296,N_19209);
and U23695 (N_23695,N_17231,N_18251);
nand U23696 (N_23696,N_17730,N_15640);
xor U23697 (N_23697,N_17623,N_15818);
or U23698 (N_23698,N_16144,N_17507);
and U23699 (N_23699,N_18185,N_19171);
and U23700 (N_23700,N_18685,N_15996);
or U23701 (N_23701,N_15488,N_16590);
or U23702 (N_23702,N_19852,N_18746);
and U23703 (N_23703,N_18550,N_17048);
or U23704 (N_23704,N_18912,N_18083);
xnor U23705 (N_23705,N_19786,N_19424);
or U23706 (N_23706,N_19107,N_16544);
nor U23707 (N_23707,N_15483,N_15754);
xor U23708 (N_23708,N_19041,N_18989);
or U23709 (N_23709,N_19250,N_19570);
xnor U23710 (N_23710,N_16022,N_15082);
and U23711 (N_23711,N_15529,N_18606);
nor U23712 (N_23712,N_18127,N_15561);
and U23713 (N_23713,N_19788,N_19768);
nor U23714 (N_23714,N_18609,N_18484);
and U23715 (N_23715,N_18182,N_17020);
xnor U23716 (N_23716,N_19487,N_15728);
nor U23717 (N_23717,N_18231,N_17465);
nor U23718 (N_23718,N_15140,N_16780);
or U23719 (N_23719,N_16861,N_18678);
nand U23720 (N_23720,N_18427,N_18407);
nand U23721 (N_23721,N_19707,N_17570);
xnor U23722 (N_23722,N_17490,N_19338);
nor U23723 (N_23723,N_18386,N_15189);
or U23724 (N_23724,N_17186,N_18854);
xnor U23725 (N_23725,N_15110,N_17948);
nor U23726 (N_23726,N_17848,N_18223);
nand U23727 (N_23727,N_17937,N_18402);
nor U23728 (N_23728,N_17478,N_18890);
nand U23729 (N_23729,N_15321,N_19909);
nand U23730 (N_23730,N_15992,N_15165);
nand U23731 (N_23731,N_16222,N_18972);
nand U23732 (N_23732,N_16304,N_19650);
or U23733 (N_23733,N_15241,N_16923);
nand U23734 (N_23734,N_16232,N_19916);
and U23735 (N_23735,N_16420,N_18794);
xor U23736 (N_23736,N_15610,N_18844);
xor U23737 (N_23737,N_15035,N_17891);
or U23738 (N_23738,N_15025,N_19598);
nand U23739 (N_23739,N_18359,N_19404);
nor U23740 (N_23740,N_15271,N_19354);
xnor U23741 (N_23741,N_19954,N_16986);
xnor U23742 (N_23742,N_16665,N_19182);
or U23743 (N_23743,N_16479,N_18284);
nand U23744 (N_23744,N_15654,N_16893);
nor U23745 (N_23745,N_18478,N_15756);
nand U23746 (N_23746,N_15771,N_19466);
or U23747 (N_23747,N_15688,N_15545);
nand U23748 (N_23748,N_18881,N_16476);
xor U23749 (N_23749,N_16804,N_18606);
nor U23750 (N_23750,N_18134,N_18663);
nand U23751 (N_23751,N_15938,N_19253);
nand U23752 (N_23752,N_17402,N_18998);
nor U23753 (N_23753,N_18214,N_19700);
xnor U23754 (N_23754,N_16558,N_16016);
nand U23755 (N_23755,N_15179,N_15826);
nand U23756 (N_23756,N_15174,N_19294);
nor U23757 (N_23757,N_15716,N_16430);
and U23758 (N_23758,N_19058,N_19957);
or U23759 (N_23759,N_15368,N_17214);
nor U23760 (N_23760,N_17494,N_16632);
nand U23761 (N_23761,N_15656,N_19018);
nor U23762 (N_23762,N_17338,N_18075);
nor U23763 (N_23763,N_15429,N_17242);
or U23764 (N_23764,N_16906,N_16395);
or U23765 (N_23765,N_18608,N_17393);
xnor U23766 (N_23766,N_15461,N_19506);
nand U23767 (N_23767,N_17610,N_15367);
nand U23768 (N_23768,N_18623,N_17356);
and U23769 (N_23769,N_16749,N_16809);
nor U23770 (N_23770,N_19310,N_16667);
or U23771 (N_23771,N_19946,N_19937);
nand U23772 (N_23772,N_16930,N_17758);
nor U23773 (N_23773,N_16107,N_15452);
and U23774 (N_23774,N_17960,N_18455);
and U23775 (N_23775,N_16804,N_17635);
xnor U23776 (N_23776,N_17765,N_16127);
xnor U23777 (N_23777,N_16069,N_18774);
or U23778 (N_23778,N_19767,N_16468);
and U23779 (N_23779,N_18233,N_17287);
xor U23780 (N_23780,N_16378,N_16766);
and U23781 (N_23781,N_16881,N_19302);
or U23782 (N_23782,N_18908,N_17285);
nand U23783 (N_23783,N_18312,N_17531);
nor U23784 (N_23784,N_18577,N_17400);
and U23785 (N_23785,N_18527,N_18291);
nand U23786 (N_23786,N_19687,N_19479);
and U23787 (N_23787,N_17310,N_18482);
nor U23788 (N_23788,N_15109,N_18650);
nand U23789 (N_23789,N_18729,N_15236);
or U23790 (N_23790,N_15724,N_15665);
nor U23791 (N_23791,N_17015,N_18251);
or U23792 (N_23792,N_18375,N_18136);
nor U23793 (N_23793,N_16105,N_18354);
nor U23794 (N_23794,N_16415,N_19593);
xor U23795 (N_23795,N_16972,N_17861);
or U23796 (N_23796,N_18224,N_16531);
nand U23797 (N_23797,N_15962,N_15873);
nand U23798 (N_23798,N_15153,N_16890);
xor U23799 (N_23799,N_17479,N_18671);
and U23800 (N_23800,N_18015,N_18746);
and U23801 (N_23801,N_16187,N_18975);
or U23802 (N_23802,N_17094,N_18230);
and U23803 (N_23803,N_15230,N_19647);
and U23804 (N_23804,N_15252,N_16897);
xnor U23805 (N_23805,N_16530,N_19091);
nand U23806 (N_23806,N_15253,N_19820);
xnor U23807 (N_23807,N_17124,N_17118);
nor U23808 (N_23808,N_19147,N_18446);
xnor U23809 (N_23809,N_17643,N_19531);
nand U23810 (N_23810,N_19224,N_19363);
and U23811 (N_23811,N_15929,N_18630);
nor U23812 (N_23812,N_19421,N_17501);
and U23813 (N_23813,N_17741,N_17559);
or U23814 (N_23814,N_15538,N_17203);
nand U23815 (N_23815,N_17645,N_17140);
nand U23816 (N_23816,N_15846,N_15810);
nor U23817 (N_23817,N_15989,N_19068);
nand U23818 (N_23818,N_19599,N_18746);
xor U23819 (N_23819,N_19907,N_17439);
and U23820 (N_23820,N_18584,N_15090);
xnor U23821 (N_23821,N_17355,N_19785);
xor U23822 (N_23822,N_16746,N_19624);
xnor U23823 (N_23823,N_15360,N_18617);
nor U23824 (N_23824,N_19844,N_19383);
nand U23825 (N_23825,N_15916,N_17219);
or U23826 (N_23826,N_16091,N_17409);
nand U23827 (N_23827,N_16556,N_18680);
xnor U23828 (N_23828,N_19555,N_18576);
nor U23829 (N_23829,N_19083,N_16526);
or U23830 (N_23830,N_18257,N_15502);
xor U23831 (N_23831,N_15193,N_18352);
nand U23832 (N_23832,N_15740,N_16304);
nor U23833 (N_23833,N_18765,N_16349);
and U23834 (N_23834,N_19250,N_19770);
or U23835 (N_23835,N_16450,N_17691);
or U23836 (N_23836,N_19772,N_15463);
nor U23837 (N_23837,N_18191,N_19989);
nand U23838 (N_23838,N_16485,N_18093);
xor U23839 (N_23839,N_18760,N_17432);
nor U23840 (N_23840,N_16989,N_18677);
and U23841 (N_23841,N_17669,N_19572);
nor U23842 (N_23842,N_16736,N_16126);
and U23843 (N_23843,N_17814,N_16071);
or U23844 (N_23844,N_15837,N_17509);
nor U23845 (N_23845,N_18079,N_16785);
and U23846 (N_23846,N_17586,N_19904);
nand U23847 (N_23847,N_19032,N_19429);
nand U23848 (N_23848,N_19337,N_17054);
xor U23849 (N_23849,N_15025,N_16591);
nor U23850 (N_23850,N_18172,N_16603);
nand U23851 (N_23851,N_15018,N_18213);
nand U23852 (N_23852,N_15068,N_18052);
xnor U23853 (N_23853,N_17368,N_18505);
and U23854 (N_23854,N_18290,N_15862);
and U23855 (N_23855,N_16779,N_17988);
nor U23856 (N_23856,N_16432,N_19767);
nand U23857 (N_23857,N_18338,N_17020);
nor U23858 (N_23858,N_17904,N_15436);
and U23859 (N_23859,N_15355,N_17514);
and U23860 (N_23860,N_16139,N_17613);
nand U23861 (N_23861,N_17601,N_18181);
xnor U23862 (N_23862,N_16791,N_16239);
and U23863 (N_23863,N_17720,N_16976);
or U23864 (N_23864,N_15874,N_15542);
and U23865 (N_23865,N_16980,N_16477);
and U23866 (N_23866,N_17802,N_17610);
nor U23867 (N_23867,N_15183,N_17311);
or U23868 (N_23868,N_15809,N_17104);
or U23869 (N_23869,N_15510,N_16879);
nor U23870 (N_23870,N_17643,N_19462);
nor U23871 (N_23871,N_17133,N_18118);
nor U23872 (N_23872,N_19103,N_15094);
xnor U23873 (N_23873,N_16091,N_15168);
or U23874 (N_23874,N_15107,N_16213);
or U23875 (N_23875,N_15993,N_16551);
xnor U23876 (N_23876,N_15601,N_18497);
nor U23877 (N_23877,N_18556,N_16974);
and U23878 (N_23878,N_15647,N_15981);
or U23879 (N_23879,N_19247,N_17220);
nand U23880 (N_23880,N_16063,N_17526);
and U23881 (N_23881,N_18942,N_16173);
and U23882 (N_23882,N_16078,N_19030);
nor U23883 (N_23883,N_19612,N_15311);
xor U23884 (N_23884,N_17361,N_16710);
nor U23885 (N_23885,N_19459,N_18179);
nor U23886 (N_23886,N_17942,N_15272);
and U23887 (N_23887,N_19911,N_15727);
and U23888 (N_23888,N_18384,N_19377);
or U23889 (N_23889,N_15784,N_16776);
nand U23890 (N_23890,N_16504,N_15918);
and U23891 (N_23891,N_17156,N_17190);
xnor U23892 (N_23892,N_17959,N_19170);
or U23893 (N_23893,N_16281,N_16124);
nor U23894 (N_23894,N_19305,N_16619);
nor U23895 (N_23895,N_17297,N_17317);
and U23896 (N_23896,N_19712,N_15162);
xnor U23897 (N_23897,N_16666,N_16979);
xor U23898 (N_23898,N_19321,N_16112);
nor U23899 (N_23899,N_17282,N_17839);
nand U23900 (N_23900,N_17228,N_17854);
or U23901 (N_23901,N_19859,N_18333);
nor U23902 (N_23902,N_16642,N_18581);
or U23903 (N_23903,N_16003,N_19233);
nand U23904 (N_23904,N_18994,N_19059);
and U23905 (N_23905,N_17391,N_16991);
nor U23906 (N_23906,N_15667,N_19534);
or U23907 (N_23907,N_17186,N_16962);
xnor U23908 (N_23908,N_18535,N_16944);
or U23909 (N_23909,N_19104,N_16551);
xnor U23910 (N_23910,N_17973,N_17600);
nand U23911 (N_23911,N_15780,N_18532);
or U23912 (N_23912,N_17710,N_15052);
nand U23913 (N_23913,N_15267,N_17705);
xnor U23914 (N_23914,N_19852,N_15564);
xnor U23915 (N_23915,N_17268,N_18659);
or U23916 (N_23916,N_16678,N_15628);
nor U23917 (N_23917,N_19261,N_15297);
or U23918 (N_23918,N_16213,N_18290);
nor U23919 (N_23919,N_18633,N_15988);
or U23920 (N_23920,N_15960,N_18581);
nor U23921 (N_23921,N_18653,N_19797);
nand U23922 (N_23922,N_19456,N_16538);
nor U23923 (N_23923,N_15478,N_17414);
or U23924 (N_23924,N_15477,N_17882);
nand U23925 (N_23925,N_17501,N_15841);
nand U23926 (N_23926,N_17278,N_15982);
nor U23927 (N_23927,N_16320,N_18979);
nor U23928 (N_23928,N_15741,N_18753);
nor U23929 (N_23929,N_16439,N_18318);
nor U23930 (N_23930,N_17536,N_19781);
or U23931 (N_23931,N_18316,N_19697);
nor U23932 (N_23932,N_19800,N_16926);
xnor U23933 (N_23933,N_18386,N_19299);
nand U23934 (N_23934,N_18195,N_16690);
nor U23935 (N_23935,N_15555,N_17789);
nand U23936 (N_23936,N_17155,N_15777);
or U23937 (N_23937,N_18222,N_15027);
and U23938 (N_23938,N_17969,N_18300);
or U23939 (N_23939,N_18895,N_18765);
or U23940 (N_23940,N_18015,N_15859);
and U23941 (N_23941,N_16884,N_17561);
nand U23942 (N_23942,N_18622,N_15640);
nand U23943 (N_23943,N_17701,N_16486);
or U23944 (N_23944,N_17525,N_18728);
nor U23945 (N_23945,N_16582,N_17720);
xnor U23946 (N_23946,N_15274,N_16744);
or U23947 (N_23947,N_17139,N_16348);
xnor U23948 (N_23948,N_15417,N_15506);
and U23949 (N_23949,N_15982,N_19327);
nand U23950 (N_23950,N_17875,N_18037);
and U23951 (N_23951,N_17006,N_17163);
nor U23952 (N_23952,N_19959,N_15153);
xor U23953 (N_23953,N_19157,N_17530);
or U23954 (N_23954,N_18449,N_17349);
xnor U23955 (N_23955,N_17319,N_17902);
nand U23956 (N_23956,N_15933,N_17901);
and U23957 (N_23957,N_15303,N_16448);
and U23958 (N_23958,N_15010,N_16375);
and U23959 (N_23959,N_16383,N_17689);
xor U23960 (N_23960,N_18562,N_17411);
or U23961 (N_23961,N_16058,N_17133);
or U23962 (N_23962,N_19188,N_18035);
nor U23963 (N_23963,N_15959,N_19557);
nor U23964 (N_23964,N_17012,N_16714);
xor U23965 (N_23965,N_19100,N_19501);
and U23966 (N_23966,N_19759,N_18849);
or U23967 (N_23967,N_16336,N_18059);
nand U23968 (N_23968,N_19251,N_19101);
xnor U23969 (N_23969,N_16110,N_15748);
nor U23970 (N_23970,N_17939,N_18062);
xnor U23971 (N_23971,N_18983,N_16354);
or U23972 (N_23972,N_19770,N_15739);
xor U23973 (N_23973,N_19047,N_15413);
nor U23974 (N_23974,N_16575,N_17816);
and U23975 (N_23975,N_15347,N_17579);
nand U23976 (N_23976,N_16236,N_19510);
nand U23977 (N_23977,N_19105,N_19895);
nor U23978 (N_23978,N_16121,N_18876);
nand U23979 (N_23979,N_15051,N_17371);
nor U23980 (N_23980,N_17547,N_16171);
and U23981 (N_23981,N_15025,N_18232);
xnor U23982 (N_23982,N_17248,N_18898);
or U23983 (N_23983,N_16909,N_19593);
nand U23984 (N_23984,N_18843,N_18735);
xnor U23985 (N_23985,N_15313,N_18005);
and U23986 (N_23986,N_15953,N_15441);
or U23987 (N_23987,N_18695,N_16953);
xor U23988 (N_23988,N_16778,N_19319);
or U23989 (N_23989,N_17886,N_19325);
nand U23990 (N_23990,N_17755,N_15296);
nand U23991 (N_23991,N_19899,N_18204);
and U23992 (N_23992,N_15817,N_16318);
xnor U23993 (N_23993,N_15323,N_19356);
nand U23994 (N_23994,N_15164,N_17265);
or U23995 (N_23995,N_19585,N_19175);
and U23996 (N_23996,N_18033,N_18824);
nand U23997 (N_23997,N_16652,N_15192);
xnor U23998 (N_23998,N_17888,N_15327);
and U23999 (N_23999,N_18079,N_18065);
xor U24000 (N_24000,N_19631,N_19139);
xnor U24001 (N_24001,N_16122,N_15529);
nor U24002 (N_24002,N_15798,N_15375);
and U24003 (N_24003,N_17168,N_16159);
and U24004 (N_24004,N_16532,N_16641);
nand U24005 (N_24005,N_17668,N_16964);
nor U24006 (N_24006,N_19984,N_15475);
and U24007 (N_24007,N_15777,N_19430);
xnor U24008 (N_24008,N_19920,N_15971);
nor U24009 (N_24009,N_17567,N_18754);
nand U24010 (N_24010,N_19104,N_15762);
nor U24011 (N_24011,N_19728,N_16728);
and U24012 (N_24012,N_15770,N_19039);
xnor U24013 (N_24013,N_16506,N_17376);
nor U24014 (N_24014,N_19173,N_18835);
or U24015 (N_24015,N_15563,N_19987);
and U24016 (N_24016,N_15776,N_19249);
nand U24017 (N_24017,N_17393,N_16602);
xnor U24018 (N_24018,N_15182,N_15031);
xnor U24019 (N_24019,N_18779,N_17134);
nor U24020 (N_24020,N_17821,N_16555);
xor U24021 (N_24021,N_18496,N_18730);
or U24022 (N_24022,N_18636,N_17079);
nand U24023 (N_24023,N_19913,N_17368);
and U24024 (N_24024,N_15834,N_16447);
xnor U24025 (N_24025,N_18620,N_16149);
nor U24026 (N_24026,N_15872,N_19707);
or U24027 (N_24027,N_19984,N_18300);
or U24028 (N_24028,N_18331,N_19511);
nor U24029 (N_24029,N_15819,N_15523);
and U24030 (N_24030,N_17111,N_17369);
xor U24031 (N_24031,N_15355,N_16654);
nor U24032 (N_24032,N_15195,N_19240);
nor U24033 (N_24033,N_19980,N_16175);
xor U24034 (N_24034,N_17144,N_18939);
xnor U24035 (N_24035,N_19775,N_19549);
and U24036 (N_24036,N_17457,N_17933);
or U24037 (N_24037,N_17974,N_15387);
nand U24038 (N_24038,N_17825,N_17470);
nand U24039 (N_24039,N_16279,N_19656);
xor U24040 (N_24040,N_17898,N_17792);
and U24041 (N_24041,N_16792,N_16864);
xnor U24042 (N_24042,N_17257,N_18587);
nor U24043 (N_24043,N_17921,N_16871);
nor U24044 (N_24044,N_16581,N_15461);
or U24045 (N_24045,N_16317,N_18640);
and U24046 (N_24046,N_17345,N_15175);
xnor U24047 (N_24047,N_16486,N_16056);
nand U24048 (N_24048,N_17399,N_19995);
nor U24049 (N_24049,N_18635,N_18890);
nor U24050 (N_24050,N_18261,N_19567);
and U24051 (N_24051,N_18822,N_19620);
nand U24052 (N_24052,N_16694,N_15696);
nor U24053 (N_24053,N_17116,N_16600);
or U24054 (N_24054,N_19617,N_15874);
and U24055 (N_24055,N_15052,N_17085);
nand U24056 (N_24056,N_15552,N_18865);
and U24057 (N_24057,N_15346,N_15444);
or U24058 (N_24058,N_16178,N_16172);
or U24059 (N_24059,N_16349,N_19384);
or U24060 (N_24060,N_18041,N_18759);
and U24061 (N_24061,N_17201,N_19577);
or U24062 (N_24062,N_17037,N_18667);
nor U24063 (N_24063,N_18976,N_19881);
nor U24064 (N_24064,N_18407,N_15998);
or U24065 (N_24065,N_18474,N_19138);
nand U24066 (N_24066,N_18096,N_15795);
xor U24067 (N_24067,N_18164,N_15097);
nand U24068 (N_24068,N_17567,N_18599);
nand U24069 (N_24069,N_17826,N_17602);
nor U24070 (N_24070,N_17593,N_16667);
and U24071 (N_24071,N_18939,N_15530);
and U24072 (N_24072,N_17970,N_18928);
nand U24073 (N_24073,N_19019,N_18716);
nor U24074 (N_24074,N_18653,N_17083);
xnor U24075 (N_24075,N_17793,N_15723);
xnor U24076 (N_24076,N_18271,N_19667);
and U24077 (N_24077,N_16962,N_16488);
nor U24078 (N_24078,N_17083,N_19202);
or U24079 (N_24079,N_19647,N_18305);
xor U24080 (N_24080,N_17924,N_17159);
nor U24081 (N_24081,N_18520,N_17169);
nand U24082 (N_24082,N_15551,N_18089);
nand U24083 (N_24083,N_18020,N_18345);
xnor U24084 (N_24084,N_15970,N_19704);
or U24085 (N_24085,N_17233,N_19307);
nor U24086 (N_24086,N_15226,N_18671);
xnor U24087 (N_24087,N_15351,N_17649);
xor U24088 (N_24088,N_18990,N_15488);
nand U24089 (N_24089,N_17846,N_15283);
nor U24090 (N_24090,N_16680,N_15899);
xnor U24091 (N_24091,N_17670,N_15698);
and U24092 (N_24092,N_17313,N_15174);
xnor U24093 (N_24093,N_17762,N_16766);
nor U24094 (N_24094,N_17865,N_18137);
xnor U24095 (N_24095,N_15750,N_15373);
nor U24096 (N_24096,N_18845,N_18733);
xor U24097 (N_24097,N_18589,N_19118);
and U24098 (N_24098,N_15345,N_16928);
xnor U24099 (N_24099,N_16617,N_18197);
nand U24100 (N_24100,N_19032,N_17816);
and U24101 (N_24101,N_18220,N_17154);
and U24102 (N_24102,N_17852,N_18822);
nand U24103 (N_24103,N_15155,N_15166);
nor U24104 (N_24104,N_19870,N_15038);
or U24105 (N_24105,N_16992,N_18545);
or U24106 (N_24106,N_17693,N_17169);
or U24107 (N_24107,N_18197,N_18858);
xor U24108 (N_24108,N_15269,N_15025);
and U24109 (N_24109,N_17655,N_15967);
and U24110 (N_24110,N_19925,N_17813);
xnor U24111 (N_24111,N_17061,N_16614);
xor U24112 (N_24112,N_15434,N_18701);
nand U24113 (N_24113,N_19705,N_17319);
nand U24114 (N_24114,N_15119,N_16805);
or U24115 (N_24115,N_16694,N_16569);
or U24116 (N_24116,N_16542,N_15804);
nor U24117 (N_24117,N_15819,N_17571);
or U24118 (N_24118,N_15358,N_16861);
xnor U24119 (N_24119,N_15192,N_17135);
xnor U24120 (N_24120,N_18963,N_16347);
or U24121 (N_24121,N_18356,N_16785);
or U24122 (N_24122,N_15428,N_16572);
xnor U24123 (N_24123,N_17510,N_19391);
or U24124 (N_24124,N_18486,N_19597);
and U24125 (N_24125,N_16161,N_19311);
nor U24126 (N_24126,N_16006,N_18896);
and U24127 (N_24127,N_18415,N_15722);
or U24128 (N_24128,N_16304,N_19620);
xor U24129 (N_24129,N_16118,N_18895);
nor U24130 (N_24130,N_15356,N_15607);
or U24131 (N_24131,N_17280,N_15855);
and U24132 (N_24132,N_15266,N_17087);
nand U24133 (N_24133,N_17726,N_19486);
nor U24134 (N_24134,N_17505,N_17628);
xor U24135 (N_24135,N_17448,N_15682);
xnor U24136 (N_24136,N_17164,N_19829);
and U24137 (N_24137,N_19170,N_17408);
nor U24138 (N_24138,N_19893,N_19113);
nor U24139 (N_24139,N_19649,N_19291);
xnor U24140 (N_24140,N_18093,N_16553);
nand U24141 (N_24141,N_17854,N_17213);
xnor U24142 (N_24142,N_16765,N_16369);
nor U24143 (N_24143,N_17251,N_15459);
or U24144 (N_24144,N_19916,N_19971);
nor U24145 (N_24145,N_18874,N_18067);
nand U24146 (N_24146,N_18241,N_15450);
nor U24147 (N_24147,N_15393,N_15352);
or U24148 (N_24148,N_16510,N_17580);
or U24149 (N_24149,N_16493,N_18871);
nand U24150 (N_24150,N_18877,N_15322);
xnor U24151 (N_24151,N_18703,N_16070);
nor U24152 (N_24152,N_17304,N_19490);
nor U24153 (N_24153,N_15008,N_18373);
or U24154 (N_24154,N_19592,N_16642);
nor U24155 (N_24155,N_19491,N_16892);
and U24156 (N_24156,N_16093,N_18175);
nor U24157 (N_24157,N_19452,N_17046);
xor U24158 (N_24158,N_19450,N_19338);
and U24159 (N_24159,N_18612,N_16432);
and U24160 (N_24160,N_17652,N_17444);
xnor U24161 (N_24161,N_17884,N_19884);
or U24162 (N_24162,N_15633,N_19130);
or U24163 (N_24163,N_16076,N_19518);
and U24164 (N_24164,N_18152,N_18557);
nand U24165 (N_24165,N_19200,N_18840);
nor U24166 (N_24166,N_17761,N_19216);
and U24167 (N_24167,N_18808,N_19546);
nor U24168 (N_24168,N_19736,N_19223);
nand U24169 (N_24169,N_16469,N_19379);
xor U24170 (N_24170,N_19172,N_17313);
nand U24171 (N_24171,N_15937,N_16718);
and U24172 (N_24172,N_15406,N_18401);
xor U24173 (N_24173,N_17253,N_15837);
or U24174 (N_24174,N_16567,N_15631);
nand U24175 (N_24175,N_16682,N_18468);
or U24176 (N_24176,N_15222,N_17771);
xor U24177 (N_24177,N_18653,N_15900);
nor U24178 (N_24178,N_15139,N_18412);
nand U24179 (N_24179,N_17027,N_17528);
or U24180 (N_24180,N_17525,N_17438);
or U24181 (N_24181,N_17527,N_19870);
xor U24182 (N_24182,N_18895,N_16745);
or U24183 (N_24183,N_16312,N_17399);
xnor U24184 (N_24184,N_16165,N_19139);
and U24185 (N_24185,N_19549,N_19499);
or U24186 (N_24186,N_15145,N_19060);
nor U24187 (N_24187,N_17141,N_15669);
nand U24188 (N_24188,N_18653,N_17983);
xor U24189 (N_24189,N_17446,N_16328);
and U24190 (N_24190,N_19656,N_19641);
or U24191 (N_24191,N_16920,N_19773);
nand U24192 (N_24192,N_18979,N_15756);
xor U24193 (N_24193,N_18000,N_16773);
nor U24194 (N_24194,N_18305,N_17547);
or U24195 (N_24195,N_16766,N_17694);
nor U24196 (N_24196,N_19300,N_19732);
xor U24197 (N_24197,N_18262,N_18249);
and U24198 (N_24198,N_19796,N_17254);
and U24199 (N_24199,N_17799,N_18273);
nand U24200 (N_24200,N_19871,N_18665);
and U24201 (N_24201,N_19057,N_18608);
nand U24202 (N_24202,N_17928,N_19041);
xnor U24203 (N_24203,N_15981,N_17999);
xnor U24204 (N_24204,N_19915,N_17460);
or U24205 (N_24205,N_16482,N_18386);
and U24206 (N_24206,N_15347,N_15177);
xnor U24207 (N_24207,N_15494,N_16857);
xor U24208 (N_24208,N_16010,N_17024);
or U24209 (N_24209,N_18757,N_19702);
xnor U24210 (N_24210,N_15609,N_15370);
nor U24211 (N_24211,N_16099,N_17060);
nand U24212 (N_24212,N_19423,N_15884);
nor U24213 (N_24213,N_15921,N_16164);
nand U24214 (N_24214,N_17509,N_19531);
nor U24215 (N_24215,N_15900,N_17470);
and U24216 (N_24216,N_16057,N_15270);
xnor U24217 (N_24217,N_16091,N_16138);
and U24218 (N_24218,N_18877,N_15469);
or U24219 (N_24219,N_15828,N_18397);
and U24220 (N_24220,N_19107,N_19417);
xor U24221 (N_24221,N_15202,N_17514);
nor U24222 (N_24222,N_17908,N_16975);
nor U24223 (N_24223,N_15980,N_18637);
nor U24224 (N_24224,N_19124,N_19663);
or U24225 (N_24225,N_16188,N_18016);
nand U24226 (N_24226,N_19756,N_15046);
and U24227 (N_24227,N_17318,N_17446);
nor U24228 (N_24228,N_17887,N_15938);
nand U24229 (N_24229,N_16729,N_18064);
nand U24230 (N_24230,N_15330,N_16566);
nand U24231 (N_24231,N_15062,N_19030);
or U24232 (N_24232,N_15400,N_17267);
or U24233 (N_24233,N_15832,N_19119);
and U24234 (N_24234,N_19426,N_16045);
and U24235 (N_24235,N_17489,N_15934);
and U24236 (N_24236,N_19986,N_18334);
and U24237 (N_24237,N_16207,N_15319);
or U24238 (N_24238,N_17927,N_18823);
nand U24239 (N_24239,N_16721,N_17491);
xor U24240 (N_24240,N_17573,N_16350);
nor U24241 (N_24241,N_17338,N_16582);
xor U24242 (N_24242,N_19565,N_18494);
xor U24243 (N_24243,N_15036,N_19016);
nor U24244 (N_24244,N_19903,N_16742);
nor U24245 (N_24245,N_17313,N_18692);
or U24246 (N_24246,N_16005,N_17499);
or U24247 (N_24247,N_15055,N_16322);
nand U24248 (N_24248,N_19631,N_16679);
nand U24249 (N_24249,N_16419,N_19735);
xor U24250 (N_24250,N_15775,N_18779);
nor U24251 (N_24251,N_18766,N_18729);
nor U24252 (N_24252,N_15286,N_17237);
or U24253 (N_24253,N_17591,N_15177);
or U24254 (N_24254,N_19295,N_16880);
nor U24255 (N_24255,N_17182,N_15889);
xnor U24256 (N_24256,N_19430,N_19751);
or U24257 (N_24257,N_16786,N_17549);
xnor U24258 (N_24258,N_17036,N_18932);
and U24259 (N_24259,N_18485,N_19858);
nand U24260 (N_24260,N_15288,N_19553);
or U24261 (N_24261,N_16319,N_17687);
xor U24262 (N_24262,N_15358,N_17220);
nand U24263 (N_24263,N_19342,N_15079);
xor U24264 (N_24264,N_15584,N_15366);
and U24265 (N_24265,N_15606,N_15255);
and U24266 (N_24266,N_18492,N_16172);
nand U24267 (N_24267,N_17593,N_15497);
xnor U24268 (N_24268,N_16683,N_19253);
nand U24269 (N_24269,N_16232,N_16174);
or U24270 (N_24270,N_17816,N_15593);
and U24271 (N_24271,N_19814,N_17186);
nor U24272 (N_24272,N_16665,N_17375);
or U24273 (N_24273,N_16329,N_17085);
nand U24274 (N_24274,N_15294,N_15841);
and U24275 (N_24275,N_19462,N_17007);
nand U24276 (N_24276,N_19542,N_16651);
and U24277 (N_24277,N_19497,N_19193);
and U24278 (N_24278,N_19604,N_19054);
nand U24279 (N_24279,N_15263,N_15382);
xnor U24280 (N_24280,N_16972,N_19050);
and U24281 (N_24281,N_19419,N_17433);
nand U24282 (N_24282,N_17079,N_17281);
nor U24283 (N_24283,N_16962,N_18010);
or U24284 (N_24284,N_18519,N_17862);
nor U24285 (N_24285,N_15284,N_16718);
nand U24286 (N_24286,N_15237,N_19416);
xnor U24287 (N_24287,N_18702,N_16593);
nor U24288 (N_24288,N_18555,N_17738);
nand U24289 (N_24289,N_18271,N_18808);
nor U24290 (N_24290,N_15927,N_19625);
nor U24291 (N_24291,N_19201,N_16723);
xor U24292 (N_24292,N_16137,N_19154);
and U24293 (N_24293,N_16486,N_17094);
nor U24294 (N_24294,N_18519,N_16424);
and U24295 (N_24295,N_15079,N_16801);
and U24296 (N_24296,N_16206,N_19536);
xor U24297 (N_24297,N_18341,N_18794);
or U24298 (N_24298,N_18554,N_16183);
and U24299 (N_24299,N_19772,N_19484);
xor U24300 (N_24300,N_17656,N_17919);
and U24301 (N_24301,N_18930,N_15575);
nor U24302 (N_24302,N_16596,N_19160);
and U24303 (N_24303,N_18195,N_18116);
nor U24304 (N_24304,N_16123,N_17036);
xnor U24305 (N_24305,N_19620,N_18622);
nand U24306 (N_24306,N_16904,N_16658);
xor U24307 (N_24307,N_17865,N_15618);
xnor U24308 (N_24308,N_16287,N_18122);
nand U24309 (N_24309,N_15035,N_18876);
nor U24310 (N_24310,N_16070,N_17694);
nand U24311 (N_24311,N_17259,N_18420);
nor U24312 (N_24312,N_16668,N_18442);
and U24313 (N_24313,N_15215,N_17617);
xnor U24314 (N_24314,N_16216,N_17538);
nand U24315 (N_24315,N_17421,N_16915);
and U24316 (N_24316,N_19564,N_16062);
nand U24317 (N_24317,N_15412,N_15361);
nor U24318 (N_24318,N_16971,N_16580);
and U24319 (N_24319,N_15490,N_18600);
or U24320 (N_24320,N_15493,N_16090);
nor U24321 (N_24321,N_16498,N_17920);
or U24322 (N_24322,N_19401,N_16842);
or U24323 (N_24323,N_15695,N_17705);
nand U24324 (N_24324,N_19014,N_19401);
nand U24325 (N_24325,N_16099,N_18885);
and U24326 (N_24326,N_17695,N_17332);
and U24327 (N_24327,N_17087,N_17781);
or U24328 (N_24328,N_18037,N_16446);
nor U24329 (N_24329,N_18100,N_15914);
xor U24330 (N_24330,N_19721,N_16415);
and U24331 (N_24331,N_16074,N_16762);
nor U24332 (N_24332,N_15036,N_17868);
nor U24333 (N_24333,N_15011,N_19000);
xnor U24334 (N_24334,N_17879,N_19730);
xnor U24335 (N_24335,N_18259,N_15594);
nor U24336 (N_24336,N_16905,N_17559);
or U24337 (N_24337,N_15877,N_15021);
or U24338 (N_24338,N_16695,N_19328);
xor U24339 (N_24339,N_17535,N_18079);
nand U24340 (N_24340,N_15982,N_17491);
or U24341 (N_24341,N_17874,N_15953);
xnor U24342 (N_24342,N_16882,N_17351);
or U24343 (N_24343,N_18433,N_15761);
or U24344 (N_24344,N_19074,N_19279);
and U24345 (N_24345,N_19639,N_19295);
xnor U24346 (N_24346,N_18306,N_18554);
nor U24347 (N_24347,N_15446,N_16896);
nor U24348 (N_24348,N_19211,N_18782);
xnor U24349 (N_24349,N_18484,N_17620);
and U24350 (N_24350,N_16723,N_19109);
and U24351 (N_24351,N_15287,N_19498);
and U24352 (N_24352,N_17563,N_18812);
xor U24353 (N_24353,N_18810,N_15172);
or U24354 (N_24354,N_15253,N_15193);
or U24355 (N_24355,N_18548,N_19342);
or U24356 (N_24356,N_16737,N_19405);
or U24357 (N_24357,N_18715,N_19925);
or U24358 (N_24358,N_17396,N_15485);
nand U24359 (N_24359,N_19943,N_17278);
nor U24360 (N_24360,N_17429,N_16082);
or U24361 (N_24361,N_19958,N_15391);
and U24362 (N_24362,N_15567,N_15526);
or U24363 (N_24363,N_17467,N_16610);
nor U24364 (N_24364,N_16521,N_17581);
and U24365 (N_24365,N_16499,N_15655);
xnor U24366 (N_24366,N_16371,N_17108);
xor U24367 (N_24367,N_16928,N_15520);
nand U24368 (N_24368,N_15373,N_19200);
xor U24369 (N_24369,N_17860,N_17992);
or U24370 (N_24370,N_16463,N_15284);
or U24371 (N_24371,N_18216,N_15276);
or U24372 (N_24372,N_17709,N_16396);
nand U24373 (N_24373,N_17326,N_15502);
nand U24374 (N_24374,N_17369,N_19199);
nor U24375 (N_24375,N_18061,N_15197);
nand U24376 (N_24376,N_17620,N_17353);
or U24377 (N_24377,N_15500,N_16600);
xnor U24378 (N_24378,N_18975,N_16232);
nand U24379 (N_24379,N_18360,N_18614);
xnor U24380 (N_24380,N_16694,N_17059);
xor U24381 (N_24381,N_17040,N_18568);
xor U24382 (N_24382,N_19841,N_15573);
and U24383 (N_24383,N_16935,N_17191);
and U24384 (N_24384,N_18906,N_19583);
xnor U24385 (N_24385,N_17616,N_19381);
xor U24386 (N_24386,N_16442,N_18357);
or U24387 (N_24387,N_17961,N_17967);
or U24388 (N_24388,N_18389,N_18051);
and U24389 (N_24389,N_17775,N_18065);
or U24390 (N_24390,N_18294,N_17421);
and U24391 (N_24391,N_19458,N_15969);
or U24392 (N_24392,N_17835,N_16013);
or U24393 (N_24393,N_16563,N_17266);
nor U24394 (N_24394,N_17866,N_16820);
nand U24395 (N_24395,N_18291,N_15714);
or U24396 (N_24396,N_15181,N_18137);
xor U24397 (N_24397,N_18415,N_19234);
xor U24398 (N_24398,N_18055,N_15874);
xor U24399 (N_24399,N_16672,N_16844);
nor U24400 (N_24400,N_17872,N_19829);
and U24401 (N_24401,N_16967,N_15178);
nor U24402 (N_24402,N_18242,N_19802);
and U24403 (N_24403,N_18003,N_17954);
and U24404 (N_24404,N_19129,N_19430);
nand U24405 (N_24405,N_15243,N_18662);
or U24406 (N_24406,N_15080,N_15157);
nand U24407 (N_24407,N_17851,N_19443);
and U24408 (N_24408,N_17857,N_19055);
and U24409 (N_24409,N_16188,N_15271);
nor U24410 (N_24410,N_19700,N_16045);
or U24411 (N_24411,N_19035,N_17387);
and U24412 (N_24412,N_15290,N_16338);
nor U24413 (N_24413,N_17157,N_17971);
and U24414 (N_24414,N_19324,N_15849);
nand U24415 (N_24415,N_18700,N_15660);
xnor U24416 (N_24416,N_19427,N_18964);
and U24417 (N_24417,N_17715,N_16805);
xor U24418 (N_24418,N_16767,N_17762);
nand U24419 (N_24419,N_17856,N_18727);
or U24420 (N_24420,N_16504,N_18682);
or U24421 (N_24421,N_17556,N_15954);
and U24422 (N_24422,N_17396,N_19661);
xor U24423 (N_24423,N_19056,N_17813);
or U24424 (N_24424,N_19924,N_16057);
nand U24425 (N_24425,N_15043,N_15652);
or U24426 (N_24426,N_15123,N_15810);
and U24427 (N_24427,N_19724,N_15392);
or U24428 (N_24428,N_15560,N_19477);
nand U24429 (N_24429,N_16857,N_18528);
xnor U24430 (N_24430,N_17423,N_19434);
nor U24431 (N_24431,N_17058,N_18172);
or U24432 (N_24432,N_16725,N_19865);
or U24433 (N_24433,N_18415,N_17417);
nor U24434 (N_24434,N_19489,N_15895);
nand U24435 (N_24435,N_18596,N_17445);
nor U24436 (N_24436,N_17178,N_17366);
nor U24437 (N_24437,N_17966,N_15164);
and U24438 (N_24438,N_19198,N_17804);
xor U24439 (N_24439,N_16033,N_18824);
or U24440 (N_24440,N_16610,N_19135);
or U24441 (N_24441,N_16894,N_15683);
nor U24442 (N_24442,N_18122,N_19620);
nor U24443 (N_24443,N_19456,N_16656);
and U24444 (N_24444,N_17023,N_18090);
nand U24445 (N_24445,N_17945,N_19186);
nand U24446 (N_24446,N_15217,N_19387);
or U24447 (N_24447,N_17945,N_19039);
nand U24448 (N_24448,N_17241,N_17024);
nand U24449 (N_24449,N_15551,N_15901);
or U24450 (N_24450,N_19805,N_16565);
xnor U24451 (N_24451,N_17390,N_15098);
nand U24452 (N_24452,N_16600,N_16935);
nand U24453 (N_24453,N_19679,N_16089);
nand U24454 (N_24454,N_17549,N_16256);
nor U24455 (N_24455,N_18737,N_16813);
nor U24456 (N_24456,N_18922,N_17099);
xor U24457 (N_24457,N_18799,N_17861);
and U24458 (N_24458,N_17642,N_18120);
or U24459 (N_24459,N_15009,N_18265);
nor U24460 (N_24460,N_17143,N_16681);
or U24461 (N_24461,N_16497,N_18555);
and U24462 (N_24462,N_15027,N_18630);
or U24463 (N_24463,N_15908,N_17428);
nand U24464 (N_24464,N_17968,N_18393);
and U24465 (N_24465,N_18738,N_19405);
and U24466 (N_24466,N_19606,N_17114);
or U24467 (N_24467,N_17382,N_15400);
or U24468 (N_24468,N_18046,N_18573);
nor U24469 (N_24469,N_17386,N_18350);
and U24470 (N_24470,N_17858,N_18508);
nand U24471 (N_24471,N_15779,N_16587);
or U24472 (N_24472,N_18046,N_19198);
or U24473 (N_24473,N_18355,N_18875);
nand U24474 (N_24474,N_19688,N_17472);
nor U24475 (N_24475,N_18568,N_15225);
nor U24476 (N_24476,N_16926,N_15534);
nand U24477 (N_24477,N_17005,N_18142);
and U24478 (N_24478,N_18305,N_17833);
and U24479 (N_24479,N_19866,N_19492);
nand U24480 (N_24480,N_17714,N_18093);
xor U24481 (N_24481,N_18819,N_15260);
and U24482 (N_24482,N_18804,N_16907);
and U24483 (N_24483,N_19582,N_18330);
or U24484 (N_24484,N_17441,N_17200);
xnor U24485 (N_24485,N_16566,N_15322);
nor U24486 (N_24486,N_16843,N_17817);
and U24487 (N_24487,N_15768,N_15764);
xnor U24488 (N_24488,N_18528,N_18588);
nand U24489 (N_24489,N_15305,N_17494);
and U24490 (N_24490,N_15731,N_19698);
and U24491 (N_24491,N_19048,N_17008);
xnor U24492 (N_24492,N_18049,N_17241);
and U24493 (N_24493,N_15275,N_19975);
xnor U24494 (N_24494,N_19604,N_15456);
and U24495 (N_24495,N_18572,N_17486);
or U24496 (N_24496,N_18078,N_19470);
or U24497 (N_24497,N_17325,N_17148);
or U24498 (N_24498,N_18131,N_17076);
or U24499 (N_24499,N_17947,N_17709);
nor U24500 (N_24500,N_16940,N_17707);
or U24501 (N_24501,N_18295,N_16820);
nor U24502 (N_24502,N_18286,N_18266);
xor U24503 (N_24503,N_19294,N_19991);
nor U24504 (N_24504,N_15304,N_18482);
nand U24505 (N_24505,N_15445,N_15105);
or U24506 (N_24506,N_16247,N_17658);
and U24507 (N_24507,N_17049,N_15344);
xnor U24508 (N_24508,N_17506,N_18799);
nor U24509 (N_24509,N_15534,N_17546);
nor U24510 (N_24510,N_18306,N_17565);
nand U24511 (N_24511,N_15606,N_19552);
or U24512 (N_24512,N_15527,N_16611);
or U24513 (N_24513,N_16048,N_17860);
nand U24514 (N_24514,N_19436,N_17685);
nor U24515 (N_24515,N_19482,N_17711);
and U24516 (N_24516,N_17044,N_19806);
or U24517 (N_24517,N_18010,N_16822);
nand U24518 (N_24518,N_17538,N_15394);
xor U24519 (N_24519,N_16913,N_19250);
nor U24520 (N_24520,N_19948,N_19445);
or U24521 (N_24521,N_15670,N_18117);
nor U24522 (N_24522,N_15329,N_18980);
and U24523 (N_24523,N_18437,N_18311);
or U24524 (N_24524,N_15113,N_17657);
xnor U24525 (N_24525,N_17167,N_19068);
and U24526 (N_24526,N_15195,N_15296);
nor U24527 (N_24527,N_18085,N_19139);
nor U24528 (N_24528,N_15705,N_15796);
nor U24529 (N_24529,N_19862,N_15212);
xor U24530 (N_24530,N_18995,N_15260);
nor U24531 (N_24531,N_19204,N_15553);
nor U24532 (N_24532,N_17874,N_18745);
nand U24533 (N_24533,N_18865,N_18502);
xor U24534 (N_24534,N_16882,N_16323);
nand U24535 (N_24535,N_18244,N_15597);
xnor U24536 (N_24536,N_17414,N_16048);
nor U24537 (N_24537,N_15241,N_16280);
nor U24538 (N_24538,N_15898,N_16711);
nor U24539 (N_24539,N_15530,N_17486);
xnor U24540 (N_24540,N_18744,N_15494);
or U24541 (N_24541,N_17423,N_15105);
or U24542 (N_24542,N_19496,N_17763);
and U24543 (N_24543,N_15841,N_16045);
xnor U24544 (N_24544,N_18815,N_18341);
xnor U24545 (N_24545,N_17052,N_17471);
and U24546 (N_24546,N_19362,N_18608);
or U24547 (N_24547,N_17190,N_15969);
and U24548 (N_24548,N_16746,N_17588);
or U24549 (N_24549,N_17982,N_19215);
nor U24550 (N_24550,N_18940,N_15327);
nor U24551 (N_24551,N_16406,N_17971);
and U24552 (N_24552,N_18161,N_15656);
or U24553 (N_24553,N_17407,N_16392);
or U24554 (N_24554,N_17028,N_15466);
nor U24555 (N_24555,N_16873,N_15621);
nand U24556 (N_24556,N_18210,N_19671);
xnor U24557 (N_24557,N_18126,N_17956);
xor U24558 (N_24558,N_16005,N_16320);
nand U24559 (N_24559,N_19966,N_17201);
xnor U24560 (N_24560,N_19896,N_16087);
xnor U24561 (N_24561,N_17029,N_15227);
xnor U24562 (N_24562,N_16304,N_16006);
xnor U24563 (N_24563,N_17187,N_19837);
and U24564 (N_24564,N_16037,N_16182);
nor U24565 (N_24565,N_16656,N_18740);
xor U24566 (N_24566,N_17084,N_15930);
nor U24567 (N_24567,N_19760,N_18038);
nand U24568 (N_24568,N_16602,N_17738);
xor U24569 (N_24569,N_18206,N_18398);
xor U24570 (N_24570,N_18095,N_16519);
or U24571 (N_24571,N_16797,N_19305);
or U24572 (N_24572,N_16827,N_16158);
xor U24573 (N_24573,N_17376,N_19434);
nand U24574 (N_24574,N_18390,N_16883);
xnor U24575 (N_24575,N_19425,N_16692);
xnor U24576 (N_24576,N_16824,N_15547);
nor U24577 (N_24577,N_18238,N_17827);
or U24578 (N_24578,N_17201,N_18418);
nand U24579 (N_24579,N_18565,N_17359);
or U24580 (N_24580,N_18326,N_18790);
xor U24581 (N_24581,N_16989,N_17898);
and U24582 (N_24582,N_17633,N_19104);
and U24583 (N_24583,N_17484,N_17238);
xnor U24584 (N_24584,N_18349,N_16850);
nor U24585 (N_24585,N_19617,N_16202);
and U24586 (N_24586,N_17347,N_17913);
and U24587 (N_24587,N_19735,N_17166);
xnor U24588 (N_24588,N_18901,N_15868);
nor U24589 (N_24589,N_17194,N_18840);
or U24590 (N_24590,N_17280,N_15386);
nand U24591 (N_24591,N_16804,N_16295);
nor U24592 (N_24592,N_19093,N_15947);
nor U24593 (N_24593,N_16396,N_15579);
or U24594 (N_24594,N_17364,N_19675);
or U24595 (N_24595,N_19285,N_18228);
and U24596 (N_24596,N_15776,N_18964);
nand U24597 (N_24597,N_17860,N_16569);
nand U24598 (N_24598,N_18606,N_18551);
nor U24599 (N_24599,N_18390,N_16319);
nand U24600 (N_24600,N_17019,N_17782);
xnor U24601 (N_24601,N_16998,N_17240);
nor U24602 (N_24602,N_16879,N_17652);
nor U24603 (N_24603,N_17553,N_16979);
nor U24604 (N_24604,N_19882,N_15633);
and U24605 (N_24605,N_17740,N_15689);
xor U24606 (N_24606,N_15834,N_19562);
and U24607 (N_24607,N_15930,N_15295);
and U24608 (N_24608,N_17031,N_16389);
nand U24609 (N_24609,N_17711,N_19102);
nor U24610 (N_24610,N_16292,N_16804);
nor U24611 (N_24611,N_19857,N_18439);
xor U24612 (N_24612,N_18348,N_17595);
xor U24613 (N_24613,N_19580,N_18005);
nand U24614 (N_24614,N_15111,N_15450);
nor U24615 (N_24615,N_19134,N_15826);
nor U24616 (N_24616,N_16382,N_16306);
nor U24617 (N_24617,N_19613,N_16298);
or U24618 (N_24618,N_18303,N_16676);
nor U24619 (N_24619,N_18554,N_16222);
nand U24620 (N_24620,N_17379,N_19862);
and U24621 (N_24621,N_15223,N_18237);
nor U24622 (N_24622,N_17861,N_17344);
xor U24623 (N_24623,N_17846,N_16125);
nor U24624 (N_24624,N_18612,N_18514);
nor U24625 (N_24625,N_18985,N_15256);
and U24626 (N_24626,N_16373,N_16335);
nor U24627 (N_24627,N_18779,N_17391);
nor U24628 (N_24628,N_15004,N_16544);
or U24629 (N_24629,N_17765,N_17098);
xor U24630 (N_24630,N_17795,N_18694);
or U24631 (N_24631,N_15274,N_18275);
xor U24632 (N_24632,N_17424,N_16356);
and U24633 (N_24633,N_19499,N_17596);
nand U24634 (N_24634,N_19374,N_15299);
xor U24635 (N_24635,N_19495,N_16618);
xnor U24636 (N_24636,N_19930,N_17962);
or U24637 (N_24637,N_19513,N_16760);
nand U24638 (N_24638,N_15701,N_15445);
and U24639 (N_24639,N_19230,N_17172);
or U24640 (N_24640,N_18372,N_15233);
nand U24641 (N_24641,N_17134,N_15840);
or U24642 (N_24642,N_17700,N_18824);
and U24643 (N_24643,N_19751,N_18998);
nand U24644 (N_24644,N_17092,N_15400);
nor U24645 (N_24645,N_15802,N_17027);
nor U24646 (N_24646,N_16310,N_18916);
xnor U24647 (N_24647,N_15410,N_15183);
or U24648 (N_24648,N_18900,N_17511);
xor U24649 (N_24649,N_18511,N_19380);
or U24650 (N_24650,N_17975,N_15788);
xnor U24651 (N_24651,N_18947,N_18148);
nor U24652 (N_24652,N_19227,N_18640);
or U24653 (N_24653,N_16542,N_15059);
and U24654 (N_24654,N_16494,N_16774);
or U24655 (N_24655,N_15864,N_19506);
or U24656 (N_24656,N_19872,N_17843);
or U24657 (N_24657,N_16333,N_16295);
and U24658 (N_24658,N_18068,N_19592);
nand U24659 (N_24659,N_17579,N_15614);
nand U24660 (N_24660,N_18950,N_19762);
and U24661 (N_24661,N_17113,N_19168);
and U24662 (N_24662,N_19768,N_15313);
or U24663 (N_24663,N_15349,N_18406);
nor U24664 (N_24664,N_15481,N_18392);
nand U24665 (N_24665,N_19076,N_18053);
nor U24666 (N_24666,N_18508,N_18525);
xnor U24667 (N_24667,N_16885,N_17584);
and U24668 (N_24668,N_19686,N_16413);
or U24669 (N_24669,N_16351,N_17564);
and U24670 (N_24670,N_17023,N_17726);
xnor U24671 (N_24671,N_19959,N_18407);
nor U24672 (N_24672,N_17485,N_17430);
or U24673 (N_24673,N_15904,N_17837);
or U24674 (N_24674,N_17257,N_15729);
nand U24675 (N_24675,N_19418,N_17145);
or U24676 (N_24676,N_16279,N_18368);
nor U24677 (N_24677,N_19396,N_15759);
or U24678 (N_24678,N_19938,N_17226);
nor U24679 (N_24679,N_16128,N_16673);
nor U24680 (N_24680,N_16184,N_18214);
and U24681 (N_24681,N_16526,N_17924);
nand U24682 (N_24682,N_15112,N_18869);
nand U24683 (N_24683,N_17250,N_19908);
nor U24684 (N_24684,N_16046,N_16352);
xnor U24685 (N_24685,N_16217,N_16501);
nand U24686 (N_24686,N_17233,N_16223);
or U24687 (N_24687,N_16902,N_17350);
xnor U24688 (N_24688,N_15982,N_19195);
or U24689 (N_24689,N_16635,N_19718);
or U24690 (N_24690,N_18196,N_15670);
and U24691 (N_24691,N_15966,N_17901);
nand U24692 (N_24692,N_19667,N_16767);
or U24693 (N_24693,N_15752,N_18711);
nor U24694 (N_24694,N_15583,N_19292);
xor U24695 (N_24695,N_15859,N_19806);
or U24696 (N_24696,N_19682,N_18394);
xor U24697 (N_24697,N_16287,N_15957);
nand U24698 (N_24698,N_19379,N_17485);
nor U24699 (N_24699,N_16239,N_18306);
and U24700 (N_24700,N_18391,N_19849);
nand U24701 (N_24701,N_15047,N_17175);
or U24702 (N_24702,N_16681,N_17687);
xnor U24703 (N_24703,N_16741,N_18269);
nand U24704 (N_24704,N_16894,N_17967);
xnor U24705 (N_24705,N_16822,N_18088);
xor U24706 (N_24706,N_18413,N_16190);
and U24707 (N_24707,N_16623,N_16638);
or U24708 (N_24708,N_16157,N_19356);
nor U24709 (N_24709,N_17717,N_15103);
nor U24710 (N_24710,N_16650,N_19743);
or U24711 (N_24711,N_18590,N_18660);
nor U24712 (N_24712,N_15175,N_19243);
or U24713 (N_24713,N_17381,N_17602);
or U24714 (N_24714,N_18965,N_17430);
xor U24715 (N_24715,N_17028,N_16497);
nand U24716 (N_24716,N_15786,N_19889);
or U24717 (N_24717,N_18341,N_15272);
nor U24718 (N_24718,N_18399,N_17977);
or U24719 (N_24719,N_16090,N_16307);
nor U24720 (N_24720,N_17148,N_16284);
and U24721 (N_24721,N_16390,N_16137);
nor U24722 (N_24722,N_18302,N_15172);
nand U24723 (N_24723,N_17736,N_15968);
nand U24724 (N_24724,N_17446,N_18544);
xnor U24725 (N_24725,N_16947,N_19448);
or U24726 (N_24726,N_17282,N_15829);
nand U24727 (N_24727,N_16791,N_17009);
and U24728 (N_24728,N_16851,N_15720);
or U24729 (N_24729,N_15844,N_17542);
nor U24730 (N_24730,N_16794,N_17384);
xor U24731 (N_24731,N_18851,N_15100);
nor U24732 (N_24732,N_18830,N_19850);
nor U24733 (N_24733,N_18609,N_17912);
nand U24734 (N_24734,N_16728,N_18142);
or U24735 (N_24735,N_17942,N_19228);
and U24736 (N_24736,N_15427,N_19903);
and U24737 (N_24737,N_16682,N_16675);
xor U24738 (N_24738,N_15308,N_15096);
nor U24739 (N_24739,N_17284,N_18074);
or U24740 (N_24740,N_16227,N_19855);
and U24741 (N_24741,N_18052,N_17015);
and U24742 (N_24742,N_18374,N_19255);
xor U24743 (N_24743,N_16773,N_19819);
nand U24744 (N_24744,N_16254,N_16895);
xor U24745 (N_24745,N_16290,N_19197);
nand U24746 (N_24746,N_17815,N_15652);
nor U24747 (N_24747,N_16272,N_18677);
and U24748 (N_24748,N_19745,N_16670);
and U24749 (N_24749,N_18362,N_19959);
and U24750 (N_24750,N_19900,N_16704);
and U24751 (N_24751,N_15126,N_17655);
or U24752 (N_24752,N_19253,N_15896);
and U24753 (N_24753,N_16394,N_15321);
or U24754 (N_24754,N_18037,N_18422);
xnor U24755 (N_24755,N_16765,N_15577);
nand U24756 (N_24756,N_19944,N_16587);
or U24757 (N_24757,N_17859,N_15633);
and U24758 (N_24758,N_18668,N_18039);
and U24759 (N_24759,N_17170,N_17491);
and U24760 (N_24760,N_18833,N_17381);
nand U24761 (N_24761,N_19739,N_18833);
xor U24762 (N_24762,N_17461,N_19907);
nand U24763 (N_24763,N_19524,N_15487);
and U24764 (N_24764,N_17772,N_15370);
nand U24765 (N_24765,N_17203,N_17117);
or U24766 (N_24766,N_17534,N_19828);
or U24767 (N_24767,N_15818,N_16199);
and U24768 (N_24768,N_16739,N_16551);
or U24769 (N_24769,N_15395,N_16613);
nand U24770 (N_24770,N_19196,N_17423);
nor U24771 (N_24771,N_16920,N_18947);
nand U24772 (N_24772,N_18637,N_16683);
xor U24773 (N_24773,N_16298,N_16106);
or U24774 (N_24774,N_15376,N_15111);
and U24775 (N_24775,N_16567,N_19097);
or U24776 (N_24776,N_19981,N_17410);
nand U24777 (N_24777,N_17534,N_17009);
nor U24778 (N_24778,N_16446,N_18360);
nor U24779 (N_24779,N_18998,N_16988);
or U24780 (N_24780,N_16881,N_15923);
and U24781 (N_24781,N_19071,N_16754);
nand U24782 (N_24782,N_15933,N_18530);
and U24783 (N_24783,N_18238,N_19258);
nor U24784 (N_24784,N_15885,N_16161);
or U24785 (N_24785,N_17623,N_19194);
and U24786 (N_24786,N_19249,N_15819);
nand U24787 (N_24787,N_19497,N_15767);
nand U24788 (N_24788,N_18423,N_17472);
and U24789 (N_24789,N_19802,N_17703);
and U24790 (N_24790,N_19702,N_19911);
or U24791 (N_24791,N_18598,N_15892);
and U24792 (N_24792,N_19312,N_17166);
xnor U24793 (N_24793,N_16649,N_18120);
nor U24794 (N_24794,N_15149,N_19352);
and U24795 (N_24795,N_19389,N_17274);
xor U24796 (N_24796,N_17775,N_17498);
nand U24797 (N_24797,N_19058,N_19381);
or U24798 (N_24798,N_17433,N_19357);
or U24799 (N_24799,N_16565,N_17714);
or U24800 (N_24800,N_16415,N_19240);
and U24801 (N_24801,N_17587,N_17939);
nand U24802 (N_24802,N_18512,N_15274);
xnor U24803 (N_24803,N_18547,N_15539);
nor U24804 (N_24804,N_17232,N_15611);
and U24805 (N_24805,N_19969,N_17577);
or U24806 (N_24806,N_19533,N_17136);
xnor U24807 (N_24807,N_16250,N_15316);
and U24808 (N_24808,N_15168,N_19397);
nor U24809 (N_24809,N_16253,N_16095);
or U24810 (N_24810,N_15336,N_15765);
or U24811 (N_24811,N_17827,N_15086);
and U24812 (N_24812,N_17701,N_19136);
or U24813 (N_24813,N_16969,N_15663);
nand U24814 (N_24814,N_17709,N_17214);
or U24815 (N_24815,N_17990,N_18854);
or U24816 (N_24816,N_16521,N_17730);
and U24817 (N_24817,N_16779,N_17101);
xor U24818 (N_24818,N_18258,N_19653);
nand U24819 (N_24819,N_15324,N_16284);
xnor U24820 (N_24820,N_16018,N_17923);
or U24821 (N_24821,N_16508,N_19558);
xor U24822 (N_24822,N_16774,N_17661);
and U24823 (N_24823,N_16135,N_17333);
nand U24824 (N_24824,N_15013,N_18615);
nor U24825 (N_24825,N_19818,N_17417);
or U24826 (N_24826,N_18059,N_15186);
nand U24827 (N_24827,N_15923,N_16529);
or U24828 (N_24828,N_16613,N_17722);
xnor U24829 (N_24829,N_16960,N_17871);
nor U24830 (N_24830,N_16505,N_19327);
and U24831 (N_24831,N_19044,N_15538);
xnor U24832 (N_24832,N_18139,N_19458);
nand U24833 (N_24833,N_17800,N_17128);
nand U24834 (N_24834,N_19111,N_16392);
nor U24835 (N_24835,N_19260,N_15732);
nor U24836 (N_24836,N_19070,N_16261);
or U24837 (N_24837,N_19329,N_18483);
nor U24838 (N_24838,N_19450,N_18702);
and U24839 (N_24839,N_15996,N_15563);
nor U24840 (N_24840,N_16254,N_15296);
nor U24841 (N_24841,N_16936,N_19629);
xor U24842 (N_24842,N_19498,N_17684);
or U24843 (N_24843,N_16839,N_16398);
and U24844 (N_24844,N_17375,N_17379);
and U24845 (N_24845,N_16929,N_16909);
xor U24846 (N_24846,N_16357,N_18452);
and U24847 (N_24847,N_19040,N_18436);
and U24848 (N_24848,N_16012,N_16362);
or U24849 (N_24849,N_15108,N_17626);
xnor U24850 (N_24850,N_19234,N_16265);
nor U24851 (N_24851,N_18500,N_19076);
or U24852 (N_24852,N_19331,N_18366);
and U24853 (N_24853,N_19858,N_18449);
or U24854 (N_24854,N_17785,N_19048);
nor U24855 (N_24855,N_16482,N_19307);
or U24856 (N_24856,N_19407,N_16773);
nor U24857 (N_24857,N_15870,N_18051);
nor U24858 (N_24858,N_18568,N_16305);
or U24859 (N_24859,N_17865,N_18922);
xnor U24860 (N_24860,N_17910,N_16295);
nor U24861 (N_24861,N_16598,N_17262);
and U24862 (N_24862,N_17561,N_17124);
xor U24863 (N_24863,N_19451,N_16331);
nand U24864 (N_24864,N_17165,N_18639);
nor U24865 (N_24865,N_15518,N_16507);
nand U24866 (N_24866,N_16661,N_19352);
nor U24867 (N_24867,N_15456,N_15376);
nand U24868 (N_24868,N_19991,N_15981);
or U24869 (N_24869,N_15934,N_16368);
xnor U24870 (N_24870,N_19475,N_17506);
nor U24871 (N_24871,N_19345,N_18676);
nor U24872 (N_24872,N_17868,N_19157);
nor U24873 (N_24873,N_16793,N_18100);
xnor U24874 (N_24874,N_15647,N_16753);
nor U24875 (N_24875,N_17778,N_17844);
xor U24876 (N_24876,N_18932,N_15103);
xor U24877 (N_24877,N_18524,N_17806);
nor U24878 (N_24878,N_19394,N_18192);
or U24879 (N_24879,N_16322,N_15631);
nand U24880 (N_24880,N_19660,N_18164);
and U24881 (N_24881,N_19063,N_19181);
or U24882 (N_24882,N_18028,N_18187);
xnor U24883 (N_24883,N_17458,N_19319);
nand U24884 (N_24884,N_18382,N_19347);
or U24885 (N_24885,N_16616,N_18101);
xnor U24886 (N_24886,N_16155,N_17607);
xor U24887 (N_24887,N_19471,N_19727);
and U24888 (N_24888,N_19405,N_17413);
nor U24889 (N_24889,N_15919,N_19071);
xor U24890 (N_24890,N_17578,N_15360);
or U24891 (N_24891,N_16991,N_18839);
nand U24892 (N_24892,N_18732,N_15600);
or U24893 (N_24893,N_15832,N_18553);
or U24894 (N_24894,N_17852,N_18652);
nand U24895 (N_24895,N_19587,N_16791);
xnor U24896 (N_24896,N_15566,N_16596);
xor U24897 (N_24897,N_15568,N_18999);
nor U24898 (N_24898,N_19992,N_16261);
xor U24899 (N_24899,N_17057,N_16724);
or U24900 (N_24900,N_17279,N_19012);
or U24901 (N_24901,N_18026,N_15473);
xor U24902 (N_24902,N_16345,N_15670);
and U24903 (N_24903,N_17110,N_18043);
and U24904 (N_24904,N_15291,N_18358);
nor U24905 (N_24905,N_19251,N_16512);
and U24906 (N_24906,N_15447,N_16442);
nor U24907 (N_24907,N_15230,N_17611);
xor U24908 (N_24908,N_17072,N_16654);
nor U24909 (N_24909,N_17872,N_17582);
and U24910 (N_24910,N_19795,N_18576);
or U24911 (N_24911,N_19731,N_19146);
xnor U24912 (N_24912,N_16574,N_19098);
nand U24913 (N_24913,N_19411,N_17126);
and U24914 (N_24914,N_17118,N_16189);
xor U24915 (N_24915,N_15449,N_17859);
xnor U24916 (N_24916,N_19343,N_16023);
xnor U24917 (N_24917,N_18711,N_15874);
or U24918 (N_24918,N_16818,N_15746);
nand U24919 (N_24919,N_15298,N_15949);
xnor U24920 (N_24920,N_19544,N_17290);
nand U24921 (N_24921,N_18881,N_15582);
and U24922 (N_24922,N_18511,N_18037);
or U24923 (N_24923,N_18131,N_19421);
xnor U24924 (N_24924,N_16907,N_19007);
or U24925 (N_24925,N_18462,N_15921);
and U24926 (N_24926,N_19866,N_17789);
and U24927 (N_24927,N_17200,N_17370);
and U24928 (N_24928,N_17797,N_18047);
xor U24929 (N_24929,N_15503,N_17182);
nand U24930 (N_24930,N_16330,N_18040);
and U24931 (N_24931,N_19348,N_16532);
and U24932 (N_24932,N_19322,N_18791);
xnor U24933 (N_24933,N_19973,N_17664);
xnor U24934 (N_24934,N_17163,N_18712);
or U24935 (N_24935,N_17005,N_19659);
nor U24936 (N_24936,N_19008,N_19944);
xnor U24937 (N_24937,N_19476,N_19341);
or U24938 (N_24938,N_18326,N_16693);
or U24939 (N_24939,N_19483,N_19612);
or U24940 (N_24940,N_17642,N_19709);
or U24941 (N_24941,N_19060,N_19716);
xor U24942 (N_24942,N_16447,N_16480);
nor U24943 (N_24943,N_15193,N_19039);
nor U24944 (N_24944,N_15659,N_18507);
and U24945 (N_24945,N_16493,N_15959);
xnor U24946 (N_24946,N_18487,N_15303);
or U24947 (N_24947,N_16033,N_16419);
and U24948 (N_24948,N_18700,N_16699);
or U24949 (N_24949,N_15340,N_19567);
and U24950 (N_24950,N_16920,N_16792);
xor U24951 (N_24951,N_19156,N_18436);
nand U24952 (N_24952,N_16003,N_18643);
nand U24953 (N_24953,N_19002,N_17729);
nand U24954 (N_24954,N_16710,N_16642);
nor U24955 (N_24955,N_15192,N_19179);
nor U24956 (N_24956,N_18557,N_15201);
and U24957 (N_24957,N_17841,N_19467);
and U24958 (N_24958,N_15873,N_16494);
or U24959 (N_24959,N_19726,N_18023);
nand U24960 (N_24960,N_15674,N_18892);
and U24961 (N_24961,N_17005,N_18013);
nor U24962 (N_24962,N_18623,N_16923);
nor U24963 (N_24963,N_17561,N_15140);
nand U24964 (N_24964,N_17349,N_19609);
nand U24965 (N_24965,N_15623,N_18047);
nor U24966 (N_24966,N_18497,N_17608);
nor U24967 (N_24967,N_19913,N_15869);
nand U24968 (N_24968,N_19412,N_16046);
xnor U24969 (N_24969,N_17146,N_15100);
nand U24970 (N_24970,N_19285,N_16661);
xnor U24971 (N_24971,N_19737,N_16957);
and U24972 (N_24972,N_16006,N_17468);
and U24973 (N_24973,N_17098,N_16344);
xnor U24974 (N_24974,N_19846,N_16947);
and U24975 (N_24975,N_19172,N_19992);
and U24976 (N_24976,N_16498,N_16270);
nand U24977 (N_24977,N_17944,N_15992);
or U24978 (N_24978,N_16413,N_19003);
xnor U24979 (N_24979,N_19889,N_15754);
and U24980 (N_24980,N_18338,N_15429);
or U24981 (N_24981,N_19731,N_17636);
xnor U24982 (N_24982,N_19835,N_18817);
nor U24983 (N_24983,N_16052,N_16152);
xor U24984 (N_24984,N_16263,N_16089);
nand U24985 (N_24985,N_19052,N_16912);
and U24986 (N_24986,N_18193,N_15956);
and U24987 (N_24987,N_17870,N_17177);
nor U24988 (N_24988,N_15743,N_15304);
nor U24989 (N_24989,N_17296,N_19443);
nand U24990 (N_24990,N_15045,N_18102);
and U24991 (N_24991,N_18813,N_16610);
or U24992 (N_24992,N_18017,N_19036);
or U24993 (N_24993,N_17439,N_15702);
or U24994 (N_24994,N_18632,N_17926);
nor U24995 (N_24995,N_18504,N_18100);
nand U24996 (N_24996,N_15601,N_15646);
and U24997 (N_24997,N_17824,N_19704);
nor U24998 (N_24998,N_19045,N_19192);
or U24999 (N_24999,N_19335,N_16885);
and U25000 (N_25000,N_21338,N_21210);
and U25001 (N_25001,N_24380,N_20343);
xnor U25002 (N_25002,N_20907,N_21701);
nand U25003 (N_25003,N_24475,N_23467);
nor U25004 (N_25004,N_23783,N_24747);
and U25005 (N_25005,N_21680,N_21780);
xnor U25006 (N_25006,N_23626,N_23725);
nor U25007 (N_25007,N_23307,N_23086);
or U25008 (N_25008,N_23497,N_20715);
or U25009 (N_25009,N_20968,N_22120);
and U25010 (N_25010,N_20679,N_23125);
nand U25011 (N_25011,N_23900,N_21905);
and U25012 (N_25012,N_24326,N_21050);
and U25013 (N_25013,N_20317,N_24110);
or U25014 (N_25014,N_20632,N_23925);
xor U25015 (N_25015,N_20155,N_23686);
xnor U25016 (N_25016,N_24846,N_22311);
or U25017 (N_25017,N_22287,N_24957);
xnor U25018 (N_25018,N_20250,N_20035);
xnor U25019 (N_25019,N_21125,N_24549);
nor U25020 (N_25020,N_20914,N_22922);
or U25021 (N_25021,N_23186,N_23773);
and U25022 (N_25022,N_24715,N_21400);
and U25023 (N_25023,N_21651,N_21201);
xor U25024 (N_25024,N_20031,N_20289);
nor U25025 (N_25025,N_22407,N_20916);
xnor U25026 (N_25026,N_20197,N_20248);
nor U25027 (N_25027,N_21037,N_24302);
nand U25028 (N_25028,N_21287,N_20404);
nand U25029 (N_25029,N_24758,N_21453);
xnor U25030 (N_25030,N_24845,N_24843);
or U25031 (N_25031,N_24648,N_20295);
nor U25032 (N_25032,N_23389,N_22813);
xor U25033 (N_25033,N_24096,N_21277);
and U25034 (N_25034,N_24201,N_24241);
nor U25035 (N_25035,N_20080,N_22435);
nor U25036 (N_25036,N_24501,N_22837);
or U25037 (N_25037,N_21447,N_20508);
or U25038 (N_25038,N_22355,N_20555);
and U25039 (N_25039,N_23145,N_20334);
nand U25040 (N_25040,N_23130,N_24239);
xor U25041 (N_25041,N_22338,N_21717);
nor U25042 (N_25042,N_21902,N_22702);
nand U25043 (N_25043,N_23939,N_21845);
xor U25044 (N_25044,N_20101,N_22686);
or U25045 (N_25045,N_23396,N_20561);
and U25046 (N_25046,N_24892,N_23463);
nand U25047 (N_25047,N_20004,N_23477);
nand U25048 (N_25048,N_20626,N_21511);
or U25049 (N_25049,N_24712,N_21278);
nand U25050 (N_25050,N_21271,N_24728);
nor U25051 (N_25051,N_24935,N_24184);
nor U25052 (N_25052,N_23311,N_24809);
or U25053 (N_25053,N_23564,N_24393);
nand U25054 (N_25054,N_21907,N_23526);
nor U25055 (N_25055,N_22981,N_22148);
nand U25056 (N_25056,N_20464,N_21268);
nor U25057 (N_25057,N_22551,N_22787);
or U25058 (N_25058,N_23269,N_20461);
and U25059 (N_25059,N_22452,N_24202);
and U25060 (N_25060,N_23177,N_24351);
nor U25061 (N_25061,N_22730,N_23092);
nor U25062 (N_25062,N_21641,N_23942);
or U25063 (N_25063,N_23046,N_21814);
xor U25064 (N_25064,N_24403,N_22073);
or U25065 (N_25065,N_24799,N_24126);
nand U25066 (N_25066,N_21023,N_22770);
nand U25067 (N_25067,N_23451,N_21851);
nor U25068 (N_25068,N_24520,N_22009);
or U25069 (N_25069,N_22137,N_24702);
nand U25070 (N_25070,N_20748,N_22823);
or U25071 (N_25071,N_22664,N_23341);
nand U25072 (N_25072,N_21529,N_20521);
nor U25073 (N_25073,N_20252,N_22558);
xor U25074 (N_25074,N_24649,N_22382);
and U25075 (N_25075,N_22843,N_21904);
or U25076 (N_25076,N_24815,N_23321);
and U25077 (N_25077,N_22964,N_21618);
nor U25078 (N_25078,N_24113,N_21620);
nor U25079 (N_25079,N_24757,N_24251);
nand U25080 (N_25080,N_22912,N_21306);
or U25081 (N_25081,N_22330,N_21549);
xnor U25082 (N_25082,N_20681,N_24144);
nor U25083 (N_25083,N_22383,N_21248);
nand U25084 (N_25084,N_24359,N_20475);
xnor U25085 (N_25085,N_20862,N_23698);
or U25086 (N_25086,N_21475,N_22515);
xnor U25087 (N_25087,N_21427,N_20222);
or U25088 (N_25088,N_20579,N_24708);
and U25089 (N_25089,N_24413,N_22871);
nor U25090 (N_25090,N_23580,N_21813);
nor U25091 (N_25091,N_22775,N_24930);
nor U25092 (N_25092,N_23587,N_22283);
and U25093 (N_25093,N_20732,N_20237);
xor U25094 (N_25094,N_24456,N_21995);
xnor U25095 (N_25095,N_20009,N_20791);
nor U25096 (N_25096,N_22602,N_23677);
xor U25097 (N_25097,N_21266,N_22965);
nand U25098 (N_25098,N_20922,N_22397);
nor U25099 (N_25099,N_23600,N_22647);
xnor U25100 (N_25100,N_24968,N_23556);
or U25101 (N_25101,N_23192,N_24292);
and U25102 (N_25102,N_20361,N_22566);
or U25103 (N_25103,N_24405,N_23780);
and U25104 (N_25104,N_24940,N_20854);
nand U25105 (N_25105,N_20801,N_22053);
nand U25106 (N_25106,N_21769,N_23143);
nor U25107 (N_25107,N_24973,N_20225);
or U25108 (N_25108,N_24162,N_22935);
or U25109 (N_25109,N_23669,N_22022);
or U25110 (N_25110,N_20757,N_20772);
or U25111 (N_25111,N_21203,N_23935);
xor U25112 (N_25112,N_20457,N_23583);
or U25113 (N_25113,N_20752,N_21703);
nor U25114 (N_25114,N_22879,N_24327);
nor U25115 (N_25115,N_20196,N_20836);
nand U25116 (N_25116,N_23338,N_23855);
and U25117 (N_25117,N_21039,N_22961);
nor U25118 (N_25118,N_23482,N_24054);
xnor U25119 (N_25119,N_24841,N_21818);
or U25120 (N_25120,N_24158,N_22160);
or U25121 (N_25121,N_23344,N_24726);
xnor U25122 (N_25122,N_22252,N_23320);
and U25123 (N_25123,N_23360,N_21080);
nand U25124 (N_25124,N_21974,N_23849);
or U25125 (N_25125,N_22521,N_22347);
xnor U25126 (N_25126,N_24568,N_21736);
and U25127 (N_25127,N_23007,N_20815);
or U25128 (N_25128,N_20362,N_21114);
and U25129 (N_25129,N_24817,N_23889);
xor U25130 (N_25130,N_22932,N_20358);
nand U25131 (N_25131,N_21344,N_21094);
xor U25132 (N_25132,N_20552,N_21381);
nand U25133 (N_25133,N_24021,N_20816);
nor U25134 (N_25134,N_20443,N_24290);
xor U25135 (N_25135,N_24873,N_24451);
nor U25136 (N_25136,N_24306,N_22171);
xor U25137 (N_25137,N_24543,N_24369);
xor U25138 (N_25138,N_22531,N_20063);
xor U25139 (N_25139,N_24874,N_22848);
xnor U25140 (N_25140,N_23891,N_24447);
xor U25141 (N_25141,N_21781,N_20079);
nor U25142 (N_25142,N_23452,N_20149);
nor U25143 (N_25143,N_24333,N_21893);
nand U25144 (N_25144,N_24638,N_24134);
nor U25145 (N_25145,N_24473,N_24354);
and U25146 (N_25146,N_23947,N_20731);
xor U25147 (N_25147,N_23040,N_21759);
xor U25148 (N_25148,N_20904,N_22485);
nand U25149 (N_25149,N_21356,N_21429);
nand U25150 (N_25150,N_20071,N_20995);
or U25151 (N_25151,N_23220,N_23206);
xor U25152 (N_25152,N_22379,N_24288);
or U25153 (N_25153,N_24065,N_23820);
and U25154 (N_25154,N_22234,N_23519);
xor U25155 (N_25155,N_24781,N_23712);
xor U25156 (N_25156,N_22825,N_21462);
and U25157 (N_25157,N_20852,N_24547);
and U25158 (N_25158,N_22470,N_23576);
nand U25159 (N_25159,N_21257,N_22141);
and U25160 (N_25160,N_23131,N_21745);
or U25161 (N_25161,N_20014,N_20513);
nand U25162 (N_25162,N_22088,N_22469);
nand U25163 (N_25163,N_20930,N_22896);
or U25164 (N_25164,N_20284,N_22432);
xor U25165 (N_25165,N_21127,N_24244);
xor U25166 (N_25166,N_24942,N_21329);
xor U25167 (N_25167,N_20835,N_24437);
nor U25168 (N_25168,N_20214,N_22914);
nor U25169 (N_25169,N_23739,N_24724);
xnor U25170 (N_25170,N_21697,N_23883);
nor U25171 (N_25171,N_20467,N_23645);
nor U25172 (N_25172,N_23454,N_22793);
nor U25173 (N_25173,N_24605,N_24682);
nor U25174 (N_25174,N_24350,N_22017);
or U25175 (N_25175,N_23475,N_24860);
and U25176 (N_25176,N_24989,N_22857);
nor U25177 (N_25177,N_23219,N_21831);
xor U25178 (N_25178,N_24165,N_23218);
or U25179 (N_25179,N_23383,N_21770);
and U25180 (N_25180,N_23678,N_21339);
xnor U25181 (N_25181,N_24213,N_24503);
nor U25182 (N_25182,N_22881,N_21839);
nor U25183 (N_25183,N_23872,N_23464);
nor U25184 (N_25184,N_23011,N_20094);
and U25185 (N_25185,N_24494,N_24342);
xnor U25186 (N_25186,N_20143,N_24234);
nor U25187 (N_25187,N_23696,N_20621);
nand U25188 (N_25188,N_22331,N_24535);
xnor U25189 (N_25189,N_21274,N_22677);
and U25190 (N_25190,N_22417,N_23730);
or U25191 (N_25191,N_23278,N_21358);
nor U25192 (N_25192,N_20178,N_22549);
nand U25193 (N_25193,N_21166,N_22937);
or U25194 (N_25194,N_22314,N_21619);
nand U25195 (N_25195,N_20190,N_20780);
nor U25196 (N_25196,N_20584,N_24705);
nor U25197 (N_25197,N_23648,N_24816);
xnor U25198 (N_25198,N_23680,N_21571);
nand U25199 (N_25199,N_21494,N_23410);
nor U25200 (N_25200,N_22082,N_21594);
and U25201 (N_25201,N_20814,N_23444);
and U25202 (N_25202,N_22643,N_24706);
xor U25203 (N_25203,N_24564,N_24627);
nand U25204 (N_25204,N_20719,N_21057);
xnor U25205 (N_25205,N_20246,N_21994);
nor U25206 (N_25206,N_24131,N_20740);
nand U25207 (N_25207,N_24878,N_23049);
xnor U25208 (N_25208,N_22633,N_22878);
and U25209 (N_25209,N_20060,N_21687);
or U25210 (N_25210,N_24842,N_20876);
or U25211 (N_25211,N_23861,N_20387);
nand U25212 (N_25212,N_21468,N_21198);
nor U25213 (N_25213,N_21647,N_24937);
xor U25214 (N_25214,N_22925,N_23215);
and U25215 (N_25215,N_23537,N_21724);
nor U25216 (N_25216,N_21150,N_22193);
nor U25217 (N_25217,N_21405,N_24242);
or U25218 (N_25218,N_21978,N_20838);
and U25219 (N_25219,N_21428,N_21586);
or U25220 (N_25220,N_20850,N_20733);
nand U25221 (N_25221,N_23166,N_22247);
and U25222 (N_25222,N_21378,N_22016);
nor U25223 (N_25223,N_20663,N_24196);
nand U25224 (N_25224,N_23352,N_24733);
or U25225 (N_25225,N_24429,N_21729);
nor U25226 (N_25226,N_21675,N_22737);
xor U25227 (N_25227,N_20722,N_21262);
nand U25228 (N_25228,N_22585,N_22797);
nand U25229 (N_25229,N_23949,N_23217);
nand U25230 (N_25230,N_21684,N_22303);
and U25231 (N_25231,N_21036,N_20753);
nor U25232 (N_25232,N_24471,N_22424);
xor U25233 (N_25233,N_21670,N_24656);
nor U25234 (N_25234,N_21744,N_21217);
and U25235 (N_25235,N_22007,N_23740);
nor U25236 (N_25236,N_20573,N_20504);
nor U25237 (N_25237,N_21304,N_21526);
and U25238 (N_25238,N_22044,N_23301);
and U25239 (N_25239,N_22213,N_22800);
nor U25240 (N_25240,N_20034,N_24880);
and U25241 (N_25241,N_22906,N_21798);
or U25242 (N_25242,N_22978,N_21895);
nand U25243 (N_25243,N_20634,N_22103);
nor U25244 (N_25244,N_24785,N_23536);
and U25245 (N_25245,N_21308,N_21275);
nand U25246 (N_25246,N_24961,N_24174);
or U25247 (N_25247,N_22526,N_21347);
nor U25248 (N_25248,N_22164,N_20028);
xor U25249 (N_25249,N_23366,N_21103);
nand U25250 (N_25250,N_21899,N_24563);
and U25251 (N_25251,N_23025,N_24170);
and U25252 (N_25252,N_23732,N_24291);
nor U25253 (N_25253,N_22298,N_22923);
or U25254 (N_25254,N_24977,N_21272);
nand U25255 (N_25255,N_22127,N_23837);
xnor U25256 (N_25256,N_22404,N_21504);
or U25257 (N_25257,N_22400,N_24743);
xnor U25258 (N_25258,N_22942,N_21202);
xor U25259 (N_25259,N_22608,N_24478);
nand U25260 (N_25260,N_22154,N_22586);
xor U25261 (N_25261,N_21528,N_21237);
xor U25262 (N_25262,N_23063,N_24792);
and U25263 (N_25263,N_20395,N_20432);
and U25264 (N_25264,N_20550,N_24427);
nor U25265 (N_25265,N_22673,N_24061);
nor U25266 (N_25266,N_23611,N_24896);
and U25267 (N_25267,N_22641,N_20773);
nand U25268 (N_25268,N_23319,N_20765);
nand U25269 (N_25269,N_22654,N_21291);
and U25270 (N_25270,N_21334,N_24252);
xnor U25271 (N_25271,N_20221,N_24830);
xnor U25272 (N_25272,N_23606,N_20761);
nand U25273 (N_25273,N_20966,N_22362);
nand U25274 (N_25274,N_20389,N_20675);
nor U25275 (N_25275,N_21354,N_23639);
or U25276 (N_25276,N_24399,N_24208);
nand U25277 (N_25277,N_22315,N_22835);
or U25278 (N_25278,N_22911,N_22372);
nand U25279 (N_25279,N_24348,N_20305);
nor U25280 (N_25280,N_20473,N_24640);
and U25281 (N_25281,N_20332,N_24551);
nand U25282 (N_25282,N_21360,N_23109);
nor U25283 (N_25283,N_23058,N_20596);
or U25284 (N_25284,N_23933,N_24668);
and U25285 (N_25285,N_22908,N_20172);
or U25286 (N_25286,N_20883,N_21757);
xor U25287 (N_25287,N_24111,N_21503);
or U25288 (N_25288,N_23555,N_23852);
and U25289 (N_25289,N_21969,N_24572);
xnor U25290 (N_25290,N_24738,N_24925);
nand U25291 (N_25291,N_24191,N_20342);
or U25292 (N_25292,N_21758,N_21194);
and U25293 (N_25293,N_21720,N_24883);
nand U25294 (N_25294,N_23857,N_21121);
or U25295 (N_25295,N_23658,N_23785);
xor U25296 (N_25296,N_21806,N_23068);
or U25297 (N_25297,N_24077,N_23767);
xnor U25298 (N_25298,N_24833,N_20266);
nor U25299 (N_25299,N_20900,N_21055);
and U25300 (N_25300,N_23834,N_21979);
and U25301 (N_25301,N_22539,N_23304);
nor U25302 (N_25302,N_23897,N_21686);
xor U25303 (N_25303,N_21398,N_22140);
xnor U25304 (N_25304,N_24772,N_23036);
nor U25305 (N_25305,N_24379,N_22324);
nand U25306 (N_25306,N_23892,N_23312);
xor U25307 (N_25307,N_22499,N_21542);
nand U25308 (N_25308,N_21653,N_24337);
and U25309 (N_25309,N_20769,N_23793);
and U25310 (N_25310,N_22429,N_24756);
and U25311 (N_25311,N_23898,N_24322);
xnor U25312 (N_25312,N_22919,N_22754);
or U25313 (N_25313,N_20228,N_22936);
nor U25314 (N_25314,N_21889,N_22883);
or U25315 (N_25315,N_20044,N_21833);
nor U25316 (N_25316,N_20264,N_21019);
or U25317 (N_25317,N_20407,N_20721);
or U25318 (N_25318,N_22996,N_24510);
and U25319 (N_25319,N_24836,N_20441);
or U25320 (N_25320,N_21578,N_24518);
xnor U25321 (N_25321,N_23581,N_22352);
nand U25322 (N_25322,N_21390,N_22126);
xnor U25323 (N_25323,N_21243,N_20446);
nand U25324 (N_25324,N_21954,N_21622);
or U25325 (N_25325,N_20460,N_23690);
or U25326 (N_25326,N_21858,N_21433);
nand U25327 (N_25327,N_22931,N_22812);
nor U25328 (N_25328,N_22547,N_24786);
or U25329 (N_25329,N_24667,N_20030);
and U25330 (N_25330,N_24876,N_20396);
and U25331 (N_25331,N_22744,N_21644);
and U25332 (N_25332,N_20352,N_21920);
nor U25333 (N_25333,N_23789,N_20986);
xnor U25334 (N_25334,N_24536,N_21442);
nand U25335 (N_25335,N_23911,N_24599);
or U25336 (N_25336,N_24979,N_24325);
or U25337 (N_25337,N_21220,N_20503);
and U25338 (N_25338,N_24683,N_21326);
xnor U25339 (N_25339,N_24624,N_23668);
nor U25340 (N_25340,N_20348,N_23745);
xor U25341 (N_25341,N_23372,N_21388);
and U25342 (N_25342,N_21149,N_23330);
xor U25343 (N_25343,N_24468,N_24051);
xor U25344 (N_25344,N_22629,N_23707);
and U25345 (N_25345,N_20819,N_22530);
xor U25346 (N_25346,N_23741,N_22060);
nand U25347 (N_25347,N_21609,N_20713);
nor U25348 (N_25348,N_24960,N_22105);
xnor U25349 (N_25349,N_22514,N_23239);
nand U25350 (N_25350,N_24114,N_21352);
or U25351 (N_25351,N_23212,N_20851);
and U25352 (N_25352,N_22944,N_20636);
and U25353 (N_25353,N_23345,N_22822);
nor U25354 (N_25354,N_24677,N_21715);
nand U25355 (N_25355,N_23017,N_24497);
nor U25356 (N_25356,N_20631,N_20232);
or U25357 (N_25357,N_20658,N_24571);
and U25358 (N_25358,N_23841,N_23647);
or U25359 (N_25359,N_21963,N_22589);
or U25360 (N_25360,N_24814,N_20877);
xnor U25361 (N_25361,N_23610,N_23569);
nand U25362 (N_25362,N_21942,N_22192);
nand U25363 (N_25363,N_21996,N_24927);
or U25364 (N_25364,N_21630,N_22880);
nand U25365 (N_25365,N_20567,N_20625);
and U25366 (N_25366,N_24514,N_21871);
xnor U25367 (N_25367,N_24856,N_24449);
nor U25368 (N_25368,N_20067,N_21659);
nor U25369 (N_25369,N_20770,N_20562);
nor U25370 (N_25370,N_20895,N_21059);
nor U25371 (N_25371,N_23674,N_24597);
nand U25372 (N_25372,N_21034,N_23000);
xnor U25373 (N_25373,N_21884,N_20173);
nand U25374 (N_25374,N_20470,N_21807);
xor U25375 (N_25375,N_22484,N_23931);
nor U25376 (N_25376,N_23609,N_20781);
nand U25377 (N_25377,N_21337,N_22697);
xnor U25378 (N_25378,N_21634,N_23198);
nand U25379 (N_25379,N_20427,N_23455);
or U25380 (N_25380,N_24688,N_24373);
and U25381 (N_25381,N_23318,N_22136);
xor U25382 (N_25382,N_22768,N_20591);
xnor U25383 (N_25383,N_24607,N_22674);
or U25384 (N_25384,N_24278,N_22885);
nor U25385 (N_25385,N_24538,N_22444);
nor U25386 (N_25386,N_23421,N_22181);
xnor U25387 (N_25387,N_23965,N_21739);
and U25388 (N_25388,N_24608,N_24911);
nand U25389 (N_25389,N_21797,N_24284);
nand U25390 (N_25390,N_21976,N_22389);
nor U25391 (N_25391,N_21345,N_23627);
xor U25392 (N_25392,N_21231,N_22257);
xnor U25393 (N_25393,N_21990,N_20527);
nor U25394 (N_25394,N_21200,N_21443);
and U25395 (N_25395,N_22058,N_21196);
and U25396 (N_25396,N_21908,N_21776);
or U25397 (N_25397,N_21108,N_22246);
nor U25398 (N_25398,N_21558,N_20202);
and U25399 (N_25399,N_20130,N_21363);
nand U25400 (N_25400,N_22190,N_20253);
or U25401 (N_25401,N_22312,N_24894);
nor U25402 (N_25402,N_20656,N_24450);
and U25403 (N_25403,N_22357,N_20614);
nor U25404 (N_25404,N_20698,N_24793);
and U25405 (N_25405,N_20365,N_21535);
nand U25406 (N_25406,N_24149,N_21302);
or U25407 (N_25407,N_20442,N_22087);
xnor U25408 (N_25408,N_24273,N_24026);
and U25409 (N_25409,N_20159,N_21449);
nand U25410 (N_25410,N_22161,N_24039);
nor U25411 (N_25411,N_21731,N_22256);
nand U25412 (N_25412,N_22745,N_24466);
nor U25413 (N_25413,N_22900,N_22591);
and U25414 (N_25414,N_22316,N_24614);
and U25415 (N_25415,N_24754,N_23187);
nand U25416 (N_25416,N_24674,N_24341);
and U25417 (N_25417,N_23866,N_23507);
nor U25418 (N_25418,N_21455,N_20008);
xnor U25419 (N_25419,N_24859,N_22143);
or U25420 (N_25420,N_23434,N_23015);
or U25421 (N_25421,N_23620,N_23742);
xor U25422 (N_25422,N_22669,N_21669);
or U25423 (N_25423,N_21877,N_22275);
nor U25424 (N_25424,N_22820,N_24981);
xor U25425 (N_25425,N_24151,N_21014);
or U25426 (N_25426,N_22508,N_22663);
xor U25427 (N_25427,N_21681,N_21683);
nand U25428 (N_25428,N_24159,N_21608);
and U25429 (N_25429,N_21250,N_20236);
nand U25430 (N_25430,N_23458,N_23332);
xor U25431 (N_25431,N_23932,N_24912);
xor U25432 (N_25432,N_23769,N_24818);
nor U25433 (N_25433,N_24179,N_23817);
and U25434 (N_25434,N_20800,N_23168);
nor U25435 (N_25435,N_21318,N_20818);
and U25436 (N_25436,N_24410,N_20022);
xnor U25437 (N_25437,N_23176,N_22267);
nand U25438 (N_25438,N_23466,N_23560);
or U25439 (N_25439,N_23847,N_22179);
xor U25440 (N_25440,N_22015,N_21525);
nand U25441 (N_25441,N_20370,N_22476);
nor U25442 (N_25442,N_23384,N_23209);
nor U25443 (N_25443,N_22985,N_22971);
xor U25444 (N_25444,N_21279,N_22755);
or U25445 (N_25445,N_24442,N_20505);
or U25446 (N_25446,N_20779,N_23542);
and U25447 (N_25447,N_22619,N_23704);
and U25448 (N_25448,N_22304,N_21434);
xor U25449 (N_25449,N_23438,N_23886);
and U25450 (N_25450,N_24691,N_22785);
or U25451 (N_25451,N_21546,N_22994);
and U25452 (N_25452,N_24370,N_23809);
nand U25453 (N_25453,N_21224,N_21154);
and U25454 (N_25454,N_22297,N_23994);
nor U25455 (N_25455,N_23548,N_24014);
nand U25456 (N_25456,N_23634,N_22263);
or U25457 (N_25457,N_20689,N_23098);
or U25458 (N_25458,N_23033,N_22278);
and U25459 (N_25459,N_20585,N_20211);
nor U25460 (N_25460,N_23349,N_22611);
or U25461 (N_25461,N_23520,N_23671);
nand U25462 (N_25462,N_23363,N_24097);
and U25463 (N_25463,N_21855,N_21496);
nor U25464 (N_25464,N_23608,N_23364);
nor U25465 (N_25465,N_23087,N_22555);
and U25466 (N_25466,N_21577,N_20472);
nand U25467 (N_25467,N_24040,N_20341);
xor U25468 (N_25468,N_20962,N_20433);
or U25469 (N_25469,N_22231,N_21973);
nor U25470 (N_25470,N_23588,N_24240);
or U25471 (N_25471,N_21104,N_23736);
nand U25472 (N_25472,N_22725,N_20996);
xnor U25473 (N_25473,N_24978,N_23916);
and U25474 (N_25474,N_23779,N_24493);
nand U25475 (N_25475,N_20247,N_20045);
nor U25476 (N_25476,N_22036,N_24323);
nor U25477 (N_25477,N_23664,N_22600);
nand U25478 (N_25478,N_22373,N_21320);
and U25479 (N_25479,N_24328,N_21408);
xor U25480 (N_25480,N_22572,N_23004);
xor U25481 (N_25481,N_20314,N_21301);
xnor U25482 (N_25482,N_20350,N_23147);
xor U25483 (N_25483,N_22112,N_20337);
nor U25484 (N_25484,N_23163,N_23371);
or U25485 (N_25485,N_23150,N_21325);
or U25486 (N_25486,N_21752,N_20351);
xnor U25487 (N_25487,N_20582,N_22237);
or U25488 (N_25488,N_20428,N_23298);
nand U25489 (N_25489,N_23061,N_21903);
and U25490 (N_25490,N_24390,N_24434);
nor U25491 (N_25491,N_23257,N_23408);
nand U25492 (N_25492,N_20360,N_21848);
nor U25493 (N_25493,N_22715,N_24005);
and U25494 (N_25494,N_23532,N_22945);
xor U25495 (N_25495,N_23182,N_23578);
or U25496 (N_25496,N_20414,N_22229);
nand U25497 (N_25497,N_23090,N_23322);
and U25498 (N_25498,N_24718,N_23012);
nand U25499 (N_25499,N_20560,N_20873);
or U25500 (N_25500,N_22228,N_21560);
or U25501 (N_25501,N_20881,N_22415);
or U25502 (N_25502,N_21095,N_24573);
xor U25503 (N_25503,N_24188,N_24559);
and U25504 (N_25504,N_24237,N_20964);
nor U25505 (N_25505,N_24676,N_22030);
nor U25506 (N_25506,N_22690,N_21371);
xor U25507 (N_25507,N_23869,N_20615);
and U25508 (N_25508,N_20323,N_22765);
xor U25509 (N_25509,N_23631,N_23735);
xor U25510 (N_25510,N_21552,N_21915);
nand U25511 (N_25511,N_20321,N_22367);
nor U25512 (N_25512,N_20794,N_21881);
xor U25513 (N_25513,N_20669,N_21621);
xnor U25514 (N_25514,N_20706,N_22013);
nor U25515 (N_25515,N_21513,N_23447);
nand U25516 (N_25516,N_21259,N_20813);
nand U25517 (N_25517,N_20339,N_22834);
xor U25518 (N_25518,N_21977,N_20758);
or U25519 (N_25519,N_23104,N_23006);
nor U25520 (N_25520,N_21501,N_23895);
xor U25521 (N_25521,N_20601,N_24049);
and U25522 (N_25522,N_24087,N_21585);
nand U25523 (N_25523,N_23411,N_22700);
nand U25524 (N_25524,N_24820,N_24224);
nor U25525 (N_25525,N_20240,N_23443);
xnor U25526 (N_25526,N_23323,N_20019);
nand U25527 (N_25527,N_21040,N_21472);
and U25528 (N_25528,N_20090,N_21256);
nor U25529 (N_25529,N_24367,N_24931);
or U25530 (N_25530,N_20534,N_24245);
and U25531 (N_25531,N_21763,N_20574);
nor U25532 (N_25532,N_21938,N_23778);
and U25533 (N_25533,N_23227,N_20647);
and U25534 (N_25534,N_20064,N_22443);
nand U25535 (N_25535,N_23175,N_24173);
nor U25536 (N_25536,N_24455,N_24336);
nor U25537 (N_25537,N_20287,N_23433);
or U25538 (N_25538,N_23416,N_22119);
nand U25539 (N_25539,N_23689,N_22040);
xor U25540 (N_25540,N_23709,N_23201);
nor U25541 (N_25541,N_20501,N_24362);
xor U25542 (N_25542,N_23409,N_22958);
nor U25543 (N_25543,N_22474,N_24382);
xor U25544 (N_25544,N_22221,N_23544);
nor U25545 (N_25545,N_23442,N_23111);
and U25546 (N_25546,N_21241,N_24117);
nand U25547 (N_25547,N_22434,N_24433);
and U25548 (N_25548,N_24834,N_20171);
and U25549 (N_25549,N_23357,N_20898);
nand U25550 (N_25550,N_21945,N_21471);
or U25551 (N_25551,N_20061,N_23602);
or U25552 (N_25552,N_21636,N_20861);
nor U25553 (N_25553,N_23010,N_20454);
nor U25554 (N_25554,N_22805,N_23285);
xor U25555 (N_25555,N_21948,N_24454);
nor U25556 (N_25556,N_24219,N_24618);
xnor U25557 (N_25557,N_22346,N_22248);
xor U25558 (N_25558,N_23958,N_22489);
nand U25559 (N_25559,N_22983,N_22081);
xor U25560 (N_25560,N_24907,N_21965);
nand U25561 (N_25561,N_20886,N_22203);
and U25562 (N_25562,N_21869,N_23469);
nand U25563 (N_25563,N_24345,N_20107);
or U25564 (N_25564,N_21239,N_21699);
nand U25565 (N_25565,N_24249,N_22209);
xor U25566 (N_25566,N_21718,N_24750);
nor U25567 (N_25567,N_23237,N_22832);
or U25568 (N_25568,N_23524,N_22128);
or U25569 (N_25569,N_23106,N_21536);
and U25570 (N_25570,N_20493,N_23595);
nor U25571 (N_25571,N_22376,N_24423);
and U25572 (N_25572,N_24589,N_20244);
xnor U25573 (N_25573,N_20548,N_20452);
nand U25574 (N_25574,N_21950,N_24787);
nor U25575 (N_25575,N_22139,N_21372);
nand U25576 (N_25576,N_22222,N_22317);
and U25577 (N_25577,N_21649,N_20313);
nor U25578 (N_25578,N_21906,N_22243);
xor U25579 (N_25579,N_24267,N_20113);
xnor U25580 (N_25580,N_23365,N_24881);
and U25581 (N_25581,N_21478,N_24698);
and U25582 (N_25582,N_20674,N_23650);
xnor U25583 (N_25583,N_22748,N_22687);
xnor U25584 (N_25584,N_20429,N_21667);
nor U25585 (N_25585,N_23770,N_23930);
and U25586 (N_25586,N_21145,N_22828);
nand U25587 (N_25587,N_20528,N_23003);
nor U25588 (N_25588,N_20609,N_21750);
nand U25589 (N_25589,N_24074,N_23851);
xor U25590 (N_25590,N_21185,N_21439);
or U25591 (N_25591,N_20078,N_20320);
nor U25592 (N_25592,N_21548,N_21107);
and U25593 (N_25593,N_20724,N_21747);
or U25594 (N_25594,N_23952,N_20939);
nor U25595 (N_25595,N_24723,N_20388);
or U25596 (N_25596,N_20541,N_20191);
nand U25597 (N_25597,N_24299,N_21297);
xor U25598 (N_25598,N_22462,N_23506);
nand U25599 (N_25599,N_21522,N_20834);
and U25600 (N_25600,N_24693,N_23204);
and U25601 (N_25601,N_23508,N_22394);
or U25602 (N_25602,N_20077,N_20771);
or U25603 (N_25603,N_21710,N_20970);
and U25604 (N_25604,N_23687,N_21580);
xnor U25605 (N_25605,N_21212,N_22109);
or U25606 (N_25606,N_24266,N_20100);
or U25607 (N_25607,N_23430,N_20976);
nor U25608 (N_25608,N_24031,N_23055);
or U25609 (N_25609,N_20529,N_23223);
and U25610 (N_25610,N_21000,N_21315);
nor U25611 (N_25611,N_22205,N_21602);
nor U25612 (N_25612,N_24182,N_21470);
nand U25613 (N_25613,N_20076,N_24807);
and U25614 (N_25614,N_24129,N_22999);
xor U25615 (N_25615,N_21702,N_24542);
or U25616 (N_25616,N_24035,N_23252);
xnor U25617 (N_25617,N_20575,N_23792);
xnor U25618 (N_25618,N_21047,N_21097);
and U25619 (N_25619,N_20782,N_24294);
or U25620 (N_25620,N_24030,N_21063);
or U25621 (N_25621,N_22532,N_20878);
or U25622 (N_25622,N_23260,N_23944);
nand U25623 (N_25623,N_22703,N_23592);
or U25624 (N_25624,N_22503,N_23636);
and U25625 (N_25625,N_24314,N_22849);
xnor U25626 (N_25626,N_21002,N_20325);
nor U25627 (N_25627,N_24163,N_24530);
xnor U25628 (N_25628,N_21033,N_22767);
nand U25629 (N_25629,N_23814,N_21090);
xnor U25630 (N_25630,N_22699,N_24938);
nor U25631 (N_25631,N_21100,N_21070);
nand U25632 (N_25632,N_22909,N_23292);
nand U25633 (N_25633,N_22414,N_22907);
or U25634 (N_25634,N_24575,N_21461);
xor U25635 (N_25635,N_20526,N_24481);
or U25636 (N_25636,N_24192,N_24967);
nand U25637 (N_25637,N_22612,N_23976);
and U25638 (N_25638,N_22374,N_23473);
or U25639 (N_25639,N_20425,N_22003);
or U25640 (N_25640,N_24849,N_22329);
xor U25641 (N_25641,N_22313,N_23406);
or U25642 (N_25642,N_22946,N_20693);
and U25643 (N_25643,N_23830,N_22803);
nand U25644 (N_25644,N_24067,N_22156);
nand U25645 (N_25645,N_23082,N_22992);
and U25646 (N_25646,N_21208,N_21537);
nand U25647 (N_25647,N_23716,N_21794);
and U25648 (N_25648,N_22893,N_22320);
and U25649 (N_25649,N_22448,N_22116);
or U25650 (N_25650,N_22439,N_20283);
xor U25651 (N_25651,N_24917,N_24516);
or U25652 (N_25652,N_20462,N_22325);
nor U25653 (N_25653,N_23954,N_20954);
or U25654 (N_25654,N_21314,N_24356);
or U25655 (N_25655,N_24524,N_24808);
or U25656 (N_25656,N_23525,N_21178);
or U25657 (N_25657,N_20670,N_21674);
or U25658 (N_25658,N_23270,N_23843);
and U25659 (N_25659,N_20495,N_22343);
xor U25660 (N_25660,N_20037,N_22777);
nand U25661 (N_25661,N_22790,N_22875);
nor U25662 (N_25662,N_22232,N_24480);
or U25663 (N_25663,N_21423,N_20416);
xor U25664 (N_25664,N_22580,N_20056);
or U25665 (N_25665,N_21303,N_22286);
xnor U25666 (N_25666,N_24922,N_24909);
xor U25667 (N_25667,N_22261,N_20619);
nor U25668 (N_25668,N_21330,N_24866);
nand U25669 (N_25669,N_22368,N_20749);
xor U25670 (N_25670,N_24238,N_21583);
or U25671 (N_25671,N_24064,N_23918);
and U25672 (N_25672,N_20597,N_21485);
or U25673 (N_25673,N_22395,N_20537);
or U25674 (N_25674,N_22063,N_23703);
and U25675 (N_25675,N_24491,N_21003);
nor U25676 (N_25676,N_24181,N_21698);
and U25677 (N_25677,N_20292,N_23240);
and U25678 (N_25678,N_21550,N_24068);
xor U25679 (N_25679,N_20857,N_22068);
nor U25680 (N_25680,N_22486,N_23005);
and U25681 (N_25681,N_21387,N_23880);
xnor U25682 (N_25682,N_22107,N_20746);
or U25683 (N_25683,N_24741,N_21713);
xor U25684 (N_25684,N_21375,N_22125);
and U25685 (N_25685,N_22818,N_23568);
nor U25686 (N_25686,N_23070,N_20400);
nand U25687 (N_25687,N_24660,N_22356);
or U25688 (N_25688,N_22218,N_23509);
nand U25689 (N_25689,N_23375,N_23995);
or U25690 (N_25690,N_21101,N_21373);
xnor U25691 (N_25691,N_23333,N_22033);
nor U25692 (N_25692,N_22288,N_22005);
or U25693 (N_25693,N_23085,N_23643);
xor U25694 (N_25694,N_21566,N_21285);
xor U25695 (N_25695,N_20750,N_23359);
xor U25696 (N_25696,N_23663,N_24377);
nor U25697 (N_25697,N_20158,N_20979);
nor U25698 (N_25698,N_21800,N_22027);
nor U25699 (N_25699,N_22548,N_23546);
nor U25700 (N_25700,N_20200,N_20271);
or U25701 (N_25701,N_21661,N_20215);
and U25702 (N_25702,N_22245,N_23361);
nand U25703 (N_25703,N_21808,N_23461);
and U25704 (N_25704,N_24598,N_21933);
xnor U25705 (N_25705,N_21891,N_21186);
nand U25706 (N_25706,N_22511,N_23051);
or U25707 (N_25707,N_21366,N_20209);
and U25708 (N_25708,N_21465,N_20081);
nand U25709 (N_25709,N_23652,N_20307);
xor U25710 (N_25710,N_23149,N_22293);
xor U25711 (N_25711,N_24424,N_24435);
nand U25712 (N_25712,N_24098,N_21159);
nor U25713 (N_25713,N_21437,N_22227);
and U25714 (N_25714,N_22170,N_24987);
xnor U25715 (N_25715,N_23392,N_20827);
or U25716 (N_25716,N_23214,N_24361);
and U25717 (N_25717,N_21993,N_24657);
and U25718 (N_25718,N_24368,N_23059);
xor U25719 (N_25719,N_21732,N_24346);
xnor U25720 (N_25720,N_21773,N_20032);
or U25721 (N_25721,N_24349,N_23381);
nand U25722 (N_25722,N_22478,N_23534);
or U25723 (N_25723,N_22761,N_20524);
nand U25724 (N_25724,N_20844,N_24882);
xnor U25725 (N_25725,N_23593,N_20789);
nand U25726 (N_25726,N_21128,N_22829);
xor U25727 (N_25727,N_23440,N_23139);
xor U25728 (N_25728,N_22197,N_23313);
xor U25729 (N_25729,N_22804,N_24633);
nand U25730 (N_25730,N_20603,N_21071);
and U25731 (N_25731,N_21746,N_23619);
xor U25732 (N_25732,N_20517,N_21207);
or U25733 (N_25733,N_22091,N_20258);
nor U25734 (N_25734,N_23997,N_23533);
nor U25735 (N_25735,N_21975,N_23230);
or U25736 (N_25736,N_24365,N_21096);
xor U25737 (N_25737,N_24689,N_21605);
nor U25738 (N_25738,N_20376,N_22831);
or U25739 (N_25739,N_20890,N_23476);
nand U25740 (N_25740,N_22578,N_23191);
or U25741 (N_25741,N_24310,N_24630);
nor U25742 (N_25742,N_23878,N_21538);
and U25743 (N_25743,N_21520,N_20357);
or U25744 (N_25744,N_23351,N_24038);
xnor U25745 (N_25745,N_20449,N_20261);
nand U25746 (N_25746,N_21436,N_20933);
nor U25747 (N_25747,N_23835,N_22163);
xor U25748 (N_25748,N_22497,N_24613);
or U25749 (N_25749,N_23398,N_23102);
nor U25750 (N_25750,N_22671,N_23823);
xnor U25751 (N_25751,N_20507,N_24444);
nor U25752 (N_25752,N_20010,N_21944);
xnor U25753 (N_25753,N_23468,N_22771);
or U25754 (N_25754,N_23799,N_21444);
and U25755 (N_25755,N_22494,N_23955);
xor U25756 (N_25756,N_24175,N_21565);
or U25757 (N_25757,N_21564,N_22451);
and U25758 (N_25758,N_23123,N_20036);
xnor U25759 (N_25759,N_20511,N_22123);
or U25760 (N_25760,N_21073,N_24000);
or U25761 (N_25761,N_24840,N_21596);
nand U25762 (N_25762,N_21650,N_20843);
nand U25763 (N_25763,N_21006,N_23500);
or U25764 (N_25764,N_21931,N_24993);
nor U25765 (N_25765,N_22199,N_23448);
nor U25766 (N_25766,N_20841,N_21861);
and U25767 (N_25767,N_22627,N_21888);
nor U25768 (N_25768,N_24763,N_24462);
xnor U25769 (N_25769,N_21812,N_24512);
nor U25770 (N_25770,N_23303,N_20269);
or U25771 (N_25771,N_24914,N_24391);
nor U25772 (N_25772,N_20075,N_22571);
nand U25773 (N_25773,N_23990,N_23749);
nor U25774 (N_25774,N_22929,N_23487);
or U25775 (N_25775,N_22752,N_23788);
xor U25776 (N_25776,N_24220,N_23894);
and U25777 (N_25777,N_23072,N_23948);
xor U25778 (N_25778,N_22728,N_20050);
and U25779 (N_25779,N_21592,N_21817);
xor U25780 (N_25780,N_22226,N_22066);
or U25781 (N_25781,N_23450,N_24602);
and U25782 (N_25782,N_24166,N_23937);
nor U25783 (N_25783,N_20199,N_24432);
nor U25784 (N_25784,N_24947,N_21819);
and U25785 (N_25785,N_22806,N_23554);
or U25786 (N_25786,N_22189,N_24190);
and U25787 (N_25787,N_24958,N_23181);
nor U25788 (N_25788,N_22817,N_21587);
or U25789 (N_25789,N_21517,N_22723);
xnor U25790 (N_25790,N_24225,N_22726);
or U25791 (N_25791,N_21838,N_23945);
xor U25792 (N_25792,N_20126,N_24171);
nand U25793 (N_25793,N_20254,N_23503);
or U25794 (N_25794,N_22024,N_24089);
nand U25795 (N_25795,N_24920,N_20047);
and U25796 (N_25796,N_23264,N_21827);
and U25797 (N_25797,N_24915,N_24470);
and U25798 (N_25798,N_21940,N_21804);
nor U25799 (N_25799,N_24483,N_21737);
nand U25800 (N_25800,N_23915,N_23453);
nand U25801 (N_25801,N_23465,N_22632);
and U25802 (N_25802,N_24015,N_20286);
nor U25803 (N_25803,N_24650,N_21678);
and U25804 (N_25804,N_23728,N_22563);
nand U25805 (N_25805,N_21119,N_24316);
nor U25806 (N_25806,N_24260,N_21043);
xnor U25807 (N_25807,N_20728,N_21643);
nor U25808 (N_25808,N_20608,N_24318);
or U25809 (N_25809,N_21021,N_24495);
and U25810 (N_25810,N_24504,N_24012);
xor U25811 (N_25811,N_21446,N_24764);
and U25812 (N_25812,N_21219,N_20532);
or U25813 (N_25813,N_24228,N_21175);
and U25814 (N_25814,N_23152,N_21980);
nand U25815 (N_25815,N_21419,N_23481);
or U25816 (N_25816,N_20088,N_21143);
nand U25817 (N_25817,N_20948,N_21755);
and U25818 (N_25818,N_20533,N_24498);
nor U25819 (N_25819,N_23327,N_20398);
nand U25820 (N_25820,N_22507,N_24945);
or U25821 (N_25821,N_24686,N_20738);
and U25822 (N_25822,N_22562,N_20089);
xnor U25823 (N_25823,N_23385,N_20542);
or U25824 (N_25824,N_23089,N_21567);
or U25825 (N_25825,N_20059,N_24643);
and U25826 (N_25826,N_23232,N_22206);
and U25827 (N_25827,N_23140,N_23665);
nor U25828 (N_25828,N_21234,N_21048);
xnor U25829 (N_25829,N_22042,N_22102);
nor U25830 (N_25830,N_22155,N_20994);
xor U25831 (N_25831,N_24212,N_20328);
nor U25832 (N_25832,N_20354,N_24687);
nand U25833 (N_25833,N_21139,N_20593);
nor U25834 (N_25834,N_23368,N_22676);
nor U25835 (N_25835,N_24477,N_24205);
or U25836 (N_25836,N_20294,N_23195);
and U25837 (N_25837,N_21012,N_20152);
nor U25838 (N_25838,N_22309,N_24593);
and U25839 (N_25839,N_20262,N_24415);
and U25840 (N_25840,N_22175,N_23585);
or U25841 (N_25841,N_20133,N_20132);
and U25842 (N_25842,N_24257,N_20563);
nand U25843 (N_25843,N_21531,N_20385);
nand U25844 (N_25844,N_23986,N_22302);
or U25845 (N_25845,N_20965,N_24558);
and U25846 (N_25846,N_21624,N_22506);
nand U25847 (N_25847,N_21440,N_21572);
nor U25848 (N_25848,N_23702,N_22061);
xor U25849 (N_25849,N_22409,N_22496);
nor U25850 (N_25850,N_23790,N_22159);
xnor U25851 (N_25851,N_20065,N_22610);
xor U25852 (N_25852,N_20445,N_21735);
or U25853 (N_25853,N_24797,N_20767);
and U25854 (N_25854,N_21309,N_23562);
nor U25855 (N_25855,N_24982,N_22386);
nor U25856 (N_25856,N_23231,N_20161);
xor U25857 (N_25857,N_24594,N_21081);
nand U25858 (N_25858,N_23504,N_21916);
nand U25859 (N_25859,N_21254,N_23906);
nor U25860 (N_25860,N_20481,N_21847);
nor U25861 (N_25861,N_20556,N_21016);
and U25862 (N_25862,N_23266,N_20399);
nor U25863 (N_25863,N_22749,N_21989);
nor U25864 (N_25864,N_23100,N_20374);
or U25865 (N_25865,N_21129,N_22930);
nor U25866 (N_25866,N_20805,N_22714);
and U25867 (N_25867,N_22370,N_24344);
xor U25868 (N_25868,N_23248,N_22705);
and U25869 (N_25869,N_20833,N_21775);
and U25870 (N_25870,N_20811,N_23484);
nor U25871 (N_25871,N_24545,N_20268);
nor U25872 (N_25872,N_22903,N_22536);
and U25873 (N_25873,N_20864,N_20616);
and U25874 (N_25874,N_23649,N_20186);
nor U25875 (N_25875,N_20496,N_22344);
xor U25876 (N_25876,N_23095,N_24279);
nor U25877 (N_25877,N_22750,N_20274);
and U25878 (N_25878,N_24851,N_23908);
and U25879 (N_25879,N_23510,N_23044);
and U25880 (N_25880,N_20847,N_21774);
xor U25881 (N_25881,N_24210,N_23300);
or U25882 (N_25882,N_21673,N_22704);
xor U25883 (N_25883,N_24672,N_24043);
nor U25884 (N_25884,N_20551,N_21987);
nor U25885 (N_25885,N_22976,N_23356);
or U25886 (N_25886,N_21679,N_24889);
and U25887 (N_25887,N_23350,N_24452);
nor U25888 (N_25888,N_21061,N_21385);
or U25889 (N_25889,N_21655,N_23822);
nor U25890 (N_25890,N_21635,N_24389);
or U25891 (N_25891,N_20899,N_22455);
nor U25892 (N_25892,N_23616,N_22020);
nand U25893 (N_25893,N_22524,N_23235);
and U25894 (N_25894,N_23567,N_20709);
xor U25895 (N_25895,N_20234,N_22729);
and U25896 (N_25896,N_24259,N_24141);
xor U25897 (N_25897,N_22262,N_22166);
xnor U25898 (N_25898,N_20666,N_21743);
nand U25899 (N_25899,N_24600,N_21654);
or U25900 (N_25900,N_23407,N_20182);
nand U25901 (N_25901,N_21335,N_21498);
xor U25902 (N_25902,N_22401,N_20412);
and U25903 (N_25903,N_21379,N_20867);
nor U25904 (N_25904,N_22588,N_22821);
nand U25905 (N_25905,N_23667,N_24078);
nand U25906 (N_25906,N_23523,N_20936);
or U25907 (N_25907,N_24888,N_24946);
and U25908 (N_25908,N_20871,N_22743);
nand U25909 (N_25909,N_22941,N_20394);
xor U25910 (N_25910,N_20417,N_24082);
xor U25911 (N_25911,N_20393,N_24254);
or U25912 (N_25912,N_24848,N_24929);
or U25913 (N_25913,N_24297,N_22609);
nand U25914 (N_25914,N_22076,N_24628);
or U25915 (N_25915,N_21102,N_21131);
and U25916 (N_25916,N_22402,N_22955);
xor U25917 (N_25917,N_23317,N_23615);
nand U25918 (N_25918,N_22393,N_23874);
and U25919 (N_25919,N_20678,N_23659);
and U25920 (N_25920,N_22235,N_23437);
xor U25921 (N_25921,N_23279,N_23165);
nor U25922 (N_25922,N_21351,N_24709);
nand U25923 (N_25923,N_20569,N_20858);
xor U25924 (N_25924,N_23846,N_20969);
and U25925 (N_25925,N_20489,N_21632);
xor U25926 (N_25926,N_21124,N_22540);
or U25927 (N_25927,N_23638,N_22322);
nand U25928 (N_25928,N_22326,N_20007);
nand U25929 (N_25929,N_23388,N_23394);
nand U25930 (N_25930,N_24264,N_21894);
nand U25931 (N_25931,N_23622,N_22590);
nor U25932 (N_25932,N_23890,N_24893);
nor U25933 (N_25933,N_23660,N_20960);
or U25934 (N_25934,N_24626,N_20549);
nand U25935 (N_25935,N_20741,N_24645);
nand U25936 (N_25936,N_22902,N_22899);
nor U25937 (N_25937,N_23579,N_22987);
or U25938 (N_25938,N_22504,N_23193);
nand U25939 (N_25939,N_21263,N_22727);
and U25940 (N_25940,N_23250,N_23572);
nor U25941 (N_25941,N_24474,N_21395);
or U25942 (N_25942,N_21728,N_21778);
and U25943 (N_25943,N_20311,N_24801);
or U25944 (N_25944,N_21183,N_20581);
nand U25945 (N_25945,N_21676,N_24570);
nor U25946 (N_25946,N_24137,N_21843);
or U25947 (N_25947,N_20998,N_24420);
or U25948 (N_25948,N_24147,N_23305);
xnor U25949 (N_25949,N_20151,N_20540);
and U25950 (N_25950,N_22388,N_24829);
or U25951 (N_25951,N_24658,N_24319);
nand U25952 (N_25952,N_24457,N_24759);
xor U25953 (N_25953,N_23733,N_21971);
nor U25954 (N_25954,N_20826,N_22480);
and U25955 (N_25955,N_24443,N_23752);
or U25956 (N_25956,N_24905,N_23013);
nand U25957 (N_25957,N_21852,N_20606);
and U25958 (N_25958,N_22233,N_21913);
nor U25959 (N_25959,N_23553,N_24387);
nor U25960 (N_25960,N_20982,N_23535);
xnor U25961 (N_25961,N_22670,N_21482);
and U25962 (N_25962,N_23575,N_22989);
nor U25963 (N_25963,N_21660,N_21109);
and U25964 (N_25964,N_24127,N_20296);
nand U25965 (N_25965,N_21300,N_23538);
nor U25966 (N_25966,N_22032,N_24928);
nor U25967 (N_25967,N_23387,N_22230);
and U25968 (N_25968,N_23956,N_23968);
and U25969 (N_25969,N_20108,N_23826);
or U25970 (N_25970,N_24421,N_21601);
nand U25971 (N_25971,N_23545,N_23970);
nand U25972 (N_25972,N_22634,N_20992);
xnor U25973 (N_25973,N_22427,N_22943);
nand U25974 (N_25974,N_21579,N_20928);
nand U25975 (N_25975,N_24554,N_20293);
or U25976 (N_25976,N_20419,N_23670);
xor U25977 (N_25977,N_20344,N_24232);
and U25978 (N_25978,N_23419,N_22887);
nor U25979 (N_25979,N_20639,N_24746);
and U25980 (N_25980,N_22988,N_23244);
and U25981 (N_25981,N_24340,N_22475);
or U25982 (N_25982,N_20822,N_23586);
or U25983 (N_25983,N_24661,N_20583);
nor U25984 (N_25984,N_21910,N_20580);
or U25985 (N_25985,N_24822,N_24751);
xor U25986 (N_25986,N_20330,N_20451);
and U25987 (N_25987,N_22465,N_20068);
nor U25988 (N_25988,N_21288,N_24321);
nand U25989 (N_25989,N_24177,N_21521);
xor U25990 (N_25990,N_21508,N_23642);
and U25991 (N_25991,N_23914,N_22463);
nand U25992 (N_25992,N_23274,N_21581);
nor U25993 (N_25993,N_23589,N_23832);
or U25994 (N_25994,N_24865,N_20853);
xor U25995 (N_25995,N_20499,N_22333);
nand U25996 (N_25996,N_24143,N_21486);
nand U25997 (N_25997,N_24867,N_23991);
nor U25998 (N_25998,N_20318,N_22072);
and U25999 (N_25999,N_23584,N_20525);
or U26000 (N_26000,N_21983,N_22963);
and U26001 (N_26001,N_23124,N_22271);
or U26002 (N_26002,N_21317,N_21075);
or U26003 (N_26003,N_23919,N_22701);
nor U26004 (N_26004,N_22212,N_22490);
and U26005 (N_26005,N_22518,N_23653);
nand U26006 (N_26006,N_20949,N_23378);
xor U26007 (N_26007,N_24167,N_20630);
or U26008 (N_26008,N_22618,N_21432);
and U26009 (N_26009,N_20256,N_20140);
nand U26010 (N_26010,N_20983,N_22290);
nand U26011 (N_26011,N_22079,N_24740);
xor U26012 (N_26012,N_20324,N_23400);
or U26013 (N_26013,N_22605,N_20944);
xnor U26014 (N_26014,N_21349,N_22795);
xnor U26015 (N_26015,N_21955,N_22108);
nand U26016 (N_26016,N_24066,N_21726);
nand U26017 (N_26017,N_22277,N_24075);
or U26018 (N_26018,N_21595,N_24303);
nor U26019 (N_26019,N_22351,N_24148);
nor U26020 (N_26020,N_22214,N_24044);
and U26021 (N_26021,N_24659,N_21087);
nor U26022 (N_26022,N_20123,N_21284);
or U26023 (N_26023,N_20298,N_24103);
nand U26024 (N_26024,N_21264,N_21790);
xor U26025 (N_26025,N_22791,N_21312);
nor U26026 (N_26026,N_22085,N_21067);
nor U26027 (N_26027,N_23179,N_24231);
and U26028 (N_26028,N_22692,N_20270);
or U26029 (N_26029,N_22816,N_22138);
xor U26030 (N_26030,N_23441,N_24317);
nor U26031 (N_26031,N_20913,N_22861);
or U26032 (N_26032,N_23295,N_21168);
and U26033 (N_26033,N_23242,N_23695);
nand U26034 (N_26034,N_20310,N_24261);
nand U26035 (N_26035,N_20547,N_22180);
xor U26036 (N_26036,N_23393,N_20477);
nor U26037 (N_26037,N_20825,N_24186);
xor U26038 (N_26038,N_21957,N_23119);
or U26039 (N_26039,N_20483,N_20338);
nor U26040 (N_26040,N_24534,N_20381);
nor U26041 (N_26041,N_21665,N_21850);
nor U26042 (N_26042,N_21140,N_22568);
nor U26043 (N_26043,N_20167,N_22915);
xnor U26044 (N_26044,N_23753,N_20622);
and U26045 (N_26045,N_23208,N_24045);
xnor U26046 (N_26046,N_24304,N_22841);
nand U26047 (N_26047,N_23802,N_20884);
nand U26048 (N_26048,N_23329,N_24305);
and U26049 (N_26049,N_21859,N_24085);
nand U26050 (N_26050,N_24651,N_24332);
nor U26051 (N_26051,N_23121,N_24145);
xor U26052 (N_26052,N_24189,N_24375);
nor U26053 (N_26053,N_21225,N_21867);
xnor U26054 (N_26054,N_22459,N_23184);
nand U26055 (N_26055,N_20418,N_20012);
or U26056 (N_26056,N_23934,N_24788);
xnor U26057 (N_26057,N_21116,N_24057);
or U26058 (N_26058,N_21172,N_24487);
xnor U26059 (N_26059,N_24198,N_24780);
nor U26060 (N_26060,N_21169,N_20423);
xnor U26061 (N_26061,N_21509,N_23893);
xnor U26062 (N_26062,N_21860,N_24532);
nand U26063 (N_26063,N_24206,N_20744);
xor U26064 (N_26064,N_21935,N_22662);
and U26065 (N_26065,N_22984,N_20198);
or U26066 (N_26066,N_23527,N_20275);
xor U26067 (N_26067,N_24722,N_20657);
nand U26068 (N_26068,N_21811,N_20903);
and U26069 (N_26069,N_21826,N_22972);
and U26070 (N_26070,N_22646,N_22450);
nor U26071 (N_26071,N_20408,N_24696);
or U26072 (N_26072,N_23748,N_24315);
or U26073 (N_26073,N_20643,N_20029);
nor U26074 (N_26074,N_22786,N_20566);
nor U26075 (N_26075,N_21953,N_23079);
xnor U26076 (N_26076,N_21582,N_24523);
xor U26077 (N_26077,N_24519,N_24301);
nor U26078 (N_26078,N_23924,N_24431);
xnor U26079 (N_26079,N_23761,N_22559);
xnor U26080 (N_26080,N_21570,N_23096);
xnor U26081 (N_26081,N_20359,N_24133);
and U26082 (N_26082,N_20764,N_21082);
xnor U26083 (N_26083,N_22062,N_21111);
xnor U26084 (N_26084,N_21421,N_22920);
nor U26085 (N_26085,N_21425,N_22974);
nand U26086 (N_26086,N_22620,N_21705);
and U26087 (N_26087,N_24070,N_21633);
xnor U26088 (N_26088,N_21384,N_20491);
nor U26089 (N_26089,N_24209,N_22651);
nor U26090 (N_26090,N_23084,N_23062);
or U26091 (N_26091,N_23249,N_20824);
xnor U26092 (N_26092,N_22440,N_23621);
xnor U26093 (N_26093,N_21193,N_22869);
and U26094 (N_26094,N_23097,N_20565);
xnor U26095 (N_26095,N_22173,N_22157);
xor U26096 (N_26096,N_22980,N_22187);
xor U26097 (N_26097,N_23864,N_22552);
nor U26098 (N_26098,N_21816,N_23076);
xnor U26099 (N_26099,N_23683,N_23644);
or U26100 (N_26100,N_20353,N_22223);
or U26101 (N_26101,N_20492,N_22874);
nor U26102 (N_26102,N_23491,N_24417);
and U26103 (N_26103,N_24953,N_20183);
xnor U26104 (N_26104,N_24274,N_21206);
nand U26105 (N_26105,N_24844,N_21348);
nor U26106 (N_26106,N_20345,N_24579);
xnor U26107 (N_26107,N_23328,N_24255);
nand U26108 (N_26108,N_23973,N_21960);
and U26109 (N_26109,N_24522,N_23921);
nand U26110 (N_26110,N_21880,N_20397);
nor U26111 (N_26111,N_24422,N_23868);
nand U26112 (N_26112,N_21885,N_21554);
nand U26113 (N_26113,N_20777,N_24974);
or U26114 (N_26114,N_21949,N_23422);
xnor U26115 (N_26115,N_22998,N_23486);
nand U26116 (N_26116,N_24666,N_23008);
nor U26117 (N_26117,N_22527,N_23805);
or U26118 (N_26118,N_24581,N_21490);
or U26119 (N_26119,N_24353,N_23386);
nand U26120 (N_26120,N_22711,N_22653);
nor U26121 (N_26121,N_20377,N_23136);
xor U26122 (N_26122,N_20879,N_24339);
nand U26123 (N_26123,N_21286,N_23699);
xnor U26124 (N_26124,N_22819,N_23662);
nand U26125 (N_26125,N_20069,N_24669);
xor U26126 (N_26126,N_20426,N_20242);
xnor U26127 (N_26127,N_20229,N_24791);
nand U26128 (N_26128,N_22405,N_21555);
nand U26129 (N_26129,N_20164,N_24187);
and U26130 (N_26130,N_20759,N_24157);
nor U26131 (N_26131,N_21401,N_20485);
nor U26132 (N_26132,N_21982,N_23777);
or U26133 (N_26133,N_22779,N_21959);
or U26134 (N_26134,N_23024,N_20568);
xor U26135 (N_26135,N_22318,N_21431);
xnor U26136 (N_26136,N_21952,N_21112);
nor U26137 (N_26137,N_24944,N_23559);
or U26138 (N_26138,N_20987,N_24539);
nor U26139 (N_26139,N_21574,N_20712);
and U26140 (N_26140,N_22661,N_22657);
or U26141 (N_26141,N_23679,N_21170);
or U26142 (N_26142,N_24169,N_22952);
nor U26143 (N_26143,N_21229,N_22467);
or U26144 (N_26144,N_21062,N_23427);
xnor U26145 (N_26145,N_22436,N_21900);
xnor U26146 (N_26146,N_24440,N_20830);
nor U26147 (N_26147,N_24936,N_20041);
and U26148 (N_26148,N_24861,N_21691);
or U26149 (N_26149,N_20710,N_21218);
xor U26150 (N_26150,N_23987,N_22954);
nor U26151 (N_26151,N_22973,N_22385);
and U26152 (N_26152,N_20023,N_21438);
or U26153 (N_26153,N_23722,N_22412);
nand U26154 (N_26154,N_20038,N_24779);
xor U26155 (N_26155,N_23905,N_23153);
xor U26156 (N_26156,N_23115,N_22731);
or U26157 (N_26157,N_23865,N_24537);
nor U26158 (N_26158,N_21041,N_23613);
and U26159 (N_26159,N_23972,N_22544);
xor U26160 (N_26160,N_21663,N_21415);
or U26161 (N_26161,N_24230,N_23528);
nand U26162 (N_26162,N_21753,N_22134);
xnor U26163 (N_26163,N_24895,N_24155);
nor U26164 (N_26164,N_22057,N_21411);
or U26165 (N_26165,N_22780,N_22348);
nand U26166 (N_26166,N_23337,N_20629);
and U26167 (N_26167,N_24577,N_21255);
xor U26168 (N_26168,N_21120,N_24472);
nor U26169 (N_26169,N_24013,N_24644);
xor U26170 (N_26170,N_23539,N_24023);
nor U26171 (N_26171,N_22152,N_20766);
and U26172 (N_26172,N_23927,N_22411);
and U26173 (N_26173,N_22560,N_21638);
nand U26174 (N_26174,N_23355,N_24641);
or U26175 (N_26175,N_22071,N_22788);
nor U26176 (N_26176,N_21018,N_24063);
nand U26177 (N_26177,N_22967,N_20235);
or U26178 (N_26178,N_22196,N_21926);
or U26179 (N_26179,N_24010,N_22259);
or U26180 (N_26180,N_24106,N_22332);
nand U26181 (N_26181,N_24102,N_22847);
nor U26182 (N_26182,N_23211,N_22365);
nor U26183 (N_26183,N_24414,N_23651);
xor U26184 (N_26184,N_21897,N_22616);
xor U26185 (N_26185,N_22041,N_24115);
or U26186 (N_26186,N_21091,N_21092);
and U26187 (N_26187,N_22886,N_23682);
xor U26188 (N_26188,N_24629,N_22517);
nor U26189 (N_26189,N_24926,N_24906);
nor U26190 (N_26190,N_20570,N_20208);
nor U26191 (N_26191,N_24794,N_21823);
nor U26192 (N_26192,N_23203,N_21377);
nand U26193 (N_26193,N_24042,N_24725);
nand U26194 (N_26194,N_24411,N_20188);
and U26195 (N_26195,N_23432,N_21122);
nand U26196 (N_26196,N_21227,N_21242);
and U26197 (N_26197,N_24060,N_22090);
and U26198 (N_26198,N_21260,N_24736);
and U26199 (N_26199,N_23963,N_23379);
and U26200 (N_26200,N_23065,N_23265);
xor U26201 (N_26201,N_20535,N_23103);
nor U26202 (N_26202,N_21730,N_20723);
and U26203 (N_26203,N_20699,N_22031);
nor U26204 (N_26204,N_20974,N_20276);
nand U26205 (N_26205,N_21840,N_20142);
nor U26206 (N_26206,N_21152,N_21209);
xnor U26207 (N_26207,N_20917,N_21222);
nand U26208 (N_26208,N_20058,N_24744);
xnor U26209 (N_26209,N_21748,N_21786);
xor U26210 (N_26210,N_22781,N_22037);
or U26211 (N_26211,N_24918,N_23325);
nor U26212 (N_26212,N_21469,N_23873);
nor U26213 (N_26213,N_22254,N_23693);
nand U26214 (N_26214,N_22734,N_20057);
and U26215 (N_26215,N_22276,N_20136);
and U26216 (N_26216,N_22255,N_21276);
xnor U26217 (N_26217,N_21042,N_22282);
or U26218 (N_26218,N_23254,N_20762);
or U26219 (N_26219,N_22421,N_21025);
nor U26220 (N_26220,N_20981,N_23833);
xnor U26221 (N_26221,N_23998,N_24505);
nor U26222 (N_26222,N_22926,N_22567);
or U26223 (N_26223,N_20282,N_23030);
or U26224 (N_26224,N_23967,N_20135);
and U26225 (N_26225,N_21591,N_24732);
xor U26226 (N_26226,N_24826,N_20255);
and U26227 (N_26227,N_20207,N_21084);
xor U26228 (N_26228,N_20941,N_24502);
xor U26229 (N_26229,N_24831,N_24385);
nand U26230 (N_26230,N_24397,N_21046);
and U26231 (N_26231,N_23200,N_24104);
nand U26232 (N_26232,N_24479,N_21502);
and U26233 (N_26233,N_22215,N_21677);
and U26234 (N_26234,N_20267,N_23088);
or U26235 (N_26235,N_20592,N_21639);
xnor U26236 (N_26236,N_23549,N_20333);
xnor U26237 (N_26237,N_24227,N_24850);
xor U26238 (N_26238,N_21992,N_24016);
nor U26239 (N_26239,N_24805,N_20046);
and U26240 (N_26240,N_24277,N_23655);
nor U26241 (N_26241,N_20440,N_21489);
xnor U26242 (N_26242,N_24128,N_21696);
xnor U26243 (N_26243,N_24970,N_24620);
nand U26244 (N_26244,N_24711,N_22772);
nand U26245 (N_26245,N_24080,N_23795);
or U26246 (N_26246,N_22718,N_24108);
xnor U26247 (N_26247,N_20720,N_24207);
nand U26248 (N_26248,N_24119,N_22576);
and U26249 (N_26249,N_24511,N_22319);
nand U26250 (N_26250,N_20300,N_21782);
nand U26251 (N_26251,N_21117,N_24615);
xor U26252 (N_26252,N_22202,N_20522);
xnor U26253 (N_26253,N_23839,N_22195);
nor U26254 (N_26254,N_23969,N_20103);
or U26255 (N_26255,N_24320,N_21045);
or U26256 (N_26256,N_20735,N_20660);
xor U26257 (N_26257,N_20204,N_22266);
nor U26258 (N_26258,N_21765,N_24366);
nand U26259 (N_26259,N_21961,N_20322);
nor U26260 (N_26260,N_24426,N_20373);
and U26261 (N_26261,N_21534,N_23543);
or U26262 (N_26262,N_24877,N_20479);
xor U26263 (N_26263,N_24465,N_23936);
nand U26264 (N_26264,N_23884,N_22537);
and U26265 (N_26265,N_22133,N_23489);
and U26266 (N_26266,N_22399,N_21497);
nor U26267 (N_26267,N_22208,N_21835);
or U26268 (N_26268,N_24124,N_24561);
xnor U26269 (N_26269,N_21085,N_22630);
nor U26270 (N_26270,N_22626,N_20536);
nor U26271 (N_26271,N_20027,N_22833);
or U26272 (N_26272,N_21130,N_20980);
xnor U26273 (N_26273,N_24076,N_20366);
and U26274 (N_26274,N_21282,N_20049);
nor U26275 (N_26275,N_21723,N_24601);
xnor U26276 (N_26276,N_20745,N_23275);
and U26277 (N_26277,N_20576,N_20807);
xnor U26278 (N_26278,N_21298,N_24533);
xnor U26279 (N_26279,N_20845,N_22165);
nor U26280 (N_26280,N_23910,N_22889);
and U26281 (N_26281,N_20848,N_24680);
or U26282 (N_26282,N_24910,N_20912);
and U26283 (N_26283,N_22991,N_22522);
nand U26284 (N_26284,N_22724,N_22488);
nor U26285 (N_26285,N_20233,N_23501);
nor U26286 (N_26286,N_20999,N_23540);
or U26287 (N_26287,N_20652,N_20985);
or U26288 (N_26288,N_21098,N_21413);
nor U26289 (N_26289,N_21013,N_24338);
xnor U26290 (N_26290,N_23018,N_22092);
nand U26291 (N_26291,N_23262,N_24448);
nor U26292 (N_26292,N_20950,N_22953);
or U26293 (N_26293,N_24546,N_22392);
and U26294 (N_26294,N_24286,N_21281);
xnor U26295 (N_26295,N_24409,N_23810);
nand U26296 (N_26296,N_21189,N_22274);
xor U26297 (N_26297,N_21789,N_20755);
xnor U26298 (N_26298,N_22099,N_21477);
or U26299 (N_26299,N_20201,N_23157);
nor U26300 (N_26300,N_22242,N_24868);
and U26301 (N_26301,N_21704,N_21590);
and U26302 (N_26302,N_23083,N_23734);
nor U26303 (N_26303,N_23261,N_24218);
nand U26304 (N_26304,N_23014,N_24036);
and U26305 (N_26305,N_22564,N_20375);
xor U26306 (N_26306,N_21230,N_24562);
nand U26307 (N_26307,N_23154,N_20648);
or U26308 (N_26308,N_24485,N_23493);
nor U26309 (N_26309,N_21754,N_20223);
xnor U26310 (N_26310,N_22917,N_21876);
or U26311 (N_26311,N_22456,N_23309);
and U26312 (N_26312,N_22305,N_20627);
nor U26313 (N_26313,N_23938,N_21296);
or U26314 (N_26314,N_22698,N_22279);
and U26315 (N_26315,N_20217,N_23917);
xor U26316 (N_26316,N_21195,N_21662);
nor U26317 (N_26317,N_20790,N_20309);
nand U26318 (N_26318,N_22584,N_22353);
nand U26319 (N_26319,N_21365,N_20888);
and U26320 (N_26320,N_23308,N_20921);
nand U26321 (N_26321,N_24720,N_24604);
or U26322 (N_26322,N_24496,N_21038);
nand U26323 (N_26323,N_21223,N_24178);
or U26324 (N_26324,N_20702,N_20520);
nor U26325 (N_26325,N_20379,N_23267);
nand U26326 (N_26326,N_23791,N_24009);
or U26327 (N_26327,N_23346,N_21947);
and U26328 (N_26328,N_22369,N_24272);
and U26329 (N_26329,N_24837,N_23713);
nor U26330 (N_26330,N_23429,N_21734);
or U26331 (N_26331,N_20763,N_23435);
nand U26332 (N_26332,N_23628,N_24357);
xnor U26333 (N_26333,N_24467,N_21069);
and U26334 (N_26334,N_21357,N_23577);
nor U26335 (N_26335,N_23798,N_21656);
or U26336 (N_26336,N_20742,N_20040);
xnor U26337 (N_26337,N_24081,N_20795);
nand U26338 (N_26338,N_21005,N_20413);
or U26339 (N_26339,N_23640,N_22891);
nand U26340 (N_26340,N_24699,N_23137);
nor U26341 (N_26341,N_23960,N_24734);
and U26342 (N_26342,N_21118,N_21901);
or U26343 (N_26343,N_20403,N_24731);
xor U26344 (N_26344,N_23514,N_22378);
or U26345 (N_26345,N_22149,N_21803);
nor U26346 (N_26346,N_21614,N_22569);
nand U26347 (N_26347,N_23977,N_24679);
xnor U26348 (N_26348,N_21246,N_24567);
xnor U26349 (N_26349,N_23080,N_24083);
or U26350 (N_26350,N_23117,N_23073);
xnor U26351 (N_26351,N_23859,N_21479);
nor U26352 (N_26352,N_22045,N_22145);
and U26353 (N_26353,N_24555,N_22425);
nand U26354 (N_26354,N_21998,N_20052);
or U26355 (N_26355,N_22308,N_20138);
nor U26356 (N_26356,N_21399,N_20018);
or U26357 (N_26357,N_21499,N_24132);
or U26358 (N_26358,N_24639,N_20265);
nand U26359 (N_26359,N_24419,N_24858);
xor U26360 (N_26360,N_22570,N_22349);
nor U26361 (N_26361,N_23756,N_24130);
nor U26362 (N_26362,N_20157,N_20870);
and U26363 (N_26363,N_24719,N_21943);
xnor U26364 (N_26364,N_24795,N_20812);
or U26365 (N_26365,N_22860,N_20924);
nor U26366 (N_26366,N_22582,N_24270);
or U26367 (N_26367,N_20048,N_23821);
and U26368 (N_26368,N_21327,N_23286);
nor U26369 (N_26369,N_24971,N_23158);
or U26370 (N_26370,N_22272,N_21457);
xor U26371 (N_26371,N_23120,N_20793);
and U26372 (N_26372,N_22681,N_20386);
xor U26373 (N_26373,N_20613,N_21988);
or U26374 (N_26374,N_21060,N_24969);
or U26375 (N_26375,N_21553,N_23081);
nor U26376 (N_26376,N_24717,N_21576);
nor U26377 (N_26377,N_24492,N_23985);
and U26378 (N_26378,N_22023,N_20111);
and U26379 (N_26379,N_22565,N_21236);
xor U26380 (N_26380,N_22975,N_22575);
or U26381 (N_26381,N_23590,N_24441);
or U26382 (N_26382,N_24897,N_24959);
nor U26383 (N_26383,N_23603,N_20169);
xor U26384 (N_26384,N_23077,N_22683);
nor U26385 (N_26385,N_22866,N_21464);
and U26386 (N_26386,N_21941,N_22799);
nand U26387 (N_26387,N_23291,N_23099);
nor U26388 (N_26388,N_20382,N_23724);
or U26389 (N_26389,N_20923,N_24821);
and U26390 (N_26390,N_20187,N_20653);
and U26391 (N_26391,N_23632,N_24486);
nand U26392 (N_26392,N_22258,N_22270);
nor U26393 (N_26393,N_23276,N_20799);
or U26394 (N_26394,N_21834,N_23414);
and U26395 (N_26395,N_22628,N_23676);
nand U26396 (N_26396,N_20952,N_23803);
xnor U26397 (N_26397,N_24285,N_22656);
xor U26398 (N_26398,N_23190,N_20887);
or U26399 (N_26399,N_20915,N_22086);
xor U26400 (N_26400,N_22993,N_23825);
and U26401 (N_26401,N_23993,N_20093);
xor U26402 (N_26402,N_23336,N_22327);
and U26403 (N_26403,N_23721,N_23920);
or U26404 (N_26404,N_23480,N_21607);
or U26405 (N_26405,N_22667,N_21467);
nand U26406 (N_26406,N_23928,N_20635);
and U26407 (N_26407,N_20514,N_23961);
nor U26408 (N_26408,N_24508,N_21369);
xor U26409 (N_26409,N_22018,N_20085);
nor U26410 (N_26410,N_24331,N_22682);
nand U26411 (N_26411,N_21192,N_22224);
nor U26412 (N_26412,N_23169,N_20645);
xor U26413 (N_26413,N_23078,N_20846);
nor U26414 (N_26414,N_21863,N_20680);
nand U26415 (N_26415,N_24086,N_23758);
xnor U26416 (N_26416,N_23151,N_24574);
nor U26417 (N_26417,N_22502,N_23162);
xor U26418 (N_26418,N_24976,N_23754);
and U26419 (N_26419,N_22850,N_24425);
nand U26420 (N_26420,N_23032,N_24665);
nor U26421 (N_26421,N_21476,N_21135);
or U26422 (N_26422,N_20977,N_24463);
nor U26423 (N_26423,N_23280,N_23402);
nor U26424 (N_26424,N_24394,N_24544);
xnor U26425 (N_26425,N_24569,N_20787);
or U26426 (N_26426,N_20304,N_21918);
xor U26427 (N_26427,N_22345,N_23786);
nor U26428 (N_26428,N_20642,N_22839);
or U26429 (N_26429,N_21510,N_23692);
nor U26430 (N_26430,N_21214,N_23558);
nor U26431 (N_26431,N_23901,N_21086);
or U26432 (N_26432,N_21575,N_20174);
nor U26433 (N_26433,N_20319,N_20016);
xnor U26434 (N_26434,N_24557,N_20516);
and U26435 (N_26435,N_23146,N_20589);
or U26436 (N_26436,N_24701,N_20195);
nor U26437 (N_26437,N_21331,N_22460);
and U26438 (N_26438,N_21299,N_20391);
nand U26439 (N_26439,N_21333,N_20005);
nand U26440 (N_26440,N_20956,N_23591);
nand U26441 (N_26441,N_24975,N_20756);
and U26442 (N_26442,N_23850,N_22774);
and U26443 (N_26443,N_23496,N_24112);
or U26444 (N_26444,N_20251,N_22756);
nor U26445 (N_26445,N_20122,N_22528);
xnor U26446 (N_26446,N_20519,N_24221);
or U26447 (N_26447,N_22239,N_22048);
xnor U26448 (N_26448,N_21221,N_24372);
nand U26449 (N_26449,N_23272,N_22769);
nor U26450 (N_26450,N_20156,N_21999);
and U26451 (N_26451,N_23729,N_22870);
or U26452 (N_26452,N_21215,N_20554);
xnor U26453 (N_26453,N_22065,N_23715);
or U26454 (N_26454,N_21708,N_24692);
or U26455 (N_26455,N_20828,N_23047);
xor U26456 (N_26456,N_20120,N_24802);
and U26457 (N_26457,N_23522,N_20902);
and U26458 (N_26458,N_24621,N_22979);
and U26459 (N_26459,N_24995,N_24295);
or U26460 (N_26460,N_23268,N_22685);
xor U26461 (N_26461,N_24875,N_24963);
xnor U26462 (N_26462,N_23255,N_22147);
nand U26463 (N_26463,N_24019,N_22337);
nand U26464 (N_26464,N_23273,N_20185);
xor U26465 (N_26465,N_20406,N_23828);
nor U26466 (N_26466,N_21937,N_24235);
xnor U26467 (N_26467,N_22390,N_24071);
and U26468 (N_26468,N_24018,N_24900);
and U26469 (N_26469,N_23617,N_20288);
and U26470 (N_26470,N_21235,N_20438);
or U26471 (N_26471,N_21652,N_20538);
or U26472 (N_26472,N_24774,N_21407);
xnor U26473 (N_26473,N_21402,N_20459);
or U26474 (N_26474,N_21197,N_23759);
and U26475 (N_26475,N_22542,N_23369);
nor U26476 (N_26476,N_24541,N_24901);
nor U26477 (N_26477,N_20523,N_22764);
nor U26478 (N_26478,N_21010,N_21158);
nand U26479 (N_26479,N_20165,N_21292);
nor U26480 (N_26480,N_20378,N_24022);
nor U26481 (N_26481,N_22798,N_22260);
and U26482 (N_26482,N_21481,N_23425);
or U26483 (N_26483,N_20610,N_24635);
nor U26484 (N_26484,N_23899,N_24287);
or U26485 (N_26485,N_22177,N_20530);
nor U26486 (N_26486,N_21664,N_22273);
nor U26487 (N_26487,N_22391,N_22419);
nand U26488 (N_26488,N_24515,N_21751);
xor U26489 (N_26489,N_22693,N_24402);
and U26490 (N_26490,N_23060,N_23367);
nand U26491 (N_26491,N_22865,N_23978);
and U26492 (N_26492,N_20925,N_21524);
and U26493 (N_26493,N_20181,N_23428);
or U26494 (N_26494,N_24161,N_20415);
and U26495 (N_26495,N_20243,N_23623);
or U26496 (N_26496,N_22639,N_21024);
nor U26497 (N_26497,N_22982,N_20127);
nor U26498 (N_26498,N_24289,N_21551);
xor U26499 (N_26499,N_20091,N_20651);
xor U26500 (N_26500,N_20894,N_22783);
nor U26501 (N_26501,N_23776,N_24592);
and U26502 (N_26502,N_24988,N_24739);
nor U26503 (N_26503,N_22253,N_22951);
nor U26504 (N_26504,N_20959,N_22144);
and U26505 (N_26505,N_22846,N_23755);
or U26506 (N_26506,N_24670,N_20671);
and U26507 (N_26507,N_24311,N_22471);
nand U26508 (N_26508,N_22481,N_22217);
nand U26509 (N_26509,N_21426,N_23829);
nand U26510 (N_26510,N_22607,N_22642);
xor U26511 (N_26511,N_22445,N_23701);
nand U26512 (N_26512,N_22933,N_21336);
nor U26513 (N_26513,N_24727,N_22097);
nand U26514 (N_26514,N_24140,N_24864);
xnor U26515 (N_26515,N_21011,N_21353);
or U26516 (N_26516,N_21606,N_23808);
nand U26517 (N_26517,N_20073,N_21792);
nor U26518 (N_26518,N_24047,N_21928);
nand U26519 (N_26519,N_22011,N_23666);
xor U26520 (N_26520,N_20020,N_21171);
nor U26521 (N_26521,N_23824,N_22446);
nand U26522 (N_26522,N_21065,N_24032);
nand U26523 (N_26523,N_24647,N_20055);
xor U26524 (N_26524,N_23499,N_24748);
nor U26525 (N_26525,N_21613,N_22713);
xnor U26526 (N_26526,N_23929,N_23057);
nor U26527 (N_26527,N_20993,N_22910);
or U26528 (N_26528,N_22492,N_24812);
xor U26529 (N_26529,N_24099,N_21791);
nor U26530 (N_26530,N_20011,N_23183);
nor U26531 (N_26531,N_20327,N_24771);
nand U26532 (N_26532,N_22852,N_21052);
nand U26533 (N_26533,N_22069,N_21165);
or U26534 (N_26534,N_21544,N_23784);
and U26535 (N_26535,N_24950,N_20218);
or U26536 (N_26536,N_24172,N_22186);
nand U26537 (N_26537,N_24072,N_21137);
or U26538 (N_26538,N_23382,N_23717);
and U26539 (N_26539,N_24678,N_20154);
nand U26540 (N_26540,N_21788,N_22901);
xnor U26541 (N_26541,N_23637,N_20474);
and U26542 (N_26542,N_22049,N_24223);
and U26543 (N_26543,N_23141,N_22321);
nor U26544 (N_26544,N_21404,N_21211);
and U26545 (N_26545,N_21179,N_24073);
nor U26546 (N_26546,N_24891,N_20856);
nand U26547 (N_26547,N_20092,N_23815);
xnor U26548 (N_26548,N_24972,N_22741);
xnor U26549 (N_26549,N_20875,N_21868);
nand U26550 (N_26550,N_22094,N_20347);
and U26551 (N_26551,N_22039,N_21422);
nand U26552 (N_26552,N_23376,N_24632);
nand U26553 (N_26553,N_22940,N_24954);
xor U26554 (N_26554,N_23256,N_20453);
or U26555 (N_26555,N_22447,N_20109);
nand U26556 (N_26556,N_23170,N_24507);
xnor U26557 (N_26557,N_21623,N_24752);
nor U26558 (N_26558,N_23045,N_24265);
or U26559 (N_26559,N_20624,N_24027);
and U26560 (N_26560,N_20184,N_20673);
or U26561 (N_26561,N_22167,N_22509);
nor U26562 (N_26562,N_24556,N_22201);
nor U26563 (N_26563,N_24646,N_22359);
or U26564 (N_26564,N_23474,N_20599);
or U26565 (N_26565,N_20633,N_20687);
nor U26566 (N_26566,N_23517,N_23711);
xor U26567 (N_26567,N_20466,N_21617);
nor U26568 (N_26568,N_20572,N_21530);
or U26569 (N_26569,N_22285,N_21836);
or U26570 (N_26570,N_20436,N_23478);
or U26571 (N_26571,N_24622,N_20588);
nand U26572 (N_26572,N_22520,N_24642);
or U26573 (N_26573,N_22052,N_20424);
nand U26574 (N_26574,N_22845,N_22055);
nor U26575 (N_26575,N_23697,N_24839);
and U26576 (N_26576,N_20910,N_22121);
nand U26577 (N_26577,N_24655,N_21716);
nor U26578 (N_26578,N_23277,N_21898);
nand U26579 (N_26579,N_20355,N_20210);
xor U26580 (N_26580,N_20971,N_20410);
or U26581 (N_26581,N_23996,N_24248);
or U26582 (N_26582,N_23957,N_24378);
nor U26583 (N_26583,N_20839,N_20498);
nand U26584 (N_26584,N_21247,N_21946);
nand U26585 (N_26585,N_22892,N_20785);
xnor U26586 (N_26586,N_23860,N_24489);
nor U26587 (N_26587,N_22413,N_21986);
nor U26588 (N_26588,N_23316,N_23075);
and U26589 (N_26589,N_21690,N_24253);
nand U26590 (N_26590,N_20259,N_24703);
or U26591 (N_26591,N_21562,N_20500);
nor U26592 (N_26592,N_22720,N_24490);
nor U26593 (N_26593,N_20026,N_21068);
nand U26594 (N_26594,N_21866,N_20192);
and U26595 (N_26595,N_20238,N_24933);
nand U26596 (N_26596,N_22622,N_24197);
and U26597 (N_26597,N_24902,N_21796);
and U26598 (N_26598,N_23113,N_24358);
and U26599 (N_26599,N_22100,N_22512);
and U26600 (N_26600,N_20809,N_22131);
xor U26601 (N_26601,N_20226,N_21784);
and U26602 (N_26602,N_24430,N_24782);
xor U26603 (N_26603,N_21370,N_23765);
nor U26604 (N_26604,N_22678,N_24226);
nor U26605 (N_26605,N_24376,N_24704);
or U26606 (N_26606,N_23657,N_24588);
xnor U26607 (N_26607,N_24800,N_21030);
nor U26608 (N_26608,N_21695,N_23391);
nor U26609 (N_26609,N_24037,N_21004);
nor U26610 (N_26610,N_20951,N_20897);
or U26611 (N_26611,N_23946,N_21563);
nand U26612 (N_26612,N_21310,N_23210);
and U26613 (N_26613,N_20372,N_22479);
nand U26614 (N_26614,N_21459,N_24985);
nand U26615 (N_26615,N_24335,N_20641);
nor U26616 (N_26616,N_24735,N_20823);
and U26617 (N_26617,N_20168,N_23395);
and U26618 (N_26618,N_22310,N_21887);
nor U26619 (N_26619,N_22652,N_24418);
nor U26620 (N_26620,N_24890,N_24271);
and U26621 (N_26621,N_23518,N_21153);
nor U26622 (N_26622,N_20125,N_23116);
xor U26623 (N_26623,N_22862,N_21289);
nor U26624 (N_26624,N_21914,N_23069);
or U26625 (N_26625,N_24033,N_20931);
or U26626 (N_26626,N_23782,N_21658);
nor U26627 (N_26627,N_20708,N_22464);
or U26628 (N_26628,N_21925,N_23999);
and U26629 (N_26629,N_20682,N_24753);
nand U26630 (N_26630,N_20147,N_21463);
or U26631 (N_26631,N_20896,N_21593);
xnor U26632 (N_26632,N_24469,N_23750);
or U26633 (N_26633,N_24552,N_22708);
or U26634 (N_26634,N_22956,N_24707);
and U26635 (N_26635,N_21685,N_20471);
xor U26636 (N_26636,N_24392,N_20659);
nor U26637 (N_26637,N_21970,N_24275);
nor U26638 (N_26638,N_24136,N_22601);
xnor U26639 (N_26639,N_20947,N_22225);
xnor U26640 (N_26640,N_22185,N_23171);
nand U26641 (N_26641,N_20874,N_23296);
nor U26642 (N_26642,N_23840,N_24330);
nor U26643 (N_26643,N_24250,N_22949);
or U26644 (N_26644,N_23923,N_21265);
nor U26645 (N_26645,N_23138,N_23243);
nor U26646 (N_26646,N_22054,N_24003);
nand U26647 (N_26647,N_20940,N_23196);
and U26648 (N_26648,N_22746,N_23718);
or U26649 (N_26649,N_20866,N_23844);
nand U26650 (N_26650,N_23485,N_21764);
xnor U26651 (N_26651,N_20798,N_23207);
nand U26652 (N_26652,N_22894,N_20935);
nor U26653 (N_26653,N_22694,N_20476);
nor U26654 (N_26654,N_20751,N_21027);
xnor U26655 (N_26655,N_24631,N_21589);
xor U26656 (N_26656,N_22084,N_20224);
nand U26657 (N_26657,N_22458,N_21533);
xor U26658 (N_26658,N_22265,N_23412);
or U26659 (N_26659,N_24919,N_22740);
xnor U26660 (N_26660,N_21872,N_24329);
xnor U26661 (N_26661,N_22709,N_23054);
and U26662 (N_26662,N_24983,N_21815);
nor U26663 (N_26663,N_23984,N_24293);
nand U26664 (N_26664,N_20306,N_24059);
xnor U26665 (N_26665,N_21343,N_22550);
nand U26666 (N_26666,N_24200,N_23390);
xor U26667 (N_26667,N_24020,N_23293);
nand U26668 (N_26668,N_21393,N_21406);
xnor U26669 (N_26669,N_20880,N_20170);
nor U26670 (N_26670,N_23189,N_22093);
and U26671 (N_26671,N_21322,N_21181);
nor U26672 (N_26672,N_24282,N_23812);
nor U26673 (N_26673,N_21177,N_23763);
and U26674 (N_26674,N_20356,N_23641);
xor U26675 (N_26675,N_23289,N_21216);
or U26676 (N_26676,N_23029,N_22466);
and U26677 (N_26677,N_20072,N_21760);
nand U26678 (N_26678,N_23966,N_20468);
or U26679 (N_26679,N_22380,N_20926);
and U26680 (N_26680,N_21714,N_21611);
nand U26681 (N_26681,N_21093,N_24401);
or U26682 (N_26682,N_22269,N_23056);
or U26683 (N_26683,N_21146,N_24855);
or U26684 (N_26684,N_24999,N_24585);
xor U26685 (N_26685,N_23306,N_24268);
xor U26686 (N_26686,N_21862,N_20760);
nand U26687 (N_26687,N_21919,N_23281);
xnor U26688 (N_26688,N_22153,N_20691);
or U26689 (N_26689,N_22840,N_24804);
nor U26690 (N_26690,N_21132,N_22890);
nand U26691 (N_26691,N_24135,N_21450);
and U26692 (N_26692,N_23258,N_21364);
nand U26693 (N_26693,N_23245,N_23028);
xor U26694 (N_26694,N_24091,N_20840);
or U26695 (N_26695,N_20946,N_24298);
nor U26696 (N_26696,N_20863,N_20213);
xnor U26697 (N_26697,N_21939,N_23684);
xnor U26698 (N_26698,N_24775,N_21240);
nand U26699 (N_26699,N_21126,N_24296);
nand U26700 (N_26700,N_24879,N_21625);
nand U26701 (N_26701,N_24662,N_24281);
xnor U26702 (N_26702,N_24386,N_21559);
or U26703 (N_26703,N_21772,N_22856);
nand U26704 (N_26704,N_23646,N_24307);
and U26705 (N_26705,N_23127,N_24587);
and U26706 (N_26706,N_23988,N_24591);
and U26707 (N_26707,N_24152,N_22573);
nor U26708 (N_26708,N_21934,N_24586);
nand U26709 (N_26709,N_24773,N_23470);
nor U26710 (N_26710,N_22583,N_20953);
and U26711 (N_26711,N_23107,N_23633);
and U26712 (N_26712,N_24459,N_23774);
nand U26713 (N_26713,N_24176,N_21612);
nor U26714 (N_26714,N_21911,N_21397);
nor U26715 (N_26715,N_20279,N_23173);
nor U26716 (N_26716,N_21383,N_23565);
nor U26717 (N_26717,N_24887,N_23953);
or U26718 (N_26718,N_24439,N_24526);
xor U26719 (N_26719,N_21380,N_22696);
nand U26720 (N_26720,N_22056,N_24308);
xnor U26721 (N_26721,N_20558,N_23598);
nor U26722 (N_26722,N_22535,N_23035);
nand U26723 (N_26723,N_21226,N_23449);
nor U26724 (N_26724,N_24084,N_23858);
and U26725 (N_26725,N_24011,N_23982);
xor U26726 (N_26726,N_24783,N_22660);
nor U26727 (N_26727,N_22501,N_24730);
xnor U26728 (N_26728,N_23570,N_20696);
xor U26729 (N_26729,N_22796,N_23512);
or U26730 (N_26730,N_21671,N_23881);
nand U26731 (N_26731,N_20070,N_20117);
and U26732 (N_26732,N_23630,N_21921);
or U26733 (N_26733,N_23870,N_24824);
xor U26734 (N_26734,N_24784,N_21480);
nand U26735 (N_26735,N_24811,N_24408);
nand U26736 (N_26736,N_22182,N_21396);
nor U26737 (N_26737,N_22268,N_20598);
xnor U26738 (N_26738,N_22350,N_22284);
nand U26739 (N_26739,N_20594,N_24347);
or U26740 (N_26740,N_21719,N_21615);
nand U26741 (N_26741,N_24404,N_20448);
nor U26742 (N_26742,N_24863,N_22557);
nand U26743 (N_26743,N_22244,N_23700);
and U26744 (N_26744,N_20604,N_23516);
xor U26745 (N_26745,N_21009,N_20205);
and U26746 (N_26746,N_24509,N_22706);
or U26747 (N_26747,N_20114,N_22637);
xor U26748 (N_26748,N_22135,N_23342);
nor U26749 (N_26749,N_22684,N_22449);
or U26750 (N_26750,N_21828,N_24778);
nand U26751 (N_26751,N_20371,N_23094);
and U26752 (N_26752,N_21341,N_22473);
or U26753 (N_26753,N_20677,N_20163);
and U26754 (N_26754,N_24406,N_23161);
xor U26755 (N_26755,N_23178,N_22898);
nand U26756 (N_26756,N_20628,N_22876);
nand U26757 (N_26757,N_24247,N_24857);
nand U26758 (N_26758,N_23594,N_20695);
and U26759 (N_26759,N_23247,N_20889);
xnor U26760 (N_26760,N_23672,N_23042);
nor U26761 (N_26761,N_24853,N_24488);
nand U26762 (N_26762,N_20892,N_20194);
or U26763 (N_26763,N_21321,N_20882);
or U26764 (N_26764,N_23071,N_22431);
and U26765 (N_26765,N_23573,N_22815);
nand U26766 (N_26766,N_21820,N_23705);
or U26767 (N_26767,N_22162,N_22493);
and U26768 (N_26768,N_21474,N_22115);
nand U26769 (N_26769,N_24164,N_20849);
nand U26770 (N_26770,N_22264,N_22340);
and U26771 (N_26771,N_24029,N_23229);
xnor U26772 (N_26772,N_22613,N_24790);
and U26773 (N_26773,N_22014,N_22977);
nand U26774 (N_26774,N_21824,N_22070);
and U26775 (N_26775,N_20967,N_22342);
xnor U26776 (N_26776,N_21584,N_21799);
xor U26777 (N_26777,N_20179,N_20260);
and U26778 (N_26778,N_24513,N_23738);
and U26779 (N_26779,N_22712,N_23288);
nor U26780 (N_26780,N_24767,N_23781);
nor U26781 (N_26781,N_23052,N_23862);
or U26782 (N_26782,N_21865,N_20349);
nor U26783 (N_26783,N_22811,N_20734);
nor U26784 (N_26784,N_20162,N_21640);
nor U26785 (N_26785,N_22220,N_23050);
nor U26786 (N_26786,N_20672,N_21051);
nand U26787 (N_26787,N_20099,N_22122);
and U26788 (N_26788,N_23353,N_22868);
nor U26789 (N_26789,N_21626,N_23726);
nand U26790 (N_26790,N_24055,N_23436);
nor U26791 (N_26791,N_24903,N_21445);
and U26792 (N_26792,N_21077,N_22008);
nor U26793 (N_26793,N_20153,N_23607);
or U26794 (N_26794,N_23037,N_20177);
or U26795 (N_26795,N_24653,N_20820);
nand U26796 (N_26796,N_24997,N_20134);
and U26797 (N_26797,N_22250,N_24553);
and U26798 (N_26798,N_21270,N_21280);
or U26799 (N_26799,N_21022,N_20683);
nor U26800 (N_26800,N_23335,N_23710);
or U26801 (N_26801,N_22597,N_20786);
and U26802 (N_26802,N_20488,N_22408);
or U26803 (N_26803,N_21886,N_21316);
xnor U26804 (N_26804,N_22948,N_24737);
nor U26805 (N_26805,N_20439,N_22025);
nor U26806 (N_26806,N_22751,N_21290);
nand U26807 (N_26807,N_20420,N_21642);
nor U26808 (N_26808,N_24374,N_23842);
or U26809 (N_26809,N_20402,N_24965);
xnor U26810 (N_26810,N_21232,N_23401);
or U26811 (N_26811,N_24180,N_23290);
and U26812 (N_26812,N_23221,N_24214);
and U26813 (N_26813,N_20039,N_24924);
or U26814 (N_26814,N_22064,N_22301);
and U26815 (N_26815,N_23719,N_23431);
nand U26816 (N_26816,N_22106,N_20098);
xnor U26817 (N_26817,N_22472,N_20024);
or U26818 (N_26818,N_22763,N_23856);
and U26819 (N_26819,N_20277,N_22672);
and U26820 (N_26820,N_24280,N_20543);
nor U26821 (N_26821,N_24203,N_23172);
xor U26822 (N_26822,N_20842,N_22561);
and U26823 (N_26823,N_23020,N_21779);
nand U26824 (N_26824,N_23550,N_20792);
and U26825 (N_26825,N_20963,N_20905);
nand U26826 (N_26826,N_21917,N_21058);
nor U26827 (N_26827,N_24770,N_22625);
nor U26828 (N_26828,N_22913,N_23762);
nand U26829 (N_26829,N_20564,N_20368);
nor U26830 (N_26830,N_23940,N_21054);
and U26831 (N_26831,N_21323,N_22853);
nor U26832 (N_26832,N_22500,N_23439);
or U26833 (N_26833,N_23992,N_24211);
or U26834 (N_26834,N_22118,N_22519);
nand U26835 (N_26835,N_21648,N_22281);
xnor U26836 (N_26836,N_21164,N_22650);
xor U26837 (N_26837,N_22851,N_22433);
and U26838 (N_26838,N_21599,N_20102);
or U26839 (N_26839,N_24453,N_20788);
or U26840 (N_26840,N_23629,N_20703);
or U26841 (N_26841,N_24671,N_23531);
nand U26842 (N_26842,N_20216,N_23031);
or U26843 (N_26843,N_24101,N_23871);
nand U26844 (N_26844,N_21878,N_21252);
or U26845 (N_26845,N_20001,N_21138);
or U26846 (N_26846,N_21892,N_20096);
or U26847 (N_26847,N_20578,N_23155);
nor U26848 (N_26848,N_24446,N_21148);
and U26849 (N_26849,N_24531,N_22002);
and U26850 (N_26850,N_21361,N_24609);
nand U26851 (N_26851,N_23134,N_22406);
xor U26852 (N_26852,N_24527,N_23397);
nand U26853 (N_26853,N_24006,N_22438);
xor U26854 (N_26854,N_23903,N_20062);
and U26855 (N_26855,N_20380,N_20920);
and U26856 (N_26856,N_22735,N_21157);
or U26857 (N_26857,N_22649,N_23417);
xnor U26858 (N_26858,N_21874,N_22491);
nor U26859 (N_26859,N_22624,N_21712);
nand U26860 (N_26860,N_21258,N_22722);
nor U26861 (N_26861,N_21414,N_24716);
nand U26862 (N_26862,N_22680,N_23460);
or U26863 (N_26863,N_23515,N_22240);
xor U26864 (N_26864,N_20465,N_23164);
nor U26865 (N_26865,N_20808,N_24869);
or U26866 (N_26866,N_22104,N_23597);
nor U26867 (N_26867,N_24729,N_22381);
nor U26868 (N_26868,N_24194,N_20685);
or U26869 (N_26869,N_23720,N_22468);
or U26870 (N_26870,N_21028,N_20083);
or U26871 (N_26871,N_20241,N_20336);
xnor U26872 (N_26872,N_22483,N_24923);
xor U26873 (N_26873,N_22710,N_24506);
nand U26874 (N_26874,N_24806,N_23216);
or U26875 (N_26875,N_24002,N_22758);
nor U26876 (N_26876,N_20458,N_23202);
nor U26877 (N_26877,N_21451,N_22990);
xor U26878 (N_26878,N_22615,N_21460);
nor U26879 (N_26879,N_20796,N_23326);
and U26880 (N_26880,N_22236,N_22241);
and U26881 (N_26881,N_24199,N_22966);
and U26882 (N_26882,N_20919,N_23913);
nor U26883 (N_26883,N_20405,N_20308);
nor U26884 (N_26884,N_24154,N_23979);
and U26885 (N_26885,N_22423,N_22487);
nand U26886 (N_26886,N_24636,N_21507);
and U26887 (N_26887,N_24560,N_21766);
nand U26888 (N_26888,N_24612,N_20885);
xnor U26889 (N_26889,N_21657,N_23251);
or U26890 (N_26890,N_23315,N_20017);
or U26891 (N_26891,N_21044,N_21163);
xor U26892 (N_26892,N_20553,N_21801);
nand U26893 (N_26893,N_20984,N_20329);
nand U26894 (N_26894,N_20707,N_23775);
or U26895 (N_26895,N_21294,N_20650);
xor U26896 (N_26896,N_24634,N_22738);
nand U26897 (N_26897,N_21089,N_20212);
and U26898 (N_26898,N_22921,N_20664);
nand U26899 (N_26899,N_24004,N_22577);
xor U26900 (N_26900,N_22635,N_23039);
nand U26901 (N_26901,N_24966,N_20997);
or U26902 (N_26902,N_23818,N_20545);
xnor U26903 (N_26903,N_20302,N_22636);
and U26904 (N_26904,N_20249,N_22089);
nand U26905 (N_26905,N_23836,N_21822);
nand U26906 (N_26906,N_23599,N_22430);
or U26907 (N_26907,N_20087,N_22739);
nand U26908 (N_26908,N_21199,N_22219);
or U26909 (N_26909,N_23423,N_23875);
nor U26910 (N_26910,N_23845,N_23226);
nand U26911 (N_26911,N_24482,N_23896);
nand U26912 (N_26912,N_23002,N_23827);
or U26913 (N_26913,N_21749,N_22810);
xor U26914 (N_26914,N_22323,N_21049);
or U26915 (N_26915,N_24312,N_24384);
and U26916 (N_26916,N_22207,N_22498);
or U26917 (N_26917,N_22553,N_20768);
xor U26918 (N_26918,N_20124,N_24625);
xor U26919 (N_26919,N_24525,N_23488);
and U26920 (N_26920,N_23283,N_20705);
or U26921 (N_26921,N_24094,N_24395);
and U26922 (N_26922,N_21767,N_20961);
nand U26923 (N_26923,N_22461,N_21929);
nor U26924 (N_26924,N_24681,N_23853);
nor U26925 (N_26925,N_20227,N_23757);
xor U26926 (N_26926,N_21389,N_20340);
xor U26927 (N_26927,N_24899,N_21603);
xnor U26928 (N_26928,N_24217,N_23128);
and U26929 (N_26929,N_23347,N_24460);
nor U26930 (N_26930,N_23975,N_22198);
nor U26931 (N_26931,N_20401,N_23253);
nand U26932 (N_26932,N_24710,N_20316);
nor U26933 (N_26933,N_23233,N_22169);
and U26934 (N_26934,N_20837,N_20700);
nand U26935 (N_26935,N_23413,N_20623);
xnor U26936 (N_26936,N_20711,N_22807);
nor U26937 (N_26937,N_21825,N_21188);
and U26938 (N_26938,N_21495,N_24885);
xor U26939 (N_26939,N_24932,N_24243);
nand U26940 (N_26940,N_24992,N_21064);
xor U26941 (N_26941,N_22124,N_24381);
nand U26942 (N_26942,N_22939,N_24813);
or U26943 (N_26943,N_20991,N_23681);
nand U26944 (N_26944,N_21527,N_20717);
or U26945 (N_26945,N_22296,N_20299);
and U26946 (N_26946,N_23807,N_20180);
or U26947 (N_26947,N_24986,N_21367);
nand U26948 (N_26948,N_21689,N_20929);
nand U26949 (N_26949,N_22191,N_20422);
or U26950 (N_26950,N_21191,N_24053);
nand U26951 (N_26951,N_22759,N_24309);
and U26952 (N_26952,N_20421,N_22210);
xnor U26953 (N_26953,N_21167,N_20335);
nand U26954 (N_26954,N_23746,N_23571);
nand U26955 (N_26955,N_20013,N_22132);
or U26956 (N_26956,N_23530,N_23563);
and U26957 (N_26957,N_20509,N_22604);
nand U26958 (N_26958,N_23904,N_23582);
nand U26959 (N_26959,N_20312,N_20434);
xnor U26960 (N_26960,N_24146,N_23926);
and U26961 (N_26961,N_21340,N_22251);
xor U26962 (N_26962,N_20829,N_22026);
nor U26963 (N_26963,N_20602,N_23816);
nor U26964 (N_26964,N_23557,N_20193);
and U26965 (N_26965,N_24262,N_20518);
nor U26966 (N_26966,N_20686,N_22877);
nand U26967 (N_26967,N_24388,N_22918);
xnor U26968 (N_26968,N_21269,N_23848);
xor U26969 (N_26969,N_22606,N_21707);
xnor U26970 (N_26970,N_22838,N_21569);
or U26971 (N_26971,N_23021,N_23907);
and U26972 (N_26972,N_24619,N_22075);
nand U26973 (N_26973,N_24760,N_23867);
xnor U26974 (N_26974,N_21162,N_23472);
nand U26975 (N_26975,N_20280,N_22012);
nand U26976 (N_26976,N_21074,N_23299);
xor U26977 (N_26977,N_24996,N_24637);
nand U26978 (N_26978,N_20021,N_21519);
or U26979 (N_26979,N_21391,N_20803);
nand U26980 (N_26980,N_22059,N_23156);
or U26981 (N_26981,N_24088,N_22645);
or U26982 (N_26982,N_23199,N_24994);
or U26983 (N_26983,N_20006,N_22534);
nor U26984 (N_26984,N_20891,N_24898);
nor U26985 (N_26985,N_24819,N_23574);
xnor U26986 (N_26986,N_21244,N_24352);
xnor U26987 (N_26987,N_21627,N_24100);
nand U26988 (N_26988,N_23043,N_24825);
xnor U26989 (N_26989,N_22525,N_24122);
and U26990 (N_26990,N_22533,N_22295);
nor U26991 (N_26991,N_20105,N_24183);
nand U26992 (N_26992,N_21879,N_20860);
or U26993 (N_26993,N_20384,N_21711);
or U26994 (N_26994,N_21742,N_23426);
nand U26995 (N_26995,N_22884,N_24685);
nor U26996 (N_26996,N_20714,N_21896);
or U26997 (N_26997,N_20571,N_20611);
nor U26998 (N_26998,N_23110,N_20668);
nor U26999 (N_26999,N_24416,N_23064);
nor U27000 (N_27000,N_22505,N_22679);
xnor U27001 (N_27001,N_21233,N_20893);
xnor U27002 (N_27002,N_24120,N_20502);
and U27003 (N_27003,N_24079,N_21972);
and U27004 (N_27004,N_20367,N_23505);
xor U27005 (N_27005,N_22855,N_21853);
nand U27006 (N_27006,N_24355,N_24584);
xor U27007 (N_27007,N_20918,N_23001);
nor U27008 (N_27008,N_20817,N_21771);
nor U27009 (N_27009,N_20447,N_24695);
xnor U27010 (N_27010,N_22688,N_21844);
nor U27011 (N_27011,N_24768,N_23284);
nand U27012 (N_27012,N_21631,N_22280);
xnor U27013 (N_27013,N_24884,N_21768);
or U27014 (N_27014,N_20942,N_22523);
and U27015 (N_27015,N_22541,N_21491);
xor U27016 (N_27016,N_24832,N_23751);
and U27017 (N_27017,N_21821,N_23370);
and U27018 (N_27018,N_22924,N_21932);
and U27019 (N_27019,N_20411,N_22864);
xnor U27020 (N_27020,N_22077,N_20278);
and U27021 (N_27021,N_20297,N_22361);
or U27022 (N_27022,N_23205,N_21927);
nor U27023 (N_27023,N_21785,N_23446);
nand U27024 (N_27024,N_24246,N_24673);
nand U27025 (N_27025,N_20662,N_23354);
nor U27026 (N_27026,N_22814,N_24745);
nor U27027 (N_27027,N_20736,N_20144);
or U27028 (N_27028,N_22640,N_23287);
nor U27029 (N_27029,N_22592,N_22695);
or U27030 (N_27030,N_23160,N_24215);
nand U27031 (N_27031,N_23404,N_22398);
xor U27032 (N_27032,N_20239,N_24623);
nand U27033 (N_27033,N_23502,N_22593);
nand U27034 (N_27034,N_22211,N_23974);
nand U27035 (N_27035,N_24093,N_22888);
nor U27036 (N_27036,N_20160,N_22078);
and U27037 (N_27037,N_20231,N_24690);
nor U27038 (N_27038,N_22334,N_21694);
nor U27039 (N_27039,N_23418,N_22719);
nor U27040 (N_27040,N_24092,N_22968);
xor U27041 (N_27041,N_23876,N_20729);
and U27042 (N_27042,N_20263,N_21985);
nor U27043 (N_27043,N_22546,N_21967);
and U27044 (N_27044,N_22778,N_20806);
or U27045 (N_27045,N_20116,N_23118);
nor U27046 (N_27046,N_21136,N_23723);
and U27047 (N_27047,N_22377,N_21597);
xor U27048 (N_27048,N_21412,N_24258);
and U27049 (N_27049,N_23529,N_20189);
or U27050 (N_27050,N_21912,N_24360);
nor U27051 (N_27051,N_20390,N_23348);
and U27052 (N_27052,N_23362,N_22867);
nand U27053 (N_27053,N_21031,N_20482);
nor U27054 (N_27054,N_21740,N_24828);
and U27055 (N_27055,N_22387,N_24445);
nand U27056 (N_27056,N_22598,N_22151);
or U27057 (N_27057,N_21267,N_22306);
nand U27058 (N_27058,N_24548,N_21761);
and U27059 (N_27059,N_22757,N_23806);
and U27060 (N_27060,N_23132,N_20115);
nand U27061 (N_27061,N_21890,N_24041);
and U27062 (N_27062,N_20661,N_21805);
or U27063 (N_27063,N_24578,N_23760);
nand U27064 (N_27064,N_23888,N_24095);
and U27065 (N_27065,N_24663,N_20972);
nor U27066 (N_27066,N_22826,N_23462);
nand U27067 (N_27067,N_20512,N_24847);
xor U27068 (N_27068,N_21386,N_23282);
nand U27069 (N_27069,N_22477,N_24276);
xnor U27070 (N_27070,N_24721,N_22442);
nor U27071 (N_27071,N_20908,N_21008);
nor U27072 (N_27072,N_20118,N_24765);
and U27073 (N_27073,N_20000,N_21293);
or U27074 (N_27074,N_20272,N_20906);
xor U27075 (N_27075,N_22529,N_23271);
nand U27076 (N_27076,N_22375,N_23066);
nor U27077 (N_27077,N_24123,N_21832);
and U27078 (N_27078,N_22595,N_23605);
nor U27079 (N_27079,N_20778,N_20932);
xnor U27080 (N_27080,N_20938,N_20855);
or U27081 (N_27081,N_23541,N_23601);
or U27082 (N_27082,N_24168,N_23511);
nor U27083 (N_27083,N_21870,N_23471);
xor U27084 (N_27084,N_21029,N_24048);
or U27085 (N_27085,N_24062,N_24984);
nand U27086 (N_27086,N_20435,N_22183);
and U27087 (N_27087,N_22801,N_23768);
and U27088 (N_27088,N_21392,N_21123);
or U27089 (N_27089,N_23238,N_21857);
xnor U27090 (N_27090,N_22950,N_21072);
or U27091 (N_27091,N_23694,N_21151);
or U27092 (N_27092,N_22453,N_24499);
nor U27093 (N_27093,N_23796,N_22080);
xnor U27094 (N_27094,N_20531,N_24517);
or U27095 (N_27095,N_23618,N_22959);
nor U27096 (N_27096,N_22644,N_22675);
or U27097 (N_27097,N_20206,N_20955);
nor U27098 (N_27098,N_24193,N_21646);
nand U27099 (N_27099,N_22336,N_21403);
nand U27100 (N_27100,N_20463,N_21628);
xnor U27101 (N_27101,N_24941,N_20605);
or U27102 (N_27102,N_24116,N_22904);
or U27103 (N_27103,N_23863,N_24675);
nor U27104 (N_27104,N_23420,N_22732);
xnor U27105 (N_27105,N_20727,N_21518);
xnor U27106 (N_27106,N_23688,N_21359);
xor U27107 (N_27107,N_24222,N_20315);
and U27108 (N_27108,N_22339,N_22970);
or U27109 (N_27109,N_24617,N_22802);
or U27110 (N_27110,N_23624,N_22428);
or U27111 (N_27111,N_23654,N_24872);
xor U27112 (N_27112,N_22307,N_21017);
or U27113 (N_27113,N_22294,N_21573);
and U27114 (N_27114,N_22872,N_20859);
and U27115 (N_27115,N_23902,N_22454);
or U27116 (N_27116,N_24464,N_21968);
and U27117 (N_27117,N_22717,N_22328);
or U27118 (N_27118,N_23294,N_24916);
nor U27119 (N_27119,N_22947,N_21435);
nor U27120 (N_27120,N_21015,N_24109);
nor U27121 (N_27121,N_21706,N_22035);
xnor U27122 (N_27122,N_22928,N_20369);
and U27123 (N_27123,N_24606,N_23343);
nor U27124 (N_27124,N_22168,N_21809);
and U27125 (N_27125,N_23377,N_20053);
nor U27126 (N_27126,N_24684,N_24952);
or U27127 (N_27127,N_22648,N_24766);
nor U27128 (N_27128,N_21787,N_22396);
or U27129 (N_27129,N_23222,N_22335);
and U27130 (N_27130,N_24363,N_21173);
or U27131 (N_27131,N_22113,N_22047);
or U27132 (N_27132,N_20958,N_23661);
nor U27133 (N_27133,N_24697,N_22441);
nor U27134 (N_27134,N_22420,N_23374);
xor U27135 (N_27135,N_24854,N_20490);
and U27136 (N_27136,N_20128,N_24458);
nand U27137 (N_27137,N_22753,N_21032);
or U27138 (N_27138,N_22882,N_22599);
and U27139 (N_27139,N_21448,N_21488);
and U27140 (N_27140,N_24964,N_20990);
nand U27141 (N_27141,N_22691,N_20450);
or U27142 (N_27142,N_21134,N_20086);
and U27143 (N_27143,N_20487,N_21923);
nor U27144 (N_27144,N_20054,N_23236);
nand U27145 (N_27145,N_24616,N_22482);
and U27146 (N_27146,N_20620,N_22581);
nand U27147 (N_27147,N_20747,N_22665);
nor U27148 (N_27148,N_21741,N_21283);
or U27149 (N_27149,N_21882,N_22291);
xor U27150 (N_27150,N_20595,N_21629);
nor U27151 (N_27151,N_21410,N_23174);
or U27152 (N_27152,N_23492,N_20726);
nand U27153 (N_27153,N_20638,N_24654);
or U27154 (N_27154,N_20121,N_21777);
or U27155 (N_27155,N_23459,N_24835);
xnor U27156 (N_27156,N_23034,N_23424);
xor U27157 (N_27157,N_22905,N_24107);
nor U27158 (N_27158,N_20804,N_21458);
or U27159 (N_27159,N_20739,N_23685);
nor U27160 (N_27160,N_20003,N_20934);
xnor U27161 (N_27161,N_23747,N_20600);
and U27162 (N_27162,N_22043,N_24749);
xnor U27163 (N_27163,N_23456,N_23604);
and U27164 (N_27164,N_21645,N_24991);
nor U27165 (N_27165,N_24949,N_24980);
and U27166 (N_27166,N_23744,N_20718);
nor U27167 (N_27167,N_24803,N_22596);
and U27168 (N_27168,N_22721,N_20655);
nand U27169 (N_27169,N_21492,N_21424);
and U27170 (N_27170,N_21682,N_23879);
nand U27171 (N_27171,N_23794,N_20245);
and U27172 (N_27172,N_21991,N_24590);
and U27173 (N_27173,N_22495,N_21783);
or U27174 (N_27174,N_22655,N_20303);
nor U27175 (N_27175,N_23596,N_21324);
nor U27176 (N_27176,N_24540,N_21355);
nand U27177 (N_27177,N_23547,N_21417);
nor U27178 (N_27178,N_21515,N_21600);
and U27179 (N_27179,N_22204,N_20285);
nor U27180 (N_27180,N_22614,N_22792);
and U27181 (N_27181,N_20667,N_20480);
xor U27182 (N_27182,N_20989,N_20486);
nand U27183 (N_27183,N_22538,N_24871);
nor U27184 (N_27184,N_24913,N_20730);
and U27185 (N_27185,N_23882,N_23673);
and U27186 (N_27186,N_21956,N_23093);
nor U27187 (N_27187,N_24034,N_22957);
or U27188 (N_27188,N_21078,N_22437);
or U27189 (N_27189,N_21141,N_24398);
xor U27190 (N_27190,N_22029,N_23552);
and U27191 (N_27191,N_22174,N_20797);
or U27192 (N_27192,N_24383,N_24582);
nor U27193 (N_27193,N_20129,N_21228);
nand U27194 (N_27194,N_21144,N_24529);
nor U27195 (N_27195,N_23358,N_21204);
nor U27196 (N_27196,N_21837,N_20775);
xor U27197 (N_27197,N_23234,N_24796);
and U27198 (N_27198,N_20456,N_20559);
xnor U27199 (N_27199,N_24436,N_21854);
or U27200 (N_27200,N_21473,N_24153);
xor U27201 (N_27201,N_21756,N_24956);
and U27202 (N_27202,N_20506,N_20716);
or U27203 (N_27203,N_21182,N_23009);
xnor U27204 (N_27204,N_22129,N_22554);
and U27205 (N_27205,N_22341,N_21545);
nor U27206 (N_27206,N_21514,N_23801);
nor U27207 (N_27207,N_22836,N_23971);
or U27208 (N_27208,N_23324,N_21466);
xnor U27209 (N_27209,N_23727,N_21692);
xnor U27210 (N_27210,N_21981,N_22689);
or U27211 (N_27211,N_23194,N_23625);
and U27212 (N_27212,N_21543,N_23737);
and U27213 (N_27213,N_24583,N_22184);
nor U27214 (N_27214,N_20497,N_23909);
xor U27215 (N_27215,N_23067,N_22006);
nand U27216 (N_27216,N_20043,N_21035);
nand U27217 (N_27217,N_23340,N_22827);
nand U27218 (N_27218,N_24001,N_20684);
nand U27219 (N_27219,N_21637,N_23026);
and U27220 (N_27220,N_23981,N_22516);
nor U27221 (N_27221,N_20774,N_20539);
nor U27222 (N_27222,N_22873,N_24755);
xnor U27223 (N_27223,N_21079,N_20137);
xor U27224 (N_27224,N_20644,N_22188);
nor U27225 (N_27225,N_23246,N_20290);
or U27226 (N_27226,N_22038,N_20166);
nand U27227 (N_27227,N_20033,N_23259);
nand U27228 (N_27228,N_24500,N_24313);
and U27229 (N_27229,N_21180,N_20515);
and U27230 (N_27230,N_23399,N_24438);
or U27231 (N_27231,N_20943,N_21487);
and U27232 (N_27232,N_21076,N_21273);
and U27233 (N_27233,N_23339,N_21007);
and U27234 (N_27234,N_23112,N_22659);
and U27235 (N_27235,N_20832,N_22371);
or U27236 (N_27236,N_20694,N_22603);
or U27237 (N_27237,N_22114,N_24236);
nand U27238 (N_27238,N_21984,N_23167);
xor U27239 (N_27239,N_21174,N_23101);
or U27240 (N_27240,N_24904,N_21418);
nand U27241 (N_27241,N_23989,N_24046);
or U27242 (N_27242,N_23838,N_24185);
and U27243 (N_27243,N_21161,N_21693);
nor U27244 (N_27244,N_20110,N_20810);
xor U27245 (N_27245,N_24028,N_21539);
or U27246 (N_27246,N_23197,N_22289);
xor U27247 (N_27247,N_22019,N_21115);
nor U27248 (N_27248,N_22858,N_22021);
nand U27249 (N_27249,N_23498,N_21500);
nor U27250 (N_27250,N_22760,N_23887);
xnor U27251 (N_27251,N_23951,N_23551);
nand U27252 (N_27252,N_22358,N_20112);
or U27253 (N_27253,N_22587,N_24762);
nor U27254 (N_27254,N_21909,N_20640);
nand U27255 (N_27255,N_20106,N_20831);
and U27256 (N_27256,N_21205,N_23053);
or U27257 (N_27257,N_22249,N_20097);
and U27258 (N_27258,N_20230,N_23656);
xor U27259 (N_27259,N_20219,N_21238);
or U27260 (N_27260,N_20203,N_20868);
and U27261 (N_27261,N_24870,N_20725);
or U27262 (N_27262,N_24943,N_24852);
and U27263 (N_27263,N_20084,N_20478);
nand U27264 (N_27264,N_24125,N_23122);
or U27265 (N_27265,N_22067,N_21253);
or U27266 (N_27266,N_24962,N_23314);
nand U27267 (N_27267,N_21846,N_20119);
and U27268 (N_27268,N_20975,N_20546);
or U27269 (N_27269,N_21483,N_24810);
and U27270 (N_27270,N_21727,N_21610);
xnor U27271 (N_27271,N_23105,N_23048);
and U27272 (N_27272,N_20978,N_22859);
and U27273 (N_27273,N_23148,N_20066);
and U27274 (N_27274,N_23959,N_22216);
or U27275 (N_27275,N_23714,N_20957);
xnor U27276 (N_27276,N_22938,N_23614);
nor U27277 (N_27277,N_20431,N_22200);
and U27278 (N_27278,N_22366,N_21604);
and U27279 (N_27279,N_23023,N_23405);
and U27280 (N_27280,N_23331,N_21725);
or U27281 (N_27281,N_24371,N_23479);
nor U27282 (N_27282,N_22742,N_23764);
and U27283 (N_27283,N_20409,N_23133);
xnor U27284 (N_27284,N_21362,N_22594);
xnor U27285 (N_27285,N_20364,N_24484);
nor U27286 (N_27286,N_20131,N_23483);
xor U27287 (N_27287,N_22986,N_23964);
nand U27288 (N_27288,N_23457,N_21762);
xnor U27289 (N_27289,N_21506,N_21307);
nor U27290 (N_27290,N_22960,N_24263);
or U27291 (N_27291,N_21245,N_20587);
and U27292 (N_27292,N_20783,N_21849);
nand U27293 (N_27293,N_22844,N_24955);
and U27294 (N_27294,N_24269,N_22895);
and U27295 (N_27295,N_23831,N_21936);
xnor U27296 (N_27296,N_24334,N_23635);
xor U27297 (N_27297,N_23912,N_20784);
xnor U27298 (N_27298,N_22083,N_22095);
nor U27299 (N_27299,N_20821,N_20607);
and U27300 (N_27300,N_21964,N_20737);
and U27301 (N_27301,N_20872,N_22510);
nand U27302 (N_27302,N_20150,N_23691);
or U27303 (N_27303,N_24364,N_20544);
nor U27304 (N_27304,N_24565,N_22545);
nor U27305 (N_27305,N_22809,N_21305);
nor U27306 (N_27306,N_21722,N_20145);
nand U27307 (N_27307,N_24407,N_23950);
nor U27308 (N_27308,N_20754,N_21350);
and U27309 (N_27309,N_24069,N_21666);
nor U27310 (N_27310,N_23513,N_24007);
or U27311 (N_27311,N_22707,N_24951);
nor U27312 (N_27312,N_21672,N_23922);
and U27313 (N_27313,N_22716,N_22354);
nor U27314 (N_27314,N_23521,N_21547);
nor U27315 (N_27315,N_21598,N_21721);
nand U27316 (N_27316,N_23185,N_23019);
nor U27317 (N_27317,N_24343,N_20945);
or U27318 (N_27318,N_22046,N_23771);
or U27319 (N_27319,N_20455,N_23415);
xnor U27320 (N_27320,N_22638,N_22098);
xor U27321 (N_27321,N_22051,N_24229);
nor U27322 (N_27322,N_24142,N_20988);
nand U27323 (N_27323,N_20273,N_20257);
nor U27324 (N_27324,N_22360,N_21523);
nand U27325 (N_27325,N_21930,N_21616);
nand U27326 (N_27326,N_20590,N_21700);
or U27327 (N_27327,N_20281,N_21251);
nor U27328 (N_27328,N_20444,N_21829);
or U27329 (N_27329,N_24396,N_23800);
nand U27330 (N_27330,N_24160,N_21368);
xor U27331 (N_27331,N_20612,N_21056);
nor U27332 (N_27332,N_23188,N_20692);
and U27333 (N_27333,N_22004,N_21793);
and U27334 (N_27334,N_22824,N_22934);
nand U27335 (N_27335,N_20025,N_22050);
or U27336 (N_27336,N_22299,N_23962);
or U27337 (N_27337,N_24939,N_20392);
xor U27338 (N_27338,N_23612,N_20646);
nand U27339 (N_27339,N_21997,N_21454);
or U27340 (N_27340,N_22010,N_24566);
or U27341 (N_27341,N_21083,N_24324);
nor U27342 (N_27342,N_20220,N_20074);
nand U27343 (N_27343,N_21688,N_23129);
xor U27344 (N_27344,N_21540,N_23126);
nand U27345 (N_27345,N_20141,N_22146);
xor U27346 (N_27346,N_22110,N_20649);
xor U27347 (N_27347,N_20095,N_22363);
nand U27348 (N_27348,N_23811,N_22403);
or U27349 (N_27349,N_22784,N_21802);
or U27350 (N_27350,N_23263,N_22842);
nand U27351 (N_27351,N_23490,N_21311);
and U27352 (N_27352,N_23980,N_24216);
or U27353 (N_27353,N_20654,N_22150);
and U27354 (N_27354,N_20437,N_23334);
or U27355 (N_27355,N_24300,N_24769);
nor U27356 (N_27356,N_22762,N_22916);
nand U27357 (N_27357,N_21441,N_21709);
and U27358 (N_27358,N_22194,N_22176);
nor U27359 (N_27359,N_22574,N_24056);
xnor U27360 (N_27360,N_24150,N_22074);
nand U27361 (N_27361,N_21951,N_21001);
nand U27362 (N_27362,N_24742,N_20484);
or U27363 (N_27363,N_20577,N_23114);
nor U27364 (N_27364,N_24761,N_21213);
or U27365 (N_27365,N_24118,N_21342);
nor U27366 (N_27366,N_24921,N_22927);
xnor U27367 (N_27367,N_24008,N_21532);
xnor U27368 (N_27368,N_20776,N_21484);
nand U27369 (N_27369,N_24777,N_23566);
nand U27370 (N_27370,N_22111,N_20909);
or U27371 (N_27371,N_23706,N_22513);
or U27372 (N_27372,N_23027,N_24652);
and U27373 (N_27373,N_24521,N_22658);
and U27374 (N_27374,N_20326,N_22579);
or U27375 (N_27375,N_23228,N_24823);
xor U27376 (N_27376,N_20301,N_21830);
nand U27377 (N_27377,N_22631,N_23142);
and U27378 (N_27378,N_21873,N_21155);
nor U27379 (N_27379,N_21842,N_22776);
nor U27380 (N_27380,N_20901,N_23091);
nand U27381 (N_27381,N_24017,N_21810);
nor U27382 (N_27382,N_24050,N_20430);
xnor U27383 (N_27383,N_22736,N_23983);
xnor U27384 (N_27384,N_20676,N_22000);
nor U27385 (N_27385,N_24461,N_23766);
nand U27386 (N_27386,N_21557,N_22962);
nand U27387 (N_27387,N_20586,N_20291);
or U27388 (N_27388,N_21883,N_24827);
nor U27389 (N_27389,N_22668,N_21313);
or U27390 (N_27390,N_23038,N_21856);
and U27391 (N_27391,N_21588,N_20911);
xnor U27392 (N_27392,N_24090,N_24948);
nor U27393 (N_27393,N_20617,N_23885);
xnor U27394 (N_27394,N_22117,N_21066);
xnor U27395 (N_27395,N_21187,N_23297);
nand U27396 (N_27396,N_23108,N_21099);
nand U27397 (N_27397,N_22028,N_22422);
xnor U27398 (N_27398,N_21110,N_24934);
and U27399 (N_27399,N_22384,N_24798);
or U27400 (N_27400,N_24256,N_20690);
or U27401 (N_27401,N_21456,N_23310);
and U27402 (N_27402,N_22034,N_22556);
or U27403 (N_27403,N_21142,N_21966);
or U27404 (N_27404,N_21319,N_24400);
nor U27405 (N_27405,N_20002,N_22364);
xnor U27406 (N_27406,N_20042,N_22142);
or U27407 (N_27407,N_21409,N_23819);
and U27408 (N_27408,N_22854,N_21113);
and U27409 (N_27409,N_21493,N_20469);
xor U27410 (N_27410,N_22789,N_23445);
nor U27411 (N_27411,N_21841,N_21962);
or U27412 (N_27412,N_24838,N_22300);
or U27413 (N_27413,N_22292,N_22410);
nand U27414 (N_27414,N_24576,N_24204);
or U27415 (N_27415,N_21176,N_22766);
or U27416 (N_27416,N_23813,N_24700);
or U27417 (N_27417,N_23225,N_22733);
nand U27418 (N_27418,N_22794,N_21249);
xor U27419 (N_27419,N_20704,N_24862);
or U27420 (N_27420,N_23941,N_20146);
and U27421 (N_27421,N_21133,N_24611);
xnor U27422 (N_27422,N_23731,N_24694);
xor U27423 (N_27423,N_24024,N_20383);
or U27424 (N_27424,N_23041,N_22623);
xor U27425 (N_27425,N_24789,N_21020);
nor U27426 (N_27426,N_22096,N_24283);
xnor U27427 (N_27427,N_23495,N_22426);
xor U27428 (N_27428,N_21864,N_20175);
nor U27429 (N_27429,N_24476,N_24412);
nor U27430 (N_27430,N_21556,N_22666);
nor U27431 (N_27431,N_21512,N_22543);
nand U27432 (N_27432,N_24105,N_21795);
nand U27433 (N_27433,N_21026,N_20937);
or U27434 (N_27434,N_20688,N_24998);
or U27435 (N_27435,N_20802,N_21053);
xnor U27436 (N_27436,N_21190,N_20697);
xor U27437 (N_27437,N_21160,N_23854);
and U27438 (N_27438,N_21374,N_24058);
nor U27439 (N_27439,N_22747,N_22101);
nand U27440 (N_27440,N_23144,N_20148);
nand U27441 (N_27441,N_22158,N_24052);
nor U27442 (N_27442,N_24595,N_21295);
and U27443 (N_27443,N_24776,N_21106);
nand U27444 (N_27444,N_21568,N_24550);
or U27445 (N_27445,N_21156,N_22897);
or U27446 (N_27446,N_23302,N_20015);
and U27447 (N_27447,N_20176,N_20927);
nor U27448 (N_27448,N_22001,N_24138);
or U27449 (N_27449,N_21541,N_23224);
xnor U27450 (N_27450,N_22782,N_23074);
and U27451 (N_27451,N_24139,N_22997);
nor U27452 (N_27452,N_23213,N_24156);
and U27453 (N_27453,N_20865,N_22172);
or U27454 (N_27454,N_22238,N_21505);
xor U27455 (N_27455,N_23943,N_22621);
and U27456 (N_27456,N_22969,N_21394);
xor U27457 (N_27457,N_24610,N_24908);
xor U27458 (N_27458,N_20618,N_21420);
nor U27459 (N_27459,N_20557,N_20637);
nand U27460 (N_27460,N_23743,N_23772);
and U27461 (N_27461,N_21924,N_24195);
nand U27462 (N_27462,N_20331,N_21922);
and U27463 (N_27463,N_21958,N_23787);
nor U27464 (N_27464,N_20082,N_23494);
xnor U27465 (N_27465,N_24664,N_22178);
and U27466 (N_27466,N_23804,N_21346);
and U27467 (N_27467,N_21105,N_23561);
and U27468 (N_27468,N_20869,N_24121);
nor U27469 (N_27469,N_20494,N_21088);
nand U27470 (N_27470,N_24580,N_22863);
and U27471 (N_27471,N_20104,N_21261);
xor U27472 (N_27472,N_23135,N_20701);
or U27473 (N_27473,N_21452,N_22808);
nand U27474 (N_27474,N_22617,N_23708);
or U27475 (N_27475,N_23797,N_20510);
nor U27476 (N_27476,N_23022,N_22830);
and U27477 (N_27477,N_21416,N_22130);
or U27478 (N_27478,N_21516,N_20973);
or U27479 (N_27479,N_21332,N_21733);
nor U27480 (N_27480,N_24886,N_23675);
nor U27481 (N_27481,N_23403,N_20743);
or U27482 (N_27482,N_21376,N_20346);
or U27483 (N_27483,N_21668,N_23180);
xor U27484 (N_27484,N_24714,N_20139);
and U27485 (N_27485,N_23373,N_21382);
and U27486 (N_27486,N_22995,N_23016);
and U27487 (N_27487,N_21184,N_24233);
and U27488 (N_27488,N_22418,N_20051);
xnor U27489 (N_27489,N_21430,N_22457);
nor U27490 (N_27490,N_21738,N_20665);
xor U27491 (N_27491,N_24603,N_23159);
and U27492 (N_27492,N_21328,N_22416);
xnor U27493 (N_27493,N_24428,N_24990);
nand U27494 (N_27494,N_23241,N_21561);
nand U27495 (N_27495,N_22773,N_23380);
xor U27496 (N_27496,N_21875,N_23877);
or U27497 (N_27497,N_24528,N_24596);
xnor U27498 (N_27498,N_24713,N_21147);
xnor U27499 (N_27499,N_24025,N_20363);
or U27500 (N_27500,N_23863,N_22497);
nand U27501 (N_27501,N_21266,N_22759);
nor U27502 (N_27502,N_22906,N_23060);
xor U27503 (N_27503,N_21523,N_22563);
or U27504 (N_27504,N_24352,N_24929);
nor U27505 (N_27505,N_20878,N_20451);
nand U27506 (N_27506,N_24761,N_20221);
or U27507 (N_27507,N_21874,N_24745);
nor U27508 (N_27508,N_24433,N_23465);
nor U27509 (N_27509,N_23467,N_24432);
nand U27510 (N_27510,N_24205,N_22706);
nor U27511 (N_27511,N_20152,N_21272);
xor U27512 (N_27512,N_23332,N_24409);
nand U27513 (N_27513,N_20572,N_24077);
and U27514 (N_27514,N_20983,N_22808);
xor U27515 (N_27515,N_20643,N_23116);
nand U27516 (N_27516,N_23495,N_21314);
xor U27517 (N_27517,N_24605,N_23193);
nor U27518 (N_27518,N_23040,N_24247);
and U27519 (N_27519,N_23495,N_22099);
and U27520 (N_27520,N_22936,N_24164);
nand U27521 (N_27521,N_20867,N_21744);
nand U27522 (N_27522,N_20584,N_21005);
xnor U27523 (N_27523,N_21763,N_24687);
nand U27524 (N_27524,N_24296,N_21700);
or U27525 (N_27525,N_24969,N_23450);
and U27526 (N_27526,N_22990,N_22879);
or U27527 (N_27527,N_21643,N_24302);
and U27528 (N_27528,N_23475,N_22754);
xor U27529 (N_27529,N_22960,N_23246);
nor U27530 (N_27530,N_21420,N_20332);
and U27531 (N_27531,N_22588,N_24434);
or U27532 (N_27532,N_22757,N_23557);
nand U27533 (N_27533,N_20920,N_20062);
or U27534 (N_27534,N_20794,N_23793);
nor U27535 (N_27535,N_21339,N_24996);
or U27536 (N_27536,N_23744,N_21066);
nor U27537 (N_27537,N_22007,N_23759);
and U27538 (N_27538,N_20621,N_23366);
nand U27539 (N_27539,N_21999,N_21667);
nand U27540 (N_27540,N_23467,N_20843);
and U27541 (N_27541,N_24813,N_24807);
xor U27542 (N_27542,N_24227,N_24546);
and U27543 (N_27543,N_23481,N_22330);
and U27544 (N_27544,N_24824,N_24062);
and U27545 (N_27545,N_21580,N_22876);
nor U27546 (N_27546,N_23511,N_21770);
and U27547 (N_27547,N_21072,N_20227);
and U27548 (N_27548,N_23305,N_20884);
nand U27549 (N_27549,N_23472,N_20780);
xnor U27550 (N_27550,N_22943,N_23569);
xor U27551 (N_27551,N_21526,N_24794);
or U27552 (N_27552,N_20092,N_21230);
nor U27553 (N_27553,N_21068,N_20923);
nor U27554 (N_27554,N_24865,N_22199);
or U27555 (N_27555,N_23875,N_20706);
and U27556 (N_27556,N_20712,N_23890);
xnor U27557 (N_27557,N_23998,N_21456);
or U27558 (N_27558,N_24954,N_21404);
or U27559 (N_27559,N_22959,N_23419);
xor U27560 (N_27560,N_22550,N_23441);
xnor U27561 (N_27561,N_22833,N_20945);
nor U27562 (N_27562,N_23731,N_20035);
xor U27563 (N_27563,N_21999,N_21097);
and U27564 (N_27564,N_22175,N_24872);
nor U27565 (N_27565,N_20399,N_22701);
and U27566 (N_27566,N_22820,N_20557);
nor U27567 (N_27567,N_22261,N_24301);
nand U27568 (N_27568,N_23713,N_23558);
nor U27569 (N_27569,N_20929,N_23302);
or U27570 (N_27570,N_23846,N_20569);
and U27571 (N_27571,N_21012,N_24073);
xor U27572 (N_27572,N_24604,N_22800);
nand U27573 (N_27573,N_24754,N_20116);
xnor U27574 (N_27574,N_24474,N_21928);
xnor U27575 (N_27575,N_23468,N_24600);
or U27576 (N_27576,N_23715,N_24554);
nand U27577 (N_27577,N_21575,N_20818);
or U27578 (N_27578,N_24695,N_20700);
nor U27579 (N_27579,N_21646,N_24322);
or U27580 (N_27580,N_24881,N_22668);
nor U27581 (N_27581,N_20806,N_24360);
nor U27582 (N_27582,N_24191,N_20214);
nand U27583 (N_27583,N_21675,N_24648);
nand U27584 (N_27584,N_23420,N_22787);
nand U27585 (N_27585,N_20463,N_20247);
or U27586 (N_27586,N_23625,N_21233);
nor U27587 (N_27587,N_22533,N_21495);
and U27588 (N_27588,N_24048,N_22819);
and U27589 (N_27589,N_23753,N_21083);
xor U27590 (N_27590,N_23178,N_21070);
or U27591 (N_27591,N_21181,N_20605);
or U27592 (N_27592,N_20283,N_22385);
xnor U27593 (N_27593,N_20749,N_20700);
nand U27594 (N_27594,N_22415,N_24790);
or U27595 (N_27595,N_24827,N_23135);
nand U27596 (N_27596,N_22468,N_22352);
nor U27597 (N_27597,N_22144,N_24952);
or U27598 (N_27598,N_24698,N_23088);
nand U27599 (N_27599,N_22164,N_20598);
and U27600 (N_27600,N_23267,N_23144);
nand U27601 (N_27601,N_24468,N_20635);
nand U27602 (N_27602,N_23446,N_23310);
xnor U27603 (N_27603,N_20960,N_21235);
nor U27604 (N_27604,N_22218,N_20793);
or U27605 (N_27605,N_20004,N_23730);
or U27606 (N_27606,N_22553,N_23643);
nand U27607 (N_27607,N_23441,N_23242);
xor U27608 (N_27608,N_22505,N_20494);
xnor U27609 (N_27609,N_23569,N_22092);
nand U27610 (N_27610,N_22790,N_24529);
nor U27611 (N_27611,N_23070,N_23175);
xor U27612 (N_27612,N_23254,N_21082);
or U27613 (N_27613,N_23653,N_20465);
and U27614 (N_27614,N_20623,N_21647);
xnor U27615 (N_27615,N_21944,N_22338);
and U27616 (N_27616,N_24673,N_24282);
xor U27617 (N_27617,N_24157,N_21703);
xor U27618 (N_27618,N_24297,N_24367);
and U27619 (N_27619,N_24182,N_21713);
and U27620 (N_27620,N_24975,N_20948);
xor U27621 (N_27621,N_21910,N_20254);
nand U27622 (N_27622,N_21715,N_24969);
or U27623 (N_27623,N_21064,N_24195);
nor U27624 (N_27624,N_24621,N_20411);
or U27625 (N_27625,N_23248,N_22563);
nor U27626 (N_27626,N_20709,N_22042);
nand U27627 (N_27627,N_21787,N_22536);
nand U27628 (N_27628,N_20399,N_21823);
xor U27629 (N_27629,N_24635,N_22973);
xnor U27630 (N_27630,N_23481,N_21546);
nor U27631 (N_27631,N_21464,N_23237);
xnor U27632 (N_27632,N_20598,N_24172);
and U27633 (N_27633,N_24250,N_24133);
nand U27634 (N_27634,N_21752,N_21574);
or U27635 (N_27635,N_21590,N_22166);
xnor U27636 (N_27636,N_20829,N_24301);
xor U27637 (N_27637,N_23034,N_20866);
or U27638 (N_27638,N_20782,N_24038);
and U27639 (N_27639,N_21018,N_22764);
nand U27640 (N_27640,N_22080,N_23349);
nor U27641 (N_27641,N_23887,N_22934);
nand U27642 (N_27642,N_23143,N_21854);
nor U27643 (N_27643,N_24465,N_21074);
and U27644 (N_27644,N_24060,N_20785);
nor U27645 (N_27645,N_20923,N_21146);
nand U27646 (N_27646,N_21994,N_23112);
nor U27647 (N_27647,N_22915,N_22599);
nand U27648 (N_27648,N_24162,N_24630);
and U27649 (N_27649,N_24774,N_20024);
or U27650 (N_27650,N_23410,N_24989);
or U27651 (N_27651,N_24132,N_23560);
and U27652 (N_27652,N_21744,N_20174);
or U27653 (N_27653,N_20003,N_20243);
nor U27654 (N_27654,N_20852,N_24723);
and U27655 (N_27655,N_23546,N_22831);
nand U27656 (N_27656,N_22453,N_23211);
nand U27657 (N_27657,N_21010,N_23258);
or U27658 (N_27658,N_20781,N_22991);
xnor U27659 (N_27659,N_21028,N_22185);
nand U27660 (N_27660,N_23024,N_20157);
and U27661 (N_27661,N_22345,N_23350);
nor U27662 (N_27662,N_22959,N_22349);
xor U27663 (N_27663,N_23629,N_24534);
nand U27664 (N_27664,N_20857,N_21519);
or U27665 (N_27665,N_23573,N_24815);
nand U27666 (N_27666,N_23195,N_24384);
nand U27667 (N_27667,N_20236,N_23402);
xnor U27668 (N_27668,N_21225,N_24300);
and U27669 (N_27669,N_24740,N_23723);
nor U27670 (N_27670,N_22533,N_23187);
or U27671 (N_27671,N_22942,N_22736);
and U27672 (N_27672,N_24112,N_21789);
or U27673 (N_27673,N_21354,N_23548);
nand U27674 (N_27674,N_24893,N_24697);
and U27675 (N_27675,N_20484,N_22881);
nand U27676 (N_27676,N_24712,N_24801);
or U27677 (N_27677,N_20690,N_23182);
and U27678 (N_27678,N_24859,N_20979);
nand U27679 (N_27679,N_23860,N_20002);
and U27680 (N_27680,N_24785,N_21745);
nor U27681 (N_27681,N_23784,N_24147);
xnor U27682 (N_27682,N_21760,N_23595);
nor U27683 (N_27683,N_23775,N_20043);
and U27684 (N_27684,N_23442,N_24017);
xor U27685 (N_27685,N_20326,N_24046);
nand U27686 (N_27686,N_22348,N_23881);
nand U27687 (N_27687,N_21174,N_21343);
nand U27688 (N_27688,N_24019,N_21347);
or U27689 (N_27689,N_22820,N_21600);
and U27690 (N_27690,N_20196,N_23031);
or U27691 (N_27691,N_24552,N_24436);
nand U27692 (N_27692,N_23572,N_22410);
or U27693 (N_27693,N_22650,N_21805);
nor U27694 (N_27694,N_23834,N_21247);
and U27695 (N_27695,N_23620,N_21017);
or U27696 (N_27696,N_24455,N_20151);
nand U27697 (N_27697,N_21981,N_21759);
and U27698 (N_27698,N_21752,N_20049);
nand U27699 (N_27699,N_22653,N_22750);
nand U27700 (N_27700,N_22028,N_21352);
or U27701 (N_27701,N_23118,N_22575);
or U27702 (N_27702,N_21444,N_22240);
nand U27703 (N_27703,N_24079,N_21021);
nor U27704 (N_27704,N_23131,N_23475);
nor U27705 (N_27705,N_22315,N_24829);
and U27706 (N_27706,N_21732,N_20009);
and U27707 (N_27707,N_23050,N_24974);
nand U27708 (N_27708,N_20390,N_22087);
xnor U27709 (N_27709,N_23523,N_24114);
xnor U27710 (N_27710,N_24543,N_23224);
nor U27711 (N_27711,N_22142,N_24000);
xor U27712 (N_27712,N_22964,N_20273);
nand U27713 (N_27713,N_21410,N_24075);
xor U27714 (N_27714,N_23670,N_20995);
nor U27715 (N_27715,N_24958,N_21672);
or U27716 (N_27716,N_23722,N_21137);
nor U27717 (N_27717,N_21880,N_20618);
and U27718 (N_27718,N_21106,N_21505);
nand U27719 (N_27719,N_24575,N_22859);
nand U27720 (N_27720,N_21861,N_21034);
xor U27721 (N_27721,N_24225,N_24818);
xor U27722 (N_27722,N_24052,N_22776);
or U27723 (N_27723,N_24849,N_20458);
nand U27724 (N_27724,N_21047,N_20624);
nor U27725 (N_27725,N_24074,N_23622);
or U27726 (N_27726,N_20266,N_24308);
xnor U27727 (N_27727,N_24840,N_20964);
xor U27728 (N_27728,N_23625,N_23069);
nor U27729 (N_27729,N_20799,N_21803);
nand U27730 (N_27730,N_20503,N_22265);
nand U27731 (N_27731,N_23808,N_21489);
xnor U27732 (N_27732,N_24253,N_20280);
and U27733 (N_27733,N_21874,N_20487);
nor U27734 (N_27734,N_20023,N_21081);
nand U27735 (N_27735,N_23873,N_22516);
or U27736 (N_27736,N_21419,N_21033);
or U27737 (N_27737,N_21602,N_21141);
or U27738 (N_27738,N_20410,N_21227);
or U27739 (N_27739,N_22036,N_21298);
nor U27740 (N_27740,N_22089,N_24014);
and U27741 (N_27741,N_21522,N_21529);
or U27742 (N_27742,N_22181,N_23990);
nand U27743 (N_27743,N_24768,N_24546);
xor U27744 (N_27744,N_23348,N_21997);
and U27745 (N_27745,N_20383,N_20688);
nor U27746 (N_27746,N_21222,N_24986);
and U27747 (N_27747,N_20553,N_24925);
nor U27748 (N_27748,N_23012,N_21912);
or U27749 (N_27749,N_21699,N_23202);
or U27750 (N_27750,N_22555,N_23688);
xor U27751 (N_27751,N_24321,N_23940);
nor U27752 (N_27752,N_24305,N_24517);
nand U27753 (N_27753,N_22325,N_21618);
nand U27754 (N_27754,N_24416,N_21392);
nor U27755 (N_27755,N_22205,N_20271);
or U27756 (N_27756,N_22193,N_23108);
nand U27757 (N_27757,N_22549,N_21964);
and U27758 (N_27758,N_20409,N_22573);
and U27759 (N_27759,N_24096,N_23752);
and U27760 (N_27760,N_21216,N_21964);
nand U27761 (N_27761,N_24110,N_21655);
nor U27762 (N_27762,N_24150,N_23506);
and U27763 (N_27763,N_24756,N_21882);
and U27764 (N_27764,N_23147,N_20783);
nand U27765 (N_27765,N_21750,N_21665);
and U27766 (N_27766,N_21035,N_20577);
or U27767 (N_27767,N_22077,N_22893);
and U27768 (N_27768,N_20480,N_24459);
nand U27769 (N_27769,N_22440,N_24311);
or U27770 (N_27770,N_24211,N_21455);
xnor U27771 (N_27771,N_24400,N_20332);
nor U27772 (N_27772,N_21905,N_22894);
nand U27773 (N_27773,N_23884,N_21868);
and U27774 (N_27774,N_20554,N_21579);
or U27775 (N_27775,N_20900,N_24545);
xor U27776 (N_27776,N_20902,N_24207);
or U27777 (N_27777,N_20509,N_22684);
or U27778 (N_27778,N_20554,N_24054);
and U27779 (N_27779,N_22472,N_23429);
or U27780 (N_27780,N_21870,N_23356);
or U27781 (N_27781,N_24966,N_21130);
nor U27782 (N_27782,N_20553,N_24427);
xnor U27783 (N_27783,N_21923,N_22241);
xnor U27784 (N_27784,N_20967,N_21506);
and U27785 (N_27785,N_21239,N_21513);
nand U27786 (N_27786,N_22245,N_23324);
and U27787 (N_27787,N_21532,N_24191);
xor U27788 (N_27788,N_20374,N_23714);
or U27789 (N_27789,N_20366,N_21997);
and U27790 (N_27790,N_20020,N_21984);
nor U27791 (N_27791,N_21506,N_20141);
or U27792 (N_27792,N_22545,N_23248);
xor U27793 (N_27793,N_22052,N_22441);
nor U27794 (N_27794,N_20410,N_20581);
nor U27795 (N_27795,N_21418,N_23809);
or U27796 (N_27796,N_23290,N_21760);
nor U27797 (N_27797,N_23280,N_24810);
nor U27798 (N_27798,N_22413,N_23586);
nor U27799 (N_27799,N_22488,N_24120);
or U27800 (N_27800,N_23481,N_23013);
and U27801 (N_27801,N_24465,N_21514);
or U27802 (N_27802,N_22784,N_21794);
xor U27803 (N_27803,N_23543,N_23926);
or U27804 (N_27804,N_22882,N_21226);
and U27805 (N_27805,N_21584,N_20665);
and U27806 (N_27806,N_20157,N_21811);
nand U27807 (N_27807,N_24467,N_24357);
nor U27808 (N_27808,N_21871,N_24226);
and U27809 (N_27809,N_22547,N_21076);
or U27810 (N_27810,N_22164,N_24766);
nor U27811 (N_27811,N_22549,N_23545);
or U27812 (N_27812,N_21256,N_22287);
or U27813 (N_27813,N_24260,N_23584);
or U27814 (N_27814,N_21510,N_20958);
or U27815 (N_27815,N_20060,N_24139);
xnor U27816 (N_27816,N_20315,N_23121);
or U27817 (N_27817,N_22332,N_22268);
xnor U27818 (N_27818,N_24980,N_22418);
nand U27819 (N_27819,N_23529,N_23847);
xor U27820 (N_27820,N_24902,N_24549);
and U27821 (N_27821,N_22446,N_22029);
nor U27822 (N_27822,N_21702,N_23227);
or U27823 (N_27823,N_24622,N_24304);
nand U27824 (N_27824,N_23727,N_24793);
xnor U27825 (N_27825,N_22346,N_23980);
nor U27826 (N_27826,N_22518,N_20668);
nor U27827 (N_27827,N_24709,N_22132);
nand U27828 (N_27828,N_23163,N_24625);
nand U27829 (N_27829,N_20840,N_23930);
xnor U27830 (N_27830,N_22490,N_20855);
nand U27831 (N_27831,N_20470,N_24379);
xnor U27832 (N_27832,N_24783,N_23115);
nand U27833 (N_27833,N_23584,N_24170);
or U27834 (N_27834,N_22596,N_24436);
or U27835 (N_27835,N_22494,N_23547);
nor U27836 (N_27836,N_22189,N_21948);
xor U27837 (N_27837,N_24059,N_23481);
nor U27838 (N_27838,N_24288,N_20844);
and U27839 (N_27839,N_21170,N_21380);
xnor U27840 (N_27840,N_24114,N_24203);
xor U27841 (N_27841,N_21536,N_24369);
or U27842 (N_27842,N_23033,N_23659);
or U27843 (N_27843,N_21233,N_22557);
nand U27844 (N_27844,N_22287,N_21100);
and U27845 (N_27845,N_20406,N_24075);
nor U27846 (N_27846,N_21827,N_24738);
xor U27847 (N_27847,N_23706,N_21547);
nand U27848 (N_27848,N_21949,N_20735);
nor U27849 (N_27849,N_21092,N_20518);
nor U27850 (N_27850,N_24934,N_24013);
xnor U27851 (N_27851,N_23658,N_23243);
nor U27852 (N_27852,N_24179,N_24831);
nor U27853 (N_27853,N_24176,N_23699);
nand U27854 (N_27854,N_20858,N_22514);
nor U27855 (N_27855,N_20422,N_20559);
nor U27856 (N_27856,N_24443,N_22838);
and U27857 (N_27857,N_22274,N_21843);
nand U27858 (N_27858,N_23220,N_21935);
nor U27859 (N_27859,N_20462,N_22575);
nor U27860 (N_27860,N_21767,N_23335);
or U27861 (N_27861,N_21594,N_22424);
xnor U27862 (N_27862,N_24464,N_24374);
nor U27863 (N_27863,N_24347,N_24430);
or U27864 (N_27864,N_22328,N_24539);
xnor U27865 (N_27865,N_23096,N_23379);
xnor U27866 (N_27866,N_21416,N_24667);
nand U27867 (N_27867,N_20176,N_20331);
nand U27868 (N_27868,N_24283,N_22981);
nand U27869 (N_27869,N_23255,N_24615);
nand U27870 (N_27870,N_23369,N_20617);
or U27871 (N_27871,N_20665,N_24464);
or U27872 (N_27872,N_24696,N_24617);
nor U27873 (N_27873,N_23183,N_23577);
and U27874 (N_27874,N_24696,N_20315);
xor U27875 (N_27875,N_24835,N_23835);
xnor U27876 (N_27876,N_23421,N_21869);
nor U27877 (N_27877,N_22411,N_21125);
nor U27878 (N_27878,N_24054,N_23461);
nand U27879 (N_27879,N_21747,N_20820);
xor U27880 (N_27880,N_24357,N_21989);
nor U27881 (N_27881,N_23529,N_22949);
and U27882 (N_27882,N_24272,N_21686);
nand U27883 (N_27883,N_24241,N_23470);
xnor U27884 (N_27884,N_24575,N_24549);
xnor U27885 (N_27885,N_21941,N_22003);
and U27886 (N_27886,N_21142,N_22350);
and U27887 (N_27887,N_21820,N_21242);
and U27888 (N_27888,N_21225,N_23737);
and U27889 (N_27889,N_23296,N_22550);
or U27890 (N_27890,N_22335,N_23589);
and U27891 (N_27891,N_22950,N_23757);
or U27892 (N_27892,N_23491,N_20660);
and U27893 (N_27893,N_24850,N_20550);
xor U27894 (N_27894,N_23462,N_20921);
and U27895 (N_27895,N_24220,N_20631);
nand U27896 (N_27896,N_24947,N_22633);
xor U27897 (N_27897,N_20682,N_24797);
and U27898 (N_27898,N_24547,N_21342);
or U27899 (N_27899,N_24031,N_20709);
xnor U27900 (N_27900,N_24589,N_21149);
nand U27901 (N_27901,N_24785,N_20258);
nand U27902 (N_27902,N_24990,N_23391);
or U27903 (N_27903,N_20362,N_22180);
or U27904 (N_27904,N_23796,N_20498);
nand U27905 (N_27905,N_21696,N_20352);
and U27906 (N_27906,N_24168,N_21155);
nor U27907 (N_27907,N_24791,N_23836);
or U27908 (N_27908,N_21840,N_23117);
xnor U27909 (N_27909,N_22364,N_22326);
or U27910 (N_27910,N_20363,N_23238);
xnor U27911 (N_27911,N_20462,N_23073);
xor U27912 (N_27912,N_20913,N_22219);
or U27913 (N_27913,N_22055,N_24645);
nand U27914 (N_27914,N_22678,N_20526);
and U27915 (N_27915,N_24944,N_22078);
and U27916 (N_27916,N_24444,N_21990);
nor U27917 (N_27917,N_23595,N_23680);
xnor U27918 (N_27918,N_21814,N_20729);
or U27919 (N_27919,N_20751,N_20983);
and U27920 (N_27920,N_23020,N_24509);
and U27921 (N_27921,N_22877,N_21278);
and U27922 (N_27922,N_22217,N_23085);
nor U27923 (N_27923,N_24918,N_22370);
nor U27924 (N_27924,N_21401,N_22417);
and U27925 (N_27925,N_20402,N_23423);
and U27926 (N_27926,N_23515,N_23424);
nand U27927 (N_27927,N_22784,N_24879);
nor U27928 (N_27928,N_20320,N_21073);
or U27929 (N_27929,N_24018,N_22364);
xnor U27930 (N_27930,N_20521,N_24718);
and U27931 (N_27931,N_21102,N_21294);
and U27932 (N_27932,N_20273,N_22000);
and U27933 (N_27933,N_23442,N_24042);
nand U27934 (N_27934,N_24389,N_24899);
xnor U27935 (N_27935,N_20597,N_22911);
and U27936 (N_27936,N_22825,N_22591);
nand U27937 (N_27937,N_23744,N_21646);
nor U27938 (N_27938,N_22990,N_24947);
nand U27939 (N_27939,N_23520,N_20876);
nor U27940 (N_27940,N_23144,N_20178);
nor U27941 (N_27941,N_22735,N_24965);
or U27942 (N_27942,N_20870,N_20540);
xor U27943 (N_27943,N_23003,N_24770);
xnor U27944 (N_27944,N_22853,N_22899);
nor U27945 (N_27945,N_22621,N_22618);
and U27946 (N_27946,N_22628,N_23450);
xor U27947 (N_27947,N_24041,N_21393);
or U27948 (N_27948,N_24647,N_24928);
and U27949 (N_27949,N_22516,N_22938);
nand U27950 (N_27950,N_20966,N_20636);
nor U27951 (N_27951,N_22140,N_22100);
xor U27952 (N_27952,N_23006,N_21914);
xor U27953 (N_27953,N_24367,N_22587);
and U27954 (N_27954,N_23266,N_20952);
nand U27955 (N_27955,N_22386,N_20385);
xor U27956 (N_27956,N_24032,N_23804);
and U27957 (N_27957,N_20432,N_22747);
nor U27958 (N_27958,N_23356,N_22775);
nand U27959 (N_27959,N_22032,N_22212);
and U27960 (N_27960,N_24079,N_24865);
nor U27961 (N_27961,N_24785,N_24121);
or U27962 (N_27962,N_20996,N_20544);
or U27963 (N_27963,N_24003,N_24714);
nand U27964 (N_27964,N_22727,N_22896);
nand U27965 (N_27965,N_24573,N_23380);
nor U27966 (N_27966,N_24585,N_23471);
xor U27967 (N_27967,N_22134,N_20193);
and U27968 (N_27968,N_23494,N_20916);
or U27969 (N_27969,N_22291,N_22156);
xnor U27970 (N_27970,N_22696,N_23285);
or U27971 (N_27971,N_24439,N_24082);
xor U27972 (N_27972,N_22221,N_22133);
or U27973 (N_27973,N_21262,N_22839);
nor U27974 (N_27974,N_24554,N_21298);
nand U27975 (N_27975,N_21247,N_21510);
nand U27976 (N_27976,N_24456,N_22163);
xor U27977 (N_27977,N_22416,N_23146);
nand U27978 (N_27978,N_21969,N_22941);
or U27979 (N_27979,N_21188,N_22190);
nand U27980 (N_27980,N_24533,N_23981);
xor U27981 (N_27981,N_23174,N_22004);
or U27982 (N_27982,N_22304,N_24285);
or U27983 (N_27983,N_23539,N_24036);
nor U27984 (N_27984,N_22736,N_24141);
or U27985 (N_27985,N_20196,N_24739);
nor U27986 (N_27986,N_24931,N_20420);
xor U27987 (N_27987,N_24589,N_21195);
or U27988 (N_27988,N_20186,N_20127);
nand U27989 (N_27989,N_23289,N_21825);
nand U27990 (N_27990,N_22364,N_22152);
or U27991 (N_27991,N_24955,N_21270);
or U27992 (N_27992,N_22604,N_23417);
and U27993 (N_27993,N_20234,N_20389);
xor U27994 (N_27994,N_23523,N_23861);
nor U27995 (N_27995,N_24206,N_21844);
nand U27996 (N_27996,N_24467,N_21356);
or U27997 (N_27997,N_23873,N_20396);
nand U27998 (N_27998,N_23272,N_24168);
and U27999 (N_27999,N_23489,N_24148);
or U28000 (N_28000,N_22738,N_20947);
and U28001 (N_28001,N_21820,N_20090);
or U28002 (N_28002,N_23917,N_21120);
or U28003 (N_28003,N_24943,N_22126);
xnor U28004 (N_28004,N_23335,N_21248);
xnor U28005 (N_28005,N_20511,N_23705);
nand U28006 (N_28006,N_24305,N_24725);
xor U28007 (N_28007,N_21960,N_21022);
and U28008 (N_28008,N_21276,N_22323);
xnor U28009 (N_28009,N_24454,N_22423);
and U28010 (N_28010,N_24673,N_20091);
or U28011 (N_28011,N_22443,N_20303);
nand U28012 (N_28012,N_20676,N_24641);
or U28013 (N_28013,N_23294,N_24759);
and U28014 (N_28014,N_20749,N_20943);
nand U28015 (N_28015,N_20646,N_20059);
nand U28016 (N_28016,N_23114,N_23599);
nand U28017 (N_28017,N_20509,N_22862);
xor U28018 (N_28018,N_21297,N_22553);
or U28019 (N_28019,N_22279,N_20599);
or U28020 (N_28020,N_21168,N_22652);
nand U28021 (N_28021,N_22182,N_20212);
nand U28022 (N_28022,N_22172,N_22831);
nand U28023 (N_28023,N_23732,N_21822);
nor U28024 (N_28024,N_23961,N_24547);
or U28025 (N_28025,N_20790,N_22525);
nor U28026 (N_28026,N_21211,N_23713);
xnor U28027 (N_28027,N_22142,N_21675);
nand U28028 (N_28028,N_24848,N_23976);
or U28029 (N_28029,N_22199,N_20997);
nor U28030 (N_28030,N_22680,N_22757);
or U28031 (N_28031,N_22451,N_21179);
nor U28032 (N_28032,N_20010,N_23293);
nor U28033 (N_28033,N_22974,N_20811);
or U28034 (N_28034,N_22583,N_22494);
or U28035 (N_28035,N_20999,N_23049);
nand U28036 (N_28036,N_21151,N_22264);
nor U28037 (N_28037,N_22014,N_23528);
nor U28038 (N_28038,N_21719,N_21327);
and U28039 (N_28039,N_23860,N_24483);
xnor U28040 (N_28040,N_22971,N_22204);
nand U28041 (N_28041,N_24040,N_21561);
or U28042 (N_28042,N_20093,N_22154);
nand U28043 (N_28043,N_23513,N_23598);
or U28044 (N_28044,N_20073,N_20265);
or U28045 (N_28045,N_23961,N_21549);
nor U28046 (N_28046,N_24979,N_24033);
xnor U28047 (N_28047,N_20628,N_24840);
xor U28048 (N_28048,N_22240,N_20151);
xor U28049 (N_28049,N_24202,N_24669);
nand U28050 (N_28050,N_23370,N_23549);
xnor U28051 (N_28051,N_21821,N_21850);
nor U28052 (N_28052,N_23494,N_23699);
or U28053 (N_28053,N_20193,N_21711);
nor U28054 (N_28054,N_23421,N_22717);
or U28055 (N_28055,N_21452,N_21194);
nor U28056 (N_28056,N_23747,N_20116);
or U28057 (N_28057,N_23109,N_20439);
or U28058 (N_28058,N_22347,N_24353);
nand U28059 (N_28059,N_23234,N_23765);
nand U28060 (N_28060,N_22036,N_20014);
or U28061 (N_28061,N_21420,N_24979);
nor U28062 (N_28062,N_24423,N_21731);
and U28063 (N_28063,N_20632,N_21394);
and U28064 (N_28064,N_23279,N_24151);
nor U28065 (N_28065,N_23079,N_22507);
or U28066 (N_28066,N_23225,N_21065);
nor U28067 (N_28067,N_21553,N_20989);
nor U28068 (N_28068,N_21023,N_20192);
nand U28069 (N_28069,N_21052,N_21757);
xnor U28070 (N_28070,N_21899,N_20769);
and U28071 (N_28071,N_20048,N_20717);
xnor U28072 (N_28072,N_23830,N_23643);
or U28073 (N_28073,N_24586,N_23106);
nand U28074 (N_28074,N_20493,N_23862);
xnor U28075 (N_28075,N_20962,N_24741);
and U28076 (N_28076,N_20350,N_22832);
nor U28077 (N_28077,N_24331,N_20450);
nor U28078 (N_28078,N_23262,N_22556);
nand U28079 (N_28079,N_20984,N_23071);
nor U28080 (N_28080,N_20663,N_24494);
xor U28081 (N_28081,N_23743,N_22187);
or U28082 (N_28082,N_24248,N_21775);
nor U28083 (N_28083,N_21070,N_21502);
or U28084 (N_28084,N_22161,N_22645);
xor U28085 (N_28085,N_23886,N_20511);
and U28086 (N_28086,N_24562,N_24738);
nor U28087 (N_28087,N_20045,N_23485);
and U28088 (N_28088,N_23293,N_21605);
nor U28089 (N_28089,N_24904,N_21483);
or U28090 (N_28090,N_20482,N_22706);
nor U28091 (N_28091,N_22346,N_21529);
or U28092 (N_28092,N_23772,N_24091);
nor U28093 (N_28093,N_22476,N_20715);
xnor U28094 (N_28094,N_23360,N_23466);
nand U28095 (N_28095,N_23299,N_24571);
or U28096 (N_28096,N_21291,N_24262);
or U28097 (N_28097,N_24312,N_21641);
nor U28098 (N_28098,N_20842,N_24712);
and U28099 (N_28099,N_20989,N_23274);
or U28100 (N_28100,N_20213,N_22650);
and U28101 (N_28101,N_24668,N_20722);
or U28102 (N_28102,N_22757,N_21615);
xor U28103 (N_28103,N_21902,N_23764);
nand U28104 (N_28104,N_23519,N_21213);
nand U28105 (N_28105,N_24162,N_22951);
nor U28106 (N_28106,N_20619,N_23539);
nor U28107 (N_28107,N_22357,N_20638);
nor U28108 (N_28108,N_22431,N_21409);
and U28109 (N_28109,N_23416,N_22474);
or U28110 (N_28110,N_22411,N_22634);
nor U28111 (N_28111,N_21567,N_21525);
nor U28112 (N_28112,N_24676,N_21596);
or U28113 (N_28113,N_23021,N_20209);
and U28114 (N_28114,N_20704,N_20318);
or U28115 (N_28115,N_24748,N_23521);
nand U28116 (N_28116,N_20520,N_22900);
or U28117 (N_28117,N_21558,N_21950);
xor U28118 (N_28118,N_20596,N_24111);
or U28119 (N_28119,N_23375,N_23014);
and U28120 (N_28120,N_20087,N_23192);
xor U28121 (N_28121,N_24798,N_22219);
and U28122 (N_28122,N_23725,N_20505);
xor U28123 (N_28123,N_22201,N_22945);
nor U28124 (N_28124,N_21587,N_23958);
nor U28125 (N_28125,N_24102,N_21335);
xor U28126 (N_28126,N_24185,N_20075);
xnor U28127 (N_28127,N_23240,N_20675);
nand U28128 (N_28128,N_22898,N_23639);
and U28129 (N_28129,N_21034,N_20458);
nand U28130 (N_28130,N_23498,N_23413);
nor U28131 (N_28131,N_24510,N_20696);
nand U28132 (N_28132,N_21410,N_23058);
nand U28133 (N_28133,N_24809,N_22874);
nand U28134 (N_28134,N_20401,N_22079);
xnor U28135 (N_28135,N_23337,N_21809);
and U28136 (N_28136,N_24049,N_22079);
nand U28137 (N_28137,N_21824,N_21825);
nor U28138 (N_28138,N_24745,N_22988);
nand U28139 (N_28139,N_21049,N_24359);
xnor U28140 (N_28140,N_20989,N_21942);
and U28141 (N_28141,N_22062,N_20556);
and U28142 (N_28142,N_20362,N_21366);
or U28143 (N_28143,N_20194,N_24612);
nand U28144 (N_28144,N_21886,N_24647);
nand U28145 (N_28145,N_20658,N_22371);
and U28146 (N_28146,N_20590,N_22637);
or U28147 (N_28147,N_22339,N_21715);
xor U28148 (N_28148,N_23886,N_20809);
nand U28149 (N_28149,N_22590,N_24822);
and U28150 (N_28150,N_24740,N_24619);
nand U28151 (N_28151,N_20725,N_20318);
nor U28152 (N_28152,N_21472,N_20878);
nand U28153 (N_28153,N_22569,N_23128);
nand U28154 (N_28154,N_23839,N_23422);
nand U28155 (N_28155,N_21693,N_22333);
nand U28156 (N_28156,N_20009,N_24107);
or U28157 (N_28157,N_21372,N_21222);
nand U28158 (N_28158,N_24229,N_23096);
nor U28159 (N_28159,N_22219,N_20083);
xnor U28160 (N_28160,N_23070,N_22595);
nor U28161 (N_28161,N_21044,N_22308);
or U28162 (N_28162,N_24119,N_23386);
xnor U28163 (N_28163,N_21805,N_23917);
nand U28164 (N_28164,N_21292,N_24673);
and U28165 (N_28165,N_24940,N_20716);
xor U28166 (N_28166,N_24779,N_23309);
nor U28167 (N_28167,N_22620,N_23492);
and U28168 (N_28168,N_21985,N_21591);
or U28169 (N_28169,N_24526,N_23592);
nor U28170 (N_28170,N_22370,N_24829);
nor U28171 (N_28171,N_24371,N_23672);
nor U28172 (N_28172,N_22499,N_22156);
xor U28173 (N_28173,N_20279,N_23467);
nor U28174 (N_28174,N_23770,N_24397);
or U28175 (N_28175,N_22274,N_21907);
and U28176 (N_28176,N_22726,N_22224);
or U28177 (N_28177,N_22137,N_21412);
nand U28178 (N_28178,N_21314,N_22967);
and U28179 (N_28179,N_22891,N_20001);
xnor U28180 (N_28180,N_20570,N_20730);
and U28181 (N_28181,N_23599,N_22082);
or U28182 (N_28182,N_21541,N_21601);
nor U28183 (N_28183,N_22221,N_23957);
xor U28184 (N_28184,N_22604,N_24380);
and U28185 (N_28185,N_21026,N_21316);
nand U28186 (N_28186,N_21767,N_24993);
nand U28187 (N_28187,N_20370,N_20955);
and U28188 (N_28188,N_20724,N_21962);
xor U28189 (N_28189,N_22693,N_20683);
nor U28190 (N_28190,N_24592,N_21051);
xor U28191 (N_28191,N_20505,N_23520);
or U28192 (N_28192,N_21699,N_22906);
nor U28193 (N_28193,N_20760,N_20886);
xnor U28194 (N_28194,N_21427,N_22475);
nand U28195 (N_28195,N_24140,N_24340);
nor U28196 (N_28196,N_20802,N_20798);
and U28197 (N_28197,N_23044,N_20574);
nand U28198 (N_28198,N_24842,N_22158);
nand U28199 (N_28199,N_24165,N_20894);
nand U28200 (N_28200,N_24133,N_21825);
and U28201 (N_28201,N_20448,N_24627);
or U28202 (N_28202,N_23605,N_20504);
and U28203 (N_28203,N_20041,N_20346);
and U28204 (N_28204,N_22160,N_21759);
xor U28205 (N_28205,N_20808,N_21235);
nand U28206 (N_28206,N_23753,N_23372);
and U28207 (N_28207,N_22431,N_21768);
nor U28208 (N_28208,N_20319,N_22045);
xor U28209 (N_28209,N_24097,N_24717);
or U28210 (N_28210,N_20998,N_21108);
nor U28211 (N_28211,N_21530,N_20785);
or U28212 (N_28212,N_21302,N_20247);
and U28213 (N_28213,N_21857,N_20369);
nand U28214 (N_28214,N_23912,N_20463);
xor U28215 (N_28215,N_20114,N_21829);
nor U28216 (N_28216,N_20833,N_22534);
nor U28217 (N_28217,N_20533,N_24120);
or U28218 (N_28218,N_23066,N_24952);
or U28219 (N_28219,N_20883,N_23137);
xor U28220 (N_28220,N_24416,N_22407);
nor U28221 (N_28221,N_22224,N_24622);
or U28222 (N_28222,N_23785,N_23503);
nor U28223 (N_28223,N_22009,N_24826);
nor U28224 (N_28224,N_22314,N_20109);
and U28225 (N_28225,N_24633,N_20815);
nor U28226 (N_28226,N_21073,N_20901);
nand U28227 (N_28227,N_21165,N_24105);
or U28228 (N_28228,N_20895,N_24402);
xor U28229 (N_28229,N_20011,N_23165);
or U28230 (N_28230,N_21453,N_24316);
nor U28231 (N_28231,N_21789,N_21710);
nor U28232 (N_28232,N_22953,N_20490);
nor U28233 (N_28233,N_22765,N_20091);
and U28234 (N_28234,N_20692,N_21395);
xor U28235 (N_28235,N_20191,N_22329);
xor U28236 (N_28236,N_24860,N_21187);
xor U28237 (N_28237,N_21274,N_22400);
nor U28238 (N_28238,N_21624,N_22050);
xnor U28239 (N_28239,N_21889,N_24172);
or U28240 (N_28240,N_20985,N_20228);
nand U28241 (N_28241,N_22154,N_21583);
nand U28242 (N_28242,N_20995,N_24382);
or U28243 (N_28243,N_21638,N_21442);
nor U28244 (N_28244,N_24313,N_24558);
or U28245 (N_28245,N_23636,N_20358);
nor U28246 (N_28246,N_24250,N_21000);
nand U28247 (N_28247,N_23295,N_20078);
and U28248 (N_28248,N_24121,N_22292);
and U28249 (N_28249,N_23289,N_22966);
nand U28250 (N_28250,N_23916,N_21653);
nand U28251 (N_28251,N_21421,N_21263);
nand U28252 (N_28252,N_24498,N_20976);
nor U28253 (N_28253,N_22238,N_23769);
nand U28254 (N_28254,N_20626,N_24441);
nor U28255 (N_28255,N_22848,N_24592);
or U28256 (N_28256,N_23761,N_20632);
nor U28257 (N_28257,N_20781,N_23946);
and U28258 (N_28258,N_20104,N_23222);
nand U28259 (N_28259,N_20264,N_22321);
xnor U28260 (N_28260,N_21189,N_22581);
nor U28261 (N_28261,N_20220,N_22566);
nand U28262 (N_28262,N_20058,N_22359);
nor U28263 (N_28263,N_24520,N_21490);
xnor U28264 (N_28264,N_21377,N_23961);
nand U28265 (N_28265,N_21873,N_21149);
nor U28266 (N_28266,N_24572,N_20419);
or U28267 (N_28267,N_23685,N_20877);
nor U28268 (N_28268,N_22902,N_21280);
and U28269 (N_28269,N_23428,N_23575);
or U28270 (N_28270,N_24569,N_24017);
and U28271 (N_28271,N_21577,N_24597);
and U28272 (N_28272,N_22411,N_20079);
xor U28273 (N_28273,N_20049,N_20277);
xor U28274 (N_28274,N_22223,N_22230);
and U28275 (N_28275,N_23151,N_23397);
xnor U28276 (N_28276,N_22900,N_22588);
and U28277 (N_28277,N_22088,N_23756);
and U28278 (N_28278,N_21927,N_21034);
nor U28279 (N_28279,N_24034,N_20492);
nand U28280 (N_28280,N_20103,N_23593);
and U28281 (N_28281,N_20321,N_22387);
xor U28282 (N_28282,N_24279,N_21495);
nand U28283 (N_28283,N_23958,N_21504);
nand U28284 (N_28284,N_21109,N_21983);
and U28285 (N_28285,N_22386,N_21645);
and U28286 (N_28286,N_20793,N_24201);
xnor U28287 (N_28287,N_20062,N_24810);
nor U28288 (N_28288,N_24897,N_22820);
or U28289 (N_28289,N_22676,N_21676);
nand U28290 (N_28290,N_21100,N_20477);
or U28291 (N_28291,N_20705,N_22284);
xnor U28292 (N_28292,N_23330,N_21812);
nand U28293 (N_28293,N_22341,N_20764);
and U28294 (N_28294,N_23637,N_21324);
nor U28295 (N_28295,N_21080,N_22015);
and U28296 (N_28296,N_22884,N_23066);
or U28297 (N_28297,N_24535,N_21549);
nand U28298 (N_28298,N_22627,N_24060);
nand U28299 (N_28299,N_23785,N_24489);
nand U28300 (N_28300,N_23556,N_20418);
or U28301 (N_28301,N_20955,N_21874);
and U28302 (N_28302,N_23981,N_24008);
xnor U28303 (N_28303,N_23383,N_24716);
or U28304 (N_28304,N_21389,N_21012);
nand U28305 (N_28305,N_23729,N_24608);
and U28306 (N_28306,N_24128,N_22442);
xor U28307 (N_28307,N_24932,N_23688);
nor U28308 (N_28308,N_24608,N_24779);
or U28309 (N_28309,N_20754,N_22440);
nor U28310 (N_28310,N_24860,N_23024);
and U28311 (N_28311,N_21637,N_22246);
or U28312 (N_28312,N_22143,N_20907);
or U28313 (N_28313,N_22800,N_20204);
nor U28314 (N_28314,N_21187,N_24755);
nor U28315 (N_28315,N_21689,N_22119);
xnor U28316 (N_28316,N_24105,N_20112);
and U28317 (N_28317,N_20303,N_24342);
nand U28318 (N_28318,N_21955,N_23039);
nor U28319 (N_28319,N_20541,N_20602);
xor U28320 (N_28320,N_20815,N_24758);
nor U28321 (N_28321,N_23056,N_22947);
and U28322 (N_28322,N_23969,N_24172);
xnor U28323 (N_28323,N_24870,N_22400);
or U28324 (N_28324,N_23562,N_20394);
or U28325 (N_28325,N_20569,N_24579);
or U28326 (N_28326,N_21985,N_20596);
or U28327 (N_28327,N_22509,N_21728);
or U28328 (N_28328,N_22079,N_23868);
xor U28329 (N_28329,N_24755,N_24696);
or U28330 (N_28330,N_24997,N_20494);
nor U28331 (N_28331,N_20169,N_24137);
nand U28332 (N_28332,N_22848,N_24710);
nand U28333 (N_28333,N_24042,N_20224);
or U28334 (N_28334,N_21090,N_23061);
xnor U28335 (N_28335,N_24864,N_20669);
nand U28336 (N_28336,N_22266,N_21059);
and U28337 (N_28337,N_24176,N_24582);
xor U28338 (N_28338,N_21166,N_21839);
or U28339 (N_28339,N_21233,N_22954);
and U28340 (N_28340,N_24309,N_22542);
nor U28341 (N_28341,N_22069,N_21326);
and U28342 (N_28342,N_22878,N_23610);
and U28343 (N_28343,N_22477,N_24280);
xnor U28344 (N_28344,N_24723,N_20802);
xnor U28345 (N_28345,N_21809,N_21617);
or U28346 (N_28346,N_21667,N_23476);
and U28347 (N_28347,N_23226,N_23491);
or U28348 (N_28348,N_23598,N_23179);
and U28349 (N_28349,N_23421,N_22743);
and U28350 (N_28350,N_24011,N_24223);
or U28351 (N_28351,N_23232,N_24163);
and U28352 (N_28352,N_22993,N_22291);
and U28353 (N_28353,N_23747,N_20553);
xnor U28354 (N_28354,N_22506,N_21381);
and U28355 (N_28355,N_24091,N_23673);
nor U28356 (N_28356,N_20447,N_24021);
xor U28357 (N_28357,N_22346,N_22577);
xor U28358 (N_28358,N_23227,N_22429);
xor U28359 (N_28359,N_23816,N_24870);
and U28360 (N_28360,N_21836,N_20071);
nor U28361 (N_28361,N_22363,N_20171);
or U28362 (N_28362,N_21189,N_24694);
nand U28363 (N_28363,N_20928,N_22977);
xnor U28364 (N_28364,N_23086,N_24932);
and U28365 (N_28365,N_23121,N_22365);
nand U28366 (N_28366,N_20385,N_23098);
nor U28367 (N_28367,N_24984,N_20639);
and U28368 (N_28368,N_21272,N_24203);
xnor U28369 (N_28369,N_22233,N_21244);
or U28370 (N_28370,N_22724,N_24320);
xor U28371 (N_28371,N_24173,N_20000);
nor U28372 (N_28372,N_24555,N_24037);
or U28373 (N_28373,N_24664,N_21500);
nand U28374 (N_28374,N_20000,N_23697);
nand U28375 (N_28375,N_21606,N_20828);
xnor U28376 (N_28376,N_24701,N_23706);
and U28377 (N_28377,N_21777,N_22955);
and U28378 (N_28378,N_20058,N_23389);
nand U28379 (N_28379,N_24893,N_22394);
xor U28380 (N_28380,N_21133,N_22271);
xnor U28381 (N_28381,N_23186,N_21657);
or U28382 (N_28382,N_22786,N_20215);
nand U28383 (N_28383,N_20534,N_21018);
nor U28384 (N_28384,N_21089,N_23807);
nand U28385 (N_28385,N_21251,N_20954);
and U28386 (N_28386,N_20188,N_22841);
and U28387 (N_28387,N_23060,N_24043);
and U28388 (N_28388,N_21524,N_21041);
or U28389 (N_28389,N_21520,N_24424);
xor U28390 (N_28390,N_20000,N_20177);
nand U28391 (N_28391,N_23643,N_21036);
nand U28392 (N_28392,N_20517,N_24606);
xor U28393 (N_28393,N_22199,N_22342);
nor U28394 (N_28394,N_20449,N_21742);
xnor U28395 (N_28395,N_23925,N_22923);
xor U28396 (N_28396,N_22912,N_21758);
and U28397 (N_28397,N_24895,N_20651);
nand U28398 (N_28398,N_21324,N_24904);
and U28399 (N_28399,N_24405,N_23587);
xnor U28400 (N_28400,N_24364,N_21326);
nor U28401 (N_28401,N_20671,N_20801);
and U28402 (N_28402,N_20693,N_24155);
nand U28403 (N_28403,N_22275,N_22351);
or U28404 (N_28404,N_21355,N_20124);
or U28405 (N_28405,N_21368,N_23843);
nor U28406 (N_28406,N_22012,N_21069);
and U28407 (N_28407,N_23691,N_23107);
xor U28408 (N_28408,N_24317,N_22855);
nor U28409 (N_28409,N_21589,N_20972);
nand U28410 (N_28410,N_24879,N_21583);
and U28411 (N_28411,N_24885,N_23322);
xor U28412 (N_28412,N_24096,N_22093);
xor U28413 (N_28413,N_21078,N_20269);
nor U28414 (N_28414,N_21682,N_22446);
and U28415 (N_28415,N_23243,N_24319);
nand U28416 (N_28416,N_20181,N_24059);
nand U28417 (N_28417,N_24265,N_20822);
or U28418 (N_28418,N_23223,N_22572);
nor U28419 (N_28419,N_21608,N_23462);
or U28420 (N_28420,N_23185,N_24742);
or U28421 (N_28421,N_21973,N_21159);
and U28422 (N_28422,N_21584,N_22802);
and U28423 (N_28423,N_23086,N_22560);
xor U28424 (N_28424,N_20823,N_21524);
and U28425 (N_28425,N_24020,N_24877);
xor U28426 (N_28426,N_21811,N_20543);
nor U28427 (N_28427,N_24668,N_22031);
nand U28428 (N_28428,N_21345,N_24993);
xnor U28429 (N_28429,N_20972,N_21784);
xnor U28430 (N_28430,N_24774,N_23644);
nor U28431 (N_28431,N_20902,N_21487);
or U28432 (N_28432,N_20904,N_24024);
or U28433 (N_28433,N_24589,N_23099);
xnor U28434 (N_28434,N_24967,N_23366);
and U28435 (N_28435,N_21208,N_20785);
xor U28436 (N_28436,N_23657,N_24807);
xnor U28437 (N_28437,N_24929,N_22332);
xor U28438 (N_28438,N_24779,N_23801);
nor U28439 (N_28439,N_23377,N_20817);
and U28440 (N_28440,N_21714,N_24260);
nand U28441 (N_28441,N_23478,N_22161);
and U28442 (N_28442,N_22245,N_20297);
and U28443 (N_28443,N_21636,N_22489);
and U28444 (N_28444,N_24613,N_21817);
xor U28445 (N_28445,N_20508,N_23980);
or U28446 (N_28446,N_22325,N_24233);
and U28447 (N_28447,N_21350,N_22340);
nand U28448 (N_28448,N_22043,N_21467);
xnor U28449 (N_28449,N_20079,N_20997);
or U28450 (N_28450,N_20682,N_23365);
or U28451 (N_28451,N_22762,N_21615);
and U28452 (N_28452,N_22217,N_22174);
or U28453 (N_28453,N_20076,N_22065);
or U28454 (N_28454,N_21246,N_20075);
nor U28455 (N_28455,N_21385,N_22388);
or U28456 (N_28456,N_20727,N_24238);
or U28457 (N_28457,N_22187,N_23592);
and U28458 (N_28458,N_20592,N_22189);
or U28459 (N_28459,N_21630,N_21475);
xnor U28460 (N_28460,N_20972,N_23515);
or U28461 (N_28461,N_24048,N_24985);
or U28462 (N_28462,N_20230,N_23848);
xnor U28463 (N_28463,N_24013,N_24660);
nand U28464 (N_28464,N_23463,N_21791);
nor U28465 (N_28465,N_20791,N_24685);
or U28466 (N_28466,N_23725,N_24442);
nand U28467 (N_28467,N_24196,N_20113);
xor U28468 (N_28468,N_24107,N_23424);
nor U28469 (N_28469,N_20236,N_23385);
nor U28470 (N_28470,N_22773,N_22400);
nand U28471 (N_28471,N_23588,N_22661);
or U28472 (N_28472,N_20296,N_21243);
nor U28473 (N_28473,N_22211,N_22834);
and U28474 (N_28474,N_23386,N_22963);
nand U28475 (N_28475,N_24258,N_22493);
nor U28476 (N_28476,N_21010,N_24021);
xor U28477 (N_28477,N_22590,N_23329);
xnor U28478 (N_28478,N_22635,N_23319);
nor U28479 (N_28479,N_20385,N_20492);
nor U28480 (N_28480,N_22253,N_20540);
nand U28481 (N_28481,N_22356,N_21245);
or U28482 (N_28482,N_21260,N_24888);
xnor U28483 (N_28483,N_22691,N_21490);
and U28484 (N_28484,N_22262,N_20239);
nor U28485 (N_28485,N_24000,N_20413);
nor U28486 (N_28486,N_24514,N_24103);
and U28487 (N_28487,N_21330,N_21975);
xor U28488 (N_28488,N_23994,N_22547);
or U28489 (N_28489,N_24024,N_20213);
or U28490 (N_28490,N_20775,N_24854);
nand U28491 (N_28491,N_23861,N_24469);
or U28492 (N_28492,N_24805,N_24839);
or U28493 (N_28493,N_22892,N_24191);
nand U28494 (N_28494,N_23950,N_22222);
and U28495 (N_28495,N_23613,N_22013);
xnor U28496 (N_28496,N_24887,N_23463);
or U28497 (N_28497,N_20413,N_20317);
nor U28498 (N_28498,N_21339,N_20864);
xor U28499 (N_28499,N_20530,N_23925);
xor U28500 (N_28500,N_21862,N_22387);
nor U28501 (N_28501,N_20245,N_20678);
xor U28502 (N_28502,N_22859,N_20502);
xor U28503 (N_28503,N_21273,N_23613);
nand U28504 (N_28504,N_24225,N_20795);
and U28505 (N_28505,N_20238,N_20752);
xnor U28506 (N_28506,N_20281,N_20955);
nand U28507 (N_28507,N_22380,N_23937);
or U28508 (N_28508,N_22340,N_24347);
nor U28509 (N_28509,N_21892,N_24892);
nor U28510 (N_28510,N_24072,N_24993);
or U28511 (N_28511,N_21192,N_23349);
nor U28512 (N_28512,N_22066,N_21415);
and U28513 (N_28513,N_20006,N_23989);
xor U28514 (N_28514,N_21662,N_21112);
nand U28515 (N_28515,N_22445,N_24432);
or U28516 (N_28516,N_21985,N_20526);
nor U28517 (N_28517,N_22974,N_23550);
nand U28518 (N_28518,N_24780,N_24270);
and U28519 (N_28519,N_21530,N_20524);
xor U28520 (N_28520,N_23952,N_23268);
xor U28521 (N_28521,N_21368,N_20813);
nor U28522 (N_28522,N_23416,N_24151);
or U28523 (N_28523,N_20143,N_22987);
xor U28524 (N_28524,N_22392,N_23709);
or U28525 (N_28525,N_20738,N_22518);
nand U28526 (N_28526,N_23973,N_21287);
or U28527 (N_28527,N_20804,N_23926);
nand U28528 (N_28528,N_21527,N_21554);
nand U28529 (N_28529,N_20457,N_24489);
xnor U28530 (N_28530,N_20207,N_21532);
and U28531 (N_28531,N_23890,N_23344);
and U28532 (N_28532,N_22169,N_24702);
nor U28533 (N_28533,N_21175,N_24372);
or U28534 (N_28534,N_20973,N_21037);
or U28535 (N_28535,N_21696,N_20674);
xnor U28536 (N_28536,N_23863,N_21125);
and U28537 (N_28537,N_22852,N_21146);
nand U28538 (N_28538,N_20632,N_23534);
nand U28539 (N_28539,N_24658,N_21583);
or U28540 (N_28540,N_24410,N_21814);
nand U28541 (N_28541,N_23683,N_20113);
nand U28542 (N_28542,N_23827,N_23683);
nor U28543 (N_28543,N_21657,N_20108);
xor U28544 (N_28544,N_24378,N_20516);
xnor U28545 (N_28545,N_20806,N_22081);
or U28546 (N_28546,N_23301,N_23522);
nand U28547 (N_28547,N_24295,N_20150);
xor U28548 (N_28548,N_23738,N_20475);
nand U28549 (N_28549,N_22653,N_24694);
nor U28550 (N_28550,N_23900,N_20184);
or U28551 (N_28551,N_23388,N_21532);
nand U28552 (N_28552,N_21412,N_20563);
nor U28553 (N_28553,N_24387,N_23645);
nand U28554 (N_28554,N_21869,N_23374);
nand U28555 (N_28555,N_21618,N_21603);
nor U28556 (N_28556,N_23765,N_21787);
and U28557 (N_28557,N_20792,N_24010);
or U28558 (N_28558,N_24210,N_22919);
nor U28559 (N_28559,N_23492,N_23357);
or U28560 (N_28560,N_24388,N_21238);
xor U28561 (N_28561,N_23824,N_23092);
or U28562 (N_28562,N_23273,N_20449);
nor U28563 (N_28563,N_22410,N_24017);
nand U28564 (N_28564,N_21290,N_24837);
nand U28565 (N_28565,N_23023,N_20751);
and U28566 (N_28566,N_20407,N_22541);
xor U28567 (N_28567,N_20527,N_21260);
nor U28568 (N_28568,N_22634,N_24921);
or U28569 (N_28569,N_20355,N_21530);
and U28570 (N_28570,N_21483,N_23785);
and U28571 (N_28571,N_24567,N_21647);
nor U28572 (N_28572,N_21036,N_24177);
nor U28573 (N_28573,N_23728,N_20904);
xnor U28574 (N_28574,N_22375,N_23176);
nand U28575 (N_28575,N_23559,N_20215);
xnor U28576 (N_28576,N_24867,N_21905);
xor U28577 (N_28577,N_20063,N_20568);
nand U28578 (N_28578,N_24247,N_23354);
nor U28579 (N_28579,N_24584,N_24781);
nand U28580 (N_28580,N_21759,N_24207);
nor U28581 (N_28581,N_24730,N_21102);
and U28582 (N_28582,N_20434,N_20509);
nand U28583 (N_28583,N_20235,N_22854);
and U28584 (N_28584,N_21145,N_23571);
or U28585 (N_28585,N_23362,N_23040);
or U28586 (N_28586,N_24126,N_23218);
xnor U28587 (N_28587,N_20938,N_21375);
or U28588 (N_28588,N_21496,N_20447);
nor U28589 (N_28589,N_23754,N_20719);
and U28590 (N_28590,N_20018,N_20249);
and U28591 (N_28591,N_24674,N_24869);
and U28592 (N_28592,N_22678,N_24090);
nand U28593 (N_28593,N_23289,N_23621);
nor U28594 (N_28594,N_21472,N_20461);
xor U28595 (N_28595,N_21996,N_22391);
or U28596 (N_28596,N_20054,N_23904);
or U28597 (N_28597,N_20084,N_24119);
nand U28598 (N_28598,N_22823,N_20210);
or U28599 (N_28599,N_23510,N_20730);
nor U28600 (N_28600,N_24713,N_24122);
and U28601 (N_28601,N_20427,N_21638);
nand U28602 (N_28602,N_20946,N_23285);
nand U28603 (N_28603,N_22649,N_21035);
or U28604 (N_28604,N_20772,N_23710);
xor U28605 (N_28605,N_21402,N_22609);
nor U28606 (N_28606,N_21862,N_23479);
or U28607 (N_28607,N_23614,N_21551);
nand U28608 (N_28608,N_22864,N_24480);
and U28609 (N_28609,N_23301,N_21725);
xor U28610 (N_28610,N_24140,N_21739);
nand U28611 (N_28611,N_20719,N_21404);
xor U28612 (N_28612,N_23306,N_20447);
nand U28613 (N_28613,N_22756,N_20871);
or U28614 (N_28614,N_22362,N_21865);
nand U28615 (N_28615,N_22028,N_21961);
and U28616 (N_28616,N_24268,N_21249);
nand U28617 (N_28617,N_22611,N_22512);
nor U28618 (N_28618,N_23301,N_20431);
or U28619 (N_28619,N_22806,N_20910);
xor U28620 (N_28620,N_20676,N_20417);
xor U28621 (N_28621,N_23212,N_24385);
nand U28622 (N_28622,N_22596,N_20071);
nor U28623 (N_28623,N_21084,N_23308);
or U28624 (N_28624,N_23525,N_20961);
xor U28625 (N_28625,N_23377,N_24419);
nor U28626 (N_28626,N_21186,N_23372);
nand U28627 (N_28627,N_22128,N_22737);
nor U28628 (N_28628,N_23603,N_22899);
and U28629 (N_28629,N_21066,N_24801);
nand U28630 (N_28630,N_21781,N_24983);
xor U28631 (N_28631,N_24660,N_21047);
nand U28632 (N_28632,N_24968,N_24561);
or U28633 (N_28633,N_22413,N_21858);
nor U28634 (N_28634,N_20953,N_22152);
xor U28635 (N_28635,N_20952,N_22735);
and U28636 (N_28636,N_23977,N_24656);
nor U28637 (N_28637,N_23308,N_21280);
or U28638 (N_28638,N_24173,N_21589);
nand U28639 (N_28639,N_22136,N_20515);
xnor U28640 (N_28640,N_24544,N_20304);
or U28641 (N_28641,N_22232,N_22778);
nand U28642 (N_28642,N_20589,N_24801);
or U28643 (N_28643,N_20289,N_24560);
and U28644 (N_28644,N_20426,N_21651);
and U28645 (N_28645,N_24828,N_21571);
nand U28646 (N_28646,N_21192,N_24787);
nand U28647 (N_28647,N_24677,N_24027);
xnor U28648 (N_28648,N_23319,N_20471);
nor U28649 (N_28649,N_20664,N_22483);
nand U28650 (N_28650,N_24941,N_23081);
or U28651 (N_28651,N_23222,N_23995);
or U28652 (N_28652,N_23747,N_22080);
or U28653 (N_28653,N_20295,N_20043);
nor U28654 (N_28654,N_22888,N_24373);
xor U28655 (N_28655,N_21789,N_24743);
nor U28656 (N_28656,N_24036,N_21809);
nand U28657 (N_28657,N_24860,N_21546);
nand U28658 (N_28658,N_21266,N_20127);
and U28659 (N_28659,N_22323,N_22230);
nand U28660 (N_28660,N_23717,N_20413);
or U28661 (N_28661,N_23771,N_24711);
or U28662 (N_28662,N_22549,N_23131);
and U28663 (N_28663,N_23399,N_24275);
nor U28664 (N_28664,N_23427,N_20707);
xnor U28665 (N_28665,N_23947,N_22556);
nor U28666 (N_28666,N_24483,N_20425);
xor U28667 (N_28667,N_20435,N_22607);
nand U28668 (N_28668,N_21661,N_21295);
or U28669 (N_28669,N_24101,N_20051);
or U28670 (N_28670,N_20509,N_23066);
or U28671 (N_28671,N_24127,N_22933);
nand U28672 (N_28672,N_24121,N_22804);
xnor U28673 (N_28673,N_20269,N_22722);
or U28674 (N_28674,N_24510,N_21872);
nor U28675 (N_28675,N_24820,N_22068);
xnor U28676 (N_28676,N_21834,N_22171);
nand U28677 (N_28677,N_23793,N_20717);
or U28678 (N_28678,N_21487,N_24094);
and U28679 (N_28679,N_23015,N_21613);
nor U28680 (N_28680,N_21456,N_23874);
xor U28681 (N_28681,N_21669,N_22968);
and U28682 (N_28682,N_24240,N_24842);
and U28683 (N_28683,N_23284,N_21182);
or U28684 (N_28684,N_20289,N_21821);
xnor U28685 (N_28685,N_23370,N_24267);
or U28686 (N_28686,N_20965,N_23205);
and U28687 (N_28687,N_23100,N_23799);
or U28688 (N_28688,N_22606,N_22191);
nor U28689 (N_28689,N_22613,N_21095);
or U28690 (N_28690,N_20225,N_22739);
nand U28691 (N_28691,N_21269,N_23175);
or U28692 (N_28692,N_23127,N_23210);
nor U28693 (N_28693,N_23356,N_20078);
nand U28694 (N_28694,N_20898,N_20044);
and U28695 (N_28695,N_20394,N_22387);
or U28696 (N_28696,N_22881,N_24379);
xor U28697 (N_28697,N_24944,N_22592);
and U28698 (N_28698,N_24115,N_21538);
and U28699 (N_28699,N_22696,N_24220);
or U28700 (N_28700,N_21281,N_23493);
nor U28701 (N_28701,N_24465,N_23553);
nand U28702 (N_28702,N_23734,N_21623);
xnor U28703 (N_28703,N_23612,N_21572);
or U28704 (N_28704,N_23755,N_23127);
xnor U28705 (N_28705,N_23478,N_21927);
nor U28706 (N_28706,N_21376,N_20499);
nand U28707 (N_28707,N_24464,N_20449);
xnor U28708 (N_28708,N_22950,N_23187);
and U28709 (N_28709,N_24862,N_21182);
xor U28710 (N_28710,N_23096,N_24832);
or U28711 (N_28711,N_22719,N_23032);
nand U28712 (N_28712,N_23464,N_20891);
nand U28713 (N_28713,N_20254,N_21940);
nor U28714 (N_28714,N_24001,N_20738);
or U28715 (N_28715,N_22785,N_23401);
and U28716 (N_28716,N_24839,N_21600);
nor U28717 (N_28717,N_22482,N_20217);
xnor U28718 (N_28718,N_24423,N_22969);
xor U28719 (N_28719,N_23126,N_24974);
or U28720 (N_28720,N_21968,N_23472);
xor U28721 (N_28721,N_23206,N_22816);
nand U28722 (N_28722,N_21404,N_20774);
and U28723 (N_28723,N_23599,N_22286);
or U28724 (N_28724,N_23436,N_24802);
and U28725 (N_28725,N_21404,N_22028);
xnor U28726 (N_28726,N_21998,N_23370);
and U28727 (N_28727,N_20307,N_20676);
xnor U28728 (N_28728,N_24804,N_21721);
and U28729 (N_28729,N_23296,N_23910);
nand U28730 (N_28730,N_23756,N_20220);
xor U28731 (N_28731,N_22254,N_24832);
nor U28732 (N_28732,N_24571,N_23767);
and U28733 (N_28733,N_22643,N_20396);
nor U28734 (N_28734,N_22769,N_23871);
xnor U28735 (N_28735,N_24782,N_20259);
nor U28736 (N_28736,N_24815,N_20487);
and U28737 (N_28737,N_22959,N_20691);
and U28738 (N_28738,N_21809,N_22269);
nand U28739 (N_28739,N_20921,N_20496);
nand U28740 (N_28740,N_22679,N_20033);
xor U28741 (N_28741,N_24959,N_24188);
and U28742 (N_28742,N_22155,N_21616);
nand U28743 (N_28743,N_24392,N_21059);
nand U28744 (N_28744,N_24442,N_22922);
nor U28745 (N_28745,N_21948,N_20212);
and U28746 (N_28746,N_20788,N_23807);
and U28747 (N_28747,N_24877,N_23813);
nor U28748 (N_28748,N_23108,N_24644);
nand U28749 (N_28749,N_21887,N_23617);
xnor U28750 (N_28750,N_20906,N_20903);
and U28751 (N_28751,N_23537,N_22833);
nand U28752 (N_28752,N_23664,N_24472);
nand U28753 (N_28753,N_20229,N_21431);
xnor U28754 (N_28754,N_23506,N_22964);
xnor U28755 (N_28755,N_21743,N_22955);
or U28756 (N_28756,N_20099,N_24433);
or U28757 (N_28757,N_21431,N_20779);
or U28758 (N_28758,N_24461,N_23980);
xor U28759 (N_28759,N_21815,N_24588);
and U28760 (N_28760,N_21522,N_23216);
xor U28761 (N_28761,N_20065,N_24164);
nor U28762 (N_28762,N_23808,N_24071);
nor U28763 (N_28763,N_21075,N_22136);
and U28764 (N_28764,N_22244,N_23189);
nand U28765 (N_28765,N_20646,N_21568);
xnor U28766 (N_28766,N_22170,N_20734);
nand U28767 (N_28767,N_21020,N_20055);
xnor U28768 (N_28768,N_23895,N_23294);
and U28769 (N_28769,N_22208,N_23260);
nand U28770 (N_28770,N_24131,N_23211);
nor U28771 (N_28771,N_21607,N_23616);
nand U28772 (N_28772,N_21718,N_21499);
nand U28773 (N_28773,N_22717,N_24780);
nand U28774 (N_28774,N_22592,N_20603);
nor U28775 (N_28775,N_22149,N_24523);
xnor U28776 (N_28776,N_21653,N_22905);
xnor U28777 (N_28777,N_24116,N_22640);
xor U28778 (N_28778,N_21099,N_24141);
or U28779 (N_28779,N_20865,N_21046);
or U28780 (N_28780,N_21770,N_24744);
nand U28781 (N_28781,N_20786,N_21981);
or U28782 (N_28782,N_22271,N_24754);
nor U28783 (N_28783,N_23974,N_24451);
xor U28784 (N_28784,N_21041,N_23656);
or U28785 (N_28785,N_20460,N_20581);
xnor U28786 (N_28786,N_21100,N_22836);
nor U28787 (N_28787,N_23700,N_20997);
nor U28788 (N_28788,N_23285,N_21806);
nand U28789 (N_28789,N_20340,N_20053);
or U28790 (N_28790,N_22815,N_20916);
xor U28791 (N_28791,N_24366,N_23395);
and U28792 (N_28792,N_21596,N_20673);
nor U28793 (N_28793,N_20931,N_24101);
or U28794 (N_28794,N_20236,N_21078);
xnor U28795 (N_28795,N_23480,N_20816);
xor U28796 (N_28796,N_20426,N_21036);
nor U28797 (N_28797,N_22154,N_24051);
or U28798 (N_28798,N_23578,N_20305);
nor U28799 (N_28799,N_24930,N_22096);
xor U28800 (N_28800,N_24932,N_22194);
or U28801 (N_28801,N_20887,N_24535);
and U28802 (N_28802,N_20483,N_22577);
or U28803 (N_28803,N_23585,N_24852);
xor U28804 (N_28804,N_22685,N_21703);
xor U28805 (N_28805,N_20656,N_21004);
xnor U28806 (N_28806,N_20531,N_22934);
or U28807 (N_28807,N_24432,N_23093);
xnor U28808 (N_28808,N_23256,N_24233);
or U28809 (N_28809,N_21119,N_23363);
nor U28810 (N_28810,N_22957,N_23243);
xor U28811 (N_28811,N_23284,N_23348);
nand U28812 (N_28812,N_24015,N_24293);
nand U28813 (N_28813,N_22948,N_21364);
xor U28814 (N_28814,N_20846,N_22211);
nand U28815 (N_28815,N_23624,N_22975);
and U28816 (N_28816,N_24962,N_21149);
and U28817 (N_28817,N_24934,N_21146);
xnor U28818 (N_28818,N_20079,N_21372);
nand U28819 (N_28819,N_22340,N_21434);
or U28820 (N_28820,N_20961,N_21289);
nor U28821 (N_28821,N_23927,N_22431);
nor U28822 (N_28822,N_24368,N_21155);
and U28823 (N_28823,N_22238,N_22777);
xnor U28824 (N_28824,N_23765,N_23480);
and U28825 (N_28825,N_20872,N_22875);
nand U28826 (N_28826,N_24758,N_23891);
or U28827 (N_28827,N_22417,N_22292);
xor U28828 (N_28828,N_23868,N_21328);
nand U28829 (N_28829,N_22487,N_24934);
and U28830 (N_28830,N_22691,N_23915);
or U28831 (N_28831,N_23130,N_20823);
and U28832 (N_28832,N_22918,N_22498);
nor U28833 (N_28833,N_20990,N_21118);
and U28834 (N_28834,N_24057,N_21370);
nor U28835 (N_28835,N_20058,N_22071);
nand U28836 (N_28836,N_22700,N_23662);
nand U28837 (N_28837,N_23696,N_23797);
xor U28838 (N_28838,N_21672,N_24597);
xor U28839 (N_28839,N_24686,N_21758);
nor U28840 (N_28840,N_22977,N_23518);
nand U28841 (N_28841,N_23190,N_20133);
and U28842 (N_28842,N_22253,N_21783);
and U28843 (N_28843,N_23532,N_20729);
nor U28844 (N_28844,N_21728,N_21900);
nor U28845 (N_28845,N_23107,N_24115);
or U28846 (N_28846,N_21500,N_22892);
nor U28847 (N_28847,N_22577,N_23990);
and U28848 (N_28848,N_22482,N_21589);
xor U28849 (N_28849,N_21306,N_20271);
or U28850 (N_28850,N_22961,N_21378);
and U28851 (N_28851,N_22374,N_22702);
and U28852 (N_28852,N_23862,N_21304);
xnor U28853 (N_28853,N_22586,N_23028);
or U28854 (N_28854,N_23259,N_21409);
and U28855 (N_28855,N_23151,N_22115);
or U28856 (N_28856,N_21292,N_22363);
and U28857 (N_28857,N_24766,N_22627);
nor U28858 (N_28858,N_20959,N_23194);
and U28859 (N_28859,N_21097,N_24022);
and U28860 (N_28860,N_20818,N_24631);
or U28861 (N_28861,N_20018,N_22793);
nor U28862 (N_28862,N_22198,N_21179);
nor U28863 (N_28863,N_24315,N_21780);
and U28864 (N_28864,N_20766,N_22489);
or U28865 (N_28865,N_20137,N_21954);
nand U28866 (N_28866,N_21561,N_23191);
nand U28867 (N_28867,N_22731,N_23770);
xor U28868 (N_28868,N_22925,N_24586);
nand U28869 (N_28869,N_21536,N_21041);
nand U28870 (N_28870,N_21859,N_20740);
nor U28871 (N_28871,N_24127,N_23584);
and U28872 (N_28872,N_22337,N_22566);
and U28873 (N_28873,N_22788,N_23681);
nand U28874 (N_28874,N_23302,N_23758);
or U28875 (N_28875,N_20418,N_20970);
nand U28876 (N_28876,N_20212,N_24958);
or U28877 (N_28877,N_20307,N_23363);
or U28878 (N_28878,N_21234,N_23113);
and U28879 (N_28879,N_21678,N_23736);
xnor U28880 (N_28880,N_22726,N_21136);
xor U28881 (N_28881,N_24413,N_20431);
nand U28882 (N_28882,N_23409,N_24835);
xnor U28883 (N_28883,N_22848,N_22095);
xnor U28884 (N_28884,N_22264,N_23876);
xor U28885 (N_28885,N_21763,N_22896);
xnor U28886 (N_28886,N_20342,N_21289);
xor U28887 (N_28887,N_20640,N_24505);
and U28888 (N_28888,N_23649,N_24222);
and U28889 (N_28889,N_22016,N_21253);
nor U28890 (N_28890,N_20416,N_21959);
xor U28891 (N_28891,N_24488,N_20851);
or U28892 (N_28892,N_23780,N_21480);
and U28893 (N_28893,N_22851,N_22237);
or U28894 (N_28894,N_21422,N_23544);
or U28895 (N_28895,N_24241,N_21567);
xnor U28896 (N_28896,N_21756,N_23264);
or U28897 (N_28897,N_24923,N_23834);
nor U28898 (N_28898,N_21705,N_20534);
nor U28899 (N_28899,N_22921,N_24822);
nand U28900 (N_28900,N_23463,N_22642);
xor U28901 (N_28901,N_21777,N_24254);
or U28902 (N_28902,N_21644,N_20409);
xor U28903 (N_28903,N_20059,N_21270);
nor U28904 (N_28904,N_21927,N_22929);
or U28905 (N_28905,N_22078,N_21042);
and U28906 (N_28906,N_24404,N_21286);
xnor U28907 (N_28907,N_20618,N_22492);
nor U28908 (N_28908,N_20867,N_23888);
or U28909 (N_28909,N_21797,N_21448);
or U28910 (N_28910,N_22407,N_21968);
xnor U28911 (N_28911,N_23370,N_23503);
and U28912 (N_28912,N_22371,N_23218);
xnor U28913 (N_28913,N_23339,N_23967);
nand U28914 (N_28914,N_22828,N_21362);
and U28915 (N_28915,N_22870,N_24838);
or U28916 (N_28916,N_21566,N_24539);
nor U28917 (N_28917,N_24303,N_20438);
and U28918 (N_28918,N_24262,N_23368);
nand U28919 (N_28919,N_21563,N_23930);
xnor U28920 (N_28920,N_21837,N_24118);
and U28921 (N_28921,N_21691,N_22439);
nor U28922 (N_28922,N_21293,N_20366);
and U28923 (N_28923,N_24128,N_23444);
nor U28924 (N_28924,N_23787,N_21801);
xor U28925 (N_28925,N_24532,N_23633);
and U28926 (N_28926,N_21471,N_21683);
or U28927 (N_28927,N_24495,N_24589);
nor U28928 (N_28928,N_24001,N_23836);
nand U28929 (N_28929,N_22133,N_20706);
nor U28930 (N_28930,N_20206,N_24155);
or U28931 (N_28931,N_24169,N_24273);
and U28932 (N_28932,N_20192,N_22847);
or U28933 (N_28933,N_23172,N_21254);
or U28934 (N_28934,N_23708,N_23301);
nor U28935 (N_28935,N_22950,N_23542);
xor U28936 (N_28936,N_24013,N_23026);
xor U28937 (N_28937,N_21484,N_22237);
nor U28938 (N_28938,N_22947,N_22497);
or U28939 (N_28939,N_22415,N_20264);
or U28940 (N_28940,N_20091,N_24987);
nor U28941 (N_28941,N_24966,N_20852);
or U28942 (N_28942,N_21798,N_22843);
xor U28943 (N_28943,N_22660,N_23088);
nor U28944 (N_28944,N_21405,N_24486);
xor U28945 (N_28945,N_21254,N_21840);
or U28946 (N_28946,N_22627,N_23359);
or U28947 (N_28947,N_22810,N_21970);
nor U28948 (N_28948,N_23975,N_20966);
xnor U28949 (N_28949,N_21308,N_20055);
nand U28950 (N_28950,N_20706,N_22459);
and U28951 (N_28951,N_20680,N_23549);
and U28952 (N_28952,N_21967,N_23311);
nand U28953 (N_28953,N_24457,N_21966);
and U28954 (N_28954,N_24445,N_23852);
xor U28955 (N_28955,N_23562,N_22706);
nor U28956 (N_28956,N_20668,N_20506);
nand U28957 (N_28957,N_21521,N_22281);
xor U28958 (N_28958,N_23030,N_24123);
and U28959 (N_28959,N_23689,N_22736);
nor U28960 (N_28960,N_22916,N_21929);
nor U28961 (N_28961,N_24786,N_22779);
nand U28962 (N_28962,N_23777,N_23616);
or U28963 (N_28963,N_20913,N_23494);
or U28964 (N_28964,N_20398,N_22785);
xor U28965 (N_28965,N_21303,N_22480);
nor U28966 (N_28966,N_21542,N_21810);
or U28967 (N_28967,N_22018,N_22346);
nor U28968 (N_28968,N_23289,N_22915);
and U28969 (N_28969,N_20407,N_23930);
nand U28970 (N_28970,N_21547,N_23069);
nand U28971 (N_28971,N_20588,N_21521);
xnor U28972 (N_28972,N_23297,N_21528);
and U28973 (N_28973,N_24757,N_22562);
and U28974 (N_28974,N_24162,N_24013);
xnor U28975 (N_28975,N_23573,N_20596);
xnor U28976 (N_28976,N_24417,N_21389);
nor U28977 (N_28977,N_20808,N_21605);
nor U28978 (N_28978,N_22777,N_23130);
nand U28979 (N_28979,N_24569,N_21123);
nand U28980 (N_28980,N_23166,N_21364);
nor U28981 (N_28981,N_23005,N_22702);
xor U28982 (N_28982,N_24475,N_22405);
or U28983 (N_28983,N_24036,N_22582);
and U28984 (N_28984,N_24390,N_24927);
nor U28985 (N_28985,N_23877,N_24215);
xnor U28986 (N_28986,N_20425,N_22910);
or U28987 (N_28987,N_22319,N_20320);
or U28988 (N_28988,N_24821,N_23565);
or U28989 (N_28989,N_21581,N_23196);
nand U28990 (N_28990,N_21138,N_20086);
or U28991 (N_28991,N_22029,N_24385);
nand U28992 (N_28992,N_23728,N_24555);
nor U28993 (N_28993,N_23260,N_24079);
nor U28994 (N_28994,N_21568,N_22497);
and U28995 (N_28995,N_22828,N_23343);
and U28996 (N_28996,N_21302,N_21688);
nor U28997 (N_28997,N_24981,N_20992);
nand U28998 (N_28998,N_24032,N_20513);
and U28999 (N_28999,N_21213,N_21375);
and U29000 (N_29000,N_20775,N_24824);
or U29001 (N_29001,N_23035,N_21423);
nand U29002 (N_29002,N_22487,N_21588);
and U29003 (N_29003,N_21083,N_21675);
or U29004 (N_29004,N_23821,N_23051);
and U29005 (N_29005,N_21779,N_23743);
xor U29006 (N_29006,N_23582,N_22501);
nand U29007 (N_29007,N_24962,N_24301);
and U29008 (N_29008,N_24593,N_23770);
nor U29009 (N_29009,N_21062,N_22659);
nand U29010 (N_29010,N_22097,N_22359);
or U29011 (N_29011,N_21649,N_22688);
nand U29012 (N_29012,N_23044,N_20000);
nor U29013 (N_29013,N_24058,N_20804);
nor U29014 (N_29014,N_21944,N_23456);
xor U29015 (N_29015,N_20456,N_22890);
nor U29016 (N_29016,N_20819,N_24833);
xnor U29017 (N_29017,N_23618,N_24963);
and U29018 (N_29018,N_22387,N_23493);
and U29019 (N_29019,N_23589,N_23543);
nand U29020 (N_29020,N_21450,N_22588);
nand U29021 (N_29021,N_22220,N_20982);
xnor U29022 (N_29022,N_24051,N_24757);
and U29023 (N_29023,N_20156,N_23455);
xnor U29024 (N_29024,N_23731,N_24355);
nor U29025 (N_29025,N_21103,N_23787);
nor U29026 (N_29026,N_23391,N_23015);
or U29027 (N_29027,N_22417,N_24568);
and U29028 (N_29028,N_20947,N_24852);
xnor U29029 (N_29029,N_22199,N_21755);
and U29030 (N_29030,N_23471,N_22621);
and U29031 (N_29031,N_22490,N_22255);
nor U29032 (N_29032,N_23460,N_24984);
nor U29033 (N_29033,N_22089,N_22238);
nand U29034 (N_29034,N_23288,N_21697);
nor U29035 (N_29035,N_20905,N_22866);
and U29036 (N_29036,N_21386,N_20824);
nor U29037 (N_29037,N_23988,N_21328);
nor U29038 (N_29038,N_21867,N_22859);
nor U29039 (N_29039,N_20122,N_22996);
and U29040 (N_29040,N_24800,N_20365);
and U29041 (N_29041,N_23737,N_24730);
and U29042 (N_29042,N_23385,N_22545);
xnor U29043 (N_29043,N_20053,N_24988);
xnor U29044 (N_29044,N_20069,N_24550);
nor U29045 (N_29045,N_20029,N_20937);
and U29046 (N_29046,N_23750,N_20484);
xor U29047 (N_29047,N_23155,N_20532);
nand U29048 (N_29048,N_23929,N_22379);
or U29049 (N_29049,N_22550,N_21146);
and U29050 (N_29050,N_24391,N_24492);
xnor U29051 (N_29051,N_24612,N_24437);
and U29052 (N_29052,N_21845,N_22917);
nor U29053 (N_29053,N_24794,N_21108);
nand U29054 (N_29054,N_23035,N_23555);
xor U29055 (N_29055,N_23013,N_21041);
or U29056 (N_29056,N_23662,N_22058);
xor U29057 (N_29057,N_22129,N_24374);
and U29058 (N_29058,N_24144,N_22784);
and U29059 (N_29059,N_21933,N_20776);
nand U29060 (N_29060,N_20771,N_20711);
or U29061 (N_29061,N_23492,N_24216);
nand U29062 (N_29062,N_22843,N_22999);
nor U29063 (N_29063,N_23197,N_21755);
nand U29064 (N_29064,N_20111,N_20615);
and U29065 (N_29065,N_20242,N_23068);
xor U29066 (N_29066,N_22290,N_22655);
nand U29067 (N_29067,N_23074,N_20223);
or U29068 (N_29068,N_22789,N_22145);
or U29069 (N_29069,N_20889,N_22370);
nor U29070 (N_29070,N_24574,N_20113);
nor U29071 (N_29071,N_20914,N_23800);
nor U29072 (N_29072,N_21239,N_23575);
and U29073 (N_29073,N_23835,N_20193);
and U29074 (N_29074,N_21665,N_21893);
nor U29075 (N_29075,N_22658,N_20889);
and U29076 (N_29076,N_21227,N_24042);
nor U29077 (N_29077,N_22541,N_21620);
nor U29078 (N_29078,N_23109,N_23101);
and U29079 (N_29079,N_23919,N_21859);
and U29080 (N_29080,N_22462,N_23966);
or U29081 (N_29081,N_20976,N_21550);
nand U29082 (N_29082,N_24593,N_20906);
nand U29083 (N_29083,N_22774,N_23493);
xor U29084 (N_29084,N_23814,N_21789);
nor U29085 (N_29085,N_23528,N_22157);
nor U29086 (N_29086,N_20898,N_24344);
nor U29087 (N_29087,N_23598,N_20173);
nor U29088 (N_29088,N_20718,N_21526);
or U29089 (N_29089,N_24882,N_22006);
nand U29090 (N_29090,N_23902,N_24669);
and U29091 (N_29091,N_23624,N_24459);
and U29092 (N_29092,N_21794,N_23394);
nor U29093 (N_29093,N_22849,N_21256);
nor U29094 (N_29094,N_24680,N_20550);
and U29095 (N_29095,N_20786,N_22163);
or U29096 (N_29096,N_23919,N_23376);
xor U29097 (N_29097,N_20899,N_23889);
or U29098 (N_29098,N_22168,N_22013);
or U29099 (N_29099,N_20822,N_23485);
nor U29100 (N_29100,N_22721,N_21800);
nand U29101 (N_29101,N_23186,N_24236);
and U29102 (N_29102,N_22007,N_20838);
nand U29103 (N_29103,N_23900,N_20311);
or U29104 (N_29104,N_24074,N_21719);
xor U29105 (N_29105,N_20592,N_24921);
nand U29106 (N_29106,N_23928,N_20829);
xnor U29107 (N_29107,N_22392,N_22555);
xor U29108 (N_29108,N_20345,N_20128);
nor U29109 (N_29109,N_23524,N_24844);
and U29110 (N_29110,N_24035,N_21234);
nand U29111 (N_29111,N_21144,N_21063);
or U29112 (N_29112,N_20662,N_24210);
and U29113 (N_29113,N_23249,N_20992);
nor U29114 (N_29114,N_24347,N_24480);
and U29115 (N_29115,N_20129,N_23157);
nand U29116 (N_29116,N_24090,N_24177);
nand U29117 (N_29117,N_24438,N_23440);
or U29118 (N_29118,N_20859,N_21738);
xnor U29119 (N_29119,N_22032,N_22634);
xor U29120 (N_29120,N_22558,N_24317);
nand U29121 (N_29121,N_24188,N_20782);
or U29122 (N_29122,N_22808,N_21211);
or U29123 (N_29123,N_22264,N_23226);
xnor U29124 (N_29124,N_22222,N_20186);
nand U29125 (N_29125,N_21261,N_22947);
nand U29126 (N_29126,N_22562,N_20017);
or U29127 (N_29127,N_22384,N_21133);
nor U29128 (N_29128,N_20785,N_21477);
or U29129 (N_29129,N_20611,N_23376);
nand U29130 (N_29130,N_24848,N_20950);
or U29131 (N_29131,N_21268,N_20129);
and U29132 (N_29132,N_23589,N_20766);
or U29133 (N_29133,N_21120,N_24820);
nand U29134 (N_29134,N_21780,N_23326);
nor U29135 (N_29135,N_20564,N_24526);
and U29136 (N_29136,N_23334,N_24564);
nand U29137 (N_29137,N_24896,N_20634);
and U29138 (N_29138,N_21328,N_24957);
or U29139 (N_29139,N_24681,N_24057);
xor U29140 (N_29140,N_24928,N_20907);
nor U29141 (N_29141,N_24709,N_22149);
or U29142 (N_29142,N_23724,N_23589);
nor U29143 (N_29143,N_23860,N_22535);
or U29144 (N_29144,N_22254,N_21311);
xnor U29145 (N_29145,N_22668,N_24789);
xnor U29146 (N_29146,N_21848,N_24095);
xnor U29147 (N_29147,N_24553,N_21121);
or U29148 (N_29148,N_22626,N_21143);
or U29149 (N_29149,N_24615,N_24704);
xor U29150 (N_29150,N_21093,N_24444);
and U29151 (N_29151,N_21040,N_22028);
nand U29152 (N_29152,N_21906,N_21673);
and U29153 (N_29153,N_24907,N_20186);
xnor U29154 (N_29154,N_20101,N_22434);
or U29155 (N_29155,N_21677,N_24230);
and U29156 (N_29156,N_23080,N_21664);
nor U29157 (N_29157,N_24560,N_21947);
xnor U29158 (N_29158,N_20421,N_23773);
xor U29159 (N_29159,N_22610,N_21831);
nand U29160 (N_29160,N_24889,N_21846);
and U29161 (N_29161,N_21020,N_24755);
or U29162 (N_29162,N_24145,N_24852);
xor U29163 (N_29163,N_24594,N_23940);
nor U29164 (N_29164,N_21527,N_23556);
xnor U29165 (N_29165,N_23531,N_23389);
nor U29166 (N_29166,N_23196,N_21146);
or U29167 (N_29167,N_21295,N_21852);
nand U29168 (N_29168,N_21211,N_24592);
nor U29169 (N_29169,N_24912,N_23885);
and U29170 (N_29170,N_22174,N_23037);
and U29171 (N_29171,N_22215,N_21225);
xnor U29172 (N_29172,N_22065,N_22919);
nor U29173 (N_29173,N_24315,N_20510);
or U29174 (N_29174,N_21298,N_23984);
or U29175 (N_29175,N_21562,N_24332);
nand U29176 (N_29176,N_20843,N_23517);
nand U29177 (N_29177,N_24732,N_22626);
nand U29178 (N_29178,N_24660,N_20993);
nand U29179 (N_29179,N_22745,N_22266);
or U29180 (N_29180,N_21041,N_20705);
or U29181 (N_29181,N_22743,N_22435);
nand U29182 (N_29182,N_24541,N_20630);
nor U29183 (N_29183,N_22641,N_22661);
or U29184 (N_29184,N_20040,N_21725);
or U29185 (N_29185,N_21062,N_21031);
nand U29186 (N_29186,N_22412,N_21687);
nor U29187 (N_29187,N_21575,N_20720);
nand U29188 (N_29188,N_20349,N_20932);
nor U29189 (N_29189,N_22157,N_21763);
and U29190 (N_29190,N_22815,N_20239);
nand U29191 (N_29191,N_23569,N_21248);
xor U29192 (N_29192,N_24692,N_21216);
nor U29193 (N_29193,N_23802,N_23063);
nand U29194 (N_29194,N_24057,N_21735);
or U29195 (N_29195,N_24756,N_21156);
or U29196 (N_29196,N_21276,N_20997);
xor U29197 (N_29197,N_21232,N_21204);
nor U29198 (N_29198,N_20353,N_21460);
or U29199 (N_29199,N_20123,N_24616);
and U29200 (N_29200,N_24000,N_20840);
and U29201 (N_29201,N_23609,N_21582);
nand U29202 (N_29202,N_20000,N_23614);
nand U29203 (N_29203,N_24069,N_22524);
nand U29204 (N_29204,N_24687,N_22015);
and U29205 (N_29205,N_21457,N_24720);
and U29206 (N_29206,N_24106,N_22701);
nand U29207 (N_29207,N_23561,N_21039);
xnor U29208 (N_29208,N_23768,N_22770);
nand U29209 (N_29209,N_22105,N_22627);
nand U29210 (N_29210,N_24171,N_22863);
or U29211 (N_29211,N_23619,N_24143);
nor U29212 (N_29212,N_20302,N_22397);
or U29213 (N_29213,N_20109,N_23932);
xnor U29214 (N_29214,N_22627,N_22242);
or U29215 (N_29215,N_20353,N_23372);
and U29216 (N_29216,N_21948,N_20539);
nand U29217 (N_29217,N_24941,N_20344);
nand U29218 (N_29218,N_20562,N_24426);
xnor U29219 (N_29219,N_24497,N_21479);
nand U29220 (N_29220,N_20715,N_22914);
xnor U29221 (N_29221,N_22746,N_21823);
nor U29222 (N_29222,N_22696,N_24200);
nor U29223 (N_29223,N_20103,N_24115);
nor U29224 (N_29224,N_24728,N_20286);
and U29225 (N_29225,N_23551,N_23774);
and U29226 (N_29226,N_22939,N_22272);
nand U29227 (N_29227,N_23880,N_23998);
or U29228 (N_29228,N_22340,N_22777);
nand U29229 (N_29229,N_23186,N_24144);
and U29230 (N_29230,N_21150,N_20615);
xnor U29231 (N_29231,N_21321,N_20051);
and U29232 (N_29232,N_24334,N_22083);
xor U29233 (N_29233,N_21588,N_24675);
nor U29234 (N_29234,N_20033,N_22759);
nand U29235 (N_29235,N_24634,N_24548);
or U29236 (N_29236,N_22594,N_23758);
nand U29237 (N_29237,N_24630,N_22280);
nand U29238 (N_29238,N_22075,N_22062);
or U29239 (N_29239,N_23930,N_23318);
xor U29240 (N_29240,N_23413,N_20638);
nand U29241 (N_29241,N_24552,N_23787);
xor U29242 (N_29242,N_23232,N_24787);
nand U29243 (N_29243,N_20699,N_22786);
xnor U29244 (N_29244,N_20178,N_21074);
xnor U29245 (N_29245,N_20811,N_20193);
and U29246 (N_29246,N_20079,N_20521);
nand U29247 (N_29247,N_20698,N_20164);
nand U29248 (N_29248,N_22111,N_20784);
and U29249 (N_29249,N_24391,N_22332);
or U29250 (N_29250,N_20736,N_23837);
nor U29251 (N_29251,N_23179,N_20482);
and U29252 (N_29252,N_24924,N_23392);
nor U29253 (N_29253,N_24237,N_21778);
or U29254 (N_29254,N_20743,N_21168);
xor U29255 (N_29255,N_23654,N_24160);
nor U29256 (N_29256,N_24046,N_22618);
xor U29257 (N_29257,N_22170,N_22785);
nor U29258 (N_29258,N_23421,N_22276);
or U29259 (N_29259,N_23756,N_20628);
or U29260 (N_29260,N_22745,N_24728);
nor U29261 (N_29261,N_24462,N_22661);
and U29262 (N_29262,N_21350,N_21359);
or U29263 (N_29263,N_22638,N_21105);
xnor U29264 (N_29264,N_22064,N_20484);
xnor U29265 (N_29265,N_21945,N_24858);
nor U29266 (N_29266,N_21783,N_24332);
and U29267 (N_29267,N_23735,N_23470);
or U29268 (N_29268,N_23139,N_20575);
nand U29269 (N_29269,N_23071,N_21663);
nor U29270 (N_29270,N_22321,N_23836);
and U29271 (N_29271,N_22712,N_20593);
nand U29272 (N_29272,N_22319,N_20738);
or U29273 (N_29273,N_22650,N_24047);
or U29274 (N_29274,N_20740,N_24552);
nor U29275 (N_29275,N_24421,N_20256);
and U29276 (N_29276,N_24574,N_24918);
or U29277 (N_29277,N_24672,N_22527);
xor U29278 (N_29278,N_24370,N_22619);
and U29279 (N_29279,N_21914,N_21179);
nor U29280 (N_29280,N_21446,N_21882);
and U29281 (N_29281,N_24310,N_22021);
xor U29282 (N_29282,N_23564,N_21662);
and U29283 (N_29283,N_23659,N_20167);
and U29284 (N_29284,N_21781,N_24516);
nor U29285 (N_29285,N_22753,N_24450);
xnor U29286 (N_29286,N_23776,N_21571);
nor U29287 (N_29287,N_20929,N_22655);
or U29288 (N_29288,N_22014,N_20738);
xnor U29289 (N_29289,N_22552,N_24019);
or U29290 (N_29290,N_22411,N_23286);
or U29291 (N_29291,N_23066,N_22880);
and U29292 (N_29292,N_23544,N_24827);
nand U29293 (N_29293,N_22491,N_24843);
nor U29294 (N_29294,N_22847,N_23595);
nor U29295 (N_29295,N_20986,N_23436);
xnor U29296 (N_29296,N_20355,N_22948);
xor U29297 (N_29297,N_21015,N_20690);
and U29298 (N_29298,N_23976,N_20906);
and U29299 (N_29299,N_24553,N_22709);
nand U29300 (N_29300,N_22835,N_23564);
nand U29301 (N_29301,N_22961,N_22259);
or U29302 (N_29302,N_20354,N_20274);
nor U29303 (N_29303,N_24091,N_20050);
nor U29304 (N_29304,N_24442,N_22335);
and U29305 (N_29305,N_21586,N_23741);
xnor U29306 (N_29306,N_22983,N_21796);
nand U29307 (N_29307,N_20113,N_20809);
and U29308 (N_29308,N_23832,N_21746);
and U29309 (N_29309,N_23691,N_20036);
or U29310 (N_29310,N_20004,N_21012);
nand U29311 (N_29311,N_22919,N_22984);
and U29312 (N_29312,N_21961,N_22250);
nor U29313 (N_29313,N_23364,N_24362);
and U29314 (N_29314,N_24612,N_24126);
nand U29315 (N_29315,N_23272,N_20878);
and U29316 (N_29316,N_22385,N_23663);
nor U29317 (N_29317,N_22253,N_20437);
or U29318 (N_29318,N_22750,N_24224);
or U29319 (N_29319,N_21809,N_20465);
nor U29320 (N_29320,N_20982,N_21646);
and U29321 (N_29321,N_20402,N_22324);
nor U29322 (N_29322,N_20251,N_20256);
and U29323 (N_29323,N_20214,N_21738);
or U29324 (N_29324,N_24668,N_21899);
nor U29325 (N_29325,N_23111,N_20785);
nand U29326 (N_29326,N_22690,N_21938);
nand U29327 (N_29327,N_24884,N_23795);
xnor U29328 (N_29328,N_21341,N_24621);
nor U29329 (N_29329,N_23438,N_22522);
and U29330 (N_29330,N_24034,N_23170);
and U29331 (N_29331,N_20107,N_23349);
nor U29332 (N_29332,N_23695,N_22053);
nand U29333 (N_29333,N_23299,N_23858);
or U29334 (N_29334,N_23405,N_22555);
xor U29335 (N_29335,N_24607,N_24328);
or U29336 (N_29336,N_21141,N_24205);
nor U29337 (N_29337,N_24754,N_20403);
nor U29338 (N_29338,N_23669,N_24969);
or U29339 (N_29339,N_24336,N_23772);
and U29340 (N_29340,N_21828,N_24287);
and U29341 (N_29341,N_23011,N_20088);
or U29342 (N_29342,N_23997,N_24607);
xor U29343 (N_29343,N_23412,N_24153);
xnor U29344 (N_29344,N_23479,N_21693);
or U29345 (N_29345,N_24159,N_21878);
xor U29346 (N_29346,N_20411,N_21095);
xor U29347 (N_29347,N_21603,N_20643);
nor U29348 (N_29348,N_20700,N_22333);
or U29349 (N_29349,N_21586,N_24740);
nor U29350 (N_29350,N_23720,N_21680);
nand U29351 (N_29351,N_22595,N_24352);
nand U29352 (N_29352,N_20805,N_22040);
nor U29353 (N_29353,N_22682,N_24278);
and U29354 (N_29354,N_20847,N_20184);
nand U29355 (N_29355,N_20269,N_23970);
and U29356 (N_29356,N_20388,N_23171);
nor U29357 (N_29357,N_22813,N_20000);
nor U29358 (N_29358,N_22871,N_23424);
and U29359 (N_29359,N_20798,N_20317);
nor U29360 (N_29360,N_22020,N_24809);
xnor U29361 (N_29361,N_23061,N_20178);
xor U29362 (N_29362,N_21559,N_24244);
or U29363 (N_29363,N_24917,N_24280);
nand U29364 (N_29364,N_22483,N_20700);
nand U29365 (N_29365,N_24786,N_21572);
or U29366 (N_29366,N_21035,N_23710);
and U29367 (N_29367,N_21025,N_23737);
xor U29368 (N_29368,N_24095,N_23900);
nor U29369 (N_29369,N_24695,N_24457);
or U29370 (N_29370,N_22327,N_23540);
xnor U29371 (N_29371,N_24665,N_23149);
xor U29372 (N_29372,N_24865,N_21007);
and U29373 (N_29373,N_24266,N_23793);
nand U29374 (N_29374,N_21555,N_24625);
nor U29375 (N_29375,N_23282,N_20560);
and U29376 (N_29376,N_22381,N_22175);
xor U29377 (N_29377,N_20907,N_20719);
nor U29378 (N_29378,N_24055,N_23510);
and U29379 (N_29379,N_20088,N_21340);
and U29380 (N_29380,N_22443,N_23855);
nand U29381 (N_29381,N_23917,N_23518);
xor U29382 (N_29382,N_21082,N_21590);
and U29383 (N_29383,N_23998,N_21759);
nor U29384 (N_29384,N_22063,N_21469);
nand U29385 (N_29385,N_22340,N_20972);
or U29386 (N_29386,N_20793,N_23121);
or U29387 (N_29387,N_21412,N_20510);
and U29388 (N_29388,N_22658,N_21355);
nand U29389 (N_29389,N_21005,N_20597);
and U29390 (N_29390,N_20294,N_22447);
xnor U29391 (N_29391,N_22578,N_24051);
nor U29392 (N_29392,N_22134,N_21940);
nor U29393 (N_29393,N_24231,N_21734);
nand U29394 (N_29394,N_23979,N_24034);
and U29395 (N_29395,N_21127,N_20943);
or U29396 (N_29396,N_20525,N_24266);
nor U29397 (N_29397,N_20440,N_20768);
or U29398 (N_29398,N_22574,N_22476);
nand U29399 (N_29399,N_20840,N_24937);
xor U29400 (N_29400,N_21578,N_23840);
xnor U29401 (N_29401,N_24472,N_21804);
nor U29402 (N_29402,N_20313,N_22210);
xor U29403 (N_29403,N_22451,N_24503);
or U29404 (N_29404,N_21069,N_22211);
and U29405 (N_29405,N_20702,N_21966);
xnor U29406 (N_29406,N_20937,N_21882);
nor U29407 (N_29407,N_22704,N_21871);
xnor U29408 (N_29408,N_24820,N_21680);
and U29409 (N_29409,N_22170,N_24552);
nor U29410 (N_29410,N_22580,N_21946);
xnor U29411 (N_29411,N_21373,N_24611);
and U29412 (N_29412,N_24866,N_23252);
nand U29413 (N_29413,N_22230,N_23753);
nand U29414 (N_29414,N_20633,N_24609);
nand U29415 (N_29415,N_20694,N_22214);
nand U29416 (N_29416,N_24046,N_23813);
nand U29417 (N_29417,N_24261,N_21034);
and U29418 (N_29418,N_22350,N_24781);
xor U29419 (N_29419,N_21799,N_20432);
nand U29420 (N_29420,N_20263,N_24260);
nor U29421 (N_29421,N_21064,N_21182);
xnor U29422 (N_29422,N_20917,N_21333);
xor U29423 (N_29423,N_23215,N_24175);
nand U29424 (N_29424,N_21489,N_20472);
or U29425 (N_29425,N_22790,N_21350);
and U29426 (N_29426,N_23602,N_24640);
or U29427 (N_29427,N_23038,N_22328);
nor U29428 (N_29428,N_22452,N_20146);
nand U29429 (N_29429,N_22657,N_22972);
and U29430 (N_29430,N_20952,N_20102);
or U29431 (N_29431,N_23754,N_24869);
xnor U29432 (N_29432,N_22035,N_22926);
and U29433 (N_29433,N_21835,N_22032);
xor U29434 (N_29434,N_22974,N_23932);
and U29435 (N_29435,N_23099,N_22384);
xnor U29436 (N_29436,N_23473,N_21537);
or U29437 (N_29437,N_23917,N_24774);
nor U29438 (N_29438,N_20222,N_23242);
and U29439 (N_29439,N_23070,N_22424);
nand U29440 (N_29440,N_24172,N_22822);
nor U29441 (N_29441,N_20067,N_24702);
or U29442 (N_29442,N_22553,N_22081);
xor U29443 (N_29443,N_23422,N_20722);
nand U29444 (N_29444,N_23031,N_23192);
or U29445 (N_29445,N_22331,N_20645);
or U29446 (N_29446,N_23576,N_21630);
nor U29447 (N_29447,N_22548,N_20077);
or U29448 (N_29448,N_23744,N_21461);
xnor U29449 (N_29449,N_21725,N_20277);
nor U29450 (N_29450,N_22866,N_21823);
xor U29451 (N_29451,N_23932,N_20607);
or U29452 (N_29452,N_24942,N_23516);
xnor U29453 (N_29453,N_22020,N_20140);
nor U29454 (N_29454,N_20803,N_20464);
nand U29455 (N_29455,N_20705,N_24453);
or U29456 (N_29456,N_24745,N_22999);
and U29457 (N_29457,N_23640,N_20442);
and U29458 (N_29458,N_24818,N_22295);
or U29459 (N_29459,N_23801,N_23470);
and U29460 (N_29460,N_21932,N_20425);
xor U29461 (N_29461,N_22729,N_21145);
nand U29462 (N_29462,N_21699,N_20197);
and U29463 (N_29463,N_24859,N_20568);
nand U29464 (N_29464,N_24197,N_23645);
nand U29465 (N_29465,N_22186,N_24287);
and U29466 (N_29466,N_24984,N_20992);
and U29467 (N_29467,N_24219,N_20828);
nand U29468 (N_29468,N_20305,N_23400);
nand U29469 (N_29469,N_24313,N_21053);
nor U29470 (N_29470,N_23474,N_20500);
xnor U29471 (N_29471,N_22731,N_20385);
and U29472 (N_29472,N_21602,N_23097);
or U29473 (N_29473,N_23013,N_23022);
or U29474 (N_29474,N_24852,N_23675);
nand U29475 (N_29475,N_22848,N_23828);
or U29476 (N_29476,N_22216,N_21117);
or U29477 (N_29477,N_20435,N_20549);
nand U29478 (N_29478,N_24006,N_23045);
nand U29479 (N_29479,N_21293,N_21775);
and U29480 (N_29480,N_21061,N_22905);
nor U29481 (N_29481,N_22104,N_24267);
and U29482 (N_29482,N_24803,N_22614);
nor U29483 (N_29483,N_23222,N_22308);
and U29484 (N_29484,N_21323,N_24149);
nand U29485 (N_29485,N_20672,N_23436);
nand U29486 (N_29486,N_24021,N_24822);
nor U29487 (N_29487,N_24880,N_20413);
and U29488 (N_29488,N_22606,N_24039);
nand U29489 (N_29489,N_22152,N_21981);
nand U29490 (N_29490,N_21392,N_21801);
or U29491 (N_29491,N_21721,N_22542);
nor U29492 (N_29492,N_21328,N_22394);
nand U29493 (N_29493,N_24090,N_20587);
nand U29494 (N_29494,N_20077,N_24957);
nand U29495 (N_29495,N_20509,N_22118);
nor U29496 (N_29496,N_24061,N_20680);
nor U29497 (N_29497,N_21807,N_20136);
xnor U29498 (N_29498,N_21396,N_23428);
nand U29499 (N_29499,N_20794,N_24090);
and U29500 (N_29500,N_23341,N_20291);
or U29501 (N_29501,N_22643,N_23639);
or U29502 (N_29502,N_20979,N_24934);
nand U29503 (N_29503,N_24152,N_21388);
or U29504 (N_29504,N_21560,N_20374);
and U29505 (N_29505,N_20127,N_20195);
nor U29506 (N_29506,N_21610,N_21810);
nor U29507 (N_29507,N_20747,N_22485);
nor U29508 (N_29508,N_21008,N_20508);
xnor U29509 (N_29509,N_21723,N_20911);
or U29510 (N_29510,N_23810,N_22120);
or U29511 (N_29511,N_20139,N_24740);
nor U29512 (N_29512,N_23162,N_24475);
nand U29513 (N_29513,N_24104,N_24462);
xor U29514 (N_29514,N_24008,N_22451);
xor U29515 (N_29515,N_24514,N_22658);
nand U29516 (N_29516,N_22416,N_20672);
nor U29517 (N_29517,N_24068,N_24631);
nor U29518 (N_29518,N_21025,N_23605);
and U29519 (N_29519,N_20832,N_22210);
or U29520 (N_29520,N_24452,N_24856);
nor U29521 (N_29521,N_24753,N_23271);
nand U29522 (N_29522,N_22175,N_20048);
or U29523 (N_29523,N_21550,N_20619);
nand U29524 (N_29524,N_20003,N_23186);
and U29525 (N_29525,N_23941,N_20121);
and U29526 (N_29526,N_20296,N_23952);
nor U29527 (N_29527,N_22826,N_22882);
or U29528 (N_29528,N_22860,N_23983);
nor U29529 (N_29529,N_20814,N_20881);
nor U29530 (N_29530,N_20001,N_21019);
or U29531 (N_29531,N_22882,N_24592);
and U29532 (N_29532,N_24640,N_23339);
or U29533 (N_29533,N_20371,N_22918);
nor U29534 (N_29534,N_24949,N_20230);
nor U29535 (N_29535,N_24408,N_20670);
xnor U29536 (N_29536,N_24921,N_22337);
or U29537 (N_29537,N_22404,N_24971);
nor U29538 (N_29538,N_21402,N_21758);
xor U29539 (N_29539,N_21636,N_21204);
nor U29540 (N_29540,N_20996,N_20847);
or U29541 (N_29541,N_22509,N_21208);
nand U29542 (N_29542,N_22882,N_23539);
nand U29543 (N_29543,N_24165,N_24052);
and U29544 (N_29544,N_24917,N_21571);
nor U29545 (N_29545,N_20311,N_24864);
or U29546 (N_29546,N_21177,N_24878);
nand U29547 (N_29547,N_21219,N_23042);
nor U29548 (N_29548,N_20168,N_24695);
and U29549 (N_29549,N_21436,N_20292);
nand U29550 (N_29550,N_23277,N_23552);
and U29551 (N_29551,N_22332,N_24309);
or U29552 (N_29552,N_20870,N_24527);
nand U29553 (N_29553,N_24764,N_20921);
nor U29554 (N_29554,N_23268,N_21693);
or U29555 (N_29555,N_23545,N_20756);
or U29556 (N_29556,N_23825,N_22359);
and U29557 (N_29557,N_20648,N_20194);
and U29558 (N_29558,N_23169,N_21025);
or U29559 (N_29559,N_22699,N_22828);
or U29560 (N_29560,N_24244,N_24008);
xor U29561 (N_29561,N_23032,N_24017);
or U29562 (N_29562,N_23574,N_20702);
xnor U29563 (N_29563,N_23132,N_22376);
nor U29564 (N_29564,N_23106,N_23130);
and U29565 (N_29565,N_21950,N_21832);
nor U29566 (N_29566,N_22373,N_22940);
xnor U29567 (N_29567,N_24692,N_20120);
or U29568 (N_29568,N_23182,N_21177);
nor U29569 (N_29569,N_22140,N_20924);
xor U29570 (N_29570,N_24202,N_24639);
or U29571 (N_29571,N_24132,N_22612);
nand U29572 (N_29572,N_20891,N_21864);
nor U29573 (N_29573,N_22906,N_20693);
xor U29574 (N_29574,N_22886,N_24589);
and U29575 (N_29575,N_24291,N_24425);
nand U29576 (N_29576,N_24690,N_21991);
xnor U29577 (N_29577,N_22173,N_24409);
and U29578 (N_29578,N_21240,N_20586);
xor U29579 (N_29579,N_20225,N_23157);
nand U29580 (N_29580,N_21319,N_21566);
nor U29581 (N_29581,N_20075,N_24965);
nor U29582 (N_29582,N_22489,N_20950);
nor U29583 (N_29583,N_23780,N_20860);
and U29584 (N_29584,N_21083,N_20955);
or U29585 (N_29585,N_24051,N_21996);
xor U29586 (N_29586,N_22102,N_22872);
xor U29587 (N_29587,N_23386,N_20734);
nand U29588 (N_29588,N_22186,N_23784);
nand U29589 (N_29589,N_24402,N_22094);
or U29590 (N_29590,N_20551,N_20353);
or U29591 (N_29591,N_22713,N_21060);
nor U29592 (N_29592,N_22236,N_21398);
nand U29593 (N_29593,N_24805,N_22797);
and U29594 (N_29594,N_24145,N_20966);
nor U29595 (N_29595,N_23309,N_20242);
xnor U29596 (N_29596,N_20204,N_24932);
xnor U29597 (N_29597,N_21351,N_22716);
nand U29598 (N_29598,N_21290,N_23064);
nor U29599 (N_29599,N_21111,N_23402);
or U29600 (N_29600,N_24368,N_24154);
nand U29601 (N_29601,N_24938,N_22460);
xor U29602 (N_29602,N_24638,N_23309);
nand U29603 (N_29603,N_24422,N_21553);
and U29604 (N_29604,N_22304,N_23844);
or U29605 (N_29605,N_20428,N_23577);
nand U29606 (N_29606,N_24053,N_22090);
nor U29607 (N_29607,N_21464,N_22191);
or U29608 (N_29608,N_24240,N_22463);
xnor U29609 (N_29609,N_21501,N_23889);
nor U29610 (N_29610,N_23904,N_20878);
and U29611 (N_29611,N_21284,N_22030);
nor U29612 (N_29612,N_20997,N_21954);
nand U29613 (N_29613,N_24295,N_20853);
xor U29614 (N_29614,N_22622,N_22425);
nor U29615 (N_29615,N_21243,N_24978);
and U29616 (N_29616,N_23378,N_20295);
xor U29617 (N_29617,N_23806,N_21529);
xnor U29618 (N_29618,N_20495,N_23140);
and U29619 (N_29619,N_23257,N_23540);
and U29620 (N_29620,N_23449,N_21428);
xnor U29621 (N_29621,N_20743,N_24377);
nand U29622 (N_29622,N_22709,N_23402);
xor U29623 (N_29623,N_21637,N_24700);
nor U29624 (N_29624,N_23438,N_23049);
or U29625 (N_29625,N_24681,N_24755);
xnor U29626 (N_29626,N_21085,N_23136);
xor U29627 (N_29627,N_21975,N_22523);
nor U29628 (N_29628,N_24688,N_22585);
and U29629 (N_29629,N_20926,N_20405);
and U29630 (N_29630,N_23838,N_22429);
or U29631 (N_29631,N_20548,N_24900);
and U29632 (N_29632,N_24148,N_23561);
xnor U29633 (N_29633,N_21727,N_20921);
nand U29634 (N_29634,N_23110,N_22934);
or U29635 (N_29635,N_24376,N_22999);
xnor U29636 (N_29636,N_20931,N_22413);
or U29637 (N_29637,N_24460,N_23185);
or U29638 (N_29638,N_21017,N_20266);
nand U29639 (N_29639,N_22068,N_22492);
nor U29640 (N_29640,N_21000,N_20320);
nand U29641 (N_29641,N_21898,N_22655);
or U29642 (N_29642,N_20311,N_20582);
nor U29643 (N_29643,N_24717,N_22665);
xor U29644 (N_29644,N_22817,N_21695);
nand U29645 (N_29645,N_23534,N_20013);
or U29646 (N_29646,N_24699,N_23938);
and U29647 (N_29647,N_22025,N_23597);
and U29648 (N_29648,N_24896,N_21895);
or U29649 (N_29649,N_21174,N_23745);
or U29650 (N_29650,N_20750,N_21916);
or U29651 (N_29651,N_24241,N_23792);
nor U29652 (N_29652,N_22294,N_24240);
or U29653 (N_29653,N_20116,N_20654);
nand U29654 (N_29654,N_21102,N_22799);
and U29655 (N_29655,N_24683,N_24606);
nand U29656 (N_29656,N_22882,N_23339);
nand U29657 (N_29657,N_20288,N_20697);
nand U29658 (N_29658,N_20678,N_20915);
nor U29659 (N_29659,N_22220,N_20625);
xor U29660 (N_29660,N_22727,N_23475);
and U29661 (N_29661,N_20905,N_20057);
nand U29662 (N_29662,N_23085,N_24048);
nand U29663 (N_29663,N_20726,N_24271);
xor U29664 (N_29664,N_20900,N_23260);
xnor U29665 (N_29665,N_21283,N_23466);
xor U29666 (N_29666,N_21579,N_20376);
nor U29667 (N_29667,N_23741,N_22669);
nand U29668 (N_29668,N_20371,N_22471);
and U29669 (N_29669,N_23535,N_23238);
nand U29670 (N_29670,N_22411,N_20040);
xnor U29671 (N_29671,N_24776,N_24091);
nand U29672 (N_29672,N_21107,N_23937);
or U29673 (N_29673,N_24885,N_21840);
xor U29674 (N_29674,N_24999,N_21558);
xnor U29675 (N_29675,N_21717,N_23039);
xnor U29676 (N_29676,N_22800,N_24339);
xnor U29677 (N_29677,N_21578,N_20401);
nand U29678 (N_29678,N_20699,N_21138);
nor U29679 (N_29679,N_20985,N_23497);
and U29680 (N_29680,N_21857,N_24091);
xor U29681 (N_29681,N_20358,N_21010);
or U29682 (N_29682,N_21188,N_22722);
nor U29683 (N_29683,N_24319,N_20058);
xor U29684 (N_29684,N_20762,N_21007);
or U29685 (N_29685,N_22000,N_21135);
nor U29686 (N_29686,N_23736,N_20800);
nor U29687 (N_29687,N_20954,N_24588);
and U29688 (N_29688,N_21731,N_21594);
xnor U29689 (N_29689,N_24562,N_21382);
nor U29690 (N_29690,N_24453,N_23464);
xor U29691 (N_29691,N_22652,N_23646);
xnor U29692 (N_29692,N_21669,N_24449);
and U29693 (N_29693,N_20094,N_24653);
nor U29694 (N_29694,N_23113,N_24868);
xnor U29695 (N_29695,N_22136,N_22168);
or U29696 (N_29696,N_22305,N_21436);
and U29697 (N_29697,N_21424,N_24751);
or U29698 (N_29698,N_20418,N_22953);
nor U29699 (N_29699,N_21206,N_24733);
xor U29700 (N_29700,N_24571,N_21798);
or U29701 (N_29701,N_20109,N_21704);
or U29702 (N_29702,N_21669,N_21517);
or U29703 (N_29703,N_21784,N_20291);
or U29704 (N_29704,N_22756,N_20269);
nor U29705 (N_29705,N_20391,N_21596);
nand U29706 (N_29706,N_23900,N_24231);
and U29707 (N_29707,N_23888,N_20342);
and U29708 (N_29708,N_21239,N_20299);
or U29709 (N_29709,N_21948,N_24845);
nand U29710 (N_29710,N_23091,N_22754);
xor U29711 (N_29711,N_21748,N_20684);
xnor U29712 (N_29712,N_21736,N_22585);
or U29713 (N_29713,N_22551,N_24701);
nor U29714 (N_29714,N_22505,N_22204);
nand U29715 (N_29715,N_22919,N_23702);
and U29716 (N_29716,N_23844,N_24305);
xor U29717 (N_29717,N_23657,N_21030);
nand U29718 (N_29718,N_23169,N_20731);
nor U29719 (N_29719,N_23693,N_22556);
and U29720 (N_29720,N_21318,N_22469);
and U29721 (N_29721,N_22436,N_22274);
or U29722 (N_29722,N_24250,N_24323);
and U29723 (N_29723,N_24767,N_23281);
or U29724 (N_29724,N_21184,N_21484);
and U29725 (N_29725,N_24821,N_23280);
or U29726 (N_29726,N_24722,N_21586);
and U29727 (N_29727,N_23903,N_20854);
xnor U29728 (N_29728,N_22109,N_22799);
or U29729 (N_29729,N_20185,N_22700);
and U29730 (N_29730,N_21958,N_24911);
and U29731 (N_29731,N_21273,N_20757);
and U29732 (N_29732,N_21697,N_24765);
nand U29733 (N_29733,N_24512,N_23956);
or U29734 (N_29734,N_20390,N_24141);
and U29735 (N_29735,N_21233,N_24030);
or U29736 (N_29736,N_24308,N_23554);
and U29737 (N_29737,N_24443,N_21292);
nand U29738 (N_29738,N_20871,N_20421);
nor U29739 (N_29739,N_23956,N_22103);
or U29740 (N_29740,N_22878,N_24916);
and U29741 (N_29741,N_22422,N_22349);
nand U29742 (N_29742,N_24545,N_23934);
and U29743 (N_29743,N_20600,N_22991);
xor U29744 (N_29744,N_21172,N_24454);
and U29745 (N_29745,N_20499,N_24569);
xor U29746 (N_29746,N_24843,N_21263);
and U29747 (N_29747,N_21534,N_21335);
nand U29748 (N_29748,N_23574,N_22414);
xor U29749 (N_29749,N_24057,N_24977);
nor U29750 (N_29750,N_24841,N_21181);
or U29751 (N_29751,N_23688,N_22962);
and U29752 (N_29752,N_21981,N_20837);
and U29753 (N_29753,N_23363,N_24176);
nor U29754 (N_29754,N_22700,N_24243);
nand U29755 (N_29755,N_22352,N_22266);
xnor U29756 (N_29756,N_24622,N_23365);
or U29757 (N_29757,N_23641,N_20399);
xnor U29758 (N_29758,N_24323,N_22495);
or U29759 (N_29759,N_22468,N_21192);
nor U29760 (N_29760,N_20530,N_22662);
xor U29761 (N_29761,N_23411,N_21462);
or U29762 (N_29762,N_24166,N_20663);
nor U29763 (N_29763,N_22442,N_21619);
and U29764 (N_29764,N_24135,N_24100);
xor U29765 (N_29765,N_22351,N_21563);
nor U29766 (N_29766,N_24470,N_24962);
or U29767 (N_29767,N_24654,N_23691);
and U29768 (N_29768,N_20364,N_20888);
nor U29769 (N_29769,N_20174,N_23084);
nor U29770 (N_29770,N_22380,N_21969);
xor U29771 (N_29771,N_24928,N_22383);
nand U29772 (N_29772,N_23918,N_23313);
or U29773 (N_29773,N_23822,N_24082);
and U29774 (N_29774,N_22203,N_22134);
xor U29775 (N_29775,N_24688,N_20275);
and U29776 (N_29776,N_21539,N_24203);
nand U29777 (N_29777,N_22995,N_21133);
nor U29778 (N_29778,N_21920,N_23616);
or U29779 (N_29779,N_24676,N_23749);
or U29780 (N_29780,N_22986,N_21363);
nand U29781 (N_29781,N_21875,N_20443);
nand U29782 (N_29782,N_21399,N_22163);
nor U29783 (N_29783,N_23024,N_23395);
or U29784 (N_29784,N_21253,N_22324);
nor U29785 (N_29785,N_23049,N_24036);
xor U29786 (N_29786,N_22246,N_23542);
nand U29787 (N_29787,N_20003,N_23973);
or U29788 (N_29788,N_24839,N_21398);
nor U29789 (N_29789,N_21667,N_20851);
or U29790 (N_29790,N_24633,N_20734);
nor U29791 (N_29791,N_22977,N_23770);
or U29792 (N_29792,N_24280,N_21076);
nand U29793 (N_29793,N_22641,N_21231);
or U29794 (N_29794,N_21763,N_21334);
nand U29795 (N_29795,N_24122,N_24929);
or U29796 (N_29796,N_22466,N_20846);
xor U29797 (N_29797,N_23481,N_22460);
nand U29798 (N_29798,N_24664,N_24798);
or U29799 (N_29799,N_20978,N_23556);
nand U29800 (N_29800,N_24817,N_23316);
or U29801 (N_29801,N_23972,N_21396);
or U29802 (N_29802,N_21283,N_24524);
xor U29803 (N_29803,N_23156,N_22172);
and U29804 (N_29804,N_21412,N_23274);
nand U29805 (N_29805,N_24972,N_21824);
or U29806 (N_29806,N_21529,N_22277);
xnor U29807 (N_29807,N_21869,N_20460);
and U29808 (N_29808,N_23208,N_22693);
nand U29809 (N_29809,N_22976,N_22534);
xor U29810 (N_29810,N_23477,N_22776);
and U29811 (N_29811,N_21530,N_24917);
nor U29812 (N_29812,N_24287,N_23655);
or U29813 (N_29813,N_24955,N_21394);
or U29814 (N_29814,N_24905,N_23244);
or U29815 (N_29815,N_21813,N_24575);
or U29816 (N_29816,N_22816,N_24758);
nor U29817 (N_29817,N_24189,N_22825);
and U29818 (N_29818,N_24051,N_20687);
or U29819 (N_29819,N_22196,N_23538);
or U29820 (N_29820,N_23129,N_22814);
nor U29821 (N_29821,N_24674,N_23491);
or U29822 (N_29822,N_21688,N_23831);
or U29823 (N_29823,N_21898,N_21595);
xor U29824 (N_29824,N_23525,N_23842);
nand U29825 (N_29825,N_21716,N_20106);
nor U29826 (N_29826,N_21593,N_21846);
and U29827 (N_29827,N_21524,N_22979);
or U29828 (N_29828,N_21323,N_20488);
and U29829 (N_29829,N_24095,N_22840);
and U29830 (N_29830,N_20170,N_21848);
and U29831 (N_29831,N_24494,N_22844);
xnor U29832 (N_29832,N_24608,N_21409);
nand U29833 (N_29833,N_21332,N_21319);
nor U29834 (N_29834,N_24731,N_21749);
nand U29835 (N_29835,N_23059,N_23622);
nor U29836 (N_29836,N_22276,N_23827);
nor U29837 (N_29837,N_21952,N_24353);
nor U29838 (N_29838,N_20768,N_20578);
and U29839 (N_29839,N_21027,N_20637);
or U29840 (N_29840,N_24839,N_20650);
nand U29841 (N_29841,N_22613,N_23022);
nor U29842 (N_29842,N_22929,N_24052);
or U29843 (N_29843,N_23644,N_21748);
xnor U29844 (N_29844,N_21293,N_20641);
nor U29845 (N_29845,N_24177,N_20537);
xnor U29846 (N_29846,N_20399,N_20456);
or U29847 (N_29847,N_24083,N_21827);
nand U29848 (N_29848,N_21981,N_20876);
nand U29849 (N_29849,N_23488,N_21067);
and U29850 (N_29850,N_24127,N_23840);
xnor U29851 (N_29851,N_23546,N_21656);
xor U29852 (N_29852,N_21883,N_20642);
or U29853 (N_29853,N_22273,N_20225);
and U29854 (N_29854,N_24828,N_21460);
nor U29855 (N_29855,N_20702,N_20164);
nor U29856 (N_29856,N_24306,N_23133);
xor U29857 (N_29857,N_23576,N_24383);
or U29858 (N_29858,N_22173,N_20712);
nor U29859 (N_29859,N_24616,N_24968);
xnor U29860 (N_29860,N_23479,N_24812);
xnor U29861 (N_29861,N_24471,N_22972);
or U29862 (N_29862,N_24913,N_23366);
or U29863 (N_29863,N_22320,N_24032);
nand U29864 (N_29864,N_21457,N_20572);
xor U29865 (N_29865,N_24771,N_21556);
or U29866 (N_29866,N_22247,N_23263);
or U29867 (N_29867,N_21653,N_23514);
or U29868 (N_29868,N_20421,N_24203);
or U29869 (N_29869,N_22747,N_22096);
nand U29870 (N_29870,N_20556,N_21634);
and U29871 (N_29871,N_20070,N_22097);
xnor U29872 (N_29872,N_21579,N_24309);
nand U29873 (N_29873,N_20512,N_23448);
nand U29874 (N_29874,N_22533,N_21489);
nand U29875 (N_29875,N_22636,N_21410);
and U29876 (N_29876,N_23453,N_22229);
nor U29877 (N_29877,N_20397,N_22812);
nor U29878 (N_29878,N_20260,N_24550);
xor U29879 (N_29879,N_22927,N_24842);
or U29880 (N_29880,N_20605,N_21582);
xor U29881 (N_29881,N_20270,N_20953);
nor U29882 (N_29882,N_21578,N_23741);
nand U29883 (N_29883,N_20115,N_22595);
xor U29884 (N_29884,N_22090,N_20335);
nand U29885 (N_29885,N_20151,N_21753);
xnor U29886 (N_29886,N_23499,N_24864);
and U29887 (N_29887,N_20460,N_23705);
nor U29888 (N_29888,N_21030,N_20020);
xnor U29889 (N_29889,N_24196,N_22407);
and U29890 (N_29890,N_21010,N_23297);
nand U29891 (N_29891,N_21087,N_22860);
nor U29892 (N_29892,N_22542,N_22643);
or U29893 (N_29893,N_20319,N_20347);
or U29894 (N_29894,N_24004,N_24448);
xor U29895 (N_29895,N_22620,N_22740);
xor U29896 (N_29896,N_22464,N_23952);
and U29897 (N_29897,N_24730,N_21242);
nor U29898 (N_29898,N_22844,N_21927);
or U29899 (N_29899,N_21323,N_22002);
nor U29900 (N_29900,N_20436,N_24420);
nor U29901 (N_29901,N_24089,N_24104);
and U29902 (N_29902,N_20847,N_22363);
xnor U29903 (N_29903,N_24806,N_20245);
nand U29904 (N_29904,N_20512,N_24004);
and U29905 (N_29905,N_21142,N_24476);
nor U29906 (N_29906,N_24488,N_24049);
xnor U29907 (N_29907,N_21111,N_20356);
nand U29908 (N_29908,N_22836,N_23900);
nand U29909 (N_29909,N_20659,N_20798);
xnor U29910 (N_29910,N_22007,N_20688);
or U29911 (N_29911,N_22177,N_20144);
nand U29912 (N_29912,N_24640,N_23242);
and U29913 (N_29913,N_24549,N_21278);
xor U29914 (N_29914,N_22955,N_24732);
xnor U29915 (N_29915,N_24142,N_23380);
or U29916 (N_29916,N_23363,N_22847);
nand U29917 (N_29917,N_20780,N_22618);
or U29918 (N_29918,N_24887,N_24682);
or U29919 (N_29919,N_24126,N_24984);
and U29920 (N_29920,N_23630,N_22474);
and U29921 (N_29921,N_23271,N_23887);
nand U29922 (N_29922,N_20945,N_22395);
nor U29923 (N_29923,N_20894,N_21064);
nand U29924 (N_29924,N_24657,N_24015);
xor U29925 (N_29925,N_21902,N_24125);
and U29926 (N_29926,N_24550,N_20724);
xor U29927 (N_29927,N_24617,N_21501);
nor U29928 (N_29928,N_21908,N_24792);
or U29929 (N_29929,N_22875,N_24250);
or U29930 (N_29930,N_21786,N_22657);
or U29931 (N_29931,N_23874,N_23847);
nor U29932 (N_29932,N_20222,N_24682);
xor U29933 (N_29933,N_23360,N_20353);
nor U29934 (N_29934,N_22978,N_22301);
nor U29935 (N_29935,N_22628,N_21665);
nor U29936 (N_29936,N_20006,N_21151);
xor U29937 (N_29937,N_21698,N_22514);
or U29938 (N_29938,N_22261,N_22349);
xnor U29939 (N_29939,N_22151,N_22780);
nand U29940 (N_29940,N_20699,N_24165);
nor U29941 (N_29941,N_24396,N_20536);
or U29942 (N_29942,N_24117,N_20934);
or U29943 (N_29943,N_23754,N_22559);
or U29944 (N_29944,N_24238,N_22819);
xor U29945 (N_29945,N_22578,N_23855);
nor U29946 (N_29946,N_23803,N_22954);
xnor U29947 (N_29947,N_22787,N_20539);
and U29948 (N_29948,N_20884,N_23668);
xnor U29949 (N_29949,N_21436,N_23568);
nor U29950 (N_29950,N_24541,N_21837);
nand U29951 (N_29951,N_21326,N_21638);
or U29952 (N_29952,N_22175,N_23696);
or U29953 (N_29953,N_22702,N_24697);
nor U29954 (N_29954,N_23993,N_23007);
and U29955 (N_29955,N_21650,N_20869);
nand U29956 (N_29956,N_23147,N_24880);
nor U29957 (N_29957,N_21683,N_24548);
xnor U29958 (N_29958,N_20050,N_23965);
or U29959 (N_29959,N_20617,N_22295);
nand U29960 (N_29960,N_21316,N_22530);
nand U29961 (N_29961,N_22353,N_22576);
xor U29962 (N_29962,N_24394,N_24930);
nand U29963 (N_29963,N_21496,N_21010);
or U29964 (N_29964,N_23398,N_21744);
xnor U29965 (N_29965,N_23881,N_20861);
and U29966 (N_29966,N_23524,N_22422);
nor U29967 (N_29967,N_23523,N_24388);
nor U29968 (N_29968,N_23652,N_24948);
nand U29969 (N_29969,N_23949,N_22692);
and U29970 (N_29970,N_24347,N_24840);
nand U29971 (N_29971,N_23648,N_20439);
or U29972 (N_29972,N_22376,N_22066);
or U29973 (N_29973,N_20273,N_20981);
or U29974 (N_29974,N_21277,N_20241);
xnor U29975 (N_29975,N_20921,N_20363);
and U29976 (N_29976,N_21241,N_24741);
or U29977 (N_29977,N_22139,N_22729);
xnor U29978 (N_29978,N_24304,N_24513);
or U29979 (N_29979,N_21411,N_20908);
and U29980 (N_29980,N_24264,N_21400);
xor U29981 (N_29981,N_22369,N_24750);
xor U29982 (N_29982,N_22257,N_22905);
and U29983 (N_29983,N_21552,N_23800);
and U29984 (N_29984,N_23606,N_23346);
nor U29985 (N_29985,N_22413,N_20664);
xor U29986 (N_29986,N_22451,N_23120);
and U29987 (N_29987,N_22244,N_24217);
xnor U29988 (N_29988,N_23178,N_20081);
and U29989 (N_29989,N_24318,N_21937);
xor U29990 (N_29990,N_22669,N_20177);
nand U29991 (N_29991,N_21346,N_20199);
and U29992 (N_29992,N_21198,N_24368);
and U29993 (N_29993,N_22332,N_23080);
and U29994 (N_29994,N_20139,N_22650);
nand U29995 (N_29995,N_22153,N_22317);
xor U29996 (N_29996,N_21423,N_22444);
nand U29997 (N_29997,N_20340,N_22729);
xor U29998 (N_29998,N_22478,N_22547);
nor U29999 (N_29999,N_22982,N_22745);
xnor UO_0 (O_0,N_28780,N_26708);
or UO_1 (O_1,N_27621,N_27736);
or UO_2 (O_2,N_28029,N_27735);
and UO_3 (O_3,N_29770,N_26466);
nor UO_4 (O_4,N_28654,N_25341);
and UO_5 (O_5,N_27538,N_27379);
nand UO_6 (O_6,N_28612,N_29323);
xnor UO_7 (O_7,N_26634,N_25193);
nand UO_8 (O_8,N_27371,N_26417);
or UO_9 (O_9,N_25442,N_26756);
xnor UO_10 (O_10,N_28599,N_25619);
nor UO_11 (O_11,N_27980,N_25074);
xor UO_12 (O_12,N_27954,N_28486);
xor UO_13 (O_13,N_29468,N_27325);
nor UO_14 (O_14,N_27017,N_28877);
nor UO_15 (O_15,N_26981,N_25661);
xor UO_16 (O_16,N_26244,N_25237);
or UO_17 (O_17,N_27543,N_26400);
or UO_18 (O_18,N_27385,N_27902);
xnor UO_19 (O_19,N_28054,N_25445);
xor UO_20 (O_20,N_29650,N_29282);
xor UO_21 (O_21,N_29987,N_29307);
and UO_22 (O_22,N_29471,N_28159);
xor UO_23 (O_23,N_29975,N_28072);
nand UO_24 (O_24,N_27337,N_27135);
xnor UO_25 (O_25,N_26998,N_25976);
xor UO_26 (O_26,N_26801,N_27530);
xor UO_27 (O_27,N_29948,N_29620);
nand UO_28 (O_28,N_27851,N_27195);
nor UO_29 (O_29,N_25657,N_28846);
xnor UO_30 (O_30,N_29377,N_28539);
nand UO_31 (O_31,N_26633,N_26074);
nand UO_32 (O_32,N_25602,N_27079);
xnor UO_33 (O_33,N_26894,N_27947);
or UO_34 (O_34,N_28785,N_29357);
or UO_35 (O_35,N_29392,N_27210);
nor UO_36 (O_36,N_28023,N_26862);
or UO_37 (O_37,N_27316,N_26975);
xnor UO_38 (O_38,N_29832,N_27144);
nor UO_39 (O_39,N_28167,N_27244);
nand UO_40 (O_40,N_29305,N_28733);
or UO_41 (O_41,N_27842,N_26486);
nor UO_42 (O_42,N_26388,N_28228);
xor UO_43 (O_43,N_28391,N_28628);
or UO_44 (O_44,N_26919,N_28001);
nand UO_45 (O_45,N_27128,N_28764);
nand UO_46 (O_46,N_26306,N_29598);
and UO_47 (O_47,N_28763,N_26700);
xor UO_48 (O_48,N_28378,N_25601);
xnor UO_49 (O_49,N_26568,N_25233);
and UO_50 (O_50,N_28296,N_29351);
xnor UO_51 (O_51,N_29244,N_26911);
nor UO_52 (O_52,N_28342,N_25090);
xor UO_53 (O_53,N_27053,N_27977);
or UO_54 (O_54,N_25021,N_29943);
xnor UO_55 (O_55,N_26235,N_25891);
nor UO_56 (O_56,N_28817,N_29743);
xor UO_57 (O_57,N_26664,N_29311);
and UO_58 (O_58,N_27141,N_26612);
and UO_59 (O_59,N_26047,N_29224);
nand UO_60 (O_60,N_27357,N_26597);
or UO_61 (O_61,N_25905,N_27000);
nor UO_62 (O_62,N_29217,N_25775);
and UO_63 (O_63,N_27092,N_27704);
or UO_64 (O_64,N_28354,N_26576);
xnor UO_65 (O_65,N_25183,N_29499);
nor UO_66 (O_66,N_25269,N_26942);
nand UO_67 (O_67,N_29691,N_27453);
xor UO_68 (O_68,N_27292,N_29378);
xor UO_69 (O_69,N_27633,N_26348);
and UO_70 (O_70,N_28884,N_26991);
xnor UO_71 (O_71,N_25926,N_25952);
or UO_72 (O_72,N_28866,N_26647);
xnor UO_73 (O_73,N_27302,N_28907);
or UO_74 (O_74,N_29081,N_25963);
or UO_75 (O_75,N_25068,N_28281);
nand UO_76 (O_76,N_28913,N_28631);
and UO_77 (O_77,N_27953,N_29602);
xor UO_78 (O_78,N_29180,N_26187);
nand UO_79 (O_79,N_29717,N_26122);
or UO_80 (O_80,N_26358,N_26219);
or UO_81 (O_81,N_27682,N_29178);
xor UO_82 (O_82,N_26176,N_28475);
nor UO_83 (O_83,N_28519,N_27611);
or UO_84 (O_84,N_25480,N_26411);
or UO_85 (O_85,N_27884,N_29623);
nand UO_86 (O_86,N_27758,N_28337);
and UO_87 (O_87,N_27235,N_29732);
nand UO_88 (O_88,N_25155,N_25300);
xor UO_89 (O_89,N_25095,N_27271);
nand UO_90 (O_90,N_28273,N_26944);
or UO_91 (O_91,N_27309,N_27662);
and UO_92 (O_92,N_28618,N_26195);
and UO_93 (O_93,N_29154,N_29285);
nand UO_94 (O_94,N_29083,N_29248);
and UO_95 (O_95,N_26101,N_26424);
and UO_96 (O_96,N_26528,N_26505);
and UO_97 (O_97,N_27679,N_26740);
xnor UO_98 (O_98,N_25538,N_29874);
nor UO_99 (O_99,N_25908,N_29540);
or UO_100 (O_100,N_29947,N_29414);
xnor UO_101 (O_101,N_28885,N_27218);
nand UO_102 (O_102,N_25889,N_25276);
and UO_103 (O_103,N_28286,N_25366);
xnor UO_104 (O_104,N_25863,N_25877);
or UO_105 (O_105,N_29904,N_28948);
and UO_106 (O_106,N_25490,N_26766);
or UO_107 (O_107,N_29761,N_27564);
nor UO_108 (O_108,N_28955,N_26444);
nor UO_109 (O_109,N_25637,N_29266);
and UO_110 (O_110,N_28129,N_29258);
and UO_111 (O_111,N_27503,N_29954);
nand UO_112 (O_112,N_27067,N_26948);
and UO_113 (O_113,N_28362,N_27544);
xnor UO_114 (O_114,N_26820,N_26720);
nand UO_115 (O_115,N_25595,N_26208);
and UO_116 (O_116,N_27264,N_26645);
nand UO_117 (O_117,N_29187,N_28711);
xor UO_118 (O_118,N_27856,N_26504);
xnor UO_119 (O_119,N_28161,N_26931);
nand UO_120 (O_120,N_26478,N_27284);
nor UO_121 (O_121,N_26330,N_26540);
or UO_122 (O_122,N_27882,N_27771);
and UO_123 (O_123,N_27938,N_27402);
nand UO_124 (O_124,N_29902,N_29641);
nand UO_125 (O_125,N_26559,N_27133);
or UO_126 (O_126,N_25029,N_26549);
or UO_127 (O_127,N_25050,N_28416);
or UO_128 (O_128,N_27197,N_28626);
nor UO_129 (O_129,N_29665,N_26300);
nor UO_130 (O_130,N_27730,N_28431);
nor UO_131 (O_131,N_29461,N_25165);
nand UO_132 (O_132,N_29853,N_29012);
nor UO_133 (O_133,N_28174,N_28484);
and UO_134 (O_134,N_29800,N_26961);
and UO_135 (O_135,N_27972,N_27295);
xnor UO_136 (O_136,N_27482,N_27762);
or UO_137 (O_137,N_26248,N_25365);
nand UO_138 (O_138,N_28392,N_28542);
nand UO_139 (O_139,N_26937,N_25784);
xnor UO_140 (O_140,N_26648,N_27510);
or UO_141 (O_141,N_26075,N_27029);
or UO_142 (O_142,N_26643,N_27504);
and UO_143 (O_143,N_29016,N_28379);
and UO_144 (O_144,N_25496,N_26027);
nor UO_145 (O_145,N_27256,N_28075);
xor UO_146 (O_146,N_28201,N_27868);
or UO_147 (O_147,N_27314,N_29385);
nor UO_148 (O_148,N_27435,N_28942);
or UO_149 (O_149,N_25427,N_29664);
and UO_150 (O_150,N_26126,N_26377);
nor UO_151 (O_151,N_28576,N_25504);
xnor UO_152 (O_152,N_28941,N_27240);
xnor UO_153 (O_153,N_29595,N_27563);
xnor UO_154 (O_154,N_25166,N_28357);
nand UO_155 (O_155,N_25060,N_26024);
or UO_156 (O_156,N_27391,N_29865);
nor UO_157 (O_157,N_26326,N_28464);
or UO_158 (O_158,N_26710,N_25779);
xor UO_159 (O_159,N_28158,N_27594);
or UO_160 (O_160,N_27843,N_27162);
xnor UO_161 (O_161,N_27072,N_28382);
nor UO_162 (O_162,N_29269,N_26726);
nand UO_163 (O_163,N_25651,N_26000);
nor UO_164 (O_164,N_27459,N_28178);
nand UO_165 (O_165,N_26673,N_26134);
xor UO_166 (O_166,N_29097,N_27702);
nand UO_167 (O_167,N_27732,N_28731);
nand UO_168 (O_168,N_27012,N_25633);
and UO_169 (O_169,N_26038,N_27927);
nor UO_170 (O_170,N_25747,N_26669);
nand UO_171 (O_171,N_25100,N_27798);
or UO_172 (O_172,N_26392,N_26930);
or UO_173 (O_173,N_26192,N_26086);
nand UO_174 (O_174,N_26216,N_26696);
and UO_175 (O_175,N_25298,N_28369);
or UO_176 (O_176,N_28441,N_26618);
or UO_177 (O_177,N_26995,N_29166);
nor UO_178 (O_178,N_26996,N_26855);
nand UO_179 (O_179,N_29809,N_28397);
nand UO_180 (O_180,N_25282,N_27440);
or UO_181 (O_181,N_29630,N_26684);
or UO_182 (O_182,N_25058,N_27929);
or UO_183 (O_183,N_26514,N_29622);
xor UO_184 (O_184,N_26167,N_25236);
xnor UO_185 (O_185,N_25857,N_25346);
and UO_186 (O_186,N_25801,N_26905);
or UO_187 (O_187,N_27962,N_26125);
and UO_188 (O_188,N_28323,N_25688);
xnor UO_189 (O_189,N_25065,N_25259);
or UO_190 (O_190,N_29241,N_28643);
nand UO_191 (O_191,N_29886,N_29485);
nor UO_192 (O_192,N_27269,N_27005);
xor UO_193 (O_193,N_28360,N_29316);
or UO_194 (O_194,N_25921,N_25798);
or UO_195 (O_195,N_28261,N_27656);
xor UO_196 (O_196,N_27196,N_28220);
or UO_197 (O_197,N_28966,N_29214);
or UO_198 (O_198,N_27461,N_27180);
and UO_199 (O_199,N_28943,N_29532);
nand UO_200 (O_200,N_25448,N_27431);
or UO_201 (O_201,N_29679,N_29420);
nor UO_202 (O_202,N_26607,N_27088);
nor UO_203 (O_203,N_26875,N_28202);
xor UO_204 (O_204,N_25609,N_26200);
xnor UO_205 (O_205,N_28083,N_27703);
or UO_206 (O_206,N_28364,N_29444);
or UO_207 (O_207,N_27267,N_26839);
and UO_208 (O_208,N_26213,N_25027);
or UO_209 (O_209,N_26882,N_26529);
xnor UO_210 (O_210,N_27599,N_26776);
and UO_211 (O_211,N_27205,N_29139);
nand UO_212 (O_212,N_27750,N_28925);
xnor UO_213 (O_213,N_29249,N_29263);
nand UO_214 (O_214,N_27400,N_28007);
or UO_215 (O_215,N_26231,N_28901);
or UO_216 (O_216,N_26480,N_25443);
nor UO_217 (O_217,N_28675,N_28127);
xnor UO_218 (O_218,N_28213,N_27266);
nor UO_219 (O_219,N_27579,N_26547);
and UO_220 (O_220,N_25834,N_26508);
nor UO_221 (O_221,N_27025,N_25208);
nand UO_222 (O_222,N_27500,N_25349);
xnor UO_223 (O_223,N_27600,N_25869);
and UO_224 (O_224,N_26396,N_26688);
xor UO_225 (O_225,N_29935,N_27939);
and UO_226 (O_226,N_28592,N_27100);
and UO_227 (O_227,N_27462,N_26941);
xnor UO_228 (O_228,N_26232,N_27700);
nor UO_229 (O_229,N_28459,N_27148);
nand UO_230 (O_230,N_29921,N_25428);
xor UO_231 (O_231,N_26381,N_28240);
nand UO_232 (O_232,N_27891,N_27399);
xor UO_233 (O_233,N_28865,N_28059);
nand UO_234 (O_234,N_25856,N_25280);
xor UO_235 (O_235,N_25936,N_25572);
or UO_236 (O_236,N_29952,N_26376);
nor UO_237 (O_237,N_29931,N_27612);
xnor UO_238 (O_238,N_29867,N_26734);
or UO_239 (O_239,N_26056,N_25948);
and UO_240 (O_240,N_25671,N_25564);
nor UO_241 (O_241,N_29728,N_26644);
xnor UO_242 (O_242,N_28221,N_28556);
and UO_243 (O_243,N_26249,N_28635);
or UO_244 (O_244,N_26347,N_26520);
xnor UO_245 (O_245,N_27265,N_25813);
nor UO_246 (O_246,N_27796,N_27499);
and UO_247 (O_247,N_28291,N_27686);
nand UO_248 (O_248,N_28175,N_25698);
nor UO_249 (O_249,N_27283,N_28722);
or UO_250 (O_250,N_27877,N_25497);
nor UO_251 (O_251,N_26405,N_29463);
xnor UO_252 (O_252,N_25518,N_28580);
or UO_253 (O_253,N_25212,N_29544);
and UO_254 (O_254,N_29346,N_26535);
and UO_255 (O_255,N_28184,N_28204);
or UO_256 (O_256,N_25329,N_29155);
nor UO_257 (O_257,N_27427,N_27623);
nor UO_258 (O_258,N_25059,N_27108);
nor UO_259 (O_259,N_27950,N_28683);
nand UO_260 (O_260,N_27675,N_29920);
xnor UO_261 (O_261,N_28041,N_27469);
or UO_262 (O_262,N_26085,N_25778);
xor UO_263 (O_263,N_28741,N_27409);
xnor UO_264 (O_264,N_29573,N_25111);
nand UO_265 (O_265,N_27974,N_25937);
xor UO_266 (O_266,N_29327,N_27691);
nand UO_267 (O_267,N_29497,N_25854);
and UO_268 (O_268,N_28619,N_25870);
nor UO_269 (O_269,N_28791,N_29852);
nand UO_270 (O_270,N_26848,N_25591);
or UO_271 (O_271,N_25780,N_28971);
or UO_272 (O_272,N_26624,N_28010);
nor UO_273 (O_273,N_28322,N_29837);
nand UO_274 (O_274,N_27782,N_28128);
or UO_275 (O_275,N_27897,N_29391);
and UO_276 (O_276,N_27414,N_25393);
xor UO_277 (O_277,N_28566,N_25684);
nand UO_278 (O_278,N_26928,N_28777);
and UO_279 (O_279,N_26403,N_27712);
xnor UO_280 (O_280,N_25682,N_29252);
nand UO_281 (O_281,N_28652,N_26357);
xor UO_282 (O_282,N_26205,N_29143);
nand UO_283 (O_283,N_28513,N_25331);
or UO_284 (O_284,N_25249,N_28815);
nor UO_285 (O_285,N_27107,N_26433);
nor UO_286 (O_286,N_25075,N_25641);
nand UO_287 (O_287,N_27213,N_27751);
or UO_288 (O_288,N_27234,N_27155);
nand UO_289 (O_289,N_26265,N_29210);
or UO_290 (O_290,N_26211,N_27262);
xor UO_291 (O_291,N_25455,N_25291);
and UO_292 (O_292,N_26678,N_28544);
and UO_293 (O_293,N_29350,N_27278);
xnor UO_294 (O_294,N_27784,N_25529);
and UO_295 (O_295,N_26215,N_26611);
nand UO_296 (O_296,N_29086,N_26191);
or UO_297 (O_297,N_26580,N_29683);
nand UO_298 (O_298,N_25051,N_29631);
nand UO_299 (O_299,N_29675,N_25524);
xor UO_300 (O_300,N_27747,N_26041);
and UO_301 (O_301,N_26453,N_25104);
and UO_302 (O_302,N_29220,N_29149);
or UO_303 (O_303,N_28000,N_25097);
and UO_304 (O_304,N_28839,N_27415);
nand UO_305 (O_305,N_29245,N_29844);
nor UO_306 (O_306,N_25719,N_25132);
and UO_307 (O_307,N_29009,N_27584);
nor UO_308 (O_308,N_28284,N_28856);
nand UO_309 (O_309,N_29708,N_26587);
and UO_310 (O_310,N_29983,N_29669);
xor UO_311 (O_311,N_29303,N_29678);
and UO_312 (O_312,N_28254,N_27721);
nor UO_313 (O_313,N_26237,N_25965);
or UO_314 (O_314,N_25628,N_28444);
nand UO_315 (O_315,N_25645,N_26033);
nor UO_316 (O_316,N_29034,N_25765);
xor UO_317 (O_317,N_28597,N_28906);
nor UO_318 (O_318,N_29317,N_25589);
nand UO_319 (O_319,N_25613,N_25328);
nor UO_320 (O_320,N_27358,N_28526);
and UO_321 (O_321,N_25211,N_28454);
and UO_322 (O_322,N_25718,N_28976);
nand UO_323 (O_323,N_27588,N_29213);
nand UO_324 (O_324,N_29854,N_28481);
and UO_325 (O_325,N_26497,N_28090);
and UO_326 (O_326,N_27438,N_26925);
and UO_327 (O_327,N_27669,N_26774);
or UO_328 (O_328,N_25762,N_29797);
nand UO_329 (O_329,N_26501,N_28225);
nor UO_330 (O_330,N_28869,N_28659);
or UO_331 (O_331,N_25109,N_29625);
xnor UO_332 (O_332,N_29528,N_25175);
xnor UO_333 (O_333,N_27236,N_26676);
and UO_334 (O_334,N_29501,N_26923);
or UO_335 (O_335,N_28922,N_29308);
or UO_336 (O_336,N_26250,N_27908);
nand UO_337 (O_337,N_25103,N_26909);
nand UO_338 (O_338,N_26110,N_25554);
and UO_339 (O_339,N_25821,N_27508);
nor UO_340 (O_340,N_25987,N_28682);
and UO_341 (O_341,N_29491,N_27695);
and UO_342 (O_342,N_25864,N_26974);
nand UO_343 (O_343,N_26990,N_28418);
or UO_344 (O_344,N_25929,N_25939);
xor UO_345 (O_345,N_29193,N_27956);
or UO_346 (O_346,N_27049,N_28716);
xor UO_347 (O_347,N_29394,N_26117);
and UO_348 (O_348,N_25954,N_29821);
nor UO_349 (O_349,N_27446,N_29747);
xnor UO_350 (O_350,N_27963,N_25322);
xor UO_351 (O_351,N_25351,N_27631);
xnor UO_352 (O_352,N_29916,N_29600);
nand UO_353 (O_353,N_25321,N_29848);
or UO_354 (O_354,N_26201,N_29341);
nor UO_355 (O_355,N_27179,N_28546);
nor UO_356 (O_356,N_25374,N_27082);
and UO_357 (O_357,N_28779,N_27451);
xnor UO_358 (O_358,N_25604,N_28149);
nor UO_359 (O_359,N_25056,N_27912);
xor UO_360 (O_360,N_26261,N_25550);
nand UO_361 (O_361,N_28867,N_26295);
xor UO_362 (O_362,N_29056,N_26838);
nand UO_363 (O_363,N_25722,N_28697);
or UO_364 (O_364,N_28782,N_25915);
and UO_365 (O_365,N_26851,N_28594);
xor UO_366 (O_366,N_29360,N_29724);
xnor UO_367 (O_367,N_28849,N_25683);
nand UO_368 (O_368,N_25787,N_29087);
or UO_369 (O_369,N_25055,N_28545);
or UO_370 (O_370,N_27450,N_27320);
or UO_371 (O_371,N_26947,N_29015);
nor UO_372 (O_372,N_28155,N_25430);
or UO_373 (O_373,N_25559,N_29570);
nand UO_374 (O_374,N_25910,N_28844);
and UO_375 (O_375,N_29319,N_27984);
or UO_376 (O_376,N_29473,N_26097);
nand UO_377 (O_377,N_25663,N_26789);
xnor UO_378 (O_378,N_29782,N_29125);
or UO_379 (O_379,N_29880,N_27576);
nor UO_380 (O_380,N_29321,N_27019);
or UO_381 (O_381,N_27015,N_25896);
or UO_382 (O_382,N_29828,N_29980);
and UO_383 (O_383,N_27952,N_29612);
nand UO_384 (O_384,N_29615,N_28403);
xnor UO_385 (O_385,N_28577,N_28356);
xor UO_386 (O_386,N_27299,N_28340);
and UO_387 (O_387,N_28050,N_29337);
xnor UO_388 (O_388,N_28570,N_25188);
nor UO_389 (O_389,N_27916,N_26890);
and UO_390 (O_390,N_29896,N_27636);
nand UO_391 (O_391,N_27670,N_25522);
nor UO_392 (O_392,N_26441,N_25899);
or UO_393 (O_393,N_26590,N_29973);
nand UO_394 (O_394,N_25770,N_25528);
nand UO_395 (O_395,N_28008,N_27160);
nand UO_396 (O_396,N_25263,N_26681);
and UO_397 (O_397,N_25403,N_27849);
nand UO_398 (O_398,N_27145,N_28666);
or UO_399 (O_399,N_29838,N_25134);
nor UO_400 (O_400,N_27059,N_29450);
nor UO_401 (O_401,N_25724,N_25961);
and UO_402 (O_402,N_27672,N_27471);
nand UO_403 (O_403,N_26221,N_29813);
nand UO_404 (O_404,N_26432,N_25515);
or UO_405 (O_405,N_29847,N_26602);
nor UO_406 (O_406,N_26218,N_29972);
and UO_407 (O_407,N_27321,N_29968);
and UO_408 (O_408,N_27800,N_27976);
and UO_409 (O_409,N_26022,N_27447);
xnor UO_410 (O_410,N_29885,N_28203);
nand UO_411 (O_411,N_26687,N_27757);
nand UO_412 (O_412,N_26521,N_26360);
and UO_413 (O_413,N_28318,N_25725);
and UO_414 (O_414,N_29026,N_25498);
xnor UO_415 (O_415,N_27467,N_27540);
and UO_416 (O_416,N_28518,N_29052);
xnor UO_417 (O_417,N_26029,N_28543);
or UO_418 (O_418,N_25118,N_26915);
or UO_419 (O_419,N_27657,N_25019);
and UO_420 (O_420,N_27456,N_27258);
or UO_421 (O_421,N_28607,N_28346);
nand UO_422 (O_422,N_28478,N_25920);
and UO_423 (O_423,N_28796,N_26577);
and UO_424 (O_424,N_25973,N_29273);
or UO_425 (O_425,N_25157,N_28048);
xnor UO_426 (O_426,N_29982,N_26365);
nand UO_427 (O_427,N_28638,N_25841);
nand UO_428 (O_428,N_27795,N_28028);
or UO_429 (O_429,N_28555,N_29676);
xnor UO_430 (O_430,N_25859,N_27822);
nand UO_431 (O_431,N_27647,N_26281);
and UO_432 (O_432,N_26062,N_25536);
nand UO_433 (O_433,N_25851,N_29764);
and UO_434 (O_434,N_25689,N_25866);
xor UO_435 (O_435,N_26876,N_25986);
and UO_436 (O_436,N_26533,N_29705);
or UO_437 (O_437,N_28406,N_29553);
or UO_438 (O_438,N_28097,N_27616);
xor UO_439 (O_439,N_28825,N_27342);
xor UO_440 (O_440,N_25481,N_29132);
and UO_441 (O_441,N_25888,N_29208);
and UO_442 (O_442,N_26435,N_26879);
nand UO_443 (O_443,N_28584,N_27310);
xnor UO_444 (O_444,N_26922,N_25826);
and UO_445 (O_445,N_25418,N_26968);
xor UO_446 (O_446,N_26494,N_29788);
or UO_447 (O_447,N_25381,N_25930);
or UO_448 (O_448,N_28929,N_29151);
or UO_449 (O_449,N_26729,N_25224);
or UO_450 (O_450,N_27537,N_28841);
or UO_451 (O_451,N_25590,N_26236);
or UO_452 (O_452,N_26270,N_26808);
or UO_453 (O_453,N_29002,N_29978);
nor UO_454 (O_454,N_27147,N_25085);
or UO_455 (O_455,N_27065,N_28949);
nor UO_456 (O_456,N_29259,N_25071);
or UO_457 (O_457,N_28095,N_28415);
or UO_458 (O_458,N_26315,N_26155);
nand UO_459 (O_459,N_26588,N_25640);
and UO_460 (O_460,N_26457,N_27628);
or UO_461 (O_461,N_29870,N_27524);
xnor UO_462 (O_462,N_26818,N_25848);
or UO_463 (O_463,N_26375,N_26571);
nand UO_464 (O_464,N_28902,N_25495);
nor UO_465 (O_465,N_26378,N_27846);
and UO_466 (O_466,N_25196,N_29068);
nand UO_467 (O_467,N_27167,N_25199);
or UO_468 (O_468,N_27031,N_28645);
xnor UO_469 (O_469,N_28992,N_26049);
nor UO_470 (O_470,N_27193,N_29267);
nor UO_471 (O_471,N_26438,N_28786);
nor UO_472 (O_472,N_25385,N_25405);
nand UO_473 (O_473,N_28238,N_25964);
xor UO_474 (O_474,N_28714,N_25159);
and UO_475 (O_475,N_26321,N_27744);
xor UO_476 (O_476,N_28848,N_25685);
and UO_477 (O_477,N_28333,N_26002);
and UO_478 (O_478,N_28689,N_29798);
and UO_479 (O_479,N_28657,N_28473);
or UO_480 (O_480,N_28193,N_27909);
or UO_481 (O_481,N_29937,N_27539);
nand UO_482 (O_482,N_27166,N_28073);
nor UO_483 (O_483,N_29201,N_29912);
nor UO_484 (O_484,N_28368,N_27046);
nor UO_485 (O_485,N_28417,N_28836);
or UO_486 (O_486,N_26667,N_29616);
or UO_487 (O_487,N_29170,N_26007);
xor UO_488 (O_488,N_26121,N_29095);
and UO_489 (O_489,N_26764,N_27637);
nand UO_490 (O_490,N_28234,N_26793);
nand UO_491 (O_491,N_25143,N_29243);
nand UO_492 (O_492,N_29587,N_28353);
or UO_493 (O_493,N_25728,N_26982);
nand UO_494 (O_494,N_29869,N_26545);
and UO_495 (O_495,N_28512,N_28781);
xor UO_496 (O_496,N_27722,N_25273);
and UO_497 (O_497,N_29368,N_29542);
and UO_498 (O_498,N_28975,N_29069);
or UO_499 (O_499,N_29951,N_25117);
nor UO_500 (O_500,N_28850,N_27787);
nor UO_501 (O_501,N_29286,N_28080);
and UO_502 (O_502,N_29707,N_25845);
nor UO_503 (O_503,N_29851,N_28939);
and UO_504 (O_504,N_26115,N_25620);
nand UO_505 (O_505,N_27815,N_29742);
and UO_506 (O_506,N_28154,N_26565);
nand UO_507 (O_507,N_28456,N_28256);
and UO_508 (O_508,N_26309,N_26900);
xor UO_509 (O_509,N_25573,N_27665);
xnor UO_510 (O_510,N_26865,N_29137);
nor UO_511 (O_511,N_29660,N_26406);
or UO_512 (O_512,N_25168,N_28712);
and UO_513 (O_513,N_25045,N_28930);
and UO_514 (O_514,N_28229,N_29129);
xor UO_515 (O_515,N_27102,N_29799);
or UO_516 (O_516,N_27098,N_27498);
nor UO_517 (O_517,N_27737,N_29596);
and UO_518 (O_518,N_28384,N_27596);
nor UO_519 (O_519,N_25755,N_27847);
and UO_520 (O_520,N_27598,N_27439);
nand UO_521 (O_521,N_27401,N_26541);
nor UO_522 (O_522,N_28687,N_27604);
nand UO_523 (O_523,N_27306,N_26495);
or UO_524 (O_524,N_26778,N_28046);
nand UO_525 (O_525,N_27634,N_29247);
and UO_526 (O_526,N_25228,N_26462);
nor UO_527 (O_527,N_26302,N_29500);
and UO_528 (O_528,N_26429,N_29618);
and UO_529 (O_529,N_28868,N_28827);
or UO_530 (O_530,N_26324,N_27632);
or UO_531 (O_531,N_27701,N_28847);
and UO_532 (O_532,N_29292,N_28275);
xor UO_533 (O_533,N_26141,N_28207);
nand UO_534 (O_534,N_27985,N_27799);
and UO_535 (O_535,N_26596,N_29924);
and UO_536 (O_536,N_26168,N_27926);
nor UO_537 (O_537,N_29067,N_27417);
and UO_538 (O_538,N_29417,N_28890);
xor UO_539 (O_539,N_28376,N_28620);
xnor UO_540 (O_540,N_29253,N_27043);
or UO_541 (O_541,N_27169,N_29588);
nand UO_542 (O_542,N_25622,N_29933);
nand UO_543 (O_543,N_28642,N_29760);
xnor UO_544 (O_544,N_25460,N_29682);
and UO_545 (O_545,N_25639,N_27416);
nor UO_546 (O_546,N_27512,N_25962);
and UO_547 (O_547,N_25789,N_29965);
and UO_548 (O_548,N_27289,N_27245);
nor UO_549 (O_549,N_27788,N_29699);
and UO_550 (O_550,N_26404,N_28598);
or UO_551 (O_551,N_27806,N_25030);
nor UO_552 (O_552,N_28798,N_28380);
or UO_553 (O_553,N_27248,N_25476);
or UO_554 (O_554,N_29156,N_27569);
xnor UO_555 (O_555,N_29049,N_29653);
nand UO_556 (O_556,N_29262,N_29116);
nor UO_557 (O_557,N_27045,N_28200);
nand UO_558 (O_558,N_27086,N_29183);
nor UO_559 (O_559,N_28957,N_25239);
xor UO_560 (O_560,N_29498,N_25478);
xor UO_561 (O_561,N_26749,N_26765);
xnor UO_562 (O_562,N_29829,N_28892);
nand UO_563 (O_563,N_27381,N_27101);
xnor UO_564 (O_564,N_27898,N_28316);
nand UO_565 (O_565,N_25776,N_29369);
nand UO_566 (O_566,N_28878,N_29458);
and UO_567 (O_567,N_29505,N_25139);
or UO_568 (O_568,N_25261,N_29594);
xnor UO_569 (O_569,N_28747,N_26585);
xor UO_570 (O_570,N_29304,N_27641);
nand UO_571 (O_571,N_25969,N_26361);
nor UO_572 (O_572,N_29452,N_25658);
and UO_573 (O_573,N_28784,N_26325);
nand UO_574 (O_574,N_25325,N_27810);
nand UO_575 (O_575,N_28426,N_25025);
nor UO_576 (O_576,N_27883,N_25985);
or UO_577 (O_577,N_27013,N_29148);
nand UO_578 (O_578,N_26864,N_28088);
nand UO_579 (O_579,N_27678,N_27738);
nor UO_580 (O_580,N_25187,N_28797);
nor UO_581 (O_581,N_27250,N_29533);
or UO_582 (O_582,N_27780,N_28259);
or UO_583 (O_583,N_26318,N_28003);
nor UO_584 (O_584,N_29758,N_26183);
or UO_585 (O_585,N_28591,N_29651);
xor UO_586 (O_586,N_27388,N_26656);
nand UO_587 (O_587,N_25842,N_28433);
nand UO_588 (O_588,N_26127,N_28181);
xnor UO_589 (O_589,N_27718,N_26222);
xor UO_590 (O_590,N_29176,N_26118);
nand UO_591 (O_591,N_26071,N_26352);
nor UO_592 (O_592,N_25177,N_27237);
nor UO_593 (O_593,N_27609,N_26952);
xnor UO_594 (O_594,N_25003,N_26706);
nor UO_595 (O_595,N_26387,N_26096);
nor UO_596 (O_596,N_27561,N_25951);
nand UO_597 (O_597,N_25753,N_25484);
and UO_598 (O_598,N_26976,N_29716);
and UO_599 (O_599,N_26735,N_29729);
xnor UO_600 (O_600,N_27685,N_27690);
or UO_601 (O_601,N_28617,N_28037);
or UO_602 (O_602,N_28452,N_28325);
nand UO_603 (O_603,N_27617,N_27714);
nand UO_604 (O_604,N_26537,N_29167);
or UO_605 (O_605,N_25711,N_26653);
nor UO_606 (O_606,N_26994,N_27465);
and UO_607 (O_607,N_26359,N_26694);
xor UO_608 (O_608,N_26052,N_28695);
and UO_609 (O_609,N_29476,N_26476);
and UO_610 (O_610,N_29223,N_27125);
xor UO_611 (O_611,N_25412,N_25015);
xor UO_612 (O_612,N_29804,N_25467);
nand UO_613 (O_613,N_25326,N_29845);
xnor UO_614 (O_614,N_28529,N_27434);
xor UO_615 (O_615,N_25486,N_27315);
xor UO_616 (O_616,N_26255,N_25284);
nor UO_617 (O_617,N_27332,N_28588);
nor UO_618 (O_618,N_29467,N_26556);
nor UO_619 (O_619,N_25472,N_25664);
nand UO_620 (O_620,N_26355,N_28537);
nand UO_621 (O_621,N_29750,N_27556);
nand UO_622 (O_622,N_27261,N_25608);
or UO_623 (O_623,N_25707,N_26093);
nand UO_624 (O_624,N_29296,N_25130);
xor UO_625 (O_625,N_28341,N_28504);
nand UO_626 (O_626,N_29073,N_27188);
nand UO_627 (O_627,N_26539,N_29915);
or UO_628 (O_628,N_28845,N_27823);
xnor UO_629 (O_629,N_25678,N_26140);
or UO_630 (O_630,N_29212,N_25947);
nand UO_631 (O_631,N_27833,N_26910);
xor UO_632 (O_632,N_26985,N_28801);
and UO_633 (O_633,N_25172,N_27116);
nand UO_634 (O_634,N_28265,N_29046);
nand UO_635 (O_635,N_28505,N_26420);
nand UO_636 (O_636,N_28699,N_29445);
and UO_637 (O_637,N_25807,N_25918);
and UO_638 (O_638,N_28448,N_26335);
xor UO_639 (O_639,N_26665,N_29158);
or UO_640 (O_640,N_25176,N_29431);
nand UO_641 (O_641,N_25756,N_27991);
and UO_642 (O_642,N_26654,N_27554);
and UO_643 (O_643,N_25454,N_25686);
nor UO_644 (O_644,N_27684,N_26697);
or UO_645 (O_645,N_25000,N_26721);
nor UO_646 (O_646,N_26847,N_26812);
nand UO_647 (O_647,N_29917,N_29860);
nand UO_648 (O_648,N_28162,N_28349);
and UO_649 (O_649,N_27478,N_25038);
nor UO_650 (O_650,N_27497,N_25674);
or UO_651 (O_651,N_27859,N_26374);
or UO_652 (O_652,N_28311,N_27352);
nand UO_653 (O_653,N_25283,N_26807);
and UO_654 (O_654,N_29523,N_28834);
or UO_655 (O_655,N_25989,N_25867);
and UO_656 (O_656,N_25413,N_25423);
nor UO_657 (O_657,N_25562,N_26574);
and UO_658 (O_658,N_27557,N_29179);
and UO_659 (O_659,N_29908,N_25927);
and UO_660 (O_660,N_25794,N_26651);
or UO_661 (O_661,N_28191,N_29106);
and UO_662 (O_662,N_28215,N_26391);
or UO_663 (O_663,N_27327,N_29996);
or UO_664 (O_664,N_26507,N_26763);
or UO_665 (O_665,N_26709,N_26560);
and UO_666 (O_666,N_28144,N_28746);
and UO_667 (O_667,N_26419,N_26434);
nor UO_668 (O_668,N_27146,N_26316);
nand UO_669 (O_669,N_25161,N_26933);
xor UO_670 (O_670,N_27343,N_25911);
nand UO_671 (O_671,N_25646,N_27058);
and UO_672 (O_672,N_28663,N_29739);
and UO_673 (O_673,N_28414,N_25360);
xor UO_674 (O_674,N_27801,N_25890);
and UO_675 (O_675,N_29988,N_27073);
and UO_676 (O_676,N_28717,N_28432);
and UO_677 (O_677,N_26436,N_27872);
or UO_678 (O_678,N_27724,N_27477);
or UO_679 (O_679,N_28899,N_28453);
nand UO_680 (O_680,N_26790,N_28068);
or UO_681 (O_681,N_25292,N_27903);
xor UO_682 (O_682,N_26761,N_28742);
or UO_683 (O_683,N_29407,N_26209);
and UO_684 (O_684,N_26017,N_28060);
nand UO_685 (O_685,N_25897,N_26522);
and UO_686 (O_686,N_26791,N_28115);
and UO_687 (O_687,N_25214,N_29925);
or UO_688 (O_688,N_27021,N_28977);
and UO_689 (O_689,N_29127,N_26011);
or UO_690 (O_690,N_26668,N_26379);
nand UO_691 (O_691,N_25675,N_28732);
nor UO_692 (O_692,N_27026,N_28172);
nor UO_693 (O_693,N_29541,N_25310);
or UO_694 (O_694,N_29521,N_29956);
or UO_695 (O_695,N_29042,N_25102);
or UO_696 (O_696,N_25617,N_27648);
nor UO_697 (O_697,N_25943,N_25493);
nor UO_698 (O_698,N_29041,N_29992);
xnor UO_699 (O_699,N_25309,N_29211);
nor UO_700 (O_700,N_27683,N_28520);
nor UO_701 (O_701,N_27990,N_29383);
nand UO_702 (O_702,N_28399,N_27163);
xnor UO_703 (O_703,N_26308,N_26967);
and UO_704 (O_704,N_26646,N_28335);
and UO_705 (O_705,N_28875,N_28319);
and UO_706 (O_706,N_25414,N_28334);
or UO_707 (O_707,N_28729,N_27033);
nand UO_708 (O_708,N_28105,N_25392);
nand UO_709 (O_709,N_26686,N_29453);
nand UO_710 (O_710,N_27729,N_25362);
or UO_711 (O_711,N_29677,N_28077);
nand UO_712 (O_712,N_27091,N_25067);
nor UO_713 (O_713,N_27231,N_25703);
nand UO_714 (O_714,N_27590,N_29637);
and UO_715 (O_715,N_27624,N_25561);
nand UO_716 (O_716,N_28525,N_27644);
nand UO_717 (O_717,N_26572,N_27591);
nand UO_718 (O_718,N_26685,N_25417);
or UO_719 (O_719,N_29111,N_25350);
nand UO_720 (O_720,N_29567,N_29215);
nor UO_721 (O_721,N_28277,N_26143);
nor UO_722 (O_722,N_25127,N_25406);
nand UO_723 (O_723,N_27666,N_28024);
or UO_724 (O_724,N_25063,N_28737);
nor UO_725 (O_725,N_27376,N_27946);
and UO_726 (O_726,N_28987,N_29538);
nand UO_727 (O_727,N_28078,N_27646);
and UO_728 (O_728,N_25881,N_29725);
nor UO_729 (O_729,N_26451,N_26510);
nor UO_730 (O_730,N_29990,N_28107);
xor UO_731 (O_731,N_28968,N_25184);
xnor UO_732 (O_732,N_29736,N_27153);
nor UO_733 (O_733,N_27552,N_27723);
nor UO_734 (O_734,N_28100,N_29159);
xnor UO_735 (O_735,N_26770,N_25610);
or UO_736 (O_736,N_29078,N_25073);
nand UO_737 (O_737,N_29063,N_25482);
or UO_738 (O_738,N_26061,N_26512);
nand UO_739 (O_739,N_29551,N_26418);
or UO_740 (O_740,N_26977,N_26103);
nor UO_741 (O_741,N_29608,N_29836);
nand UO_742 (O_742,N_29873,N_28678);
or UO_743 (O_743,N_25934,N_25377);
nor UO_744 (O_744,N_28548,N_25824);
xor UO_745 (O_745,N_27515,N_28605);
or UO_746 (O_746,N_29994,N_28749);
and UO_747 (O_747,N_28124,N_29367);
and UO_748 (O_748,N_25483,N_27494);
or UO_749 (O_749,N_27699,N_26005);
xor UO_750 (O_750,N_26058,N_25838);
and UO_751 (O_751,N_27081,N_28015);
xor UO_752 (O_752,N_25654,N_26532);
nand UO_753 (O_753,N_27194,N_27192);
xor UO_754 (O_754,N_27054,N_28049);
or UO_755 (O_755,N_25694,N_28690);
nor UO_756 (O_756,N_26133,N_28231);
and UO_757 (O_757,N_29007,N_28084);
and UO_758 (O_758,N_26935,N_27037);
nand UO_759 (O_759,N_29435,N_27206);
nand UO_760 (O_760,N_26286,N_28062);
and UO_761 (O_761,N_28226,N_28727);
xnor UO_762 (O_762,N_29926,N_26344);
and UO_763 (O_763,N_25978,N_28163);
and UO_764 (O_764,N_25267,N_29218);
nor UO_765 (O_765,N_28960,N_29181);
xnor UO_766 (O_766,N_27571,N_25505);
and UO_767 (O_767,N_25565,N_25129);
nand UO_768 (O_768,N_26616,N_25795);
xor UO_769 (O_769,N_28551,N_28411);
nor UO_770 (O_770,N_25627,N_25861);
nor UO_771 (O_771,N_27513,N_28183);
nor UO_772 (O_772,N_26692,N_26262);
nor UO_773 (O_773,N_28569,N_26733);
and UO_774 (O_774,N_26305,N_27746);
nand UO_775 (O_775,N_29816,N_25110);
or UO_776 (O_776,N_26670,N_28070);
or UO_777 (O_777,N_25148,N_27587);
and UO_778 (O_778,N_26257,N_28314);
xnor UO_779 (O_779,N_29353,N_25031);
and UO_780 (O_780,N_26186,N_28171);
nand UO_781 (O_781,N_27774,N_25582);
or UO_782 (O_782,N_25342,N_28713);
nor UO_783 (O_783,N_26500,N_29493);
nor UO_784 (O_784,N_27115,N_29028);
nand UO_785 (O_785,N_25796,N_29328);
nor UO_786 (O_786,N_29470,N_27254);
or UO_787 (O_787,N_27429,N_27535);
or UO_788 (O_788,N_27981,N_27836);
and UO_789 (O_789,N_27386,N_29923);
or UO_790 (O_790,N_26267,N_26997);
nand UO_791 (O_791,N_29374,N_27362);
nand UO_792 (O_792,N_27663,N_29361);
and UO_793 (O_793,N_27472,N_25234);
or UO_794 (O_794,N_26785,N_26567);
or UO_795 (O_795,N_29457,N_25123);
nor UO_796 (O_796,N_29513,N_29636);
or UO_797 (O_797,N_25944,N_27159);
or UO_798 (O_798,N_27992,N_25942);
or UO_799 (O_799,N_27649,N_28517);
or UO_800 (O_800,N_28532,N_25040);
and UO_801 (O_801,N_26819,N_27126);
nand UO_802 (O_802,N_29864,N_26349);
and UO_803 (O_803,N_28536,N_25421);
and UO_804 (O_804,N_27252,N_26707);
nand UO_805 (O_805,N_26001,N_27495);
xor UO_806 (O_806,N_28246,N_25875);
or UO_807 (O_807,N_26336,N_29197);
or UO_808 (O_808,N_28696,N_27001);
xnor UO_809 (O_809,N_28224,N_25556);
nand UO_810 (O_810,N_27999,N_29586);
xnor UO_811 (O_811,N_28725,N_25717);
xor UO_812 (O_812,N_29393,N_27793);
xor UO_813 (O_813,N_26965,N_28460);
nand UO_814 (O_814,N_27770,N_26714);
xnor UO_815 (O_815,N_25532,N_28019);
xnor UO_816 (O_816,N_25708,N_26130);
or UO_817 (O_817,N_26102,N_29101);
or UO_818 (O_818,N_27792,N_25988);
nand UO_819 (O_819,N_28744,N_26446);
xor UO_820 (O_820,N_28662,N_28701);
and UO_821 (O_821,N_25024,N_27889);
or UO_822 (O_822,N_27454,N_27233);
or UO_823 (O_823,N_28236,N_25049);
xor UO_824 (O_824,N_25347,N_27111);
xnor UO_825 (O_825,N_28004,N_28561);
nand UO_826 (O_826,N_28489,N_26384);
nand UO_827 (O_827,N_28936,N_26897);
nand UO_828 (O_828,N_26491,N_27601);
or UO_829 (O_829,N_29585,N_29072);
or UO_830 (O_830,N_26342,N_26842);
nand UO_831 (O_831,N_25474,N_28112);
xor UO_832 (O_832,N_27363,N_28851);
or UO_833 (O_833,N_28534,N_27660);
nand UO_834 (O_834,N_26456,N_25169);
xor UO_835 (O_835,N_28616,N_29107);
nor UO_836 (O_836,N_25540,N_25083);
and UO_837 (O_837,N_25048,N_26962);
nand UO_838 (O_838,N_26885,N_25053);
or UO_839 (O_839,N_26650,N_29710);
nand UO_840 (O_840,N_29840,N_25285);
and UO_841 (O_841,N_26546,N_29577);
and UO_842 (O_842,N_25398,N_26775);
xnor UO_843 (O_843,N_26924,N_26803);
or UO_844 (O_844,N_28595,N_26426);
nor UO_845 (O_845,N_29079,N_29597);
or UO_846 (O_846,N_25140,N_27214);
or UO_847 (O_847,N_26279,N_26260);
nand UO_848 (O_848,N_26169,N_27650);
nand UO_849 (O_849,N_29958,N_27406);
xnor UO_850 (O_850,N_29380,N_29726);
nand UO_851 (O_851,N_26832,N_29757);
and UO_852 (O_852,N_25709,N_27551);
or UO_853 (O_853,N_28671,N_29657);
xor UO_854 (O_854,N_26723,N_29238);
or UO_855 (O_855,N_28298,N_25774);
or UO_856 (O_856,N_29720,N_28887);
xor UO_857 (O_857,N_26196,N_26291);
xor UO_858 (O_858,N_25151,N_28921);
nand UO_859 (O_859,N_27773,N_25205);
or UO_860 (O_860,N_27921,N_27297);
nand UO_861 (O_861,N_27520,N_26869);
nand UO_862 (O_862,N_25981,N_28412);
nor UO_863 (O_863,N_27533,N_26263);
and UO_864 (O_864,N_29647,N_28153);
xor UO_865 (O_865,N_29753,N_25732);
or UO_866 (O_866,N_29986,N_26171);
nor UO_867 (O_867,N_26100,N_29163);
or UO_868 (O_868,N_25967,N_25315);
nor UO_869 (O_869,N_28371,N_28715);
or UO_870 (O_870,N_28123,N_29820);
xor UO_871 (O_871,N_27090,N_28043);
nand UO_872 (O_872,N_29347,N_29057);
nand UO_873 (O_873,N_29496,N_27209);
nor UO_874 (O_874,N_25666,N_26053);
or UO_875 (O_875,N_26698,N_25547);
and UO_876 (O_876,N_28272,N_28157);
and UO_877 (O_877,N_26292,N_25008);
and UO_878 (O_878,N_26943,N_28549);
nor UO_879 (O_879,N_29202,N_27789);
and UO_880 (O_880,N_27693,N_25793);
nor UO_881 (O_881,N_28165,N_29581);
or UO_882 (O_882,N_25240,N_27216);
nand UO_883 (O_883,N_28299,N_29607);
xor UO_884 (O_884,N_27989,N_28754);
nor UO_885 (O_885,N_25659,N_27501);
and UO_886 (O_886,N_28728,N_28860);
nand UO_887 (O_887,N_28956,N_29900);
and UO_888 (O_888,N_28541,N_29849);
xnor UO_889 (O_889,N_28071,N_28313);
nor UO_890 (O_890,N_29324,N_27536);
nand UO_891 (O_891,N_27474,N_29693);
or UO_892 (O_892,N_25201,N_28248);
nor UO_893 (O_893,N_28720,N_25064);
and UO_894 (O_894,N_25307,N_26239);
or UO_895 (O_895,N_26859,N_26428);
or UO_896 (O_896,N_27442,N_28709);
xor UO_897 (O_897,N_27064,N_25380);
or UO_898 (O_898,N_25402,N_25054);
or UO_899 (O_899,N_29235,N_27577);
or UO_900 (O_900,N_26802,N_25082);
nor UO_901 (O_901,N_28708,N_26028);
or UO_902 (O_902,N_27642,N_27445);
and UO_903 (O_903,N_29254,N_29783);
or UO_904 (O_904,N_28710,N_27835);
and UO_905 (O_905,N_28982,N_29939);
nor UO_906 (O_906,N_29053,N_27251);
nand UO_907 (O_907,N_28169,N_29370);
or UO_908 (O_908,N_29556,N_29746);
and UO_909 (O_909,N_29070,N_26278);
nand UO_910 (O_910,N_28324,N_29227);
and UO_911 (O_911,N_26475,N_27692);
nand UO_912 (O_912,N_26119,N_28624);
nor UO_913 (O_913,N_25806,N_29325);
nor UO_914 (O_914,N_27331,N_26402);
nor UO_915 (O_915,N_27667,N_27760);
xor UO_916 (O_916,N_27466,N_28658);
nand UO_917 (O_917,N_28745,N_28496);
nor UO_918 (O_918,N_25710,N_28895);
xor UO_919 (O_919,N_29349,N_25598);
or UO_920 (O_920,N_26662,N_25539);
or UO_921 (O_921,N_26020,N_26334);
xnor UO_922 (O_922,N_28765,N_29005);
nor UO_923 (O_923,N_28199,N_29010);
nand UO_924 (O_924,N_28790,N_25142);
xor UO_925 (O_925,N_28672,N_27680);
nand UO_926 (O_926,N_29702,N_25179);
nor UO_927 (O_927,N_28276,N_29177);
xor UO_928 (O_928,N_27296,N_28030);
or UO_929 (O_929,N_26247,N_29440);
nand UO_930 (O_930,N_29017,N_29893);
xnor UO_931 (O_931,N_26206,N_28122);
nor UO_932 (O_932,N_27355,N_29433);
and UO_933 (O_933,N_29510,N_29422);
nand UO_934 (O_934,N_29089,N_29140);
nor UO_935 (O_935,N_28400,N_25318);
and UO_936 (O_936,N_29226,N_26068);
nand UO_937 (O_937,N_27925,N_29606);
nor UO_938 (O_938,N_28422,N_28034);
or UO_939 (O_939,N_27971,N_29464);
or UO_940 (O_940,N_25147,N_28301);
and UO_941 (O_941,N_29108,N_27074);
nor UO_942 (O_942,N_29564,N_28094);
or UO_943 (O_943,N_27275,N_29356);
nor UO_944 (O_944,N_29727,N_26181);
nor UO_945 (O_945,N_26786,N_25670);
nand UO_946 (O_946,N_27928,N_25805);
nor UO_947 (O_947,N_29756,N_25923);
or UO_948 (O_948,N_29898,N_27791);
or UO_949 (O_949,N_29401,N_29745);
or UO_950 (O_950,N_27915,N_28533);
or UO_951 (O_951,N_26254,N_29998);
nor UO_952 (O_952,N_26088,N_28615);
and UO_953 (O_953,N_25337,N_26442);
xnor UO_954 (O_954,N_27328,N_26304);
nand UO_955 (O_955,N_25216,N_28893);
xnor UO_956 (O_956,N_25026,N_28247);
xor UO_957 (O_957,N_28563,N_29550);
nor UO_958 (O_958,N_25191,N_27523);
xor UO_959 (O_959,N_27452,N_26652);
or UO_960 (O_960,N_29776,N_28994);
nor UO_961 (O_961,N_29999,N_25946);
or UO_962 (O_962,N_28021,N_27048);
and UO_963 (O_963,N_27689,N_29681);
nor UO_964 (O_964,N_29090,N_25116);
nor UO_965 (O_965,N_27444,N_25232);
xor UO_966 (O_966,N_28510,N_28446);
and UO_967 (O_967,N_29738,N_27769);
xor UO_968 (O_968,N_25372,N_28651);
nor UO_969 (O_969,N_27268,N_28788);
or UO_970 (O_970,N_27725,N_29288);
and UO_971 (O_971,N_29927,N_28211);
xnor UO_972 (O_972,N_29246,N_28562);
xnor UO_973 (O_973,N_28274,N_25679);
nor UO_974 (O_974,N_26730,N_25832);
xor UO_975 (O_975,N_29576,N_26988);
xor UO_976 (O_976,N_26946,N_28358);
and UO_977 (O_977,N_29913,N_28560);
or UO_978 (O_978,N_28036,N_28343);
or UO_979 (O_979,N_29668,N_28898);
nand UO_980 (O_980,N_25812,N_25457);
nand UO_981 (O_981,N_25681,N_28470);
or UO_982 (O_982,N_29780,N_26016);
nor UO_983 (O_983,N_28758,N_29115);
nand UO_984 (O_984,N_25091,N_28531);
xnor UO_985 (O_985,N_29817,N_29878);
nor UO_986 (O_986,N_25788,N_25189);
nand UO_987 (O_987,N_26164,N_25904);
xnor UO_988 (O_988,N_26617,N_25563);
nand UO_989 (O_989,N_25013,N_28586);
or UO_990 (O_990,N_28833,N_27841);
or UO_991 (O_991,N_27198,N_26973);
nand UO_992 (O_992,N_29735,N_26256);
or UO_993 (O_993,N_27368,N_28092);
or UO_994 (O_994,N_25037,N_29520);
nor UO_995 (O_995,N_29082,N_26630);
and UO_996 (O_996,N_27437,N_26312);
and UO_997 (O_997,N_25886,N_25435);
and UO_998 (O_998,N_26212,N_25072);
xnor UO_999 (O_999,N_25734,N_28862);
and UO_1000 (O_1000,N_28130,N_29099);
or UO_1001 (O_1001,N_27668,N_25729);
or UO_1002 (O_1002,N_28738,N_29946);
nor UO_1003 (O_1003,N_28794,N_27460);
nand UO_1004 (O_1004,N_29460,N_27565);
nand UO_1005 (O_1005,N_28640,N_25882);
and UO_1006 (O_1006,N_25933,N_29013);
xnor UO_1007 (O_1007,N_26955,N_29436);
nor UO_1008 (O_1008,N_27983,N_26674);
nand UO_1009 (O_1009,N_25182,N_27906);
xnor UO_1010 (O_1010,N_25348,N_27931);
nand UO_1011 (O_1011,N_27455,N_26912);
and UO_1012 (O_1012,N_27177,N_28109);
nor UO_1013 (O_1013,N_28434,N_25131);
and UO_1014 (O_1014,N_28550,N_26180);
or UO_1015 (O_1015,N_25652,N_25126);
nand UO_1016 (O_1016,N_28006,N_25420);
and UO_1017 (O_1017,N_27221,N_25568);
nor UO_1018 (O_1018,N_29519,N_29001);
or UO_1019 (O_1019,N_27138,N_25022);
and UO_1020 (O_1020,N_29967,N_27945);
and UO_1021 (O_1021,N_27246,N_26054);
or UO_1022 (O_1022,N_25431,N_26104);
xnor UO_1023 (O_1023,N_27865,N_26156);
or UO_1024 (O_1024,N_29811,N_29278);
nor UO_1025 (O_1025,N_28967,N_28888);
or UO_1026 (O_1026,N_26124,N_29762);
xnor UO_1027 (O_1027,N_27532,N_27281);
and UO_1028 (O_1028,N_29807,N_28150);
nand UO_1029 (O_1029,N_29569,N_29071);
or UO_1030 (O_1030,N_28194,N_26666);
xnor UO_1031 (O_1031,N_29387,N_25530);
and UO_1032 (O_1032,N_27940,N_25209);
nor UO_1033 (O_1033,N_25593,N_26227);
xor UO_1034 (O_1034,N_28096,N_29779);
xnor UO_1035 (O_1035,N_29275,N_26956);
and UO_1036 (O_1036,N_25636,N_26311);
and UO_1037 (O_1037,N_27011,N_26179);
nor UO_1038 (O_1038,N_27028,N_28926);
and UO_1039 (O_1039,N_28748,N_29152);
nor UO_1040 (O_1040,N_29640,N_27473);
and UO_1041 (O_1041,N_29604,N_28824);
nor UO_1042 (O_1042,N_25512,N_29748);
and UO_1043 (O_1043,N_25466,N_27639);
or UO_1044 (O_1044,N_26613,N_29029);
xor UO_1045 (O_1045,N_29634,N_29455);
and UO_1046 (O_1046,N_28168,N_27397);
nor UO_1047 (O_1047,N_26273,N_25735);
or UO_1048 (O_1048,N_26903,N_25194);
and UO_1049 (O_1049,N_29366,N_26702);
nand UO_1050 (O_1050,N_26683,N_25740);
and UO_1051 (O_1051,N_26896,N_28692);
or UO_1052 (O_1052,N_29442,N_25763);
or UO_1053 (O_1053,N_29033,N_25108);
or UO_1054 (O_1054,N_29684,N_26422);
xnor UO_1055 (O_1055,N_26189,N_27651);
nand UO_1056 (O_1056,N_26437,N_27080);
xnor UO_1057 (O_1057,N_27249,N_25144);
and UO_1058 (O_1058,N_26868,N_28195);
nand UO_1059 (O_1059,N_28074,N_25260);
nor UO_1060 (O_1060,N_29555,N_28217);
and UO_1061 (O_1061,N_25804,N_28385);
and UO_1062 (O_1062,N_29793,N_27139);
and UO_1063 (O_1063,N_27652,N_25043);
xnor UO_1064 (O_1064,N_27307,N_26363);
nor UO_1065 (O_1065,N_26809,N_26578);
xor UO_1066 (O_1066,N_27226,N_27345);
and UO_1067 (O_1067,N_27852,N_28771);
or UO_1068 (O_1068,N_26979,N_28182);
nor UO_1069 (O_1069,N_26188,N_28972);
or UO_1070 (O_1070,N_27560,N_25621);
and UO_1071 (O_1071,N_27134,N_28212);
or UO_1072 (O_1072,N_25585,N_26095);
nand UO_1073 (O_1073,N_25676,N_27492);
or UO_1074 (O_1074,N_29314,N_28661);
nand UO_1075 (O_1075,N_25492,N_25761);
or UO_1076 (O_1076,N_29580,N_28552);
nor UO_1077 (O_1077,N_27318,N_28302);
and UO_1078 (O_1078,N_26109,N_29236);
nand UO_1079 (O_1079,N_26628,N_28953);
and UO_1080 (O_1080,N_28056,N_27227);
nand UO_1081 (O_1081,N_25754,N_28608);
nor UO_1082 (O_1082,N_26246,N_28753);
nand UO_1083 (O_1083,N_27761,N_25584);
or UO_1084 (O_1084,N_27071,N_29552);
nand UO_1085 (O_1085,N_29237,N_28035);
xor UO_1086 (O_1086,N_25324,N_25907);
or UO_1087 (O_1087,N_29768,N_28700);
nand UO_1088 (O_1088,N_27225,N_26746);
nand UO_1089 (O_1089,N_29945,N_27277);
or UO_1090 (O_1090,N_25358,N_29881);
nand UO_1091 (O_1091,N_26725,N_29088);
xor UO_1092 (O_1092,N_29400,N_29336);
or UO_1093 (O_1093,N_26949,N_26660);
xor UO_1094 (O_1094,N_26025,N_27741);
nor UO_1095 (O_1095,N_27413,N_27060);
nand UO_1096 (O_1096,N_26899,N_25052);
xor UO_1097 (O_1097,N_25340,N_27077);
xor UO_1098 (O_1098,N_29066,N_25566);
nor UO_1099 (O_1099,N_26455,N_28674);
or UO_1100 (O_1100,N_25458,N_25894);
xor UO_1101 (O_1101,N_29448,N_26407);
xnor UO_1102 (O_1102,N_25928,N_25632);
and UO_1103 (O_1103,N_26680,N_28912);
and UO_1104 (O_1104,N_27619,N_26252);
nand UO_1105 (O_1105,N_25970,N_26513);
nand UO_1106 (O_1106,N_28131,N_27781);
nand UO_1107 (O_1107,N_27303,N_25386);
nand UO_1108 (O_1108,N_28653,N_25535);
xnor UO_1109 (O_1109,N_27428,N_26224);
nand UO_1110 (O_1110,N_26019,N_29562);
or UO_1111 (O_1111,N_29479,N_29685);
and UO_1112 (O_1112,N_29601,N_25809);
nor UO_1113 (O_1113,N_26471,N_26518);
or UO_1114 (O_1114,N_25296,N_27542);
and UO_1115 (O_1115,N_28920,N_27305);
or UO_1116 (O_1116,N_28463,N_29949);
nand UO_1117 (O_1117,N_26467,N_29628);
nand UO_1118 (O_1118,N_27410,N_26519);
or UO_1119 (O_1119,N_28826,N_29114);
nor UO_1120 (O_1120,N_28799,N_26310);
xnor UO_1121 (O_1121,N_27645,N_28621);
and UO_1122 (O_1122,N_28492,N_25407);
nor UO_1123 (O_1123,N_29363,N_27286);
nor UO_1124 (O_1124,N_29941,N_25833);
and UO_1125 (O_1125,N_28429,N_27276);
nor UO_1126 (O_1126,N_27004,N_28983);
and UO_1127 (O_1127,N_29781,N_29787);
nand UO_1128 (O_1128,N_25146,N_25257);
and UO_1129 (O_1129,N_25500,N_29642);
or UO_1130 (O_1130,N_25959,N_26177);
and UO_1131 (O_1131,N_28558,N_28872);
or UO_1132 (O_1132,N_29940,N_25011);
xnor UO_1133 (O_1133,N_28079,N_27824);
and UO_1134 (O_1134,N_28623,N_25932);
nand UO_1135 (O_1135,N_25925,N_26886);
xor UO_1136 (O_1136,N_28033,N_29613);
nor UO_1137 (O_1137,N_26328,N_27242);
or UO_1138 (O_1138,N_25668,N_25468);
nor UO_1139 (O_1139,N_26008,N_27910);
xor UO_1140 (O_1140,N_27185,N_28723);
xor UO_1141 (O_1141,N_28515,N_25772);
and UO_1142 (O_1142,N_26893,N_28681);
and UO_1143 (O_1143,N_26920,N_29955);
nor UO_1144 (O_1144,N_25306,N_28879);
nand UO_1145 (O_1145,N_28477,N_25438);
nor UO_1146 (O_1146,N_26506,N_27698);
or UO_1147 (O_1147,N_26069,N_29866);
nand UO_1148 (O_1148,N_27586,N_25543);
xnor UO_1149 (O_1149,N_25879,N_27887);
nor UO_1150 (O_1150,N_26006,N_28606);
nand UO_1151 (O_1151,N_29737,N_28377);
or UO_1152 (O_1152,N_25919,N_26470);
and UO_1153 (O_1153,N_28889,N_25950);
xnor UO_1154 (O_1154,N_28933,N_28413);
or UO_1155 (O_1155,N_25819,N_27605);
xor UO_1156 (O_1156,N_26190,N_25265);
and UO_1157 (O_1157,N_25373,N_27635);
or UO_1158 (O_1158,N_29721,N_29135);
nor UO_1159 (O_1159,N_26736,N_26751);
and UO_1160 (O_1160,N_27136,N_25145);
xnor UO_1161 (O_1161,N_28842,N_28630);
or UO_1162 (O_1162,N_29671,N_25459);
and UO_1163 (O_1163,N_29290,N_27171);
or UO_1164 (O_1164,N_25995,N_28506);
and UO_1165 (O_1165,N_26498,N_28924);
nand UO_1166 (O_1166,N_28677,N_25094);
nand UO_1167 (O_1167,N_28904,N_25369);
and UO_1168 (O_1168,N_25429,N_28991);
nand UO_1169 (O_1169,N_25700,N_29522);
and UO_1170 (O_1170,N_26830,N_29754);
nand UO_1171 (O_1171,N_26815,N_28022);
or UO_1172 (O_1172,N_28268,N_28381);
nand UO_1173 (O_1173,N_27676,N_28609);
or UO_1174 (O_1174,N_29150,N_26502);
xnor UO_1175 (O_1175,N_27055,N_26695);
nor UO_1176 (O_1176,N_26153,N_28990);
nor UO_1177 (O_1177,N_28571,N_29959);
or UO_1178 (O_1178,N_26798,N_25643);
or UO_1179 (O_1179,N_27794,N_26081);
nand UO_1180 (O_1180,N_27677,N_26794);
or UO_1181 (O_1181,N_25757,N_29240);
or UO_1182 (O_1182,N_27629,N_25370);
nor UO_1183 (O_1183,N_27920,N_29424);
nand UO_1184 (O_1184,N_27570,N_28134);
or UO_1185 (O_1185,N_26883,N_28025);
and UO_1186 (O_1186,N_27739,N_27715);
xor UO_1187 (O_1187,N_25378,N_25570);
xor UO_1188 (O_1188,N_27821,N_25016);
or UO_1189 (O_1189,N_27052,N_26743);
and UO_1190 (O_1190,N_27405,N_25968);
nand UO_1191 (O_1191,N_26927,N_28114);
xnor UO_1192 (O_1192,N_25873,N_25983);
or UO_1193 (O_1193,N_26701,N_25552);
and UO_1194 (O_1194,N_27009,N_26579);
nand UO_1195 (O_1195,N_25371,N_29919);
nor UO_1196 (O_1196,N_25509,N_25312);
nor UO_1197 (O_1197,N_27581,N_26430);
and UO_1198 (O_1198,N_26663,N_28487);
nand UO_1199 (O_1199,N_25949,N_29888);
and UO_1200 (O_1200,N_28602,N_26795);
xor UO_1201 (O_1201,N_25264,N_29842);
xnor UO_1202 (O_1202,N_28650,N_28861);
xor UO_1203 (O_1203,N_28116,N_25508);
nor UO_1204 (O_1204,N_28611,N_27830);
nand UO_1205 (O_1205,N_27260,N_26157);
nand UO_1206 (O_1206,N_25009,N_29810);
nand UO_1207 (O_1207,N_27259,N_27607);
or UO_1208 (O_1208,N_28279,N_28491);
or UO_1209 (O_1209,N_29584,N_28012);
or UO_1210 (O_1210,N_28110,N_26293);
nor UO_1211 (O_1211,N_28835,N_29373);
nor UO_1212 (O_1212,N_26561,N_28614);
and UO_1213 (O_1213,N_27566,N_26040);
or UO_1214 (O_1214,N_26123,N_25957);
nor UO_1215 (O_1215,N_28011,N_27164);
nor UO_1216 (O_1216,N_26479,N_29991);
xor UO_1217 (O_1217,N_28282,N_26163);
xor UO_1218 (O_1218,N_26821,N_29985);
and UO_1219 (O_1219,N_25626,N_26999);
nand UO_1220 (O_1220,N_27802,N_29666);
and UO_1221 (O_1221,N_28498,N_26824);
xor UO_1222 (O_1222,N_29494,N_25317);
and UO_1223 (O_1223,N_27186,N_28813);
or UO_1224 (O_1224,N_29279,N_28998);
nor UO_1225 (O_1225,N_29997,N_26800);
or UO_1226 (O_1226,N_29661,N_29503);
and UO_1227 (O_1227,N_29413,N_29929);
nor UO_1228 (O_1228,N_27973,N_27075);
nor UO_1229 (O_1229,N_29318,N_26591);
nor UO_1230 (O_1230,N_26489,N_29877);
or UO_1231 (O_1231,N_28721,N_27364);
nor UO_1232 (O_1232,N_28180,N_28679);
and UO_1233 (O_1233,N_29709,N_27378);
xnor UO_1234 (O_1234,N_29795,N_27516);
nand UO_1235 (O_1235,N_29094,N_27688);
and UO_1236 (O_1236,N_26337,N_26584);
nor UO_1237 (O_1237,N_25773,N_29343);
or UO_1238 (O_1238,N_29592,N_27487);
or UO_1239 (O_1239,N_27567,N_27966);
xnor UO_1240 (O_1240,N_28857,N_26816);
xor UO_1241 (O_1241,N_27395,N_27740);
or UO_1242 (O_1242,N_25439,N_28767);
or UO_1243 (O_1243,N_29696,N_26892);
xor UO_1244 (O_1244,N_29322,N_28365);
and UO_1245 (O_1245,N_26116,N_29014);
nand UO_1246 (O_1246,N_28294,N_28997);
xnor UO_1247 (O_1247,N_27280,N_26570);
xor UO_1248 (O_1248,N_28244,N_26303);
and UO_1249 (O_1249,N_29031,N_26880);
or UO_1250 (O_1250,N_25416,N_27965);
xor UO_1251 (O_1251,N_26691,N_28837);
nor UO_1252 (O_1252,N_26938,N_27944);
nor UO_1253 (O_1253,N_27151,N_28047);
xnor UO_1254 (O_1254,N_29011,N_26145);
nand UO_1255 (O_1255,N_25665,N_29517);
and UO_1256 (O_1256,N_27959,N_29188);
or UO_1257 (O_1257,N_28476,N_27433);
nand UO_1258 (O_1258,N_26760,N_25047);
nor UO_1259 (O_1259,N_25803,N_29697);
nand UO_1260 (O_1260,N_29936,N_28374);
and UO_1261 (O_1261,N_28233,N_25990);
and UO_1262 (O_1262,N_29144,N_25791);
or UO_1263 (O_1263,N_27820,N_28409);
or UO_1264 (O_1264,N_27349,N_25569);
or UO_1265 (O_1265,N_27593,N_29335);
or UO_1266 (O_1266,N_25855,N_25287);
or UO_1267 (O_1267,N_25792,N_26583);
or UO_1268 (O_1268,N_28593,N_28138);
xor UO_1269 (O_1269,N_27340,N_27103);
or UO_1270 (O_1270,N_25425,N_28423);
nor UO_1271 (O_1271,N_27942,N_27354);
and UO_1272 (O_1272,N_25611,N_25313);
nand UO_1273 (O_1273,N_29568,N_26689);
nand UO_1274 (O_1274,N_29766,N_29355);
nor UO_1275 (O_1275,N_27754,N_27020);
nor UO_1276 (O_1276,N_26964,N_28772);
nor UO_1277 (O_1277,N_27888,N_29198);
nand UO_1278 (O_1278,N_25463,N_27664);
nand UO_1279 (O_1279,N_26450,N_25511);
xor UO_1280 (O_1280,N_28241,N_27997);
xnor UO_1281 (O_1281,N_29830,N_25874);
nand UO_1282 (O_1282,N_27957,N_29040);
xnor UO_1283 (O_1283,N_27809,N_25885);
nor UO_1284 (O_1284,N_29953,N_26184);
nand UO_1285 (O_1285,N_28809,N_28081);
nand UO_1286 (O_1286,N_28553,N_29603);
or UO_1287 (O_1287,N_28336,N_28442);
nand UO_1288 (O_1288,N_29294,N_26881);
and UO_1289 (O_1289,N_26043,N_29609);
nor UO_1290 (O_1290,N_29784,N_26814);
xor UO_1291 (O_1291,N_27867,N_29104);
nand UO_1292 (O_1292,N_25716,N_27489);
nor UO_1293 (O_1293,N_29371,N_28355);
and UO_1294 (O_1294,N_25844,N_25220);
and UO_1295 (O_1295,N_25782,N_25739);
and UO_1296 (O_1296,N_27862,N_28828);
nor UO_1297 (O_1297,N_27424,N_28601);
nor UO_1298 (O_1298,N_27755,N_29352);
and UO_1299 (O_1299,N_25254,N_29667);
xor UO_1300 (O_1300,N_29964,N_25014);
nand UO_1301 (O_1301,N_27734,N_29610);
and UO_1302 (O_1302,N_26269,N_25375);
nand UO_1303 (O_1303,N_29526,N_26055);
nor UO_1304 (O_1304,N_27117,N_26867);
xnor UO_1305 (O_1305,N_26932,N_26290);
or UO_1306 (O_1306,N_29591,N_27673);
and UO_1307 (O_1307,N_27458,N_29537);
nand UO_1308 (O_1308,N_25195,N_27035);
or UO_1309 (O_1309,N_27178,N_26454);
nor UO_1310 (O_1310,N_29792,N_25138);
nor UO_1311 (O_1311,N_27603,N_25042);
nand UO_1312 (O_1312,N_27420,N_29887);
and UO_1313 (O_1313,N_27559,N_26511);
nand UO_1314 (O_1314,N_28166,N_26079);
or UO_1315 (O_1315,N_27076,N_26185);
nor UO_1316 (O_1316,N_26902,N_25537);
nor UO_1317 (O_1317,N_26332,N_28916);
or UO_1318 (O_1318,N_29345,N_28042);
nand UO_1319 (O_1319,N_26620,N_29740);
nor UO_1320 (O_1320,N_26146,N_27964);
nor UO_1321 (O_1321,N_25853,N_27710);
xnor UO_1322 (O_1322,N_28053,N_27348);
or UO_1323 (O_1323,N_28572,N_28345);
xnor UO_1324 (O_1324,N_25940,N_27767);
xnor UO_1325 (O_1325,N_25150,N_27421);
and UO_1326 (O_1326,N_27211,N_26251);
nand UO_1327 (O_1327,N_27215,N_25900);
and UO_1328 (O_1328,N_28538,N_26026);
and UO_1329 (O_1329,N_28326,N_27720);
nand UO_1330 (O_1330,N_26277,N_29659);
nand UO_1331 (O_1331,N_29423,N_26635);
xor UO_1332 (O_1332,N_28501,N_26493);
or UO_1333 (O_1333,N_28740,N_25648);
nor UO_1334 (O_1334,N_28810,N_27346);
xor UO_1335 (O_1335,N_25909,N_26193);
xnor UO_1336 (O_1336,N_29624,N_28117);
nand UO_1337 (O_1337,N_26913,N_25615);
or UO_1338 (O_1338,N_25241,N_27068);
xor UO_1339 (O_1339,N_29121,N_26958);
xor UO_1340 (O_1340,N_26609,N_27706);
nand UO_1341 (O_1341,N_27517,N_29298);
nand UO_1342 (O_1342,N_29402,N_25379);
or UO_1343 (O_1343,N_28260,N_26509);
nor UO_1344 (O_1344,N_25462,N_27157);
nor UO_1345 (O_1345,N_26468,N_27786);
xnor UO_1346 (O_1346,N_25680,N_25811);
xnor UO_1347 (O_1347,N_25122,N_27087);
nor UO_1348 (O_1348,N_26657,N_26340);
nand UO_1349 (O_1349,N_27137,N_29514);
xnor UO_1350 (O_1350,N_25850,N_26137);
or UO_1351 (O_1351,N_25749,N_26073);
or UO_1352 (O_1352,N_27083,N_26057);
nand UO_1353 (O_1353,N_28684,N_26395);
and UO_1354 (O_1354,N_25449,N_26836);
nor UO_1355 (O_1355,N_27027,N_27273);
nor UO_1356 (O_1356,N_29543,N_26878);
and UO_1357 (O_1357,N_27014,N_25002);
nand UO_1358 (O_1358,N_25820,N_28093);
nor UO_1359 (O_1359,N_26658,N_25797);
and UO_1360 (O_1360,N_26159,N_29117);
nor UO_1361 (O_1361,N_26229,N_27764);
or UO_1362 (O_1362,N_25120,N_29814);
or UO_1363 (O_1363,N_29984,N_27998);
and UO_1364 (O_1364,N_26039,N_26174);
nor UO_1365 (O_1365,N_27893,N_27335);
xnor UO_1366 (O_1366,N_28575,N_29695);
nand UO_1367 (O_1367,N_26526,N_26351);
nor UO_1368 (O_1368,N_29418,N_28970);
xnor UO_1369 (O_1369,N_27034,N_29113);
nand UO_1370 (O_1370,N_26037,N_25815);
or UO_1371 (O_1371,N_28853,N_26021);
or UO_1372 (O_1372,N_26951,N_25156);
or UO_1373 (O_1373,N_27149,N_26870);
or UO_1374 (O_1374,N_29589,N_29861);
or UO_1375 (O_1375,N_25079,N_25084);
and UO_1376 (O_1376,N_27113,N_25411);
and UO_1377 (O_1377,N_25255,N_25353);
and UO_1378 (O_1378,N_28443,N_26615);
and UO_1379 (O_1379,N_26013,N_27407);
nor UO_1380 (O_1380,N_29239,N_26114);
and UO_1381 (O_1381,N_26841,N_28644);
xnor UO_1382 (O_1382,N_25913,N_29334);
and UO_1383 (O_1383,N_25764,N_26094);
or UO_1384 (O_1384,N_27592,N_27804);
or UO_1385 (O_1385,N_26884,N_29030);
or UO_1386 (O_1386,N_29525,N_25594);
xor UO_1387 (O_1387,N_29824,N_28783);
xor UO_1388 (O_1388,N_28359,N_25289);
nand UO_1389 (O_1389,N_29487,N_28386);
and UO_1390 (O_1390,N_28013,N_25319);
or UO_1391 (O_1391,N_28141,N_26203);
nand UO_1392 (O_1392,N_26722,N_27084);
or UO_1393 (O_1393,N_27069,N_25868);
xor UO_1394 (O_1394,N_29644,N_27969);
and UO_1395 (O_1395,N_26517,N_29808);
nor UO_1396 (O_1396,N_27961,N_25799);
nor UO_1397 (O_1397,N_29396,N_26371);
and UO_1398 (O_1398,N_29061,N_29131);
and UO_1399 (O_1399,N_26264,N_29044);
nand UO_1400 (O_1400,N_27614,N_26158);
xor UO_1401 (O_1401,N_28320,N_26065);
nand UO_1402 (O_1402,N_28789,N_29405);
or UO_1403 (O_1403,N_27707,N_28329);
nor UO_1404 (O_1404,N_29340,N_25507);
nor UO_1405 (O_1405,N_28216,N_27301);
or UO_1406 (O_1406,N_29856,N_26148);
or UO_1407 (O_1407,N_29372,N_29579);
or UO_1408 (O_1408,N_28668,N_26861);
nor UO_1409 (O_1409,N_28148,N_28146);
nor UO_1410 (O_1410,N_28069,N_27658);
nand UO_1411 (O_1411,N_28309,N_28283);
or UO_1412 (O_1412,N_29331,N_26175);
and UO_1413 (O_1413,N_26835,N_26621);
and UO_1414 (O_1414,N_29404,N_25771);
and UO_1415 (O_1415,N_27766,N_27057);
and UO_1416 (O_1416,N_25839,N_27448);
nand UO_1417 (O_1417,N_26690,N_25692);
and UO_1418 (O_1418,N_29118,N_25687);
nand UO_1419 (O_1419,N_25447,N_28038);
nor UO_1420 (O_1420,N_28903,N_25993);
or UO_1421 (O_1421,N_29415,N_25941);
and UO_1422 (O_1422,N_26555,N_25399);
nor UO_1423 (O_1423,N_27238,N_27063);
nand UO_1424 (O_1424,N_25311,N_26268);
or UO_1425 (O_1425,N_27627,N_28648);
nor UO_1426 (O_1426,N_25041,N_28214);
xor UO_1427 (O_1427,N_25984,N_27713);
and UO_1428 (O_1428,N_27339,N_26779);
nor UO_1429 (O_1429,N_26503,N_29055);
nand UO_1430 (O_1430,N_26346,N_27104);
nand UO_1431 (O_1431,N_26087,N_29428);
or UO_1432 (O_1432,N_27935,N_27232);
nor UO_1433 (O_1433,N_29398,N_26112);
nand UO_1434 (O_1434,N_29674,N_25320);
nor UO_1435 (O_1435,N_27595,N_28295);
or UO_1436 (O_1436,N_29186,N_27423);
and UO_1437 (O_1437,N_25070,N_27430);
nor UO_1438 (O_1438,N_26853,N_28307);
or UO_1439 (O_1439,N_26160,N_26036);
or UO_1440 (O_1440,N_27528,N_27502);
and UO_1441 (O_1441,N_29558,N_25088);
xnor UO_1442 (O_1442,N_26739,N_26837);
nor UO_1443 (O_1443,N_27812,N_29819);
nand UO_1444 (O_1444,N_26178,N_27896);
xor UO_1445 (O_1445,N_26044,N_28145);
nand UO_1446 (O_1446,N_27808,N_29456);
nor UO_1447 (O_1447,N_29283,N_25956);
xnor UO_1448 (O_1448,N_28428,N_29348);
nor UO_1449 (O_1449,N_28331,N_28132);
or UO_1450 (O_1450,N_29330,N_27338);
nor UO_1451 (O_1451,N_26230,N_27322);
nand UO_1452 (O_1452,N_26367,N_25434);
nand UO_1453 (O_1453,N_28002,N_28944);
or UO_1454 (O_1454,N_27003,N_28255);
nand UO_1455 (O_1455,N_27312,N_27425);
nor UO_1456 (O_1456,N_27408,N_25945);
xnor UO_1457 (O_1457,N_29454,N_25914);
or UO_1458 (O_1458,N_25389,N_25401);
nand UO_1459 (O_1459,N_28946,N_25790);
and UO_1460 (O_1460,N_28055,N_29060);
and UO_1461 (O_1461,N_27937,N_26129);
and UO_1462 (O_1462,N_25098,N_29643);
and UO_1463 (O_1463,N_28969,N_28482);
nor UO_1464 (O_1464,N_29098,N_28993);
or UO_1465 (O_1465,N_27525,N_26301);
nor UO_1466 (O_1466,N_26515,N_28881);
nor UO_1467 (O_1467,N_25502,N_29771);
or UO_1468 (O_1468,N_29714,N_27803);
or UO_1469 (O_1469,N_27618,N_29509);
xor UO_1470 (O_1470,N_26866,N_27894);
xnor UO_1471 (O_1471,N_27097,N_27857);
nor UO_1472 (O_1472,N_29539,N_26914);
and UO_1473 (O_1473,N_29395,N_28121);
and UO_1474 (O_1474,N_27522,N_28757);
xor UO_1475 (O_1475,N_26898,N_25759);
xor UO_1476 (O_1476,N_28883,N_26329);
nand UO_1477 (O_1477,N_25316,N_27654);
and UO_1478 (O_1478,N_29895,N_28500);
nand UO_1479 (O_1479,N_27024,N_28137);
or UO_1480 (O_1480,N_27863,N_29397);
nand UO_1481 (O_1481,N_27838,N_27899);
xor UO_1482 (O_1482,N_25391,N_25436);
xor UO_1483 (O_1483,N_25527,N_26966);
nand UO_1484 (O_1484,N_29850,N_27879);
xor UO_1485 (O_1485,N_26655,N_25293);
nand UO_1486 (O_1486,N_28974,N_28739);
nor UO_1487 (O_1487,N_26682,N_29216);
xnor UO_1488 (O_1488,N_25364,N_25210);
nand UO_1489 (O_1489,N_25802,N_29003);
nand UO_1490 (O_1490,N_29548,N_26461);
nand UO_1491 (O_1491,N_28152,N_28366);
or UO_1492 (O_1492,N_26527,N_27881);
nor UO_1493 (O_1493,N_28126,N_28535);
and UO_1494 (O_1494,N_29711,N_25592);
nor UO_1495 (O_1495,N_29701,N_27041);
nor UO_1496 (O_1496,N_29635,N_26242);
xor UO_1497 (O_1497,N_26131,N_28761);
xor UO_1498 (O_1498,N_28402,N_28461);
nand UO_1499 (O_1499,N_28133,N_26317);
nand UO_1500 (O_1500,N_25723,N_25966);
or UO_1501 (O_1501,N_28205,N_25501);
and UO_1502 (O_1502,N_27727,N_26319);
or UO_1503 (O_1503,N_28113,N_28425);
nand UO_1504 (O_1504,N_26015,N_28242);
nand UO_1505 (O_1505,N_27172,N_29563);
nor UO_1506 (O_1506,N_29103,N_28565);
nand UO_1507 (O_1507,N_25768,N_28410);
nor UO_1508 (O_1508,N_29723,N_29791);
and UO_1509 (O_1509,N_26197,N_27638);
nand UO_1510 (O_1510,N_27625,N_26439);
nor UO_1511 (O_1511,N_26431,N_25731);
and UO_1512 (O_1512,N_25800,N_27597);
or UO_1513 (O_1513,N_28762,N_28503);
xnor UO_1514 (O_1514,N_29443,N_29478);
nand UO_1515 (O_1515,N_28760,N_29670);
nand UO_1516 (O_1516,N_25387,N_27610);
nor UO_1517 (O_1517,N_29297,N_29504);
nand UO_1518 (O_1518,N_26338,N_28466);
nand UO_1519 (O_1519,N_27132,N_29006);
nand UO_1520 (O_1520,N_26496,N_27333);
nand UO_1521 (O_1521,N_29566,N_29164);
or UO_1522 (O_1522,N_29614,N_26139);
nand UO_1523 (O_1523,N_28389,N_27967);
nor UO_1524 (O_1524,N_27839,N_28179);
and UO_1525 (O_1525,N_26728,N_26797);
nand UO_1526 (O_1526,N_26945,N_29855);
nand UO_1527 (O_1527,N_29142,N_26589);
nor UO_1528 (O_1528,N_29038,N_29466);
or UO_1529 (O_1529,N_27123,N_26050);
or UO_1530 (O_1530,N_28736,N_25023);
nor UO_1531 (O_1531,N_27933,N_28805);
or UO_1532 (O_1532,N_28082,N_25575);
or UO_1533 (O_1533,N_27418,N_28951);
nand UO_1534 (O_1534,N_27175,N_28880);
or UO_1535 (O_1535,N_29629,N_29230);
and UO_1536 (O_1536,N_26099,N_28935);
nand UO_1537 (O_1537,N_28218,N_29549);
or UO_1538 (O_1538,N_27521,N_28395);
nand UO_1539 (O_1539,N_28390,N_27960);
xnor UO_1540 (O_1540,N_25513,N_26226);
nor UO_1541 (O_1541,N_26857,N_26772);
xnor UO_1542 (O_1542,N_26032,N_29574);
xnor UO_1543 (O_1543,N_25600,N_28637);
and UO_1544 (O_1544,N_27785,N_25077);
and UO_1545 (O_1545,N_29561,N_27490);
or UO_1546 (O_1546,N_25112,N_28447);
and UO_1547 (O_1547,N_27630,N_29823);
nand UO_1548 (O_1548,N_26210,N_28823);
xnor UO_1549 (O_1549,N_28573,N_29611);
nor UO_1550 (O_1550,N_26382,N_27023);
nand UO_1551 (O_1551,N_25746,N_29191);
or UO_1552 (O_1552,N_28057,N_29767);
xnor UO_1553 (O_1553,N_29863,N_27114);
nand UO_1554 (O_1554,N_27904,N_29022);
and UO_1555 (O_1555,N_25213,N_26173);
nor UO_1556 (O_1556,N_25695,N_28031);
and UO_1557 (O_1557,N_29134,N_25227);
and UO_1558 (O_1558,N_27257,N_27687);
and UO_1559 (O_1559,N_27457,N_26769);
xnor UO_1560 (O_1560,N_25714,N_25977);
nor UO_1561 (O_1561,N_27220,N_25816);
xor UO_1562 (O_1562,N_27511,N_27574);
nor UO_1563 (O_1563,N_25491,N_28830);
xnor UO_1564 (O_1564,N_29871,N_27911);
nand UO_1565 (O_1565,N_27212,N_26524);
nand UO_1566 (O_1566,N_29169,N_25395);
nor UO_1567 (O_1567,N_26592,N_27002);
and UO_1568 (O_1568,N_27105,N_25823);
nand UO_1569 (O_1569,N_25733,N_26731);
xnor UO_1570 (O_1570,N_27042,N_29225);
or UO_1571 (O_1571,N_26566,N_27152);
or UO_1572 (O_1572,N_25777,N_28039);
nor UO_1573 (O_1573,N_28208,N_25410);
and UO_1574 (O_1574,N_28627,N_25367);
nand UO_1575 (O_1575,N_28328,N_29617);
and UO_1576 (O_1576,N_25514,N_28330);
nor UO_1577 (O_1577,N_26813,N_29302);
xor UO_1578 (O_1578,N_29715,N_26718);
nand UO_1579 (O_1579,N_26238,N_27805);
and UO_1580 (O_1580,N_25057,N_28051);
nor UO_1581 (O_1581,N_29242,N_27241);
or UO_1582 (O_1582,N_28494,N_27970);
nand UO_1583 (O_1583,N_27099,N_27553);
nand UO_1584 (O_1584,N_29333,N_29384);
nand UO_1585 (O_1585,N_25858,N_27124);
nor UO_1586 (O_1586,N_28262,N_28250);
or UO_1587 (O_1587,N_25893,N_27016);
nand UO_1588 (O_1588,N_25419,N_25567);
nand UO_1589 (O_1589,N_28027,N_28106);
or UO_1590 (O_1590,N_27653,N_25650);
and UO_1591 (O_1591,N_25546,N_25489);
or UO_1592 (O_1592,N_27039,N_26389);
xnor UO_1593 (O_1593,N_26543,N_29411);
nand UO_1594 (O_1594,N_29375,N_29441);
and UO_1595 (O_1595,N_28269,N_25297);
and UO_1596 (O_1596,N_25262,N_25355);
xor UO_1597 (O_1597,N_26712,N_25701);
or UO_1598 (O_1598,N_28766,N_25999);
xnor UO_1599 (O_1599,N_28522,N_28321);
nand UO_1600 (O_1600,N_27223,N_26787);
nor UO_1601 (O_1601,N_29219,N_27527);
nand UO_1602 (O_1602,N_29957,N_26170);
xnor UO_1603 (O_1603,N_28176,N_26408);
and UO_1604 (O_1604,N_28928,N_29133);
nor UO_1605 (O_1605,N_27848,N_28811);
nor UO_1606 (O_1606,N_26472,N_29110);
nor UO_1607 (O_1607,N_28020,N_26601);
nor UO_1608 (O_1608,N_26362,N_25256);
and UO_1609 (O_1609,N_29206,N_28436);
nor UO_1610 (O_1610,N_29502,N_25400);
and UO_1611 (O_1611,N_27207,N_29080);
nand UO_1612 (O_1612,N_29105,N_29123);
xnor UO_1613 (O_1613,N_26804,N_26823);
xor UO_1614 (O_1614,N_29299,N_26485);
nand UO_1615 (O_1615,N_28981,N_29076);
or UO_1616 (O_1616,N_29802,N_27341);
and UO_1617 (O_1617,N_28954,N_28251);
xnor UO_1618 (O_1618,N_29203,N_25953);
xnor UO_1619 (O_1619,N_29803,N_27519);
and UO_1620 (O_1620,N_26298,N_25441);
nand UO_1621 (O_1621,N_29529,N_28373);
nand UO_1622 (O_1622,N_26553,N_28404);
xor UO_1623 (O_1623,N_27534,N_26240);
nand UO_1624 (O_1624,N_26120,N_26199);
or UO_1625 (O_1625,N_25250,N_28061);
nor UO_1626 (O_1626,N_27255,N_29037);
xnor UO_1627 (O_1627,N_28688,N_29338);
or UO_1628 (O_1628,N_26926,N_29694);
xor UO_1629 (O_1629,N_29483,N_26581);
and UO_1630 (O_1630,N_26525,N_28923);
and UO_1631 (O_1631,N_25629,N_26551);
and UO_1632 (O_1632,N_28297,N_26483);
xor UO_1633 (O_1633,N_26563,N_28656);
or UO_1634 (O_1634,N_29024,N_25583);
and UO_1635 (O_1635,N_25624,N_25078);
nand UO_1636 (O_1636,N_28032,N_27066);
and UO_1637 (O_1637,N_29147,N_26593);
or UO_1638 (O_1638,N_29755,N_27613);
or UO_1639 (O_1639,N_27986,N_27813);
or UO_1640 (O_1640,N_25862,N_28622);
nand UO_1641 (O_1641,N_26161,N_28237);
and UO_1642 (O_1642,N_28206,N_26045);
nand UO_1643 (O_1643,N_28673,N_28308);
nand UO_1644 (O_1644,N_27062,N_26844);
and UO_1645 (O_1645,N_29490,N_25517);
or UO_1646 (O_1646,N_25018,N_29329);
xor UO_1647 (O_1647,N_29627,N_25271);
xnor UO_1648 (O_1648,N_26753,N_26871);
or UO_1649 (O_1649,N_25614,N_25830);
or UO_1650 (O_1650,N_27875,N_26752);
xnor UO_1651 (O_1651,N_27131,N_27323);
nor UO_1652 (O_1652,N_27756,N_26490);
and UO_1653 (O_1653,N_25817,N_25916);
or UO_1654 (O_1654,N_29656,N_28227);
or UO_1655 (O_1655,N_27716,N_28219);
or UO_1656 (O_1656,N_25124,N_29277);
and UO_1657 (O_1657,N_28187,N_28239);
and UO_1658 (O_1658,N_28469,N_26889);
nand UO_1659 (O_1659,N_26464,N_25137);
nor UO_1660 (O_1660,N_26012,N_26423);
and UO_1661 (O_1661,N_25330,N_29438);
and UO_1662 (O_1662,N_26447,N_25503);
xnor UO_1663 (O_1663,N_25376,N_26727);
and UO_1664 (O_1664,N_28245,N_25141);
or UO_1665 (O_1665,N_25715,N_28439);
nand UO_1666 (O_1666,N_26271,N_29621);
nand UO_1667 (O_1667,N_29638,N_25231);
or UO_1668 (O_1668,N_26091,N_29064);
nor UO_1669 (O_1669,N_25836,N_25440);
nand UO_1670 (O_1670,N_26777,N_25294);
nand UO_1671 (O_1671,N_26758,N_28800);
nor UO_1672 (O_1672,N_26757,N_25523);
nand UO_1673 (O_1673,N_26009,N_29276);
nor UO_1674 (O_1674,N_27272,N_26594);
nand UO_1675 (O_1675,N_27040,N_25314);
xor UO_1676 (O_1676,N_25290,N_26014);
and UO_1677 (O_1677,N_25506,N_29228);
or UO_1678 (O_1678,N_28698,N_27229);
or UO_1679 (O_1679,N_28458,N_27622);
and UO_1680 (O_1680,N_25743,N_28263);
or UO_1681 (O_1681,N_26642,N_25548);
nand UO_1682 (O_1682,N_25133,N_26929);
nand UO_1683 (O_1683,N_25616,N_25656);
nand UO_1684 (O_1684,N_27344,N_29075);
nor UO_1685 (O_1685,N_29554,N_26274);
or UO_1686 (O_1686,N_29019,N_25557);
or UO_1687 (O_1687,N_27643,N_29633);
nor UO_1688 (O_1688,N_27387,N_27864);
or UO_1689 (O_1689,N_26142,N_28908);
nor UO_1690 (O_1690,N_26383,N_25001);
nand UO_1691 (O_1691,N_27366,N_25192);
nor UO_1692 (O_1692,N_29962,N_27922);
or UO_1693 (O_1693,N_27886,N_27753);
xnor UO_1694 (O_1694,N_28686,N_26412);
nand UO_1695 (O_1695,N_28058,N_26172);
or UO_1696 (O_1696,N_28667,N_29136);
nor UO_1697 (O_1697,N_26768,N_27779);
xnor UO_1698 (O_1698,N_27085,N_25308);
or UO_1699 (O_1699,N_26386,N_29050);
or UO_1700 (O_1700,N_25525,N_29465);
nor UO_1701 (O_1701,N_29534,N_25487);
and UO_1702 (O_1702,N_29100,N_28820);
or UO_1703 (O_1703,N_25494,N_28516);
and UO_1704 (O_1704,N_25880,N_28911);
xnor UO_1705 (O_1705,N_27347,N_26980);
nand UO_1706 (O_1706,N_27817,N_27943);
or UO_1707 (O_1707,N_29389,N_29744);
xnor UO_1708 (O_1708,N_25545,N_29310);
and UO_1709 (O_1709,N_29172,N_29835);
nor UO_1710 (O_1710,N_28814,N_26850);
or UO_1711 (O_1711,N_28685,N_25588);
and UO_1712 (O_1712,N_28915,N_26970);
or UO_1713 (O_1713,N_25357,N_25720);
and UO_1714 (O_1714,N_29639,N_25012);
nand UO_1715 (O_1715,N_25741,N_26107);
or UO_1716 (O_1716,N_28832,N_29173);
and UO_1717 (O_1717,N_29085,N_26076);
nor UO_1718 (O_1718,N_25035,N_28177);
and UO_1719 (O_1719,N_25062,N_27506);
or UO_1720 (O_1720,N_28367,N_26266);
and UO_1721 (O_1721,N_27871,N_26872);
and UO_1722 (O_1722,N_28052,N_25303);
xor UO_1723 (O_1723,N_27200,N_29182);
nand UO_1724 (O_1724,N_26783,N_26599);
and UO_1725 (O_1725,N_25278,N_25516);
and UO_1726 (O_1726,N_28769,N_28424);
or UO_1727 (O_1727,N_28085,N_26953);
nor UO_1728 (O_1728,N_29419,N_28554);
or UO_1729 (O_1729,N_28646,N_29232);
nand UO_1730 (O_1730,N_25225,N_25433);
xnor UO_1731 (O_1731,N_27850,N_25253);
or UO_1732 (O_1732,N_26416,N_27743);
nand UO_1733 (O_1733,N_29763,N_25248);
nor UO_1734 (O_1734,N_29362,N_26253);
xnor UO_1735 (O_1735,N_28315,N_28419);
or UO_1736 (O_1736,N_27876,N_28488);
or UO_1737 (O_1737,N_26873,N_26604);
or UO_1738 (O_1738,N_26649,N_26415);
xnor UO_1739 (O_1739,N_28985,N_27370);
xnor UO_1740 (O_1740,N_29091,N_25107);
and UO_1741 (O_1741,N_25424,N_28787);
or UO_1742 (O_1742,N_27994,N_25974);
xor UO_1743 (O_1743,N_29565,N_25991);
nand UO_1744 (O_1744,N_27187,N_28530);
or UO_1745 (O_1745,N_26987,N_28189);
and UO_1746 (O_1746,N_29995,N_26831);
or UO_1747 (O_1747,N_25828,N_25119);
and UO_1748 (O_1748,N_29261,N_26151);
or UO_1749 (O_1749,N_25114,N_25152);
nand UO_1750 (O_1750,N_25221,N_29271);
xor UO_1751 (O_1751,N_29879,N_28770);
and UO_1752 (O_1752,N_28147,N_27367);
nand UO_1753 (O_1753,N_25781,N_26064);
xor UO_1754 (O_1754,N_28198,N_29293);
and UO_1755 (O_1755,N_28958,N_26368);
xor UO_1756 (O_1756,N_29839,N_29205);
nor UO_1757 (O_1757,N_29284,N_28705);
xor UO_1758 (O_1758,N_27095,N_26034);
nand UO_1759 (O_1759,N_26715,N_25975);
and UO_1760 (O_1760,N_29184,N_29096);
or UO_1761 (O_1761,N_28457,N_27996);
or UO_1762 (O_1762,N_26631,N_26354);
or UO_1763 (O_1763,N_25246,N_28370);
xor UO_1764 (O_1764,N_28718,N_25277);
nand UO_1765 (O_1765,N_25396,N_28959);
nand UO_1766 (O_1766,N_28963,N_29654);
nor UO_1767 (O_1767,N_25810,N_25200);
nand UO_1768 (O_1768,N_26460,N_27777);
and UO_1769 (O_1769,N_28394,N_28589);
nand UO_1770 (O_1770,N_26098,N_26399);
nor UO_1771 (O_1771,N_26421,N_27118);
and UO_1772 (O_1772,N_25153,N_27768);
nand UO_1773 (O_1773,N_26458,N_25302);
nand UO_1774 (O_1774,N_28102,N_29773);
nand UO_1775 (O_1775,N_28596,N_29673);
xnor UO_1776 (O_1776,N_29381,N_28310);
nand UO_1777 (O_1777,N_29841,N_25274);
or UO_1778 (O_1778,N_25335,N_29036);
xor UO_1779 (O_1779,N_27150,N_25586);
xnor UO_1780 (O_1780,N_25883,N_29250);
or UO_1781 (O_1781,N_25901,N_25163);
or UO_1782 (O_1782,N_27204,N_27913);
nand UO_1783 (O_1783,N_27948,N_26636);
nor UO_1784 (O_1784,N_26372,N_29827);
nand UO_1785 (O_1785,N_27183,N_26992);
or UO_1786 (O_1786,N_26136,N_29209);
nor UO_1787 (O_1787,N_29112,N_28350);
nand UO_1788 (O_1788,N_25549,N_29777);
xnor UO_1789 (O_1789,N_25258,N_27389);
or UO_1790 (O_1790,N_25394,N_29619);
nor UO_1791 (O_1791,N_29690,N_25574);
or UO_1792 (O_1792,N_25935,N_25464);
and UO_1793 (O_1793,N_26390,N_26198);
and UO_1794 (O_1794,N_26484,N_25338);
nand UO_1795 (O_1795,N_27978,N_26738);
and UO_1796 (O_1796,N_27056,N_27165);
or UO_1797 (O_1797,N_26031,N_29560);
xnor UO_1798 (O_1798,N_29765,N_26380);
nand UO_1799 (O_1799,N_28703,N_29257);
nand UO_1800 (O_1800,N_28694,N_28938);
or UO_1801 (O_1801,N_29426,N_25631);
or UO_1802 (O_1802,N_25697,N_27485);
xor UO_1803 (O_1803,N_26385,N_25576);
and UO_1804 (O_1804,N_26538,N_26182);
and UO_1805 (O_1805,N_26846,N_26826);
nand UO_1806 (O_1806,N_26799,N_28344);
and UO_1807 (O_1807,N_25361,N_28280);
nand UO_1808 (O_1808,N_25207,N_26477);
nand UO_1809 (O_1809,N_26605,N_29386);
and UO_1810 (O_1810,N_27742,N_27070);
or UO_1811 (O_1811,N_28691,N_25808);
xor UO_1812 (O_1812,N_26350,N_25004);
xor UO_1813 (O_1813,N_25304,N_26849);
and UO_1814 (O_1814,N_26782,N_25096);
nor UO_1815 (O_1815,N_25526,N_28897);
or UO_1816 (O_1816,N_26465,N_29035);
nand UO_1817 (O_1817,N_26716,N_29427);
xor UO_1818 (O_1818,N_27291,N_26345);
xor UO_1819 (O_1819,N_28910,N_26105);
xor UO_1820 (O_1820,N_28870,N_28590);
nand UO_1821 (O_1821,N_27731,N_27222);
or UO_1822 (O_1822,N_28502,N_26603);
xor UO_1823 (O_1823,N_27890,N_26366);
or UO_1824 (O_1824,N_25180,N_27170);
or UO_1825 (O_1825,N_28064,N_28164);
and UO_1826 (O_1826,N_27326,N_25305);
nor UO_1827 (O_1827,N_26939,N_29825);
xor UO_1828 (O_1828,N_28305,N_29801);
nand UO_1829 (O_1829,N_25479,N_27526);
xnor UO_1830 (O_1830,N_27078,N_27051);
nand UO_1831 (O_1831,N_25635,N_26969);
xor UO_1832 (O_1832,N_26600,N_26569);
nor UO_1833 (O_1833,N_27361,N_27541);
nor UO_1834 (O_1834,N_29451,N_29032);
nand UO_1835 (O_1835,N_26834,N_29289);
xor UO_1836 (O_1836,N_28235,N_29687);
xor UO_1837 (O_1837,N_26672,N_26111);
and UO_1838 (O_1838,N_25903,N_29047);
xnor UO_1839 (O_1839,N_26916,N_25852);
nand UO_1840 (O_1840,N_25247,N_28257);
xnor UO_1841 (O_1841,N_28804,N_26272);
nor UO_1842 (O_1842,N_28792,N_28574);
nand UO_1843 (O_1843,N_25185,N_27719);
nand UO_1844 (O_1844,N_29406,N_25473);
nor UO_1845 (O_1845,N_28332,N_26223);
nand UO_1846 (O_1846,N_25242,N_27156);
nand UO_1847 (O_1847,N_26552,N_29268);
and UO_1848 (O_1848,N_26887,N_29119);
or UO_1849 (O_1849,N_26840,N_25115);
or UO_1850 (O_1850,N_26626,N_26080);
xor UO_1851 (O_1851,N_26972,N_28775);
nand UO_1852 (O_1852,N_28793,N_29648);
and UO_1853 (O_1853,N_29806,N_25699);
nor UO_1854 (O_1854,N_25164,N_25544);
nor UO_1855 (O_1855,N_26082,N_29309);
nand UO_1856 (O_1856,N_27130,N_28435);
and UO_1857 (O_1857,N_26356,N_26829);
xnor UO_1858 (O_1858,N_28490,N_27319);
nor UO_1859 (O_1859,N_28751,N_29339);
xnor UO_1860 (O_1860,N_26784,N_28044);
or UO_1861 (O_1861,N_27270,N_28303);
nand UO_1862 (O_1862,N_27036,N_29281);
nor UO_1863 (O_1863,N_27507,N_26138);
xor UO_1864 (O_1864,N_28821,N_28831);
nor UO_1865 (O_1865,N_27606,N_27411);
or UO_1866 (O_1866,N_27110,N_29672);
or UO_1867 (O_1867,N_29048,N_26833);
and UO_1868 (O_1868,N_28547,N_27562);
nand UO_1869 (O_1869,N_25270,N_29876);
or UO_1870 (O_1870,N_25206,N_29903);
or UO_1871 (O_1871,N_25878,N_25997);
xnor UO_1872 (O_1872,N_27483,N_27353);
or UO_1873 (O_1873,N_25125,N_29796);
nand UO_1874 (O_1874,N_26748,N_25388);
and UO_1875 (O_1875,N_25898,N_28891);
nand UO_1876 (O_1876,N_29265,N_28634);
xor UO_1877 (O_1877,N_28934,N_25876);
xnor UO_1878 (O_1878,N_29979,N_28375);
nand UO_1879 (O_1879,N_26106,N_26983);
or UO_1880 (O_1880,N_25069,N_28188);
nor UO_1881 (O_1881,N_25580,N_29645);
or UO_1882 (O_1882,N_26469,N_26220);
or UO_1883 (O_1883,N_29547,N_27190);
and UO_1884 (O_1884,N_27202,N_29698);
nor UO_1885 (O_1885,N_27288,N_25542);
and UO_1886 (O_1886,N_25599,N_28988);
xor UO_1887 (O_1887,N_26713,N_29264);
and UO_1888 (O_1888,N_29507,N_29231);
nand UO_1889 (O_1889,N_25275,N_27050);
xnor UO_1890 (O_1890,N_26341,N_27626);
xnor UO_1891 (O_1891,N_27873,N_26629);
and UO_1892 (O_1892,N_29515,N_25587);
or UO_1893 (O_1893,N_28372,N_27360);
nand UO_1894 (O_1894,N_27918,N_27311);
or UO_1895 (O_1895,N_28521,N_26827);
nand UO_1896 (O_1896,N_28919,N_25702);
xor UO_1897 (O_1897,N_28564,N_27917);
nand UO_1898 (O_1898,N_25160,N_27496);
nor UO_1899 (O_1899,N_25581,N_29910);
xnor UO_1900 (O_1900,N_29495,N_28479);
nand UO_1901 (O_1901,N_27479,N_25902);
and UO_1902 (O_1902,N_28405,N_26904);
xor UO_1903 (O_1903,N_26516,N_26542);
nor UO_1904 (O_1904,N_27294,N_29043);
nor UO_1905 (O_1905,N_27853,N_29704);
nor UO_1906 (O_1906,N_25281,N_26092);
or UO_1907 (O_1907,N_26825,N_27422);
nor UO_1908 (O_1908,N_26241,N_29944);
xor UO_1909 (O_1909,N_26327,N_27140);
xnor UO_1910 (O_1910,N_27369,N_29145);
and UO_1911 (O_1911,N_28312,N_26084);
nor UO_1912 (O_1912,N_25383,N_27112);
xor UO_1913 (O_1913,N_25245,N_26233);
nand UO_1914 (O_1914,N_28636,N_27568);
nor UO_1915 (O_1915,N_28514,N_27860);
nor UO_1916 (O_1916,N_26440,N_27022);
and UO_1917 (O_1917,N_26747,N_25327);
and UO_1918 (O_1918,N_29062,N_25551);
xnor UO_1919 (O_1919,N_28863,N_29430);
and UO_1920 (O_1920,N_25334,N_27578);
or UO_1921 (O_1921,N_26413,N_26901);
and UO_1922 (O_1922,N_27096,N_29312);
nor UO_1923 (O_1923,N_25036,N_25996);
nor UO_1924 (O_1924,N_25061,N_25579);
or UO_1925 (O_1925,N_26564,N_29379);
nor UO_1926 (O_1926,N_26004,N_28632);
nand UO_1927 (O_1927,N_27300,N_29759);
nor UO_1928 (O_1928,N_26963,N_29918);
xor UO_1929 (O_1929,N_29712,N_27555);
nand UO_1930 (O_1930,N_28099,N_25235);
xor UO_1931 (O_1931,N_27208,N_28756);
nand UO_1932 (O_1932,N_26443,N_26595);
xor UO_1933 (O_1933,N_27463,N_25691);
xnor UO_1934 (O_1934,N_29189,N_28587);
and UO_1935 (O_1935,N_28876,N_27694);
xnor UO_1936 (O_1936,N_27129,N_26906);
nor UO_1937 (O_1937,N_26089,N_28838);
nand UO_1938 (O_1938,N_29439,N_26679);
and UO_1939 (O_1939,N_28719,N_28882);
nor UO_1940 (O_1940,N_28603,N_28387);
or UO_1941 (O_1941,N_25301,N_25089);
nor UO_1942 (O_1942,N_25994,N_26888);
and UO_1943 (O_1943,N_28304,N_25712);
nor UO_1944 (O_1944,N_27919,N_27840);
and UO_1945 (O_1945,N_28140,N_25972);
or UO_1946 (O_1946,N_29272,N_26523);
xor UO_1947 (O_1947,N_27380,N_26030);
and UO_1948 (O_1948,N_29489,N_27733);
nor UO_1949 (O_1949,N_29474,N_29410);
or UO_1950 (O_1950,N_27293,N_26575);
nand UO_1951 (O_1951,N_29059,N_25605);
nand UO_1952 (O_1952,N_27828,N_28557);
and UO_1953 (O_1953,N_25642,N_26228);
nand UO_1954 (O_1954,N_28773,N_25662);
nor UO_1955 (O_1955,N_25171,N_27094);
xnor UO_1956 (O_1956,N_26671,N_27182);
and UO_1957 (O_1957,N_27661,N_25846);
or UO_1958 (O_1958,N_28306,N_27298);
xor UO_1959 (O_1959,N_29021,N_27772);
xor UO_1960 (O_1960,N_25835,N_26950);
and UO_1961 (O_1961,N_25343,N_26796);
or UO_1962 (O_1962,N_26744,N_25553);
nor UO_1963 (O_1963,N_25006,N_26573);
xnor UO_1964 (O_1964,N_25713,N_29812);
and UO_1965 (O_1965,N_26638,N_28965);
nor UO_1966 (O_1966,N_25488,N_27351);
nor UO_1967 (O_1967,N_28665,N_28351);
nor UO_1968 (O_1968,N_27674,N_28629);
and UO_1969 (O_1969,N_25426,N_25742);
xor UO_1970 (O_1970,N_26487,N_26530);
nand UO_1971 (O_1971,N_25895,N_25295);
or UO_1972 (O_1972,N_28600,N_25603);
or UO_1973 (O_1973,N_27393,N_25093);
nor UO_1974 (O_1974,N_26562,N_29907);
xor UO_1975 (O_1975,N_25751,N_25005);
xor UO_1976 (O_1976,N_27885,N_26320);
and UO_1977 (O_1977,N_25992,N_25034);
nor UO_1978 (O_1978,N_25485,N_27549);
or UO_1979 (O_1979,N_25113,N_28437);
or UO_1980 (O_1980,N_29857,N_29882);
and UO_1981 (O_1981,N_27189,N_27659);
and UO_1982 (O_1982,N_25451,N_26917);
or UO_1983 (O_1983,N_28854,N_25660);
xnor UO_1984 (O_1984,N_28894,N_27726);
or UO_1985 (O_1985,N_26641,N_29421);
and UO_1986 (O_1986,N_29932,N_27547);
nor UO_1987 (O_1987,N_25998,N_29741);
and UO_1988 (O_1988,N_28271,N_27861);
and UO_1989 (O_1989,N_28451,N_29772);
or UO_1990 (O_1990,N_26283,N_25461);
nor UO_1991 (O_1991,N_27184,N_28984);
nand UO_1992 (O_1992,N_27765,N_26737);
and UO_1993 (O_1993,N_28352,N_25840);
xnor UO_1994 (O_1994,N_28173,N_27403);
nand UO_1995 (O_1995,N_28528,N_27486);
nand UO_1996 (O_1996,N_29652,N_29899);
and UO_1997 (O_1997,N_25186,N_27573);
nand UO_1998 (O_1998,N_29175,N_29583);
and UO_1999 (O_1999,N_29557,N_29578);
or UO_2000 (O_2000,N_25092,N_28524);
nor UO_2001 (O_2001,N_28973,N_29020);
or UO_2002 (O_2002,N_26150,N_25390);
nand UO_2003 (O_2003,N_27158,N_28408);
and UO_2004 (O_2004,N_26488,N_28440);
or UO_2005 (O_2005,N_29778,N_28445);
nand UO_2006 (O_2006,N_28726,N_29141);
nor UO_2007 (O_2007,N_26445,N_27995);
nor UO_2008 (O_2008,N_28999,N_26750);
nand UO_2009 (O_2009,N_28005,N_27061);
and UO_2010 (O_2010,N_25534,N_26792);
nor UO_2011 (O_2011,N_25223,N_25409);
xor UO_2012 (O_2012,N_25704,N_28527);
nor UO_2013 (O_2013,N_25044,N_27191);
nand UO_2014 (O_2014,N_28812,N_26401);
xor UO_2015 (O_2015,N_27514,N_29412);
xor UO_2016 (O_2016,N_25649,N_28693);
and UO_2017 (O_2017,N_27509,N_29162);
or UO_2018 (O_2018,N_28759,N_25229);
nand UO_2019 (O_2019,N_28287,N_25750);
and UO_2020 (O_2020,N_28497,N_27941);
nand UO_2021 (O_2021,N_26614,N_27382);
and UO_2022 (O_2022,N_27818,N_25721);
nand UO_2023 (O_2023,N_26558,N_25033);
or UO_2024 (O_2024,N_27955,N_27173);
nand UO_2025 (O_2025,N_29897,N_25299);
or UO_2026 (O_2026,N_27476,N_28932);
nand UO_2027 (O_2027,N_25818,N_27006);
nor UO_2028 (O_2028,N_26194,N_25673);
nand UO_2029 (O_2029,N_29858,N_29805);
and UO_2030 (O_2030,N_26165,N_26023);
nand UO_2031 (O_2031,N_27287,N_27290);
and UO_2032 (O_2032,N_29481,N_27365);
nor UO_2033 (O_2033,N_29785,N_29425);
xnor UO_2034 (O_2034,N_28420,N_29530);
or UO_2035 (O_2035,N_25046,N_28816);
or UO_2036 (O_2036,N_29449,N_27121);
and UO_2037 (O_2037,N_29971,N_29535);
xnor UO_2038 (O_2038,N_29901,N_27988);
nand UO_2039 (O_2039,N_26144,N_25106);
xnor UO_2040 (O_2040,N_29160,N_27671);
nor UO_2041 (O_2041,N_27219,N_26427);
xor UO_2042 (O_2042,N_27949,N_26762);
and UO_2043 (O_2043,N_26845,N_26307);
xnor UO_2044 (O_2044,N_26852,N_28523);
xnor UO_2045 (O_2045,N_29482,N_27032);
nand UO_2046 (O_2046,N_27350,N_25625);
nor UO_2047 (O_2047,N_27468,N_28752);
nand UO_2048 (O_2048,N_25758,N_26860);
and UO_2049 (O_2049,N_26397,N_29734);
xnor UO_2050 (O_2050,N_28493,N_28170);
nor UO_2051 (O_2051,N_26767,N_27247);
nor UO_2052 (O_2052,N_29274,N_26741);
nand UO_2053 (O_2053,N_28730,N_26280);
nand UO_2054 (O_2054,N_25938,N_25368);
nand UO_2055 (O_2055,N_27154,N_25767);
or UO_2056 (O_2056,N_27982,N_28859);
or UO_2057 (O_2057,N_28625,N_27870);
or UO_2058 (O_2058,N_27529,N_25578);
nor UO_2059 (O_2059,N_27394,N_25577);
and UO_2060 (O_2060,N_28873,N_26811);
xor UO_2061 (O_2061,N_29993,N_28676);
nor UO_2062 (O_2062,N_26936,N_29831);
nand UO_2063 (O_2063,N_25149,N_26135);
or UO_2064 (O_2064,N_25032,N_29190);
xor UO_2065 (O_2065,N_25437,N_28063);
nand UO_2066 (O_2066,N_27217,N_28270);
and UO_2067 (O_2067,N_29222,N_28190);
xnor UO_2068 (O_2068,N_25744,N_26755);
or UO_2069 (O_2069,N_28156,N_26287);
and UO_2070 (O_2070,N_26225,N_26289);
or UO_2071 (O_2071,N_25696,N_29545);
xor UO_2072 (O_2072,N_28087,N_29102);
and UO_2073 (O_2073,N_25219,N_25066);
nor UO_2074 (O_2074,N_29130,N_29981);
xnor UO_2075 (O_2075,N_25076,N_28210);
or UO_2076 (O_2076,N_25087,N_28610);
and UO_2077 (O_2077,N_29713,N_27708);
nor UO_2078 (O_2078,N_26473,N_29590);
and UO_2079 (O_2079,N_27404,N_29074);
nor UO_2080 (O_2080,N_26217,N_29093);
nand UO_2081 (O_2081,N_26364,N_29905);
nor UO_2082 (O_2082,N_27122,N_28289);
nand UO_2083 (O_2083,N_25634,N_27831);
nor UO_2084 (O_2084,N_29185,N_25268);
or UO_2085 (O_2085,N_25667,N_26481);
xor UO_2086 (O_2086,N_25422,N_27373);
nor UO_2087 (O_2087,N_25198,N_28568);
nor UO_2088 (O_2088,N_29524,N_26152);
or UO_2089 (O_2089,N_28931,N_26828);
or UO_2090 (O_2090,N_26854,N_29688);
and UO_2091 (O_2091,N_29960,N_28669);
xnor UO_2092 (O_2092,N_26070,N_28252);
xor UO_2093 (O_2093,N_29722,N_28338);
nor UO_2094 (O_2094,N_25354,N_28807);
and UO_2095 (O_2095,N_29572,N_28819);
nand UO_2096 (O_2096,N_29051,N_25669);
nand UO_2097 (O_2097,N_26806,N_25204);
and UO_2098 (O_2098,N_29536,N_28430);
nand UO_2099 (O_2099,N_27550,N_26482);
xnor UO_2100 (O_2100,N_28750,N_28471);
nor UO_2101 (O_2101,N_26940,N_26677);
or UO_2102 (O_2102,N_25849,N_26067);
xor UO_2103 (O_2103,N_26619,N_27752);
or UO_2104 (O_2104,N_28209,N_29437);
xnor UO_2105 (O_2105,N_29300,N_26046);
or UO_2106 (O_2106,N_29516,N_29733);
nor UO_2107 (O_2107,N_25105,N_25222);
or UO_2108 (O_2108,N_26492,N_25408);
or UO_2109 (O_2109,N_29390,N_28808);
and UO_2110 (O_2110,N_29730,N_25672);
nor UO_2111 (O_2111,N_28300,N_28886);
nor UO_2112 (O_2112,N_25452,N_26934);
nand UO_2113 (O_2113,N_29388,N_26204);
or UO_2114 (O_2114,N_29477,N_29122);
xor UO_2115 (O_2115,N_28076,N_25475);
nor UO_2116 (O_2116,N_28578,N_25748);
nand UO_2117 (O_2117,N_27493,N_26051);
nor UO_2118 (O_2118,N_28285,N_27834);
nor UO_2119 (O_2119,N_26704,N_27044);
or UO_2120 (O_2120,N_29894,N_25266);
nor UO_2121 (O_2121,N_27924,N_29492);
nor UO_2122 (O_2122,N_29199,N_28196);
nor UO_2123 (O_2123,N_25499,N_29818);
nor UO_2124 (O_2124,N_28927,N_25010);
nor UO_2125 (O_2125,N_29658,N_28120);
nand UO_2126 (O_2126,N_25453,N_25906);
or UO_2127 (O_2127,N_27580,N_27176);
or UO_2128 (O_2128,N_28806,N_25892);
nor UO_2129 (O_2129,N_29429,N_25477);
xor UO_2130 (O_2130,N_25158,N_27372);
nor UO_2131 (O_2131,N_26623,N_27968);
and UO_2132 (O_2132,N_26954,N_28103);
or UO_2133 (O_2133,N_26282,N_26394);
xnor UO_2134 (O_2134,N_25769,N_25017);
or UO_2135 (O_2135,N_29157,N_27008);
nor UO_2136 (O_2136,N_28918,N_27336);
xnor UO_2137 (O_2137,N_26393,N_28986);
nor UO_2138 (O_2138,N_29146,N_26276);
xor UO_2139 (O_2139,N_25470,N_26719);
nand UO_2140 (O_2140,N_29769,N_26693);
or UO_2141 (O_2141,N_28485,N_28267);
nor UO_2142 (O_2142,N_28559,N_27558);
or UO_2143 (O_2143,N_27377,N_25173);
or UO_2144 (O_2144,N_28540,N_25081);
and UO_2145 (O_2145,N_26554,N_25217);
nor UO_2146 (O_2146,N_27443,N_25814);
and UO_2147 (O_2147,N_29124,N_25979);
xnor UO_2148 (O_2148,N_29165,N_29434);
and UO_2149 (O_2149,N_26285,N_27441);
and UO_2150 (O_2150,N_25251,N_28026);
and UO_2151 (O_2151,N_25982,N_26333);
or UO_2152 (O_2152,N_28185,N_28339);
and UO_2153 (O_2153,N_26331,N_25162);
or UO_2154 (O_2154,N_29774,N_27545);
nand UO_2155 (O_2155,N_29974,N_27811);
and UO_2156 (O_2156,N_27093,N_26788);
nand UO_2157 (O_2157,N_28583,N_29472);
nor UO_2158 (O_2158,N_26759,N_27620);
nand UO_2159 (O_2159,N_27711,N_27230);
and UO_2160 (O_2160,N_28664,N_27832);
and UO_2161 (O_2161,N_25135,N_28104);
xor UO_2162 (O_2162,N_26637,N_27907);
nand UO_2163 (O_2163,N_26202,N_26323);
and UO_2164 (O_2164,N_28724,N_27375);
nor UO_2165 (O_2165,N_27308,N_28582);
nor UO_2166 (O_2166,N_28407,N_28401);
nand UO_2167 (O_2167,N_29480,N_29582);
and UO_2168 (O_2168,N_25333,N_28118);
or UO_2169 (O_2169,N_29789,N_28223);
nor UO_2170 (O_2170,N_26544,N_26699);
nand UO_2171 (O_2171,N_29906,N_29989);
xnor UO_2172 (O_2172,N_27480,N_29909);
or UO_2173 (O_2173,N_28142,N_28290);
or UO_2174 (O_2174,N_27583,N_28101);
nor UO_2175 (O_2175,N_29084,N_29126);
and UO_2176 (O_2176,N_27816,N_27951);
xnor UO_2177 (O_2177,N_25647,N_28670);
and UO_2178 (O_2178,N_29194,N_26703);
or UO_2179 (O_2179,N_25471,N_29287);
nand UO_2180 (O_2180,N_29488,N_26474);
and UO_2181 (O_2181,N_29706,N_27705);
or UO_2182 (O_2182,N_27763,N_29004);
nor UO_2183 (O_2183,N_25871,N_26622);
nand UO_2184 (O_2184,N_27007,N_27829);
nor UO_2185 (O_2185,N_28474,N_28264);
nand UO_2186 (O_2186,N_25737,N_27263);
xnor UO_2187 (O_2187,N_26090,N_26659);
or UO_2188 (O_2188,N_28232,N_29039);
and UO_2189 (O_2189,N_29306,N_28018);
nor UO_2190 (O_2190,N_25510,N_25086);
xnor UO_2191 (O_2191,N_28266,N_29511);
nand UO_2192 (O_2192,N_29655,N_25922);
nand UO_2193 (O_2193,N_27845,N_25766);
nor UO_2194 (O_2194,N_25630,N_26078);
or UO_2195 (O_2195,N_27987,N_27585);
and UO_2196 (O_2196,N_26077,N_29922);
nor UO_2197 (O_2197,N_26245,N_28905);
nor UO_2198 (O_2198,N_26149,N_29527);
xnor UO_2199 (O_2199,N_29291,N_25352);
xor UO_2200 (O_2200,N_29662,N_28864);
nor UO_2201 (O_2201,N_27491,N_26627);
and UO_2202 (O_2202,N_29966,N_29506);
nand UO_2203 (O_2203,N_28961,N_28086);
xor UO_2204 (O_2204,N_26984,N_28499);
nand UO_2205 (O_2205,N_25653,N_28009);
and UO_2206 (O_2206,N_27436,N_28317);
and UO_2207 (O_2207,N_25190,N_25384);
nand UO_2208 (O_2208,N_25596,N_25336);
or UO_2209 (O_2209,N_27120,N_26993);
and UO_2210 (O_2210,N_26921,N_29409);
nor UO_2211 (O_2211,N_29161,N_25786);
xor UO_2212 (O_2212,N_28680,N_27900);
nand UO_2213 (O_2213,N_25170,N_25203);
nand UO_2214 (O_2214,N_26113,N_28581);
and UO_2215 (O_2215,N_27655,N_28778);
or UO_2216 (O_2216,N_29313,N_26059);
xor UO_2217 (O_2217,N_26745,N_26259);
xnor UO_2218 (O_2218,N_25693,N_29207);
xor UO_2219 (O_2219,N_25727,N_28940);
nand UO_2220 (O_2220,N_26296,N_25339);
and UO_2221 (O_2221,N_27383,N_26162);
nand UO_2222 (O_2222,N_27589,N_26843);
nand UO_2223 (O_2223,N_27334,N_29934);
xor UO_2224 (O_2224,N_27932,N_26297);
xor UO_2225 (O_2225,N_28393,N_26284);
nor UO_2226 (O_2226,N_27869,N_26724);
nand UO_2227 (O_2227,N_26858,N_28388);
nor UO_2228 (O_2228,N_25345,N_26459);
and UO_2229 (O_2229,N_25007,N_29459);
and UO_2230 (O_2230,N_26891,N_28734);
or UO_2231 (O_2231,N_26810,N_29486);
xor UO_2232 (O_2232,N_29403,N_29447);
xor UO_2233 (O_2233,N_26353,N_29462);
or UO_2234 (O_2234,N_25822,N_29599);
and UO_2235 (O_2235,N_27464,N_26717);
or UO_2236 (O_2236,N_26610,N_25197);
nor UO_2237 (O_2237,N_27392,N_28243);
xor UO_2238 (O_2238,N_25829,N_29256);
or UO_2239 (O_2239,N_29890,N_25444);
nor UO_2240 (O_2240,N_28108,N_26234);
nand UO_2241 (O_2241,N_25706,N_27640);
nand UO_2242 (O_2242,N_25955,N_25404);
or UO_2243 (O_2243,N_29531,N_28768);
xnor UO_2244 (O_2244,N_28776,N_26339);
nor UO_2245 (O_2245,N_26639,N_26410);
or UO_2246 (O_2246,N_26299,N_29834);
nand UO_2247 (O_2247,N_29229,N_29359);
or UO_2248 (O_2248,N_27819,N_29469);
nor UO_2249 (O_2249,N_27892,N_27390);
or UO_2250 (O_2250,N_29786,N_28045);
or UO_2251 (O_2251,N_29794,N_25783);
nand UO_2252 (O_2252,N_27874,N_26780);
and UO_2253 (O_2253,N_29692,N_27697);
or UO_2254 (O_2254,N_29911,N_26536);
and UO_2255 (O_2255,N_27878,N_27481);
or UO_2256 (O_2256,N_28427,N_28917);
nor UO_2257 (O_2257,N_27398,N_28495);
or UO_2258 (O_2258,N_28293,N_26373);
nand UO_2259 (O_2259,N_25606,N_29128);
or UO_2260 (O_2260,N_29432,N_25618);
xnor UO_2261 (O_2261,N_25244,N_28421);
and UO_2262 (O_2262,N_28347,N_27143);
and UO_2263 (O_2263,N_28660,N_26369);
nand UO_2264 (O_2264,N_27790,N_26732);
nor UO_2265 (O_2265,N_26550,N_25174);
or UO_2266 (O_2266,N_26010,N_28258);
or UO_2267 (O_2267,N_26207,N_29342);
and UO_2268 (O_2268,N_25243,N_28755);
xor UO_2269 (O_2269,N_25837,N_25752);
and UO_2270 (O_2270,N_28119,N_26586);
or UO_2271 (O_2271,N_29446,N_26661);
and UO_2272 (O_2272,N_27582,N_25238);
and UO_2273 (O_2273,N_28467,N_28707);
xor UO_2274 (O_2274,N_28125,N_28647);
and UO_2275 (O_2275,N_28914,N_27127);
nor UO_2276 (O_2276,N_25887,N_29416);
nor UO_2277 (O_2277,N_26072,N_29008);
xnor UO_2278 (O_2278,N_29077,N_26856);
nand UO_2279 (O_2279,N_29065,N_28952);
or UO_2280 (O_2280,N_25136,N_26343);
nor UO_2281 (O_2281,N_28361,N_28396);
or UO_2282 (O_2282,N_26214,N_25397);
nor UO_2283 (O_2283,N_29376,N_29892);
and UO_2284 (O_2284,N_29775,N_28843);
nor UO_2285 (O_2285,N_25382,N_28840);
or UO_2286 (O_2286,N_26398,N_29977);
nor UO_2287 (O_2287,N_28900,N_29251);
or UO_2288 (O_2288,N_29686,N_29045);
and UO_2289 (O_2289,N_25705,N_25154);
or UO_2290 (O_2290,N_28383,N_29942);
nor UO_2291 (O_2291,N_28472,N_28197);
nand UO_2292 (O_2292,N_25020,N_27855);
and UO_2293 (O_2293,N_27979,N_27745);
or UO_2294 (O_2294,N_28995,N_28135);
nor UO_2295 (O_2295,N_25560,N_29970);
nand UO_2296 (O_2296,N_29270,N_25519);
nand UO_2297 (O_2297,N_28655,N_26608);
or UO_2298 (O_2298,N_29120,N_26258);
nand UO_2299 (O_2299,N_29846,N_29822);
nor UO_2300 (O_2300,N_25924,N_28066);
or UO_2301 (O_2301,N_28253,N_27575);
or UO_2302 (O_2302,N_29196,N_26132);
xnor UO_2303 (O_2303,N_29255,N_26313);
nor UO_2304 (O_2304,N_25760,N_29875);
or UO_2305 (O_2305,N_27783,N_27228);
nand UO_2306 (O_2306,N_27317,N_29518);
or UO_2307 (O_2307,N_29833,N_25272);
or UO_2308 (O_2308,N_28143,N_26742);
or UO_2309 (O_2309,N_25099,N_28089);
xnor UO_2310 (O_2310,N_26018,N_27531);
nand UO_2311 (O_2311,N_28649,N_29058);
xnor UO_2312 (O_2312,N_27426,N_26035);
or UO_2313 (O_2313,N_25738,N_27797);
nand UO_2314 (O_2314,N_29484,N_25931);
nor UO_2315 (O_2315,N_28874,N_28348);
nand UO_2316 (O_2316,N_29358,N_28585);
nor UO_2317 (O_2317,N_28613,N_28855);
or UO_2318 (O_2318,N_25323,N_28462);
xnor UO_2319 (O_2319,N_27359,N_29320);
nand UO_2320 (O_2320,N_28398,N_25178);
and UO_2321 (O_2321,N_28950,N_29171);
nor UO_2322 (O_2322,N_28288,N_27018);
nor UO_2323 (O_2323,N_25958,N_25128);
xnor UO_2324 (O_2324,N_27329,N_26908);
or UO_2325 (O_2325,N_26754,N_28136);
nor UO_2326 (O_2326,N_28962,N_26598);
nor UO_2327 (O_2327,N_29649,N_29295);
xnor UO_2328 (O_2328,N_27837,N_26288);
nand UO_2329 (O_2329,N_25726,N_27608);
nand UO_2330 (O_2330,N_26063,N_25831);
nand UO_2331 (O_2331,N_25730,N_27827);
xor UO_2332 (O_2332,N_27324,N_25465);
or UO_2333 (O_2333,N_28040,N_28465);
or UO_2334 (O_2334,N_26452,N_26166);
and UO_2335 (O_2335,N_25785,N_26083);
nand UO_2336 (O_2336,N_27930,N_29092);
and UO_2337 (O_2337,N_25884,N_27161);
nor UO_2338 (O_2338,N_28704,N_28978);
xor UO_2339 (O_2339,N_27181,N_29195);
and UO_2340 (O_2340,N_26711,N_27412);
and UO_2341 (O_2341,N_28222,N_28230);
and UO_2342 (O_2342,N_27681,N_27047);
nor UO_2343 (O_2343,N_28091,N_29054);
nor UO_2344 (O_2344,N_29632,N_26877);
nor UO_2345 (O_2345,N_28483,N_25101);
or UO_2346 (O_2346,N_25252,N_26959);
and UO_2347 (O_2347,N_25363,N_27282);
and UO_2348 (O_2348,N_28480,N_27201);
nor UO_2349 (O_2349,N_27224,N_25167);
or UO_2350 (O_2350,N_27449,N_29718);
xnor UO_2351 (O_2351,N_29950,N_29752);
or UO_2352 (O_2352,N_26448,N_26705);
and UO_2353 (O_2353,N_26957,N_28945);
xor UO_2354 (O_2354,N_29703,N_27880);
nand UO_2355 (O_2355,N_27505,N_27923);
nand UO_2356 (O_2356,N_28871,N_26918);
and UO_2357 (O_2357,N_29872,N_29399);
xor UO_2358 (O_2358,N_26582,N_26294);
and UO_2359 (O_2359,N_27142,N_29301);
or UO_2360 (O_2360,N_27243,N_27106);
nor UO_2361 (O_2361,N_25827,N_25432);
and UO_2362 (O_2362,N_26874,N_25971);
xnor UO_2363 (O_2363,N_25356,N_25872);
or UO_2364 (O_2364,N_29969,N_28735);
and UO_2365 (O_2365,N_29546,N_27615);
xor UO_2366 (O_2366,N_29689,N_27572);
nand UO_2367 (O_2367,N_27432,N_28067);
and UO_2368 (O_2368,N_28803,N_27814);
and UO_2369 (O_2369,N_28449,N_26322);
nand UO_2370 (O_2370,N_26048,N_25638);
nand UO_2371 (O_2371,N_29204,N_26425);
nand UO_2372 (O_2372,N_25607,N_25080);
and UO_2373 (O_2373,N_26817,N_28509);
or UO_2374 (O_2374,N_26895,N_27038);
or UO_2375 (O_2375,N_28511,N_29508);
and UO_2376 (O_2376,N_26463,N_29976);
and UO_2377 (O_2377,N_25960,N_27854);
nand UO_2378 (O_2378,N_25181,N_29928);
nor UO_2379 (O_2379,N_25218,N_27914);
xor UO_2380 (O_2380,N_29884,N_27895);
nor UO_2381 (O_2381,N_26409,N_28438);
and UO_2382 (O_2382,N_28639,N_26640);
nor UO_2383 (O_2383,N_26243,N_29883);
nor UO_2384 (O_2384,N_27119,N_29326);
nand UO_2385 (O_2385,N_27174,N_28822);
and UO_2386 (O_2386,N_28979,N_27778);
nand UO_2387 (O_2387,N_26548,N_26606);
nor UO_2388 (O_2388,N_26771,N_27776);
nand UO_2389 (O_2389,N_25745,N_25215);
or UO_2390 (O_2390,N_27109,N_29512);
nand UO_2391 (O_2391,N_29354,N_25359);
xnor UO_2392 (O_2392,N_27958,N_26042);
nor UO_2393 (O_2393,N_28706,N_27330);
and UO_2394 (O_2394,N_25520,N_27728);
or UO_2395 (O_2395,N_29023,N_25843);
nor UO_2396 (O_2396,N_25571,N_25521);
or UO_2397 (O_2397,N_25202,N_28468);
and UO_2398 (O_2398,N_27696,N_28567);
xor UO_2399 (O_2399,N_27396,N_29938);
nand UO_2400 (O_2400,N_25917,N_29559);
nor UO_2401 (O_2401,N_28186,N_25860);
or UO_2402 (O_2402,N_25847,N_25655);
xor UO_2403 (O_2403,N_29843,N_28947);
nand UO_2404 (O_2404,N_27901,N_29382);
and UO_2405 (O_2405,N_27304,N_26822);
or UO_2406 (O_2406,N_26632,N_26275);
or UO_2407 (O_2407,N_25332,N_28852);
nor UO_2408 (O_2408,N_25456,N_25028);
xor UO_2409 (O_2409,N_29575,N_25690);
or UO_2410 (O_2410,N_26781,N_29751);
nand UO_2411 (O_2411,N_25344,N_25039);
nand UO_2412 (O_2412,N_27866,N_28292);
and UO_2413 (O_2413,N_28641,N_26557);
or UO_2414 (O_2414,N_27602,N_28450);
nor UO_2415 (O_2415,N_27475,N_27975);
and UO_2416 (O_2416,N_28795,N_25279);
nand UO_2417 (O_2417,N_25865,N_27488);
or UO_2418 (O_2418,N_29027,N_29605);
xor UO_2419 (O_2419,N_27356,N_29663);
nand UO_2420 (O_2420,N_28014,N_26625);
and UO_2421 (O_2421,N_29731,N_29365);
nand UO_2422 (O_2422,N_29889,N_27384);
or UO_2423 (O_2423,N_26989,N_29961);
or UO_2424 (O_2424,N_28633,N_27709);
or UO_2425 (O_2425,N_25446,N_25415);
or UO_2426 (O_2426,N_27030,N_27548);
nand UO_2427 (O_2427,N_26370,N_25555);
nor UO_2428 (O_2428,N_28802,N_29168);
or UO_2429 (O_2429,N_25736,N_28964);
or UO_2430 (O_2430,N_27374,N_29109);
nor UO_2431 (O_2431,N_25623,N_29930);
xor UO_2432 (O_2432,N_29626,N_28016);
xor UO_2433 (O_2433,N_29174,N_27807);
xor UO_2434 (O_2434,N_26805,N_29344);
nand UO_2435 (O_2435,N_28065,N_26003);
and UO_2436 (O_2436,N_26108,N_27253);
nor UO_2437 (O_2437,N_27905,N_25612);
nor UO_2438 (O_2438,N_26863,N_25230);
xnor UO_2439 (O_2439,N_25644,N_29914);
xnor UO_2440 (O_2440,N_29862,N_29891);
nand UO_2441 (O_2441,N_29826,N_29332);
and UO_2442 (O_2442,N_27518,N_27993);
xnor UO_2443 (O_2443,N_27844,N_28455);
nor UO_2444 (O_2444,N_27279,N_25533);
nand UO_2445 (O_2445,N_29815,N_26534);
or UO_2446 (O_2446,N_26499,N_28829);
nor UO_2447 (O_2447,N_28507,N_28579);
and UO_2448 (O_2448,N_26986,N_25121);
and UO_2449 (O_2449,N_26154,N_28996);
nand UO_2450 (O_2450,N_26414,N_26066);
or UO_2451 (O_2451,N_29749,N_27274);
nor UO_2452 (O_2452,N_28818,N_28508);
nor UO_2453 (O_2453,N_25980,N_28896);
nand UO_2454 (O_2454,N_27010,N_29315);
or UO_2455 (O_2455,N_26960,N_25531);
nand UO_2456 (O_2456,N_27089,N_27470);
xnor UO_2457 (O_2457,N_25912,N_27749);
and UO_2458 (O_2458,N_29963,N_26449);
nand UO_2459 (O_2459,N_28909,N_26675);
xnor UO_2460 (O_2460,N_28098,N_26314);
nor UO_2461 (O_2461,N_29868,N_25226);
xnor UO_2462 (O_2462,N_28192,N_28937);
or UO_2463 (O_2463,N_29646,N_29233);
nor UO_2464 (O_2464,N_27199,N_29025);
nor UO_2465 (O_2465,N_28980,N_28151);
nand UO_2466 (O_2466,N_29221,N_27484);
xnor UO_2467 (O_2467,N_26060,N_27313);
or UO_2468 (O_2468,N_25558,N_28363);
and UO_2469 (O_2469,N_29680,N_29018);
or UO_2470 (O_2470,N_25541,N_25450);
and UO_2471 (O_2471,N_27934,N_25469);
xor UO_2472 (O_2472,N_27203,N_29000);
or UO_2473 (O_2473,N_28249,N_28111);
and UO_2474 (O_2474,N_28604,N_28774);
or UO_2475 (O_2475,N_27168,N_29719);
xor UO_2476 (O_2476,N_29593,N_27239);
nand UO_2477 (O_2477,N_29859,N_27717);
xnor UO_2478 (O_2478,N_28139,N_26978);
and UO_2479 (O_2479,N_29364,N_29200);
nor UO_2480 (O_2480,N_28017,N_25597);
nand UO_2481 (O_2481,N_26531,N_29260);
and UO_2482 (O_2482,N_29234,N_29700);
and UO_2483 (O_2483,N_27825,N_29475);
xor UO_2484 (O_2484,N_26773,N_27775);
nand UO_2485 (O_2485,N_26971,N_29153);
nand UO_2486 (O_2486,N_28989,N_25677);
nand UO_2487 (O_2487,N_29280,N_28858);
xnor UO_2488 (O_2488,N_28743,N_28278);
nor UO_2489 (O_2489,N_27759,N_26147);
and UO_2490 (O_2490,N_28702,N_27748);
and UO_2491 (O_2491,N_29571,N_29408);
nor UO_2492 (O_2492,N_25288,N_29790);
or UO_2493 (O_2493,N_27419,N_26907);
nand UO_2494 (O_2494,N_27546,N_25286);
and UO_2495 (O_2495,N_25825,N_27936);
or UO_2496 (O_2496,N_28327,N_28160);
nor UO_2497 (O_2497,N_27858,N_29192);
nand UO_2498 (O_2498,N_26128,N_27285);
nand UO_2499 (O_2499,N_29138,N_27826);
nor UO_2500 (O_2500,N_25543,N_29527);
and UO_2501 (O_2501,N_27060,N_26044);
nor UO_2502 (O_2502,N_27932,N_25858);
and UO_2503 (O_2503,N_29203,N_29326);
and UO_2504 (O_2504,N_29268,N_26730);
nand UO_2505 (O_2505,N_28385,N_25862);
or UO_2506 (O_2506,N_29517,N_28524);
or UO_2507 (O_2507,N_28068,N_25696);
xor UO_2508 (O_2508,N_29503,N_29009);
nor UO_2509 (O_2509,N_29456,N_25106);
xnor UO_2510 (O_2510,N_27040,N_29772);
nand UO_2511 (O_2511,N_27772,N_27207);
or UO_2512 (O_2512,N_27753,N_28637);
nand UO_2513 (O_2513,N_27985,N_28305);
and UO_2514 (O_2514,N_25405,N_28465);
nor UO_2515 (O_2515,N_26216,N_28921);
xor UO_2516 (O_2516,N_29229,N_27064);
nor UO_2517 (O_2517,N_27323,N_27748);
or UO_2518 (O_2518,N_29131,N_27552);
xor UO_2519 (O_2519,N_29831,N_25395);
nor UO_2520 (O_2520,N_27949,N_28099);
xnor UO_2521 (O_2521,N_27592,N_26231);
or UO_2522 (O_2522,N_26929,N_27610);
xor UO_2523 (O_2523,N_26208,N_25544);
or UO_2524 (O_2524,N_29474,N_27216);
or UO_2525 (O_2525,N_28390,N_25149);
xor UO_2526 (O_2526,N_28245,N_26893);
or UO_2527 (O_2527,N_29045,N_28220);
or UO_2528 (O_2528,N_29471,N_25681);
xor UO_2529 (O_2529,N_28303,N_28851);
xor UO_2530 (O_2530,N_26321,N_29894);
nor UO_2531 (O_2531,N_25316,N_29792);
nand UO_2532 (O_2532,N_27592,N_27163);
nand UO_2533 (O_2533,N_26699,N_25569);
or UO_2534 (O_2534,N_26425,N_29581);
nand UO_2535 (O_2535,N_27119,N_29024);
nor UO_2536 (O_2536,N_26064,N_25282);
nor UO_2537 (O_2537,N_26164,N_26877);
nor UO_2538 (O_2538,N_28882,N_28299);
or UO_2539 (O_2539,N_27433,N_26760);
or UO_2540 (O_2540,N_28892,N_26031);
and UO_2541 (O_2541,N_29511,N_25425);
or UO_2542 (O_2542,N_27545,N_26996);
and UO_2543 (O_2543,N_25170,N_27469);
nor UO_2544 (O_2544,N_27309,N_28019);
and UO_2545 (O_2545,N_27071,N_26493);
nand UO_2546 (O_2546,N_27309,N_29311);
nand UO_2547 (O_2547,N_29420,N_25122);
nand UO_2548 (O_2548,N_25330,N_26936);
or UO_2549 (O_2549,N_27631,N_27707);
xor UO_2550 (O_2550,N_26296,N_26408);
or UO_2551 (O_2551,N_29555,N_28856);
xnor UO_2552 (O_2552,N_29394,N_27372);
and UO_2553 (O_2553,N_29044,N_26325);
or UO_2554 (O_2554,N_27851,N_27059);
and UO_2555 (O_2555,N_28476,N_29653);
nor UO_2556 (O_2556,N_25843,N_26123);
or UO_2557 (O_2557,N_27937,N_29562);
and UO_2558 (O_2558,N_28085,N_28185);
nor UO_2559 (O_2559,N_27102,N_27948);
or UO_2560 (O_2560,N_25019,N_29794);
nand UO_2561 (O_2561,N_25865,N_25565);
nand UO_2562 (O_2562,N_27497,N_28869);
xnor UO_2563 (O_2563,N_29575,N_29673);
or UO_2564 (O_2564,N_29507,N_25746);
or UO_2565 (O_2565,N_29300,N_29161);
or UO_2566 (O_2566,N_29437,N_27927);
xor UO_2567 (O_2567,N_29305,N_25969);
xor UO_2568 (O_2568,N_27471,N_25085);
nor UO_2569 (O_2569,N_29921,N_29289);
nor UO_2570 (O_2570,N_26498,N_26933);
and UO_2571 (O_2571,N_27615,N_28235);
or UO_2572 (O_2572,N_26003,N_26259);
nand UO_2573 (O_2573,N_27708,N_25436);
and UO_2574 (O_2574,N_29589,N_29919);
nand UO_2575 (O_2575,N_29327,N_28993);
nand UO_2576 (O_2576,N_28755,N_25869);
nor UO_2577 (O_2577,N_25532,N_26863);
nand UO_2578 (O_2578,N_26935,N_28983);
nand UO_2579 (O_2579,N_25346,N_26465);
nor UO_2580 (O_2580,N_29315,N_25482);
xor UO_2581 (O_2581,N_27858,N_27086);
nor UO_2582 (O_2582,N_28311,N_27266);
xor UO_2583 (O_2583,N_28766,N_27908);
or UO_2584 (O_2584,N_25844,N_29429);
nand UO_2585 (O_2585,N_29985,N_28671);
nor UO_2586 (O_2586,N_26098,N_29499);
xnor UO_2587 (O_2587,N_25241,N_26087);
xor UO_2588 (O_2588,N_26611,N_25264);
nor UO_2589 (O_2589,N_25432,N_28684);
xnor UO_2590 (O_2590,N_29538,N_27154);
nor UO_2591 (O_2591,N_27779,N_29406);
xnor UO_2592 (O_2592,N_27339,N_29372);
xor UO_2593 (O_2593,N_29629,N_28496);
nand UO_2594 (O_2594,N_27692,N_27326);
nor UO_2595 (O_2595,N_29336,N_25893);
nor UO_2596 (O_2596,N_28922,N_27962);
xor UO_2597 (O_2597,N_27722,N_25042);
and UO_2598 (O_2598,N_28892,N_26230);
or UO_2599 (O_2599,N_26729,N_26400);
nor UO_2600 (O_2600,N_28817,N_25173);
and UO_2601 (O_2601,N_29141,N_27623);
or UO_2602 (O_2602,N_25798,N_29383);
xnor UO_2603 (O_2603,N_26048,N_25223);
xor UO_2604 (O_2604,N_28856,N_25972);
nand UO_2605 (O_2605,N_25709,N_28953);
nor UO_2606 (O_2606,N_27440,N_28222);
or UO_2607 (O_2607,N_29310,N_28321);
xor UO_2608 (O_2608,N_26078,N_29761);
and UO_2609 (O_2609,N_27275,N_27413);
xor UO_2610 (O_2610,N_26374,N_27043);
xnor UO_2611 (O_2611,N_25789,N_26220);
or UO_2612 (O_2612,N_29180,N_26240);
or UO_2613 (O_2613,N_25428,N_28524);
and UO_2614 (O_2614,N_27713,N_29611);
nor UO_2615 (O_2615,N_25424,N_29760);
and UO_2616 (O_2616,N_29589,N_27593);
nand UO_2617 (O_2617,N_26444,N_26389);
nor UO_2618 (O_2618,N_29246,N_26003);
xor UO_2619 (O_2619,N_27359,N_29270);
and UO_2620 (O_2620,N_27324,N_27541);
xnor UO_2621 (O_2621,N_27252,N_25840);
nand UO_2622 (O_2622,N_25672,N_26210);
or UO_2623 (O_2623,N_27432,N_27466);
nor UO_2624 (O_2624,N_26878,N_26042);
and UO_2625 (O_2625,N_29421,N_29823);
nor UO_2626 (O_2626,N_27229,N_28326);
nor UO_2627 (O_2627,N_27897,N_25006);
xor UO_2628 (O_2628,N_29156,N_25178);
and UO_2629 (O_2629,N_27737,N_29212);
nand UO_2630 (O_2630,N_26592,N_26238);
xor UO_2631 (O_2631,N_25703,N_28562);
nor UO_2632 (O_2632,N_29031,N_28670);
or UO_2633 (O_2633,N_25300,N_28128);
or UO_2634 (O_2634,N_26411,N_29438);
or UO_2635 (O_2635,N_26957,N_28922);
xnor UO_2636 (O_2636,N_29633,N_29876);
xnor UO_2637 (O_2637,N_26040,N_26676);
and UO_2638 (O_2638,N_27798,N_25983);
or UO_2639 (O_2639,N_28914,N_25579);
or UO_2640 (O_2640,N_27659,N_25889);
and UO_2641 (O_2641,N_28853,N_26143);
nand UO_2642 (O_2642,N_25545,N_26443);
nand UO_2643 (O_2643,N_26053,N_27371);
nor UO_2644 (O_2644,N_26758,N_28636);
and UO_2645 (O_2645,N_26085,N_26099);
or UO_2646 (O_2646,N_25038,N_26559);
and UO_2647 (O_2647,N_25902,N_26471);
nor UO_2648 (O_2648,N_29581,N_29971);
and UO_2649 (O_2649,N_25371,N_29774);
nor UO_2650 (O_2650,N_26425,N_26128);
and UO_2651 (O_2651,N_25678,N_26644);
nor UO_2652 (O_2652,N_25600,N_29532);
or UO_2653 (O_2653,N_27900,N_29202);
nor UO_2654 (O_2654,N_28420,N_28705);
xor UO_2655 (O_2655,N_26668,N_27672);
nand UO_2656 (O_2656,N_29186,N_29174);
nor UO_2657 (O_2657,N_26963,N_29118);
and UO_2658 (O_2658,N_26988,N_26586);
xor UO_2659 (O_2659,N_25471,N_29378);
nor UO_2660 (O_2660,N_29702,N_28770);
nand UO_2661 (O_2661,N_29547,N_29169);
or UO_2662 (O_2662,N_27415,N_27203);
or UO_2663 (O_2663,N_25175,N_26049);
nand UO_2664 (O_2664,N_25215,N_27140);
and UO_2665 (O_2665,N_28500,N_27748);
nor UO_2666 (O_2666,N_29174,N_27799);
or UO_2667 (O_2667,N_25674,N_29181);
nand UO_2668 (O_2668,N_26260,N_26055);
nor UO_2669 (O_2669,N_26253,N_25657);
nor UO_2670 (O_2670,N_27697,N_27457);
xor UO_2671 (O_2671,N_27025,N_29873);
xnor UO_2672 (O_2672,N_29573,N_29532);
nand UO_2673 (O_2673,N_26480,N_25194);
nand UO_2674 (O_2674,N_25161,N_29130);
and UO_2675 (O_2675,N_29365,N_29001);
or UO_2676 (O_2676,N_25733,N_29650);
and UO_2677 (O_2677,N_29931,N_25372);
nor UO_2678 (O_2678,N_28815,N_28434);
nor UO_2679 (O_2679,N_25078,N_29369);
nand UO_2680 (O_2680,N_27176,N_27598);
nor UO_2681 (O_2681,N_26481,N_26612);
nor UO_2682 (O_2682,N_27671,N_29332);
xnor UO_2683 (O_2683,N_26117,N_26835);
nor UO_2684 (O_2684,N_27507,N_27070);
nor UO_2685 (O_2685,N_25723,N_26846);
nand UO_2686 (O_2686,N_28794,N_25544);
and UO_2687 (O_2687,N_26574,N_26153);
xnor UO_2688 (O_2688,N_28483,N_29892);
xnor UO_2689 (O_2689,N_29466,N_28889);
nor UO_2690 (O_2690,N_26678,N_29992);
or UO_2691 (O_2691,N_29908,N_28545);
nand UO_2692 (O_2692,N_26038,N_28706);
nor UO_2693 (O_2693,N_28997,N_27061);
xor UO_2694 (O_2694,N_25076,N_26408);
and UO_2695 (O_2695,N_29927,N_26050);
and UO_2696 (O_2696,N_28801,N_28045);
and UO_2697 (O_2697,N_26643,N_27846);
nand UO_2698 (O_2698,N_29030,N_29647);
nand UO_2699 (O_2699,N_25930,N_26920);
xor UO_2700 (O_2700,N_27881,N_25800);
nor UO_2701 (O_2701,N_28626,N_25661);
and UO_2702 (O_2702,N_25467,N_27197);
or UO_2703 (O_2703,N_29392,N_27639);
xnor UO_2704 (O_2704,N_29977,N_28454);
nand UO_2705 (O_2705,N_25854,N_25920);
and UO_2706 (O_2706,N_25608,N_28175);
and UO_2707 (O_2707,N_26005,N_28903);
xnor UO_2708 (O_2708,N_28307,N_29015);
and UO_2709 (O_2709,N_27842,N_27311);
or UO_2710 (O_2710,N_29979,N_28350);
nand UO_2711 (O_2711,N_28255,N_28611);
nand UO_2712 (O_2712,N_25457,N_25751);
xnor UO_2713 (O_2713,N_25609,N_28999);
and UO_2714 (O_2714,N_27662,N_26188);
xor UO_2715 (O_2715,N_25914,N_27956);
nor UO_2716 (O_2716,N_28846,N_26011);
or UO_2717 (O_2717,N_29359,N_26448);
nand UO_2718 (O_2718,N_27330,N_26041);
and UO_2719 (O_2719,N_29720,N_27811);
and UO_2720 (O_2720,N_28057,N_28357);
nor UO_2721 (O_2721,N_25405,N_26560);
and UO_2722 (O_2722,N_26004,N_29173);
nand UO_2723 (O_2723,N_29802,N_28378);
nor UO_2724 (O_2724,N_28504,N_27833);
nand UO_2725 (O_2725,N_27630,N_28684);
xnor UO_2726 (O_2726,N_29788,N_26329);
xor UO_2727 (O_2727,N_27868,N_25958);
or UO_2728 (O_2728,N_27432,N_28567);
or UO_2729 (O_2729,N_28865,N_29023);
or UO_2730 (O_2730,N_28212,N_29552);
or UO_2731 (O_2731,N_27377,N_25983);
nor UO_2732 (O_2732,N_25107,N_26991);
nor UO_2733 (O_2733,N_27077,N_28185);
nor UO_2734 (O_2734,N_28746,N_29771);
xor UO_2735 (O_2735,N_29015,N_27537);
nor UO_2736 (O_2736,N_26572,N_29979);
and UO_2737 (O_2737,N_28087,N_25152);
or UO_2738 (O_2738,N_26413,N_25883);
and UO_2739 (O_2739,N_26935,N_27359);
nor UO_2740 (O_2740,N_28014,N_27487);
and UO_2741 (O_2741,N_27808,N_25881);
nor UO_2742 (O_2742,N_25870,N_25597);
nand UO_2743 (O_2743,N_28294,N_25514);
or UO_2744 (O_2744,N_29589,N_25814);
xnor UO_2745 (O_2745,N_29195,N_29425);
and UO_2746 (O_2746,N_29948,N_27136);
nor UO_2747 (O_2747,N_27695,N_26112);
nor UO_2748 (O_2748,N_25716,N_26232);
or UO_2749 (O_2749,N_26584,N_28987);
nand UO_2750 (O_2750,N_29801,N_25324);
and UO_2751 (O_2751,N_25440,N_26682);
or UO_2752 (O_2752,N_25960,N_25071);
nor UO_2753 (O_2753,N_28587,N_29931);
or UO_2754 (O_2754,N_28218,N_25307);
nand UO_2755 (O_2755,N_29944,N_29921);
or UO_2756 (O_2756,N_25357,N_25555);
or UO_2757 (O_2757,N_26361,N_25377);
nand UO_2758 (O_2758,N_26097,N_25419);
or UO_2759 (O_2759,N_26082,N_27559);
nand UO_2760 (O_2760,N_27149,N_26455);
xnor UO_2761 (O_2761,N_27438,N_29316);
xnor UO_2762 (O_2762,N_26283,N_25668);
and UO_2763 (O_2763,N_29360,N_27347);
xor UO_2764 (O_2764,N_28633,N_25576);
and UO_2765 (O_2765,N_29086,N_27778);
or UO_2766 (O_2766,N_25546,N_29123);
and UO_2767 (O_2767,N_28345,N_25774);
or UO_2768 (O_2768,N_28843,N_29858);
or UO_2769 (O_2769,N_29640,N_29616);
and UO_2770 (O_2770,N_29807,N_28720);
xor UO_2771 (O_2771,N_26303,N_28111);
xor UO_2772 (O_2772,N_25218,N_28735);
nand UO_2773 (O_2773,N_27313,N_27714);
xnor UO_2774 (O_2774,N_25689,N_28648);
nor UO_2775 (O_2775,N_27738,N_28482);
xnor UO_2776 (O_2776,N_27726,N_28367);
and UO_2777 (O_2777,N_28420,N_26225);
xnor UO_2778 (O_2778,N_28527,N_26544);
or UO_2779 (O_2779,N_26326,N_25191);
nor UO_2780 (O_2780,N_27682,N_28814);
and UO_2781 (O_2781,N_29690,N_29538);
or UO_2782 (O_2782,N_29798,N_26422);
nor UO_2783 (O_2783,N_27178,N_26702);
or UO_2784 (O_2784,N_28290,N_27583);
nand UO_2785 (O_2785,N_29898,N_25178);
or UO_2786 (O_2786,N_29617,N_28687);
or UO_2787 (O_2787,N_26013,N_25003);
and UO_2788 (O_2788,N_27532,N_25448);
and UO_2789 (O_2789,N_28878,N_27429);
or UO_2790 (O_2790,N_27288,N_28578);
and UO_2791 (O_2791,N_26347,N_29137);
nand UO_2792 (O_2792,N_29551,N_27997);
nor UO_2793 (O_2793,N_27322,N_27798);
xnor UO_2794 (O_2794,N_28721,N_29777);
and UO_2795 (O_2795,N_29904,N_27957);
nand UO_2796 (O_2796,N_29343,N_25994);
and UO_2797 (O_2797,N_26442,N_28131);
nand UO_2798 (O_2798,N_26905,N_29136);
xor UO_2799 (O_2799,N_27305,N_29917);
and UO_2800 (O_2800,N_25591,N_29829);
or UO_2801 (O_2801,N_27540,N_25261);
xnor UO_2802 (O_2802,N_27524,N_29366);
nor UO_2803 (O_2803,N_27553,N_25983);
xnor UO_2804 (O_2804,N_29445,N_28757);
and UO_2805 (O_2805,N_26156,N_27866);
nor UO_2806 (O_2806,N_27105,N_28283);
nor UO_2807 (O_2807,N_27200,N_27315);
nand UO_2808 (O_2808,N_27305,N_26527);
xor UO_2809 (O_2809,N_27058,N_28474);
and UO_2810 (O_2810,N_29883,N_29995);
or UO_2811 (O_2811,N_25130,N_29552);
nand UO_2812 (O_2812,N_25795,N_25078);
and UO_2813 (O_2813,N_26973,N_25447);
or UO_2814 (O_2814,N_28871,N_29515);
and UO_2815 (O_2815,N_28488,N_26692);
nor UO_2816 (O_2816,N_29589,N_29196);
nor UO_2817 (O_2817,N_27703,N_25210);
or UO_2818 (O_2818,N_29311,N_28645);
nor UO_2819 (O_2819,N_28252,N_28429);
nor UO_2820 (O_2820,N_28063,N_27679);
and UO_2821 (O_2821,N_26524,N_28844);
nand UO_2822 (O_2822,N_26576,N_27984);
nand UO_2823 (O_2823,N_27529,N_28159);
nor UO_2824 (O_2824,N_29347,N_28322);
nand UO_2825 (O_2825,N_27222,N_27739);
or UO_2826 (O_2826,N_29393,N_26096);
xor UO_2827 (O_2827,N_26482,N_28125);
or UO_2828 (O_2828,N_25119,N_27373);
nor UO_2829 (O_2829,N_28335,N_26470);
nor UO_2830 (O_2830,N_29216,N_29242);
nor UO_2831 (O_2831,N_27304,N_26619);
and UO_2832 (O_2832,N_25243,N_27673);
nor UO_2833 (O_2833,N_26783,N_28683);
nor UO_2834 (O_2834,N_29556,N_26858);
nor UO_2835 (O_2835,N_25101,N_26866);
or UO_2836 (O_2836,N_25746,N_29147);
nor UO_2837 (O_2837,N_25522,N_25857);
and UO_2838 (O_2838,N_29717,N_28634);
xor UO_2839 (O_2839,N_25071,N_29430);
nor UO_2840 (O_2840,N_28742,N_27915);
nor UO_2841 (O_2841,N_26859,N_28573);
xnor UO_2842 (O_2842,N_28606,N_27735);
and UO_2843 (O_2843,N_29414,N_29235);
xor UO_2844 (O_2844,N_29479,N_29239);
nor UO_2845 (O_2845,N_26630,N_27259);
and UO_2846 (O_2846,N_28907,N_28553);
nand UO_2847 (O_2847,N_27041,N_29935);
and UO_2848 (O_2848,N_29899,N_27790);
or UO_2849 (O_2849,N_25537,N_26667);
or UO_2850 (O_2850,N_25305,N_25955);
or UO_2851 (O_2851,N_27089,N_29732);
xor UO_2852 (O_2852,N_27948,N_27738);
xnor UO_2853 (O_2853,N_27364,N_26026);
or UO_2854 (O_2854,N_26169,N_27407);
or UO_2855 (O_2855,N_28359,N_29612);
nor UO_2856 (O_2856,N_28322,N_25831);
nor UO_2857 (O_2857,N_29252,N_27771);
nor UO_2858 (O_2858,N_25790,N_27892);
and UO_2859 (O_2859,N_25057,N_27757);
nand UO_2860 (O_2860,N_26084,N_26397);
nor UO_2861 (O_2861,N_28292,N_26114);
xor UO_2862 (O_2862,N_29266,N_27924);
and UO_2863 (O_2863,N_27717,N_29786);
and UO_2864 (O_2864,N_28500,N_27363);
nand UO_2865 (O_2865,N_26028,N_26833);
nor UO_2866 (O_2866,N_25738,N_29400);
and UO_2867 (O_2867,N_28954,N_29479);
nor UO_2868 (O_2868,N_28600,N_27395);
or UO_2869 (O_2869,N_25109,N_26947);
nand UO_2870 (O_2870,N_28063,N_26082);
and UO_2871 (O_2871,N_28691,N_27284);
nor UO_2872 (O_2872,N_28196,N_28758);
nor UO_2873 (O_2873,N_27360,N_25772);
or UO_2874 (O_2874,N_25934,N_29870);
and UO_2875 (O_2875,N_29053,N_28283);
nor UO_2876 (O_2876,N_25871,N_29198);
or UO_2877 (O_2877,N_27067,N_26067);
or UO_2878 (O_2878,N_29803,N_26029);
or UO_2879 (O_2879,N_28744,N_28098);
nor UO_2880 (O_2880,N_28289,N_27887);
nor UO_2881 (O_2881,N_26462,N_25170);
or UO_2882 (O_2882,N_26606,N_25108);
and UO_2883 (O_2883,N_26550,N_25720);
nor UO_2884 (O_2884,N_29617,N_27514);
nand UO_2885 (O_2885,N_26787,N_29145);
and UO_2886 (O_2886,N_28335,N_29544);
xor UO_2887 (O_2887,N_25817,N_26459);
nand UO_2888 (O_2888,N_27793,N_29463);
nand UO_2889 (O_2889,N_28678,N_25347);
xnor UO_2890 (O_2890,N_28106,N_26678);
xnor UO_2891 (O_2891,N_27000,N_27372);
nand UO_2892 (O_2892,N_29365,N_25015);
xnor UO_2893 (O_2893,N_25061,N_26799);
nor UO_2894 (O_2894,N_27535,N_25381);
nor UO_2895 (O_2895,N_27786,N_29069);
xnor UO_2896 (O_2896,N_29683,N_28983);
and UO_2897 (O_2897,N_25798,N_29990);
nand UO_2898 (O_2898,N_29427,N_25256);
or UO_2899 (O_2899,N_26714,N_27325);
xnor UO_2900 (O_2900,N_28563,N_25206);
and UO_2901 (O_2901,N_29511,N_26128);
or UO_2902 (O_2902,N_29113,N_26406);
nor UO_2903 (O_2903,N_26975,N_28344);
and UO_2904 (O_2904,N_25378,N_26709);
or UO_2905 (O_2905,N_27620,N_26470);
xnor UO_2906 (O_2906,N_26684,N_28899);
and UO_2907 (O_2907,N_28897,N_25198);
and UO_2908 (O_2908,N_25618,N_25882);
and UO_2909 (O_2909,N_29522,N_26414);
nand UO_2910 (O_2910,N_25658,N_26842);
nor UO_2911 (O_2911,N_25835,N_26974);
xor UO_2912 (O_2912,N_28179,N_27828);
nand UO_2913 (O_2913,N_27759,N_28386);
or UO_2914 (O_2914,N_25701,N_29404);
xor UO_2915 (O_2915,N_27459,N_28558);
nand UO_2916 (O_2916,N_28608,N_28648);
xnor UO_2917 (O_2917,N_27865,N_25389);
nand UO_2918 (O_2918,N_28196,N_27175);
xor UO_2919 (O_2919,N_29011,N_27003);
and UO_2920 (O_2920,N_29515,N_28096);
nand UO_2921 (O_2921,N_27703,N_27782);
xnor UO_2922 (O_2922,N_28933,N_27969);
nand UO_2923 (O_2923,N_26024,N_25729);
nand UO_2924 (O_2924,N_29601,N_28340);
or UO_2925 (O_2925,N_27327,N_29511);
and UO_2926 (O_2926,N_28530,N_27654);
xnor UO_2927 (O_2927,N_27495,N_27050);
nor UO_2928 (O_2928,N_27522,N_27693);
or UO_2929 (O_2929,N_29584,N_26565);
nor UO_2930 (O_2930,N_28730,N_27775);
nor UO_2931 (O_2931,N_27587,N_26966);
nor UO_2932 (O_2932,N_26672,N_29706);
xnor UO_2933 (O_2933,N_25595,N_28121);
and UO_2934 (O_2934,N_26235,N_25573);
or UO_2935 (O_2935,N_28968,N_25859);
and UO_2936 (O_2936,N_29346,N_27351);
nand UO_2937 (O_2937,N_29666,N_25729);
nor UO_2938 (O_2938,N_29636,N_28954);
nor UO_2939 (O_2939,N_29596,N_28507);
and UO_2940 (O_2940,N_26378,N_25343);
xor UO_2941 (O_2941,N_26872,N_29813);
nand UO_2942 (O_2942,N_28560,N_28545);
and UO_2943 (O_2943,N_26367,N_29138);
and UO_2944 (O_2944,N_29915,N_25276);
nand UO_2945 (O_2945,N_29100,N_26818);
and UO_2946 (O_2946,N_25662,N_29483);
and UO_2947 (O_2947,N_28065,N_29077);
nand UO_2948 (O_2948,N_25967,N_25380);
nor UO_2949 (O_2949,N_26862,N_25803);
xor UO_2950 (O_2950,N_29615,N_28427);
nor UO_2951 (O_2951,N_27223,N_25212);
xor UO_2952 (O_2952,N_29604,N_25604);
xnor UO_2953 (O_2953,N_26796,N_28135);
nand UO_2954 (O_2954,N_28279,N_25838);
nand UO_2955 (O_2955,N_27711,N_28633);
and UO_2956 (O_2956,N_28229,N_27991);
nand UO_2957 (O_2957,N_26033,N_28146);
nand UO_2958 (O_2958,N_25963,N_26269);
and UO_2959 (O_2959,N_26127,N_27653);
nor UO_2960 (O_2960,N_26265,N_28503);
or UO_2961 (O_2961,N_26579,N_26573);
nand UO_2962 (O_2962,N_29855,N_29227);
nor UO_2963 (O_2963,N_25697,N_25515);
nor UO_2964 (O_2964,N_25317,N_26042);
and UO_2965 (O_2965,N_28538,N_25144);
xnor UO_2966 (O_2966,N_25332,N_29566);
nor UO_2967 (O_2967,N_25464,N_29093);
xnor UO_2968 (O_2968,N_28069,N_27936);
xnor UO_2969 (O_2969,N_27805,N_25092);
or UO_2970 (O_2970,N_26242,N_29163);
or UO_2971 (O_2971,N_28306,N_29804);
nand UO_2972 (O_2972,N_27796,N_27433);
nand UO_2973 (O_2973,N_25429,N_26224);
nand UO_2974 (O_2974,N_26356,N_28095);
nor UO_2975 (O_2975,N_26631,N_28460);
nor UO_2976 (O_2976,N_28838,N_29841);
and UO_2977 (O_2977,N_27108,N_29764);
or UO_2978 (O_2978,N_29082,N_28064);
or UO_2979 (O_2979,N_27059,N_29120);
nand UO_2980 (O_2980,N_27122,N_26260);
or UO_2981 (O_2981,N_28962,N_26335);
and UO_2982 (O_2982,N_26867,N_25052);
nor UO_2983 (O_2983,N_27538,N_28856);
or UO_2984 (O_2984,N_27459,N_28163);
xor UO_2985 (O_2985,N_27488,N_27520);
and UO_2986 (O_2986,N_29694,N_29608);
xnor UO_2987 (O_2987,N_26980,N_27658);
or UO_2988 (O_2988,N_26826,N_26148);
xnor UO_2989 (O_2989,N_27721,N_28589);
nor UO_2990 (O_2990,N_26173,N_25477);
xor UO_2991 (O_2991,N_25381,N_25726);
or UO_2992 (O_2992,N_26322,N_25686);
xor UO_2993 (O_2993,N_29883,N_25082);
or UO_2994 (O_2994,N_28495,N_25486);
or UO_2995 (O_2995,N_26902,N_26712);
nand UO_2996 (O_2996,N_25788,N_25633);
xnor UO_2997 (O_2997,N_27781,N_27818);
nor UO_2998 (O_2998,N_27835,N_25849);
or UO_2999 (O_2999,N_27345,N_25398);
or UO_3000 (O_3000,N_25802,N_29498);
and UO_3001 (O_3001,N_28595,N_28092);
or UO_3002 (O_3002,N_26226,N_27429);
nand UO_3003 (O_3003,N_28201,N_26648);
nor UO_3004 (O_3004,N_26737,N_28346);
nor UO_3005 (O_3005,N_25517,N_27269);
and UO_3006 (O_3006,N_28523,N_28672);
and UO_3007 (O_3007,N_25086,N_25298);
xnor UO_3008 (O_3008,N_29330,N_28199);
nand UO_3009 (O_3009,N_25501,N_26000);
nand UO_3010 (O_3010,N_27245,N_29977);
or UO_3011 (O_3011,N_25562,N_27989);
nor UO_3012 (O_3012,N_25429,N_27529);
and UO_3013 (O_3013,N_28725,N_29174);
or UO_3014 (O_3014,N_28858,N_28723);
xnor UO_3015 (O_3015,N_27006,N_27579);
nand UO_3016 (O_3016,N_28443,N_28631);
nand UO_3017 (O_3017,N_29810,N_29917);
and UO_3018 (O_3018,N_25786,N_25658);
and UO_3019 (O_3019,N_28940,N_28380);
xor UO_3020 (O_3020,N_27205,N_28647);
and UO_3021 (O_3021,N_26427,N_28080);
nand UO_3022 (O_3022,N_26448,N_28380);
nor UO_3023 (O_3023,N_28208,N_29703);
nand UO_3024 (O_3024,N_29499,N_28997);
nor UO_3025 (O_3025,N_26908,N_28528);
nand UO_3026 (O_3026,N_26268,N_26683);
and UO_3027 (O_3027,N_26859,N_28661);
nor UO_3028 (O_3028,N_28568,N_27323);
and UO_3029 (O_3029,N_29783,N_28981);
xor UO_3030 (O_3030,N_27946,N_28838);
nor UO_3031 (O_3031,N_25016,N_25582);
or UO_3032 (O_3032,N_27204,N_29740);
xor UO_3033 (O_3033,N_29309,N_27478);
xor UO_3034 (O_3034,N_27865,N_29727);
nor UO_3035 (O_3035,N_27335,N_29448);
xor UO_3036 (O_3036,N_25746,N_26516);
nor UO_3037 (O_3037,N_28899,N_29379);
and UO_3038 (O_3038,N_26727,N_26502);
xor UO_3039 (O_3039,N_29768,N_26907);
or UO_3040 (O_3040,N_26165,N_28662);
or UO_3041 (O_3041,N_26135,N_25372);
and UO_3042 (O_3042,N_25054,N_27230);
nor UO_3043 (O_3043,N_28403,N_26601);
nor UO_3044 (O_3044,N_29079,N_25882);
xnor UO_3045 (O_3045,N_26401,N_26072);
xnor UO_3046 (O_3046,N_27682,N_27373);
nor UO_3047 (O_3047,N_26554,N_25232);
nor UO_3048 (O_3048,N_29843,N_28624);
and UO_3049 (O_3049,N_29315,N_29476);
or UO_3050 (O_3050,N_26813,N_27109);
nor UO_3051 (O_3051,N_27362,N_27806);
xnor UO_3052 (O_3052,N_29378,N_25836);
and UO_3053 (O_3053,N_28140,N_25015);
xor UO_3054 (O_3054,N_27843,N_29272);
or UO_3055 (O_3055,N_26138,N_26177);
xnor UO_3056 (O_3056,N_26199,N_29334);
or UO_3057 (O_3057,N_28426,N_25638);
nand UO_3058 (O_3058,N_27982,N_25323);
nor UO_3059 (O_3059,N_27139,N_25542);
and UO_3060 (O_3060,N_29724,N_28399);
nor UO_3061 (O_3061,N_29517,N_28241);
and UO_3062 (O_3062,N_25113,N_25728);
nand UO_3063 (O_3063,N_28636,N_26841);
xor UO_3064 (O_3064,N_26050,N_26874);
or UO_3065 (O_3065,N_26593,N_25135);
nand UO_3066 (O_3066,N_29371,N_29327);
nand UO_3067 (O_3067,N_28414,N_28957);
and UO_3068 (O_3068,N_27194,N_26077);
or UO_3069 (O_3069,N_26428,N_29490);
and UO_3070 (O_3070,N_28251,N_26618);
xnor UO_3071 (O_3071,N_25751,N_26606);
xnor UO_3072 (O_3072,N_25130,N_28650);
and UO_3073 (O_3073,N_29878,N_27369);
and UO_3074 (O_3074,N_28709,N_27750);
nand UO_3075 (O_3075,N_28738,N_26324);
nand UO_3076 (O_3076,N_25213,N_28456);
nor UO_3077 (O_3077,N_29947,N_26914);
nor UO_3078 (O_3078,N_28933,N_25733);
or UO_3079 (O_3079,N_28308,N_27158);
nor UO_3080 (O_3080,N_28538,N_25884);
nor UO_3081 (O_3081,N_26417,N_25705);
xnor UO_3082 (O_3082,N_27401,N_29363);
or UO_3083 (O_3083,N_28360,N_26433);
xnor UO_3084 (O_3084,N_29854,N_28054);
nand UO_3085 (O_3085,N_26247,N_29134);
or UO_3086 (O_3086,N_27148,N_27600);
or UO_3087 (O_3087,N_27167,N_27444);
or UO_3088 (O_3088,N_27407,N_29093);
nand UO_3089 (O_3089,N_28384,N_28507);
xnor UO_3090 (O_3090,N_28901,N_28233);
and UO_3091 (O_3091,N_29856,N_28116);
and UO_3092 (O_3092,N_25692,N_29473);
and UO_3093 (O_3093,N_28856,N_29870);
xor UO_3094 (O_3094,N_26806,N_28049);
and UO_3095 (O_3095,N_27903,N_29736);
nor UO_3096 (O_3096,N_26587,N_27317);
xor UO_3097 (O_3097,N_29563,N_26427);
or UO_3098 (O_3098,N_26757,N_25587);
xor UO_3099 (O_3099,N_27492,N_26151);
xor UO_3100 (O_3100,N_26355,N_26231);
xor UO_3101 (O_3101,N_27997,N_27726);
and UO_3102 (O_3102,N_27816,N_29679);
or UO_3103 (O_3103,N_26924,N_25078);
and UO_3104 (O_3104,N_29759,N_26701);
or UO_3105 (O_3105,N_28339,N_25172);
or UO_3106 (O_3106,N_25357,N_28912);
and UO_3107 (O_3107,N_26935,N_25823);
xnor UO_3108 (O_3108,N_27082,N_27658);
nor UO_3109 (O_3109,N_28899,N_29222);
xor UO_3110 (O_3110,N_28656,N_26508);
xnor UO_3111 (O_3111,N_26789,N_26418);
xnor UO_3112 (O_3112,N_28698,N_25400);
xnor UO_3113 (O_3113,N_25757,N_25470);
nor UO_3114 (O_3114,N_26155,N_29692);
or UO_3115 (O_3115,N_26673,N_28399);
nand UO_3116 (O_3116,N_26841,N_25695);
nand UO_3117 (O_3117,N_25681,N_28445);
or UO_3118 (O_3118,N_26252,N_25344);
and UO_3119 (O_3119,N_26637,N_29002);
xor UO_3120 (O_3120,N_27303,N_25513);
and UO_3121 (O_3121,N_29224,N_25481);
nor UO_3122 (O_3122,N_25440,N_29651);
xor UO_3123 (O_3123,N_26048,N_27930);
xor UO_3124 (O_3124,N_29117,N_26228);
and UO_3125 (O_3125,N_29157,N_29212);
and UO_3126 (O_3126,N_25848,N_26546);
or UO_3127 (O_3127,N_27168,N_25999);
and UO_3128 (O_3128,N_29233,N_26093);
or UO_3129 (O_3129,N_25072,N_27432);
and UO_3130 (O_3130,N_26418,N_25642);
and UO_3131 (O_3131,N_28041,N_27395);
and UO_3132 (O_3132,N_28160,N_29525);
nor UO_3133 (O_3133,N_28821,N_26835);
nor UO_3134 (O_3134,N_26088,N_28329);
or UO_3135 (O_3135,N_25616,N_27412);
or UO_3136 (O_3136,N_27795,N_26362);
and UO_3137 (O_3137,N_28593,N_26195);
xnor UO_3138 (O_3138,N_25238,N_28950);
nor UO_3139 (O_3139,N_26538,N_26788);
and UO_3140 (O_3140,N_29806,N_25870);
nor UO_3141 (O_3141,N_25154,N_26455);
and UO_3142 (O_3142,N_26027,N_27415);
nor UO_3143 (O_3143,N_26646,N_28053);
or UO_3144 (O_3144,N_25002,N_25220);
nand UO_3145 (O_3145,N_26168,N_29283);
nor UO_3146 (O_3146,N_27594,N_26865);
or UO_3147 (O_3147,N_28246,N_25793);
nand UO_3148 (O_3148,N_27169,N_27451);
xor UO_3149 (O_3149,N_27003,N_25755);
nand UO_3150 (O_3150,N_27763,N_29330);
nor UO_3151 (O_3151,N_26326,N_28300);
or UO_3152 (O_3152,N_25988,N_28297);
or UO_3153 (O_3153,N_29723,N_25275);
xnor UO_3154 (O_3154,N_25709,N_28323);
nor UO_3155 (O_3155,N_26884,N_25874);
nor UO_3156 (O_3156,N_29570,N_28544);
xor UO_3157 (O_3157,N_27001,N_27053);
nor UO_3158 (O_3158,N_28645,N_25559);
or UO_3159 (O_3159,N_25671,N_25387);
or UO_3160 (O_3160,N_29048,N_26609);
nand UO_3161 (O_3161,N_29188,N_28563);
nand UO_3162 (O_3162,N_26608,N_28679);
nand UO_3163 (O_3163,N_25524,N_27382);
and UO_3164 (O_3164,N_25506,N_25944);
or UO_3165 (O_3165,N_25712,N_29852);
nand UO_3166 (O_3166,N_29891,N_25244);
or UO_3167 (O_3167,N_27036,N_29458);
nor UO_3168 (O_3168,N_26983,N_29893);
nor UO_3169 (O_3169,N_29851,N_28385);
nand UO_3170 (O_3170,N_26109,N_27785);
or UO_3171 (O_3171,N_27401,N_28389);
nand UO_3172 (O_3172,N_26303,N_25858);
and UO_3173 (O_3173,N_29036,N_26688);
and UO_3174 (O_3174,N_27426,N_26277);
and UO_3175 (O_3175,N_28698,N_25295);
nor UO_3176 (O_3176,N_27141,N_29918);
xnor UO_3177 (O_3177,N_29444,N_26563);
and UO_3178 (O_3178,N_28083,N_25179);
xor UO_3179 (O_3179,N_27254,N_28289);
and UO_3180 (O_3180,N_26613,N_27491);
xor UO_3181 (O_3181,N_26087,N_25372);
nand UO_3182 (O_3182,N_29767,N_27510);
nor UO_3183 (O_3183,N_26647,N_25403);
and UO_3184 (O_3184,N_25980,N_28555);
nand UO_3185 (O_3185,N_27757,N_29302);
or UO_3186 (O_3186,N_26272,N_29904);
xnor UO_3187 (O_3187,N_26146,N_28227);
nand UO_3188 (O_3188,N_27190,N_27049);
nor UO_3189 (O_3189,N_29075,N_25195);
or UO_3190 (O_3190,N_28032,N_27086);
nand UO_3191 (O_3191,N_25221,N_28794);
nand UO_3192 (O_3192,N_26795,N_29794);
nand UO_3193 (O_3193,N_26332,N_27731);
nor UO_3194 (O_3194,N_28864,N_27852);
and UO_3195 (O_3195,N_26240,N_28460);
or UO_3196 (O_3196,N_29585,N_26876);
xnor UO_3197 (O_3197,N_27661,N_27447);
or UO_3198 (O_3198,N_28306,N_25101);
and UO_3199 (O_3199,N_26486,N_28682);
xor UO_3200 (O_3200,N_28224,N_28178);
or UO_3201 (O_3201,N_28581,N_25876);
xnor UO_3202 (O_3202,N_27112,N_27170);
xor UO_3203 (O_3203,N_26404,N_29106);
nor UO_3204 (O_3204,N_28305,N_29823);
xor UO_3205 (O_3205,N_28287,N_27904);
or UO_3206 (O_3206,N_29716,N_27517);
and UO_3207 (O_3207,N_26181,N_26433);
nor UO_3208 (O_3208,N_27642,N_26541);
and UO_3209 (O_3209,N_25366,N_28335);
and UO_3210 (O_3210,N_29908,N_28532);
xnor UO_3211 (O_3211,N_26226,N_26873);
nor UO_3212 (O_3212,N_27873,N_27938);
or UO_3213 (O_3213,N_29156,N_29111);
nor UO_3214 (O_3214,N_28639,N_28747);
xnor UO_3215 (O_3215,N_27921,N_26818);
nor UO_3216 (O_3216,N_25103,N_29875);
nand UO_3217 (O_3217,N_29250,N_28285);
nor UO_3218 (O_3218,N_29745,N_28004);
xnor UO_3219 (O_3219,N_27471,N_27587);
nor UO_3220 (O_3220,N_27926,N_28429);
and UO_3221 (O_3221,N_27557,N_28636);
xnor UO_3222 (O_3222,N_28183,N_28367);
nor UO_3223 (O_3223,N_26516,N_28079);
nand UO_3224 (O_3224,N_27980,N_29730);
or UO_3225 (O_3225,N_26267,N_29929);
and UO_3226 (O_3226,N_26726,N_26814);
and UO_3227 (O_3227,N_29263,N_29507);
nand UO_3228 (O_3228,N_29595,N_29123);
or UO_3229 (O_3229,N_26599,N_25821);
nand UO_3230 (O_3230,N_29901,N_27038);
xor UO_3231 (O_3231,N_25314,N_28983);
and UO_3232 (O_3232,N_27162,N_28691);
nand UO_3233 (O_3233,N_25423,N_28414);
and UO_3234 (O_3234,N_27148,N_25142);
and UO_3235 (O_3235,N_28612,N_25220);
or UO_3236 (O_3236,N_28605,N_29871);
nand UO_3237 (O_3237,N_26088,N_25077);
nor UO_3238 (O_3238,N_29743,N_29201);
xor UO_3239 (O_3239,N_26474,N_28685);
nor UO_3240 (O_3240,N_25266,N_27074);
nand UO_3241 (O_3241,N_27167,N_28615);
and UO_3242 (O_3242,N_29384,N_26780);
nand UO_3243 (O_3243,N_27309,N_26779);
nor UO_3244 (O_3244,N_27395,N_28346);
xnor UO_3245 (O_3245,N_29782,N_28125);
nand UO_3246 (O_3246,N_26271,N_26429);
xor UO_3247 (O_3247,N_26453,N_29775);
nand UO_3248 (O_3248,N_27666,N_26195);
xor UO_3249 (O_3249,N_25903,N_29850);
and UO_3250 (O_3250,N_27880,N_29047);
and UO_3251 (O_3251,N_25322,N_25452);
nand UO_3252 (O_3252,N_26096,N_27695);
nor UO_3253 (O_3253,N_25129,N_28661);
nor UO_3254 (O_3254,N_26089,N_25921);
xnor UO_3255 (O_3255,N_29661,N_27792);
nor UO_3256 (O_3256,N_27178,N_28865);
and UO_3257 (O_3257,N_27200,N_27902);
xnor UO_3258 (O_3258,N_28075,N_25249);
and UO_3259 (O_3259,N_25152,N_26399);
or UO_3260 (O_3260,N_28510,N_27870);
nand UO_3261 (O_3261,N_27452,N_27509);
and UO_3262 (O_3262,N_27945,N_26124);
nand UO_3263 (O_3263,N_29458,N_29408);
nor UO_3264 (O_3264,N_26651,N_28720);
nand UO_3265 (O_3265,N_29885,N_27355);
xnor UO_3266 (O_3266,N_27754,N_28096);
xnor UO_3267 (O_3267,N_29171,N_29091);
xnor UO_3268 (O_3268,N_29349,N_29744);
nand UO_3269 (O_3269,N_27945,N_26801);
nor UO_3270 (O_3270,N_29881,N_25822);
and UO_3271 (O_3271,N_28704,N_25146);
nand UO_3272 (O_3272,N_27413,N_25356);
nor UO_3273 (O_3273,N_27531,N_28835);
and UO_3274 (O_3274,N_26666,N_25849);
and UO_3275 (O_3275,N_28166,N_27536);
and UO_3276 (O_3276,N_28526,N_27191);
nand UO_3277 (O_3277,N_25090,N_26875);
and UO_3278 (O_3278,N_26747,N_25122);
xor UO_3279 (O_3279,N_29111,N_26868);
xor UO_3280 (O_3280,N_29859,N_25815);
nor UO_3281 (O_3281,N_25941,N_25001);
nor UO_3282 (O_3282,N_26674,N_28666);
or UO_3283 (O_3283,N_26860,N_27884);
and UO_3284 (O_3284,N_29262,N_27923);
nor UO_3285 (O_3285,N_27067,N_27946);
xnor UO_3286 (O_3286,N_27036,N_27520);
xor UO_3287 (O_3287,N_26707,N_27433);
xnor UO_3288 (O_3288,N_29493,N_27564);
nor UO_3289 (O_3289,N_26496,N_27823);
nand UO_3290 (O_3290,N_27608,N_27915);
or UO_3291 (O_3291,N_25382,N_27012);
nor UO_3292 (O_3292,N_27144,N_28430);
nor UO_3293 (O_3293,N_27759,N_29790);
nand UO_3294 (O_3294,N_29373,N_26594);
nand UO_3295 (O_3295,N_29216,N_29202);
nand UO_3296 (O_3296,N_26063,N_27205);
or UO_3297 (O_3297,N_26788,N_28440);
or UO_3298 (O_3298,N_27022,N_25857);
or UO_3299 (O_3299,N_26504,N_27827);
or UO_3300 (O_3300,N_25201,N_25564);
or UO_3301 (O_3301,N_28848,N_25065);
nor UO_3302 (O_3302,N_25095,N_29747);
nand UO_3303 (O_3303,N_28440,N_28026);
nor UO_3304 (O_3304,N_29528,N_28900);
nand UO_3305 (O_3305,N_25810,N_28820);
or UO_3306 (O_3306,N_26805,N_26885);
xor UO_3307 (O_3307,N_26396,N_29741);
nor UO_3308 (O_3308,N_26324,N_27647);
nand UO_3309 (O_3309,N_25449,N_28699);
nand UO_3310 (O_3310,N_26082,N_25074);
nand UO_3311 (O_3311,N_26927,N_29789);
and UO_3312 (O_3312,N_27090,N_29076);
nand UO_3313 (O_3313,N_29332,N_29293);
nand UO_3314 (O_3314,N_25189,N_26077);
xnor UO_3315 (O_3315,N_27303,N_26450);
xor UO_3316 (O_3316,N_29619,N_28465);
xor UO_3317 (O_3317,N_26596,N_29442);
nand UO_3318 (O_3318,N_25499,N_29587);
nor UO_3319 (O_3319,N_27430,N_29039);
or UO_3320 (O_3320,N_25743,N_25005);
or UO_3321 (O_3321,N_25318,N_25032);
nand UO_3322 (O_3322,N_28474,N_28681);
xnor UO_3323 (O_3323,N_26403,N_26897);
nand UO_3324 (O_3324,N_29213,N_29018);
nor UO_3325 (O_3325,N_28967,N_25900);
nand UO_3326 (O_3326,N_29625,N_26418);
and UO_3327 (O_3327,N_26417,N_28733);
nor UO_3328 (O_3328,N_28167,N_25015);
and UO_3329 (O_3329,N_27665,N_26940);
and UO_3330 (O_3330,N_25476,N_27890);
nand UO_3331 (O_3331,N_29642,N_28320);
nand UO_3332 (O_3332,N_26263,N_27724);
and UO_3333 (O_3333,N_29450,N_27063);
nand UO_3334 (O_3334,N_29256,N_25507);
nor UO_3335 (O_3335,N_28293,N_28096);
nor UO_3336 (O_3336,N_29226,N_28814);
xnor UO_3337 (O_3337,N_28885,N_27780);
nor UO_3338 (O_3338,N_28073,N_27050);
or UO_3339 (O_3339,N_27192,N_26151);
nor UO_3340 (O_3340,N_28447,N_28262);
xnor UO_3341 (O_3341,N_25711,N_25091);
xnor UO_3342 (O_3342,N_27087,N_29841);
and UO_3343 (O_3343,N_29804,N_28461);
xnor UO_3344 (O_3344,N_26579,N_28834);
nand UO_3345 (O_3345,N_28570,N_29392);
xnor UO_3346 (O_3346,N_29832,N_26065);
nor UO_3347 (O_3347,N_29722,N_26623);
xor UO_3348 (O_3348,N_27916,N_26419);
xor UO_3349 (O_3349,N_26584,N_27327);
xor UO_3350 (O_3350,N_27105,N_26495);
xor UO_3351 (O_3351,N_28026,N_26803);
or UO_3352 (O_3352,N_29353,N_25434);
xnor UO_3353 (O_3353,N_25226,N_25234);
nor UO_3354 (O_3354,N_27821,N_29038);
or UO_3355 (O_3355,N_27050,N_25889);
nor UO_3356 (O_3356,N_25589,N_28335);
and UO_3357 (O_3357,N_25545,N_27211);
and UO_3358 (O_3358,N_27678,N_28635);
nand UO_3359 (O_3359,N_28142,N_29102);
nor UO_3360 (O_3360,N_26135,N_25742);
and UO_3361 (O_3361,N_27816,N_29425);
or UO_3362 (O_3362,N_27710,N_25518);
xor UO_3363 (O_3363,N_26014,N_26936);
or UO_3364 (O_3364,N_25628,N_28770);
or UO_3365 (O_3365,N_29540,N_29074);
xnor UO_3366 (O_3366,N_28260,N_27786);
nand UO_3367 (O_3367,N_28078,N_28638);
or UO_3368 (O_3368,N_27007,N_28107);
xnor UO_3369 (O_3369,N_26684,N_28444);
nand UO_3370 (O_3370,N_27435,N_27814);
or UO_3371 (O_3371,N_25360,N_25557);
xor UO_3372 (O_3372,N_25955,N_25458);
nand UO_3373 (O_3373,N_28517,N_27819);
nor UO_3374 (O_3374,N_27625,N_27162);
nor UO_3375 (O_3375,N_29353,N_29440);
nand UO_3376 (O_3376,N_27066,N_25947);
nor UO_3377 (O_3377,N_26159,N_26403);
nor UO_3378 (O_3378,N_27802,N_26693);
xor UO_3379 (O_3379,N_28784,N_25620);
xnor UO_3380 (O_3380,N_29407,N_25634);
xnor UO_3381 (O_3381,N_27669,N_29719);
and UO_3382 (O_3382,N_26728,N_28243);
and UO_3383 (O_3383,N_29571,N_25174);
nor UO_3384 (O_3384,N_27788,N_26449);
nor UO_3385 (O_3385,N_26737,N_27759);
or UO_3386 (O_3386,N_25766,N_26518);
or UO_3387 (O_3387,N_27077,N_25841);
nand UO_3388 (O_3388,N_27501,N_27697);
nand UO_3389 (O_3389,N_27980,N_29594);
and UO_3390 (O_3390,N_28346,N_29257);
xor UO_3391 (O_3391,N_28852,N_27277);
and UO_3392 (O_3392,N_26524,N_26392);
or UO_3393 (O_3393,N_26173,N_27192);
nor UO_3394 (O_3394,N_28010,N_29384);
and UO_3395 (O_3395,N_26868,N_28225);
or UO_3396 (O_3396,N_26597,N_28002);
nand UO_3397 (O_3397,N_26711,N_28502);
xor UO_3398 (O_3398,N_28233,N_28401);
nor UO_3399 (O_3399,N_27247,N_28447);
nand UO_3400 (O_3400,N_26752,N_27744);
or UO_3401 (O_3401,N_28260,N_25725);
xor UO_3402 (O_3402,N_28201,N_28148);
nor UO_3403 (O_3403,N_27673,N_25319);
and UO_3404 (O_3404,N_29447,N_27134);
or UO_3405 (O_3405,N_27993,N_28991);
xnor UO_3406 (O_3406,N_29036,N_26005);
nand UO_3407 (O_3407,N_28443,N_27031);
or UO_3408 (O_3408,N_26098,N_25115);
nor UO_3409 (O_3409,N_29625,N_29966);
nor UO_3410 (O_3410,N_26783,N_26966);
or UO_3411 (O_3411,N_29060,N_25799);
nand UO_3412 (O_3412,N_26086,N_28905);
nor UO_3413 (O_3413,N_28710,N_25607);
or UO_3414 (O_3414,N_29107,N_29670);
and UO_3415 (O_3415,N_29125,N_26667);
xnor UO_3416 (O_3416,N_27339,N_29837);
nand UO_3417 (O_3417,N_25101,N_25799);
or UO_3418 (O_3418,N_29660,N_29715);
xor UO_3419 (O_3419,N_27422,N_28454);
or UO_3420 (O_3420,N_29296,N_28930);
nand UO_3421 (O_3421,N_26737,N_25863);
xor UO_3422 (O_3422,N_28350,N_25445);
xnor UO_3423 (O_3423,N_29998,N_25212);
and UO_3424 (O_3424,N_26230,N_27640);
xnor UO_3425 (O_3425,N_27742,N_28574);
nor UO_3426 (O_3426,N_27818,N_26572);
nand UO_3427 (O_3427,N_27326,N_28840);
nor UO_3428 (O_3428,N_26908,N_25224);
xor UO_3429 (O_3429,N_28469,N_27112);
nand UO_3430 (O_3430,N_25093,N_26189);
or UO_3431 (O_3431,N_29622,N_25289);
nand UO_3432 (O_3432,N_27532,N_25439);
xnor UO_3433 (O_3433,N_28227,N_29691);
xor UO_3434 (O_3434,N_29866,N_29907);
nor UO_3435 (O_3435,N_27807,N_29240);
nor UO_3436 (O_3436,N_25555,N_26341);
xor UO_3437 (O_3437,N_29855,N_27674);
and UO_3438 (O_3438,N_28085,N_29694);
nand UO_3439 (O_3439,N_29117,N_25194);
nor UO_3440 (O_3440,N_29627,N_28784);
xor UO_3441 (O_3441,N_28727,N_27285);
nand UO_3442 (O_3442,N_27107,N_25915);
nand UO_3443 (O_3443,N_27702,N_26454);
nand UO_3444 (O_3444,N_26724,N_26026);
nand UO_3445 (O_3445,N_27394,N_28002);
xnor UO_3446 (O_3446,N_25244,N_26713);
or UO_3447 (O_3447,N_26435,N_28827);
xnor UO_3448 (O_3448,N_27881,N_27481);
nand UO_3449 (O_3449,N_28597,N_25926);
xor UO_3450 (O_3450,N_26485,N_29640);
or UO_3451 (O_3451,N_29588,N_25473);
nor UO_3452 (O_3452,N_26381,N_25442);
and UO_3453 (O_3453,N_29414,N_25021);
and UO_3454 (O_3454,N_26731,N_25160);
xor UO_3455 (O_3455,N_28369,N_28072);
xor UO_3456 (O_3456,N_29249,N_28423);
or UO_3457 (O_3457,N_27228,N_28590);
and UO_3458 (O_3458,N_27747,N_27886);
nand UO_3459 (O_3459,N_27087,N_29110);
nor UO_3460 (O_3460,N_25603,N_25591);
or UO_3461 (O_3461,N_26828,N_27173);
nor UO_3462 (O_3462,N_25937,N_28963);
and UO_3463 (O_3463,N_25225,N_27895);
nor UO_3464 (O_3464,N_25077,N_29588);
nand UO_3465 (O_3465,N_29865,N_29717);
nand UO_3466 (O_3466,N_29521,N_26088);
or UO_3467 (O_3467,N_27428,N_29831);
nand UO_3468 (O_3468,N_25590,N_27112);
nand UO_3469 (O_3469,N_29306,N_27478);
or UO_3470 (O_3470,N_28154,N_29894);
xnor UO_3471 (O_3471,N_29511,N_27853);
and UO_3472 (O_3472,N_28094,N_26914);
nor UO_3473 (O_3473,N_26787,N_28571);
nand UO_3474 (O_3474,N_27103,N_29477);
or UO_3475 (O_3475,N_26931,N_26777);
and UO_3476 (O_3476,N_29695,N_26487);
nor UO_3477 (O_3477,N_29297,N_29235);
xor UO_3478 (O_3478,N_29854,N_29561);
nor UO_3479 (O_3479,N_27207,N_26152);
xor UO_3480 (O_3480,N_27061,N_26464);
nand UO_3481 (O_3481,N_26385,N_28323);
and UO_3482 (O_3482,N_27876,N_26235);
xor UO_3483 (O_3483,N_27915,N_28872);
or UO_3484 (O_3484,N_29810,N_29139);
or UO_3485 (O_3485,N_28214,N_25038);
and UO_3486 (O_3486,N_25496,N_26885);
nor UO_3487 (O_3487,N_25883,N_29503);
nor UO_3488 (O_3488,N_27656,N_28331);
nand UO_3489 (O_3489,N_26499,N_29862);
nand UO_3490 (O_3490,N_26340,N_27123);
or UO_3491 (O_3491,N_26310,N_28831);
and UO_3492 (O_3492,N_27922,N_27490);
xor UO_3493 (O_3493,N_29810,N_28141);
xor UO_3494 (O_3494,N_28707,N_27892);
or UO_3495 (O_3495,N_29498,N_28507);
or UO_3496 (O_3496,N_28651,N_26455);
nor UO_3497 (O_3497,N_29464,N_29156);
or UO_3498 (O_3498,N_27958,N_25331);
or UO_3499 (O_3499,N_28213,N_29760);
endmodule